module dtc_split05_bm61 (
	input  wire [12-1:0] inp,
	output wire [11-1:0] outp
);

	wire [11-1:0] node1;
	wire [11-1:0] node2;
	wire [11-1:0] node3;
	wire [11-1:0] node4;
	wire [11-1:0] node5;
	wire [11-1:0] node8;
	wire [11-1:0] node9;
	wire [11-1:0] node10;
	wire [11-1:0] node14;
	wire [11-1:0] node15;
	wire [11-1:0] node19;
	wire [11-1:0] node20;
	wire [11-1:0] node22;
	wire [11-1:0] node23;
	wire [11-1:0] node27;
	wire [11-1:0] node29;
	wire [11-1:0] node30;
	wire [11-1:0] node33;
	wire [11-1:0] node36;
	wire [11-1:0] node37;
	wire [11-1:0] node38;
	wire [11-1:0] node39;
	wire [11-1:0] node40;
	wire [11-1:0] node43;
	wire [11-1:0] node46;
	wire [11-1:0] node48;
	wire [11-1:0] node51;
	wire [11-1:0] node52;
	wire [11-1:0] node55;
	wire [11-1:0] node58;
	wire [11-1:0] node59;
	wire [11-1:0] node60;
	wire [11-1:0] node63;
	wire [11-1:0] node64;
	wire [11-1:0] node68;
	wire [11-1:0] node69;
	wire [11-1:0] node70;
	wire [11-1:0] node73;
	wire [11-1:0] node76;
	wire [11-1:0] node77;
	wire [11-1:0] node80;
	wire [11-1:0] node83;
	wire [11-1:0] node84;
	wire [11-1:0] node85;
	wire [11-1:0] node86;
	wire [11-1:0] node87;
	wire [11-1:0] node89;
	wire [11-1:0] node93;
	wire [11-1:0] node94;
	wire [11-1:0] node95;
	wire [11-1:0] node98;
	wire [11-1:0] node101;
	wire [11-1:0] node102;
	wire [11-1:0] node106;
	wire [11-1:0] node107;
	wire [11-1:0] node108;
	wire [11-1:0] node109;
	wire [11-1:0] node112;
	wire [11-1:0] node115;
	wire [11-1:0] node116;
	wire [11-1:0] node120;
	wire [11-1:0] node121;
	wire [11-1:0] node122;
	wire [11-1:0] node125;
	wire [11-1:0] node128;
	wire [11-1:0] node129;
	wire [11-1:0] node133;
	wire [11-1:0] node134;
	wire [11-1:0] node135;
	wire [11-1:0] node136;
	wire [11-1:0] node137;
	wire [11-1:0] node141;
	wire [11-1:0] node142;
	wire [11-1:0] node146;
	wire [11-1:0] node147;
	wire [11-1:0] node148;
	wire [11-1:0] node151;
	wire [11-1:0] node154;
	wire [11-1:0] node155;
	wire [11-1:0] node159;
	wire [11-1:0] node160;
	wire [11-1:0] node161;
	wire [11-1:0] node165;
	wire [11-1:0] node166;
	wire [11-1:0] node168;
	wire [11-1:0] node171;
	wire [11-1:0] node172;
	wire [11-1:0] node176;
	wire [11-1:0] node177;
	wire [11-1:0] node178;
	wire [11-1:0] node179;
	wire [11-1:0] node180;
	wire [11-1:0] node181;
	wire [11-1:0] node182;
	wire [11-1:0] node186;
	wire [11-1:0] node187;
	wire [11-1:0] node191;
	wire [11-1:0] node192;
	wire [11-1:0] node196;
	wire [11-1:0] node197;
	wire [11-1:0] node198;
	wire [11-1:0] node201;
	wire [11-1:0] node202;
	wire [11-1:0] node205;
	wire [11-1:0] node208;
	wire [11-1:0] node209;
	wire [11-1:0] node212;
	wire [11-1:0] node213;
	wire [11-1:0] node216;
	wire [11-1:0] node219;
	wire [11-1:0] node220;
	wire [11-1:0] node221;
	wire [11-1:0] node222;
	wire [11-1:0] node224;
	wire [11-1:0] node227;
	wire [11-1:0] node228;
	wire [11-1:0] node232;
	wire [11-1:0] node233;
	wire [11-1:0] node235;
	wire [11-1:0] node238;
	wire [11-1:0] node240;
	wire [11-1:0] node243;
	wire [11-1:0] node244;
	wire [11-1:0] node245;
	wire [11-1:0] node248;
	wire [11-1:0] node249;
	wire [11-1:0] node252;
	wire [11-1:0] node255;
	wire [11-1:0] node256;
	wire [11-1:0] node257;
	wire [11-1:0] node260;
	wire [11-1:0] node263;
	wire [11-1:0] node266;
	wire [11-1:0] node267;
	wire [11-1:0] node268;
	wire [11-1:0] node269;
	wire [11-1:0] node270;
	wire [11-1:0] node271;
	wire [11-1:0] node275;
	wire [11-1:0] node277;
	wire [11-1:0] node280;
	wire [11-1:0] node281;
	wire [11-1:0] node285;
	wire [11-1:0] node286;
	wire [11-1:0] node287;
	wire [11-1:0] node288;
	wire [11-1:0] node292;
	wire [11-1:0] node295;
	wire [11-1:0] node297;
	wire [11-1:0] node300;
	wire [11-1:0] node301;
	wire [11-1:0] node302;
	wire [11-1:0] node304;
	wire [11-1:0] node307;
	wire [11-1:0] node310;
	wire [11-1:0] node311;
	wire [11-1:0] node312;
	wire [11-1:0] node313;
	wire [11-1:0] node316;
	wire [11-1:0] node319;
	wire [11-1:0] node320;
	wire [11-1:0] node323;
	wire [11-1:0] node326;
	wire [11-1:0] node327;
	wire [11-1:0] node328;
	wire [11-1:0] node331;
	wire [11-1:0] node334;

	assign outp = (inp[1]) ? node176 : node1;
		assign node1 = (inp[7]) ? node83 : node2;
			assign node2 = (inp[2]) ? node36 : node3;
				assign node3 = (inp[6]) ? node19 : node4;
					assign node4 = (inp[5]) ? node8 : node5;
						assign node5 = (inp[3]) ? 11'b01101111101 : 11'b01101011101;
						assign node8 = (inp[8]) ? node14 : node9;
							assign node9 = (inp[10]) ? 11'b11010001110 : node10;
								assign node10 = (inp[9]) ? 11'b01011111010 : 11'b01011011110;
							assign node14 = (inp[3]) ? 11'b01101101100 : node15;
								assign node15 = (inp[0]) ? 11'b01001111010 : 11'b01001011010;
					assign node19 = (inp[10]) ? node27 : node20;
						assign node20 = (inp[3]) ? node22 : 11'b01011011001;
							assign node22 = (inp[4]) ? 11'b11101001001 : node23;
								assign node23 = (inp[5]) ? 11'b11000111001 : 11'b11101111000;
						assign node27 = (inp[3]) ? node29 : 11'b01101111111;
							assign node29 = (inp[5]) ? node33 : node30;
								assign node30 = (inp[0]) ? 11'b01000001010 : 11'b01110000010;
								assign node33 = (inp[11]) ? 11'b01001001001 : 11'b01010001011;
				assign node36 = (inp[0]) ? node58 : node37;
					assign node37 = (inp[6]) ? node51 : node38;
						assign node38 = (inp[11]) ? node46 : node39;
							assign node39 = (inp[10]) ? node43 : node40;
								assign node40 = (inp[8]) ? 11'b11101010101 : 11'b01111110100;
								assign node43 = (inp[3]) ? 11'b01000110001 : 11'b11011010000;
							assign node46 = (inp[8]) ? node48 : 11'b01100000011;
								assign node48 = (inp[4]) ? 11'b11010010101 : 11'b11010110001;
						assign node51 = (inp[10]) ? node55 : node52;
							assign node52 = (inp[8]) ? 11'b11100100111 : 11'b01100101100;
							assign node55 = (inp[4]) ? 11'b01011101010 : 11'b11110001011;
					assign node58 = (inp[8]) ? node68 : node59;
						assign node59 = (inp[5]) ? node63 : node60;
							assign node60 = (inp[3]) ? 11'b01001101000 : 11'b01001100011;
							assign node63 = (inp[9]) ? 11'b01000100011 : node64;
								assign node64 = (inp[6]) ? 11'b01111100001 : 11'b01110000001;
						assign node68 = (inp[11]) ? node76 : node69;
							assign node69 = (inp[10]) ? node73 : node70;
								assign node70 = (inp[5]) ? 11'b01100010010 : 11'b01010110001;
								assign node73 = (inp[3]) ? 11'b01111000011 : 11'b01101110011;
							assign node76 = (inp[9]) ? node80 : node77;
								assign node77 = (inp[4]) ? 11'b01100010010 : 11'b01100100000;
								assign node80 = (inp[3]) ? 11'b01000000000 : 11'b01000100000;
			assign node83 = (inp[6]) ? node133 : node84;
				assign node84 = (inp[2]) ? node106 : node85;
					assign node85 = (inp[4]) ? node93 : node86;
						assign node86 = (inp[9]) ? 11'b01000000111 : node87;
							assign node87 = (inp[10]) ? node89 : 11'b01001110010;
								assign node89 = (inp[8]) ? 11'b01001010100 : 11'b11011000001;
						assign node93 = (inp[11]) ? node101 : node94;
							assign node94 = (inp[3]) ? node98 : node95;
								assign node95 = (inp[9]) ? 11'b01101110100 : 11'b11110110100;
								assign node98 = (inp[9]) ? 11'b01110010010 : 11'b01110100000;
							assign node101 = (inp[8]) ? 11'b10101001111 : node102;
								assign node102 = (inp[10]) ? 11'b01100000000 : 11'b11110010110;
					assign node106 = (inp[8]) ? node120 : node107;
						assign node107 = (inp[11]) ? node115 : node108;
							assign node108 = (inp[4]) ? node112 : node109;
								assign node109 = (inp[10]) ? 11'b00101111110 : 11'b00111111000;
								assign node112 = (inp[10]) ? 11'b00010111000 : 11'b10001111010;
							assign node115 = (inp[4]) ? 11'b00000001100 : node116;
								assign node116 = (inp[10]) ? 11'b00111011110 : 11'b00011001010;
						assign node120 = (inp[3]) ? node128 : node121;
							assign node121 = (inp[9]) ? node125 : node122;
								assign node122 = (inp[0]) ? 11'b00001001101 : 11'b10001011101;
								assign node125 = (inp[4]) ? 11'b10010011001 : 11'b00110011001;
							assign node128 = (inp[5]) ? 11'b10100101000 : node129;
								assign node129 = (inp[9]) ? 11'b00101101011 : 11'b00000101001;
				assign node133 = (inp[8]) ? node159 : node134;
					assign node134 = (inp[2]) ? node146 : node135;
						assign node135 = (inp[5]) ? node141 : node136;
							assign node136 = (inp[9]) ? 11'b00101011000 : node137;
								assign node137 = (inp[0]) ? 11'b00011101000 : 11'b00011101010;
							assign node141 = (inp[0]) ? 11'b00011110011 : node142;
								assign node142 = (inp[9]) ? 11'b10001110101 : 11'b00000010001;
						assign node146 = (inp[4]) ? node154 : node147;
							assign node147 = (inp[0]) ? node151 : node148;
								assign node148 = (inp[5]) ? 11'b10000100011 : 11'b00101100011;
								assign node151 = (inp[11]) ? 11'b00011000011 : 11'b00110000001;
							assign node154 = (inp[9]) ? 11'b00001110001 : node155;
								assign node155 = (inp[5]) ? 11'b00110010111 : 11'b00010010011;
					assign node159 = (inp[9]) ? node165 : node160;
						assign node160 = (inp[3]) ? 11'b00111010110 : node161;
							assign node161 = (inp[2]) ? 11'b00111100100 : 11'b00001100000;
						assign node165 = (inp[0]) ? node171 : node166;
							assign node166 = (inp[5]) ? node168 : 11'b00100010111;
								assign node168 = (inp[10]) ? 11'b00000000000 : 11'b00000110110;
							assign node171 = (inp[4]) ? 11'b00011110100 : node172;
								assign node172 = (inp[2]) ? 11'b00000100010 : 11'b00011100010;
		assign node176 = (inp[7]) ? node266 : node177;
			assign node177 = (inp[6]) ? node219 : node178;
				assign node178 = (inp[8]) ? node196 : node179;
					assign node179 = (inp[11]) ? node191 : node180;
						assign node180 = (inp[2]) ? node186 : node181;
							assign node181 = (inp[5]) ? 11'b00111111101 : node182;
								assign node182 = (inp[4]) ? 11'b00001111001 : 11'b00000111001;
							assign node186 = (inp[9]) ? 11'b00100011001 : node187;
								assign node187 = (inp[3]) ? 11'b00011001000 : 11'b10111001010;
						assign node191 = (inp[3]) ? 11'b10010011001 : node192;
							assign node192 = (inp[10]) ? 11'b10000111111 : 11'b00010111011;
					assign node196 = (inp[4]) ? node208 : node197;
						assign node197 = (inp[10]) ? node201 : node198;
							assign node198 = (inp[3]) ? 11'b10000011010 : 11'b00100011010;
							assign node201 = (inp[11]) ? node205 : node202;
								assign node202 = (inp[2]) ? 11'b00000101100 : 11'b00001111000;
								assign node205 = (inp[9]) ? 11'b10001001110 : 11'b00011011110;
						assign node208 = (inp[2]) ? node212 : node209;
							assign node209 = (inp[5]) ? 11'b00111111100 : 11'b00100101100;
							assign node212 = (inp[5]) ? node216 : node213;
								assign node213 = (inp[10]) ? 11'b00110001001 : 11'b00011001100;
								assign node216 = (inp[3]) ? 11'b00001001000 : 11'b00000001100;
				assign node219 = (inp[3]) ? node243 : node220;
					assign node220 = (inp[2]) ? node232 : node221;
						assign node221 = (inp[0]) ? node227 : node222;
							assign node222 = (inp[4]) ? node224 : 11'b00011011010;
								assign node224 = (inp[10]) ? 11'b10000001110 : 11'b00000011110;
							assign node227 = (inp[5]) ? 11'b00111110001 : node228;
								assign node228 = (inp[4]) ? 11'b00001011010 : 11'b00110111100;
						assign node232 = (inp[5]) ? node238 : node233;
							assign node233 = (inp[0]) ? node235 : 11'b10001110100;
								assign node235 = (inp[10]) ? 11'b00110000100 : 11'b00100100100;
							assign node238 = (inp[8]) ? node240 : 11'b00000000000;
								assign node240 = (inp[11]) ? 11'b00010000110 : 11'b00000010110;
					assign node243 = (inp[2]) ? node255 : node244;
						assign node244 = (inp[5]) ? node248 : node245;
							assign node245 = (inp[9]) ? 11'b10111111010 : 11'b10011101000;
							assign node248 = (inp[0]) ? node252 : node249;
								assign node249 = (inp[10]) ? 11'b00100000001 : 11'b10101010101;
								assign node252 = (inp[11]) ? 11'b00010110001 : 11'b00100110001;
						assign node255 = (inp[10]) ? node263 : node256;
							assign node256 = (inp[0]) ? node260 : node257;
								assign node257 = (inp[11]) ? 11'b10111000010 : 11'b10101000011;
								assign node260 = (inp[11]) ? 11'b00011010010 : 11'b00111000010;
							assign node263 = (inp[0]) ? 11'b00000000000 : 11'b00111000100;
			assign node266 = (inp[2]) ? node300 : node267;
				assign node267 = (inp[6]) ? node285 : node268;
					assign node268 = (inp[11]) ? node280 : node269;
						assign node269 = (inp[8]) ? node275 : node270;
							assign node270 = (inp[0]) ? 11'b00001110001 : node271;
								assign node271 = (inp[3]) ? 11'b00110110001 : 11'b00010110001;
							assign node275 = (inp[10]) ? node277 : 11'b10011100111;
								assign node277 = (inp[3]) ? 11'b00000100001 : 11'b10010000001;
						assign node280 = (inp[9]) ? 11'b00101000011 : node281;
							assign node281 = (inp[10]) ? 11'b00101100001 : 11'b00111110001;
					assign node285 = (inp[5]) ? node295 : node286;
						assign node286 = (inp[9]) ? node292 : node287;
							assign node287 = (inp[0]) ? 11'b00000100010 : node288;
								assign node288 = (inp[11]) ? 11'b00001100000 : 11'b00101100010;
							assign node292 = (inp[3]) ? 11'b00000100000 : 11'b10010110100;
						assign node295 = (inp[11]) ? node297 : 11'b00000010100;
							assign node297 = (inp[9]) ? 11'b10110000000 : 11'b10010010010;
				assign node300 = (inp[5]) ? node310 : node301;
					assign node301 = (inp[11]) ? node307 : node302;
						assign node302 = (inp[10]) ? node304 : 11'b00010000111;
							assign node304 = (inp[3]) ? 11'b00101010110 : 11'b10101000011;
						assign node307 = (inp[10]) ? 11'b00001110000 : 11'b00111000000;
					assign node310 = (inp[3]) ? node326 : node311;
						assign node311 = (inp[0]) ? node319 : node312;
							assign node312 = (inp[4]) ? node316 : node313;
								assign node313 = (inp[10]) ? 11'b10110010010 : 11'b00100010000;
								assign node316 = (inp[9]) ? 11'b00010010110 : 11'b10110000100;
							assign node319 = (inp[6]) ? node323 : node320;
								assign node320 = (inp[9]) ? 11'b00110100100 : 11'b00001110100;
								assign node323 = (inp[11]) ? 11'b00000010000 : 11'b00100000100;
						assign node326 = (inp[9]) ? node334 : node327;
							assign node327 = (inp[6]) ? node331 : node328;
								assign node328 = (inp[4]) ? 11'b00000010010 : 11'b00100000110;
								assign node331 = (inp[10]) ? 11'b00010010100 : 11'b10000010110;
							assign node334 = (inp[0]) ? 11'b00001000000 : 11'b00000000000;

endmodule