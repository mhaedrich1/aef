module dtc_split5_bm22 (
	input  wire [11-1:0] inp,
	output wire [11-1:0] outp
);

	wire [11-1:0] node1;
	wire [11-1:0] node2;
	wire [11-1:0] node3;
	wire [11-1:0] node4;
	wire [11-1:0] node5;
	wire [11-1:0] node6;
	wire [11-1:0] node7;
	wire [11-1:0] node8;
	wire [11-1:0] node11;
	wire [11-1:0] node14;
	wire [11-1:0] node15;
	wire [11-1:0] node18;
	wire [11-1:0] node21;
	wire [11-1:0] node22;
	wire [11-1:0] node23;
	wire [11-1:0] node26;
	wire [11-1:0] node29;
	wire [11-1:0] node30;
	wire [11-1:0] node33;
	wire [11-1:0] node36;
	wire [11-1:0] node37;
	wire [11-1:0] node38;
	wire [11-1:0] node39;
	wire [11-1:0] node42;
	wire [11-1:0] node45;
	wire [11-1:0] node46;
	wire [11-1:0] node49;
	wire [11-1:0] node52;
	wire [11-1:0] node53;
	wire [11-1:0] node54;
	wire [11-1:0] node57;
	wire [11-1:0] node60;
	wire [11-1:0] node61;
	wire [11-1:0] node64;
	wire [11-1:0] node67;
	wire [11-1:0] node68;
	wire [11-1:0] node69;
	wire [11-1:0] node70;
	wire [11-1:0] node71;
	wire [11-1:0] node75;
	wire [11-1:0] node76;
	wire [11-1:0] node79;
	wire [11-1:0] node82;
	wire [11-1:0] node83;
	wire [11-1:0] node84;
	wire [11-1:0] node87;
	wire [11-1:0] node90;
	wire [11-1:0] node91;
	wire [11-1:0] node94;
	wire [11-1:0] node97;
	wire [11-1:0] node98;
	wire [11-1:0] node99;
	wire [11-1:0] node100;
	wire [11-1:0] node103;
	wire [11-1:0] node106;
	wire [11-1:0] node107;
	wire [11-1:0] node110;
	wire [11-1:0] node113;
	wire [11-1:0] node114;
	wire [11-1:0] node116;
	wire [11-1:0] node119;
	wire [11-1:0] node120;
	wire [11-1:0] node123;
	wire [11-1:0] node126;
	wire [11-1:0] node127;
	wire [11-1:0] node128;
	wire [11-1:0] node129;
	wire [11-1:0] node130;
	wire [11-1:0] node131;
	wire [11-1:0] node134;
	wire [11-1:0] node137;
	wire [11-1:0] node138;
	wire [11-1:0] node141;
	wire [11-1:0] node144;
	wire [11-1:0] node145;
	wire [11-1:0] node146;
	wire [11-1:0] node149;
	wire [11-1:0] node152;
	wire [11-1:0] node153;
	wire [11-1:0] node156;
	wire [11-1:0] node159;
	wire [11-1:0] node160;
	wire [11-1:0] node161;
	wire [11-1:0] node162;
	wire [11-1:0] node165;
	wire [11-1:0] node168;
	wire [11-1:0] node169;
	wire [11-1:0] node172;
	wire [11-1:0] node175;
	wire [11-1:0] node176;
	wire [11-1:0] node177;
	wire [11-1:0] node180;
	wire [11-1:0] node183;
	wire [11-1:0] node184;
	wire [11-1:0] node187;
	wire [11-1:0] node190;
	wire [11-1:0] node191;
	wire [11-1:0] node192;
	wire [11-1:0] node194;
	wire [11-1:0] node195;
	wire [11-1:0] node198;
	wire [11-1:0] node201;
	wire [11-1:0] node202;
	wire [11-1:0] node203;
	wire [11-1:0] node206;
	wire [11-1:0] node209;
	wire [11-1:0] node210;
	wire [11-1:0] node213;
	wire [11-1:0] node216;
	wire [11-1:0] node217;
	wire [11-1:0] node218;
	wire [11-1:0] node219;
	wire [11-1:0] node222;
	wire [11-1:0] node225;
	wire [11-1:0] node226;
	wire [11-1:0] node229;
	wire [11-1:0] node232;
	wire [11-1:0] node233;
	wire [11-1:0] node234;
	wire [11-1:0] node237;
	wire [11-1:0] node240;
	wire [11-1:0] node241;
	wire [11-1:0] node244;
	wire [11-1:0] node247;
	wire [11-1:0] node248;
	wire [11-1:0] node249;
	wire [11-1:0] node250;
	wire [11-1:0] node251;
	wire [11-1:0] node252;
	wire [11-1:0] node253;
	wire [11-1:0] node256;
	wire [11-1:0] node259;
	wire [11-1:0] node260;
	wire [11-1:0] node263;
	wire [11-1:0] node266;
	wire [11-1:0] node267;
	wire [11-1:0] node268;
	wire [11-1:0] node271;
	wire [11-1:0] node274;
	wire [11-1:0] node275;
	wire [11-1:0] node278;
	wire [11-1:0] node281;
	wire [11-1:0] node282;
	wire [11-1:0] node283;
	wire [11-1:0] node284;
	wire [11-1:0] node287;
	wire [11-1:0] node290;
	wire [11-1:0] node291;
	wire [11-1:0] node294;
	wire [11-1:0] node297;
	wire [11-1:0] node298;
	wire [11-1:0] node299;
	wire [11-1:0] node302;
	wire [11-1:0] node305;
	wire [11-1:0] node306;
	wire [11-1:0] node309;
	wire [11-1:0] node312;
	wire [11-1:0] node313;
	wire [11-1:0] node314;
	wire [11-1:0] node315;
	wire [11-1:0] node316;
	wire [11-1:0] node319;
	wire [11-1:0] node322;
	wire [11-1:0] node323;
	wire [11-1:0] node326;
	wire [11-1:0] node329;
	wire [11-1:0] node330;
	wire [11-1:0] node332;
	wire [11-1:0] node335;
	wire [11-1:0] node336;
	wire [11-1:0] node340;
	wire [11-1:0] node341;
	wire [11-1:0] node342;
	wire [11-1:0] node343;
	wire [11-1:0] node346;
	wire [11-1:0] node349;
	wire [11-1:0] node350;
	wire [11-1:0] node354;
	wire [11-1:0] node355;
	wire [11-1:0] node356;
	wire [11-1:0] node359;
	wire [11-1:0] node362;
	wire [11-1:0] node363;
	wire [11-1:0] node366;
	wire [11-1:0] node369;
	wire [11-1:0] node370;
	wire [11-1:0] node371;
	wire [11-1:0] node372;
	wire [11-1:0] node373;
	wire [11-1:0] node374;
	wire [11-1:0] node377;
	wire [11-1:0] node380;
	wire [11-1:0] node381;
	wire [11-1:0] node384;
	wire [11-1:0] node387;
	wire [11-1:0] node388;
	wire [11-1:0] node389;
	wire [11-1:0] node392;
	wire [11-1:0] node395;
	wire [11-1:0] node396;
	wire [11-1:0] node399;
	wire [11-1:0] node402;
	wire [11-1:0] node403;
	wire [11-1:0] node404;
	wire [11-1:0] node405;
	wire [11-1:0] node408;
	wire [11-1:0] node411;
	wire [11-1:0] node412;
	wire [11-1:0] node415;
	wire [11-1:0] node418;
	wire [11-1:0] node419;
	wire [11-1:0] node420;
	wire [11-1:0] node423;
	wire [11-1:0] node426;
	wire [11-1:0] node427;
	wire [11-1:0] node430;
	wire [11-1:0] node433;
	wire [11-1:0] node434;
	wire [11-1:0] node435;
	wire [11-1:0] node436;
	wire [11-1:0] node437;
	wire [11-1:0] node440;
	wire [11-1:0] node443;
	wire [11-1:0] node444;
	wire [11-1:0] node447;
	wire [11-1:0] node450;
	wire [11-1:0] node451;
	wire [11-1:0] node452;
	wire [11-1:0] node455;
	wire [11-1:0] node458;
	wire [11-1:0] node459;
	wire [11-1:0] node462;
	wire [11-1:0] node465;
	wire [11-1:0] node466;
	wire [11-1:0] node467;
	wire [11-1:0] node468;
	wire [11-1:0] node471;
	wire [11-1:0] node474;
	wire [11-1:0] node475;
	wire [11-1:0] node478;
	wire [11-1:0] node481;
	wire [11-1:0] node482;
	wire [11-1:0] node483;
	wire [11-1:0] node486;
	wire [11-1:0] node489;
	wire [11-1:0] node490;
	wire [11-1:0] node493;
	wire [11-1:0] node496;
	wire [11-1:0] node497;
	wire [11-1:0] node498;
	wire [11-1:0] node499;
	wire [11-1:0] node500;
	wire [11-1:0] node501;
	wire [11-1:0] node502;
	wire [11-1:0] node503;
	wire [11-1:0] node506;
	wire [11-1:0] node509;
	wire [11-1:0] node510;
	wire [11-1:0] node513;
	wire [11-1:0] node516;
	wire [11-1:0] node517;
	wire [11-1:0] node518;
	wire [11-1:0] node521;
	wire [11-1:0] node524;
	wire [11-1:0] node525;
	wire [11-1:0] node528;
	wire [11-1:0] node531;
	wire [11-1:0] node532;
	wire [11-1:0] node533;
	wire [11-1:0] node534;
	wire [11-1:0] node537;
	wire [11-1:0] node540;
	wire [11-1:0] node541;
	wire [11-1:0] node544;
	wire [11-1:0] node547;
	wire [11-1:0] node548;
	wire [11-1:0] node549;
	wire [11-1:0] node552;
	wire [11-1:0] node555;
	wire [11-1:0] node556;
	wire [11-1:0] node559;
	wire [11-1:0] node562;
	wire [11-1:0] node563;
	wire [11-1:0] node564;
	wire [11-1:0] node565;
	wire [11-1:0] node566;
	wire [11-1:0] node569;
	wire [11-1:0] node572;
	wire [11-1:0] node573;
	wire [11-1:0] node576;
	wire [11-1:0] node579;
	wire [11-1:0] node580;
	wire [11-1:0] node581;
	wire [11-1:0] node584;
	wire [11-1:0] node587;
	wire [11-1:0] node588;
	wire [11-1:0] node591;
	wire [11-1:0] node594;
	wire [11-1:0] node595;
	wire [11-1:0] node596;
	wire [11-1:0] node597;
	wire [11-1:0] node600;
	wire [11-1:0] node603;
	wire [11-1:0] node604;
	wire [11-1:0] node607;
	wire [11-1:0] node610;
	wire [11-1:0] node611;
	wire [11-1:0] node612;
	wire [11-1:0] node615;
	wire [11-1:0] node618;
	wire [11-1:0] node619;
	wire [11-1:0] node622;
	wire [11-1:0] node625;
	wire [11-1:0] node626;
	wire [11-1:0] node627;
	wire [11-1:0] node628;
	wire [11-1:0] node629;
	wire [11-1:0] node630;
	wire [11-1:0] node633;
	wire [11-1:0] node636;
	wire [11-1:0] node637;
	wire [11-1:0] node640;
	wire [11-1:0] node643;
	wire [11-1:0] node644;
	wire [11-1:0] node645;
	wire [11-1:0] node648;
	wire [11-1:0] node651;
	wire [11-1:0] node652;
	wire [11-1:0] node655;
	wire [11-1:0] node658;
	wire [11-1:0] node659;
	wire [11-1:0] node660;
	wire [11-1:0] node661;
	wire [11-1:0] node664;
	wire [11-1:0] node667;
	wire [11-1:0] node668;
	wire [11-1:0] node671;
	wire [11-1:0] node674;
	wire [11-1:0] node675;
	wire [11-1:0] node676;
	wire [11-1:0] node679;
	wire [11-1:0] node682;
	wire [11-1:0] node683;
	wire [11-1:0] node686;
	wire [11-1:0] node689;
	wire [11-1:0] node690;
	wire [11-1:0] node691;
	wire [11-1:0] node692;
	wire [11-1:0] node693;
	wire [11-1:0] node696;
	wire [11-1:0] node699;
	wire [11-1:0] node700;
	wire [11-1:0] node703;
	wire [11-1:0] node706;
	wire [11-1:0] node707;
	wire [11-1:0] node709;
	wire [11-1:0] node712;
	wire [11-1:0] node714;
	wire [11-1:0] node717;
	wire [11-1:0] node718;
	wire [11-1:0] node719;
	wire [11-1:0] node720;
	wire [11-1:0] node723;
	wire [11-1:0] node726;
	wire [11-1:0] node727;
	wire [11-1:0] node730;
	wire [11-1:0] node733;
	wire [11-1:0] node734;
	wire [11-1:0] node736;
	wire [11-1:0] node739;
	wire [11-1:0] node741;
	wire [11-1:0] node744;
	wire [11-1:0] node745;
	wire [11-1:0] node746;
	wire [11-1:0] node747;
	wire [11-1:0] node748;
	wire [11-1:0] node749;
	wire [11-1:0] node750;
	wire [11-1:0] node753;
	wire [11-1:0] node756;
	wire [11-1:0] node757;
	wire [11-1:0] node761;
	wire [11-1:0] node762;
	wire [11-1:0] node763;
	wire [11-1:0] node766;
	wire [11-1:0] node769;
	wire [11-1:0] node770;
	wire [11-1:0] node773;
	wire [11-1:0] node776;
	wire [11-1:0] node777;
	wire [11-1:0] node778;
	wire [11-1:0] node779;
	wire [11-1:0] node783;
	wire [11-1:0] node784;
	wire [11-1:0] node787;
	wire [11-1:0] node790;
	wire [11-1:0] node791;
	wire [11-1:0] node793;
	wire [11-1:0] node796;
	wire [11-1:0] node797;
	wire [11-1:0] node800;
	wire [11-1:0] node803;
	wire [11-1:0] node804;
	wire [11-1:0] node805;
	wire [11-1:0] node806;
	wire [11-1:0] node807;
	wire [11-1:0] node810;
	wire [11-1:0] node813;
	wire [11-1:0] node814;
	wire [11-1:0] node817;
	wire [11-1:0] node820;
	wire [11-1:0] node821;
	wire [11-1:0] node822;
	wire [11-1:0] node825;
	wire [11-1:0] node828;
	wire [11-1:0] node829;
	wire [11-1:0] node832;
	wire [11-1:0] node835;
	wire [11-1:0] node836;
	wire [11-1:0] node837;
	wire [11-1:0] node838;
	wire [11-1:0] node841;
	wire [11-1:0] node844;
	wire [11-1:0] node845;
	wire [11-1:0] node849;
	wire [11-1:0] node850;
	wire [11-1:0] node851;
	wire [11-1:0] node854;
	wire [11-1:0] node857;
	wire [11-1:0] node858;
	wire [11-1:0] node861;
	wire [11-1:0] node864;
	wire [11-1:0] node865;
	wire [11-1:0] node866;
	wire [11-1:0] node867;
	wire [11-1:0] node868;
	wire [11-1:0] node869;
	wire [11-1:0] node872;
	wire [11-1:0] node875;
	wire [11-1:0] node876;
	wire [11-1:0] node879;
	wire [11-1:0] node882;
	wire [11-1:0] node883;
	wire [11-1:0] node885;
	wire [11-1:0] node888;
	wire [11-1:0] node889;
	wire [11-1:0] node892;
	wire [11-1:0] node895;
	wire [11-1:0] node896;
	wire [11-1:0] node897;
	wire [11-1:0] node898;
	wire [11-1:0] node901;
	wire [11-1:0] node904;
	wire [11-1:0] node905;
	wire [11-1:0] node908;
	wire [11-1:0] node911;
	wire [11-1:0] node912;
	wire [11-1:0] node913;
	wire [11-1:0] node916;
	wire [11-1:0] node919;
	wire [11-1:0] node920;
	wire [11-1:0] node923;
	wire [11-1:0] node926;
	wire [11-1:0] node927;
	wire [11-1:0] node928;
	wire [11-1:0] node929;
	wire [11-1:0] node930;
	wire [11-1:0] node933;
	wire [11-1:0] node936;
	wire [11-1:0] node937;
	wire [11-1:0] node940;
	wire [11-1:0] node943;
	wire [11-1:0] node944;
	wire [11-1:0] node945;
	wire [11-1:0] node948;
	wire [11-1:0] node951;
	wire [11-1:0] node952;
	wire [11-1:0] node955;
	wire [11-1:0] node958;
	wire [11-1:0] node959;
	wire [11-1:0] node960;
	wire [11-1:0] node961;
	wire [11-1:0] node964;
	wire [11-1:0] node967;
	wire [11-1:0] node968;
	wire [11-1:0] node971;
	wire [11-1:0] node974;
	wire [11-1:0] node975;
	wire [11-1:0] node976;
	wire [11-1:0] node979;
	wire [11-1:0] node982;
	wire [11-1:0] node984;

	assign outp = (inp[0]) ? node496 : node1;
		assign node1 = (inp[2]) ? node247 : node2;
			assign node2 = (inp[9]) ? node126 : node3;
				assign node3 = (inp[1]) ? node67 : node4;
					assign node4 = (inp[10]) ? node36 : node5;
						assign node5 = (inp[7]) ? node21 : node6;
							assign node6 = (inp[4]) ? node14 : node7;
								assign node7 = (inp[3]) ? node11 : node8;
									assign node8 = (inp[8]) ? 11'b00111111111 : 11'b01111111111;
									assign node11 = (inp[5]) ? 11'b00011111111 : 11'b00111111111;
								assign node14 = (inp[8]) ? node18 : node15;
									assign node15 = (inp[6]) ? 11'b00011111111 : 11'b00011111111;
									assign node18 = (inp[3]) ? 11'b00001111111 : 11'b00001111111;
							assign node21 = (inp[8]) ? node29 : node22;
								assign node22 = (inp[6]) ? node26 : node23;
									assign node23 = (inp[4]) ? 11'b00011111111 : 11'b00111111111;
									assign node26 = (inp[5]) ? 11'b00001111111 : 11'b00011111111;
								assign node29 = (inp[5]) ? node33 : node30;
									assign node30 = (inp[3]) ? 11'b00001111111 : 11'b00111111111;
									assign node33 = (inp[3]) ? 11'b00000111111 : 11'b00001111111;
						assign node36 = (inp[8]) ? node52 : node37;
							assign node37 = (inp[3]) ? node45 : node38;
								assign node38 = (inp[5]) ? node42 : node39;
									assign node39 = (inp[4]) ? 11'b00011111111 : 11'b00111111111;
									assign node42 = (inp[4]) ? 11'b00001111111 : 11'b00011111111;
								assign node45 = (inp[6]) ? node49 : node46;
									assign node46 = (inp[7]) ? 11'b00001111111 : 11'b00011111111;
									assign node49 = (inp[4]) ? 11'b00000111111 : 11'b00001111111;
							assign node52 = (inp[6]) ? node60 : node53;
								assign node53 = (inp[3]) ? node57 : node54;
									assign node54 = (inp[5]) ? 11'b00001111111 : 11'b00011111111;
									assign node57 = (inp[7]) ? 11'b00000111111 : 11'b00001111111;
								assign node60 = (inp[4]) ? node64 : node61;
									assign node61 = (inp[3]) ? 11'b00000111111 : 11'b00001111111;
									assign node64 = (inp[7]) ? 11'b00000011111 : 11'b00000111111;
					assign node67 = (inp[4]) ? node97 : node68;
						assign node68 = (inp[3]) ? node82 : node69;
							assign node69 = (inp[10]) ? node75 : node70;
								assign node70 = (inp[6]) ? 11'b00011111111 : node71;
									assign node71 = (inp[7]) ? 11'b00011111111 : 11'b00111111111;
								assign node75 = (inp[7]) ? node79 : node76;
									assign node76 = (inp[8]) ? 11'b00001111111 : 11'b00011111111;
									assign node79 = (inp[8]) ? 11'b00000111111 : 11'b00001111111;
							assign node82 = (inp[7]) ? node90 : node83;
								assign node83 = (inp[5]) ? node87 : node84;
									assign node84 = (inp[10]) ? 11'b00001111111 : 11'b00011111111;
									assign node87 = (inp[6]) ? 11'b00000111111 : 11'b00001111111;
								assign node90 = (inp[8]) ? node94 : node91;
									assign node91 = (inp[6]) ? 11'b00000111111 : 11'b00000111111;
									assign node94 = (inp[10]) ? 11'b00000011111 : 11'b00000111111;
						assign node97 = (inp[6]) ? node113 : node98;
							assign node98 = (inp[5]) ? node106 : node99;
								assign node99 = (inp[3]) ? node103 : node100;
									assign node100 = (inp[8]) ? 11'b00001111111 : 11'b00011111111;
									assign node103 = (inp[7]) ? 11'b00000111111 : 11'b00001111111;
								assign node106 = (inp[10]) ? node110 : node107;
									assign node107 = (inp[8]) ? 11'b00000111111 : 11'b00001111111;
									assign node110 = (inp[7]) ? 11'b00000011111 : 11'b00000111111;
							assign node113 = (inp[3]) ? node119 : node114;
								assign node114 = (inp[10]) ? node116 : 11'b00000111111;
									assign node116 = (inp[8]) ? 11'b00000011111 : 11'b00000111111;
								assign node119 = (inp[10]) ? node123 : node120;
									assign node120 = (inp[7]) ? 11'b00000011111 : 11'b00000111111;
									assign node123 = (inp[5]) ? 11'b00000000111 : 11'b00000011111;
				assign node126 = (inp[1]) ? node190 : node127;
					assign node127 = (inp[4]) ? node159 : node128;
						assign node128 = (inp[10]) ? node144 : node129;
							assign node129 = (inp[3]) ? node137 : node130;
								assign node130 = (inp[6]) ? node134 : node131;
									assign node131 = (inp[8]) ? 11'b00011111111 : 11'b00111111111;
									assign node134 = (inp[7]) ? 11'b00000111111 : 11'b00011111111;
								assign node137 = (inp[7]) ? node141 : node138;
									assign node138 = (inp[6]) ? 11'b00001111111 : 11'b00011111111;
									assign node141 = (inp[8]) ? 11'b00000111111 : 11'b00001111111;
							assign node144 = (inp[3]) ? node152 : node145;
								assign node145 = (inp[5]) ? node149 : node146;
									assign node146 = (inp[6]) ? 11'b00001111111 : 11'b00011111111;
									assign node149 = (inp[7]) ? 11'b00000111111 : 11'b00001111111;
								assign node152 = (inp[8]) ? node156 : node153;
									assign node153 = (inp[7]) ? 11'b00000011111 : 11'b00000111111;
									assign node156 = (inp[7]) ? 11'b00000111111 : 11'b00000111111;
						assign node159 = (inp[6]) ? node175 : node160;
							assign node160 = (inp[8]) ? node168 : node161;
								assign node161 = (inp[3]) ? node165 : node162;
									assign node162 = (inp[7]) ? 11'b00001111111 : 11'b00011111111;
									assign node165 = (inp[5]) ? 11'b00000011111 : 11'b00001111111;
								assign node168 = (inp[10]) ? node172 : node169;
									assign node169 = (inp[7]) ? 11'b00000111111 : 11'b00001111111;
									assign node172 = (inp[3]) ? 11'b00000011111 : 11'b00000111111;
							assign node175 = (inp[3]) ? node183 : node176;
								assign node176 = (inp[10]) ? node180 : node177;
									assign node177 = (inp[8]) ? 11'b00000111111 : 11'b00001111111;
									assign node180 = (inp[8]) ? 11'b00000011111 : 11'b00000111111;
								assign node183 = (inp[7]) ? node187 : node184;
									assign node184 = (inp[8]) ? 11'b00000011111 : 11'b00000111111;
									assign node187 = (inp[10]) ? 11'b00000001111 : 11'b00000011111;
					assign node190 = (inp[8]) ? node216 : node191;
						assign node191 = (inp[4]) ? node201 : node192;
							assign node192 = (inp[7]) ? node194 : 11'b00001111111;
								assign node194 = (inp[3]) ? node198 : node195;
									assign node195 = (inp[5]) ? 11'b00000111111 : 11'b00001111111;
									assign node198 = (inp[5]) ? 11'b00000011111 : 11'b00000111111;
							assign node201 = (inp[5]) ? node209 : node202;
								assign node202 = (inp[7]) ? node206 : node203;
									assign node203 = (inp[6]) ? 11'b00000111111 : 11'b00001111111;
									assign node206 = (inp[3]) ? 11'b00000011111 : 11'b00000111111;
								assign node209 = (inp[3]) ? node213 : node210;
									assign node210 = (inp[6]) ? 11'b00000011111 : 11'b00000111111;
									assign node213 = (inp[7]) ? 11'b00000000111 : 11'b00000001111;
						assign node216 = (inp[3]) ? node232 : node217;
							assign node217 = (inp[7]) ? node225 : node218;
								assign node218 = (inp[4]) ? node222 : node219;
									assign node219 = (inp[6]) ? 11'b00000111111 : 11'b00000111111;
									assign node222 = (inp[6]) ? 11'b00000011111 : 11'b00000111111;
								assign node225 = (inp[4]) ? node229 : node226;
									assign node226 = (inp[6]) ? 11'b00000011111 : 11'b00001111111;
									assign node229 = (inp[5]) ? 11'b00000001111 : 11'b00000011111;
							assign node232 = (inp[10]) ? node240 : node233;
								assign node233 = (inp[4]) ? node237 : node234;
									assign node234 = (inp[6]) ? 11'b00000011111 : 11'b00000111111;
									assign node237 = (inp[7]) ? 11'b00000001111 : 11'b00000011111;
								assign node240 = (inp[5]) ? node244 : node241;
									assign node241 = (inp[4]) ? 11'b00000001111 : 11'b00000001111;
									assign node244 = (inp[4]) ? 11'b00000000011 : 11'b00000000111;
			assign node247 = (inp[5]) ? node369 : node248;
				assign node248 = (inp[3]) ? node312 : node249;
					assign node249 = (inp[6]) ? node281 : node250;
						assign node250 = (inp[10]) ? node266 : node251;
							assign node251 = (inp[8]) ? node259 : node252;
								assign node252 = (inp[4]) ? node256 : node253;
									assign node253 = (inp[1]) ? 11'b00011111111 : 11'b00111111111;
									assign node256 = (inp[1]) ? 11'b00000111111 : 11'b00011111111;
								assign node259 = (inp[1]) ? node263 : node260;
									assign node260 = (inp[4]) ? 11'b00001111111 : 11'b00001111111;
									assign node263 = (inp[9]) ? 11'b00000111111 : 11'b00001111111;
							assign node266 = (inp[4]) ? node274 : node267;
								assign node267 = (inp[9]) ? node271 : node268;
									assign node268 = (inp[8]) ? 11'b00001111111 : 11'b00001111111;
									assign node271 = (inp[7]) ? 11'b00001111111 : 11'b00001111111;
								assign node274 = (inp[9]) ? node278 : node275;
									assign node275 = (inp[8]) ? 11'b00000111111 : 11'b00001111111;
									assign node278 = (inp[7]) ? 11'b00000011111 : 11'b00000111111;
						assign node281 = (inp[1]) ? node297 : node282;
							assign node282 = (inp[10]) ? node290 : node283;
								assign node283 = (inp[8]) ? node287 : node284;
									assign node284 = (inp[7]) ? 11'b00001111111 : 11'b00111111111;
									assign node287 = (inp[4]) ? 11'b00000111111 : 11'b00001111111;
								assign node290 = (inp[7]) ? node294 : node291;
									assign node291 = (inp[8]) ? 11'b00000111111 : 11'b00011111111;
									assign node294 = (inp[8]) ? 11'b00000011111 : 11'b00000111111;
							assign node297 = (inp[4]) ? node305 : node298;
								assign node298 = (inp[7]) ? node302 : node299;
									assign node299 = (inp[10]) ? 11'b00000111111 : 11'b00001111111;
									assign node302 = (inp[8]) ? 11'b00000011111 : 11'b00000111111;
								assign node305 = (inp[10]) ? node309 : node306;
									assign node306 = (inp[9]) ? 11'b00000011111 : 11'b00000111111;
									assign node309 = (inp[8]) ? 11'b00000001111 : 11'b00000011111;
					assign node312 = (inp[7]) ? node340 : node313;
						assign node313 = (inp[9]) ? node329 : node314;
							assign node314 = (inp[1]) ? node322 : node315;
								assign node315 = (inp[6]) ? node319 : node316;
									assign node316 = (inp[8]) ? 11'b00001111111 : 11'b00011111111;
									assign node319 = (inp[8]) ? 11'b00000111111 : 11'b00001111111;
								assign node322 = (inp[4]) ? node326 : node323;
									assign node323 = (inp[6]) ? 11'b00000111111 : 11'b00001111111;
									assign node326 = (inp[6]) ? 11'b00000011111 : 11'b00000111111;
							assign node329 = (inp[6]) ? node335 : node330;
								assign node330 = (inp[4]) ? node332 : 11'b00001111111;
									assign node332 = (inp[8]) ? 11'b00000011111 : 11'b00000111111;
								assign node335 = (inp[10]) ? 11'b00000011111 : node336;
									assign node336 = (inp[4]) ? 11'b00000011111 : 11'b00000111111;
						assign node340 = (inp[4]) ? node354 : node341;
							assign node341 = (inp[1]) ? node349 : node342;
								assign node342 = (inp[6]) ? node346 : node343;
									assign node343 = (inp[9]) ? 11'b00000111111 : 11'b00001111111;
									assign node346 = (inp[9]) ? 11'b00000011111 : 11'b00000111111;
								assign node349 = (inp[9]) ? 11'b00000001111 : node350;
									assign node350 = (inp[10]) ? 11'b00000011111 : 11'b00000111111;
							assign node354 = (inp[8]) ? node362 : node355;
								assign node355 = (inp[1]) ? node359 : node356;
									assign node356 = (inp[6]) ? 11'b00000001111 : 11'b00000111111;
									assign node359 = (inp[9]) ? 11'b00000001111 : 11'b00000011111;
								assign node362 = (inp[10]) ? node366 : node363;
									assign node363 = (inp[6]) ? 11'b00000001111 : 11'b00000011111;
									assign node366 = (inp[6]) ? 11'b00000000111 : 11'b00000001111;
				assign node369 = (inp[9]) ? node433 : node370;
					assign node370 = (inp[10]) ? node402 : node371;
						assign node371 = (inp[8]) ? node387 : node372;
							assign node372 = (inp[6]) ? node380 : node373;
								assign node373 = (inp[1]) ? node377 : node374;
									assign node374 = (inp[3]) ? 11'b00001111111 : 11'b00001111111;
									assign node377 = (inp[7]) ? 11'b00000111111 : 11'b00001111111;
								assign node380 = (inp[4]) ? node384 : node381;
									assign node381 = (inp[3]) ? 11'b00000111111 : 11'b00001111111;
									assign node384 = (inp[1]) ? 11'b00000001111 : 11'b00000111111;
							assign node387 = (inp[6]) ? node395 : node388;
								assign node388 = (inp[4]) ? node392 : node389;
									assign node389 = (inp[1]) ? 11'b00000111111 : 11'b00001111111;
									assign node392 = (inp[3]) ? 11'b00000011111 : 11'b00000011111;
								assign node395 = (inp[7]) ? node399 : node396;
									assign node396 = (inp[3]) ? 11'b00000011111 : 11'b00000111111;
									assign node399 = (inp[3]) ? 11'b00000001111 : 11'b00000011111;
						assign node402 = (inp[3]) ? node418 : node403;
							assign node403 = (inp[1]) ? node411 : node404;
								assign node404 = (inp[7]) ? node408 : node405;
									assign node405 = (inp[6]) ? 11'b00000111111 : 11'b00000111111;
									assign node408 = (inp[4]) ? 11'b00000011111 : 11'b00000111111;
								assign node411 = (inp[7]) ? node415 : node412;
									assign node412 = (inp[8]) ? 11'b00000001111 : 11'b00000111111;
									assign node415 = (inp[4]) ? 11'b00000001111 : 11'b00000011111;
							assign node418 = (inp[7]) ? node426 : node419;
								assign node419 = (inp[8]) ? node423 : node420;
									assign node420 = (inp[1]) ? 11'b00000011111 : 11'b00000111111;
									assign node423 = (inp[4]) ? 11'b00000001111 : 11'b00000011111;
								assign node426 = (inp[6]) ? node430 : node427;
									assign node427 = (inp[1]) ? 11'b00000011111 : 11'b00000001111;
									assign node430 = (inp[1]) ? 11'b00000000111 : 11'b00000001111;
					assign node433 = (inp[10]) ? node465 : node434;
						assign node434 = (inp[8]) ? node450 : node435;
							assign node435 = (inp[4]) ? node443 : node436;
								assign node436 = (inp[3]) ? node440 : node437;
									assign node437 = (inp[1]) ? 11'b00001111111 : 11'b00011111111;
									assign node440 = (inp[7]) ? 11'b00000011111 : 11'b00000111111;
								assign node443 = (inp[3]) ? node447 : node444;
									assign node444 = (inp[1]) ? 11'b00000011111 : 11'b00000111111;
									assign node447 = (inp[7]) ? 11'b00000001111 : 11'b00000011111;
							assign node450 = (inp[7]) ? node458 : node451;
								assign node451 = (inp[1]) ? node455 : node452;
									assign node452 = (inp[3]) ? 11'b00000011111 : 11'b00000111111;
									assign node455 = (inp[4]) ? 11'b00000001111 : 11'b00000011111;
								assign node458 = (inp[4]) ? node462 : node459;
									assign node459 = (inp[3]) ? 11'b00000001111 : 11'b00000011111;
									assign node462 = (inp[1]) ? 11'b00000000111 : 11'b00000001111;
						assign node465 = (inp[3]) ? node481 : node466;
							assign node466 = (inp[6]) ? node474 : node467;
								assign node467 = (inp[7]) ? node471 : node468;
									assign node468 = (inp[1]) ? 11'b00000011111 : 11'b00000111111;
									assign node471 = (inp[8]) ? 11'b00000001111 : 11'b00000011111;
								assign node474 = (inp[1]) ? node478 : node475;
									assign node475 = (inp[4]) ? 11'b00000001111 : 11'b00000011111;
									assign node478 = (inp[4]) ? 11'b00000000011 : 11'b00000001111;
							assign node481 = (inp[1]) ? node489 : node482;
								assign node482 = (inp[4]) ? node486 : node483;
									assign node483 = (inp[7]) ? 11'b00000001111 : 11'b00000001111;
									assign node486 = (inp[6]) ? 11'b00000000111 : 11'b00000000111;
								assign node489 = (inp[8]) ? node493 : node490;
									assign node490 = (inp[6]) ? 11'b00000000111 : 11'b00000001111;
									assign node493 = (inp[7]) ? 11'b00000000011 : 11'b00000000011;
		assign node496 = (inp[10]) ? node744 : node497;
			assign node497 = (inp[4]) ? node625 : node498;
				assign node498 = (inp[7]) ? node562 : node499;
					assign node499 = (inp[2]) ? node531 : node500;
						assign node500 = (inp[8]) ? node516 : node501;
							assign node501 = (inp[1]) ? node509 : node502;
								assign node502 = (inp[3]) ? node506 : node503;
									assign node503 = (inp[6]) ? 11'b00011111111 : 11'b00111111111;
									assign node506 = (inp[6]) ? 11'b00001111111 : 11'b00011111111;
								assign node509 = (inp[6]) ? node513 : node510;
									assign node510 = (inp[3]) ? 11'b00001111111 : 11'b00011111111;
									assign node513 = (inp[9]) ? 11'b00000111111 : 11'b00001111111;
							assign node516 = (inp[5]) ? node524 : node517;
								assign node517 = (inp[9]) ? node521 : node518;
									assign node518 = (inp[6]) ? 11'b00001111111 : 11'b00011111111;
									assign node521 = (inp[3]) ? 11'b00000111111 : 11'b00001111111;
								assign node524 = (inp[1]) ? node528 : node525;
									assign node525 = (inp[6]) ? 11'b00000111111 : 11'b00001111111;
									assign node528 = (inp[3]) ? 11'b00000011111 : 11'b00000111111;
						assign node531 = (inp[9]) ? node547 : node532;
							assign node532 = (inp[3]) ? node540 : node533;
								assign node533 = (inp[1]) ? node537 : node534;
									assign node534 = (inp[6]) ? 11'b00001111111 : 11'b00011111111;
									assign node537 = (inp[8]) ? 11'b00000111111 : 11'b00001111111;
								assign node540 = (inp[5]) ? node544 : node541;
									assign node541 = (inp[8]) ? 11'b00000111111 : 11'b00001111111;
									assign node544 = (inp[6]) ? 11'b00000011111 : 11'b00000111111;
							assign node547 = (inp[1]) ? node555 : node548;
								assign node548 = (inp[5]) ? node552 : node549;
									assign node549 = (inp[3]) ? 11'b00000111111 : 11'b00001111111;
									assign node552 = (inp[8]) ? 11'b00000001111 : 11'b00000111111;
								assign node555 = (inp[5]) ? node559 : node556;
									assign node556 = (inp[8]) ? 11'b00000011111 : 11'b00000011111;
									assign node559 = (inp[6]) ? 11'b00000001111 : 11'b00000011111;
					assign node562 = (inp[3]) ? node594 : node563;
						assign node563 = (inp[5]) ? node579 : node564;
							assign node564 = (inp[9]) ? node572 : node565;
								assign node565 = (inp[6]) ? node569 : node566;
									assign node566 = (inp[8]) ? 11'b00001111111 : 11'b00011111111;
									assign node569 = (inp[1]) ? 11'b00000111111 : 11'b00001111111;
								assign node572 = (inp[1]) ? node576 : node573;
									assign node573 = (inp[2]) ? 11'b00000111111 : 11'b00001111111;
									assign node576 = (inp[6]) ? 11'b00000011111 : 11'b00000111111;
							assign node579 = (inp[8]) ? node587 : node580;
								assign node580 = (inp[9]) ? node584 : node581;
									assign node581 = (inp[1]) ? 11'b00000111111 : 11'b00001111111;
									assign node584 = (inp[2]) ? 11'b00000011111 : 11'b00000111111;
								assign node587 = (inp[1]) ? node591 : node588;
									assign node588 = (inp[6]) ? 11'b00000011111 : 11'b00000111111;
									assign node591 = (inp[9]) ? 11'b00000001111 : 11'b00000011111;
						assign node594 = (inp[2]) ? node610 : node595;
							assign node595 = (inp[5]) ? node603 : node596;
								assign node596 = (inp[9]) ? node600 : node597;
									assign node597 = (inp[1]) ? 11'b00000111111 : 11'b00001111111;
									assign node600 = (inp[8]) ? 11'b00000011111 : 11'b00000111111;
								assign node603 = (inp[8]) ? node607 : node604;
									assign node604 = (inp[1]) ? 11'b00000011111 : 11'b00000111111;
									assign node607 = (inp[9]) ? 11'b00000001111 : 11'b00000001111;
							assign node610 = (inp[9]) ? node618 : node611;
								assign node611 = (inp[6]) ? node615 : node612;
									assign node612 = (inp[5]) ? 11'b00000011111 : 11'b00001111111;
									assign node615 = (inp[5]) ? 11'b00000001111 : 11'b00000011111;
								assign node618 = (inp[5]) ? node622 : node619;
									assign node619 = (inp[8]) ? 11'b00000001111 : 11'b00000011111;
									assign node622 = (inp[8]) ? 11'b00000000011 : 11'b00000001111;
				assign node625 = (inp[5]) ? node689 : node626;
					assign node626 = (inp[6]) ? node658 : node627;
						assign node627 = (inp[9]) ? node643 : node628;
							assign node628 = (inp[1]) ? node636 : node629;
								assign node629 = (inp[2]) ? node633 : node630;
									assign node630 = (inp[7]) ? 11'b00001111111 : 11'b00011111111;
									assign node633 = (inp[3]) ? 11'b00000111111 : 11'b00001111111;
								assign node636 = (inp[8]) ? node640 : node637;
									assign node637 = (inp[3]) ? 11'b00000111111 : 11'b00001111111;
									assign node640 = (inp[7]) ? 11'b00000011111 : 11'b00000111111;
							assign node643 = (inp[1]) ? node651 : node644;
								assign node644 = (inp[2]) ? node648 : node645;
									assign node645 = (inp[8]) ? 11'b00000111111 : 11'b00001111111;
									assign node648 = (inp[3]) ? 11'b00000011111 : 11'b00000011111;
								assign node651 = (inp[7]) ? node655 : node652;
									assign node652 = (inp[8]) ? 11'b00000111111 : 11'b00000011111;
									assign node655 = (inp[3]) ? 11'b00000001111 : 11'b00000011111;
						assign node658 = (inp[3]) ? node674 : node659;
							assign node659 = (inp[7]) ? node667 : node660;
								assign node660 = (inp[8]) ? node664 : node661;
									assign node661 = (inp[1]) ? 11'b00000111111 : 11'b00001111111;
									assign node664 = (inp[1]) ? 11'b00000011111 : 11'b00000111111;
								assign node667 = (inp[1]) ? node671 : node668;
									assign node668 = (inp[9]) ? 11'b00000011111 : 11'b00000111111;
									assign node671 = (inp[2]) ? 11'b00000001111 : 11'b00000011111;
							assign node674 = (inp[1]) ? node682 : node675;
								assign node675 = (inp[7]) ? node679 : node676;
									assign node676 = (inp[8]) ? 11'b00000011111 : 11'b00000011111;
									assign node679 = (inp[9]) ? 11'b00000001111 : 11'b00000011111;
								assign node682 = (inp[9]) ? node686 : node683;
									assign node683 = (inp[7]) ? 11'b00000001111 : 11'b00000011111;
									assign node686 = (inp[2]) ? 11'b00000000111 : 11'b00000000111;
					assign node689 = (inp[1]) ? node717 : node690;
						assign node690 = (inp[9]) ? node706 : node691;
							assign node691 = (inp[7]) ? node699 : node692;
								assign node692 = (inp[8]) ? node696 : node693;
									assign node693 = (inp[3]) ? 11'b00000111111 : 11'b00001111111;
									assign node696 = (inp[6]) ? 11'b00000001111 : 11'b00000111111;
								assign node699 = (inp[2]) ? node703 : node700;
									assign node700 = (inp[6]) ? 11'b00000011111 : 11'b00000111111;
									assign node703 = (inp[8]) ? 11'b00000001111 : 11'b00000001111;
							assign node706 = (inp[6]) ? node712 : node707;
								assign node707 = (inp[2]) ? node709 : 11'b00000011111;
									assign node709 = (inp[8]) ? 11'b00000000111 : 11'b00000011111;
								assign node712 = (inp[8]) ? node714 : 11'b00000001111;
									assign node714 = (inp[3]) ? 11'b00000000111 : 11'b00000001111;
						assign node717 = (inp[2]) ? node733 : node718;
							assign node718 = (inp[6]) ? node726 : node719;
								assign node719 = (inp[8]) ? node723 : node720;
									assign node720 = (inp[7]) ? 11'b00000011111 : 11'b00000111111;
									assign node723 = (inp[9]) ? 11'b00000001111 : 11'b00000011111;
								assign node726 = (inp[3]) ? node730 : node727;
									assign node727 = (inp[7]) ? 11'b00000001111 : 11'b00000011111;
									assign node730 = (inp[9]) ? 11'b00000000111 : 11'b00000001111;
							assign node733 = (inp[9]) ? node739 : node734;
								assign node734 = (inp[7]) ? node736 : 11'b00000011111;
									assign node736 = (inp[6]) ? 11'b00000000111 : 11'b00000000111;
								assign node739 = (inp[6]) ? node741 : 11'b00000000111;
									assign node741 = (inp[7]) ? 11'b00000000001 : 11'b00000000111;
			assign node744 = (inp[5]) ? node864 : node745;
				assign node745 = (inp[3]) ? node803 : node746;
					assign node746 = (inp[8]) ? node776 : node747;
						assign node747 = (inp[7]) ? node761 : node748;
							assign node748 = (inp[2]) ? node756 : node749;
								assign node749 = (inp[1]) ? node753 : node750;
									assign node750 = (inp[9]) ? 11'b00001111111 : 11'b00011111111;
									assign node753 = (inp[9]) ? 11'b00000011111 : 11'b00001111111;
								assign node756 = (inp[6]) ? 11'b00000111111 : node757;
									assign node757 = (inp[1]) ? 11'b00000111111 : 11'b00001111111;
							assign node761 = (inp[2]) ? node769 : node762;
								assign node762 = (inp[9]) ? node766 : node763;
									assign node763 = (inp[1]) ? 11'b00000111111 : 11'b00001111111;
									assign node766 = (inp[6]) ? 11'b00000011111 : 11'b00000111111;
								assign node769 = (inp[1]) ? node773 : node770;
									assign node770 = (inp[6]) ? 11'b00000011111 : 11'b00000111111;
									assign node773 = (inp[9]) ? 11'b00000000111 : 11'b00000011111;
						assign node776 = (inp[6]) ? node790 : node777;
							assign node777 = (inp[9]) ? node783 : node778;
								assign node778 = (inp[2]) ? 11'b00000111111 : node779;
									assign node779 = (inp[7]) ? 11'b00000111111 : 11'b00000111111;
								assign node783 = (inp[1]) ? node787 : node784;
									assign node784 = (inp[7]) ? 11'b00000011111 : 11'b00000111111;
									assign node787 = (inp[2]) ? 11'b00000000111 : 11'b00000011111;
							assign node790 = (inp[9]) ? node796 : node791;
								assign node791 = (inp[2]) ? node793 : 11'b00000011111;
									assign node793 = (inp[1]) ? 11'b00000001111 : 11'b00000011111;
								assign node796 = (inp[4]) ? node800 : node797;
									assign node797 = (inp[7]) ? 11'b00000001111 : 11'b00000011111;
									assign node800 = (inp[2]) ? 11'b00000000111 : 11'b00000000111;
					assign node803 = (inp[9]) ? node835 : node804;
						assign node804 = (inp[2]) ? node820 : node805;
							assign node805 = (inp[4]) ? node813 : node806;
								assign node806 = (inp[1]) ? node810 : node807;
									assign node807 = (inp[7]) ? 11'b00000111111 : 11'b00001111111;
									assign node810 = (inp[6]) ? 11'b00000011111 : 11'b00000111111;
								assign node813 = (inp[6]) ? node817 : node814;
									assign node814 = (inp[8]) ? 11'b00000011111 : 11'b00000111111;
									assign node817 = (inp[7]) ? 11'b00000001111 : 11'b00000011111;
							assign node820 = (inp[6]) ? node828 : node821;
								assign node821 = (inp[1]) ? node825 : node822;
									assign node822 = (inp[7]) ? 11'b00000011111 : 11'b00000111111;
									assign node825 = (inp[8]) ? 11'b00000001111 : 11'b00000011111;
								assign node828 = (inp[1]) ? node832 : node829;
									assign node829 = (inp[7]) ? 11'b00000001111 : 11'b00000011111;
									assign node832 = (inp[4]) ? 11'b00000000111 : 11'b00000001111;
						assign node835 = (inp[4]) ? node849 : node836;
							assign node836 = (inp[6]) ? node844 : node837;
								assign node837 = (inp[2]) ? node841 : node838;
									assign node838 = (inp[1]) ? 11'b00000011111 : 11'b00000011111;
									assign node841 = (inp[7]) ? 11'b00000001111 : 11'b00000011111;
								assign node844 = (inp[2]) ? 11'b00000000111 : node845;
									assign node845 = (inp[1]) ? 11'b00000001111 : 11'b00000001111;
							assign node849 = (inp[8]) ? node857 : node850;
								assign node850 = (inp[6]) ? node854 : node851;
									assign node851 = (inp[2]) ? 11'b00000001111 : 11'b00000011111;
									assign node854 = (inp[7]) ? 11'b00000000111 : 11'b00000001111;
								assign node857 = (inp[7]) ? node861 : node858;
									assign node858 = (inp[2]) ? 11'b00000000111 : 11'b00000001111;
									assign node861 = (inp[2]) ? 11'b00000000011 : 11'b00000000111;
				assign node864 = (inp[2]) ? node926 : node865;
					assign node865 = (inp[7]) ? node895 : node866;
						assign node866 = (inp[8]) ? node882 : node867;
							assign node867 = (inp[3]) ? node875 : node868;
								assign node868 = (inp[6]) ? node872 : node869;
									assign node869 = (inp[9]) ? 11'b00000111111 : 11'b00001111111;
									assign node872 = (inp[4]) ? 11'b00000011111 : 11'b00000111111;
								assign node875 = (inp[1]) ? node879 : node876;
									assign node876 = (inp[6]) ? 11'b00000011111 : 11'b00000111111;
									assign node879 = (inp[6]) ? 11'b00000001111 : 11'b00000011111;
							assign node882 = (inp[3]) ? node888 : node883;
								assign node883 = (inp[4]) ? node885 : 11'b00000111111;
									assign node885 = (inp[1]) ? 11'b00000001111 : 11'b00000011111;
								assign node888 = (inp[4]) ? node892 : node889;
									assign node889 = (inp[9]) ? 11'b00000001111 : 11'b00000001111;
									assign node892 = (inp[1]) ? 11'b00000000111 : 11'b00000001111;
						assign node895 = (inp[9]) ? node911 : node896;
							assign node896 = (inp[1]) ? node904 : node897;
								assign node897 = (inp[8]) ? node901 : node898;
									assign node898 = (inp[3]) ? 11'b00000011111 : 11'b00000111111;
									assign node901 = (inp[4]) ? 11'b00000001111 : 11'b00000011111;
								assign node904 = (inp[4]) ? node908 : node905;
									assign node905 = (inp[6]) ? 11'b00000001111 : 11'b00000011111;
									assign node908 = (inp[3]) ? 11'b00000000111 : 11'b00000001111;
							assign node911 = (inp[3]) ? node919 : node912;
								assign node912 = (inp[1]) ? node916 : node913;
									assign node913 = (inp[4]) ? 11'b00000001111 : 11'b00000011111;
									assign node916 = (inp[4]) ? 11'b00000000111 : 11'b00000001111;
								assign node919 = (inp[1]) ? node923 : node920;
									assign node920 = (inp[4]) ? 11'b00000000111 : 11'b00000000111;
									assign node923 = (inp[8]) ? 11'b00000000011 : 11'b00000000111;
					assign node926 = (inp[7]) ? node958 : node927;
						assign node927 = (inp[8]) ? node943 : node928;
							assign node928 = (inp[3]) ? node936 : node929;
								assign node929 = (inp[6]) ? node933 : node930;
									assign node930 = (inp[4]) ? 11'b00000011111 : 11'b00000011111;
									assign node933 = (inp[1]) ? 11'b00000001111 : 11'b00000011111;
								assign node936 = (inp[4]) ? node940 : node937;
									assign node937 = (inp[9]) ? 11'b00000001111 : 11'b00000011111;
									assign node940 = (inp[6]) ? 11'b00000000111 : 11'b00000000111;
							assign node943 = (inp[1]) ? node951 : node944;
								assign node944 = (inp[9]) ? node948 : node945;
									assign node945 = (inp[3]) ? 11'b00000001111 : 11'b00000011111;
									assign node948 = (inp[6]) ? 11'b00000000111 : 11'b00000001111;
								assign node951 = (inp[6]) ? node955 : node952;
									assign node952 = (inp[9]) ? 11'b00000000111 : 11'b00000000111;
									assign node955 = (inp[4]) ? 11'b00000000011 : 11'b00000000111;
						assign node958 = (inp[1]) ? node974 : node959;
							assign node959 = (inp[9]) ? node967 : node960;
								assign node960 = (inp[6]) ? node964 : node961;
									assign node961 = (inp[4]) ? 11'b00000001111 : 11'b00000111111;
									assign node964 = (inp[8]) ? 11'b00000000111 : 11'b00000001111;
								assign node967 = (inp[6]) ? node971 : node968;
									assign node968 = (inp[3]) ? 11'b00000000111 : 11'b00000001111;
									assign node971 = (inp[4]) ? 11'b00000000001 : 11'b00000000111;
							assign node974 = (inp[8]) ? node982 : node975;
								assign node975 = (inp[9]) ? node979 : node976;
									assign node976 = (inp[3]) ? 11'b00000000011 : 11'b00000001111;
									assign node979 = (inp[6]) ? 11'b00000000001 : 11'b00000000111;
								assign node982 = (inp[3]) ? node984 : 11'b00000000011;
									assign node984 = (inp[9]) ? 11'b00000000001 : 11'b00000000001;

endmodule