module dtc_split66_bm64 (
	input  wire [16-1:0] inp,
	output wire [4-1:0] outp
);

	wire [4-1:0] node2;
	wire [4-1:0] node3;
	wire [4-1:0] node4;
	wire [4-1:0] node5;
	wire [4-1:0] node6;
	wire [4-1:0] node7;
	wire [4-1:0] node8;
	wire [4-1:0] node9;
	wire [4-1:0] node10;
	wire [4-1:0] node11;
	wire [4-1:0] node12;
	wire [4-1:0] node14;
	wire [4-1:0] node16;
	wire [4-1:0] node17;
	wire [4-1:0] node22;
	wire [4-1:0] node24;
	wire [4-1:0] node25;
	wire [4-1:0] node26;
	wire [4-1:0] node30;
	wire [4-1:0] node32;
	wire [4-1:0] node34;
	wire [4-1:0] node38;
	wire [4-1:0] node40;
	wire [4-1:0] node41;
	wire [4-1:0] node42;
	wire [4-1:0] node43;
	wire [4-1:0] node45;
	wire [4-1:0] node48;
	wire [4-1:0] node50;
	wire [4-1:0] node52;
	wire [4-1:0] node56;
	wire [4-1:0] node58;
	wire [4-1:0] node59;
	wire [4-1:0] node60;
	wire [4-1:0] node64;
	wire [4-1:0] node66;
	wire [4-1:0] node67;
	wire [4-1:0] node72;
	wire [4-1:0] node74;
	wire [4-1:0] node75;
	wire [4-1:0] node76;
	wire [4-1:0] node77;
	wire [4-1:0] node78;
	wire [4-1:0] node79;
	wire [4-1:0] node80;
	wire [4-1:0] node82;
	wire [4-1:0] node86;
	wire [4-1:0] node88;
	wire [4-1:0] node89;
	wire [4-1:0] node94;
	wire [4-1:0] node96;
	wire [4-1:0] node97;
	wire [4-1:0] node98;
	wire [4-1:0] node100;
	wire [4-1:0] node104;
	wire [4-1:0] node106;
	wire [4-1:0] node107;
	wire [4-1:0] node112;
	wire [4-1:0] node114;
	wire [4-1:0] node115;
	wire [4-1:0] node116;
	wire [4-1:0] node117;
	wire [4-1:0] node118;
	wire [4-1:0] node119;
	wire [4-1:0] node124;
	wire [4-1:0] node126;
	wire [4-1:0] node127;
	wire [4-1:0] node132;
	wire [4-1:0] node134;
	wire [4-1:0] node135;
	wire [4-1:0] node136;
	wire [4-1:0] node137;
	wire [4-1:0] node142;
	wire [4-1:0] node144;
	wire [4-1:0] node148;
	wire [4-1:0] node149;
	wire [4-1:0] node150;
	wire [4-1:0] node151;
	wire [4-1:0] node152;
	wire [4-1:0] node153;
	wire [4-1:0] node154;
	wire [4-1:0] node155;
	wire [4-1:0] node156;
	wire [4-1:0] node158;
	wire [4-1:0] node162;
	wire [4-1:0] node164;
	wire [4-1:0] node168;
	wire [4-1:0] node170;
	wire [4-1:0] node171;
	wire [4-1:0] node172;
	wire [4-1:0] node173;
	wire [4-1:0] node178;
	wire [4-1:0] node179;
	wire [4-1:0] node181;
	wire [4-1:0] node186;
	wire [4-1:0] node188;
	wire [4-1:0] node189;
	wire [4-1:0] node190;
	wire [4-1:0] node191;
	wire [4-1:0] node193;
	wire [4-1:0] node194;
	wire [4-1:0] node198;
	wire [4-1:0] node200;
	wire [4-1:0] node201;
	wire [4-1:0] node206;
	wire [4-1:0] node208;
	wire [4-1:0] node209;
	wire [4-1:0] node210;
	wire [4-1:0] node214;
	wire [4-1:0] node216;
	wire [4-1:0] node218;
	wire [4-1:0] node221;
	wire [4-1:0] node222;
	wire [4-1:0] node223;
	wire [4-1:0] node225;
	wire [4-1:0] node226;
	wire [4-1:0] node227;
	wire [4-1:0] node229;
	wire [4-1:0] node230;
	wire [4-1:0] node234;
	wire [4-1:0] node235;
	wire [4-1:0] node237;
	wire [4-1:0] node238;
	wire [4-1:0] node245;
	wire [4-1:0] node246;
	wire [4-1:0] node248;
	wire [4-1:0] node249;
	wire [4-1:0] node250;
	wire [4-1:0] node251;
	wire [4-1:0] node253;
	wire [4-1:0] node255;
	wire [4-1:0] node258;
	wire [4-1:0] node260;
	wire [4-1:0] node265;
	wire [4-1:0] node266;
	wire [4-1:0] node267;
	wire [4-1:0] node269;
	wire [4-1:0] node270;
	wire [4-1:0] node271;
	wire [4-1:0] node272;
	wire [4-1:0] node279;
	wire [4-1:0] node280;
	wire [4-1:0] node282;
	wire [4-1:0] node284;
	wire [4-1:0] node286;
	wire [4-1:0] node289;
	wire [4-1:0] node290;
	wire [4-1:0] node291;
	wire [4-1:0] node293;
	wire [4-1:0] node297;
	wire [4-1:0] node299;
	wire [4-1:0] node300;
	wire [4-1:0] node301;
	wire [4-1:0] node306;
	wire [4-1:0] node308;
	wire [4-1:0] node309;
	wire [4-1:0] node310;
	wire [4-1:0] node311;
	wire [4-1:0] node312;
	wire [4-1:0] node313;
	wire [4-1:0] node314;
	wire [4-1:0] node315;
	wire [4-1:0] node320;
	wire [4-1:0] node322;
	wire [4-1:0] node324;
	wire [4-1:0] node328;
	wire [4-1:0] node330;
	wire [4-1:0] node331;
	wire [4-1:0] node332;
	wire [4-1:0] node334;
	wire [4-1:0] node338;
	wire [4-1:0] node340;
	wire [4-1:0] node341;
	wire [4-1:0] node346;
	wire [4-1:0] node348;
	wire [4-1:0] node349;
	wire [4-1:0] node350;
	wire [4-1:0] node351;
	wire [4-1:0] node352;
	wire [4-1:0] node353;
	wire [4-1:0] node358;
	wire [4-1:0] node360;
	wire [4-1:0] node362;
	wire [4-1:0] node366;
	wire [4-1:0] node368;
	wire [4-1:0] node369;
	wire [4-1:0] node370;
	wire [4-1:0] node371;
	wire [4-1:0] node376;
	wire [4-1:0] node377;
	wire [4-1:0] node379;
	wire [4-1:0] node383;
	wire [4-1:0] node384;
	wire [4-1:0] node386;
	wire [4-1:0] node387;
	wire [4-1:0] node388;
	wire [4-1:0] node389;
	wire [4-1:0] node390;
	wire [4-1:0] node391;
	wire [4-1:0] node392;
	wire [4-1:0] node393;
	wire [4-1:0] node394;
	wire [4-1:0] node395;
	wire [4-1:0] node402;
	wire [4-1:0] node404;
	wire [4-1:0] node405;
	wire [4-1:0] node406;
	wire [4-1:0] node408;
	wire [4-1:0] node412;
	wire [4-1:0] node413;
	wire [4-1:0] node415;
	wire [4-1:0] node420;
	wire [4-1:0] node422;
	wire [4-1:0] node423;
	wire [4-1:0] node424;
	wire [4-1:0] node425;
	wire [4-1:0] node426;
	wire [4-1:0] node430;
	wire [4-1:0] node432;
	wire [4-1:0] node436;
	wire [4-1:0] node438;
	wire [4-1:0] node439;
	wire [4-1:0] node440;
	wire [4-1:0] node444;
	wire [4-1:0] node446;
	wire [4-1:0] node447;
	wire [4-1:0] node452;
	wire [4-1:0] node454;
	wire [4-1:0] node455;
	wire [4-1:0] node456;
	wire [4-1:0] node457;
	wire [4-1:0] node458;
	wire [4-1:0] node459;
	wire [4-1:0] node460;
	wire [4-1:0] node466;
	wire [4-1:0] node468;
	wire [4-1:0] node469;
	wire [4-1:0] node471;
	wire [4-1:0] node474;
	wire [4-1:0] node476;
	wire [4-1:0] node480;
	wire [4-1:0] node482;
	wire [4-1:0] node483;
	wire [4-1:0] node484;
	wire [4-1:0] node485;
	wire [4-1:0] node486;
	wire [4-1:0] node487;
	wire [4-1:0] node492;
	wire [4-1:0] node494;
	wire [4-1:0] node496;
	wire [4-1:0] node500;
	wire [4-1:0] node502;
	wire [4-1:0] node503;
	wire [4-1:0] node505;
	wire [4-1:0] node508;
	wire [4-1:0] node509;
	wire [4-1:0] node510;
	wire [4-1:0] node514;
	wire [4-1:0] node516;
	wire [4-1:0] node519;
	wire [4-1:0] node520;
	wire [4-1:0] node521;
	wire [4-1:0] node522;
	wire [4-1:0] node523;
	wire [4-1:0] node524;
	wire [4-1:0] node525;
	wire [4-1:0] node526;
	wire [4-1:0] node527;
	wire [4-1:0] node532;
	wire [4-1:0] node534;
	wire [4-1:0] node536;
	wire [4-1:0] node539;
	wire [4-1:0] node540;
	wire [4-1:0] node542;
	wire [4-1:0] node543;
	wire [4-1:0] node548;
	wire [4-1:0] node550;
	wire [4-1:0] node551;
	wire [4-1:0] node552;
	wire [4-1:0] node554;
	wire [4-1:0] node558;
	wire [4-1:0] node560;
	wire [4-1:0] node562;
	wire [4-1:0] node565;
	wire [4-1:0] node566;
	wire [4-1:0] node567;
	wire [4-1:0] node568;
	wire [4-1:0] node569;
	wire [4-1:0] node570;
	wire [4-1:0] node572;
	wire [4-1:0] node574;
	wire [4-1:0] node577;
	wire [4-1:0] node578;
	wire [4-1:0] node583;
	wire [4-1:0] node585;
	wire [4-1:0] node586;
	wire [4-1:0] node587;
	wire [4-1:0] node592;
	wire [4-1:0] node594;
	wire [4-1:0] node595;
	wire [4-1:0] node596;
	wire [4-1:0] node598;
	wire [4-1:0] node603;
	wire [4-1:0] node605;
	wire [4-1:0] node606;
	wire [4-1:0] node607;
	wire [4-1:0] node609;
	wire [4-1:0] node610;
	wire [4-1:0] node615;
	wire [4-1:0] node616;
	wire [4-1:0] node618;
	wire [4-1:0] node619;
	wire [4-1:0] node624;
	wire [4-1:0] node625;
	wire [4-1:0] node626;
	wire [4-1:0] node627;
	wire [4-1:0] node628;
	wire [4-1:0] node629;
	wire [4-1:0] node632;
	wire [4-1:0] node634;
	wire [4-1:0] node635;
	wire [4-1:0] node639;
	wire [4-1:0] node640;
	wire [4-1:0] node641;
	wire [4-1:0] node642;
	wire [4-1:0] node647;
	wire [4-1:0] node650;
	wire [4-1:0] node651;
	wire [4-1:0] node652;
	wire [4-1:0] node654;
	wire [4-1:0] node656;
	wire [4-1:0] node657;
	wire [4-1:0] node661;
	wire [4-1:0] node663;
	wire [4-1:0] node665;
	wire [4-1:0] node668;
	wire [4-1:0] node669;
	wire [4-1:0] node672;
	wire [4-1:0] node673;
	wire [4-1:0] node677;
	wire [4-1:0] node678;
	wire [4-1:0] node679;
	wire [4-1:0] node680;
	wire [4-1:0] node682;
	wire [4-1:0] node685;
	wire [4-1:0] node687;
	wire [4-1:0] node689;
	wire [4-1:0] node692;
	wire [4-1:0] node693;
	wire [4-1:0] node695;
	wire [4-1:0] node698;
	wire [4-1:0] node699;
	wire [4-1:0] node701;
	wire [4-1:0] node705;
	wire [4-1:0] node706;
	wire [4-1:0] node707;
	wire [4-1:0] node708;
	wire [4-1:0] node709;
	wire [4-1:0] node710;
	wire [4-1:0] node713;
	wire [4-1:0] node716;
	wire [4-1:0] node717;
	wire [4-1:0] node719;
	wire [4-1:0] node723;
	wire [4-1:0] node724;
	wire [4-1:0] node726;
	wire [4-1:0] node729;
	wire [4-1:0] node730;
	wire [4-1:0] node733;
	wire [4-1:0] node736;
	wire [4-1:0] node737;
	wire [4-1:0] node738;
	wire [4-1:0] node739;
	wire [4-1:0] node741;
	wire [4-1:0] node745;
	wire [4-1:0] node748;
	wire [4-1:0] node749;
	wire [4-1:0] node751;
	wire [4-1:0] node752;
	wire [4-1:0] node756;
	wire [4-1:0] node758;
	wire [4-1:0] node759;
	wire [4-1:0] node763;
	wire [4-1:0] node764;
	wire [4-1:0] node765;
	wire [4-1:0] node767;
	wire [4-1:0] node768;
	wire [4-1:0] node770;
	wire [4-1:0] node773;
	wire [4-1:0] node776;
	wire [4-1:0] node778;
	wire [4-1:0] node779;
	wire [4-1:0] node782;
	wire [4-1:0] node783;
	wire [4-1:0] node787;
	wire [4-1:0] node788;
	wire [4-1:0] node790;
	wire [4-1:0] node793;
	wire [4-1:0] node794;
	wire [4-1:0] node797;
	wire [4-1:0] node798;
	wire [4-1:0] node802;
	wire [4-1:0] node803;
	wire [4-1:0] node804;
	wire [4-1:0] node805;
	wire [4-1:0] node806;
	wire [4-1:0] node807;
	wire [4-1:0] node808;
	wire [4-1:0] node809;
	wire [4-1:0] node814;
	wire [4-1:0] node815;
	wire [4-1:0] node817;
	wire [4-1:0] node820;
	wire [4-1:0] node821;
	wire [4-1:0] node825;
	wire [4-1:0] node826;
	wire [4-1:0] node827;
	wire [4-1:0] node831;
	wire [4-1:0] node834;
	wire [4-1:0] node835;
	wire [4-1:0] node837;
	wire [4-1:0] node838;
	wire [4-1:0] node840;
	wire [4-1:0] node844;
	wire [4-1:0] node846;
	wire [4-1:0] node848;
	wire [4-1:0] node851;
	wire [4-1:0] node852;
	wire [4-1:0] node853;
	wire [4-1:0] node855;
	wire [4-1:0] node856;
	wire [4-1:0] node861;
	wire [4-1:0] node862;
	wire [4-1:0] node864;
	wire [4-1:0] node865;
	wire [4-1:0] node869;
	wire [4-1:0] node872;
	wire [4-1:0] node873;
	wire [4-1:0] node874;
	wire [4-1:0] node875;
	wire [4-1:0] node877;
	wire [4-1:0] node880;
	wire [4-1:0] node882;
	wire [4-1:0] node883;
	wire [4-1:0] node887;
	wire [4-1:0] node888;
	wire [4-1:0] node890;
	wire [4-1:0] node892;
	wire [4-1:0] node894;
	wire [4-1:0] node897;
	wire [4-1:0] node898;
	wire [4-1:0] node900;
	wire [4-1:0] node904;
	wire [4-1:0] node905;
	wire [4-1:0] node906;
	wire [4-1:0] node907;
	wire [4-1:0] node911;
	wire [4-1:0] node913;
	wire [4-1:0] node914;
	wire [4-1:0] node918;
	wire [4-1:0] node921;
	wire [4-1:0] node922;
	wire [4-1:0] node923;
	wire [4-1:0] node924;
	wire [4-1:0] node925;
	wire [4-1:0] node926;
	wire [4-1:0] node928;
	wire [4-1:0] node930;
	wire [4-1:0] node933;
	wire [4-1:0] node934;
	wire [4-1:0] node935;
	wire [4-1:0] node936;
	wire [4-1:0] node942;
	wire [4-1:0] node943;
	wire [4-1:0] node944;
	wire [4-1:0] node945;
	wire [4-1:0] node947;
	wire [4-1:0] node948;
	wire [4-1:0] node952;
	wire [4-1:0] node953;
	wire [4-1:0] node955;
	wire [4-1:0] node959;
	wire [4-1:0] node960;
	wire [4-1:0] node962;
	wire [4-1:0] node963;
	wire [4-1:0] node967;
	wire [4-1:0] node969;
	wire [4-1:0] node971;
	wire [4-1:0] node974;
	wire [4-1:0] node975;
	wire [4-1:0] node977;
	wire [4-1:0] node978;
	wire [4-1:0] node979;
	wire [4-1:0] node985;
	wire [4-1:0] node986;
	wire [4-1:0] node987;
	wire [4-1:0] node989;
	wire [4-1:0] node990;
	wire [4-1:0] node991;
	wire [4-1:0] node996;
	wire [4-1:0] node997;
	wire [4-1:0] node999;
	wire [4-1:0] node1000;
	wire [4-1:0] node1004;
	wire [4-1:0] node1006;
	wire [4-1:0] node1009;
	wire [4-1:0] node1010;
	wire [4-1:0] node1012;
	wire [4-1:0] node1013;
	wire [4-1:0] node1017;
	wire [4-1:0] node1018;
	wire [4-1:0] node1020;
	wire [4-1:0] node1021;
	wire [4-1:0] node1026;
	wire [4-1:0] node1027;
	wire [4-1:0] node1028;
	wire [4-1:0] node1029;
	wire [4-1:0] node1030;
	wire [4-1:0] node1031;
	wire [4-1:0] node1036;
	wire [4-1:0] node1038;
	wire [4-1:0] node1039;
	wire [4-1:0] node1043;
	wire [4-1:0] node1044;
	wire [4-1:0] node1045;
	wire [4-1:0] node1046;
	wire [4-1:0] node1047;
	wire [4-1:0] node1048;
	wire [4-1:0] node1053;
	wire [4-1:0] node1055;
	wire [4-1:0] node1059;
	wire [4-1:0] node1061;
	wire [4-1:0] node1062;
	wire [4-1:0] node1063;
	wire [4-1:0] node1068;
	wire [4-1:0] node1069;
	wire [4-1:0] node1070;
	wire [4-1:0] node1072;
	wire [4-1:0] node1073;
	wire [4-1:0] node1074;
	wire [4-1:0] node1078;
	wire [4-1:0] node1080;
	wire [4-1:0] node1084;
	wire [4-1:0] node1085;
	wire [4-1:0] node1087;
	wire [4-1:0] node1088;
	wire [4-1:0] node1092;
	wire [4-1:0] node1094;
	wire [4-1:0] node1096;
	wire [4-1:0] node1099;
	wire [4-1:0] node1100;
	wire [4-1:0] node1101;
	wire [4-1:0] node1102;
	wire [4-1:0] node1103;
	wire [4-1:0] node1104;
	wire [4-1:0] node1105;
	wire [4-1:0] node1107;
	wire [4-1:0] node1110;
	wire [4-1:0] node1111;
	wire [4-1:0] node1113;
	wire [4-1:0] node1117;
	wire [4-1:0] node1118;
	wire [4-1:0] node1121;
	wire [4-1:0] node1122;
	wire [4-1:0] node1126;
	wire [4-1:0] node1127;
	wire [4-1:0] node1128;
	wire [4-1:0] node1129;
	wire [4-1:0] node1134;
	wire [4-1:0] node1135;
	wire [4-1:0] node1136;
	wire [4-1:0] node1141;
	wire [4-1:0] node1142;
	wire [4-1:0] node1143;
	wire [4-1:0] node1144;
	wire [4-1:0] node1147;
	wire [4-1:0] node1149;
	wire [4-1:0] node1152;
	wire [4-1:0] node1153;
	wire [4-1:0] node1156;
	wire [4-1:0] node1157;
	wire [4-1:0] node1159;
	wire [4-1:0] node1163;
	wire [4-1:0] node1164;
	wire [4-1:0] node1165;
	wire [4-1:0] node1167;
	wire [4-1:0] node1171;
	wire [4-1:0] node1172;
	wire [4-1:0] node1176;
	wire [4-1:0] node1177;
	wire [4-1:0] node1178;
	wire [4-1:0] node1179;
	wire [4-1:0] node1181;
	wire [4-1:0] node1182;
	wire [4-1:0] node1184;
	wire [4-1:0] node1186;
	wire [4-1:0] node1190;
	wire [4-1:0] node1192;
	wire [4-1:0] node1195;
	wire [4-1:0] node1196;
	wire [4-1:0] node1197;
	wire [4-1:0] node1198;
	wire [4-1:0] node1200;
	wire [4-1:0] node1204;
	wire [4-1:0] node1205;
	wire [4-1:0] node1209;
	wire [4-1:0] node1210;
	wire [4-1:0] node1212;
	wire [4-1:0] node1214;
	wire [4-1:0] node1217;
	wire [4-1:0] node1218;
	wire [4-1:0] node1219;
	wire [4-1:0] node1223;
	wire [4-1:0] node1226;
	wire [4-1:0] node1227;
	wire [4-1:0] node1228;
	wire [4-1:0] node1229;
	wire [4-1:0] node1230;
	wire [4-1:0] node1231;
	wire [4-1:0] node1235;
	wire [4-1:0] node1236;
	wire [4-1:0] node1241;
	wire [4-1:0] node1242;
	wire [4-1:0] node1243;
	wire [4-1:0] node1248;
	wire [4-1:0] node1249;
	wire [4-1:0] node1250;
	wire [4-1:0] node1252;
	wire [4-1:0] node1255;
	wire [4-1:0] node1256;
	wire [4-1:0] node1257;
	wire [4-1:0] node1261;
	wire [4-1:0] node1263;
	wire [4-1:0] node1266;
	wire [4-1:0] node1269;
	wire [4-1:0] node1270;
	wire [4-1:0] node1271;
	wire [4-1:0] node1272;
	wire [4-1:0] node1273;
	wire [4-1:0] node1274;
	wire [4-1:0] node1275;
	wire [4-1:0] node1278;
	wire [4-1:0] node1281;
	wire [4-1:0] node1282;
	wire [4-1:0] node1283;
	wire [4-1:0] node1287;
	wire [4-1:0] node1290;
	wire [4-1:0] node1291;
	wire [4-1:0] node1292;
	wire [4-1:0] node1295;
	wire [4-1:0] node1297;
	wire [4-1:0] node1300;
	wire [4-1:0] node1301;
	wire [4-1:0] node1304;
	wire [4-1:0] node1305;
	wire [4-1:0] node1309;
	wire [4-1:0] node1310;
	wire [4-1:0] node1311;
	wire [4-1:0] node1312;
	wire [4-1:0] node1316;
	wire [4-1:0] node1317;
	wire [4-1:0] node1318;
	wire [4-1:0] node1322;
	wire [4-1:0] node1324;
	wire [4-1:0] node1327;
	wire [4-1:0] node1328;
	wire [4-1:0] node1329;
	wire [4-1:0] node1330;
	wire [4-1:0] node1334;
	wire [4-1:0] node1335;
	wire [4-1:0] node1339;
	wire [4-1:0] node1340;
	wire [4-1:0] node1342;
	wire [4-1:0] node1345;
	wire [4-1:0] node1348;
	wire [4-1:0] node1349;
	wire [4-1:0] node1350;
	wire [4-1:0] node1353;
	wire [4-1:0] node1356;
	wire [4-1:0] node1357;
	wire [4-1:0] node1360;
	wire [4-1:0] node1363;
	wire [4-1:0] node1364;
	wire [4-1:0] node1365;
	wire [4-1:0] node1366;
	wire [4-1:0] node1369;
	wire [4-1:0] node1372;
	wire [4-1:0] node1373;
	wire [4-1:0] node1376;
	wire [4-1:0] node1380;
	wire [4-1:0] node1382;
	wire [4-1:0] node1383;
	wire [4-1:0] node1384;
	wire [4-1:0] node1385;
	wire [4-1:0] node1386;
	wire [4-1:0] node1387;
	wire [4-1:0] node1388;
	wire [4-1:0] node1389;
	wire [4-1:0] node1390;
	wire [4-1:0] node1391;
	wire [4-1:0] node1392;
	wire [4-1:0] node1393;
	wire [4-1:0] node1398;
	wire [4-1:0] node1400;
	wire [4-1:0] node1404;
	wire [4-1:0] node1406;
	wire [4-1:0] node1407;
	wire [4-1:0] node1408;
	wire [4-1:0] node1410;
	wire [4-1:0] node1414;
	wire [4-1:0] node1416;
	wire [4-1:0] node1417;
	wire [4-1:0] node1422;
	wire [4-1:0] node1424;
	wire [4-1:0] node1425;
	wire [4-1:0] node1426;
	wire [4-1:0] node1427;
	wire [4-1:0] node1428;
	wire [4-1:0] node1430;
	wire [4-1:0] node1433;
	wire [4-1:0] node1434;
	wire [4-1:0] node1440;
	wire [4-1:0] node1442;
	wire [4-1:0] node1443;
	wire [4-1:0] node1445;
	wire [4-1:0] node1446;
	wire [4-1:0] node1450;
	wire [4-1:0] node1452;
	wire [4-1:0] node1456;
	wire [4-1:0] node1457;
	wire [4-1:0] node1458;
	wire [4-1:0] node1459;
	wire [4-1:0] node1460;
	wire [4-1:0] node1461;
	wire [4-1:0] node1462;
	wire [4-1:0] node1464;
	wire [4-1:0] node1468;
	wire [4-1:0] node1470;
	wire [4-1:0] node1472;
	wire [4-1:0] node1476;
	wire [4-1:0] node1477;
	wire [4-1:0] node1479;
	wire [4-1:0] node1480;
	wire [4-1:0] node1481;
	wire [4-1:0] node1487;
	wire [4-1:0] node1488;
	wire [4-1:0] node1490;
	wire [4-1:0] node1491;
	wire [4-1:0] node1492;
	wire [4-1:0] node1494;
	wire [4-1:0] node1498;
	wire [4-1:0] node1499;
	wire [4-1:0] node1501;
	wire [4-1:0] node1505;
	wire [4-1:0] node1506;
	wire [4-1:0] node1507;
	wire [4-1:0] node1509;
	wire [4-1:0] node1510;
	wire [4-1:0] node1512;
	wire [4-1:0] node1517;
	wire [4-1:0] node1518;
	wire [4-1:0] node1519;
	wire [4-1:0] node1520;
	wire [4-1:0] node1525;
	wire [4-1:0] node1527;
	wire [4-1:0] node1528;
	wire [4-1:0] node1529;
	wire [4-1:0] node1534;
	wire [4-1:0] node1536;
	wire [4-1:0] node1537;
	wire [4-1:0] node1538;
	wire [4-1:0] node1539;
	wire [4-1:0] node1540;
	wire [4-1:0] node1542;
	wire [4-1:0] node1546;
	wire [4-1:0] node1548;
	wire [4-1:0] node1550;
	wire [4-1:0] node1554;
	wire [4-1:0] node1555;
	wire [4-1:0] node1556;
	wire [4-1:0] node1557;
	wire [4-1:0] node1559;
	wire [4-1:0] node1564;
	wire [4-1:0] node1566;
	wire [4-1:0] node1568;
	wire [4-1:0] node1569;
	wire [4-1:0] node1573;
	wire [4-1:0] node1574;
	wire [4-1:0] node1576;
	wire [4-1:0] node1577;
	wire [4-1:0] node1578;
	wire [4-1:0] node1579;
	wire [4-1:0] node1580;
	wire [4-1:0] node1581;
	wire [4-1:0] node1582;
	wire [4-1:0] node1583;
	wire [4-1:0] node1588;
	wire [4-1:0] node1590;
	wire [4-1:0] node1592;
	wire [4-1:0] node1596;
	wire [4-1:0] node1598;
	wire [4-1:0] node1599;
	wire [4-1:0] node1600;
	wire [4-1:0] node1601;
	wire [4-1:0] node1608;
	wire [4-1:0] node1610;
	wire [4-1:0] node1611;
	wire [4-1:0] node1612;
	wire [4-1:0] node1613;
	wire [4-1:0] node1614;
	wire [4-1:0] node1615;
	wire [4-1:0] node1620;
	wire [4-1:0] node1621;
	wire [4-1:0] node1626;
	wire [4-1:0] node1628;
	wire [4-1:0] node1629;
	wire [4-1:0] node1630;
	wire [4-1:0] node1634;
	wire [4-1:0] node1636;
	wire [4-1:0] node1639;
	wire [4-1:0] node1640;
	wire [4-1:0] node1641;
	wire [4-1:0] node1642;
	wire [4-1:0] node1643;
	wire [4-1:0] node1644;
	wire [4-1:0] node1645;
	wire [4-1:0] node1649;
	wire [4-1:0] node1651;
	wire [4-1:0] node1654;
	wire [4-1:0] node1656;
	wire [4-1:0] node1658;
	wire [4-1:0] node1661;
	wire [4-1:0] node1662;
	wire [4-1:0] node1663;
	wire [4-1:0] node1664;
	wire [4-1:0] node1666;
	wire [4-1:0] node1667;
	wire [4-1:0] node1671;
	wire [4-1:0] node1673;
	wire [4-1:0] node1677;
	wire [4-1:0] node1679;
	wire [4-1:0] node1680;
	wire [4-1:0] node1681;
	wire [4-1:0] node1682;
	wire [4-1:0] node1688;
	wire [4-1:0] node1689;
	wire [4-1:0] node1690;
	wire [4-1:0] node1691;
	wire [4-1:0] node1692;
	wire [4-1:0] node1693;
	wire [4-1:0] node1694;
	wire [4-1:0] node1699;
	wire [4-1:0] node1701;
	wire [4-1:0] node1704;
	wire [4-1:0] node1705;
	wire [4-1:0] node1707;
	wire [4-1:0] node1708;
	wire [4-1:0] node1713;
	wire [4-1:0] node1714;
	wire [4-1:0] node1715;
	wire [4-1:0] node1716;
	wire [4-1:0] node1717;
	wire [4-1:0] node1720;
	wire [4-1:0] node1723;
	wire [4-1:0] node1724;
	wire [4-1:0] node1727;
	wire [4-1:0] node1730;
	wire [4-1:0] node1732;
	wire [4-1:0] node1733;
	wire [4-1:0] node1736;
	wire [4-1:0] node1739;
	wire [4-1:0] node1740;
	wire [4-1:0] node1741;
	wire [4-1:0] node1743;
	wire [4-1:0] node1747;
	wire [4-1:0] node1750;
	wire [4-1:0] node1751;
	wire [4-1:0] node1752;
	wire [4-1:0] node1753;
	wire [4-1:0] node1756;
	wire [4-1:0] node1757;
	wire [4-1:0] node1759;
	wire [4-1:0] node1763;
	wire [4-1:0] node1764;
	wire [4-1:0] node1765;
	wire [4-1:0] node1767;
	wire [4-1:0] node1770;
	wire [4-1:0] node1773;
	wire [4-1:0] node1774;
	wire [4-1:0] node1778;
	wire [4-1:0] node1779;
	wire [4-1:0] node1780;
	wire [4-1:0] node1782;
	wire [4-1:0] node1786;
	wire [4-1:0] node1787;
	wire [4-1:0] node1789;
	wire [4-1:0] node1791;
	wire [4-1:0] node1795;
	wire [4-1:0] node1796;
	wire [4-1:0] node1797;
	wire [4-1:0] node1798;
	wire [4-1:0] node1799;
	wire [4-1:0] node1801;
	wire [4-1:0] node1802;
	wire [4-1:0] node1803;
	wire [4-1:0] node1808;
	wire [4-1:0] node1809;
	wire [4-1:0] node1813;
	wire [4-1:0] node1814;
	wire [4-1:0] node1815;
	wire [4-1:0] node1816;
	wire [4-1:0] node1817;
	wire [4-1:0] node1822;
	wire [4-1:0] node1823;
	wire [4-1:0] node1827;
	wire [4-1:0] node1828;
	wire [4-1:0] node1830;
	wire [4-1:0] node1834;
	wire [4-1:0] node1835;
	wire [4-1:0] node1836;
	wire [4-1:0] node1837;
	wire [4-1:0] node1841;
	wire [4-1:0] node1843;
	wire [4-1:0] node1845;
	wire [4-1:0] node1847;
	wire [4-1:0] node1850;
	wire [4-1:0] node1851;
	wire [4-1:0] node1852;
	wire [4-1:0] node1853;
	wire [4-1:0] node1858;
	wire [4-1:0] node1860;
	wire [4-1:0] node1863;
	wire [4-1:0] node1864;
	wire [4-1:0] node1865;
	wire [4-1:0] node1866;
	wire [4-1:0] node1867;
	wire [4-1:0] node1868;
	wire [4-1:0] node1869;
	wire [4-1:0] node1873;
	wire [4-1:0] node1877;
	wire [4-1:0] node1878;
	wire [4-1:0] node1879;
	wire [4-1:0] node1882;
	wire [4-1:0] node1886;
	wire [4-1:0] node1887;
	wire [4-1:0] node1888;
	wire [4-1:0] node1889;
	wire [4-1:0] node1891;
	wire [4-1:0] node1894;
	wire [4-1:0] node1897;
	wire [4-1:0] node1898;
	wire [4-1:0] node1899;
	wire [4-1:0] node1903;
	wire [4-1:0] node1905;
	wire [4-1:0] node1908;
	wire [4-1:0] node1911;
	wire [4-1:0] node1912;
	wire [4-1:0] node1913;
	wire [4-1:0] node1914;
	wire [4-1:0] node1917;
	wire [4-1:0] node1920;
	wire [4-1:0] node1921;
	wire [4-1:0] node1924;
	wire [4-1:0] node1928;
	wire [4-1:0] node1930;
	wire [4-1:0] node1931;
	wire [4-1:0] node1932;
	wire [4-1:0] node1933;
	wire [4-1:0] node1934;
	wire [4-1:0] node1935;
	wire [4-1:0] node1936;
	wire [4-1:0] node1937;
	wire [4-1:0] node1938;
	wire [4-1:0] node1940;
	wire [4-1:0] node1944;
	wire [4-1:0] node1946;
	wire [4-1:0] node1950;
	wire [4-1:0] node1952;
	wire [4-1:0] node1953;
	wire [4-1:0] node1954;
	wire [4-1:0] node1955;
	wire [4-1:0] node1960;
	wire [4-1:0] node1962;
	wire [4-1:0] node1964;
	wire [4-1:0] node1968;
	wire [4-1:0] node1969;
	wire [4-1:0] node1970;
	wire [4-1:0] node1971;
	wire [4-1:0] node1973;
	wire [4-1:0] node1974;
	wire [4-1:0] node1975;
	wire [4-1:0] node1980;
	wire [4-1:0] node1982;
	wire [4-1:0] node1983;
	wire [4-1:0] node1988;
	wire [4-1:0] node1989;
	wire [4-1:0] node1990;
	wire [4-1:0] node1991;
	wire [4-1:0] node1993;
	wire [4-1:0] node1997;
	wire [4-1:0] node1998;
	wire [4-1:0] node2000;
	wire [4-1:0] node2004;
	wire [4-1:0] node2005;
	wire [4-1:0] node2007;
	wire [4-1:0] node2008;
	wire [4-1:0] node2009;
	wire [4-1:0] node2014;
	wire [4-1:0] node2016;
	wire [4-1:0] node2018;
	wire [4-1:0] node2021;
	wire [4-1:0] node2022;
	wire [4-1:0] node2024;
	wire [4-1:0] node2025;
	wire [4-1:0] node2027;
	wire [4-1:0] node2028;
	wire [4-1:0] node2030;
	wire [4-1:0] node2031;
	wire [4-1:0] node2036;
	wire [4-1:0] node2038;
	wire [4-1:0] node2039;
	wire [4-1:0] node2041;
	wire [4-1:0] node2042;
	wire [4-1:0] node2046;
	wire [4-1:0] node2048;
	wire [4-1:0] node2049;
	wire [4-1:0] node2053;
	wire [4-1:0] node2054;
	wire [4-1:0] node2055;
	wire [4-1:0] node2056;
	wire [4-1:0] node2057;
	wire [4-1:0] node2059;
	wire [4-1:0] node2062;
	wire [4-1:0] node2064;
	wire [4-1:0] node2066;
	wire [4-1:0] node2069;
	wire [4-1:0] node2070;
	wire [4-1:0] node2072;
	wire [4-1:0] node2076;
	wire [4-1:0] node2077;
	wire [4-1:0] node2078;
	wire [4-1:0] node2079;
	wire [4-1:0] node2081;
	wire [4-1:0] node2085;
	wire [4-1:0] node2086;
	wire [4-1:0] node2090;
	wire [4-1:0] node2091;
	wire [4-1:0] node2094;
	wire [4-1:0] node2097;
	wire [4-1:0] node2098;
	wire [4-1:0] node2099;
	wire [4-1:0] node2100;
	wire [4-1:0] node2101;
	wire [4-1:0] node2104;
	wire [4-1:0] node2107;
	wire [4-1:0] node2109;
	wire [4-1:0] node2111;
	wire [4-1:0] node2114;
	wire [4-1:0] node2115;
	wire [4-1:0] node2118;
	wire [4-1:0] node2121;
	wire [4-1:0] node2122;
	wire [4-1:0] node2123;
	wire [4-1:0] node2126;
	wire [4-1:0] node2130;
	wire [4-1:0] node2132;
	wire [4-1:0] node2133;
	wire [4-1:0] node2134;
	wire [4-1:0] node2135;
	wire [4-1:0] node2136;
	wire [4-1:0] node2137;
	wire [4-1:0] node2138;
	wire [4-1:0] node2139;
	wire [4-1:0] node2142;
	wire [4-1:0] node2143;
	wire [4-1:0] node2148;
	wire [4-1:0] node2149;
	wire [4-1:0] node2151;
	wire [4-1:0] node2155;
	wire [4-1:0] node2156;
	wire [4-1:0] node2157;
	wire [4-1:0] node2159;
	wire [4-1:0] node2162;
	wire [4-1:0] node2163;
	wire [4-1:0] node2168;
	wire [4-1:0] node2170;
	wire [4-1:0] node2172;
	wire [4-1:0] node2173;
	wire [4-1:0] node2177;
	wire [4-1:0] node2178;
	wire [4-1:0] node2180;
	wire [4-1:0] node2181;
	wire [4-1:0] node2182;
	wire [4-1:0] node2187;
	wire [4-1:0] node2188;
	wire [4-1:0] node2189;
	wire [4-1:0] node2190;
	wire [4-1:0] node2192;
	wire [4-1:0] node2196;
	wire [4-1:0] node2197;
	wire [4-1:0] node2201;
	wire [4-1:0] node2202;
	wire [4-1:0] node2204;
	wire [4-1:0] node2205;
	wire [4-1:0] node2209;
	wire [4-1:0] node2210;
	wire [4-1:0] node2214;
	wire [4-1:0] node2216;
	wire [4-1:0] node2217;
	wire [4-1:0] node2218;
	wire [4-1:0] node2219;
	wire [4-1:0] node2221;
	wire [4-1:0] node2224;
	wire [4-1:0] node2225;
	wire [4-1:0] node2226;
	wire [4-1:0] node2230;
	wire [4-1:0] node2231;
	wire [4-1:0] node2235;
	wire [4-1:0] node2236;
	wire [4-1:0] node2237;
	wire [4-1:0] node2239;
	wire [4-1:0] node2242;
	wire [4-1:0] node2245;
	wire [4-1:0] node2246;
	wire [4-1:0] node2248;
	wire [4-1:0] node2251;
	wire [4-1:0] node2252;
	wire [4-1:0] node2256;
	wire [4-1:0] node2258;
	wire [4-1:0] node2259;
	wire [4-1:0] node2260;
	wire [4-1:0] node2261;
	wire [4-1:0] node2266;
	wire [4-1:0] node2267;

	assign outp = (inp[14]) ? node2 : 4'b0000;
		assign node2 = (inp[12]) ? node1380 : node3;
			assign node3 = (inp[3]) ? node383 : node4;
				assign node4 = (inp[0]) ? node148 : node5;
					assign node5 = (inp[4]) ? 4'b0000 : node6;
						assign node6 = (inp[11]) ? node72 : node7;
							assign node7 = (inp[7]) ? 4'b0010 : node8;
								assign node8 = (inp[9]) ? node38 : node9;
									assign node9 = (inp[5]) ? 4'b0000 : node10;
										assign node10 = (inp[15]) ? node22 : node11;
											assign node11 = (inp[13]) ? 4'b0010 : node12;
												assign node12 = (inp[8]) ? node14 : 4'b0010;
													assign node14 = (inp[1]) ? node16 : 4'b0000;
														assign node16 = (inp[6]) ? 4'b0010 : node17;
															assign node17 = (inp[10]) ? 4'b0000 : 4'b0010;
											assign node22 = (inp[13]) ? node24 : 4'b0000;
												assign node24 = (inp[1]) ? node30 : node25;
													assign node25 = (inp[8]) ? 4'b0000 : node26;
														assign node26 = (inp[6]) ? 4'b0010 : 4'b0000;
													assign node30 = (inp[10]) ? node32 : 4'b0010;
														assign node32 = (inp[8]) ? node34 : 4'b0010;
															assign node34 = (inp[6]) ? 4'b0010 : 4'b0000;
									assign node38 = (inp[5]) ? node40 : 4'b0010;
										assign node40 = (inp[15]) ? node56 : node41;
											assign node41 = (inp[13]) ? 4'b0010 : node42;
												assign node42 = (inp[10]) ? node48 : node43;
													assign node43 = (inp[8]) ? node45 : 4'b0010;
														assign node45 = (inp[1]) ? 4'b0010 : 4'b0000;
													assign node48 = (inp[6]) ? node50 : 4'b0000;
														assign node50 = (inp[8]) ? node52 : 4'b0010;
															assign node52 = (inp[2]) ? 4'b0010 : 4'b0000;
											assign node56 = (inp[13]) ? node58 : 4'b0000;
												assign node58 = (inp[1]) ? node64 : node59;
													assign node59 = (inp[8]) ? 4'b0000 : node60;
														assign node60 = (inp[6]) ? 4'b0010 : 4'b0000;
													assign node64 = (inp[10]) ? node66 : 4'b0010;
														assign node66 = (inp[6]) ? 4'b0010 : node67;
															assign node67 = (inp[8]) ? 4'b0000 : 4'b0010;
							assign node72 = (inp[7]) ? node74 : 4'b0000;
								assign node74 = (inp[9]) ? node112 : node75;
									assign node75 = (inp[5]) ? 4'b0000 : node76;
										assign node76 = (inp[13]) ? node94 : node77;
											assign node77 = (inp[15]) ? 4'b0000 : node78;
												assign node78 = (inp[8]) ? node86 : node79;
													assign node79 = (inp[1]) ? 4'b0010 : node80;
														assign node80 = (inp[10]) ? node82 : 4'b0010;
															assign node82 = (inp[2]) ? 4'b0010 : 4'b0000;
													assign node86 = (inp[1]) ? node88 : 4'b0000;
														assign node88 = (inp[6]) ? 4'b0010 : node89;
															assign node89 = (inp[10]) ? 4'b0000 : 4'b0010;
											assign node94 = (inp[15]) ? node96 : 4'b0010;
												assign node96 = (inp[1]) ? node104 : node97;
													assign node97 = (inp[8]) ? 4'b0000 : node98;
														assign node98 = (inp[10]) ? node100 : 4'b0010;
															assign node100 = (inp[2]) ? 4'b0000 : 4'b0010;
													assign node104 = (inp[10]) ? node106 : 4'b0010;
														assign node106 = (inp[6]) ? 4'b0010 : node107;
															assign node107 = (inp[8]) ? 4'b0000 : 4'b0010;
									assign node112 = (inp[5]) ? node114 : 4'b0010;
										assign node114 = (inp[15]) ? node132 : node115;
											assign node115 = (inp[13]) ? 4'b0010 : node116;
												assign node116 = (inp[8]) ? node124 : node117;
													assign node117 = (inp[6]) ? 4'b0010 : node118;
														assign node118 = (inp[1]) ? 4'b0010 : node119;
															assign node119 = (inp[2]) ? 4'b0000 : 4'b0010;
													assign node124 = (inp[1]) ? node126 : 4'b0000;
														assign node126 = (inp[6]) ? 4'b0010 : node127;
															assign node127 = (inp[10]) ? 4'b0000 : 4'b0010;
											assign node132 = (inp[13]) ? node134 : 4'b0000;
												assign node134 = (inp[8]) ? node142 : node135;
													assign node135 = (inp[1]) ? 4'b0010 : node136;
														assign node136 = (inp[6]) ? 4'b0010 : node137;
															assign node137 = (inp[10]) ? 4'b0000 : 4'b0010;
													assign node142 = (inp[1]) ? node144 : 4'b0000;
														assign node144 = (inp[10]) ? 4'b0000 : 4'b0010;
					assign node148 = (inp[4]) ? node306 : node149;
						assign node149 = (inp[7]) ? node221 : node150;
							assign node150 = (inp[11]) ? node186 : node151;
								assign node151 = (inp[9]) ? 4'b0000 : node152;
									assign node152 = (inp[5]) ? node168 : node153;
										assign node153 = (inp[13]) ? 4'b0000 : node154;
											assign node154 = (inp[15]) ? node162 : node155;
												assign node155 = (inp[6]) ? 4'b0000 : node156;
													assign node156 = (inp[8]) ? node158 : 4'b0000;
														assign node158 = (inp[1]) ? 4'b0000 : 4'b0010;
												assign node162 = (inp[1]) ? node164 : 4'b0010;
													assign node164 = (inp[8]) ? 4'b0010 : 4'b0000;
										assign node168 = (inp[13]) ? node170 : 4'b0010;
											assign node170 = (inp[1]) ? node178 : node171;
												assign node171 = (inp[15]) ? 4'b0010 : node172;
													assign node172 = (inp[6]) ? 4'b0000 : node173;
														assign node173 = (inp[8]) ? 4'b0010 : 4'b0000;
												assign node178 = (inp[6]) ? 4'b0000 : node179;
													assign node179 = (inp[15]) ? node181 : 4'b0000;
														assign node181 = (inp[8]) ? 4'b0010 : 4'b0000;
								assign node186 = (inp[9]) ? node188 : 4'b0010;
									assign node188 = (inp[13]) ? node206 : node189;
										assign node189 = (inp[5]) ? 4'b0010 : node190;
											assign node190 = (inp[15]) ? node198 : node191;
												assign node191 = (inp[8]) ? node193 : 4'b0000;
													assign node193 = (inp[6]) ? 4'b0000 : node194;
														assign node194 = (inp[1]) ? 4'b0000 : 4'b0010;
												assign node198 = (inp[1]) ? node200 : 4'b0010;
													assign node200 = (inp[6]) ? 4'b0000 : node201;
														assign node201 = (inp[8]) ? 4'b0010 : 4'b0000;
										assign node206 = (inp[5]) ? node208 : 4'b0000;
											assign node208 = (inp[1]) ? node214 : node209;
												assign node209 = (inp[15]) ? 4'b0010 : node210;
													assign node210 = (inp[8]) ? 4'b0010 : 4'b0000;
												assign node214 = (inp[15]) ? node216 : 4'b0000;
													assign node216 = (inp[8]) ? node218 : 4'b0000;
														assign node218 = (inp[6]) ? 4'b0000 : 4'b0010;
							assign node221 = (inp[9]) ? node245 : node222;
								assign node222 = (inp[11]) ? 4'b0000 : node223;
									assign node223 = (inp[13]) ? node225 : 4'b0000;
										assign node225 = (inp[5]) ? 4'b0000 : node226;
											assign node226 = (inp[1]) ? node234 : node227;
												assign node227 = (inp[6]) ? node229 : 4'b0000;
													assign node229 = (inp[15]) ? 4'b0000 : node230;
														assign node230 = (inp[8]) ? 4'b0000 : 4'b0010;
												assign node234 = (inp[6]) ? 4'b0010 : node235;
													assign node235 = (inp[15]) ? node237 : 4'b0010;
														assign node237 = (inp[8]) ? 4'b0000 : node238;
															assign node238 = (inp[10]) ? 4'b0000 : 4'b0010;
								assign node245 = (inp[11]) ? node265 : node246;
									assign node246 = (inp[5]) ? node248 : 4'b0010;
										assign node248 = (inp[1]) ? 4'b0010 : node249;
											assign node249 = (inp[13]) ? 4'b0010 : node250;
												assign node250 = (inp[15]) ? node258 : node251;
													assign node251 = (inp[10]) ? node253 : 4'b0010;
														assign node253 = (inp[8]) ? node255 : 4'b0010;
															assign node255 = (inp[6]) ? 4'b0010 : 4'b0000;
													assign node258 = (inp[6]) ? node260 : 4'b0000;
														assign node260 = (inp[8]) ? 4'b0000 : 4'b0010;
									assign node265 = (inp[13]) ? node279 : node266;
										assign node266 = (inp[5]) ? 4'b0000 : node267;
											assign node267 = (inp[1]) ? node269 : 4'b0000;
												assign node269 = (inp[15]) ? 4'b0000 : node270;
													assign node270 = (inp[6]) ? 4'b0010 : node271;
														assign node271 = (inp[8]) ? 4'b0000 : node272;
															assign node272 = (inp[2]) ? 4'b0000 : 4'b0010;
										assign node279 = (inp[5]) ? node289 : node280;
											assign node280 = (inp[2]) ? node282 : 4'b0010;
												assign node282 = (inp[10]) ? node284 : 4'b0010;
													assign node284 = (inp[8]) ? node286 : 4'b0010;
														assign node286 = (inp[6]) ? 4'b0010 : 4'b0000;
											assign node289 = (inp[1]) ? node297 : node290;
												assign node290 = (inp[8]) ? 4'b0000 : node291;
													assign node291 = (inp[6]) ? node293 : 4'b0000;
														assign node293 = (inp[15]) ? 4'b0000 : 4'b0010;
												assign node297 = (inp[15]) ? node299 : 4'b0010;
													assign node299 = (inp[6]) ? 4'b0010 : node300;
														assign node300 = (inp[10]) ? 4'b0000 : node301;
															assign node301 = (inp[8]) ? 4'b0000 : 4'b0010;
						assign node306 = (inp[7]) ? node308 : 4'b0010;
							assign node308 = (inp[11]) ? node346 : node309;
								assign node309 = (inp[9]) ? 4'b0000 : node310;
									assign node310 = (inp[13]) ? node328 : node311;
										assign node311 = (inp[5]) ? 4'b0010 : node312;
											assign node312 = (inp[15]) ? node320 : node313;
												assign node313 = (inp[1]) ? 4'b0000 : node314;
													assign node314 = (inp[6]) ? 4'b0000 : node315;
														assign node315 = (inp[10]) ? 4'b0000 : 4'b0010;
												assign node320 = (inp[1]) ? node322 : 4'b0010;
													assign node322 = (inp[8]) ? node324 : 4'b0000;
														assign node324 = (inp[6]) ? 4'b0000 : 4'b0010;
										assign node328 = (inp[5]) ? node330 : 4'b0000;
											assign node330 = (inp[15]) ? node338 : node331;
												assign node331 = (inp[6]) ? 4'b0000 : node332;
													assign node332 = (inp[8]) ? node334 : 4'b0000;
														assign node334 = (inp[1]) ? 4'b0000 : 4'b0010;
												assign node338 = (inp[1]) ? node340 : 4'b0010;
													assign node340 = (inp[6]) ? 4'b0000 : node341;
														assign node341 = (inp[8]) ? 4'b0010 : 4'b0000;
								assign node346 = (inp[9]) ? node348 : 4'b0010;
									assign node348 = (inp[5]) ? node366 : node349;
										assign node349 = (inp[13]) ? 4'b0000 : node350;
											assign node350 = (inp[15]) ? node358 : node351;
												assign node351 = (inp[6]) ? 4'b0000 : node352;
													assign node352 = (inp[1]) ? 4'b0000 : node353;
														assign node353 = (inp[8]) ? 4'b0010 : 4'b0000;
												assign node358 = (inp[1]) ? node360 : 4'b0010;
													assign node360 = (inp[8]) ? node362 : 4'b0000;
														assign node362 = (inp[6]) ? 4'b0000 : 4'b0010;
										assign node366 = (inp[13]) ? node368 : 4'b0010;
											assign node368 = (inp[1]) ? node376 : node369;
												assign node369 = (inp[15]) ? 4'b0010 : node370;
													assign node370 = (inp[6]) ? 4'b0000 : node371;
														assign node371 = (inp[8]) ? 4'b0010 : 4'b0000;
												assign node376 = (inp[6]) ? 4'b0000 : node377;
													assign node377 = (inp[15]) ? node379 : 4'b0000;
														assign node379 = (inp[8]) ? 4'b0010 : 4'b0000;
				assign node383 = (inp[0]) ? node519 : node384;
					assign node384 = (inp[4]) ? node386 : 4'b0010;
						assign node386 = (inp[11]) ? node452 : node387;
							assign node387 = (inp[7]) ? 4'b0010 : node388;
								assign node388 = (inp[5]) ? node420 : node389;
									assign node389 = (inp[9]) ? 4'b0010 : node390;
										assign node390 = (inp[15]) ? node402 : node391;
											assign node391 = (inp[13]) ? 4'b0010 : node392;
												assign node392 = (inp[1]) ? 4'b0010 : node393;
													assign node393 = (inp[8]) ? 4'b0000 : node394;
														assign node394 = (inp[6]) ? 4'b0010 : node395;
															assign node395 = (inp[10]) ? 4'b0000 : 4'b0010;
											assign node402 = (inp[13]) ? node404 : 4'b0000;
												assign node404 = (inp[1]) ? node412 : node405;
													assign node405 = (inp[8]) ? 4'b0000 : node406;
														assign node406 = (inp[10]) ? node408 : 4'b0010;
															assign node408 = (inp[6]) ? 4'b0010 : 4'b0000;
													assign node412 = (inp[6]) ? 4'b0010 : node413;
														assign node413 = (inp[10]) ? node415 : 4'b0010;
															assign node415 = (inp[8]) ? 4'b0000 : 4'b0010;
									assign node420 = (inp[9]) ? node422 : 4'b0000;
										assign node422 = (inp[13]) ? node436 : node423;
											assign node423 = (inp[15]) ? 4'b0000 : node424;
												assign node424 = (inp[1]) ? node430 : node425;
													assign node425 = (inp[8]) ? 4'b0000 : node426;
														assign node426 = (inp[10]) ? 4'b0000 : 4'b0010;
													assign node430 = (inp[10]) ? node432 : 4'b0010;
														assign node432 = (inp[6]) ? 4'b0010 : 4'b0000;
											assign node436 = (inp[15]) ? node438 : 4'b0010;
												assign node438 = (inp[8]) ? node444 : node439;
													assign node439 = (inp[6]) ? 4'b0010 : node440;
														assign node440 = (inp[10]) ? 4'b0000 : 4'b0010;
													assign node444 = (inp[1]) ? node446 : 4'b0000;
														assign node446 = (inp[6]) ? 4'b0010 : node447;
															assign node447 = (inp[10]) ? 4'b0000 : 4'b0010;
							assign node452 = (inp[7]) ? node454 : 4'b0000;
								assign node454 = (inp[9]) ? node480 : node455;
									assign node455 = (inp[5]) ? 4'b0000 : node456;
										assign node456 = (inp[15]) ? node466 : node457;
											assign node457 = (inp[13]) ? 4'b0010 : node458;
												assign node458 = (inp[1]) ? 4'b0010 : node459;
													assign node459 = (inp[8]) ? 4'b0000 : node460;
														assign node460 = (inp[6]) ? 4'b0010 : 4'b0000;
											assign node466 = (inp[13]) ? node468 : 4'b0000;
												assign node468 = (inp[8]) ? node474 : node469;
													assign node469 = (inp[10]) ? node471 : 4'b0010;
														assign node471 = (inp[6]) ? 4'b0010 : 4'b0000;
													assign node474 = (inp[1]) ? node476 : 4'b0000;
														assign node476 = (inp[6]) ? 4'b0010 : 4'b0000;
									assign node480 = (inp[5]) ? node482 : 4'b0010;
										assign node482 = (inp[13]) ? node500 : node483;
											assign node483 = (inp[15]) ? 4'b0000 : node484;
												assign node484 = (inp[8]) ? node492 : node485;
													assign node485 = (inp[6]) ? 4'b0010 : node486;
														assign node486 = (inp[2]) ? 4'b0010 : node487;
															assign node487 = (inp[1]) ? 4'b0010 : 4'b0000;
													assign node492 = (inp[1]) ? node494 : 4'b0000;
														assign node494 = (inp[10]) ? node496 : 4'b0010;
															assign node496 = (inp[6]) ? 4'b0010 : 4'b0000;
											assign node500 = (inp[15]) ? node502 : 4'b0010;
												assign node502 = (inp[10]) ? node508 : node503;
													assign node503 = (inp[8]) ? node505 : 4'b0010;
														assign node505 = (inp[1]) ? 4'b0010 : 4'b0000;
													assign node508 = (inp[1]) ? node514 : node509;
														assign node509 = (inp[8]) ? 4'b0000 : node510;
															assign node510 = (inp[2]) ? 4'b0010 : 4'b0000;
														assign node514 = (inp[2]) ? node516 : 4'b0010;
															assign node516 = (inp[6]) ? 4'b0010 : 4'b0000;
					assign node519 = (inp[9]) ? node921 : node520;
						assign node520 = (inp[7]) ? node624 : node521;
							assign node521 = (inp[4]) ? node565 : node522;
								assign node522 = (inp[11]) ? node548 : node523;
									assign node523 = (inp[13]) ? node539 : node524;
										assign node524 = (inp[1]) ? node532 : node525;
											assign node525 = (inp[5]) ? 4'b0010 : node526;
												assign node526 = (inp[6]) ? 4'b1000 : node527;
													assign node527 = (inp[15]) ? 4'b0010 : 4'b1000;
											assign node532 = (inp[5]) ? node534 : 4'b1000;
												assign node534 = (inp[15]) ? node536 : 4'b1000;
													assign node536 = (inp[6]) ? 4'b1000 : 4'b0010;
										assign node539 = (inp[5]) ? 4'b1000 : node540;
											assign node540 = (inp[1]) ? node542 : 4'b1000;
												assign node542 = (inp[6]) ? 4'b1010 : node543;
													assign node543 = (inp[15]) ? 4'b1000 : 4'b1010;
									assign node548 = (inp[13]) ? node550 : 4'b0010;
										assign node550 = (inp[1]) ? node558 : node551;
											assign node551 = (inp[5]) ? 4'b0010 : node552;
												assign node552 = (inp[15]) ? node554 : 4'b1000;
													assign node554 = (inp[6]) ? 4'b1000 : 4'b0010;
											assign node558 = (inp[5]) ? node560 : 4'b1000;
												assign node560 = (inp[15]) ? node562 : 4'b1000;
													assign node562 = (inp[6]) ? 4'b1000 : 4'b0010;
								assign node565 = (inp[11]) ? node603 : node566;
									assign node566 = (inp[13]) ? node592 : node567;
										assign node567 = (inp[5]) ? node583 : node568;
											assign node568 = (inp[1]) ? 4'b0010 : node569;
												assign node569 = (inp[15]) ? node577 : node570;
													assign node570 = (inp[10]) ? node572 : 4'b0010;
														assign node572 = (inp[8]) ? node574 : 4'b0010;
															assign node574 = (inp[2]) ? 4'b0000 : 4'b0010;
													assign node577 = (inp[8]) ? 4'b0000 : node578;
														assign node578 = (inp[6]) ? 4'b0010 : 4'b0000;
											assign node583 = (inp[1]) ? node585 : 4'b0000;
												assign node585 = (inp[15]) ? 4'b0000 : node586;
													assign node586 = (inp[6]) ? 4'b0010 : node587;
														assign node587 = (inp[8]) ? 4'b0000 : 4'b0010;
										assign node592 = (inp[10]) ? node594 : 4'b0010;
											assign node594 = (inp[6]) ? 4'b0010 : node595;
												assign node595 = (inp[1]) ? 4'b0010 : node596;
													assign node596 = (inp[5]) ? node598 : 4'b0010;
														assign node598 = (inp[15]) ? 4'b0000 : 4'b0010;
									assign node603 = (inp[13]) ? node605 : 4'b0000;
										assign node605 = (inp[1]) ? node615 : node606;
											assign node606 = (inp[15]) ? 4'b0000 : node607;
												assign node607 = (inp[6]) ? node609 : 4'b0000;
													assign node609 = (inp[5]) ? 4'b0000 : node610;
														assign node610 = (inp[8]) ? 4'b0000 : 4'b0010;
											assign node615 = (inp[5]) ? 4'b0000 : node616;
												assign node616 = (inp[15]) ? node618 : 4'b0010;
													assign node618 = (inp[6]) ? 4'b0010 : node619;
														assign node619 = (inp[8]) ? 4'b0000 : 4'b0010;
							assign node624 = (inp[13]) ? node802 : node625;
								assign node625 = (inp[4]) ? node677 : node626;
									assign node626 = (inp[11]) ? node650 : node627;
										assign node627 = (inp[6]) ? node639 : node628;
											assign node628 = (inp[1]) ? node632 : node629;
												assign node629 = (inp[5]) ? 4'b1010 : 4'b0000;
												assign node632 = (inp[5]) ? node634 : 4'b0010;
													assign node634 = (inp[15]) ? 4'b0000 : node635;
														assign node635 = (inp[10]) ? 4'b0000 : 4'b0010;
											assign node639 = (inp[1]) ? node647 : node640;
												assign node640 = (inp[15]) ? 4'b0000 : node641;
													assign node641 = (inp[5]) ? 4'b0000 : node642;
														assign node642 = (inp[8]) ? 4'b0000 : 4'b0010;
												assign node647 = (inp[5]) ? 4'b0010 : 4'b0000;
										assign node650 = (inp[1]) ? node668 : node651;
											assign node651 = (inp[5]) ? node661 : node652;
												assign node652 = (inp[10]) ? node654 : 4'b1010;
													assign node654 = (inp[8]) ? node656 : 4'b1010;
														assign node656 = (inp[6]) ? 4'b1010 : node657;
															assign node657 = (inp[15]) ? 4'b1000 : 4'b1010;
												assign node661 = (inp[6]) ? node663 : 4'b1000;
													assign node663 = (inp[8]) ? node665 : 4'b1010;
														assign node665 = (inp[15]) ? 4'b1000 : 4'b1010;
											assign node668 = (inp[6]) ? node672 : node669;
												assign node669 = (inp[5]) ? 4'b1010 : 4'b0000;
												assign node672 = (inp[15]) ? 4'b0000 : node673;
													assign node673 = (inp[5]) ? 4'b0000 : 4'b0010;
									assign node677 = (inp[15]) ? node705 : node678;
										assign node678 = (inp[1]) ? node692 : node679;
											assign node679 = (inp[11]) ? node685 : node680;
												assign node680 = (inp[5]) ? node682 : 4'b1000;
													assign node682 = (inp[6]) ? 4'b1000 : 4'b1010;
												assign node685 = (inp[5]) ? node687 : 4'b1010;
													assign node687 = (inp[6]) ? node689 : 4'b1000;
														assign node689 = (inp[8]) ? 4'b1000 : 4'b1010;
											assign node692 = (inp[11]) ? node698 : node693;
												assign node693 = (inp[5]) ? node695 : 4'b1010;
													assign node695 = (inp[6]) ? 4'b1010 : 4'b1000;
												assign node698 = (inp[5]) ? 4'b1010 : node699;
													assign node699 = (inp[8]) ? node701 : 4'b1000;
														assign node701 = (inp[6]) ? 4'b1000 : 4'b1010;
										assign node705 = (inp[10]) ? node763 : node706;
											assign node706 = (inp[8]) ? node736 : node707;
												assign node707 = (inp[6]) ? node723 : node708;
													assign node708 = (inp[1]) ? node716 : node709;
														assign node709 = (inp[11]) ? node713 : node710;
															assign node710 = (inp[5]) ? 4'b1010 : 4'b1000;
															assign node713 = (inp[5]) ? 4'b1000 : 4'b1010;
														assign node716 = (inp[2]) ? 4'b1010 : node717;
															assign node717 = (inp[5]) ? node719 : 4'b1010;
																assign node719 = (inp[11]) ? 4'b1010 : 4'b1000;
													assign node723 = (inp[11]) ? node729 : node724;
														assign node724 = (inp[5]) ? node726 : 4'b1000;
															assign node726 = (inp[1]) ? 4'b1000 : 4'b1010;
														assign node729 = (inp[5]) ? node733 : node730;
															assign node730 = (inp[1]) ? 4'b1000 : 4'b1010;
															assign node733 = (inp[1]) ? 4'b1010 : 4'b1000;
												assign node736 = (inp[6]) ? node748 : node737;
													assign node737 = (inp[5]) ? node745 : node738;
														assign node738 = (inp[2]) ? 4'b1000 : node739;
															assign node739 = (inp[1]) ? node741 : 4'b1010;
																assign node741 = (inp[11]) ? 4'b1010 : 4'b1000;
														assign node745 = (inp[2]) ? 4'b1010 : 4'b1000;
													assign node748 = (inp[1]) ? node756 : node749;
														assign node749 = (inp[2]) ? node751 : 4'b1000;
															assign node751 = (inp[5]) ? 4'b1000 : node752;
																assign node752 = (inp[11]) ? 4'b1010 : 4'b1000;
														assign node756 = (inp[2]) ? node758 : 4'b1010;
															assign node758 = (inp[11]) ? 4'b1000 : node759;
																assign node759 = (inp[5]) ? 4'b1000 : 4'b1010;
											assign node763 = (inp[1]) ? node787 : node764;
												assign node764 = (inp[8]) ? node776 : node765;
													assign node765 = (inp[6]) ? node767 : 4'b1000;
														assign node767 = (inp[2]) ? node773 : node768;
															assign node768 = (inp[11]) ? node770 : 4'b1010;
																assign node770 = (inp[5]) ? 4'b1000 : 4'b1010;
															assign node773 = (inp[5]) ? 4'b1010 : 4'b1000;
													assign node776 = (inp[2]) ? node778 : 4'b1010;
														assign node778 = (inp[6]) ? node782 : node779;
															assign node779 = (inp[11]) ? 4'b1000 : 4'b1010;
															assign node782 = (inp[5]) ? 4'b1000 : node783;
																assign node783 = (inp[11]) ? 4'b1010 : 4'b1000;
												assign node787 = (inp[11]) ? node793 : node788;
													assign node788 = (inp[6]) ? node790 : 4'b1000;
														assign node790 = (inp[5]) ? 4'b1000 : 4'b1010;
													assign node793 = (inp[5]) ? node797 : node794;
														assign node794 = (inp[6]) ? 4'b1000 : 4'b1010;
														assign node797 = (inp[6]) ? 4'b1010 : node798;
															assign node798 = (inp[8]) ? 4'b1000 : 4'b1010;
								assign node802 = (inp[5]) ? node872 : node803;
									assign node803 = (inp[6]) ? node851 : node804;
										assign node804 = (inp[4]) ? node834 : node805;
											assign node805 = (inp[1]) ? node825 : node806;
												assign node806 = (inp[10]) ? node814 : node807;
													assign node807 = (inp[15]) ? 4'b0010 : node808;
														assign node808 = (inp[8]) ? 4'b0010 : node809;
															assign node809 = (inp[11]) ? 4'b0000 : 4'b0010;
													assign node814 = (inp[8]) ? node820 : node815;
														assign node815 = (inp[11]) ? node817 : 4'b0010;
															assign node817 = (inp[2]) ? 4'b0010 : 4'b0000;
														assign node820 = (inp[11]) ? 4'b0010 : node821;
															assign node821 = (inp[15]) ? 4'b0000 : 4'b0010;
												assign node825 = (inp[15]) ? node831 : node826;
													assign node826 = (inp[11]) ? 4'b1000 : node827;
														assign node827 = (inp[8]) ? 4'b1010 : 4'b1000;
													assign node831 = (inp[11]) ? 4'b0010 : 4'b1010;
											assign node834 = (inp[1]) ? node844 : node835;
												assign node835 = (inp[11]) ? node837 : 4'b0000;
													assign node837 = (inp[15]) ? 4'b1000 : node838;
														assign node838 = (inp[8]) ? node840 : 4'b1010;
															assign node840 = (inp[10]) ? 4'b1000 : 4'b1010;
												assign node844 = (inp[8]) ? node846 : 4'b0000;
													assign node846 = (inp[15]) ? node848 : 4'b0000;
														assign node848 = (inp[11]) ? 4'b0000 : 4'b0010;
										assign node851 = (inp[4]) ? node861 : node852;
											assign node852 = (inp[1]) ? 4'b1010 : node853;
												assign node853 = (inp[11]) ? node855 : 4'b1000;
													assign node855 = (inp[8]) ? 4'b0000 : node856;
														assign node856 = (inp[15]) ? 4'b0000 : 4'b0010;
											assign node861 = (inp[11]) ? node869 : node862;
												assign node862 = (inp[8]) ? node864 : 4'b0010;
													assign node864 = (inp[1]) ? 4'b0010 : node865;
														assign node865 = (inp[15]) ? 4'b0000 : 4'b0010;
												assign node869 = (inp[1]) ? 4'b0010 : 4'b1010;
									assign node872 = (inp[6]) ? node904 : node873;
										assign node873 = (inp[4]) ? node887 : node874;
											assign node874 = (inp[11]) ? node880 : node875;
												assign node875 = (inp[1]) ? node877 : 4'b0000;
													assign node877 = (inp[15]) ? 4'b1000 : 4'b1010;
												assign node880 = (inp[15]) ? node882 : 4'b0010;
													assign node882 = (inp[10]) ? 4'b0000 : node883;
														assign node883 = (inp[8]) ? 4'b0000 : 4'b0010;
											assign node887 = (inp[11]) ? node897 : node888;
												assign node888 = (inp[1]) ? node890 : 4'b1010;
													assign node890 = (inp[10]) ? node892 : 4'b0010;
														assign node892 = (inp[15]) ? node894 : 4'b0010;
															assign node894 = (inp[8]) ? 4'b0000 : 4'b0010;
												assign node897 = (inp[1]) ? 4'b1010 : node898;
													assign node898 = (inp[8]) ? node900 : 4'b1000;
														assign node900 = (inp[15]) ? 4'b1010 : 4'b1000;
										assign node904 = (inp[1]) ? node918 : node905;
											assign node905 = (inp[4]) ? node911 : node906;
												assign node906 = (inp[15]) ? 4'b0010 : node907;
													assign node907 = (inp[11]) ? 4'b0000 : 4'b0010;
												assign node911 = (inp[11]) ? node913 : 4'b0000;
													assign node913 = (inp[8]) ? 4'b1000 : node914;
														assign node914 = (inp[15]) ? 4'b1000 : 4'b1010;
											assign node918 = (inp[4]) ? 4'b0000 : 4'b1000;
						assign node921 = (inp[7]) ? node1099 : node922;
							assign node922 = (inp[4]) ? node1026 : node923;
								assign node923 = (inp[11]) ? node985 : node924;
									assign node924 = (inp[13]) ? node942 : node925;
										assign node925 = (inp[1]) ? node933 : node926;
											assign node926 = (inp[5]) ? node928 : 4'b1010;
												assign node928 = (inp[15]) ? node930 : 4'b1010;
													assign node930 = (inp[6]) ? 4'b1010 : 4'b1000;
											assign node933 = (inp[5]) ? 4'b1010 : node934;
												assign node934 = (inp[6]) ? 4'b1000 : node935;
													assign node935 = (inp[8]) ? 4'b1010 : node936;
														assign node936 = (inp[15]) ? 4'b1010 : 4'b1000;
										assign node942 = (inp[1]) ? node974 : node943;
											assign node943 = (inp[2]) ? node959 : node944;
												assign node944 = (inp[15]) ? node952 : node945;
													assign node945 = (inp[6]) ? node947 : 4'b1000;
														assign node947 = (inp[8]) ? 4'b1000 : node948;
															assign node948 = (inp[5]) ? 4'b1000 : 4'b1010;
													assign node952 = (inp[6]) ? 4'b1000 : node953;
														assign node953 = (inp[8]) ? node955 : 4'b1000;
															assign node955 = (inp[5]) ? 4'b1010 : 4'b1000;
												assign node959 = (inp[8]) ? node967 : node960;
													assign node960 = (inp[6]) ? node962 : 4'b1000;
														assign node962 = (inp[5]) ? 4'b1000 : node963;
															assign node963 = (inp[15]) ? 4'b1000 : 4'b1010;
													assign node967 = (inp[5]) ? node969 : 4'b1000;
														assign node969 = (inp[15]) ? node971 : 4'b1000;
															assign node971 = (inp[6]) ? 4'b1000 : 4'b1010;
											assign node974 = (inp[6]) ? 4'b1010 : node975;
												assign node975 = (inp[5]) ? node977 : 4'b1010;
													assign node977 = (inp[15]) ? 4'b1000 : node978;
														assign node978 = (inp[10]) ? 4'b1000 : node979;
															assign node979 = (inp[8]) ? 4'b1000 : 4'b1010;
									assign node985 = (inp[13]) ? node1009 : node986;
										assign node986 = (inp[1]) ? node996 : node987;
											assign node987 = (inp[6]) ? node989 : 4'b1000;
												assign node989 = (inp[5]) ? 4'b1000 : node990;
													assign node990 = (inp[15]) ? 4'b1000 : node991;
														assign node991 = (inp[8]) ? 4'b1000 : 4'b1010;
											assign node996 = (inp[5]) ? node1004 : node997;
												assign node997 = (inp[8]) ? node999 : 4'b1010;
													assign node999 = (inp[6]) ? 4'b1010 : node1000;
														assign node1000 = (inp[15]) ? 4'b1000 : 4'b1010;
												assign node1004 = (inp[6]) ? node1006 : 4'b1000;
													assign node1006 = (inp[15]) ? 4'b1000 : 4'b1010;
										assign node1009 = (inp[1]) ? node1017 : node1010;
											assign node1010 = (inp[6]) ? node1012 : 4'b1010;
												assign node1012 = (inp[5]) ? 4'b1010 : node1013;
													assign node1013 = (inp[15]) ? 4'b1010 : 4'b1000;
											assign node1017 = (inp[6]) ? 4'b1000 : node1018;
												assign node1018 = (inp[5]) ? node1020 : 4'b1000;
													assign node1020 = (inp[15]) ? 4'b1010 : node1021;
														assign node1021 = (inp[8]) ? 4'b1010 : 4'b1000;
								assign node1026 = (inp[11]) ? node1068 : node1027;
									assign node1027 = (inp[13]) ? node1043 : node1028;
										assign node1028 = (inp[5]) ? node1036 : node1029;
											assign node1029 = (inp[6]) ? 4'b1000 : node1030;
												assign node1030 = (inp[1]) ? 4'b1000 : node1031;
													assign node1031 = (inp[15]) ? 4'b0010 : 4'b1000;
											assign node1036 = (inp[1]) ? node1038 : 4'b0010;
												assign node1038 = (inp[6]) ? 4'b1000 : node1039;
													assign node1039 = (inp[15]) ? 4'b0010 : 4'b1000;
										assign node1043 = (inp[1]) ? node1059 : node1044;
											assign node1044 = (inp[5]) ? 4'b1000 : node1045;
												assign node1045 = (inp[6]) ? node1053 : node1046;
													assign node1046 = (inp[15]) ? 4'b1000 : node1047;
														assign node1047 = (inp[10]) ? 4'b1000 : node1048;
															assign node1048 = (inp[8]) ? 4'b1000 : 4'b1010;
													assign node1053 = (inp[8]) ? node1055 : 4'b1010;
														assign node1055 = (inp[15]) ? 4'b1000 : 4'b1010;
											assign node1059 = (inp[5]) ? node1061 : 4'b1010;
												assign node1061 = (inp[6]) ? 4'b1010 : node1062;
													assign node1062 = (inp[15]) ? 4'b1000 : node1063;
														assign node1063 = (inp[10]) ? 4'b1000 : 4'b1010;
									assign node1068 = (inp[13]) ? node1084 : node1069;
										assign node1069 = (inp[1]) ? 4'b0010 : node1070;
											assign node1070 = (inp[5]) ? node1072 : 4'b0010;
												assign node1072 = (inp[6]) ? node1078 : node1073;
													assign node1073 = (inp[15]) ? 4'b0000 : node1074;
														assign node1074 = (inp[8]) ? 4'b0000 : 4'b0010;
													assign node1078 = (inp[15]) ? node1080 : 4'b0010;
														assign node1080 = (inp[8]) ? 4'b0000 : 4'b0010;
										assign node1084 = (inp[5]) ? node1092 : node1085;
											assign node1085 = (inp[15]) ? node1087 : 4'b1000;
												assign node1087 = (inp[6]) ? 4'b1000 : node1088;
													assign node1088 = (inp[1]) ? 4'b1000 : 4'b0010;
											assign node1092 = (inp[1]) ? node1094 : 4'b0010;
												assign node1094 = (inp[15]) ? node1096 : 4'b1000;
													assign node1096 = (inp[6]) ? 4'b1000 : 4'b0010;
							assign node1099 = (inp[13]) ? node1269 : node1100;
								assign node1100 = (inp[4]) ? node1176 : node1101;
									assign node1101 = (inp[15]) ? node1141 : node1102;
										assign node1102 = (inp[6]) ? node1126 : node1103;
											assign node1103 = (inp[11]) ? node1117 : node1104;
												assign node1104 = (inp[1]) ? node1110 : node1105;
													assign node1105 = (inp[8]) ? node1107 : 4'b0001;
														assign node1107 = (inp[5]) ? 4'b0001 : 4'b0011;
													assign node1110 = (inp[5]) ? 4'b1011 : node1111;
														assign node1111 = (inp[8]) ? node1113 : 4'b0011;
															assign node1113 = (inp[10]) ? 4'b0001 : 4'b0011;
												assign node1117 = (inp[1]) ? node1121 : node1118;
													assign node1118 = (inp[5]) ? 4'b1000 : 4'b1010;
													assign node1121 = (inp[5]) ? 4'b1001 : node1122;
														assign node1122 = (inp[8]) ? 4'b1011 : 4'b1001;
											assign node1126 = (inp[11]) ? node1134 : node1127;
												assign node1127 = (inp[1]) ? 4'b1011 : node1128;
													assign node1128 = (inp[5]) ? 4'b0011 : node1129;
														assign node1129 = (inp[8]) ? 4'b1001 : 4'b1011;
												assign node1134 = (inp[1]) ? 4'b0011 : node1135;
													assign node1135 = (inp[8]) ? 4'b0001 : node1136;
														assign node1136 = (inp[5]) ? 4'b0011 : 4'b0001;
										assign node1141 = (inp[6]) ? node1163 : node1142;
											assign node1142 = (inp[11]) ? node1152 : node1143;
												assign node1143 = (inp[5]) ? node1147 : node1144;
													assign node1144 = (inp[1]) ? 4'b0001 : 4'b0011;
													assign node1147 = (inp[1]) ? node1149 : 4'b0001;
														assign node1149 = (inp[8]) ? 4'b1001 : 4'b1011;
												assign node1152 = (inp[1]) ? node1156 : node1153;
													assign node1153 = (inp[10]) ? 4'b1000 : 4'b1010;
													assign node1156 = (inp[5]) ? 4'b0011 : node1157;
														assign node1157 = (inp[8]) ? node1159 : 4'b1011;
															assign node1159 = (inp[10]) ? 4'b1001 : 4'b1011;
											assign node1163 = (inp[11]) ? node1171 : node1164;
												assign node1164 = (inp[1]) ? 4'b1001 : node1165;
													assign node1165 = (inp[5]) ? node1167 : 4'b1001;
														assign node1167 = (inp[8]) ? 4'b0001 : 4'b0011;
												assign node1171 = (inp[1]) ? 4'b0001 : node1172;
													assign node1172 = (inp[5]) ? 4'b0001 : 4'b0011;
									assign node1176 = (inp[1]) ? node1226 : node1177;
										assign node1177 = (inp[11]) ? node1195 : node1178;
											assign node1178 = (inp[5]) ? node1190 : node1179;
												assign node1179 = (inp[15]) ? node1181 : 4'b1010;
													assign node1181 = (inp[8]) ? 4'b1000 : node1182;
														assign node1182 = (inp[2]) ? node1184 : 4'b1010;
															assign node1184 = (inp[10]) ? node1186 : 4'b1010;
																assign node1186 = (inp[6]) ? 4'b1010 : 4'b1000;
												assign node1190 = (inp[15]) ? node1192 : 4'b1000;
													assign node1192 = (inp[6]) ? 4'b1010 : 4'b0010;
											assign node1195 = (inp[5]) ? node1209 : node1196;
												assign node1196 = (inp[6]) ? node1204 : node1197;
													assign node1197 = (inp[15]) ? 4'b0000 : node1198;
														assign node1198 = (inp[10]) ? node1200 : 4'b0010;
															assign node1200 = (inp[8]) ? 4'b0000 : 4'b0010;
													assign node1204 = (inp[8]) ? 4'b1000 : node1205;
														assign node1205 = (inp[15]) ? 4'b1000 : 4'b1010;
												assign node1209 = (inp[2]) ? node1217 : node1210;
													assign node1210 = (inp[8]) ? node1212 : 4'b0010;
														assign node1212 = (inp[15]) ? node1214 : 4'b0010;
															assign node1214 = (inp[6]) ? 4'b0000 : 4'b0010;
													assign node1217 = (inp[10]) ? node1223 : node1218;
														assign node1218 = (inp[15]) ? 4'b0010 : node1219;
															assign node1219 = (inp[6]) ? 4'b0010 : 4'b0000;
														assign node1223 = (inp[15]) ? 4'b0000 : 4'b0010;
										assign node1226 = (inp[15]) ? node1248 : node1227;
											assign node1227 = (inp[11]) ? node1241 : node1228;
												assign node1228 = (inp[6]) ? 4'b1011 : node1229;
													assign node1229 = (inp[8]) ? node1235 : node1230;
														assign node1230 = (inp[5]) ? 4'b0011 : node1231;
															assign node1231 = (inp[2]) ? 4'b0001 : 4'b0011;
														assign node1235 = (inp[10]) ? 4'b0001 : node1236;
															assign node1236 = (inp[5]) ? 4'b0011 : 4'b0001;
												assign node1241 = (inp[6]) ? 4'b0011 : node1242;
													assign node1242 = (inp[8]) ? 4'b1010 : node1243;
														assign node1243 = (inp[5]) ? 4'b1000 : 4'b1010;
											assign node1248 = (inp[6]) ? node1266 : node1249;
												assign node1249 = (inp[11]) ? node1255 : node1250;
													assign node1250 = (inp[8]) ? node1252 : 4'b0001;
														assign node1252 = (inp[5]) ? 4'b0001 : 4'b0011;
													assign node1255 = (inp[2]) ? node1261 : node1256;
														assign node1256 = (inp[10]) ? 4'b1000 : node1257;
															assign node1257 = (inp[8]) ? 4'b1000 : 4'b1010;
														assign node1261 = (inp[8]) ? node1263 : 4'b1010;
															assign node1263 = (inp[10]) ? 4'b1000 : 4'b1010;
												assign node1266 = (inp[11]) ? 4'b0001 : 4'b1001;
								assign node1269 = (inp[6]) ? node1363 : node1270;
									assign node1270 = (inp[1]) ? node1348 : node1271;
										assign node1271 = (inp[4]) ? node1309 : node1272;
											assign node1272 = (inp[5]) ? node1290 : node1273;
												assign node1273 = (inp[11]) ? node1281 : node1274;
													assign node1274 = (inp[15]) ? node1278 : node1275;
														assign node1275 = (inp[8]) ? 4'b0010 : 4'b0000;
														assign node1278 = (inp[8]) ? 4'b0000 : 4'b0010;
													assign node1281 = (inp[15]) ? node1287 : node1282;
														assign node1282 = (inp[8]) ? 4'b1000 : node1283;
															assign node1283 = (inp[10]) ? 4'b1000 : 4'b1010;
														assign node1287 = (inp[8]) ? 4'b0000 : 4'b0010;
												assign node1290 = (inp[11]) ? node1300 : node1291;
													assign node1291 = (inp[8]) ? node1295 : node1292;
														assign node1292 = (inp[15]) ? 4'b1000 : 4'b1010;
														assign node1295 = (inp[10]) ? node1297 : 4'b1010;
															assign node1297 = (inp[15]) ? 4'b1010 : 4'b1000;
													assign node1300 = (inp[15]) ? node1304 : node1301;
														assign node1301 = (inp[8]) ? 4'b0010 : 4'b0000;
														assign node1304 = (inp[8]) ? 4'b0000 : node1305;
															assign node1305 = (inp[10]) ? 4'b0000 : 4'b0010;
											assign node1309 = (inp[5]) ? node1327 : node1310;
												assign node1310 = (inp[11]) ? node1316 : node1311;
													assign node1311 = (inp[8]) ? 4'b1011 : node1312;
														assign node1312 = (inp[15]) ? 4'b1001 : 4'b1011;
													assign node1316 = (inp[10]) ? node1322 : node1317;
														assign node1317 = (inp[8]) ? 4'b0001 : node1318;
															assign node1318 = (inp[15]) ? 4'b0011 : 4'b0001;
														assign node1322 = (inp[8]) ? node1324 : 4'b0001;
															assign node1324 = (inp[15]) ? 4'b0001 : 4'b0011;
												assign node1327 = (inp[15]) ? node1339 : node1328;
													assign node1328 = (inp[8]) ? node1334 : node1329;
														assign node1329 = (inp[11]) ? 4'b1011 : node1330;
															assign node1330 = (inp[10]) ? 4'b1001 : 4'b1011;
														assign node1334 = (inp[10]) ? 4'b1001 : node1335;
															assign node1335 = (inp[11]) ? 4'b1011 : 4'b1001;
													assign node1339 = (inp[11]) ? node1345 : node1340;
														assign node1340 = (inp[10]) ? node1342 : 4'b0011;
															assign node1342 = (inp[8]) ? 4'b0001 : 4'b0011;
														assign node1345 = (inp[8]) ? 4'b1011 : 4'b1001;
										assign node1348 = (inp[10]) ? node1356 : node1349;
											assign node1349 = (inp[15]) ? node1353 : node1350;
												assign node1350 = (inp[11]) ? 4'b1110 : 4'b1111;
												assign node1353 = (inp[11]) ? 4'b0110 : 4'b0111;
											assign node1356 = (inp[15]) ? node1360 : node1357;
												assign node1357 = (inp[11]) ? 4'b1100 : 4'b1101;
												assign node1360 = (inp[11]) ? 4'b0100 : 4'b0101;
									assign node1363 = (inp[1]) ? 4'b0000 : node1364;
										assign node1364 = (inp[4]) ? node1372 : node1365;
											assign node1365 = (inp[8]) ? node1369 : node1366;
												assign node1366 = (inp[5]) ? 4'b0011 : 4'b1011;
												assign node1369 = (inp[5]) ? 4'b0001 : 4'b1001;
											assign node1372 = (inp[5]) ? node1376 : node1373;
												assign node1373 = (inp[8]) ? 4'b1000 : 4'b1010;
												assign node1376 = (inp[8]) ? 4'b0000 : 4'b0010;
			assign node1380 = (inp[0]) ? node1382 : 4'b0000;
				assign node1382 = (inp[4]) ? node1928 : node1383;
					assign node1383 = (inp[7]) ? node1573 : node1384;
						assign node1384 = (inp[3]) ? node1456 : node1385;
							assign node1385 = (inp[11]) ? 4'b0000 : node1386;
								assign node1386 = (inp[9]) ? node1422 : node1387;
									assign node1387 = (inp[5]) ? 4'b0000 : node1388;
										assign node1388 = (inp[13]) ? node1404 : node1389;
											assign node1389 = (inp[15]) ? 4'b0000 : node1390;
												assign node1390 = (inp[1]) ? node1398 : node1391;
													assign node1391 = (inp[8]) ? 4'b0000 : node1392;
														assign node1392 = (inp[6]) ? 4'b0010 : node1393;
															assign node1393 = (inp[10]) ? 4'b0000 : 4'b0010;
													assign node1398 = (inp[10]) ? node1400 : 4'b0010;
														assign node1400 = (inp[6]) ? 4'b0010 : 4'b0000;
											assign node1404 = (inp[15]) ? node1406 : 4'b0010;
												assign node1406 = (inp[1]) ? node1414 : node1407;
													assign node1407 = (inp[8]) ? 4'b0000 : node1408;
														assign node1408 = (inp[10]) ? node1410 : 4'b0010;
															assign node1410 = (inp[6]) ? 4'b0010 : 4'b0000;
													assign node1414 = (inp[8]) ? node1416 : 4'b0010;
														assign node1416 = (inp[6]) ? 4'b0010 : node1417;
															assign node1417 = (inp[10]) ? 4'b0000 : 4'b0010;
									assign node1422 = (inp[5]) ? node1424 : 4'b0010;
										assign node1424 = (inp[15]) ? node1440 : node1425;
											assign node1425 = (inp[13]) ? 4'b0010 : node1426;
												assign node1426 = (inp[6]) ? 4'b0010 : node1427;
													assign node1427 = (inp[10]) ? node1433 : node1428;
														assign node1428 = (inp[8]) ? node1430 : 4'b0010;
															assign node1430 = (inp[1]) ? 4'b0010 : 4'b0000;
														assign node1433 = (inp[8]) ? 4'b0000 : node1434;
															assign node1434 = (inp[1]) ? 4'b0010 : 4'b0000;
											assign node1440 = (inp[13]) ? node1442 : 4'b0000;
												assign node1442 = (inp[8]) ? node1450 : node1443;
													assign node1443 = (inp[10]) ? node1445 : 4'b0010;
														assign node1445 = (inp[1]) ? 4'b0010 : node1446;
															assign node1446 = (inp[6]) ? 4'b0010 : 4'b0000;
													assign node1450 = (inp[1]) ? node1452 : 4'b0000;
														assign node1452 = (inp[6]) ? 4'b0010 : 4'b0000;
							assign node1456 = (inp[11]) ? node1534 : node1457;
								assign node1457 = (inp[13]) ? node1487 : node1458;
									assign node1458 = (inp[9]) ? node1476 : node1459;
										assign node1459 = (inp[5]) ? 4'b0010 : node1460;
											assign node1460 = (inp[15]) ? node1468 : node1461;
												assign node1461 = (inp[6]) ? 4'b0000 : node1462;
													assign node1462 = (inp[8]) ? node1464 : 4'b0000;
														assign node1464 = (inp[1]) ? 4'b0000 : 4'b0010;
												assign node1468 = (inp[1]) ? node1470 : 4'b0010;
													assign node1470 = (inp[8]) ? node1472 : 4'b0000;
														assign node1472 = (inp[6]) ? 4'b0000 : 4'b0010;
										assign node1476 = (inp[15]) ? 4'b0000 : node1477;
											assign node1477 = (inp[1]) ? node1479 : 4'b0000;
												assign node1479 = (inp[5]) ? 4'b0000 : node1480;
													assign node1480 = (inp[6]) ? 4'b0010 : node1481;
														assign node1481 = (inp[10]) ? 4'b0000 : 4'b0010;
									assign node1487 = (inp[9]) ? node1505 : node1488;
										assign node1488 = (inp[5]) ? node1490 : 4'b0000;
											assign node1490 = (inp[1]) ? node1498 : node1491;
												assign node1491 = (inp[15]) ? 4'b0010 : node1492;
													assign node1492 = (inp[8]) ? node1494 : 4'b0000;
														assign node1494 = (inp[6]) ? 4'b0000 : 4'b0010;
												assign node1498 = (inp[6]) ? 4'b0000 : node1499;
													assign node1499 = (inp[15]) ? node1501 : 4'b0000;
														assign node1501 = (inp[8]) ? 4'b0010 : 4'b0000;
										assign node1505 = (inp[5]) ? node1517 : node1506;
											assign node1506 = (inp[1]) ? 4'b0010 : node1507;
												assign node1507 = (inp[15]) ? node1509 : 4'b0010;
													assign node1509 = (inp[6]) ? 4'b0010 : node1510;
														assign node1510 = (inp[10]) ? node1512 : 4'b0010;
															assign node1512 = (inp[8]) ? 4'b0000 : 4'b0010;
											assign node1517 = (inp[1]) ? node1525 : node1518;
												assign node1518 = (inp[8]) ? 4'b0000 : node1519;
													assign node1519 = (inp[15]) ? 4'b0000 : node1520;
														assign node1520 = (inp[6]) ? 4'b0010 : 4'b0000;
												assign node1525 = (inp[15]) ? node1527 : 4'b0010;
													assign node1527 = (inp[6]) ? 4'b0010 : node1528;
														assign node1528 = (inp[10]) ? 4'b0000 : node1529;
															assign node1529 = (inp[8]) ? 4'b0000 : 4'b0010;
								assign node1534 = (inp[9]) ? node1536 : 4'b0010;
									assign node1536 = (inp[13]) ? node1554 : node1537;
										assign node1537 = (inp[5]) ? 4'b0010 : node1538;
											assign node1538 = (inp[15]) ? node1546 : node1539;
												assign node1539 = (inp[6]) ? 4'b0000 : node1540;
													assign node1540 = (inp[8]) ? node1542 : 4'b0000;
														assign node1542 = (inp[1]) ? 4'b0000 : 4'b0010;
												assign node1546 = (inp[1]) ? node1548 : 4'b0010;
													assign node1548 = (inp[8]) ? node1550 : 4'b0000;
														assign node1550 = (inp[6]) ? 4'b0000 : 4'b0010;
										assign node1554 = (inp[15]) ? node1564 : node1555;
											assign node1555 = (inp[6]) ? 4'b0000 : node1556;
												assign node1556 = (inp[1]) ? 4'b0000 : node1557;
													assign node1557 = (inp[5]) ? node1559 : 4'b0000;
														assign node1559 = (inp[8]) ? 4'b0010 : 4'b0000;
											assign node1564 = (inp[5]) ? node1566 : 4'b0000;
												assign node1566 = (inp[1]) ? node1568 : 4'b0010;
													assign node1568 = (inp[6]) ? 4'b0000 : node1569;
														assign node1569 = (inp[8]) ? 4'b0010 : 4'b0000;
						assign node1573 = (inp[3]) ? node1639 : node1574;
							assign node1574 = (inp[11]) ? node1576 : 4'b0010;
								assign node1576 = (inp[5]) ? node1608 : node1577;
									assign node1577 = (inp[9]) ? 4'b0010 : node1578;
										assign node1578 = (inp[15]) ? node1596 : node1579;
											assign node1579 = (inp[13]) ? 4'b0010 : node1580;
												assign node1580 = (inp[8]) ? node1588 : node1581;
													assign node1581 = (inp[1]) ? 4'b0010 : node1582;
														assign node1582 = (inp[6]) ? 4'b0010 : node1583;
															assign node1583 = (inp[10]) ? 4'b0000 : 4'b0010;
													assign node1588 = (inp[1]) ? node1590 : 4'b0000;
														assign node1590 = (inp[10]) ? node1592 : 4'b0010;
															assign node1592 = (inp[6]) ? 4'b0010 : 4'b0000;
											assign node1596 = (inp[13]) ? node1598 : 4'b0000;
												assign node1598 = (inp[1]) ? 4'b0010 : node1599;
													assign node1599 = (inp[8]) ? 4'b0000 : node1600;
														assign node1600 = (inp[6]) ? 4'b0010 : node1601;
															assign node1601 = (inp[10]) ? 4'b0000 : 4'b0010;
									assign node1608 = (inp[9]) ? node1610 : 4'b0000;
										assign node1610 = (inp[15]) ? node1626 : node1611;
											assign node1611 = (inp[13]) ? 4'b0010 : node1612;
												assign node1612 = (inp[6]) ? node1620 : node1613;
													assign node1613 = (inp[10]) ? 4'b0000 : node1614;
														assign node1614 = (inp[1]) ? 4'b0010 : node1615;
															assign node1615 = (inp[8]) ? 4'b0000 : 4'b0010;
													assign node1620 = (inp[1]) ? 4'b0010 : node1621;
														assign node1621 = (inp[8]) ? 4'b0000 : 4'b0010;
											assign node1626 = (inp[13]) ? node1628 : 4'b0000;
												assign node1628 = (inp[8]) ? node1634 : node1629;
													assign node1629 = (inp[6]) ? 4'b0010 : node1630;
														assign node1630 = (inp[10]) ? 4'b0000 : 4'b0010;
													assign node1634 = (inp[1]) ? node1636 : 4'b0000;
														assign node1636 = (inp[10]) ? 4'b0000 : 4'b0010;
							assign node1639 = (inp[13]) ? node1795 : node1640;
								assign node1640 = (inp[9]) ? node1688 : node1641;
									assign node1641 = (inp[11]) ? node1661 : node1642;
										assign node1642 = (inp[5]) ? node1654 : node1643;
											assign node1643 = (inp[6]) ? node1649 : node1644;
												assign node1644 = (inp[1]) ? 4'b1000 : node1645;
													assign node1645 = (inp[15]) ? 4'b0010 : 4'b1000;
												assign node1649 = (inp[1]) ? node1651 : 4'b1000;
													assign node1651 = (inp[15]) ? 4'b1000 : 4'b1010;
											assign node1654 = (inp[1]) ? node1656 : 4'b0010;
												assign node1656 = (inp[15]) ? node1658 : 4'b1000;
													assign node1658 = (inp[6]) ? 4'b1000 : 4'b0010;
										assign node1661 = (inp[5]) ? node1677 : node1662;
											assign node1662 = (inp[1]) ? 4'b0010 : node1663;
												assign node1663 = (inp[15]) ? node1671 : node1664;
													assign node1664 = (inp[8]) ? node1666 : 4'b0010;
														assign node1666 = (inp[2]) ? 4'b0010 : node1667;
															assign node1667 = (inp[10]) ? 4'b0000 : 4'b0010;
													assign node1671 = (inp[6]) ? node1673 : 4'b0000;
														assign node1673 = (inp[8]) ? 4'b0000 : 4'b0010;
											assign node1677 = (inp[1]) ? node1679 : 4'b0000;
												assign node1679 = (inp[15]) ? 4'b0000 : node1680;
													assign node1680 = (inp[6]) ? 4'b0010 : node1681;
														assign node1681 = (inp[8]) ? 4'b0000 : node1682;
															assign node1682 = (inp[10]) ? 4'b0000 : 4'b0010;
									assign node1688 = (inp[15]) ? node1750 : node1689;
										assign node1689 = (inp[11]) ? node1713 : node1690;
											assign node1690 = (inp[1]) ? node1704 : node1691;
												assign node1691 = (inp[5]) ? node1699 : node1692;
													assign node1692 = (inp[8]) ? 4'b0000 : node1693;
														assign node1693 = (inp[2]) ? 4'b0000 : node1694;
															assign node1694 = (inp[6]) ? 4'b0000 : 4'b0010;
													assign node1699 = (inp[6]) ? node1701 : 4'b1010;
														assign node1701 = (inp[8]) ? 4'b0000 : 4'b0010;
												assign node1704 = (inp[6]) ? 4'b1010 : node1705;
													assign node1705 = (inp[5]) ? node1707 : 4'b1000;
														assign node1707 = (inp[10]) ? 4'b0000 : node1708;
															assign node1708 = (inp[8]) ? 4'b0000 : 4'b0010;
											assign node1713 = (inp[1]) ? node1739 : node1714;
												assign node1714 = (inp[10]) ? node1730 : node1715;
													assign node1715 = (inp[8]) ? node1723 : node1716;
														assign node1716 = (inp[5]) ? node1720 : node1717;
															assign node1717 = (inp[6]) ? 4'b1010 : 4'b1000;
															assign node1720 = (inp[6]) ? 4'b1000 : 4'b1010;
														assign node1723 = (inp[5]) ? node1727 : node1724;
															assign node1724 = (inp[6]) ? 4'b1010 : 4'b1000;
															assign node1727 = (inp[6]) ? 4'b1000 : 4'b1010;
													assign node1730 = (inp[8]) ? node1732 : 4'b1010;
														assign node1732 = (inp[6]) ? node1736 : node1733;
															assign node1733 = (inp[5]) ? 4'b1010 : 4'b1000;
															assign node1736 = (inp[5]) ? 4'b1000 : 4'b1010;
												assign node1739 = (inp[5]) ? node1747 : node1740;
													assign node1740 = (inp[6]) ? 4'b0010 : node1741;
														assign node1741 = (inp[10]) ? node1743 : 4'b0010;
															assign node1743 = (inp[8]) ? 4'b0000 : 4'b0010;
													assign node1747 = (inp[6]) ? 4'b0010 : 4'b1010;
										assign node1750 = (inp[1]) ? node1778 : node1751;
											assign node1751 = (inp[11]) ? node1763 : node1752;
												assign node1752 = (inp[5]) ? node1756 : node1753;
													assign node1753 = (inp[6]) ? 4'b0010 : 4'b0000;
													assign node1756 = (inp[6]) ? 4'b0000 : node1757;
														assign node1757 = (inp[10]) ? node1759 : 4'b1010;
															assign node1759 = (inp[8]) ? 4'b1000 : 4'b1010;
												assign node1763 = (inp[6]) ? node1773 : node1764;
													assign node1764 = (inp[8]) ? node1770 : node1765;
														assign node1765 = (inp[5]) ? node1767 : 4'b1000;
															assign node1767 = (inp[10]) ? 4'b1000 : 4'b1010;
														assign node1770 = (inp[5]) ? 4'b1000 : 4'b1010;
													assign node1773 = (inp[5]) ? 4'b1010 : node1774;
														assign node1774 = (inp[8]) ? 4'b1000 : 4'b1010;
											assign node1778 = (inp[11]) ? node1786 : node1779;
												assign node1779 = (inp[6]) ? 4'b1000 : node1780;
													assign node1780 = (inp[5]) ? node1782 : 4'b0010;
														assign node1782 = (inp[8]) ? 4'b0010 : 4'b0000;
												assign node1786 = (inp[6]) ? 4'b0000 : node1787;
													assign node1787 = (inp[5]) ? node1789 : 4'b0000;
														assign node1789 = (inp[2]) ? node1791 : 4'b1000;
															assign node1791 = (inp[10]) ? 4'b1000 : 4'b1010;
								assign node1795 = (inp[9]) ? node1863 : node1796;
									assign node1796 = (inp[11]) ? node1834 : node1797;
										assign node1797 = (inp[5]) ? node1813 : node1798;
											assign node1798 = (inp[6]) ? node1808 : node1799;
												assign node1799 = (inp[1]) ? node1801 : 4'b1010;
													assign node1801 = (inp[10]) ? 4'b1000 : node1802;
														assign node1802 = (inp[8]) ? 4'b1000 : node1803;
															assign node1803 = (inp[15]) ? 4'b1000 : 4'b1010;
												assign node1808 = (inp[1]) ? 4'b1010 : node1809;
													assign node1809 = (inp[15]) ? 4'b1010 : 4'b1000;
											assign node1813 = (inp[6]) ? node1827 : node1814;
												assign node1814 = (inp[1]) ? node1822 : node1815;
													assign node1815 = (inp[8]) ? 4'b1000 : node1816;
														assign node1816 = (inp[15]) ? 4'b1000 : node1817;
															assign node1817 = (inp[10]) ? 4'b1000 : 4'b1010;
													assign node1822 = (inp[8]) ? 4'b1010 : node1823;
														assign node1823 = (inp[15]) ? 4'b1010 : 4'b1000;
												assign node1827 = (inp[1]) ? 4'b1000 : node1828;
													assign node1828 = (inp[15]) ? node1830 : 4'b1010;
														assign node1830 = (inp[8]) ? 4'b1000 : 4'b1010;
										assign node1834 = (inp[1]) ? node1850 : node1835;
											assign node1835 = (inp[5]) ? node1841 : node1836;
												assign node1836 = (inp[6]) ? 4'b1000 : node1837;
													assign node1837 = (inp[15]) ? 4'b0010 : 4'b1000;
												assign node1841 = (inp[8]) ? node1843 : 4'b0010;
													assign node1843 = (inp[10]) ? node1845 : 4'b0010;
														assign node1845 = (inp[15]) ? node1847 : 4'b0010;
															assign node1847 = (inp[6]) ? 4'b0010 : 4'b0000;
											assign node1850 = (inp[5]) ? node1858 : node1851;
												assign node1851 = (inp[6]) ? 4'b1010 : node1852;
													assign node1852 = (inp[15]) ? 4'b1000 : node1853;
														assign node1853 = (inp[10]) ? 4'b1000 : 4'b1010;
												assign node1858 = (inp[15]) ? node1860 : 4'b1000;
													assign node1860 = (inp[6]) ? 4'b1000 : 4'b0010;
									assign node1863 = (inp[1]) ? node1911 : node1864;
										assign node1864 = (inp[5]) ? node1886 : node1865;
											assign node1865 = (inp[8]) ? node1877 : node1866;
												assign node1866 = (inp[6]) ? 4'b1011 : node1867;
													assign node1867 = (inp[11]) ? node1873 : node1868;
														assign node1868 = (inp[15]) ? 4'b0011 : node1869;
															assign node1869 = (inp[10]) ? 4'b1001 : 4'b1011;
														assign node1873 = (inp[15]) ? 4'b1000 : 4'b1010;
												assign node1877 = (inp[6]) ? 4'b1001 : node1878;
													assign node1878 = (inp[15]) ? node1882 : node1879;
														assign node1879 = (inp[11]) ? 4'b1000 : 4'b1001;
														assign node1882 = (inp[11]) ? 4'b1010 : 4'b0011;
											assign node1886 = (inp[6]) ? node1908 : node1887;
												assign node1887 = (inp[11]) ? node1897 : node1888;
													assign node1888 = (inp[8]) ? node1894 : node1889;
														assign node1889 = (inp[15]) ? node1891 : 4'b0001;
															assign node1891 = (inp[10]) ? 4'b0001 : 4'b0011;
														assign node1894 = (inp[15]) ? 4'b0001 : 4'b0011;
													assign node1897 = (inp[15]) ? node1903 : node1898;
														assign node1898 = (inp[8]) ? 4'b1000 : node1899;
															assign node1899 = (inp[10]) ? 4'b1000 : 4'b1010;
														assign node1903 = (inp[10]) ? node1905 : 4'b0010;
															assign node1905 = (inp[8]) ? 4'b0000 : 4'b0010;
												assign node1908 = (inp[8]) ? 4'b0001 : 4'b0011;
										assign node1911 = (inp[6]) ? 4'b0000 : node1912;
											assign node1912 = (inp[10]) ? node1920 : node1913;
												assign node1913 = (inp[15]) ? node1917 : node1914;
													assign node1914 = (inp[11]) ? 4'b1010 : 4'b1011;
													assign node1917 = (inp[11]) ? 4'b0010 : 4'b0011;
												assign node1920 = (inp[11]) ? node1924 : node1921;
													assign node1921 = (inp[15]) ? 4'b0001 : 4'b1001;
													assign node1924 = (inp[15]) ? 4'b0000 : 4'b1000;
					assign node1928 = (inp[3]) ? node1930 : 4'b0000;
						assign node1930 = (inp[11]) ? node2130 : node1931;
							assign node1931 = (inp[9]) ? node2021 : node1932;
								assign node1932 = (inp[7]) ? node1968 : node1933;
									assign node1933 = (inp[5]) ? 4'b0000 : node1934;
										assign node1934 = (inp[13]) ? node1950 : node1935;
											assign node1935 = (inp[15]) ? 4'b0000 : node1936;
												assign node1936 = (inp[8]) ? node1944 : node1937;
													assign node1937 = (inp[6]) ? 4'b0010 : node1938;
														assign node1938 = (inp[10]) ? node1940 : 4'b0010;
															assign node1940 = (inp[1]) ? 4'b0010 : 4'b0000;
													assign node1944 = (inp[1]) ? node1946 : 4'b0000;
														assign node1946 = (inp[6]) ? 4'b0010 : 4'b0000;
											assign node1950 = (inp[15]) ? node1952 : 4'b0010;
												assign node1952 = (inp[8]) ? node1960 : node1953;
													assign node1953 = (inp[6]) ? 4'b0010 : node1954;
														assign node1954 = (inp[1]) ? 4'b0010 : node1955;
															assign node1955 = (inp[10]) ? 4'b0000 : 4'b0010;
													assign node1960 = (inp[1]) ? node1962 : 4'b0000;
														assign node1962 = (inp[10]) ? node1964 : 4'b0010;
															assign node1964 = (inp[6]) ? 4'b0010 : 4'b0000;
									assign node1968 = (inp[13]) ? node1988 : node1969;
										assign node1969 = (inp[5]) ? 4'b0010 : node1970;
											assign node1970 = (inp[15]) ? node1980 : node1971;
												assign node1971 = (inp[2]) ? node1973 : 4'b0000;
													assign node1973 = (inp[1]) ? 4'b0000 : node1974;
														assign node1974 = (inp[6]) ? 4'b0000 : node1975;
															assign node1975 = (inp[8]) ? 4'b0010 : 4'b0000;
												assign node1980 = (inp[1]) ? node1982 : 4'b0010;
													assign node1982 = (inp[6]) ? 4'b0000 : node1983;
														assign node1983 = (inp[8]) ? 4'b0010 : 4'b0000;
										assign node1988 = (inp[15]) ? node2004 : node1989;
											assign node1989 = (inp[5]) ? node1997 : node1990;
												assign node1990 = (inp[1]) ? 4'b0010 : node1991;
													assign node1991 = (inp[6]) ? node1993 : 4'b0000;
														assign node1993 = (inp[8]) ? 4'b0000 : 4'b0010;
												assign node1997 = (inp[1]) ? 4'b0000 : node1998;
													assign node1998 = (inp[8]) ? node2000 : 4'b0000;
														assign node2000 = (inp[6]) ? 4'b0000 : 4'b0010;
											assign node2004 = (inp[5]) ? node2014 : node2005;
												assign node2005 = (inp[1]) ? node2007 : 4'b0000;
													assign node2007 = (inp[6]) ? 4'b0010 : node2008;
														assign node2008 = (inp[10]) ? 4'b0000 : node2009;
															assign node2009 = (inp[8]) ? 4'b0000 : 4'b0010;
												assign node2014 = (inp[1]) ? node2016 : 4'b0010;
													assign node2016 = (inp[8]) ? node2018 : 4'b0000;
														assign node2018 = (inp[6]) ? 4'b0000 : 4'b0010;
								assign node2021 = (inp[7]) ? node2053 : node2022;
									assign node2022 = (inp[5]) ? node2024 : 4'b0010;
										assign node2024 = (inp[15]) ? node2036 : node2025;
											assign node2025 = (inp[8]) ? node2027 : 4'b0010;
												assign node2027 = (inp[13]) ? 4'b0010 : node2028;
													assign node2028 = (inp[1]) ? node2030 : 4'b0000;
														assign node2030 = (inp[6]) ? 4'b0010 : node2031;
															assign node2031 = (inp[10]) ? 4'b0000 : 4'b0010;
											assign node2036 = (inp[13]) ? node2038 : 4'b0000;
												assign node2038 = (inp[8]) ? node2046 : node2039;
													assign node2039 = (inp[10]) ? node2041 : 4'b0010;
														assign node2041 = (inp[6]) ? 4'b0010 : node2042;
															assign node2042 = (inp[1]) ? 4'b0010 : 4'b0000;
													assign node2046 = (inp[1]) ? node2048 : 4'b0000;
														assign node2048 = (inp[6]) ? 4'b0010 : node2049;
															assign node2049 = (inp[10]) ? 4'b0000 : 4'b0010;
									assign node2053 = (inp[13]) ? node2097 : node2054;
										assign node2054 = (inp[5]) ? node2076 : node2055;
											assign node2055 = (inp[6]) ? node2069 : node2056;
												assign node2056 = (inp[15]) ? node2062 : node2057;
													assign node2057 = (inp[1]) ? node2059 : 4'b1000;
														assign node2059 = (inp[8]) ? 4'b1010 : 4'b1000;
													assign node2062 = (inp[1]) ? node2064 : 4'b0010;
														assign node2064 = (inp[8]) ? node2066 : 4'b1010;
															assign node2066 = (inp[10]) ? 4'b1000 : 4'b1010;
												assign node2069 = (inp[15]) ? 4'b1000 : node2070;
													assign node2070 = (inp[8]) ? node2072 : 4'b1010;
														assign node2072 = (inp[1]) ? 4'b1010 : 4'b1000;
											assign node2076 = (inp[1]) ? node2090 : node2077;
												assign node2077 = (inp[15]) ? node2085 : node2078;
													assign node2078 = (inp[6]) ? 4'b0010 : node2079;
														assign node2079 = (inp[10]) ? node2081 : 4'b0010;
															assign node2081 = (inp[8]) ? 4'b0000 : 4'b0010;
													assign node2085 = (inp[8]) ? 4'b0000 : node2086;
														assign node2086 = (inp[6]) ? 4'b0010 : 4'b0000;
												assign node2090 = (inp[15]) ? node2094 : node2091;
													assign node2091 = (inp[6]) ? 4'b1010 : 4'b1000;
													assign node2094 = (inp[6]) ? 4'b1000 : 4'b0010;
										assign node2097 = (inp[6]) ? node2121 : node2098;
											assign node2098 = (inp[1]) ? node2114 : node2099;
												assign node2099 = (inp[5]) ? node2107 : node2100;
													assign node2100 = (inp[8]) ? node2104 : node2101;
														assign node2101 = (inp[15]) ? 4'b0010 : 4'b0000;
														assign node2104 = (inp[15]) ? 4'b0000 : 4'b0010;
													assign node2107 = (inp[10]) ? node2109 : 4'b1010;
														assign node2109 = (inp[15]) ? node2111 : 4'b1000;
															assign node2111 = (inp[8]) ? 4'b1010 : 4'b1000;
												assign node2114 = (inp[10]) ? node2118 : node2115;
													assign node2115 = (inp[15]) ? 4'b0011 : 4'b1011;
													assign node2118 = (inp[15]) ? 4'b0001 : 4'b1001;
											assign node2121 = (inp[1]) ? 4'b0000 : node2122;
												assign node2122 = (inp[5]) ? node2126 : node2123;
													assign node2123 = (inp[8]) ? 4'b1000 : 4'b1010;
													assign node2126 = (inp[8]) ? 4'b0000 : 4'b0010;
							assign node2130 = (inp[7]) ? node2132 : 4'b0000;
								assign node2132 = (inp[5]) ? node2214 : node2133;
									assign node2133 = (inp[13]) ? node2177 : node2134;
										assign node2134 = (inp[15]) ? node2168 : node2135;
											assign node2135 = (inp[1]) ? node2155 : node2136;
												assign node2136 = (inp[10]) ? node2148 : node2137;
													assign node2137 = (inp[2]) ? 4'b0010 : node2138;
														assign node2138 = (inp[8]) ? node2142 : node2139;
															assign node2139 = (inp[9]) ? 4'b0000 : 4'b0010;
															assign node2142 = (inp[6]) ? 4'b0000 : node2143;
																assign node2143 = (inp[9]) ? 4'b0010 : 4'b0000;
													assign node2148 = (inp[9]) ? 4'b0000 : node2149;
														assign node2149 = (inp[6]) ? node2151 : 4'b0000;
															assign node2151 = (inp[8]) ? 4'b0000 : 4'b0010;
												assign node2155 = (inp[6]) ? 4'b0010 : node2156;
													assign node2156 = (inp[9]) ? node2162 : node2157;
														assign node2157 = (inp[8]) ? node2159 : 4'b0010;
															assign node2159 = (inp[10]) ? 4'b0000 : 4'b0010;
														assign node2162 = (inp[10]) ? 4'b0000 : node2163;
															assign node2163 = (inp[8]) ? 4'b0000 : 4'b0010;
											assign node2168 = (inp[9]) ? node2170 : 4'b0000;
												assign node2170 = (inp[1]) ? node2172 : 4'b0010;
													assign node2172 = (inp[6]) ? 4'b0000 : node2173;
														assign node2173 = (inp[8]) ? 4'b0010 : 4'b0000;
										assign node2177 = (inp[9]) ? node2187 : node2178;
											assign node2178 = (inp[15]) ? node2180 : 4'b0010;
												assign node2180 = (inp[1]) ? 4'b0010 : node2181;
													assign node2181 = (inp[8]) ? 4'b0000 : node2182;
														assign node2182 = (inp[10]) ? 4'b0000 : 4'b0010;
											assign node2187 = (inp[15]) ? node2201 : node2188;
												assign node2188 = (inp[6]) ? node2196 : node2189;
													assign node2189 = (inp[10]) ? 4'b1000 : node2190;
														assign node2190 = (inp[8]) ? node2192 : 4'b1010;
															assign node2192 = (inp[1]) ? 4'b1010 : 4'b1000;
													assign node2196 = (inp[1]) ? 4'b0000 : node2197;
														assign node2197 = (inp[8]) ? 4'b1000 : 4'b1010;
												assign node2201 = (inp[6]) ? node2209 : node2202;
													assign node2202 = (inp[10]) ? node2204 : 4'b0010;
														assign node2204 = (inp[1]) ? 4'b0000 : node2205;
															assign node2205 = (inp[8]) ? 4'b0000 : 4'b0010;
													assign node2209 = (inp[1]) ? 4'b0000 : node2210;
														assign node2210 = (inp[8]) ? 4'b1000 : 4'b1010;
									assign node2214 = (inp[9]) ? node2216 : 4'b0000;
										assign node2216 = (inp[15]) ? node2256 : node2217;
											assign node2217 = (inp[10]) ? node2235 : node2218;
												assign node2218 = (inp[13]) ? node2224 : node2219;
													assign node2219 = (inp[8]) ? node2221 : 4'b0010;
														assign node2221 = (inp[1]) ? 4'b0010 : 4'b0000;
													assign node2224 = (inp[6]) ? node2230 : node2225;
														assign node2225 = (inp[1]) ? 4'b1010 : node2226;
															assign node2226 = (inp[8]) ? 4'b0010 : 4'b0000;
														assign node2230 = (inp[1]) ? 4'b0000 : node2231;
															assign node2231 = (inp[8]) ? 4'b0000 : 4'b0010;
												assign node2235 = (inp[6]) ? node2245 : node2236;
													assign node2236 = (inp[1]) ? node2242 : node2237;
														assign node2237 = (inp[8]) ? node2239 : 4'b0000;
															assign node2239 = (inp[13]) ? 4'b0010 : 4'b0000;
														assign node2242 = (inp[13]) ? 4'b1000 : 4'b0000;
													assign node2245 = (inp[8]) ? node2251 : node2246;
														assign node2246 = (inp[1]) ? node2248 : 4'b0010;
															assign node2248 = (inp[13]) ? 4'b0000 : 4'b0010;
														assign node2251 = (inp[13]) ? 4'b0000 : node2252;
															assign node2252 = (inp[1]) ? 4'b0010 : 4'b0000;
											assign node2256 = (inp[13]) ? node2258 : 4'b0000;
												assign node2258 = (inp[6]) ? node2266 : node2259;
													assign node2259 = (inp[10]) ? 4'b0000 : node2260;
														assign node2260 = (inp[1]) ? 4'b0010 : node2261;
															assign node2261 = (inp[8]) ? 4'b0000 : 4'b0010;
													assign node2266 = (inp[1]) ? 4'b0000 : node2267;
														assign node2267 = (inp[8]) ? 4'b0000 : 4'b0010;

endmodule