module dtc_split125_bm39 (
	input  wire [14-1:0] inp,
	output wire [14-1:0] outp
);

	wire [14-1:0] node1;
	wire [14-1:0] node3;
	wire [14-1:0] node4;
	wire [14-1:0] node5;
	wire [14-1:0] node6;
	wire [14-1:0] node7;
	wire [14-1:0] node8;
	wire [14-1:0] node9;
	wire [14-1:0] node10;
	wire [14-1:0] node11;
	wire [14-1:0] node16;
	wire [14-1:0] node17;
	wire [14-1:0] node19;
	wire [14-1:0] node20;
	wire [14-1:0] node24;
	wire [14-1:0] node27;
	wire [14-1:0] node28;
	wire [14-1:0] node30;
	wire [14-1:0] node31;
	wire [14-1:0] node34;
	wire [14-1:0] node35;
	wire [14-1:0] node39;
	wire [14-1:0] node40;
	wire [14-1:0] node42;
	wire [14-1:0] node46;
	wire [14-1:0] node47;
	wire [14-1:0] node48;
	wire [14-1:0] node49;
	wire [14-1:0] node50;
	wire [14-1:0] node52;
	wire [14-1:0] node56;
	wire [14-1:0] node57;
	wire [14-1:0] node60;
	wire [14-1:0] node61;
	wire [14-1:0] node65;
	wire [14-1:0] node67;
	wire [14-1:0] node70;
	wire [14-1:0] node71;
	wire [14-1:0] node72;
	wire [14-1:0] node73;
	wire [14-1:0] node77;
	wire [14-1:0] node79;
	wire [14-1:0] node80;
	wire [14-1:0] node84;
	wire [14-1:0] node85;
	wire [14-1:0] node86;
	wire [14-1:0] node87;
	wire [14-1:0] node90;
	wire [14-1:0] node91;
	wire [14-1:0] node95;
	wire [14-1:0] node99;
	wire [14-1:0] node100;
	wire [14-1:0] node101;
	wire [14-1:0] node102;
	wire [14-1:0] node103;
	wire [14-1:0] node104;
	wire [14-1:0] node106;
	wire [14-1:0] node109;
	wire [14-1:0] node112;
	wire [14-1:0] node113;
	wire [14-1:0] node117;
	wire [14-1:0] node118;
	wire [14-1:0] node120;
	wire [14-1:0] node123;
	wire [14-1:0] node124;
	wire [14-1:0] node127;
	wire [14-1:0] node131;
	wire [14-1:0] node133;
	wire [14-1:0] node134;
	wire [14-1:0] node135;
	wire [14-1:0] node137;
	wire [14-1:0] node138;
	wire [14-1:0] node142;
	wire [14-1:0] node144;
	wire [14-1:0] node148;
	wire [14-1:0] node149;
	wire [14-1:0] node150;
	wire [14-1:0] node151;
	wire [14-1:0] node152;
	wire [14-1:0] node155;
	wire [14-1:0] node156;
	wire [14-1:0] node157;
	wire [14-1:0] node158;
	wire [14-1:0] node163;
	wire [14-1:0] node166;
	wire [14-1:0] node167;
	wire [14-1:0] node168;
	wire [14-1:0] node169;
	wire [14-1:0] node171;
	wire [14-1:0] node175;
	wire [14-1:0] node176;
	wire [14-1:0] node180;
	wire [14-1:0] node181;
	wire [14-1:0] node184;
	wire [14-1:0] node186;
	wire [14-1:0] node187;
	wire [14-1:0] node191;
	wire [14-1:0] node192;
	wire [14-1:0] node193;
	wire [14-1:0] node195;
	wire [14-1:0] node196;
	wire [14-1:0] node197;
	wire [14-1:0] node200;
	wire [14-1:0] node207;
	wire [14-1:0] node208;
	wire [14-1:0] node209;
	wire [14-1:0] node210;
	wire [14-1:0] node211;
	wire [14-1:0] node212;
	wire [14-1:0] node213;
	wire [14-1:0] node216;
	wire [14-1:0] node219;
	wire [14-1:0] node220;
	wire [14-1:0] node222;
	wire [14-1:0] node223;
	wire [14-1:0] node227;
	wire [14-1:0] node230;
	wire [14-1:0] node231;
	wire [14-1:0] node232;
	wire [14-1:0] node233;
	wire [14-1:0] node234;
	wire [14-1:0] node237;
	wire [14-1:0] node241;
	wire [14-1:0] node242;
	wire [14-1:0] node247;
	wire [14-1:0] node248;
	wire [14-1:0] node249;
	wire [14-1:0] node250;
	wire [14-1:0] node251;
	wire [14-1:0] node254;
	wire [14-1:0] node255;
	wire [14-1:0] node259;
	wire [14-1:0] node260;
	wire [14-1:0] node264;
	wire [14-1:0] node265;
	wire [14-1:0] node267;
	wire [14-1:0] node272;
	wire [14-1:0] node273;
	wire [14-1:0] node274;
	wire [14-1:0] node275;
	wire [14-1:0] node276;
	wire [14-1:0] node279;
	wire [14-1:0] node280;
	wire [14-1:0] node283;
	wire [14-1:0] node287;
	wire [14-1:0] node288;
	wire [14-1:0] node289;
	wire [14-1:0] node291;
	wire [14-1:0] node296;
	wire [14-1:0] node298;
	wire [14-1:0] node299;
	wire [14-1:0] node300;
	wire [14-1:0] node305;
	wire [14-1:0] node306;
	wire [14-1:0] node307;
	wire [14-1:0] node308;
	wire [14-1:0] node309;
	wire [14-1:0] node311;
	wire [14-1:0] node318;
	wire [14-1:0] node319;
	wire [14-1:0] node320;
	wire [14-1:0] node321;
	wire [14-1:0] node322;
	wire [14-1:0] node323;
	wire [14-1:0] node324;
	wire [14-1:0] node325;
	wire [14-1:0] node326;
	wire [14-1:0] node329;
	wire [14-1:0] node330;
	wire [14-1:0] node332;
	wire [14-1:0] node335;
	wire [14-1:0] node336;
	wire [14-1:0] node337;
	wire [14-1:0] node342;
	wire [14-1:0] node343;
	wire [14-1:0] node345;
	wire [14-1:0] node348;
	wire [14-1:0] node349;
	wire [14-1:0] node352;
	wire [14-1:0] node355;
	wire [14-1:0] node356;
	wire [14-1:0] node357;
	wire [14-1:0] node358;
	wire [14-1:0] node359;
	wire [14-1:0] node363;
	wire [14-1:0] node365;
	wire [14-1:0] node370;
	wire [14-1:0] node371;
	wire [14-1:0] node372;
	wire [14-1:0] node373;
	wire [14-1:0] node375;
	wire [14-1:0] node379;
	wire [14-1:0] node381;
	wire [14-1:0] node382;
	wire [14-1:0] node385;
	wire [14-1:0] node388;
	wire [14-1:0] node389;
	wire [14-1:0] node390;
	wire [14-1:0] node391;
	wire [14-1:0] node395;
	wire [14-1:0] node396;
	wire [14-1:0] node399;
	wire [14-1:0] node400;
	wire [14-1:0] node403;
	wire [14-1:0] node406;
	wire [14-1:0] node407;
	wire [14-1:0] node409;
	wire [14-1:0] node412;
	wire [14-1:0] node413;
	wire [14-1:0] node416;
	wire [14-1:0] node418;
	wire [14-1:0] node421;
	wire [14-1:0] node422;
	wire [14-1:0] node423;
	wire [14-1:0] node424;
	wire [14-1:0] node425;
	wire [14-1:0] node428;
	wire [14-1:0] node430;
	wire [14-1:0] node432;
	wire [14-1:0] node435;
	wire [14-1:0] node436;
	wire [14-1:0] node437;
	wire [14-1:0] node440;
	wire [14-1:0] node443;
	wire [14-1:0] node444;
	wire [14-1:0] node447;
	wire [14-1:0] node448;
	wire [14-1:0] node449;
	wire [14-1:0] node453;
	wire [14-1:0] node454;
	wire [14-1:0] node457;
	wire [14-1:0] node460;
	wire [14-1:0] node461;
	wire [14-1:0] node462;
	wire [14-1:0] node465;
	wire [14-1:0] node467;
	wire [14-1:0] node471;
	wire [14-1:0] node472;
	wire [14-1:0] node473;
	wire [14-1:0] node474;
	wire [14-1:0] node477;
	wire [14-1:0] node480;
	wire [14-1:0] node481;
	wire [14-1:0] node483;
	wire [14-1:0] node488;
	wire [14-1:0] node489;
	wire [14-1:0] node490;
	wire [14-1:0] node491;
	wire [14-1:0] node492;
	wire [14-1:0] node494;
	wire [14-1:0] node497;
	wire [14-1:0] node498;
	wire [14-1:0] node500;
	wire [14-1:0] node504;
	wire [14-1:0] node505;
	wire [14-1:0] node506;
	wire [14-1:0] node507;
	wire [14-1:0] node510;
	wire [14-1:0] node511;
	wire [14-1:0] node516;
	wire [14-1:0] node517;
	wire [14-1:0] node518;
	wire [14-1:0] node521;
	wire [14-1:0] node523;
	wire [14-1:0] node527;
	wire [14-1:0] node528;
	wire [14-1:0] node529;
	wire [14-1:0] node530;
	wire [14-1:0] node533;
	wire [14-1:0] node534;
	wire [14-1:0] node535;
	wire [14-1:0] node539;
	wire [14-1:0] node542;
	wire [14-1:0] node543;
	wire [14-1:0] node544;
	wire [14-1:0] node546;
	wire [14-1:0] node550;
	wire [14-1:0] node552;
	wire [14-1:0] node554;
	wire [14-1:0] node557;
	wire [14-1:0] node558;
	wire [14-1:0] node559;
	wire [14-1:0] node560;
	wire [14-1:0] node563;
	wire [14-1:0] node566;
	wire [14-1:0] node568;
	wire [14-1:0] node569;
	wire [14-1:0] node574;
	wire [14-1:0] node575;
	wire [14-1:0] node576;
	wire [14-1:0] node577;
	wire [14-1:0] node578;
	wire [14-1:0] node579;
	wire [14-1:0] node582;
	wire [14-1:0] node585;
	wire [14-1:0] node586;
	wire [14-1:0] node590;
	wire [14-1:0] node591;
	wire [14-1:0] node592;
	wire [14-1:0] node595;
	wire [14-1:0] node599;
	wire [14-1:0] node600;
	wire [14-1:0] node602;
	wire [14-1:0] node603;
	wire [14-1:0] node608;
	wire [14-1:0] node609;
	wire [14-1:0] node611;
	wire [14-1:0] node612;
	wire [14-1:0] node617;
	wire [14-1:0] node618;
	wire [14-1:0] node619;
	wire [14-1:0] node620;
	wire [14-1:0] node621;
	wire [14-1:0] node622;
	wire [14-1:0] node623;
	wire [14-1:0] node624;
	wire [14-1:0] node628;
	wire [14-1:0] node629;
	wire [14-1:0] node632;
	wire [14-1:0] node635;
	wire [14-1:0] node636;
	wire [14-1:0] node637;
	wire [14-1:0] node640;
	wire [14-1:0] node642;
	wire [14-1:0] node646;
	wire [14-1:0] node647;
	wire [14-1:0] node648;
	wire [14-1:0] node652;
	wire [14-1:0] node653;
	wire [14-1:0] node655;
	wire [14-1:0] node659;
	wire [14-1:0] node660;
	wire [14-1:0] node661;
	wire [14-1:0] node662;
	wire [14-1:0] node663;
	wire [14-1:0] node667;
	wire [14-1:0] node668;
	wire [14-1:0] node671;
	wire [14-1:0] node674;
	wire [14-1:0] node675;
	wire [14-1:0] node677;
	wire [14-1:0] node681;
	wire [14-1:0] node683;
	wire [14-1:0] node685;
	wire [14-1:0] node688;
	wire [14-1:0] node690;
	wire [14-1:0] node691;
	wire [14-1:0] node692;
	wire [14-1:0] node693;
	wire [14-1:0] node695;
	wire [14-1:0] node698;
	wire [14-1:0] node701;
	wire [14-1:0] node702;
	wire [14-1:0] node706;
	wire [14-1:0] node707;
	wire [14-1:0] node708;
	wire [14-1:0] node710;
	wire [14-1:0] node715;
	wire [14-1:0] node716;
	wire [14-1:0] node717;
	wire [14-1:0] node718;
	wire [14-1:0] node720;
	wire [14-1:0] node721;
	wire [14-1:0] node722;
	wire [14-1:0] node726;
	wire [14-1:0] node727;
	wire [14-1:0] node730;
	wire [14-1:0] node733;
	wire [14-1:0] node734;
	wire [14-1:0] node735;
	wire [14-1:0] node737;
	wire [14-1:0] node740;
	wire [14-1:0] node743;
	wire [14-1:0] node745;
	wire [14-1:0] node746;
	wire [14-1:0] node750;
	wire [14-1:0] node751;
	wire [14-1:0] node752;
	wire [14-1:0] node758;
	wire [14-1:0] node759;
	wire [14-1:0] node760;
	wire [14-1:0] node761;
	wire [14-1:0] node762;
	wire [14-1:0] node763;
	wire [14-1:0] node764;
	wire [14-1:0] node765;
	wire [14-1:0] node767;
	wire [14-1:0] node768;
	wire [14-1:0] node773;
	wire [14-1:0] node774;
	wire [14-1:0] node775;
	wire [14-1:0] node778;
	wire [14-1:0] node782;
	wire [14-1:0] node783;
	wire [14-1:0] node784;
	wire [14-1:0] node787;
	wire [14-1:0] node788;
	wire [14-1:0] node790;
	wire [14-1:0] node796;
	wire [14-1:0] node797;
	wire [14-1:0] node798;
	wire [14-1:0] node799;
	wire [14-1:0] node800;
	wire [14-1:0] node801;
	wire [14-1:0] node804;
	wire [14-1:0] node805;
	wire [14-1:0] node810;
	wire [14-1:0] node811;
	wire [14-1:0] node812;
	wire [14-1:0] node814;
	wire [14-1:0] node818;
	wire [14-1:0] node819;
	wire [14-1:0] node823;
	wire [14-1:0] node824;
	wire [14-1:0] node825;
	wire [14-1:0] node827;
	wire [14-1:0] node829;
	wire [14-1:0] node832;
	wire [14-1:0] node833;
	wire [14-1:0] node835;
	wire [14-1:0] node839;
	wire [14-1:0] node840;
	wire [14-1:0] node841;
	wire [14-1:0] node843;
	wire [14-1:0] node848;
	wire [14-1:0] node849;
	wire [14-1:0] node850;
	wire [14-1:0] node851;
	wire [14-1:0] node853;
	wire [14-1:0] node856;
	wire [14-1:0] node860;
	wire [14-1:0] node861;
	wire [14-1:0] node862;
	wire [14-1:0] node864;
	wire [14-1:0] node869;
	wire [14-1:0] node870;
	wire [14-1:0] node871;
	wire [14-1:0] node872;
	wire [14-1:0] node873;
	wire [14-1:0] node874;
	wire [14-1:0] node876;
	wire [14-1:0] node879;
	wire [14-1:0] node881;
	wire [14-1:0] node884;
	wire [14-1:0] node886;
	wire [14-1:0] node888;
	wire [14-1:0] node889;
	wire [14-1:0] node893;
	wire [14-1:0] node894;
	wire [14-1:0] node896;
	wire [14-1:0] node900;
	wire [14-1:0] node902;
	wire [14-1:0] node904;
	wire [14-1:0] node905;
	wire [14-1:0] node906;
	wire [14-1:0] node912;
	wire [14-1:0] node913;
	wire [14-1:0] node914;
	wire [14-1:0] node915;
	wire [14-1:0] node916;
	wire [14-1:0] node917;
	wire [14-1:0] node918;
	wire [14-1:0] node919;
	wire [14-1:0] node920;
	wire [14-1:0] node924;
	wire [14-1:0] node927;
	wire [14-1:0] node929;
	wire [14-1:0] node931;
	wire [14-1:0] node934;
	wire [14-1:0] node935;
	wire [14-1:0] node937;
	wire [14-1:0] node941;
	wire [14-1:0] node943;
	wire [14-1:0] node944;
	wire [14-1:0] node946;
	wire [14-1:0] node947;
	wire [14-1:0] node952;
	wire [14-1:0] node953;
	wire [14-1:0] node954;
	wire [14-1:0] node956;
	wire [14-1:0] node957;
	wire [14-1:0] node958;
	wire [14-1:0] node962;
	wire [14-1:0] node965;
	wire [14-1:0] node967;
	wire [14-1:0] node971;
	wire [14-1:0] node972;
	wire [14-1:0] node973;
	wire [14-1:0] node975;
	wire [14-1:0] node976;
	wire [14-1:0] node982;
	wire [14-1:0] node984;
	wire [14-1:0] node986;
	wire [14-1:0] node987;
	wire [14-1:0] node989;

	assign outp = (inp[8]) ? node318 : node1;
		assign node1 = (inp[13]) ? node3 : 14'b00000000000000;
			assign node3 = (inp[1]) ? node207 : node4;
				assign node4 = (inp[10]) ? node148 : node5;
					assign node5 = (inp[3]) ? node99 : node6;
						assign node6 = (inp[6]) ? node46 : node7;
							assign node7 = (inp[0]) ? node27 : node8;
								assign node8 = (inp[9]) ? node16 : node9;
									assign node9 = (inp[2]) ? 14'b00000000000001 : node10;
										assign node10 = (inp[4]) ? 14'b00000000000001 : node11;
											assign node11 = (inp[11]) ? 14'b00000000000001 : 14'b10000000001000;
									assign node16 = (inp[7]) ? node24 : node17;
										assign node17 = (inp[2]) ? node19 : 14'b01000000000100;
											assign node19 = (inp[12]) ? 14'b01000100000000 : node20;
												assign node20 = (inp[11]) ? 14'b01000000000010 : 14'b01000100000010;
										assign node24 = (inp[2]) ? 14'b00000000000001 : 14'b00000000000110;
								assign node27 = (inp[4]) ? node39 : node28;
									assign node28 = (inp[9]) ? node30 : 14'b01000010110000;
										assign node30 = (inp[5]) ? node34 : node31;
											assign node31 = (inp[12]) ? 14'b01000010010100 : 14'b01100010010110;
											assign node34 = (inp[2]) ? 14'b01000110010010 : node35;
												assign node35 = (inp[7]) ? 14'b01000010010110 : 14'b01000110010110;
									assign node39 = (inp[2]) ? 14'b00000000000001 : node40;
										assign node40 = (inp[11]) ? node42 : 14'b00100110010110;
											assign node42 = (inp[7]) ? 14'b00000010110110 : 14'b00000110110110;
							assign node46 = (inp[0]) ? node70 : node47;
								assign node47 = (inp[9]) ? node65 : node48;
									assign node48 = (inp[11]) ? node56 : node49;
										assign node49 = (inp[4]) ? 14'b00000000000001 : node50;
											assign node50 = (inp[2]) ? node52 : 14'b00000000000001;
												assign node52 = (inp[5]) ? 14'b01010100110010 : 14'b01110000110110;
										assign node56 = (inp[5]) ? node60 : node57;
											assign node57 = (inp[7]) ? 14'b01110000110100 : 14'b01110100110100;
											assign node60 = (inp[7]) ? 14'b01010000110000 : node61;
												assign node61 = (inp[4]) ? 14'b01010000110010 : 14'b01010100110010;
									assign node65 = (inp[4]) ? node67 : 14'b01110100010110;
										assign node67 = (inp[2]) ? 14'b01010000010010 : 14'b00010100010110;
								assign node70 = (inp[7]) ? node84 : node71;
									assign node71 = (inp[9]) ? node77 : node72;
										assign node72 = (inp[4]) ? 14'b00000100110110 : node73;
											assign node73 = (inp[12]) ? 14'b01100100110100 : 14'b01100100110110;
										assign node77 = (inp[12]) ? node79 : 14'b00000000000001;
											assign node79 = (inp[11]) ? 14'b01000100010100 : node80;
												assign node80 = (inp[5]) ? 14'b00000000000001 : 14'b00100100010100;
									assign node84 = (inp[2]) ? 14'b00000000000001 : node85;
										assign node85 = (inp[12]) ? node95 : node86;
											assign node86 = (inp[5]) ? node90 : node87;
												assign node87 = (inp[11]) ? 14'b00000000110010 : 14'b00000000010010;
												assign node90 = (inp[11]) ? 14'b00000000010110 : node91;
													assign node91 = (inp[4]) ? 14'b00000000110110 : 14'b01000000110110;
											assign node95 = (inp[5]) ? 14'b00000000000001 : 14'b00000000010000;
						assign node99 = (inp[6]) ? node131 : node100;
							assign node100 = (inp[0]) ? 14'b00000000000001 : node101;
								assign node101 = (inp[12]) ? node117 : node102;
									assign node102 = (inp[9]) ? node112 : node103;
										assign node103 = (inp[2]) ? node109 : node104;
											assign node104 = (inp[7]) ? node106 : 14'b00010110110110;
												assign node106 = (inp[5]) ? 14'b00010010110110 : 14'b00010010110010;
											assign node109 = (inp[11]) ? 14'b00000000000001 : 14'b01010010110010;
										assign node112 = (inp[2]) ? 14'b01110110010110 : node113;
											assign node113 = (inp[11]) ? 14'b00110010010110 : 14'b00010010010010;
									assign node117 = (inp[4]) ? node123 : node118;
										assign node118 = (inp[2]) ? node120 : 14'b01010110010100;
											assign node120 = (inp[9]) ? 14'b01010010010000 : 14'b01010110110000;
										assign node123 = (inp[11]) ? node127 : node124;
											assign node124 = (inp[2]) ? 14'b00000000000001 : 14'b00010010010100;
											assign node127 = (inp[9]) ? 14'b00010110010100 : 14'b00010110110100;
							assign node131 = (inp[0]) ? node133 : 14'b00000000000001;
								assign node133 = (inp[9]) ? 14'b00000000000001 : node134;
									assign node134 = (inp[4]) ? node142 : node135;
										assign node135 = (inp[11]) ? node137 : 14'b01000000100000;
											assign node137 = (inp[7]) ? 14'b01100000100110 : node138;
												assign node138 = (inp[5]) ? 14'b01000100100110 : 14'b01100100100100;
										assign node142 = (inp[12]) ? node144 : 14'b00000000000001;
											assign node144 = (inp[11]) ? 14'b00100100100100 : 14'b00000000100100;
					assign node148 = (inp[5]) ? 14'b00000000000001 : node149;
						assign node149 = (inp[2]) ? node191 : node150;
							assign node150 = (inp[12]) ? node166 : node151;
								assign node151 = (inp[0]) ? node155 : node152;
									assign node152 = (inp[9]) ? 14'b00110000010010 : 14'b00000000000001;
									assign node155 = (inp[7]) ? node163 : node156;
										assign node156 = (inp[3]) ? 14'b01100100100010 : node157;
											assign node157 = (inp[6]) ? 14'b00100100110010 : node158;
												assign node158 = (inp[4]) ? 14'b00100110110010 : 14'b01100110110010;
										assign node163 = (inp[6]) ? 14'b01100000010010 : 14'b01100010110010;
								assign node166 = (inp[3]) ? node180 : node167;
									assign node167 = (inp[6]) ? node175 : node168;
										assign node168 = (inp[0]) ? 14'b01100110110000 : node169;
											assign node169 = (inp[9]) ? node171 : 14'b00000000000001;
												assign node171 = (inp[4]) ? 14'b00100100000000 : 14'b01100100000000;
										assign node175 = (inp[9]) ? 14'b01100000010000 : node176;
											assign node176 = (inp[11]) ? 14'b01110000110000 : 14'b01110100110000;
									assign node180 = (inp[6]) ? node184 : node181;
										assign node181 = (inp[0]) ? 14'b00000000000001 : 14'b00110010010000;
										assign node184 = (inp[0]) ? node186 : 14'b00000000000001;
											assign node186 = (inp[7]) ? 14'b00100000100000 : node187;
												assign node187 = (inp[4]) ? 14'b00100100100000 : 14'b01100100100000;
							assign node191 = (inp[0]) ? 14'b00000000000001 : node192;
								assign node192 = (inp[7]) ? 14'b00000000000001 : node193;
									assign node193 = (inp[4]) ? node195 : 14'b00000000000001;
										assign node195 = (inp[11]) ? 14'b00000100000000 : node196;
											assign node196 = (inp[9]) ? node200 : node197;
												assign node197 = (inp[12]) ? 14'b00010100110000 : 14'b00010100110010;
												assign node200 = (inp[6]) ? 14'b00010100010010 : 14'b00010110010010;
				assign node207 = (inp[0]) ? node305 : node208;
					assign node208 = (inp[2]) ? node272 : node209;
						assign node209 = (inp[3]) ? node247 : node210;
							assign node210 = (inp[5]) ? node230 : node211;
								assign node211 = (inp[7]) ? node219 : node212;
									assign node212 = (inp[6]) ? node216 : node213;
										assign node213 = (inp[4]) ? 14'b00110110000010 : 14'b01110110000010;
										assign node216 = (inp[12]) ? 14'b01110100000000 : 14'b00110100000110;
									assign node219 = (inp[6]) ? node227 : node220;
										assign node220 = (inp[4]) ? node222 : 14'b00010010000010;
											assign node222 = (inp[9]) ? 14'b00110010000100 : node223;
												assign node223 = (inp[10]) ? 14'b00110010100000 : 14'b00110010100100;
										assign node227 = (inp[4]) ? 14'b00110000100110 : 14'b01110000100000;
								assign node230 = (inp[10]) ? 14'b00000000000001 : node231;
									assign node231 = (inp[12]) ? node241 : node232;
										assign node232 = (inp[4]) ? 14'b00010000100110 : node233;
											assign node233 = (inp[7]) ? node237 : node234;
												assign node234 = (inp[11]) ? 14'b01010100000110 : 14'b01010110000110;
												assign node237 = (inp[6]) ? 14'b01010000000110 : 14'b01010010000110;
										assign node241 = (inp[11]) ? 14'b00000000000001 : node242;
											assign node242 = (inp[4]) ? 14'b00010010000100 : 14'b01010110000100;
							assign node247 = (inp[6]) ? 14'b00000000000001 : node248;
								assign node248 = (inp[5]) ? node264 : node249;
									assign node249 = (inp[9]) ? node259 : node250;
										assign node250 = (inp[10]) ? node254 : node251;
											assign node251 = (inp[12]) ? 14'b01000010100100 : 14'b00000000000001;
											assign node254 = (inp[7]) ? 14'b00100010100000 : node255;
												assign node255 = (inp[11]) ? 14'b01100110100000 : 14'b01100110100010;
										assign node259 = (inp[12]) ? 14'b00100110000000 : node260;
											assign node260 = (inp[10]) ? 14'b01100110000010 : 14'b00100110000110;
									assign node264 = (inp[10]) ? 14'b00000000000001 : node265;
										assign node265 = (inp[9]) ? node267 : 14'b01000010100110;
											assign node267 = (inp[12]) ? 14'b00000010000100 : 14'b00000010000110;
						assign node272 = (inp[10]) ? node296 : node273;
							assign node273 = (inp[7]) ? node287 : node274;
								assign node274 = (inp[6]) ? 14'b00000000000001 : node275;
									assign node275 = (inp[12]) ? node279 : node276;
										assign node276 = (inp[5]) ? 14'b01000010000010 : 14'b00000000000001;
										assign node279 = (inp[3]) ? node283 : node280;
											assign node280 = (inp[4]) ? 14'b00010110100100 : 14'b01110110100100;
											assign node283 = (inp[11]) ? 14'b00000110000100 : 14'b01000110100000;
								assign node287 = (inp[4]) ? 14'b00000000000001 : node288;
									assign node288 = (inp[3]) ? 14'b00000000000001 : node289;
										assign node289 = (inp[6]) ? node291 : 14'b00000000000001;
											assign node291 = (inp[9]) ? 14'b01110000000110 : 14'b01010000100000;
							assign node296 = (inp[4]) ? node298 : 14'b00000000000001;
								assign node298 = (inp[7]) ? 14'b00000000000001 : node299;
									assign node299 = (inp[5]) ? 14'b00000000000001 : node300;
										assign node300 = (inp[6]) ? 14'b00000000000001 : 14'b00010110000010;
					assign node305 = (inp[6]) ? 14'b00000000000001 : node306;
						assign node306 = (inp[11]) ? 14'b00000000000001 : node307;
							assign node307 = (inp[12]) ? 14'b00000000000001 : node308;
								assign node308 = (inp[4]) ? 14'b00000000000001 : node309;
									assign node309 = (inp[3]) ? node311 : 14'b00000000000001;
										assign node311 = (inp[10]) ? 14'b00000000000001 : 14'b10000000000010;
		assign node318 = (inp[0]) ? node758 : node319;
			assign node319 = (inp[3]) ? node617 : node320;
				assign node320 = (inp[12]) ? node488 : node321;
					assign node321 = (inp[2]) ? node421 : node322;
						assign node322 = (inp[13]) ? node370 : node323;
							assign node323 = (inp[11]) ? node355 : node324;
								assign node324 = (inp[4]) ? node342 : node325;
									assign node325 = (inp[5]) ? node329 : node326;
										assign node326 = (inp[10]) ? 14'b01101000000010 : 14'b00000000000001;
										assign node329 = (inp[6]) ? node335 : node330;
											assign node330 = (inp[9]) ? node332 : 14'b01110010000010;
												assign node332 = (inp[1]) ? 14'b00100000000010 : 14'b01100100000010;
											assign node335 = (inp[7]) ? 14'b01100000110010 : node336;
												assign node336 = (inp[1]) ? 14'b00110000110010 : node337;
													assign node337 = (inp[10]) ? 14'b01110100110010 : 14'b00110100110010;
									assign node342 = (inp[7]) ? node348 : node343;
										assign node343 = (inp[5]) ? node345 : 14'b01111100110000;
											assign node345 = (inp[1]) ? 14'b01110000010000 : 14'b01110100010000;
										assign node348 = (inp[10]) ? node352 : node349;
											assign node349 = (inp[9]) ? 14'b01101010010110 : 14'b01100010110110;
											assign node352 = (inp[5]) ? 14'b01100110010000 : 14'b01101010110000;
								assign node355 = (inp[10]) ? 14'b00000000000001 : node356;
									assign node356 = (inp[4]) ? 14'b00000000000001 : node357;
										assign node357 = (inp[7]) ? node363 : node358;
											assign node358 = (inp[1]) ? 14'b01110010000100 : node359;
												assign node359 = (inp[5]) ? 14'b01110100010100 : 14'b01111100010100;
											assign node363 = (inp[1]) ? node365 : 14'b01101110110100;
												assign node365 = (inp[5]) ? 14'b01100010110100 : 14'b01101010110100;
							assign node370 = (inp[6]) ? node388 : node371;
								assign node371 = (inp[5]) ? node379 : node372;
									assign node372 = (inp[11]) ? 14'b00000000000001 : node373;
										assign node373 = (inp[9]) ? node375 : 14'b00010010100000;
											assign node375 = (inp[7]) ? 14'b00100000000100 : 14'b00000000000001;
									assign node379 = (inp[1]) ? node381 : 14'b00000000000001;
										assign node381 = (inp[9]) ? node385 : node382;
											assign node382 = (inp[7]) ? 14'b00110010100000 : 14'b01110110100000;
											assign node385 = (inp[7]) ? 14'b01110010000000 : 14'b01110110000000;
								assign node388 = (inp[9]) ? node406 : node389;
									assign node389 = (inp[4]) ? node395 : node390;
										assign node390 = (inp[7]) ? 14'b01110000110000 : node391;
											assign node391 = (inp[1]) ? 14'b01110100100000 : 14'b01110100110000;
										assign node395 = (inp[1]) ? node399 : node396;
											assign node396 = (inp[7]) ? 14'b00110000110100 : 14'b00110100110100;
											assign node399 = (inp[5]) ? node403 : node400;
												assign node400 = (inp[7]) ? 14'b00110000100100 : 14'b00110100100100;
												assign node403 = (inp[7]) ? 14'b00110000100000 : 14'b00110100100000;
									assign node406 = (inp[1]) ? node412 : node407;
										assign node407 = (inp[4]) ? node409 : 14'b01110100010000;
											assign node409 = (inp[7]) ? 14'b00110000010100 : 14'b00110100010100;
										assign node412 = (inp[5]) ? node416 : node413;
											assign node413 = (inp[10]) ? 14'b00000000000001 : 14'b00010000000000;
											assign node416 = (inp[4]) ? node418 : 14'b01110000000000;
												assign node418 = (inp[7]) ? 14'b00110000000000 : 14'b00110100000000;
						assign node421 = (inp[11]) ? node471 : node422;
							assign node422 = (inp[13]) ? node460 : node423;
								assign node423 = (inp[9]) ? node435 : node424;
									assign node424 = (inp[10]) ? node428 : node425;
										assign node425 = (inp[7]) ? 14'b00001100110000 : 14'b00011100110000;
										assign node428 = (inp[5]) ? node430 : 14'b00000000000001;
											assign node430 = (inp[7]) ? node432 : 14'b00000000000001;
												assign node432 = (inp[6]) ? 14'b00100100110000 : 14'b00100110110000;
									assign node435 = (inp[5]) ? node443 : node436;
										assign node436 = (inp[7]) ? node440 : node437;
											assign node437 = (inp[1]) ? 14'b00011000010000 : 14'b00111100010010;
											assign node440 = (inp[6]) ? 14'b00101100010110 : 14'b00101010010110;
										assign node443 = (inp[1]) ? node447 : node444;
											assign node444 = (inp[10]) ? 14'b00000000000001 : 14'b00000100000000;
											assign node447 = (inp[10]) ? node453 : node448;
												assign node448 = (inp[6]) ? 14'b00110000010110 : node449;
													assign node449 = (inp[7]) ? 14'b00100010010110 : 14'b00100000000110;
												assign node453 = (inp[7]) ? node457 : node454;
													assign node454 = (inp[6]) ? 14'b00110000010000 : 14'b00100000000000;
													assign node457 = (inp[6]) ? 14'b00100000010000 : 14'b00100010010000;
								assign node460 = (inp[7]) ? 14'b00000000000001 : node461;
									assign node461 = (inp[5]) ? node465 : node462;
										assign node462 = (inp[10]) ? 14'b01100100000100 : 14'b01110100100100;
										assign node465 = (inp[9]) ? node467 : 14'b00010110100000;
											assign node467 = (inp[4]) ? 14'b00000100000000 : 14'b00000000000001;
							assign node471 = (inp[4]) ? 14'b00000000000001 : node472;
								assign node472 = (inp[10]) ? node480 : node473;
									assign node473 = (inp[6]) ? node477 : node474;
										assign node474 = (inp[5]) ? 14'b00100100000100 : 14'b00101100000100;
										assign node477 = (inp[1]) ? 14'b00110000010100 : 14'b01110000010100;
									assign node480 = (inp[5]) ? 14'b00000000000001 : node481;
										assign node481 = (inp[13]) ? node483 : 14'b00000000000001;
											assign node483 = (inp[6]) ? 14'b01110000010100 : 14'b01100100000100;
					assign node488 = (inp[5]) ? node574 : node489;
						assign node489 = (inp[13]) ? node527 : node490;
							assign node490 = (inp[6]) ? node504 : node491;
								assign node491 = (inp[11]) ? node497 : node492;
									assign node492 = (inp[1]) ? node494 : 14'b00000000000001;
										assign node494 = (inp[7]) ? 14'b00001010110110 : 14'b00011010000010;
									assign node497 = (inp[10]) ? 14'b00000000000001 : node498;
										assign node498 = (inp[7]) ? node500 : 14'b00000000000001;
											assign node500 = (inp[2]) ? 14'b00000000000001 : 14'b01001110110000;
								assign node504 = (inp[11]) ? node516 : node505;
									assign node505 = (inp[4]) ? 14'b00000000000001 : node506;
										assign node506 = (inp[1]) ? node510 : node507;
											assign node507 = (inp[2]) ? 14'b00011100010110 : 14'b01011100010010;
											assign node510 = (inp[7]) ? 14'b00001000010010 : node511;
												assign node511 = (inp[2]) ? 14'b00011000110010 : 14'b01011000110010;
									assign node516 = (inp[10]) ? 14'b00000000000001 : node517;
										assign node517 = (inp[9]) ? node521 : node518;
											assign node518 = (inp[7]) ? 14'b01001000110100 : 14'b00011000110100;
											assign node521 = (inp[7]) ? node523 : 14'b01011000010000;
												assign node523 = (inp[4]) ? 14'b01001100010000 : 14'b01001100010100;
							assign node527 = (inp[4]) ? node557 : node528;
								assign node528 = (inp[1]) ? node542 : node529;
									assign node529 = (inp[6]) ? node533 : node530;
										assign node530 = (inp[9]) ? 14'b01000100000000 : 14'b00000000000001;
										assign node533 = (inp[7]) ? node539 : node534;
											assign node534 = (inp[9]) ? 14'b01010100010000 : node535;
												assign node535 = (inp[11]) ? 14'b01010100110000 : 14'b01010100110100;
											assign node539 = (inp[2]) ? 14'b01010000010000 : 14'b01010000010100;
									assign node542 = (inp[9]) ? node550 : node543;
										assign node543 = (inp[6]) ? 14'b01010100100000 : node544;
											assign node544 = (inp[7]) ? node546 : 14'b01010110100100;
												assign node546 = (inp[2]) ? 14'b01010010100000 : 14'b01010010100100;
										assign node550 = (inp[7]) ? node552 : 14'b01010110000000;
											assign node552 = (inp[2]) ? node554 : 14'b01010010000100;
												assign node554 = (inp[6]) ? 14'b01010000000000 : 14'b01010010000000;
								assign node557 = (inp[2]) ? 14'b00000000000001 : node558;
									assign node558 = (inp[7]) ? node566 : node559;
										assign node559 = (inp[9]) ? node563 : node560;
											assign node560 = (inp[6]) ? 14'b00010100100100 : 14'b00010110100100;
											assign node563 = (inp[11]) ? 14'b00010100000100 : 14'b00000100000100;
										assign node566 = (inp[6]) ? node568 : 14'b00000000000001;
											assign node568 = (inp[9]) ? 14'b00010000000100 : node569;
												assign node569 = (inp[11]) ? 14'b00010000110100 : 14'b00010000100100;
						assign node574 = (inp[13]) ? node608 : node575;
							assign node575 = (inp[10]) ? node599 : node576;
								assign node576 = (inp[2]) ? node590 : node577;
									assign node577 = (inp[11]) ? node585 : node578;
										assign node578 = (inp[7]) ? node582 : node579;
											assign node579 = (inp[4]) ? 14'b01010010000010 : 14'b01000000000110;
											assign node582 = (inp[6]) ? 14'b01000000010010 : 14'b01000010010010;
										assign node585 = (inp[6]) ? 14'b01010100010000 : node586;
											assign node586 = (inp[4]) ? 14'b01000010110000 : 14'b01000010110100;
									assign node590 = (inp[7]) ? 14'b00000000000001 : node591;
										assign node591 = (inp[6]) ? node595 : node592;
											assign node592 = (inp[9]) ? 14'b00000000000100 : 14'b00010010000100;
											assign node595 = (inp[9]) ? 14'b00010000010110 : 14'b00010000110110;
								assign node599 = (inp[4]) ? 14'b00000000000001 : node600;
									assign node600 = (inp[7]) ? node602 : 14'b00000000000001;
										assign node602 = (inp[11]) ? 14'b00000000000001 : node603;
											assign node603 = (inp[9]) ? 14'b00000010010010 : 14'b00000000110010;
							assign node608 = (inp[9]) ? 14'b00000000000001 : node609;
								assign node609 = (inp[2]) ? node611 : 14'b00000000000001;
									assign node611 = (inp[6]) ? 14'b00000000000001 : node612;
										assign node612 = (inp[7]) ? 14'b10001000001000 : 14'b00000000000001;
				assign node617 = (inp[6]) ? node715 : node618;
					assign node618 = (inp[7]) ? node688 : node619;
						assign node619 = (inp[11]) ? node659 : node620;
							assign node620 = (inp[13]) ? node646 : node621;
								assign node621 = (inp[4]) ? node635 : node622;
									assign node622 = (inp[12]) ? node628 : node623;
										assign node623 = (inp[2]) ? 14'b00111010110010 : node624;
											assign node624 = (inp[1]) ? 14'b00110010110010 : 14'b00110110110010;
										assign node628 = (inp[2]) ? node632 : node629;
											assign node629 = (inp[5]) ? 14'b01010110110110 : 14'b01011110110110;
											assign node632 = (inp[1]) ? 14'b00011010010110 : 14'b00011110010110;
									assign node635 = (inp[2]) ? 14'b00000000000001 : node636;
										assign node636 = (inp[10]) ? node640 : node637;
											assign node637 = (inp[1]) ? 14'b01010010010010 : 14'b00000000000001;
											assign node640 = (inp[12]) ? node642 : 14'b01110110110000;
												assign node642 = (inp[1]) ? 14'b00111010010000 : 14'b00111110110000;
								assign node646 = (inp[5]) ? node652 : node647;
									assign node647 = (inp[9]) ? 14'b00000110000100 : node648;
										assign node648 = (inp[4]) ? 14'b00100110100100 : 14'b01100110100100;
									assign node652 = (inp[12]) ? 14'b00000000000001 : node653;
										assign node653 = (inp[4]) ? node655 : 14'b01100110000000;
											assign node655 = (inp[1]) ? 14'b00000110100000 : 14'b00010110110000;
							assign node659 = (inp[10]) ? node681 : node660;
								assign node660 = (inp[4]) ? node674 : node661;
									assign node661 = (inp[13]) ? node667 : node662;
										assign node662 = (inp[9]) ? 14'b01111110010100 : node663;
											assign node663 = (inp[12]) ? 14'b01010010110100 : 14'b01110110110100;
										assign node667 = (inp[5]) ? node671 : node668;
											assign node668 = (inp[1]) ? 14'b01100110100100 : 14'b01110110010100;
											assign node671 = (inp[2]) ? 14'b00000000000001 : 14'b01100110000000;
									assign node674 = (inp[2]) ? 14'b00000000000001 : node675;
										assign node675 = (inp[5]) ? node677 : 14'b00110110010100;
											assign node677 = (inp[12]) ? 14'b01010110110000 : 14'b00000000000001;
								assign node681 = (inp[12]) ? node683 : 14'b00000000000001;
									assign node683 = (inp[13]) ? node685 : 14'b00000000000001;
										assign node685 = (inp[1]) ? 14'b01000110100100 : 14'b00000000000001;
						assign node688 = (inp[13]) ? node690 : 14'b00000000000001;
							assign node690 = (inp[4]) ? node706 : node691;
								assign node691 = (inp[5]) ? node701 : node692;
									assign node692 = (inp[1]) ? node698 : node693;
										assign node693 = (inp[11]) ? node695 : 14'b01110010110100;
											assign node695 = (inp[2]) ? 14'b01010010110000 : 14'b01010010110100;
										assign node698 = (inp[12]) ? 14'b01000010000100 : 14'b01100010000100;
									assign node701 = (inp[12]) ? 14'b00000000000001 : node702;
										assign node702 = (inp[9]) ? 14'b01100010000000 : 14'b01110010110000;
								assign node706 = (inp[2]) ? 14'b00000000000001 : node707;
									assign node707 = (inp[1]) ? 14'b00000000000001 : node708;
										assign node708 = (inp[9]) ? node710 : 14'b00110010110000;
											assign node710 = (inp[10]) ? 14'b00110010010000 : 14'b00110010010100;
					assign node715 = (inp[9]) ? 14'b00000000000001 : node716;
						assign node716 = (inp[13]) ? node750 : node717;
							assign node717 = (inp[7]) ? node733 : node718;
								assign node718 = (inp[1]) ? node720 : 14'b00000000000001;
									assign node720 = (inp[12]) ? node726 : node721;
										assign node721 = (inp[11]) ? 14'b00000000000001 : node722;
											assign node722 = (inp[10]) ? 14'b00000000000001 : 14'b00110000100010;
										assign node726 = (inp[10]) ? node730 : node727;
											assign node727 = (inp[5]) ? 14'b01010000100100 : 14'b00011000100100;
											assign node730 = (inp[11]) ? 14'b00000000000001 : 14'b00111000100000;
								assign node733 = (inp[1]) ? node743 : node734;
									assign node734 = (inp[4]) ? node740 : node735;
										assign node735 = (inp[10]) ? node737 : 14'b01001100100110;
											assign node737 = (inp[12]) ? 14'b00000100100010 : 14'b01100100100010;
										assign node740 = (inp[5]) ? 14'b00100100100000 : 14'b00101100100000;
									assign node743 = (inp[10]) ? node745 : 14'b00001000100100;
										assign node745 = (inp[4]) ? 14'b00000000000001 : node746;
											assign node746 = (inp[12]) ? 14'b00000000000001 : 14'b00101000100010;
							assign node750 = (inp[12]) ? 14'b00000000000001 : node751;
								assign node751 = (inp[10]) ? 14'b00000000000001 : node752;
									assign node752 = (inp[5]) ? 14'b00000000000001 : 14'b10000000000000;
			assign node758 = (inp[1]) ? node912 : node759;
				assign node759 = (inp[3]) ? node869 : node760;
					assign node760 = (inp[13]) ? node796 : node761;
						assign node761 = (inp[7]) ? 14'b00000000000001 : node762;
							assign node762 = (inp[11]) ? node782 : node763;
								assign node763 = (inp[9]) ? node773 : node764;
									assign node764 = (inp[10]) ? 14'b00000000000001 : node765;
										assign node765 = (inp[12]) ? node767 : 14'b00000000000001;
											assign node767 = (inp[2]) ? 14'b00010100100110 : node768;
												assign node768 = (inp[6]) ? 14'b01010100100110 : 14'b01010110100110;
									assign node773 = (inp[5]) ? 14'b00010100000000 : node774;
										assign node774 = (inp[6]) ? node778 : node775;
											assign node775 = (inp[12]) ? 14'b00111110000000 : 14'b01111110000000;
											assign node778 = (inp[10]) ? 14'b01111100000010 : 14'b00111100000110;
								assign node782 = (inp[10]) ? 14'b00000000000001 : node783;
									assign node783 = (inp[4]) ? node787 : node784;
										assign node784 = (inp[9]) ? 14'b00010100000100 : 14'b00111100100100;
										assign node787 = (inp[2]) ? 14'b00000000000001 : node788;
											assign node788 = (inp[12]) ? node790 : 14'b00000000000001;
												assign node790 = (inp[5]) ? 14'b01010110100000 : 14'b01011100000000;
						assign node796 = (inp[2]) ? node848 : node797;
							assign node797 = (inp[4]) ? node823 : node798;
								assign node798 = (inp[6]) ? node810 : node799;
									assign node799 = (inp[12]) ? 14'b00000000000001 : node800;
										assign node800 = (inp[5]) ? node804 : node801;
											assign node801 = (inp[7]) ? 14'b00000010110000 : 14'b00000000000001;
											assign node804 = (inp[11]) ? 14'b01100010010000 : node805;
												assign node805 = (inp[10]) ? 14'b01100110110000 : 14'b01100010110000;
									assign node810 = (inp[12]) ? node818 : node811;
										assign node811 = (inp[5]) ? 14'b01100100110000 : node812;
											assign node812 = (inp[7]) ? node814 : 14'b00000000000001;
												assign node814 = (inp[9]) ? 14'b00000000010000 : 14'b00000000110000;
										assign node818 = (inp[5]) ? 14'b00000000000001 : node819;
											assign node819 = (inp[7]) ? 14'b01000000110100 : 14'b01000100110100;
								assign node823 = (inp[5]) ? node839 : node824;
									assign node824 = (inp[12]) ? node832 : node825;
										assign node825 = (inp[9]) ? node827 : 14'b00100100110100;
											assign node827 = (inp[7]) ? node829 : 14'b00100110010100;
												assign node829 = (inp[6]) ? 14'b00100000010100 : 14'b00100010010100;
										assign node832 = (inp[7]) ? 14'b00000000110100 : node833;
											assign node833 = (inp[9]) ? node835 : 14'b00000110110100;
												assign node835 = (inp[6]) ? 14'b00000100010100 : 14'b00000110010100;
									assign node839 = (inp[12]) ? 14'b00000000000001 : node840;
										assign node840 = (inp[10]) ? 14'b00100110010000 : node841;
											assign node841 = (inp[9]) ? node843 : 14'b00100100110000;
												assign node843 = (inp[7]) ? 14'b00100000010000 : 14'b00100100010000;
							assign node848 = (inp[5]) ? node860 : node849;
								assign node849 = (inp[4]) ? 14'b00000000000001 : node850;
									assign node850 = (inp[12]) ? node856 : node851;
										assign node851 = (inp[9]) ? node853 : 14'b01100110110100;
											assign node853 = (inp[6]) ? 14'b01100000010100 : 14'b01100010010100;
										assign node856 = (inp[9]) ? 14'b01000010010000 : 14'b01000000110000;
								assign node860 = (inp[7]) ? 14'b00000000000001 : node861;
									assign node861 = (inp[12]) ? 14'b00000000000001 : node862;
										assign node862 = (inp[11]) ? node864 : 14'b00000000000001;
											assign node864 = (inp[10]) ? 14'b00000100110000 : 14'b00000110010000;
					assign node869 = (inp[9]) ? 14'b00000000000001 : node870;
						assign node870 = (inp[7]) ? node900 : node871;
							assign node871 = (inp[11]) ? node893 : node872;
								assign node872 = (inp[13]) ? node884 : node873;
									assign node873 = (inp[4]) ? node879 : node874;
										assign node874 = (inp[10]) ? node876 : 14'b01001110100110;
											assign node876 = (inp[12]) ? 14'b00000110100010 : 14'b01100110100010;
										assign node879 = (inp[10]) ? node881 : 14'b00000000000001;
											assign node881 = (inp[2]) ? 14'b00000000000001 : 14'b00101110100000;
									assign node884 = (inp[2]) ? node886 : 14'b00000000000001;
										assign node886 = (inp[6]) ? node888 : 14'b00000000000001;
											assign node888 = (inp[10]) ? 14'b01100100100100 : node889;
												assign node889 = (inp[12]) ? 14'b01000100100000 : 14'b00000100100000;
								assign node893 = (inp[10]) ? 14'b00000000000001 : node894;
									assign node894 = (inp[6]) ? node896 : 14'b00000000000001;
										assign node896 = (inp[5]) ? 14'b00100100100000 : 14'b01001110000000;
							assign node900 = (inp[6]) ? node902 : 14'b00000000000001;
								assign node902 = (inp[13]) ? node904 : 14'b00000000000001;
									assign node904 = (inp[2]) ? 14'b00000000000001 : node905;
										assign node905 = (inp[12]) ? 14'b01000000100100 : node906;
											assign node906 = (inp[5]) ? 14'b01100000100000 : 14'b00000000100000;
				assign node912 = (inp[7]) ? node982 : node913;
					assign node913 = (inp[13]) ? node971 : node914;
						assign node914 = (inp[6]) ? node952 : node915;
							assign node915 = (inp[9]) ? node941 : node916;
								assign node916 = (inp[10]) ? node934 : node917;
									assign node917 = (inp[4]) ? node927 : node918;
										assign node918 = (inp[2]) ? node924 : node919;
											assign node919 = (inp[5]) ? 14'b01010010100110 : node920;
												assign node920 = (inp[11]) ? 14'b01011010100100 : 14'b01011010100110;
											assign node924 = (inp[5]) ? 14'b00010010100000 : 14'b00011010100100;
										assign node927 = (inp[5]) ? node929 : 14'b00000000000001;
											assign node929 = (inp[12]) ? node931 : 14'b01100010100110;
												assign node931 = (inp[11]) ? 14'b01000010100000 : 14'b01000010100010;
									assign node934 = (inp[11]) ? 14'b00000000000001 : node935;
										assign node935 = (inp[3]) ? node937 : 14'b00111010100000;
											assign node937 = (inp[12]) ? 14'b00000000000001 : 14'b00100010100000;
								assign node941 = (inp[3]) ? node943 : 14'b00000000000001;
									assign node943 = (inp[2]) ? 14'b00000000000001 : node944;
										assign node944 = (inp[12]) ? node946 : 14'b01101010000110;
											assign node946 = (inp[10]) ? 14'b01001010000010 : node947;
												assign node947 = (inp[11]) ? 14'b01001010000000 : 14'b00000000000001;
							assign node952 = (inp[3]) ? 14'b00000000000001 : node953;
								assign node953 = (inp[4]) ? node965 : node954;
									assign node954 = (inp[9]) ? node956 : 14'b00000000000001;
										assign node956 = (inp[5]) ? node962 : node957;
											assign node957 = (inp[12]) ? 14'b00011000000100 : node958;
												assign node958 = (inp[11]) ? 14'b01111000000100 : 14'b01111000000010;
											assign node962 = (inp[11]) ? 14'b00000000000001 : 14'b00010000000000;
									assign node965 = (inp[12]) ? node967 : 14'b00000000000001;
										assign node967 = (inp[9]) ? 14'b00000000000001 : 14'b10000000000000;
						assign node971 = (inp[2]) ? 14'b00000000000001 : node972;
							assign node972 = (inp[12]) ? 14'b00000000000001 : node973;
								assign node973 = (inp[3]) ? node975 : 14'b00000000000001;
									assign node975 = (inp[6]) ? 14'b00000000000001 : node976;
										assign node976 = (inp[4]) ? 14'b00000000000001 : 14'b10000000000010;
					assign node982 = (inp[13]) ? node984 : 14'b00000000000001;
						assign node984 = (inp[3]) ? node986 : 14'b00000000000001;
							assign node986 = (inp[6]) ? 14'b00000000000001 : node987;
								assign node987 = (inp[2]) ? node989 : 14'b00000000000001;
									assign node989 = (inp[11]) ? 14'b10001000001010 : 14'b00000000000001;

endmodule