module dtc_split5_bm59 (
	input  wire [12-1:0] inp,
	output wire [3-1:0] outp
);

	wire [3-1:0] node1;
	wire [3-1:0] node2;
	wire [3-1:0] node3;
	wire [3-1:0] node4;
	wire [3-1:0] node5;
	wire [3-1:0] node6;
	wire [3-1:0] node7;
	wire [3-1:0] node8;
	wire [3-1:0] node10;
	wire [3-1:0] node12;
	wire [3-1:0] node16;
	wire [3-1:0] node17;
	wire [3-1:0] node19;
	wire [3-1:0] node20;
	wire [3-1:0] node24;
	wire [3-1:0] node25;
	wire [3-1:0] node26;
	wire [3-1:0] node29;
	wire [3-1:0] node31;
	wire [3-1:0] node34;
	wire [3-1:0] node38;
	wire [3-1:0] node39;
	wire [3-1:0] node40;
	wire [3-1:0] node41;
	wire [3-1:0] node43;
	wire [3-1:0] node45;
	wire [3-1:0] node48;
	wire [3-1:0] node49;
	wire [3-1:0] node53;
	wire [3-1:0] node54;
	wire [3-1:0] node55;
	wire [3-1:0] node57;
	wire [3-1:0] node60;
	wire [3-1:0] node63;
	wire [3-1:0] node65;
	wire [3-1:0] node68;
	wire [3-1:0] node69;
	wire [3-1:0] node70;
	wire [3-1:0] node72;
	wire [3-1:0] node75;
	wire [3-1:0] node77;
	wire [3-1:0] node78;
	wire [3-1:0] node82;
	wire [3-1:0] node83;
	wire [3-1:0] node84;
	wire [3-1:0] node88;
	wire [3-1:0] node90;
	wire [3-1:0] node92;
	wire [3-1:0] node96;
	wire [3-1:0] node97;
	wire [3-1:0] node98;
	wire [3-1:0] node99;
	wire [3-1:0] node100;
	wire [3-1:0] node102;
	wire [3-1:0] node104;
	wire [3-1:0] node107;
	wire [3-1:0] node108;
	wire [3-1:0] node109;
	wire [3-1:0] node110;
	wire [3-1:0] node113;
	wire [3-1:0] node114;
	wire [3-1:0] node118;
	wire [3-1:0] node119;
	wire [3-1:0] node122;
	wire [3-1:0] node125;
	wire [3-1:0] node126;
	wire [3-1:0] node127;
	wire [3-1:0] node131;
	wire [3-1:0] node134;
	wire [3-1:0] node135;
	wire [3-1:0] node136;
	wire [3-1:0] node138;
	wire [3-1:0] node140;
	wire [3-1:0] node142;
	wire [3-1:0] node145;
	wire [3-1:0] node146;
	wire [3-1:0] node148;
	wire [3-1:0] node151;
	wire [3-1:0] node152;
	wire [3-1:0] node153;
	wire [3-1:0] node158;
	wire [3-1:0] node159;
	wire [3-1:0] node161;
	wire [3-1:0] node163;
	wire [3-1:0] node167;
	wire [3-1:0] node168;
	wire [3-1:0] node169;
	wire [3-1:0] node170;
	wire [3-1:0] node173;
	wire [3-1:0] node174;
	wire [3-1:0] node177;
	wire [3-1:0] node178;
	wire [3-1:0] node182;
	wire [3-1:0] node183;
	wire [3-1:0] node184;
	wire [3-1:0] node185;
	wire [3-1:0] node189;
	wire [3-1:0] node190;
	wire [3-1:0] node192;
	wire [3-1:0] node196;
	wire [3-1:0] node197;
	wire [3-1:0] node199;
	wire [3-1:0] node202;
	wire [3-1:0] node204;
	wire [3-1:0] node208;
	wire [3-1:0] node209;
	wire [3-1:0] node210;
	wire [3-1:0] node211;
	wire [3-1:0] node212;
	wire [3-1:0] node213;
	wire [3-1:0] node215;
	wire [3-1:0] node218;
	wire [3-1:0] node219;
	wire [3-1:0] node223;
	wire [3-1:0] node225;
	wire [3-1:0] node226;
	wire [3-1:0] node227;
	wire [3-1:0] node231;
	wire [3-1:0] node233;
	wire [3-1:0] node236;
	wire [3-1:0] node237;
	wire [3-1:0] node238;
	wire [3-1:0] node239;
	wire [3-1:0] node240;
	wire [3-1:0] node244;
	wire [3-1:0] node247;
	wire [3-1:0] node249;
	wire [3-1:0] node252;
	wire [3-1:0] node253;
	wire [3-1:0] node254;
	wire [3-1:0] node256;
	wire [3-1:0] node260;
	wire [3-1:0] node261;
	wire [3-1:0] node264;
	wire [3-1:0] node267;
	wire [3-1:0] node268;
	wire [3-1:0] node269;
	wire [3-1:0] node270;
	wire [3-1:0] node272;
	wire [3-1:0] node276;
	wire [3-1:0] node277;
	wire [3-1:0] node280;
	wire [3-1:0] node281;
	wire [3-1:0] node282;
	wire [3-1:0] node286;
	wire [3-1:0] node287;
	wire [3-1:0] node291;
	wire [3-1:0] node292;
	wire [3-1:0] node293;
	wire [3-1:0] node295;
	wire [3-1:0] node298;
	wire [3-1:0] node300;
	wire [3-1:0] node304;
	wire [3-1:0] node305;
	wire [3-1:0] node306;
	wire [3-1:0] node307;
	wire [3-1:0] node308;
	wire [3-1:0] node311;
	wire [3-1:0] node314;
	wire [3-1:0] node315;
	wire [3-1:0] node319;
	wire [3-1:0] node320;
	wire [3-1:0] node322;
	wire [3-1:0] node324;
	wire [3-1:0] node328;
	wire [3-1:0] node329;
	wire [3-1:0] node330;
	wire [3-1:0] node331;
	wire [3-1:0] node334;
	wire [3-1:0] node335;
	wire [3-1:0] node336;
	wire [3-1:0] node339;
	wire [3-1:0] node345;
	wire [3-1:0] node346;
	wire [3-1:0] node347;
	wire [3-1:0] node348;
	wire [3-1:0] node350;
	wire [3-1:0] node351;
	wire [3-1:0] node352;
	wire [3-1:0] node354;
	wire [3-1:0] node356;
	wire [3-1:0] node359;
	wire [3-1:0] node361;
	wire [3-1:0] node365;
	wire [3-1:0] node366;
	wire [3-1:0] node367;
	wire [3-1:0] node368;
	wire [3-1:0] node369;
	wire [3-1:0] node370;
	wire [3-1:0] node372;
	wire [3-1:0] node376;
	wire [3-1:0] node379;
	wire [3-1:0] node380;
	wire [3-1:0] node381;
	wire [3-1:0] node385;
	wire [3-1:0] node386;
	wire [3-1:0] node390;
	wire [3-1:0] node391;
	wire [3-1:0] node392;
	wire [3-1:0] node395;
	wire [3-1:0] node396;
	wire [3-1:0] node398;
	wire [3-1:0] node401;
	wire [3-1:0] node402;
	wire [3-1:0] node406;
	wire [3-1:0] node407;
	wire [3-1:0] node409;
	wire [3-1:0] node412;
	wire [3-1:0] node415;
	wire [3-1:0] node417;
	wire [3-1:0] node418;
	wire [3-1:0] node419;
	wire [3-1:0] node421;
	wire [3-1:0] node424;
	wire [3-1:0] node426;
	wire [3-1:0] node429;
	wire [3-1:0] node431;
	wire [3-1:0] node435;
	wire [3-1:0] node436;
	wire [3-1:0] node437;
	wire [3-1:0] node438;
	wire [3-1:0] node439;
	wire [3-1:0] node440;
	wire [3-1:0] node441;
	wire [3-1:0] node442;
	wire [3-1:0] node447;
	wire [3-1:0] node448;
	wire [3-1:0] node450;
	wire [3-1:0] node453;
	wire [3-1:0] node454;
	wire [3-1:0] node456;
	wire [3-1:0] node460;
	wire [3-1:0] node461;
	wire [3-1:0] node462;
	wire [3-1:0] node464;
	wire [3-1:0] node466;
	wire [3-1:0] node469;
	wire [3-1:0] node470;
	wire [3-1:0] node472;
	wire [3-1:0] node475;
	wire [3-1:0] node478;
	wire [3-1:0] node479;
	wire [3-1:0] node480;
	wire [3-1:0] node485;
	wire [3-1:0] node486;
	wire [3-1:0] node487;
	wire [3-1:0] node488;
	wire [3-1:0] node490;
	wire [3-1:0] node491;
	wire [3-1:0] node496;
	wire [3-1:0] node497;
	wire [3-1:0] node498;
	wire [3-1:0] node501;
	wire [3-1:0] node503;
	wire [3-1:0] node507;
	wire [3-1:0] node508;
	wire [3-1:0] node509;
	wire [3-1:0] node513;
	wire [3-1:0] node515;
	wire [3-1:0] node518;
	wire [3-1:0] node519;
	wire [3-1:0] node520;
	wire [3-1:0] node521;
	wire [3-1:0] node522;
	wire [3-1:0] node524;
	wire [3-1:0] node526;
	wire [3-1:0] node530;
	wire [3-1:0] node531;
	wire [3-1:0] node532;
	wire [3-1:0] node536;
	wire [3-1:0] node539;
	wire [3-1:0] node540;
	wire [3-1:0] node541;
	wire [3-1:0] node543;
	wire [3-1:0] node547;
	wire [3-1:0] node549;
	wire [3-1:0] node552;
	wire [3-1:0] node553;
	wire [3-1:0] node555;
	wire [3-1:0] node556;
	wire [3-1:0] node560;
	wire [3-1:0] node561;
	wire [3-1:0] node563;
	wire [3-1:0] node564;
	wire [3-1:0] node566;
	wire [3-1:0] node571;
	wire [3-1:0] node572;
	wire [3-1:0] node573;
	wire [3-1:0] node575;
	wire [3-1:0] node576;
	wire [3-1:0] node578;
	wire [3-1:0] node579;
	wire [3-1:0] node582;
	wire [3-1:0] node585;
	wire [3-1:0] node587;
	wire [3-1:0] node591;
	wire [3-1:0] node592;
	wire [3-1:0] node593;
	wire [3-1:0] node594;
	wire [3-1:0] node595;
	wire [3-1:0] node599;
	wire [3-1:0] node602;
	wire [3-1:0] node603;
	wire [3-1:0] node604;
	wire [3-1:0] node608;
	wire [3-1:0] node609;
	wire [3-1:0] node610;
	wire [3-1:0] node613;
	wire [3-1:0] node617;
	wire [3-1:0] node618;
	wire [3-1:0] node619;
	wire [3-1:0] node620;
	wire [3-1:0] node622;
	wire [3-1:0] node627;
	wire [3-1:0] node629;
	wire [3-1:0] node631;
	wire [3-1:0] node633;
	wire [3-1:0] node636;
	wire [3-1:0] node637;
	wire [3-1:0] node638;
	wire [3-1:0] node639;
	wire [3-1:0] node640;
	wire [3-1:0] node641;
	wire [3-1:0] node642;
	wire [3-1:0] node643;
	wire [3-1:0] node644;
	wire [3-1:0] node647;
	wire [3-1:0] node650;
	wire [3-1:0] node652;
	wire [3-1:0] node655;
	wire [3-1:0] node656;
	wire [3-1:0] node658;
	wire [3-1:0] node661;
	wire [3-1:0] node662;
	wire [3-1:0] node664;
	wire [3-1:0] node669;
	wire [3-1:0] node670;
	wire [3-1:0] node671;
	wire [3-1:0] node672;
	wire [3-1:0] node673;
	wire [3-1:0] node676;
	wire [3-1:0] node679;
	wire [3-1:0] node680;
	wire [3-1:0] node681;
	wire [3-1:0] node686;
	wire [3-1:0] node687;
	wire [3-1:0] node689;
	wire [3-1:0] node691;
	wire [3-1:0] node694;
	wire [3-1:0] node696;
	wire [3-1:0] node699;
	wire [3-1:0] node700;
	wire [3-1:0] node701;
	wire [3-1:0] node702;
	wire [3-1:0] node704;
	wire [3-1:0] node707;
	wire [3-1:0] node708;
	wire [3-1:0] node709;
	wire [3-1:0] node712;
	wire [3-1:0] node716;
	wire [3-1:0] node718;
	wire [3-1:0] node721;
	wire [3-1:0] node722;
	wire [3-1:0] node723;
	wire [3-1:0] node726;
	wire [3-1:0] node728;
	wire [3-1:0] node731;
	wire [3-1:0] node732;
	wire [3-1:0] node733;
	wire [3-1:0] node737;
	wire [3-1:0] node738;
	wire [3-1:0] node743;
	wire [3-1:0] node744;
	wire [3-1:0] node745;
	wire [3-1:0] node746;
	wire [3-1:0] node747;
	wire [3-1:0] node748;
	wire [3-1:0] node749;
	wire [3-1:0] node752;
	wire [3-1:0] node755;
	wire [3-1:0] node756;
	wire [3-1:0] node759;
	wire [3-1:0] node760;
	wire [3-1:0] node761;
	wire [3-1:0] node766;
	wire [3-1:0] node767;
	wire [3-1:0] node768;
	wire [3-1:0] node769;
	wire [3-1:0] node772;
	wire [3-1:0] node776;
	wire [3-1:0] node777;
	wire [3-1:0] node778;
	wire [3-1:0] node782;
	wire [3-1:0] node784;
	wire [3-1:0] node787;
	wire [3-1:0] node788;
	wire [3-1:0] node789;
	wire [3-1:0] node790;
	wire [3-1:0] node791;
	wire [3-1:0] node794;
	wire [3-1:0] node798;
	wire [3-1:0] node799;
	wire [3-1:0] node801;
	wire [3-1:0] node804;
	wire [3-1:0] node807;
	wire [3-1:0] node808;
	wire [3-1:0] node810;
	wire [3-1:0] node812;
	wire [3-1:0] node815;
	wire [3-1:0] node816;
	wire [3-1:0] node820;
	wire [3-1:0] node821;
	wire [3-1:0] node822;
	wire [3-1:0] node823;
	wire [3-1:0] node824;
	wire [3-1:0] node826;
	wire [3-1:0] node828;
	wire [3-1:0] node831;
	wire [3-1:0] node834;
	wire [3-1:0] node835;
	wire [3-1:0] node839;
	wire [3-1:0] node840;
	wire [3-1:0] node842;
	wire [3-1:0] node844;
	wire [3-1:0] node846;
	wire [3-1:0] node849;
	wire [3-1:0] node851;
	wire [3-1:0] node853;
	wire [3-1:0] node857;
	wire [3-1:0] node858;
	wire [3-1:0] node859;
	wire [3-1:0] node860;
	wire [3-1:0] node861;
	wire [3-1:0] node863;
	wire [3-1:0] node864;
	wire [3-1:0] node867;
	wire [3-1:0] node870;
	wire [3-1:0] node871;
	wire [3-1:0] node872;
	wire [3-1:0] node874;
	wire [3-1:0] node878;
	wire [3-1:0] node879;
	wire [3-1:0] node883;
	wire [3-1:0] node884;
	wire [3-1:0] node885;
	wire [3-1:0] node886;
	wire [3-1:0] node890;
	wire [3-1:0] node891;
	wire [3-1:0] node893;
	wire [3-1:0] node897;
	wire [3-1:0] node898;
	wire [3-1:0] node899;
	wire [3-1:0] node904;
	wire [3-1:0] node905;
	wire [3-1:0] node907;
	wire [3-1:0] node908;
	wire [3-1:0] node912;
	wire [3-1:0] node913;
	wire [3-1:0] node914;
	wire [3-1:0] node915;
	wire [3-1:0] node920;
	wire [3-1:0] node921;
	wire [3-1:0] node923;
	wire [3-1:0] node925;
	wire [3-1:0] node928;
	wire [3-1:0] node930;
	wire [3-1:0] node933;
	wire [3-1:0] node934;
	wire [3-1:0] node935;
	wire [3-1:0] node936;
	wire [3-1:0] node937;
	wire [3-1:0] node939;
	wire [3-1:0] node941;
	wire [3-1:0] node944;
	wire [3-1:0] node945;
	wire [3-1:0] node949;
	wire [3-1:0] node950;
	wire [3-1:0] node951;
	wire [3-1:0] node955;
	wire [3-1:0] node957;
	wire [3-1:0] node958;
	wire [3-1:0] node961;
	wire [3-1:0] node964;
	wire [3-1:0] node965;
	wire [3-1:0] node966;
	wire [3-1:0] node967;
	wire [3-1:0] node970;
	wire [3-1:0] node972;
	wire [3-1:0] node977;
	wire [3-1:0] node978;
	wire [3-1:0] node979;
	wire [3-1:0] node980;
	wire [3-1:0] node982;
	wire [3-1:0] node985;
	wire [3-1:0] node986;
	wire [3-1:0] node989;
	wire [3-1:0] node994;
	wire [3-1:0] node995;
	wire [3-1:0] node996;
	wire [3-1:0] node997;
	wire [3-1:0] node999;
	wire [3-1:0] node1000;
	wire [3-1:0] node1001;
	wire [3-1:0] node1003;
	wire [3-1:0] node1008;
	wire [3-1:0] node1009;
	wire [3-1:0] node1010;
	wire [3-1:0] node1011;
	wire [3-1:0] node1012;
	wire [3-1:0] node1015;
	wire [3-1:0] node1018;
	wire [3-1:0] node1019;
	wire [3-1:0] node1022;
	wire [3-1:0] node1024;
	wire [3-1:0] node1027;
	wire [3-1:0] node1028;
	wire [3-1:0] node1030;
	wire [3-1:0] node1031;
	wire [3-1:0] node1034;
	wire [3-1:0] node1037;
	wire [3-1:0] node1039;
	wire [3-1:0] node1040;
	wire [3-1:0] node1043;
	wire [3-1:0] node1046;
	wire [3-1:0] node1048;
	wire [3-1:0] node1049;
	wire [3-1:0] node1051;
	wire [3-1:0] node1053;
	wire [3-1:0] node1056;
	wire [3-1:0] node1058;
	wire [3-1:0] node1061;
	wire [3-1:0] node1062;
	wire [3-1:0] node1063;
	wire [3-1:0] node1064;
	wire [3-1:0] node1065;
	wire [3-1:0] node1066;
	wire [3-1:0] node1070;
	wire [3-1:0] node1071;
	wire [3-1:0] node1072;
	wire [3-1:0] node1075;
	wire [3-1:0] node1078;
	wire [3-1:0] node1080;
	wire [3-1:0] node1083;
	wire [3-1:0] node1084;
	wire [3-1:0] node1085;
	wire [3-1:0] node1086;
	wire [3-1:0] node1090;
	wire [3-1:0] node1092;
	wire [3-1:0] node1093;
	wire [3-1:0] node1096;
	wire [3-1:0] node1099;
	wire [3-1:0] node1100;
	wire [3-1:0] node1102;
	wire [3-1:0] node1105;
	wire [3-1:0] node1106;
	wire [3-1:0] node1110;
	wire [3-1:0] node1111;
	wire [3-1:0] node1112;
	wire [3-1:0] node1113;
	wire [3-1:0] node1116;
	wire [3-1:0] node1117;
	wire [3-1:0] node1121;
	wire [3-1:0] node1122;
	wire [3-1:0] node1124;
	wire [3-1:0] node1127;
	wire [3-1:0] node1129;
	wire [3-1:0] node1132;
	wire [3-1:0] node1133;
	wire [3-1:0] node1134;
	wire [3-1:0] node1138;
	wire [3-1:0] node1139;
	wire [3-1:0] node1141;
	wire [3-1:0] node1144;
	wire [3-1:0] node1146;
	wire [3-1:0] node1149;
	wire [3-1:0] node1150;
	wire [3-1:0] node1151;
	wire [3-1:0] node1152;
	wire [3-1:0] node1153;
	wire [3-1:0] node1154;
	wire [3-1:0] node1158;
	wire [3-1:0] node1159;
	wire [3-1:0] node1163;
	wire [3-1:0] node1164;
	wire [3-1:0] node1167;
	wire [3-1:0] node1168;
	wire [3-1:0] node1172;
	wire [3-1:0] node1174;
	wire [3-1:0] node1175;
	wire [3-1:0] node1176;
	wire [3-1:0] node1177;
	wire [3-1:0] node1181;
	wire [3-1:0] node1184;
	wire [3-1:0] node1185;
	wire [3-1:0] node1189;
	wire [3-1:0] node1190;
	wire [3-1:0] node1191;
	wire [3-1:0] node1192;
	wire [3-1:0] node1196;
	wire [3-1:0] node1197;
	wire [3-1:0] node1199;
	wire [3-1:0] node1202;
	wire [3-1:0] node1203;
	wire [3-1:0] node1207;
	wire [3-1:0] node1208;
	wire [3-1:0] node1209;
	wire [3-1:0] node1210;
	wire [3-1:0] node1213;
	wire [3-1:0] node1218;
	wire [3-1:0] node1220;
	wire [3-1:0] node1221;
	wire [3-1:0] node1222;
	wire [3-1:0] node1224;
	wire [3-1:0] node1225;
	wire [3-1:0] node1229;
	wire [3-1:0] node1230;
	wire [3-1:0] node1231;
	wire [3-1:0] node1232;
	wire [3-1:0] node1233;
	wire [3-1:0] node1237;
	wire [3-1:0] node1238;
	wire [3-1:0] node1242;
	wire [3-1:0] node1245;
	wire [3-1:0] node1246;
	wire [3-1:0] node1247;
	wire [3-1:0] node1252;
	wire [3-1:0] node1253;
	wire [3-1:0] node1254;
	wire [3-1:0] node1255;

	assign outp = (inp[10]) ? node636 : node1;
		assign node1 = (inp[9]) ? node345 : node2;
			assign node2 = (inp[2]) ? node96 : node3;
				assign node3 = (inp[0]) ? 3'b110 : node4;
					assign node4 = (inp[1]) ? node38 : node5;
						assign node5 = (inp[3]) ? 3'b111 : node6;
							assign node6 = (inp[7]) ? node16 : node7;
								assign node7 = (inp[8]) ? 3'b111 : node8;
									assign node8 = (inp[5]) ? node10 : 3'b000;
										assign node10 = (inp[6]) ? node12 : 3'b010;
											assign node12 = (inp[11]) ? 3'b010 : 3'b000;
								assign node16 = (inp[8]) ? node24 : node17;
									assign node17 = (inp[5]) ? node19 : 3'b100;
										assign node19 = (inp[11]) ? 3'b110 : node20;
											assign node20 = (inp[6]) ? 3'b100 : 3'b110;
									assign node24 = (inp[4]) ? node34 : node25;
										assign node25 = (inp[5]) ? node29 : node26;
											assign node26 = (inp[11]) ? 3'b000 : 3'b010;
											assign node29 = (inp[6]) ? node31 : 3'b010;
												assign node31 = (inp[11]) ? 3'b010 : 3'b000;
										assign node34 = (inp[6]) ? 3'b100 : 3'b110;
						assign node38 = (inp[5]) ? node68 : node39;
							assign node39 = (inp[6]) ? node53 : node40;
								assign node40 = (inp[7]) ? node48 : node41;
									assign node41 = (inp[11]) ? node43 : 3'b000;
										assign node43 = (inp[3]) ? node45 : 3'b000;
											assign node45 = (inp[8]) ? 3'b111 : 3'b000;
									assign node48 = (inp[4]) ? 3'b100 : node49;
										assign node49 = (inp[8]) ? 3'b000 : 3'b100;
								assign node53 = (inp[11]) ? node63 : node54;
									assign node54 = (inp[7]) ? node60 : node55;
										assign node55 = (inp[3]) ? node57 : 3'b110;
											assign node57 = (inp[4]) ? 3'b010 : 3'b111;
										assign node60 = (inp[8]) ? 3'b010 : 3'b110;
									assign node63 = (inp[7]) ? node65 : 3'b000;
										assign node65 = (inp[4]) ? 3'b100 : 3'b000;
							assign node68 = (inp[7]) ? node82 : node69;
								assign node69 = (inp[8]) ? node75 : node70;
									assign node70 = (inp[6]) ? node72 : 3'b010;
										assign node72 = (inp[11]) ? 3'b010 : 3'b000;
									assign node75 = (inp[4]) ? node77 : 3'b111;
										assign node77 = (inp[11]) ? 3'b010 : node78;
											assign node78 = (inp[6]) ? 3'b000 : 3'b010;
								assign node82 = (inp[6]) ? node88 : node83;
									assign node83 = (inp[4]) ? 3'b110 : node84;
										assign node84 = (inp[8]) ? 3'b010 : 3'b110;
									assign node88 = (inp[11]) ? node90 : 3'b100;
										assign node90 = (inp[8]) ? node92 : 3'b110;
											assign node92 = (inp[4]) ? 3'b110 : 3'b010;
				assign node96 = (inp[1]) ? node208 : node97;
					assign node97 = (inp[0]) ? node167 : node98;
						assign node98 = (inp[11]) ? node134 : node99;
							assign node99 = (inp[4]) ? node107 : node100;
								assign node100 = (inp[8]) ? node102 : 3'b000;
									assign node102 = (inp[7]) ? node104 : 3'b110;
										assign node104 = (inp[5]) ? 3'b000 : 3'b100;
								assign node107 = (inp[6]) ? node125 : node108;
									assign node108 = (inp[8]) ? node118 : node109;
										assign node109 = (inp[3]) ? node113 : node110;
											assign node110 = (inp[7]) ? 3'b010 : 3'b100;
											assign node113 = (inp[5]) ? 3'b010 : node114;
												assign node114 = (inp[7]) ? 3'b100 : 3'b000;
										assign node118 = (inp[5]) ? node122 : node119;
											assign node119 = (inp[7]) ? 3'b010 : 3'b000;
											assign node122 = (inp[7]) ? 3'b100 : 3'b010;
									assign node125 = (inp[3]) ? node131 : node126;
										assign node126 = (inp[5]) ? 3'b100 : node127;
											assign node127 = (inp[8]) ? 3'b000 : 3'b100;
										assign node131 = (inp[5]) ? 3'b100 : 3'b110;
							assign node134 = (inp[5]) ? node158 : node135;
								assign node135 = (inp[8]) ? node145 : node136;
									assign node136 = (inp[4]) ? node138 : 3'b010;
										assign node138 = (inp[6]) ? node140 : 3'b100;
											assign node140 = (inp[3]) ? node142 : 3'b110;
												assign node142 = (inp[7]) ? 3'b110 : 3'b000;
									assign node145 = (inp[4]) ? node151 : node146;
										assign node146 = (inp[7]) ? node148 : 3'b100;
											assign node148 = (inp[3]) ? 3'b000 : 3'b110;
										assign node151 = (inp[6]) ? 3'b010 : node152;
											assign node152 = (inp[3]) ? 3'b000 : node153;
												assign node153 = (inp[7]) ? 3'b000 : 3'b010;
								assign node158 = (inp[4]) ? 3'b110 : node159;
									assign node159 = (inp[3]) ? node161 : 3'b010;
										assign node161 = (inp[8]) ? node163 : 3'b010;
											assign node163 = (inp[7]) ? 3'b010 : 3'b110;
						assign node167 = (inp[3]) ? 3'b110 : node168;
							assign node168 = (inp[5]) ? node182 : node169;
								assign node169 = (inp[11]) ? node173 : node170;
									assign node170 = (inp[6]) ? 3'b010 : 3'b000;
									assign node173 = (inp[7]) ? node177 : node174;
										assign node174 = (inp[4]) ? 3'b000 : 3'b110;
										assign node177 = (inp[4]) ? 3'b100 : node178;
											assign node178 = (inp[8]) ? 3'b000 : 3'b100;
								assign node182 = (inp[11]) ? node196 : node183;
									assign node183 = (inp[6]) ? node189 : node184;
										assign node184 = (inp[4]) ? 3'b110 : node185;
											assign node185 = (inp[8]) ? 3'b110 : 3'b010;
										assign node189 = (inp[4]) ? 3'b000 : node190;
											assign node190 = (inp[7]) ? node192 : 3'b110;
												assign node192 = (inp[8]) ? 3'b000 : 3'b100;
									assign node196 = (inp[7]) ? node202 : node197;
										assign node197 = (inp[8]) ? node199 : 3'b010;
											assign node199 = (inp[4]) ? 3'b010 : 3'b110;
										assign node202 = (inp[8]) ? node204 : 3'b110;
											assign node204 = (inp[4]) ? 3'b110 : 3'b010;
					assign node208 = (inp[7]) ? node304 : node209;
						assign node209 = (inp[11]) ? node267 : node210;
							assign node210 = (inp[3]) ? node236 : node211;
								assign node211 = (inp[0]) ? node223 : node212;
									assign node212 = (inp[5]) ? node218 : node213;
										assign node213 = (inp[6]) ? node215 : 3'b100;
											assign node215 = (inp[4]) ? 3'b010 : 3'b100;
										assign node218 = (inp[4]) ? 3'b000 : node219;
											assign node219 = (inp[8]) ? 3'b010 : 3'b110;
									assign node223 = (inp[6]) ? node225 : 3'b000;
										assign node225 = (inp[4]) ? node231 : node226;
											assign node226 = (inp[5]) ? 3'b000 : node227;
												assign node227 = (inp[8]) ? 3'b110 : 3'b000;
											assign node231 = (inp[8]) ? node233 : 3'b100;
												assign node233 = (inp[5]) ? 3'b100 : 3'b000;
								assign node236 = (inp[8]) ? node252 : node237;
									assign node237 = (inp[4]) ? node247 : node238;
										assign node238 = (inp[5]) ? node244 : node239;
											assign node239 = (inp[6]) ? 3'b000 : node240;
												assign node240 = (inp[0]) ? 3'b000 : 3'b010;
											assign node244 = (inp[0]) ? 3'b010 : 3'b100;
										assign node247 = (inp[6]) ? node249 : 3'b010;
											assign node249 = (inp[5]) ? 3'b000 : 3'b010;
									assign node252 = (inp[5]) ? node260 : node253;
										assign node253 = (inp[0]) ? 3'b110 : node254;
											assign node254 = (inp[4]) ? node256 : 3'b100;
												assign node256 = (inp[6]) ? 3'b100 : 3'b110;
										assign node260 = (inp[4]) ? node264 : node261;
											assign node261 = (inp[0]) ? 3'b110 : 3'b010;
											assign node264 = (inp[0]) ? 3'b000 : 3'b010;
							assign node267 = (inp[5]) ? node291 : node268;
								assign node268 = (inp[8]) ? node276 : node269;
									assign node269 = (inp[3]) ? 3'b000 : node270;
										assign node270 = (inp[4]) ? node272 : 3'b010;
											assign node272 = (inp[0]) ? 3'b000 : 3'b010;
									assign node276 = (inp[6]) ? node280 : node277;
										assign node277 = (inp[4]) ? 3'b010 : 3'b110;
										assign node280 = (inp[3]) ? node286 : node281;
											assign node281 = (inp[4]) ? 3'b100 : node282;
												assign node282 = (inp[0]) ? 3'b100 : 3'b010;
											assign node286 = (inp[0]) ? 3'b000 : node287;
												assign node287 = (inp[4]) ? 3'b010 : 3'b000;
								assign node291 = (inp[4]) ? 3'b010 : node292;
									assign node292 = (inp[6]) ? node298 : node293;
										assign node293 = (inp[3]) ? node295 : 3'b010;
											assign node295 = (inp[8]) ? 3'b010 : 3'b110;
										assign node298 = (inp[0]) ? node300 : 3'b110;
											assign node300 = (inp[3]) ? 3'b110 : 3'b010;
						assign node304 = (inp[4]) ? node328 : node305;
							assign node305 = (inp[11]) ? node319 : node306;
								assign node306 = (inp[0]) ? node314 : node307;
									assign node307 = (inp[5]) ? node311 : node308;
										assign node308 = (inp[3]) ? 3'b000 : 3'b010;
										assign node311 = (inp[3]) ? 3'b010 : 3'b000;
									assign node314 = (inp[5]) ? 3'b000 : node315;
										assign node315 = (inp[6]) ? 3'b010 : 3'b000;
								assign node319 = (inp[5]) ? 3'b010 : node320;
									assign node320 = (inp[0]) ? node322 : 3'b010;
										assign node322 = (inp[8]) ? node324 : 3'b000;
											assign node324 = (inp[6]) ? 3'b000 : 3'b010;
							assign node328 = (inp[11]) ? 3'b000 : node329;
								assign node329 = (inp[5]) ? 3'b000 : node330;
									assign node330 = (inp[6]) ? node334 : node331;
										assign node331 = (inp[3]) ? 3'b010 : 3'b000;
										assign node334 = (inp[3]) ? 3'b000 : node335;
											assign node335 = (inp[0]) ? node339 : node336;
												assign node336 = (inp[8]) ? 3'b000 : 3'b010;
												assign node339 = (inp[8]) ? 3'b010 : 3'b000;
			assign node345 = (inp[2]) ? node435 : node346;
				assign node346 = (inp[0]) ? 3'b010 : node347;
					assign node347 = (inp[1]) ? node365 : node348;
						assign node348 = (inp[7]) ? node350 : 3'b011;
							assign node350 = (inp[3]) ? 3'b011 : node351;
								assign node351 = (inp[8]) ? node359 : node352;
									assign node352 = (inp[5]) ? node354 : 3'b000;
										assign node354 = (inp[6]) ? node356 : 3'b010;
											assign node356 = (inp[4]) ? 3'b010 : 3'b000;
									assign node359 = (inp[4]) ? node361 : 3'b011;
										assign node361 = (inp[5]) ? 3'b010 : 3'b000;
						assign node365 = (inp[3]) ? node415 : node366;
							assign node366 = (inp[5]) ? node390 : node367;
								assign node367 = (inp[11]) ? node379 : node368;
									assign node368 = (inp[6]) ? node376 : node369;
										assign node369 = (inp[4]) ? 3'b000 : node370;
											assign node370 = (inp[8]) ? node372 : 3'b100;
												assign node372 = (inp[7]) ? 3'b100 : 3'b000;
										assign node376 = (inp[7]) ? 3'b110 : 3'b010;
									assign node379 = (inp[7]) ? node385 : node380;
										assign node380 = (inp[4]) ? 3'b100 : node381;
											assign node381 = (inp[8]) ? 3'b000 : 3'b100;
										assign node385 = (inp[6]) ? 3'b000 : node386;
											assign node386 = (inp[8]) ? 3'b100 : 3'b000;
								assign node390 = (inp[6]) ? node406 : node391;
									assign node391 = (inp[8]) ? node395 : node392;
										assign node392 = (inp[7]) ? 3'b010 : 3'b110;
										assign node395 = (inp[11]) ? node401 : node396;
											assign node396 = (inp[7]) ? node398 : 3'b010;
												assign node398 = (inp[4]) ? 3'b010 : 3'b110;
											assign node401 = (inp[7]) ? 3'b110 : node402;
												assign node402 = (inp[4]) ? 3'b110 : 3'b010;
									assign node406 = (inp[11]) ? node412 : node407;
										assign node407 = (inp[4]) ? node409 : 3'b100;
											assign node409 = (inp[7]) ? 3'b000 : 3'b100;
										assign node412 = (inp[7]) ? 3'b010 : 3'b110;
							assign node415 = (inp[7]) ? node417 : 3'b011;
								assign node417 = (inp[8]) ? node429 : node418;
									assign node418 = (inp[5]) ? node424 : node419;
										assign node419 = (inp[6]) ? node421 : 3'b000;
											assign node421 = (inp[11]) ? 3'b000 : 3'b010;
										assign node424 = (inp[6]) ? node426 : 3'b010;
											assign node426 = (inp[11]) ? 3'b010 : 3'b000;
									assign node429 = (inp[4]) ? node431 : 3'b011;
										assign node431 = (inp[5]) ? 3'b010 : 3'b000;
				assign node435 = (inp[0]) ? node571 : node436;
					assign node436 = (inp[1]) ? node518 : node437;
						assign node437 = (inp[5]) ? node485 : node438;
							assign node438 = (inp[6]) ? node460 : node439;
								assign node439 = (inp[7]) ? node447 : node440;
									assign node440 = (inp[8]) ? 3'b000 : node441;
										assign node441 = (inp[3]) ? 3'b100 : node442;
											assign node442 = (inp[4]) ? 3'b000 : 3'b100;
									assign node447 = (inp[8]) ? node453 : node448;
										assign node448 = (inp[11]) ? node450 : 3'b000;
											assign node450 = (inp[3]) ? 3'b010 : 3'b000;
										assign node453 = (inp[3]) ? 3'b100 : node454;
											assign node454 = (inp[4]) ? node456 : 3'b010;
												assign node456 = (inp[11]) ? 3'b110 : 3'b100;
								assign node460 = (inp[3]) ? node478 : node461;
									assign node461 = (inp[7]) ? node469 : node462;
										assign node462 = (inp[8]) ? node464 : 3'b010;
											assign node464 = (inp[11]) ? node466 : 3'b010;
												assign node466 = (inp[4]) ? 3'b100 : 3'b000;
										assign node469 = (inp[11]) ? node475 : node470;
											assign node470 = (inp[8]) ? node472 : 3'b000;
												assign node472 = (inp[4]) ? 3'b100 : 3'b000;
											assign node475 = (inp[8]) ? 3'b010 : 3'b000;
									assign node478 = (inp[11]) ? 3'b010 : node479;
										assign node479 = (inp[4]) ? 3'b110 : node480;
											assign node480 = (inp[7]) ? 3'b110 : 3'b010;
							assign node485 = (inp[11]) ? node507 : node486;
								assign node486 = (inp[6]) ? node496 : node487;
									assign node487 = (inp[4]) ? 3'b000 : node488;
										assign node488 = (inp[3]) ? node490 : 3'b010;
											assign node490 = (inp[8]) ? 3'b110 : node491;
												assign node491 = (inp[7]) ? 3'b010 : 3'b110;
									assign node496 = (inp[8]) ? 3'b100 : node497;
										assign node497 = (inp[4]) ? node501 : node498;
											assign node498 = (inp[3]) ? 3'b000 : 3'b100;
											assign node501 = (inp[7]) ? node503 : 3'b000;
												assign node503 = (inp[3]) ? 3'b000 : 3'b010;
								assign node507 = (inp[4]) ? node513 : node508;
									assign node508 = (inp[7]) ? 3'b110 : node509;
										assign node509 = (inp[8]) ? 3'b010 : 3'b110;
									assign node513 = (inp[3]) ? node515 : 3'b010;
										assign node515 = (inp[7]) ? 3'b010 : 3'b110;
						assign node518 = (inp[7]) ? node552 : node519;
							assign node519 = (inp[11]) ? node539 : node520;
								assign node520 = (inp[3]) ? node530 : node521;
									assign node521 = (inp[5]) ? 3'b000 : node522;
										assign node522 = (inp[8]) ? node524 : 3'b110;
											assign node524 = (inp[6]) ? node526 : 3'b010;
												assign node526 = (inp[4]) ? 3'b010 : 3'b000;
									assign node530 = (inp[5]) ? node536 : node531;
										assign node531 = (inp[8]) ? 3'b000 : node532;
											assign node532 = (inp[4]) ? 3'b000 : 3'b100;
										assign node536 = (inp[8]) ? 3'b100 : 3'b000;
								assign node539 = (inp[5]) ? node547 : node540;
									assign node540 = (inp[4]) ? 3'b000 : node541;
										assign node541 = (inp[3]) ? node543 : 3'b100;
											assign node543 = (inp[8]) ? 3'b010 : 3'b110;
									assign node547 = (inp[3]) ? node549 : 3'b010;
										assign node549 = (inp[4]) ? 3'b010 : 3'b110;
							assign node552 = (inp[4]) ? node560 : node553;
								assign node553 = (inp[11]) ? node555 : 3'b000;
									assign node555 = (inp[5]) ? 3'b010 : node556;
										assign node556 = (inp[3]) ? 3'b010 : 3'b000;
								assign node560 = (inp[11]) ? 3'b000 : node561;
									assign node561 = (inp[6]) ? node563 : 3'b000;
										assign node563 = (inp[5]) ? 3'b000 : node564;
											assign node564 = (inp[3]) ? node566 : 3'b010;
												assign node566 = (inp[8]) ? 3'b000 : 3'b010;
					assign node571 = (inp[1]) ? node591 : node572;
						assign node572 = (inp[3]) ? 3'b010 : node573;
							assign node573 = (inp[7]) ? node575 : 3'b010;
								assign node575 = (inp[8]) ? node585 : node576;
									assign node576 = (inp[6]) ? node578 : 3'b000;
										assign node578 = (inp[4]) ? node582 : node579;
											assign node579 = (inp[5]) ? 3'b000 : 3'b010;
											assign node582 = (inp[5]) ? 3'b010 : 3'b000;
									assign node585 = (inp[4]) ? node587 : 3'b010;
										assign node587 = (inp[5]) ? 3'b010 : 3'b000;
						assign node591 = (inp[4]) ? node617 : node592;
							assign node592 = (inp[5]) ? node602 : node593;
								assign node593 = (inp[6]) ? node599 : node594;
									assign node594 = (inp[11]) ? 3'b000 : node595;
										assign node595 = (inp[3]) ? 3'b000 : 3'b100;
									assign node599 = (inp[3]) ? 3'b010 : 3'b000;
								assign node602 = (inp[7]) ? node608 : node603;
									assign node603 = (inp[3]) ? 3'b010 : node604;
										assign node604 = (inp[8]) ? 3'b010 : 3'b110;
									assign node608 = (inp[11]) ? 3'b010 : node609;
										assign node609 = (inp[3]) ? node613 : node610;
											assign node610 = (inp[6]) ? 3'b010 : 3'b000;
											assign node613 = (inp[6]) ? 3'b000 : 3'b010;
							assign node617 = (inp[7]) ? node627 : node618;
								assign node618 = (inp[3]) ? 3'b010 : node619;
									assign node619 = (inp[11]) ? 3'b010 : node620;
										assign node620 = (inp[8]) ? node622 : 3'b000;
											assign node622 = (inp[6]) ? 3'b000 : 3'b100;
								assign node627 = (inp[8]) ? node629 : 3'b000;
									assign node629 = (inp[3]) ? node631 : 3'b000;
										assign node631 = (inp[6]) ? node633 : 3'b000;
											assign node633 = (inp[11]) ? 3'b000 : 3'b010;
		assign node636 = (inp[9]) ? node994 : node637;
			assign node637 = (inp[2]) ? node743 : node638;
				assign node638 = (inp[0]) ? 3'b100 : node639;
					assign node639 = (inp[1]) ? node669 : node640;
						assign node640 = (inp[3]) ? 3'b101 : node641;
							assign node641 = (inp[7]) ? node655 : node642;
								assign node642 = (inp[8]) ? node650 : node643;
									assign node643 = (inp[4]) ? node647 : node644;
										assign node644 = (inp[5]) ? 3'b000 : 3'b101;
										assign node647 = (inp[6]) ? 3'b000 : 3'b010;
									assign node650 = (inp[5]) ? node652 : 3'b101;
										assign node652 = (inp[6]) ? 3'b101 : 3'b000;
								assign node655 = (inp[5]) ? node661 : node656;
									assign node656 = (inp[4]) ? node658 : 3'b010;
										assign node658 = (inp[8]) ? 3'b000 : 3'b110;
									assign node661 = (inp[11]) ? 3'b100 : node662;
										assign node662 = (inp[6]) ? node664 : 3'b100;
											assign node664 = (inp[8]) ? 3'b010 : 3'b110;
						assign node669 = (inp[3]) ? node699 : node670;
							assign node670 = (inp[5]) ? node686 : node671;
								assign node671 = (inp[11]) ? node679 : node672;
									assign node672 = (inp[6]) ? node676 : node673;
										assign node673 = (inp[7]) ? 3'b110 : 3'b010;
										assign node676 = (inp[8]) ? 3'b000 : 3'b100;
									assign node679 = (inp[7]) ? 3'b010 : node680;
										assign node680 = (inp[8]) ? 3'b110 : node681;
											assign node681 = (inp[6]) ? 3'b010 : 3'b110;
								assign node686 = (inp[11]) ? node694 : node687;
									assign node687 = (inp[6]) ? node689 : 3'b000;
										assign node689 = (inp[7]) ? node691 : 3'b110;
											assign node691 = (inp[4]) ? 3'b110 : 3'b010;
									assign node694 = (inp[7]) ? node696 : 3'b000;
										assign node696 = (inp[4]) ? 3'b100 : 3'b000;
							assign node699 = (inp[7]) ? node721 : node700;
								assign node700 = (inp[8]) ? node716 : node701;
									assign node701 = (inp[4]) ? node707 : node702;
										assign node702 = (inp[5]) ? node704 : 3'b101;
											assign node704 = (inp[6]) ? 3'b101 : 3'b000;
										assign node707 = (inp[11]) ? 3'b010 : node708;
											assign node708 = (inp[5]) ? node712 : node709;
												assign node709 = (inp[6]) ? 3'b000 : 3'b010;
												assign node712 = (inp[6]) ? 3'b010 : 3'b000;
									assign node716 = (inp[4]) ? node718 : 3'b101;
										assign node718 = (inp[5]) ? 3'b000 : 3'b101;
								assign node721 = (inp[4]) ? node731 : node722;
									assign node722 = (inp[5]) ? node726 : node723;
										assign node723 = (inp[6]) ? 3'b000 : 3'b010;
										assign node726 = (inp[6]) ? node728 : 3'b000;
											assign node728 = (inp[11]) ? 3'b000 : 3'b010;
									assign node731 = (inp[8]) ? node737 : node732;
										assign node732 = (inp[6]) ? 3'b100 : node733;
											assign node733 = (inp[5]) ? 3'b100 : 3'b110;
										assign node737 = (inp[11]) ? 3'b100 : node738;
											assign node738 = (inp[5]) ? 3'b010 : 3'b000;
				assign node743 = (inp[1]) ? node857 : node744;
					assign node744 = (inp[0]) ? node820 : node745;
						assign node745 = (inp[11]) ? node787 : node746;
							assign node746 = (inp[7]) ? node766 : node747;
								assign node747 = (inp[4]) ? node755 : node748;
									assign node748 = (inp[6]) ? node752 : node749;
										assign node749 = (inp[5]) ? 3'b000 : 3'b110;
										assign node752 = (inp[5]) ? 3'b110 : 3'b100;
									assign node755 = (inp[3]) ? node759 : node756;
										assign node756 = (inp[5]) ? 3'b110 : 3'b010;
										assign node759 = (inp[8]) ? 3'b100 : node760;
											assign node760 = (inp[5]) ? 3'b000 : node761;
												assign node761 = (inp[6]) ? 3'b000 : 3'b010;
								assign node766 = (inp[8]) ? node776 : node767;
									assign node767 = (inp[3]) ? 3'b110 : node768;
										assign node768 = (inp[4]) ? node772 : node769;
											assign node769 = (inp[5]) ? 3'b010 : 3'b110;
											assign node772 = (inp[5]) ? 3'b110 : 3'b000;
									assign node776 = (inp[6]) ? node782 : node777;
										assign node777 = (inp[4]) ? 3'b010 : node778;
											assign node778 = (inp[3]) ? 3'b010 : 3'b110;
										assign node782 = (inp[4]) ? node784 : 3'b010;
											assign node784 = (inp[5]) ? 3'b000 : 3'b010;
							assign node787 = (inp[5]) ? node807 : node788;
								assign node788 = (inp[7]) ? node798 : node789;
									assign node789 = (inp[8]) ? 3'b110 : node790;
										assign node790 = (inp[3]) ? node794 : node791;
											assign node791 = (inp[4]) ? 3'b100 : 3'b000;
											assign node794 = (inp[4]) ? 3'b010 : 3'b110;
									assign node798 = (inp[8]) ? node804 : node799;
										assign node799 = (inp[4]) ? node801 : 3'b000;
											assign node801 = (inp[6]) ? 3'b100 : 3'b010;
										assign node804 = (inp[6]) ? 3'b010 : 3'b000;
								assign node807 = (inp[4]) ? node815 : node808;
									assign node808 = (inp[3]) ? node810 : 3'b000;
										assign node810 = (inp[8]) ? node812 : 3'b000;
											assign node812 = (inp[7]) ? 3'b000 : 3'b100;
									assign node815 = (inp[7]) ? 3'b100 : node816;
										assign node816 = (inp[3]) ? 3'b000 : 3'b100;
						assign node820 = (inp[3]) ? 3'b100 : node821;
							assign node821 = (inp[8]) ? node839 : node822;
								assign node822 = (inp[5]) ? node834 : node823;
									assign node823 = (inp[7]) ? node831 : node824;
										assign node824 = (inp[4]) ? node826 : 3'b100;
											assign node826 = (inp[6]) ? node828 : 3'b010;
												assign node828 = (inp[11]) ? 3'b010 : 3'b000;
										assign node831 = (inp[4]) ? 3'b110 : 3'b010;
									assign node834 = (inp[7]) ? 3'b100 : node835;
										assign node835 = (inp[4]) ? 3'b010 : 3'b000;
								assign node839 = (inp[7]) ? node849 : node840;
									assign node840 = (inp[5]) ? node842 : 3'b100;
										assign node842 = (inp[4]) ? node844 : 3'b100;
											assign node844 = (inp[6]) ? node846 : 3'b000;
												assign node846 = (inp[11]) ? 3'b000 : 3'b100;
									assign node849 = (inp[5]) ? node851 : 3'b010;
										assign node851 = (inp[11]) ? node853 : 3'b010;
											assign node853 = (inp[4]) ? 3'b100 : 3'b000;
					assign node857 = (inp[7]) ? node933 : node858;
						assign node858 = (inp[4]) ? node904 : node859;
							assign node859 = (inp[0]) ? node883 : node860;
								assign node860 = (inp[3]) ? node870 : node861;
									assign node861 = (inp[5]) ? node863 : 3'b000;
										assign node863 = (inp[8]) ? node867 : node864;
											assign node864 = (inp[6]) ? 3'b000 : 3'b100;
											assign node867 = (inp[6]) ? 3'b100 : 3'b000;
									assign node870 = (inp[5]) ? node878 : node871;
										assign node871 = (inp[8]) ? 3'b110 : node872;
											assign node872 = (inp[6]) ? node874 : 3'b000;
												assign node874 = (inp[11]) ? 3'b010 : 3'b110;
										assign node878 = (inp[11]) ? 3'b100 : node879;
											assign node879 = (inp[6]) ? 3'b000 : 3'b010;
								assign node883 = (inp[3]) ? node897 : node884;
									assign node884 = (inp[8]) ? node890 : node885;
										assign node885 = (inp[11]) ? 3'b000 : node886;
											assign node886 = (inp[5]) ? 3'b010 : 3'b110;
										assign node890 = (inp[11]) ? 3'b110 : node891;
											assign node891 = (inp[6]) ? node893 : 3'b100;
												assign node893 = (inp[5]) ? 3'b110 : 3'b100;
									assign node897 = (inp[6]) ? 3'b100 : node898;
										assign node898 = (inp[8]) ? 3'b100 : node899;
											assign node899 = (inp[5]) ? 3'b000 : 3'b100;
							assign node904 = (inp[3]) ? node912 : node905;
								assign node905 = (inp[11]) ? node907 : 3'b010;
									assign node907 = (inp[5]) ? 3'b000 : node908;
										assign node908 = (inp[0]) ? 3'b000 : 3'b010;
								assign node912 = (inp[8]) ? node920 : node913;
									assign node913 = (inp[6]) ? 3'b000 : node914;
										assign node914 = (inp[5]) ? 3'b000 : node915;
											assign node915 = (inp[0]) ? 3'b010 : 3'b000;
									assign node920 = (inp[11]) ? node928 : node921;
										assign node921 = (inp[5]) ? node923 : 3'b100;
											assign node923 = (inp[0]) ? node925 : 3'b000;
												assign node925 = (inp[6]) ? 3'b100 : 3'b000;
										assign node928 = (inp[0]) ? node930 : 3'b000;
											assign node930 = (inp[5]) ? 3'b000 : 3'b100;
						assign node933 = (inp[11]) ? node977 : node934;
							assign node934 = (inp[4]) ? node964 : node935;
								assign node935 = (inp[3]) ? node949 : node936;
									assign node936 = (inp[8]) ? node944 : node937;
										assign node937 = (inp[0]) ? node939 : 3'b000;
											assign node939 = (inp[6]) ? node941 : 3'b000;
												assign node941 = (inp[5]) ? 3'b010 : 3'b000;
										assign node944 = (inp[0]) ? 3'b010 : node945;
											assign node945 = (inp[6]) ? 3'b000 : 3'b010;
									assign node949 = (inp[8]) ? node955 : node950;
										assign node950 = (inp[0]) ? 3'b010 : node951;
											assign node951 = (inp[5]) ? 3'b000 : 3'b010;
										assign node955 = (inp[0]) ? node957 : 3'b000;
											assign node957 = (inp[6]) ? node961 : node958;
												assign node958 = (inp[5]) ? 3'b000 : 3'b010;
												assign node961 = (inp[5]) ? 3'b010 : 3'b000;
								assign node964 = (inp[5]) ? 3'b000 : node965;
									assign node965 = (inp[3]) ? 3'b010 : node966;
										assign node966 = (inp[6]) ? node970 : node967;
											assign node967 = (inp[8]) ? 3'b000 : 3'b010;
											assign node970 = (inp[8]) ? node972 : 3'b000;
												assign node972 = (inp[0]) ? 3'b000 : 3'b010;
							assign node977 = (inp[4]) ? 3'b000 : node978;
								assign node978 = (inp[5]) ? 3'b000 : node979;
									assign node979 = (inp[8]) ? node985 : node980;
										assign node980 = (inp[6]) ? node982 : 3'b000;
											assign node982 = (inp[0]) ? 3'b000 : 3'b010;
										assign node985 = (inp[0]) ? node989 : node986;
											assign node986 = (inp[3]) ? 3'b000 : 3'b010;
											assign node989 = (inp[3]) ? 3'b010 : 3'b000;
			assign node994 = (inp[0]) ? node1218 : node995;
				assign node995 = (inp[2]) ? node1061 : node996;
					assign node996 = (inp[1]) ? node1008 : node997;
						assign node997 = (inp[7]) ? node999 : 3'b001;
							assign node999 = (inp[3]) ? 3'b001 : node1000;
								assign node1000 = (inp[5]) ? 3'b000 : node1001;
									assign node1001 = (inp[4]) ? node1003 : 3'b001;
										assign node1003 = (inp[8]) ? 3'b001 : 3'b010;
						assign node1008 = (inp[3]) ? node1046 : node1009;
							assign node1009 = (inp[5]) ? node1027 : node1010;
								assign node1010 = (inp[7]) ? node1018 : node1011;
									assign node1011 = (inp[6]) ? node1015 : node1012;
										assign node1012 = (inp[8]) ? 3'b010 : 3'b110;
										assign node1015 = (inp[11]) ? 3'b010 : 3'b000;
									assign node1018 = (inp[8]) ? node1022 : node1019;
										assign node1019 = (inp[4]) ? 3'b010 : 3'b110;
										assign node1022 = (inp[6]) ? node1024 : 3'b110;
											assign node1024 = (inp[11]) ? 3'b110 : 3'b100;
								assign node1027 = (inp[11]) ? node1037 : node1028;
									assign node1028 = (inp[6]) ? node1030 : 3'b100;
										assign node1030 = (inp[4]) ? node1034 : node1031;
											assign node1031 = (inp[7]) ? 3'b110 : 3'b010;
											assign node1034 = (inp[7]) ? 3'b010 : 3'b110;
									assign node1037 = (inp[6]) ? node1039 : 3'b100;
										assign node1039 = (inp[4]) ? node1043 : node1040;
											assign node1040 = (inp[7]) ? 3'b100 : 3'b000;
											assign node1043 = (inp[7]) ? 3'b000 : 3'b100;
							assign node1046 = (inp[7]) ? node1048 : 3'b001;
								assign node1048 = (inp[8]) ? node1056 : node1049;
									assign node1049 = (inp[5]) ? node1051 : 3'b010;
										assign node1051 = (inp[6]) ? node1053 : 3'b000;
											assign node1053 = (inp[11]) ? 3'b000 : 3'b010;
									assign node1056 = (inp[4]) ? node1058 : 3'b001;
										assign node1058 = (inp[5]) ? 3'b000 : 3'b001;
					assign node1061 = (inp[1]) ? node1149 : node1062;
						assign node1062 = (inp[11]) ? node1110 : node1063;
							assign node1063 = (inp[4]) ? node1083 : node1064;
								assign node1064 = (inp[3]) ? node1070 : node1065;
									assign node1065 = (inp[8]) ? 3'b010 : node1066;
										assign node1066 = (inp[5]) ? 3'b100 : 3'b010;
									assign node1070 = (inp[7]) ? node1078 : node1071;
										assign node1071 = (inp[6]) ? node1075 : node1072;
											assign node1072 = (inp[5]) ? 3'b100 : 3'b010;
											assign node1075 = (inp[5]) ? 3'b010 : 3'b000;
										assign node1078 = (inp[8]) ? node1080 : 3'b110;
											assign node1080 = (inp[5]) ? 3'b100 : 3'b110;
								assign node1083 = (inp[6]) ? node1099 : node1084;
									assign node1084 = (inp[5]) ? node1090 : node1085;
										assign node1085 = (inp[7]) ? 3'b110 : node1086;
											assign node1086 = (inp[8]) ? 3'b010 : 3'b110;
										assign node1090 = (inp[8]) ? node1092 : 3'b010;
											assign node1092 = (inp[3]) ? node1096 : node1093;
												assign node1093 = (inp[7]) ? 3'b110 : 3'b100;
												assign node1096 = (inp[7]) ? 3'b000 : 3'b100;
									assign node1099 = (inp[5]) ? node1105 : node1100;
										assign node1100 = (inp[8]) ? node1102 : 3'b100;
											assign node1102 = (inp[7]) ? 3'b100 : 3'b000;
										assign node1105 = (inp[3]) ? 3'b010 : node1106;
											assign node1106 = (inp[8]) ? 3'b110 : 3'b000;
							assign node1110 = (inp[5]) ? node1132 : node1111;
								assign node1111 = (inp[7]) ? node1121 : node1112;
									assign node1112 = (inp[3]) ? node1116 : node1113;
										assign node1113 = (inp[8]) ? 3'b010 : 3'b000;
										assign node1116 = (inp[8]) ? 3'b010 : node1117;
											assign node1117 = (inp[4]) ? 3'b110 : 3'b010;
									assign node1121 = (inp[3]) ? node1127 : node1122;
										assign node1122 = (inp[8]) ? node1124 : 3'b100;
											assign node1124 = (inp[4]) ? 3'b100 : 3'b000;
										assign node1127 = (inp[4]) ? node1129 : 3'b110;
											assign node1129 = (inp[8]) ? 3'b110 : 3'b000;
								assign node1132 = (inp[3]) ? node1138 : node1133;
									assign node1133 = (inp[4]) ? 3'b000 : node1134;
										assign node1134 = (inp[8]) ? 3'b000 : 3'b100;
									assign node1138 = (inp[7]) ? node1144 : node1139;
										assign node1139 = (inp[8]) ? node1141 : 3'b100;
											assign node1141 = (inp[4]) ? 3'b100 : 3'b000;
										assign node1144 = (inp[8]) ? node1146 : 3'b000;
											assign node1146 = (inp[4]) ? 3'b000 : 3'b100;
						assign node1149 = (inp[7]) ? node1189 : node1150;
							assign node1150 = (inp[5]) ? node1172 : node1151;
								assign node1151 = (inp[3]) ? node1163 : node1152;
									assign node1152 = (inp[4]) ? node1158 : node1153;
										assign node1153 = (inp[8]) ? 3'b010 : node1154;
											assign node1154 = (inp[11]) ? 3'b110 : 3'b010;
										assign node1158 = (inp[8]) ? 3'b100 : node1159;
											assign node1159 = (inp[11]) ? 3'b010 : 3'b100;
									assign node1163 = (inp[11]) ? node1167 : node1164;
										assign node1164 = (inp[4]) ? 3'b000 : 3'b010;
										assign node1167 = (inp[4]) ? 3'b010 : node1168;
											assign node1168 = (inp[8]) ? 3'b000 : 3'b100;
								assign node1172 = (inp[8]) ? node1174 : 3'b000;
									assign node1174 = (inp[4]) ? node1184 : node1175;
										assign node1175 = (inp[11]) ? node1181 : node1176;
											assign node1176 = (inp[3]) ? 3'b010 : node1177;
												assign node1177 = (inp[6]) ? 3'b100 : 3'b110;
											assign node1181 = (inp[3]) ? 3'b100 : 3'b000;
										assign node1184 = (inp[11]) ? 3'b000 : node1185;
											assign node1185 = (inp[3]) ? 3'b010 : 3'b000;
							assign node1189 = (inp[4]) ? node1207 : node1190;
								assign node1190 = (inp[8]) ? node1196 : node1191;
									assign node1191 = (inp[11]) ? 3'b000 : node1192;
										assign node1192 = (inp[3]) ? 3'b000 : 3'b010;
									assign node1196 = (inp[3]) ? node1202 : node1197;
										assign node1197 = (inp[6]) ? node1199 : 3'b000;
											assign node1199 = (inp[11]) ? 3'b000 : 3'b010;
										assign node1202 = (inp[5]) ? 3'b010 : node1203;
											assign node1203 = (inp[11]) ? 3'b010 : 3'b000;
								assign node1207 = (inp[11]) ? 3'b000 : node1208;
									assign node1208 = (inp[5]) ? 3'b000 : node1209;
										assign node1209 = (inp[6]) ? node1213 : node1210;
											assign node1210 = (inp[3]) ? 3'b000 : 3'b010;
											assign node1213 = (inp[3]) ? 3'b010 : 3'b000;
				assign node1218 = (inp[2]) ? node1220 : 3'b000;
					assign node1220 = (inp[3]) ? node1252 : node1221;
						assign node1221 = (inp[1]) ? node1229 : node1222;
							assign node1222 = (inp[4]) ? node1224 : 3'b000;
								assign node1224 = (inp[5]) ? 3'b000 : node1225;
									assign node1225 = (inp[8]) ? 3'b000 : 3'b010;
							assign node1229 = (inp[7]) ? node1245 : node1230;
								assign node1230 = (inp[8]) ? node1242 : node1231;
									assign node1231 = (inp[11]) ? node1237 : node1232;
										assign node1232 = (inp[6]) ? 3'b100 : node1233;
											assign node1233 = (inp[4]) ? 3'b010 : 3'b100;
										assign node1237 = (inp[4]) ? 3'b000 : node1238;
											assign node1238 = (inp[5]) ? 3'b100 : 3'b010;
									assign node1242 = (inp[11]) ? 3'b000 : 3'b010;
								assign node1245 = (inp[5]) ? 3'b000 : node1246;
									assign node1246 = (inp[11]) ? 3'b000 : node1247;
										assign node1247 = (inp[4]) ? 3'b000 : 3'b010;
						assign node1252 = (inp[5]) ? 3'b000 : node1253;
							assign node1253 = (inp[8]) ? 3'b000 : node1254;
								assign node1254 = (inp[6]) ? 3'b000 : node1255;
									assign node1255 = (inp[11]) ? 3'b000 : 3'b010;

endmodule