module dtc_split5_bm83 (
	input  wire [12-1:0] inp,
	output wire [3-1:0] outp
);

	wire [3-1:0] node1;
	wire [3-1:0] node2;
	wire [3-1:0] node3;
	wire [3-1:0] node4;
	wire [3-1:0] node5;
	wire [3-1:0] node6;
	wire [3-1:0] node7;
	wire [3-1:0] node8;
	wire [3-1:0] node9;
	wire [3-1:0] node10;
	wire [3-1:0] node15;
	wire [3-1:0] node16;
	wire [3-1:0] node17;
	wire [3-1:0] node20;
	wire [3-1:0] node23;
	wire [3-1:0] node24;
	wire [3-1:0] node28;
	wire [3-1:0] node29;
	wire [3-1:0] node31;
	wire [3-1:0] node33;
	wire [3-1:0] node36;
	wire [3-1:0] node37;
	wire [3-1:0] node38;
	wire [3-1:0] node42;
	wire [3-1:0] node43;
	wire [3-1:0] node46;
	wire [3-1:0] node49;
	wire [3-1:0] node50;
	wire [3-1:0] node51;
	wire [3-1:0] node52;
	wire [3-1:0] node53;
	wire [3-1:0] node57;
	wire [3-1:0] node59;
	wire [3-1:0] node62;
	wire [3-1:0] node64;
	wire [3-1:0] node67;
	wire [3-1:0] node68;
	wire [3-1:0] node69;
	wire [3-1:0] node70;
	wire [3-1:0] node73;
	wire [3-1:0] node77;
	wire [3-1:0] node78;
	wire [3-1:0] node81;
	wire [3-1:0] node82;
	wire [3-1:0] node86;
	wire [3-1:0] node87;
	wire [3-1:0] node88;
	wire [3-1:0] node89;
	wire [3-1:0] node90;
	wire [3-1:0] node94;
	wire [3-1:0] node97;
	wire [3-1:0] node98;
	wire [3-1:0] node102;
	wire [3-1:0] node103;
	wire [3-1:0] node104;
	wire [3-1:0] node105;
	wire [3-1:0] node107;
	wire [3-1:0] node111;
	wire [3-1:0] node112;
	wire [3-1:0] node114;
	wire [3-1:0] node117;
	wire [3-1:0] node118;
	wire [3-1:0] node123;
	wire [3-1:0] node124;
	wire [3-1:0] node125;
	wire [3-1:0] node126;
	wire [3-1:0] node128;
	wire [3-1:0] node132;
	wire [3-1:0] node134;
	wire [3-1:0] node135;
	wire [3-1:0] node136;
	wire [3-1:0] node138;
	wire [3-1:0] node141;
	wire [3-1:0] node145;
	wire [3-1:0] node146;
	wire [3-1:0] node147;
	wire [3-1:0] node148;
	wire [3-1:0] node149;
	wire [3-1:0] node153;
	wire [3-1:0] node154;
	wire [3-1:0] node155;
	wire [3-1:0] node158;
	wire [3-1:0] node162;
	wire [3-1:0] node164;
	wire [3-1:0] node165;
	wire [3-1:0] node169;
	wire [3-1:0] node170;
	wire [3-1:0] node174;
	wire [3-1:0] node175;
	wire [3-1:0] node176;
	wire [3-1:0] node177;
	wire [3-1:0] node178;
	wire [3-1:0] node179;
	wire [3-1:0] node180;
	wire [3-1:0] node181;
	wire [3-1:0] node184;
	wire [3-1:0] node187;
	wire [3-1:0] node188;
	wire [3-1:0] node192;
	wire [3-1:0] node193;
	wire [3-1:0] node195;
	wire [3-1:0] node198;
	wire [3-1:0] node199;
	wire [3-1:0] node203;
	wire [3-1:0] node204;
	wire [3-1:0] node206;
	wire [3-1:0] node209;
	wire [3-1:0] node210;
	wire [3-1:0] node212;
	wire [3-1:0] node215;
	wire [3-1:0] node218;
	wire [3-1:0] node219;
	wire [3-1:0] node220;
	wire [3-1:0] node221;
	wire [3-1:0] node222;
	wire [3-1:0] node226;
	wire [3-1:0] node227;
	wire [3-1:0] node231;
	wire [3-1:0] node232;
	wire [3-1:0] node233;
	wire [3-1:0] node238;
	wire [3-1:0] node240;
	wire [3-1:0] node241;
	wire [3-1:0] node242;
	wire [3-1:0] node247;
	wire [3-1:0] node248;
	wire [3-1:0] node249;
	wire [3-1:0] node250;
	wire [3-1:0] node251;
	wire [3-1:0] node252;
	wire [3-1:0] node255;
	wire [3-1:0] node258;
	wire [3-1:0] node259;
	wire [3-1:0] node263;
	wire [3-1:0] node264;
	wire [3-1:0] node265;
	wire [3-1:0] node269;
	wire [3-1:0] node272;
	wire [3-1:0] node273;
	wire [3-1:0] node274;
	wire [3-1:0] node275;
	wire [3-1:0] node278;
	wire [3-1:0] node282;
	wire [3-1:0] node283;
	wire [3-1:0] node284;
	wire [3-1:0] node288;
	wire [3-1:0] node289;
	wire [3-1:0] node293;
	wire [3-1:0] node294;
	wire [3-1:0] node295;
	wire [3-1:0] node297;
	wire [3-1:0] node298;
	wire [3-1:0] node302;
	wire [3-1:0] node303;
	wire [3-1:0] node304;
	wire [3-1:0] node307;
	wire [3-1:0] node310;
	wire [3-1:0] node312;
	wire [3-1:0] node315;
	wire [3-1:0] node316;
	wire [3-1:0] node318;
	wire [3-1:0] node321;
	wire [3-1:0] node322;
	wire [3-1:0] node324;
	wire [3-1:0] node327;
	wire [3-1:0] node330;
	wire [3-1:0] node331;
	wire [3-1:0] node332;
	wire [3-1:0] node333;
	wire [3-1:0] node334;
	wire [3-1:0] node337;
	wire [3-1:0] node339;
	wire [3-1:0] node342;
	wire [3-1:0] node343;
	wire [3-1:0] node344;
	wire [3-1:0] node346;
	wire [3-1:0] node349;
	wire [3-1:0] node350;
	wire [3-1:0] node353;
	wire [3-1:0] node356;
	wire [3-1:0] node357;
	wire [3-1:0] node358;
	wire [3-1:0] node361;
	wire [3-1:0] node364;
	wire [3-1:0] node365;
	wire [3-1:0] node369;
	wire [3-1:0] node370;
	wire [3-1:0] node371;
	wire [3-1:0] node372;
	wire [3-1:0] node373;
	wire [3-1:0] node377;
	wire [3-1:0] node378;
	wire [3-1:0] node382;
	wire [3-1:0] node383;
	wire [3-1:0] node385;
	wire [3-1:0] node388;
	wire [3-1:0] node390;
	wire [3-1:0] node393;
	wire [3-1:0] node394;
	wire [3-1:0] node395;
	wire [3-1:0] node396;
	wire [3-1:0] node400;
	wire [3-1:0] node401;
	wire [3-1:0] node405;
	wire [3-1:0] node406;
	wire [3-1:0] node408;
	wire [3-1:0] node411;
	wire [3-1:0] node413;
	wire [3-1:0] node416;
	wire [3-1:0] node417;
	wire [3-1:0] node418;
	wire [3-1:0] node419;
	wire [3-1:0] node420;
	wire [3-1:0] node421;
	wire [3-1:0] node426;
	wire [3-1:0] node427;
	wire [3-1:0] node431;
	wire [3-1:0] node432;
	wire [3-1:0] node433;
	wire [3-1:0] node434;
	wire [3-1:0] node438;
	wire [3-1:0] node440;
	wire [3-1:0] node443;
	wire [3-1:0] node444;
	wire [3-1:0] node446;
	wire [3-1:0] node449;
	wire [3-1:0] node452;
	wire [3-1:0] node454;
	wire [3-1:0] node455;
	wire [3-1:0] node458;
	wire [3-1:0] node459;
	wire [3-1:0] node463;
	wire [3-1:0] node464;
	wire [3-1:0] node465;
	wire [3-1:0] node466;
	wire [3-1:0] node467;
	wire [3-1:0] node468;
	wire [3-1:0] node469;
	wire [3-1:0] node470;
	wire [3-1:0] node471;
	wire [3-1:0] node475;
	wire [3-1:0] node476;
	wire [3-1:0] node480;
	wire [3-1:0] node481;
	wire [3-1:0] node482;
	wire [3-1:0] node486;
	wire [3-1:0] node488;
	wire [3-1:0] node491;
	wire [3-1:0] node492;
	wire [3-1:0] node493;
	wire [3-1:0] node494;
	wire [3-1:0] node498;
	wire [3-1:0] node501;
	wire [3-1:0] node502;
	wire [3-1:0] node505;
	wire [3-1:0] node507;
	wire [3-1:0] node510;
	wire [3-1:0] node511;
	wire [3-1:0] node512;
	wire [3-1:0] node514;
	wire [3-1:0] node516;
	wire [3-1:0] node519;
	wire [3-1:0] node520;
	wire [3-1:0] node521;
	wire [3-1:0] node525;
	wire [3-1:0] node527;
	wire [3-1:0] node530;
	wire [3-1:0] node531;
	wire [3-1:0] node532;
	wire [3-1:0] node533;
	wire [3-1:0] node536;
	wire [3-1:0] node539;
	wire [3-1:0] node540;
	wire [3-1:0] node544;
	wire [3-1:0] node545;
	wire [3-1:0] node546;
	wire [3-1:0] node549;
	wire [3-1:0] node552;
	wire [3-1:0] node555;
	wire [3-1:0] node556;
	wire [3-1:0] node557;
	wire [3-1:0] node558;
	wire [3-1:0] node559;
	wire [3-1:0] node561;
	wire [3-1:0] node564;
	wire [3-1:0] node565;
	wire [3-1:0] node569;
	wire [3-1:0] node571;
	wire [3-1:0] node573;
	wire [3-1:0] node576;
	wire [3-1:0] node577;
	wire [3-1:0] node580;
	wire [3-1:0] node581;
	wire [3-1:0] node583;
	wire [3-1:0] node586;
	wire [3-1:0] node587;
	wire [3-1:0] node591;
	wire [3-1:0] node592;
	wire [3-1:0] node593;
	wire [3-1:0] node596;
	wire [3-1:0] node597;
	wire [3-1:0] node599;
	wire [3-1:0] node602;
	wire [3-1:0] node604;
	wire [3-1:0] node607;
	wire [3-1:0] node608;
	wire [3-1:0] node609;
	wire [3-1:0] node612;
	wire [3-1:0] node614;
	wire [3-1:0] node617;
	wire [3-1:0] node619;
	wire [3-1:0] node620;
	wire [3-1:0] node623;
	wire [3-1:0] node626;
	wire [3-1:0] node627;
	wire [3-1:0] node628;
	wire [3-1:0] node629;
	wire [3-1:0] node630;
	wire [3-1:0] node631;
	wire [3-1:0] node633;
	wire [3-1:0] node636;
	wire [3-1:0] node637;
	wire [3-1:0] node641;
	wire [3-1:0] node642;
	wire [3-1:0] node645;
	wire [3-1:0] node648;
	wire [3-1:0] node649;
	wire [3-1:0] node650;
	wire [3-1:0] node651;
	wire [3-1:0] node654;
	wire [3-1:0] node657;
	wire [3-1:0] node658;
	wire [3-1:0] node661;
	wire [3-1:0] node664;
	wire [3-1:0] node665;
	wire [3-1:0] node666;
	wire [3-1:0] node670;
	wire [3-1:0] node673;
	wire [3-1:0] node674;
	wire [3-1:0] node675;
	wire [3-1:0] node676;
	wire [3-1:0] node677;
	wire [3-1:0] node681;
	wire [3-1:0] node682;
	wire [3-1:0] node686;
	wire [3-1:0] node688;
	wire [3-1:0] node691;
	wire [3-1:0] node692;
	wire [3-1:0] node693;
	wire [3-1:0] node694;
	wire [3-1:0] node697;
	wire [3-1:0] node700;
	wire [3-1:0] node702;
	wire [3-1:0] node705;
	wire [3-1:0] node706;
	wire [3-1:0] node707;
	wire [3-1:0] node710;
	wire [3-1:0] node713;
	wire [3-1:0] node714;
	wire [3-1:0] node717;
	wire [3-1:0] node720;
	wire [3-1:0] node721;
	wire [3-1:0] node722;
	wire [3-1:0] node723;
	wire [3-1:0] node724;
	wire [3-1:0] node725;
	wire [3-1:0] node730;
	wire [3-1:0] node732;
	wire [3-1:0] node735;
	wire [3-1:0] node736;
	wire [3-1:0] node737;
	wire [3-1:0] node740;
	wire [3-1:0] node744;
	wire [3-1:0] node745;
	wire [3-1:0] node746;
	wire [3-1:0] node747;
	wire [3-1:0] node751;
	wire [3-1:0] node752;
	wire [3-1:0] node753;
	wire [3-1:0] node758;
	wire [3-1:0] node759;
	wire [3-1:0] node760;
	wire [3-1:0] node762;
	wire [3-1:0] node765;
	wire [3-1:0] node768;
	wire [3-1:0] node769;
	wire [3-1:0] node770;
	wire [3-1:0] node775;
	wire [3-1:0] node776;
	wire [3-1:0] node777;
	wire [3-1:0] node778;
	wire [3-1:0] node779;
	wire [3-1:0] node781;
	wire [3-1:0] node782;
	wire [3-1:0] node784;
	wire [3-1:0] node788;
	wire [3-1:0] node789;
	wire [3-1:0] node790;
	wire [3-1:0] node792;
	wire [3-1:0] node795;
	wire [3-1:0] node798;
	wire [3-1:0] node799;
	wire [3-1:0] node800;
	wire [3-1:0] node805;
	wire [3-1:0] node806;
	wire [3-1:0] node807;
	wire [3-1:0] node809;
	wire [3-1:0] node810;
	wire [3-1:0] node814;
	wire [3-1:0] node815;
	wire [3-1:0] node816;
	wire [3-1:0] node820;
	wire [3-1:0] node821;
	wire [3-1:0] node825;
	wire [3-1:0] node826;
	wire [3-1:0] node827;
	wire [3-1:0] node829;
	wire [3-1:0] node832;
	wire [3-1:0] node834;
	wire [3-1:0] node837;
	wire [3-1:0] node838;
	wire [3-1:0] node842;
	wire [3-1:0] node843;
	wire [3-1:0] node844;
	wire [3-1:0] node845;
	wire [3-1:0] node846;
	wire [3-1:0] node850;
	wire [3-1:0] node851;
	wire [3-1:0] node853;
	wire [3-1:0] node856;
	wire [3-1:0] node858;
	wire [3-1:0] node861;
	wire [3-1:0] node862;
	wire [3-1:0] node863;
	wire [3-1:0] node867;
	wire [3-1:0] node869;
	wire [3-1:0] node872;
	wire [3-1:0] node873;
	wire [3-1:0] node874;
	wire [3-1:0] node875;
	wire [3-1:0] node876;
	wire [3-1:0] node880;
	wire [3-1:0] node883;
	wire [3-1:0] node884;
	wire [3-1:0] node886;
	wire [3-1:0] node889;
	wire [3-1:0] node890;
	wire [3-1:0] node893;
	wire [3-1:0] node896;
	wire [3-1:0] node897;
	wire [3-1:0] node898;
	wire [3-1:0] node902;
	wire [3-1:0] node903;
	wire [3-1:0] node906;
	wire [3-1:0] node909;
	wire [3-1:0] node910;
	wire [3-1:0] node911;
	wire [3-1:0] node912;
	wire [3-1:0] node913;
	wire [3-1:0] node914;
	wire [3-1:0] node915;
	wire [3-1:0] node919;
	wire [3-1:0] node920;
	wire [3-1:0] node923;
	wire [3-1:0] node926;
	wire [3-1:0] node928;
	wire [3-1:0] node929;
	wire [3-1:0] node933;
	wire [3-1:0] node934;
	wire [3-1:0] node935;
	wire [3-1:0] node936;
	wire [3-1:0] node940;
	wire [3-1:0] node942;
	wire [3-1:0] node945;
	wire [3-1:0] node946;
	wire [3-1:0] node947;
	wire [3-1:0] node951;
	wire [3-1:0] node952;
	wire [3-1:0] node956;
	wire [3-1:0] node957;
	wire [3-1:0] node958;
	wire [3-1:0] node959;
	wire [3-1:0] node960;
	wire [3-1:0] node963;
	wire [3-1:0] node966;
	wire [3-1:0] node968;
	wire [3-1:0] node971;
	wire [3-1:0] node972;
	wire [3-1:0] node973;
	wire [3-1:0] node977;
	wire [3-1:0] node979;
	wire [3-1:0] node982;
	wire [3-1:0] node983;
	wire [3-1:0] node984;
	wire [3-1:0] node985;
	wire [3-1:0] node989;
	wire [3-1:0] node991;
	wire [3-1:0] node994;
	wire [3-1:0] node995;
	wire [3-1:0] node996;
	wire [3-1:0] node1000;
	wire [3-1:0] node1001;
	wire [3-1:0] node1004;
	wire [3-1:0] node1007;
	wire [3-1:0] node1008;
	wire [3-1:0] node1009;
	wire [3-1:0] node1010;
	wire [3-1:0] node1011;
	wire [3-1:0] node1013;
	wire [3-1:0] node1016;
	wire [3-1:0] node1017;
	wire [3-1:0] node1020;
	wire [3-1:0] node1023;
	wire [3-1:0] node1024;
	wire [3-1:0] node1025;
	wire [3-1:0] node1028;
	wire [3-1:0] node1031;
	wire [3-1:0] node1032;
	wire [3-1:0] node1035;
	wire [3-1:0] node1038;
	wire [3-1:0] node1039;
	wire [3-1:0] node1040;
	wire [3-1:0] node1041;
	wire [3-1:0] node1045;
	wire [3-1:0] node1046;
	wire [3-1:0] node1049;
	wire [3-1:0] node1052;
	wire [3-1:0] node1053;
	wire [3-1:0] node1057;
	wire [3-1:0] node1058;
	wire [3-1:0] node1059;
	wire [3-1:0] node1060;
	wire [3-1:0] node1062;
	wire [3-1:0] node1065;
	wire [3-1:0] node1068;
	wire [3-1:0] node1069;
	wire [3-1:0] node1070;
	wire [3-1:0] node1074;
	wire [3-1:0] node1075;
	wire [3-1:0] node1078;
	wire [3-1:0] node1081;
	wire [3-1:0] node1082;
	wire [3-1:0] node1085;
	wire [3-1:0] node1086;
	wire [3-1:0] node1088;
	wire [3-1:0] node1091;
	wire [3-1:0] node1092;
	wire [3-1:0] node1096;
	wire [3-1:0] node1097;
	wire [3-1:0] node1098;
	wire [3-1:0] node1099;
	wire [3-1:0] node1100;
	wire [3-1:0] node1101;
	wire [3-1:0] node1102;
	wire [3-1:0] node1103;
	wire [3-1:0] node1104;
	wire [3-1:0] node1105;
	wire [3-1:0] node1109;
	wire [3-1:0] node1111;
	wire [3-1:0] node1114;
	wire [3-1:0] node1115;
	wire [3-1:0] node1119;
	wire [3-1:0] node1120;
	wire [3-1:0] node1121;
	wire [3-1:0] node1122;
	wire [3-1:0] node1125;
	wire [3-1:0] node1129;
	wire [3-1:0] node1130;
	wire [3-1:0] node1132;
	wire [3-1:0] node1135;
	wire [3-1:0] node1136;
	wire [3-1:0] node1140;
	wire [3-1:0] node1141;
	wire [3-1:0] node1142;
	wire [3-1:0] node1143;
	wire [3-1:0] node1146;
	wire [3-1:0] node1149;
	wire [3-1:0] node1150;
	wire [3-1:0] node1151;
	wire [3-1:0] node1156;
	wire [3-1:0] node1157;
	wire [3-1:0] node1158;
	wire [3-1:0] node1161;
	wire [3-1:0] node1162;
	wire [3-1:0] node1166;
	wire [3-1:0] node1167;
	wire [3-1:0] node1170;
	wire [3-1:0] node1172;
	wire [3-1:0] node1175;
	wire [3-1:0] node1176;
	wire [3-1:0] node1177;
	wire [3-1:0] node1178;
	wire [3-1:0] node1180;
	wire [3-1:0] node1182;
	wire [3-1:0] node1185;
	wire [3-1:0] node1186;
	wire [3-1:0] node1189;
	wire [3-1:0] node1191;
	wire [3-1:0] node1194;
	wire [3-1:0] node1195;
	wire [3-1:0] node1196;
	wire [3-1:0] node1199;
	wire [3-1:0] node1202;
	wire [3-1:0] node1203;
	wire [3-1:0] node1204;
	wire [3-1:0] node1207;
	wire [3-1:0] node1210;
	wire [3-1:0] node1212;
	wire [3-1:0] node1215;
	wire [3-1:0] node1216;
	wire [3-1:0] node1217;
	wire [3-1:0] node1219;
	wire [3-1:0] node1220;
	wire [3-1:0] node1225;
	wire [3-1:0] node1226;
	wire [3-1:0] node1227;
	wire [3-1:0] node1228;
	wire [3-1:0] node1232;
	wire [3-1:0] node1233;
	wire [3-1:0] node1237;
	wire [3-1:0] node1238;
	wire [3-1:0] node1241;
	wire [3-1:0] node1243;
	wire [3-1:0] node1246;
	wire [3-1:0] node1247;
	wire [3-1:0] node1248;
	wire [3-1:0] node1249;
	wire [3-1:0] node1250;
	wire [3-1:0] node1252;
	wire [3-1:0] node1254;
	wire [3-1:0] node1257;
	wire [3-1:0] node1259;
	wire [3-1:0] node1260;
	wire [3-1:0] node1264;
	wire [3-1:0] node1265;
	wire [3-1:0] node1266;
	wire [3-1:0] node1267;
	wire [3-1:0] node1271;
	wire [3-1:0] node1272;
	wire [3-1:0] node1275;
	wire [3-1:0] node1278;
	wire [3-1:0] node1279;
	wire [3-1:0] node1281;
	wire [3-1:0] node1285;
	wire [3-1:0] node1286;
	wire [3-1:0] node1287;
	wire [3-1:0] node1288;
	wire [3-1:0] node1292;
	wire [3-1:0] node1293;
	wire [3-1:0] node1297;
	wire [3-1:0] node1298;
	wire [3-1:0] node1299;
	wire [3-1:0] node1300;
	wire [3-1:0] node1304;
	wire [3-1:0] node1306;
	wire [3-1:0] node1309;
	wire [3-1:0] node1310;
	wire [3-1:0] node1312;
	wire [3-1:0] node1316;
	wire [3-1:0] node1317;
	wire [3-1:0] node1318;
	wire [3-1:0] node1319;
	wire [3-1:0] node1320;
	wire [3-1:0] node1322;
	wire [3-1:0] node1325;
	wire [3-1:0] node1328;
	wire [3-1:0] node1329;
	wire [3-1:0] node1332;
	wire [3-1:0] node1334;
	wire [3-1:0] node1337;
	wire [3-1:0] node1338;
	wire [3-1:0] node1340;
	wire [3-1:0] node1341;
	wire [3-1:0] node1345;
	wire [3-1:0] node1346;
	wire [3-1:0] node1349;
	wire [3-1:0] node1352;
	wire [3-1:0] node1353;
	wire [3-1:0] node1354;
	wire [3-1:0] node1355;
	wire [3-1:0] node1357;
	wire [3-1:0] node1360;
	wire [3-1:0] node1363;
	wire [3-1:0] node1364;
	wire [3-1:0] node1365;
	wire [3-1:0] node1369;
	wire [3-1:0] node1372;
	wire [3-1:0] node1373;
	wire [3-1:0] node1374;
	wire [3-1:0] node1376;
	wire [3-1:0] node1379;
	wire [3-1:0] node1380;
	wire [3-1:0] node1384;
	wire [3-1:0] node1385;
	wire [3-1:0] node1388;
	wire [3-1:0] node1390;
	wire [3-1:0] node1393;
	wire [3-1:0] node1394;
	wire [3-1:0] node1395;
	wire [3-1:0] node1397;
	wire [3-1:0] node1399;
	wire [3-1:0] node1400;
	wire [3-1:0] node1402;
	wire [3-1:0] node1405;
	wire [3-1:0] node1406;
	wire [3-1:0] node1410;
	wire [3-1:0] node1411;
	wire [3-1:0] node1412;
	wire [3-1:0] node1413;
	wire [3-1:0] node1415;
	wire [3-1:0] node1416;
	wire [3-1:0] node1420;
	wire [3-1:0] node1423;
	wire [3-1:0] node1424;
	wire [3-1:0] node1426;
	wire [3-1:0] node1427;
	wire [3-1:0] node1431;
	wire [3-1:0] node1433;
	wire [3-1:0] node1435;
	wire [3-1:0] node1438;
	wire [3-1:0] node1439;
	wire [3-1:0] node1441;
	wire [3-1:0] node1443;
	wire [3-1:0] node1446;
	wire [3-1:0] node1447;
	wire [3-1:0] node1448;
	wire [3-1:0] node1449;
	wire [3-1:0] node1452;
	wire [3-1:0] node1455;
	wire [3-1:0] node1457;
	wire [3-1:0] node1460;
	wire [3-1:0] node1462;
	wire [3-1:0] node1465;
	wire [3-1:0] node1466;
	wire [3-1:0] node1467;
	wire [3-1:0] node1468;
	wire [3-1:0] node1469;
	wire [3-1:0] node1471;
	wire [3-1:0] node1472;
	wire [3-1:0] node1475;
	wire [3-1:0] node1478;
	wire [3-1:0] node1479;
	wire [3-1:0] node1483;
	wire [3-1:0] node1484;
	wire [3-1:0] node1485;
	wire [3-1:0] node1486;
	wire [3-1:0] node1489;
	wire [3-1:0] node1492;
	wire [3-1:0] node1493;
	wire [3-1:0] node1496;
	wire [3-1:0] node1499;
	wire [3-1:0] node1502;
	wire [3-1:0] node1503;
	wire [3-1:0] node1504;
	wire [3-1:0] node1505;
	wire [3-1:0] node1506;
	wire [3-1:0] node1509;
	wire [3-1:0] node1513;
	wire [3-1:0] node1514;
	wire [3-1:0] node1516;
	wire [3-1:0] node1519;
	wire [3-1:0] node1522;
	wire [3-1:0] node1524;
	wire [3-1:0] node1526;
	wire [3-1:0] node1528;
	wire [3-1:0] node1531;
	wire [3-1:0] node1532;
	wire [3-1:0] node1533;
	wire [3-1:0] node1534;
	wire [3-1:0] node1535;
	wire [3-1:0] node1538;
	wire [3-1:0] node1539;
	wire [3-1:0] node1543;
	wire [3-1:0] node1544;
	wire [3-1:0] node1545;
	wire [3-1:0] node1550;
	wire [3-1:0] node1551;
	wire [3-1:0] node1552;
	wire [3-1:0] node1553;
	wire [3-1:0] node1556;
	wire [3-1:0] node1560;
	wire [3-1:0] node1561;
	wire [3-1:0] node1563;
	wire [3-1:0] node1566;
	wire [3-1:0] node1567;
	wire [3-1:0] node1570;
	wire [3-1:0] node1573;
	wire [3-1:0] node1574;
	wire [3-1:0] node1575;
	wire [3-1:0] node1578;
	wire [3-1:0] node1579;
	wire [3-1:0] node1580;
	wire [3-1:0] node1584;
	wire [3-1:0] node1586;
	wire [3-1:0] node1589;
	wire [3-1:0] node1590;
	wire [3-1:0] node1591;
	wire [3-1:0] node1592;
	wire [3-1:0] node1596;
	wire [3-1:0] node1599;
	wire [3-1:0] node1600;
	wire [3-1:0] node1604;
	wire [3-1:0] node1605;
	wire [3-1:0] node1606;
	wire [3-1:0] node1607;
	wire [3-1:0] node1608;
	wire [3-1:0] node1610;
	wire [3-1:0] node1611;
	wire [3-1:0] node1613;
	wire [3-1:0] node1618;
	wire [3-1:0] node1619;
	wire [3-1:0] node1621;
	wire [3-1:0] node1622;
	wire [3-1:0] node1624;
	wire [3-1:0] node1627;
	wire [3-1:0] node1628;
	wire [3-1:0] node1629;
	wire [3-1:0] node1634;
	wire [3-1:0] node1635;
	wire [3-1:0] node1636;
	wire [3-1:0] node1637;
	wire [3-1:0] node1639;
	wire [3-1:0] node1643;
	wire [3-1:0] node1644;
	wire [3-1:0] node1646;
	wire [3-1:0] node1650;
	wire [3-1:0] node1651;
	wire [3-1:0] node1652;
	wire [3-1:0] node1653;
	wire [3-1:0] node1657;
	wire [3-1:0] node1658;
	wire [3-1:0] node1662;
	wire [3-1:0] node1663;
	wire [3-1:0] node1664;
	wire [3-1:0] node1668;
	wire [3-1:0] node1670;
	wire [3-1:0] node1673;
	wire [3-1:0] node1674;
	wire [3-1:0] node1675;
	wire [3-1:0] node1676;
	wire [3-1:0] node1677;
	wire [3-1:0] node1678;
	wire [3-1:0] node1680;
	wire [3-1:0] node1684;
	wire [3-1:0] node1685;
	wire [3-1:0] node1686;
	wire [3-1:0] node1691;
	wire [3-1:0] node1692;
	wire [3-1:0] node1693;
	wire [3-1:0] node1695;
	wire [3-1:0] node1698;
	wire [3-1:0] node1699;
	wire [3-1:0] node1702;
	wire [3-1:0] node1705;
	wire [3-1:0] node1706;
	wire [3-1:0] node1708;
	wire [3-1:0] node1711;
	wire [3-1:0] node1712;
	wire [3-1:0] node1716;
	wire [3-1:0] node1717;
	wire [3-1:0] node1719;
	wire [3-1:0] node1720;
	wire [3-1:0] node1721;
	wire [3-1:0] node1726;
	wire [3-1:0] node1727;
	wire [3-1:0] node1729;
	wire [3-1:0] node1730;
	wire [3-1:0] node1735;
	wire [3-1:0] node1736;
	wire [3-1:0] node1737;
	wire [3-1:0] node1738;
	wire [3-1:0] node1739;
	wire [3-1:0] node1742;
	wire [3-1:0] node1745;
	wire [3-1:0] node1746;
	wire [3-1:0] node1749;
	wire [3-1:0] node1751;
	wire [3-1:0] node1754;
	wire [3-1:0] node1755;
	wire [3-1:0] node1757;
	wire [3-1:0] node1758;
	wire [3-1:0] node1762;
	wire [3-1:0] node1763;
	wire [3-1:0] node1764;
	wire [3-1:0] node1769;
	wire [3-1:0] node1770;
	wire [3-1:0] node1771;
	wire [3-1:0] node1772;
	wire [3-1:0] node1774;
	wire [3-1:0] node1777;
	wire [3-1:0] node1780;
	wire [3-1:0] node1781;
	wire [3-1:0] node1783;
	wire [3-1:0] node1786;
	wire [3-1:0] node1787;
	wire [3-1:0] node1791;
	wire [3-1:0] node1792;
	wire [3-1:0] node1794;
	wire [3-1:0] node1797;
	wire [3-1:0] node1798;
	wire [3-1:0] node1800;
	wire [3-1:0] node1803;
	wire [3-1:0] node1805;
	wire [3-1:0] node1808;
	wire [3-1:0] node1809;
	wire [3-1:0] node1810;
	wire [3-1:0] node1811;
	wire [3-1:0] node1813;
	wire [3-1:0] node1815;
	wire [3-1:0] node1820;
	wire [3-1:0] node1821;
	wire [3-1:0] node1823;
	wire [3-1:0] node1824;
	wire [3-1:0] node1825;
	wire [3-1:0] node1829;
	wire [3-1:0] node1831;
	wire [3-1:0] node1833;
	wire [3-1:0] node1836;
	wire [3-1:0] node1837;
	wire [3-1:0] node1838;
	wire [3-1:0] node1839;
	wire [3-1:0] node1841;
	wire [3-1:0] node1846;
	wire [3-1:0] node1847;
	wire [3-1:0] node1848;
	wire [3-1:0] node1849;
	wire [3-1:0] node1851;
	wire [3-1:0] node1854;
	wire [3-1:0] node1856;
	wire [3-1:0] node1859;
	wire [3-1:0] node1860;
	wire [3-1:0] node1861;
	wire [3-1:0] node1865;
	wire [3-1:0] node1866;
	wire [3-1:0] node1870;
	wire [3-1:0] node1871;

	assign outp = (inp[3]) ? node1096 : node1;
		assign node1 = (inp[4]) ? node463 : node2;
			assign node2 = (inp[9]) ? node174 : node3;
				assign node3 = (inp[7]) ? node123 : node4;
					assign node4 = (inp[0]) ? node86 : node5;
						assign node5 = (inp[6]) ? node49 : node6;
							assign node6 = (inp[5]) ? node28 : node7;
								assign node7 = (inp[1]) ? node15 : node8;
									assign node8 = (inp[2]) ? 3'b101 : node9;
										assign node9 = (inp[11]) ? 3'b001 : node10;
											assign node10 = (inp[10]) ? 3'b101 : 3'b001;
									assign node15 = (inp[11]) ? node23 : node16;
										assign node16 = (inp[2]) ? node20 : node17;
											assign node17 = (inp[10]) ? 3'b001 : 3'b011;
											assign node20 = (inp[10]) ? 3'b011 : 3'b001;
										assign node23 = (inp[2]) ? 3'b101 : node24;
											assign node24 = (inp[8]) ? 3'b111 : 3'b101;
								assign node28 = (inp[2]) ? node36 : node29;
									assign node29 = (inp[8]) ? node31 : 3'b001;
										assign node31 = (inp[1]) ? node33 : 3'b001;
											assign node33 = (inp[11]) ? 3'b001 : 3'b101;
									assign node36 = (inp[1]) ? node42 : node37;
										assign node37 = (inp[11]) ? 3'b110 : node38;
											assign node38 = (inp[10]) ? 3'b001 : 3'b101;
										assign node42 = (inp[10]) ? node46 : node43;
											assign node43 = (inp[11]) ? 3'b001 : 3'b011;
											assign node46 = (inp[8]) ? 3'b001 : 3'b001;
							assign node49 = (inp[10]) ? node67 : node50;
								assign node50 = (inp[5]) ? node62 : node51;
									assign node51 = (inp[8]) ? node57 : node52;
										assign node52 = (inp[11]) ? 3'b111 : node53;
											assign node53 = (inp[1]) ? 3'b001 : 3'b101;
										assign node57 = (inp[11]) ? node59 : 3'b001;
											assign node59 = (inp[2]) ? 3'b001 : 3'b011;
									assign node62 = (inp[8]) ? node64 : 3'b011;
										assign node64 = (inp[2]) ? 3'b011 : 3'b111;
								assign node67 = (inp[5]) ? node77 : node68;
									assign node68 = (inp[8]) ? 3'b111 : node69;
										assign node69 = (inp[1]) ? node73 : node70;
											assign node70 = (inp[11]) ? 3'b011 : 3'b111;
											assign node73 = (inp[11]) ? 3'b111 : 3'b011;
									assign node77 = (inp[8]) ? node81 : node78;
										assign node78 = (inp[2]) ? 3'b011 : 3'b001;
										assign node81 = (inp[2]) ? 3'b011 : node82;
											assign node82 = (inp[11]) ? 3'b011 : 3'b111;
						assign node86 = (inp[1]) ? node102 : node87;
							assign node87 = (inp[5]) ? node97 : node88;
								assign node88 = (inp[10]) ? node94 : node89;
									assign node89 = (inp[2]) ? 3'b111 : node90;
										assign node90 = (inp[8]) ? 3'b111 : 3'b011;
									assign node94 = (inp[11]) ? 3'b111 : 3'b011;
								assign node97 = (inp[2]) ? 3'b101 : node98;
									assign node98 = (inp[8]) ? 3'b101 : 3'b001;
							assign node102 = (inp[6]) ? 3'b111 : node103;
								assign node103 = (inp[5]) ? node111 : node104;
									assign node104 = (inp[8]) ? 3'b111 : node105;
										assign node105 = (inp[11]) ? node107 : 3'b111;
											assign node107 = (inp[2]) ? 3'b111 : 3'b011;
									assign node111 = (inp[10]) ? node117 : node112;
										assign node112 = (inp[2]) ? node114 : 3'b111;
											assign node114 = (inp[8]) ? 3'b111 : 3'b011;
										assign node117 = (inp[11]) ? 3'b011 : node118;
											assign node118 = (inp[8]) ? 3'b011 : 3'b011;
					assign node123 = (inp[5]) ? node145 : node124;
						assign node124 = (inp[8]) ? node132 : node125;
							assign node125 = (inp[6]) ? 3'b111 : node126;
								assign node126 = (inp[1]) ? node128 : 3'b111;
									assign node128 = (inp[2]) ? 3'b111 : 3'b011;
							assign node132 = (inp[2]) ? node134 : 3'b111;
								assign node134 = (inp[11]) ? 3'b111 : node135;
									assign node135 = (inp[0]) ? node141 : node136;
										assign node136 = (inp[1]) ? node138 : 3'b101;
											assign node138 = (inp[6]) ? 3'b101 : 3'b001;
										assign node141 = (inp[6]) ? 3'b111 : 3'b011;
						assign node145 = (inp[6]) ? node169 : node146;
							assign node146 = (inp[0]) ? node162 : node147;
								assign node147 = (inp[1]) ? node153 : node148;
									assign node148 = (inp[8]) ? 3'b111 : node149;
										assign node149 = (inp[2]) ? 3'b111 : 3'b101;
									assign node153 = (inp[10]) ? 3'b011 : node154;
										assign node154 = (inp[2]) ? node158 : node155;
											assign node155 = (inp[8]) ? 3'b011 : 3'b101;
											assign node158 = (inp[8]) ? 3'b111 : 3'b011;
								assign node162 = (inp[1]) ? node164 : 3'b011;
									assign node164 = (inp[2]) ? 3'b011 : node165;
										assign node165 = (inp[8]) ? 3'b011 : 3'b111;
							assign node169 = (inp[1]) ? 3'b111 : node170;
								assign node170 = (inp[0]) ? 3'b011 : 3'b111;
				assign node174 = (inp[6]) ? node330 : node175;
					assign node175 = (inp[0]) ? node247 : node176;
						assign node176 = (inp[5]) ? node218 : node177;
							assign node177 = (inp[1]) ? node203 : node178;
								assign node178 = (inp[11]) ? node192 : node179;
									assign node179 = (inp[8]) ? node187 : node180;
										assign node180 = (inp[2]) ? node184 : node181;
											assign node181 = (inp[10]) ? 3'b110 : 3'b000;
											assign node184 = (inp[10]) ? 3'b001 : 3'b101;
										assign node187 = (inp[10]) ? 3'b001 : node188;
											assign node188 = (inp[7]) ? 3'b101 : 3'b001;
									assign node192 = (inp[10]) ? node198 : node193;
										assign node193 = (inp[7]) ? node195 : 3'b110;
											assign node195 = (inp[8]) ? 3'b101 : 3'b001;
										assign node198 = (inp[7]) ? 3'b110 : node199;
											assign node199 = (inp[8]) ? 3'b010 : 3'b010;
								assign node203 = (inp[10]) ? node209 : node204;
									assign node204 = (inp[11]) ? node206 : 3'b101;
										assign node206 = (inp[7]) ? 3'b101 : 3'b001;
									assign node209 = (inp[11]) ? node215 : node210;
										assign node210 = (inp[7]) ? node212 : 3'b001;
											assign node212 = (inp[2]) ? 3'b101 : 3'b001;
										assign node215 = (inp[7]) ? 3'b001 : 3'b110;
							assign node218 = (inp[10]) ? node238 : node219;
								assign node219 = (inp[7]) ? node231 : node220;
									assign node220 = (inp[11]) ? node226 : node221;
										assign node221 = (inp[8]) ? 3'b001 : node222;
											assign node222 = (inp[2]) ? 3'b110 : 3'b010;
										assign node226 = (inp[1]) ? 3'b110 : node227;
											assign node227 = (inp[2]) ? 3'b010 : 3'b010;
									assign node231 = (inp[1]) ? 3'b001 : node232;
										assign node232 = (inp[2]) ? 3'b001 : node233;
											assign node233 = (inp[8]) ? 3'b000 : 3'b110;
								assign node238 = (inp[7]) ? node240 : 3'b010;
									assign node240 = (inp[8]) ? 3'b110 : node241;
										assign node241 = (inp[2]) ? 3'b110 : node242;
											assign node242 = (inp[11]) ? 3'b010 : 3'b010;
						assign node247 = (inp[5]) ? node293 : node248;
							assign node248 = (inp[1]) ? node272 : node249;
								assign node249 = (inp[11]) ? node263 : node250;
									assign node250 = (inp[10]) ? node258 : node251;
										assign node251 = (inp[7]) ? node255 : node252;
											assign node252 = (inp[8]) ? 3'b000 : 3'b101;
											assign node255 = (inp[8]) ? 3'b001 : 3'b011;
										assign node258 = (inp[7]) ? 3'b101 : node259;
											assign node259 = (inp[2]) ? 3'b101 : 3'b001;
									assign node263 = (inp[10]) ? node269 : node264;
										assign node264 = (inp[8]) ? 3'b101 : node265;
											assign node265 = (inp[7]) ? 3'b101 : 3'b001;
										assign node269 = (inp[7]) ? 3'b101 : 3'b110;
								assign node272 = (inp[10]) ? node282 : node273;
									assign node273 = (inp[2]) ? 3'b011 : node274;
										assign node274 = (inp[7]) ? node278 : node275;
											assign node275 = (inp[11]) ? 3'b101 : 3'b011;
											assign node278 = (inp[11]) ? 3'b011 : 3'b111;
									assign node282 = (inp[2]) ? node288 : node283;
										assign node283 = (inp[7]) ? 3'b101 : node284;
											assign node284 = (inp[8]) ? 3'b101 : 3'b001;
										assign node288 = (inp[8]) ? 3'b011 : node289;
											assign node289 = (inp[7]) ? 3'b101 : 3'b001;
							assign node293 = (inp[10]) ? node315 : node294;
								assign node294 = (inp[11]) ? node302 : node295;
									assign node295 = (inp[2]) ? node297 : 3'b101;
										assign node297 = (inp[8]) ? 3'b101 : node298;
											assign node298 = (inp[7]) ? 3'b101 : 3'b001;
									assign node302 = (inp[2]) ? node310 : node303;
										assign node303 = (inp[1]) ? node307 : node304;
											assign node304 = (inp[7]) ? 3'b011 : 3'b110;
											assign node307 = (inp[8]) ? 3'b101 : 3'b001;
										assign node310 = (inp[8]) ? node312 : 3'b101;
											assign node312 = (inp[1]) ? 3'b011 : 3'b001;
								assign node315 = (inp[1]) ? node321 : node316;
									assign node316 = (inp[8]) ? node318 : 3'b110;
										assign node318 = (inp[7]) ? 3'b001 : 3'b110;
									assign node321 = (inp[11]) ? node327 : node322;
										assign node322 = (inp[7]) ? node324 : 3'b001;
											assign node324 = (inp[2]) ? 3'b101 : 3'b001;
										assign node327 = (inp[7]) ? 3'b001 : 3'b110;
					assign node330 = (inp[0]) ? node416 : node331;
						assign node331 = (inp[1]) ? node369 : node332;
							assign node332 = (inp[10]) ? node342 : node333;
								assign node333 = (inp[7]) ? node337 : node334;
									assign node334 = (inp[5]) ? 3'b001 : 3'b101;
									assign node337 = (inp[8]) ? node339 : 3'b101;
										assign node339 = (inp[5]) ? 3'b101 : 3'b111;
								assign node342 = (inp[5]) ? node356 : node343;
									assign node343 = (inp[7]) ? node349 : node344;
										assign node344 = (inp[2]) ? node346 : 3'b001;
											assign node346 = (inp[8]) ? 3'b101 : 3'b001;
										assign node349 = (inp[11]) ? node353 : node350;
											assign node350 = (inp[8]) ? 3'b001 : 3'b101;
											assign node353 = (inp[8]) ? 3'b101 : 3'b001;
									assign node356 = (inp[7]) ? node364 : node357;
										assign node357 = (inp[8]) ? node361 : node358;
											assign node358 = (inp[2]) ? 3'b110 : 3'b010;
											assign node361 = (inp[11]) ? 3'b110 : 3'b010;
										assign node364 = (inp[2]) ? 3'b001 : node365;
											assign node365 = (inp[11]) ? 3'b110 : 3'b001;
							assign node369 = (inp[10]) ? node393 : node370;
								assign node370 = (inp[7]) ? node382 : node371;
									assign node371 = (inp[5]) ? node377 : node372;
										assign node372 = (inp[8]) ? 3'b011 : node373;
											assign node373 = (inp[11]) ? 3'b001 : 3'b011;
										assign node377 = (inp[11]) ? 3'b101 : node378;
											assign node378 = (inp[8]) ? 3'b001 : 3'b101;
									assign node382 = (inp[5]) ? node388 : node383;
										assign node383 = (inp[8]) ? node385 : 3'b111;
											assign node385 = (inp[11]) ? 3'b111 : 3'b001;
										assign node388 = (inp[11]) ? node390 : 3'b011;
											assign node390 = (inp[8]) ? 3'b011 : 3'b001;
								assign node393 = (inp[5]) ? node405 : node394;
									assign node394 = (inp[11]) ? node400 : node395;
										assign node395 = (inp[7]) ? 3'b011 : node396;
											assign node396 = (inp[2]) ? 3'b011 : 3'b101;
										assign node400 = (inp[7]) ? 3'b101 : node401;
											assign node401 = (inp[8]) ? 3'b101 : 3'b001;
									assign node405 = (inp[7]) ? node411 : node406;
										assign node406 = (inp[2]) ? node408 : 3'b001;
											assign node408 = (inp[11]) ? 3'b001 : 3'b101;
										assign node411 = (inp[11]) ? node413 : 3'b101;
											assign node413 = (inp[8]) ? 3'b101 : 3'b001;
						assign node416 = (inp[7]) ? node452 : node417;
							assign node417 = (inp[5]) ? node431 : node418;
								assign node418 = (inp[11]) ? node426 : node419;
									assign node419 = (inp[1]) ? 3'b111 : node420;
										assign node420 = (inp[10]) ? 3'b011 : node421;
											assign node421 = (inp[2]) ? 3'b111 : 3'b011;
									assign node426 = (inp[1]) ? 3'b011 : node427;
										assign node427 = (inp[10]) ? 3'b101 : 3'b011;
								assign node431 = (inp[1]) ? node443 : node432;
									assign node432 = (inp[11]) ? node438 : node433;
										assign node433 = (inp[10]) ? 3'b101 : node434;
											assign node434 = (inp[8]) ? 3'b011 : 3'b001;
										assign node438 = (inp[10]) ? node440 : 3'b101;
											assign node440 = (inp[8]) ? 3'b001 : 3'b001;
									assign node443 = (inp[2]) ? node449 : node444;
										assign node444 = (inp[10]) ? node446 : 3'b011;
											assign node446 = (inp[11]) ? 3'b101 : 3'b001;
										assign node449 = (inp[10]) ? 3'b011 : 3'b111;
							assign node452 = (inp[5]) ? node454 : 3'b111;
								assign node454 = (inp[8]) ? node458 : node455;
									assign node455 = (inp[2]) ? 3'b111 : 3'b011;
									assign node458 = (inp[1]) ? 3'b111 : node459;
										assign node459 = (inp[10]) ? 3'b011 : 3'b111;
			assign node463 = (inp[0]) ? node775 : node464;
				assign node464 = (inp[11]) ? node626 : node465;
					assign node465 = (inp[5]) ? node555 : node466;
						assign node466 = (inp[9]) ? node510 : node467;
							assign node467 = (inp[2]) ? node491 : node468;
								assign node468 = (inp[1]) ? node480 : node469;
									assign node469 = (inp[6]) ? node475 : node470;
										assign node470 = (inp[7]) ? 3'b001 : node471;
											assign node471 = (inp[8]) ? 3'b001 : 3'b100;
										assign node475 = (inp[10]) ? 3'b101 : node476;
											assign node476 = (inp[7]) ? 3'b001 : 3'b101;
									assign node480 = (inp[7]) ? node486 : node481;
										assign node481 = (inp[10]) ? 3'b001 : node482;
											assign node482 = (inp[8]) ? 3'b101 : 3'b001;
										assign node486 = (inp[10]) ? node488 : 3'b000;
											assign node488 = (inp[6]) ? 3'b011 : 3'b001;
								assign node491 = (inp[10]) ? node501 : node492;
									assign node492 = (inp[1]) ? node498 : node493;
										assign node493 = (inp[7]) ? 3'b101 : node494;
											assign node494 = (inp[6]) ? 3'b011 : 3'b001;
										assign node498 = (inp[7]) ? 3'b100 : 3'b101;
									assign node501 = (inp[1]) ? node505 : node502;
										assign node502 = (inp[6]) ? 3'b101 : 3'b110;
										assign node505 = (inp[7]) ? node507 : 3'b001;
											assign node507 = (inp[8]) ? 3'b110 : 3'b001;
							assign node510 = (inp[6]) ? node530 : node511;
								assign node511 = (inp[1]) ? node519 : node512;
									assign node512 = (inp[8]) ? node514 : 3'b100;
										assign node514 = (inp[2]) ? node516 : 3'b010;
											assign node516 = (inp[7]) ? 3'b000 : 3'b000;
									assign node519 = (inp[7]) ? node525 : node520;
										assign node520 = (inp[2]) ? 3'b010 : node521;
											assign node521 = (inp[10]) ? 3'b100 : 3'b010;
										assign node525 = (inp[8]) ? node527 : 3'b010;
											assign node527 = (inp[2]) ? 3'b001 : 3'b010;
								assign node530 = (inp[1]) ? node544 : node531;
									assign node531 = (inp[7]) ? node539 : node532;
										assign node532 = (inp[8]) ? node536 : node533;
											assign node533 = (inp[10]) ? 3'b010 : 3'b110;
											assign node536 = (inp[10]) ? 3'b010 : 3'b000;
										assign node539 = (inp[10]) ? 3'b110 : node540;
											assign node540 = (inp[8]) ? 3'b001 : 3'b011;
									assign node544 = (inp[10]) ? node552 : node545;
										assign node545 = (inp[8]) ? node549 : node546;
											assign node546 = (inp[2]) ? 3'b001 : 3'b010;
											assign node549 = (inp[7]) ? 3'b101 : 3'b001;
										assign node552 = (inp[7]) ? 3'b001 : 3'b010;
						assign node555 = (inp[9]) ? node591 : node556;
							assign node556 = (inp[7]) ? node576 : node557;
								assign node557 = (inp[2]) ? node569 : node558;
									assign node558 = (inp[6]) ? node564 : node559;
										assign node559 = (inp[10]) ? node561 : 3'b110;
											assign node561 = (inp[8]) ? 3'b110 : 3'b100;
										assign node564 = (inp[8]) ? 3'b110 : node565;
											assign node565 = (inp[1]) ? 3'b010 : 3'b110;
									assign node569 = (inp[8]) ? node571 : 3'b010;
										assign node571 = (inp[10]) ? node573 : 3'b010;
											assign node573 = (inp[1]) ? 3'b110 : 3'b010;
								assign node576 = (inp[1]) ? node580 : node577;
									assign node577 = (inp[10]) ? 3'b101 : 3'b001;
									assign node580 = (inp[6]) ? node586 : node581;
										assign node581 = (inp[10]) ? node583 : 3'b001;
											assign node583 = (inp[2]) ? 3'b000 : 3'b110;
										assign node586 = (inp[10]) ? 3'b101 : node587;
											assign node587 = (inp[8]) ? 3'b110 : 3'b011;
							assign node591 = (inp[6]) ? node607 : node592;
								assign node592 = (inp[1]) ? node596 : node593;
									assign node593 = (inp[10]) ? 3'b000 : 3'b100;
									assign node596 = (inp[8]) ? node602 : node597;
										assign node597 = (inp[2]) ? node599 : 3'b100;
											assign node599 = (inp[7]) ? 3'b000 : 3'b000;
										assign node602 = (inp[2]) ? node604 : 3'b010;
											assign node604 = (inp[10]) ? 3'b010 : 3'b000;
								assign node607 = (inp[10]) ? node617 : node608;
									assign node608 = (inp[8]) ? node612 : node609;
										assign node609 = (inp[1]) ? 3'b110 : 3'b010;
										assign node612 = (inp[1]) ? node614 : 3'b110;
											assign node614 = (inp[7]) ? 3'b001 : 3'b000;
									assign node617 = (inp[7]) ? node619 : 3'b010;
										assign node619 = (inp[8]) ? node623 : node620;
											assign node620 = (inp[1]) ? 3'b010 : 3'b010;
											assign node623 = (inp[2]) ? 3'b110 : 3'b010;
					assign node626 = (inp[9]) ? node720 : node627;
						assign node627 = (inp[7]) ? node673 : node628;
							assign node628 = (inp[1]) ? node648 : node629;
								assign node629 = (inp[6]) ? node641 : node630;
									assign node630 = (inp[8]) ? node636 : node631;
										assign node631 = (inp[5]) ? node633 : 3'b010;
											assign node633 = (inp[10]) ? 3'b100 : 3'b010;
										assign node636 = (inp[10]) ? 3'b010 : node637;
											assign node637 = (inp[2]) ? 3'b110 : 3'b010;
									assign node641 = (inp[10]) ? node645 : node642;
										assign node642 = (inp[5]) ? 3'b001 : 3'b101;
										assign node645 = (inp[5]) ? 3'b110 : 3'b001;
								assign node648 = (inp[2]) ? node664 : node649;
									assign node649 = (inp[6]) ? node657 : node650;
										assign node650 = (inp[10]) ? node654 : node651;
											assign node651 = (inp[5]) ? 3'b110 : 3'b010;
											assign node654 = (inp[5]) ? 3'b010 : 3'b110;
										assign node657 = (inp[8]) ? node661 : node658;
											assign node658 = (inp[5]) ? 3'b010 : 3'b110;
											assign node661 = (inp[5]) ? 3'b110 : 3'b010;
									assign node664 = (inp[5]) ? node670 : node665;
										assign node665 = (inp[10]) ? 3'b110 : node666;
											assign node666 = (inp[8]) ? 3'b110 : 3'b010;
										assign node670 = (inp[10]) ? 3'b010 : 3'b110;
							assign node673 = (inp[1]) ? node691 : node674;
								assign node674 = (inp[10]) ? node686 : node675;
									assign node675 = (inp[5]) ? node681 : node676;
										assign node676 = (inp[8]) ? 3'b010 : node677;
											assign node677 = (inp[6]) ? 3'b010 : 3'b010;
										assign node681 = (inp[2]) ? 3'b110 : node682;
											assign node682 = (inp[6]) ? 3'b010 : 3'b110;
									assign node686 = (inp[5]) ? node688 : 3'b110;
										assign node688 = (inp[6]) ? 3'b010 : 3'b110;
								assign node691 = (inp[8]) ? node705 : node692;
									assign node692 = (inp[5]) ? node700 : node693;
										assign node693 = (inp[6]) ? node697 : node694;
											assign node694 = (inp[10]) ? 3'b000 : 3'b101;
											assign node697 = (inp[10]) ? 3'b101 : 3'b000;
										assign node700 = (inp[6]) ? node702 : 3'b000;
											assign node702 = (inp[10]) ? 3'b000 : 3'b001;
									assign node705 = (inp[2]) ? node713 : node706;
										assign node706 = (inp[6]) ? node710 : node707;
											assign node707 = (inp[5]) ? 3'b000 : 3'b000;
											assign node710 = (inp[10]) ? 3'b001 : 3'b100;
										assign node713 = (inp[6]) ? node717 : node714;
											assign node714 = (inp[5]) ? 3'b110 : 3'b001;
											assign node717 = (inp[5]) ? 3'b111 : 3'b110;
						assign node720 = (inp[6]) ? node744 : node721;
							assign node721 = (inp[1]) ? node735 : node722;
								assign node722 = (inp[5]) ? node730 : node723;
									assign node723 = (inp[10]) ? 3'b100 : node724;
										assign node724 = (inp[7]) ? 3'b010 : node725;
											assign node725 = (inp[8]) ? 3'b000 : 3'b100;
									assign node730 = (inp[8]) ? node732 : 3'b000;
										assign node732 = (inp[2]) ? 3'b100 : 3'b000;
								assign node735 = (inp[10]) ? 3'b100 : node736;
									assign node736 = (inp[7]) ? node740 : node737;
										assign node737 = (inp[5]) ? 3'b100 : 3'b010;
										assign node740 = (inp[5]) ? 3'b010 : 3'b110;
							assign node744 = (inp[5]) ? node758 : node745;
								assign node745 = (inp[10]) ? node751 : node746;
									assign node746 = (inp[7]) ? 3'b001 : node747;
										assign node747 = (inp[8]) ? 3'b110 : 3'b111;
									assign node751 = (inp[7]) ? 3'b110 : node752;
										assign node752 = (inp[8]) ? 3'b010 : node753;
											assign node753 = (inp[1]) ? 3'b010 : 3'b100;
								assign node758 = (inp[7]) ? node768 : node759;
									assign node759 = (inp[10]) ? node765 : node760;
										assign node760 = (inp[8]) ? node762 : 3'b110;
											assign node762 = (inp[1]) ? 3'b000 : 3'b010;
										assign node765 = (inp[2]) ? 3'b100 : 3'b000;
									assign node768 = (inp[10]) ? 3'b010 : node769;
										assign node769 = (inp[1]) ? 3'b001 : node770;
											assign node770 = (inp[2]) ? 3'b110 : 3'b010;
				assign node775 = (inp[6]) ? node909 : node776;
					assign node776 = (inp[9]) ? node842 : node777;
						assign node777 = (inp[5]) ? node805 : node778;
							assign node778 = (inp[7]) ? node788 : node779;
								assign node779 = (inp[8]) ? node781 : 3'b101;
									assign node781 = (inp[10]) ? 3'b001 : node782;
										assign node782 = (inp[1]) ? node784 : 3'b101;
											assign node784 = (inp[11]) ? 3'b101 : 3'b001;
								assign node788 = (inp[11]) ? node798 : node789;
									assign node789 = (inp[8]) ? node795 : node790;
										assign node790 = (inp[2]) ? node792 : 3'b011;
											assign node792 = (inp[10]) ? 3'b011 : 3'b111;
										assign node795 = (inp[1]) ? 3'b011 : 3'b001;
									assign node798 = (inp[8]) ? 3'b111 : node799;
										assign node799 = (inp[1]) ? 3'b101 : node800;
											assign node800 = (inp[2]) ? 3'b111 : 3'b000;
							assign node805 = (inp[7]) ? node825 : node806;
								assign node806 = (inp[10]) ? node814 : node807;
									assign node807 = (inp[1]) ? node809 : 3'b011;
										assign node809 = (inp[2]) ? 3'b001 : node810;
											assign node810 = (inp[8]) ? 3'b001 : 3'b000;
									assign node814 = (inp[8]) ? node820 : node815;
										assign node815 = (inp[2]) ? 3'b110 : node816;
											assign node816 = (inp[1]) ? 3'b000 : 3'b110;
										assign node820 = (inp[1]) ? 3'b001 : node821;
											assign node821 = (inp[2]) ? 3'b000 : 3'b110;
								assign node825 = (inp[10]) ? node837 : node826;
									assign node826 = (inp[1]) ? node832 : node827;
										assign node827 = (inp[11]) ? node829 : 3'b101;
											assign node829 = (inp[8]) ? 3'b101 : 3'b010;
										assign node832 = (inp[2]) ? node834 : 3'b101;
											assign node834 = (inp[8]) ? 3'b011 : 3'b011;
									assign node837 = (inp[11]) ? 3'b001 : node838;
										assign node838 = (inp[1]) ? 3'b101 : 3'b001;
						assign node842 = (inp[7]) ? node872 : node843;
							assign node843 = (inp[5]) ? node861 : node844;
								assign node844 = (inp[10]) ? node850 : node845;
									assign node845 = (inp[11]) ? 3'b110 : node846;
										assign node846 = (inp[1]) ? 3'b001 : 3'b110;
									assign node850 = (inp[1]) ? node856 : node851;
										assign node851 = (inp[11]) ? node853 : 3'b010;
											assign node853 = (inp[2]) ? 3'b010 : 3'b100;
										assign node856 = (inp[11]) ? node858 : 3'b110;
											assign node858 = (inp[2]) ? 3'b010 : 3'b010;
								assign node861 = (inp[10]) ? node867 : node862;
									assign node862 = (inp[11]) ? 3'b010 : node863;
										assign node863 = (inp[2]) ? 3'b110 : 3'b010;
									assign node867 = (inp[8]) ? node869 : 3'b100;
										assign node869 = (inp[1]) ? 3'b010 : 3'b100;
							assign node872 = (inp[1]) ? node896 : node873;
								assign node873 = (inp[11]) ? node883 : node874;
									assign node874 = (inp[10]) ? node880 : node875;
										assign node875 = (inp[5]) ? 3'b110 : node876;
											assign node876 = (inp[2]) ? 3'b110 : 3'b001;
										assign node880 = (inp[5]) ? 3'b010 : 3'b110;
									assign node883 = (inp[2]) ? node889 : node884;
										assign node884 = (inp[8]) ? node886 : 3'b100;
											assign node886 = (inp[10]) ? 3'b010 : 3'b001;
										assign node889 = (inp[8]) ? node893 : node890;
											assign node890 = (inp[5]) ? 3'b100 : 3'b010;
											assign node893 = (inp[10]) ? 3'b010 : 3'b110;
								assign node896 = (inp[2]) ? node902 : node897;
									assign node897 = (inp[8]) ? 3'b010 : node898;
										assign node898 = (inp[10]) ? 3'b110 : 3'b010;
									assign node902 = (inp[10]) ? node906 : node903;
										assign node903 = (inp[8]) ? 3'b001 : 3'b101;
										assign node906 = (inp[11]) ? 3'b010 : 3'b001;
					assign node909 = (inp[10]) ? node1007 : node910;
						assign node910 = (inp[9]) ? node956 : node911;
							assign node911 = (inp[5]) ? node933 : node912;
								assign node912 = (inp[2]) ? node926 : node913;
									assign node913 = (inp[8]) ? node919 : node914;
										assign node914 = (inp[1]) ? 3'b101 : node915;
											assign node915 = (inp[7]) ? 3'b111 : 3'b001;
										assign node919 = (inp[1]) ? node923 : node920;
											assign node920 = (inp[11]) ? 3'b101 : 3'b011;
											assign node923 = (inp[7]) ? 3'b001 : 3'b011;
									assign node926 = (inp[7]) ? node928 : 3'b011;
										assign node928 = (inp[1]) ? 3'b101 : node929;
											assign node929 = (inp[11]) ? 3'b011 : 3'b001;
								assign node933 = (inp[11]) ? node945 : node934;
									assign node934 = (inp[7]) ? node940 : node935;
										assign node935 = (inp[2]) ? 3'b011 : node936;
											assign node936 = (inp[1]) ? 3'b101 : 3'b011;
										assign node940 = (inp[1]) ? node942 : 3'b101;
											assign node942 = (inp[8]) ? 3'b011 : 3'b111;
									assign node945 = (inp[7]) ? node951 : node946;
										assign node946 = (inp[1]) ? 3'b101 : node947;
											assign node947 = (inp[8]) ? 3'b111 : 3'b101;
										assign node951 = (inp[1]) ? 3'b111 : node952;
											assign node952 = (inp[8]) ? 3'b001 : 3'b010;
							assign node956 = (inp[2]) ? node982 : node957;
								assign node957 = (inp[5]) ? node971 : node958;
									assign node958 = (inp[8]) ? node966 : node959;
										assign node959 = (inp[1]) ? node963 : node960;
											assign node960 = (inp[7]) ? 3'b101 : 3'b011;
											assign node963 = (inp[7]) ? 3'b011 : 3'b001;
										assign node966 = (inp[11]) ? node968 : 3'b011;
											assign node968 = (inp[7]) ? 3'b011 : 3'b001;
									assign node971 = (inp[7]) ? node977 : node972;
										assign node972 = (inp[1]) ? 3'b001 : node973;
											assign node973 = (inp[11]) ? 3'b111 : 3'b011;
										assign node977 = (inp[1]) ? node979 : 3'b001;
											assign node979 = (inp[8]) ? 3'b101 : 3'b001;
								assign node982 = (inp[5]) ? node994 : node983;
									assign node983 = (inp[1]) ? node989 : node984;
										assign node984 = (inp[8]) ? 3'b101 : node985;
											assign node985 = (inp[11]) ? 3'b001 : 3'b101;
										assign node989 = (inp[11]) ? node991 : 3'b011;
											assign node991 = (inp[8]) ? 3'b111 : 3'b101;
									assign node994 = (inp[7]) ? node1000 : node995;
										assign node995 = (inp[1]) ? 3'b001 : node996;
											assign node996 = (inp[8]) ? 3'b011 : 3'b111;
										assign node1000 = (inp[1]) ? node1004 : node1001;
											assign node1001 = (inp[11]) ? 3'b001 : 3'b101;
											assign node1004 = (inp[8]) ? 3'b011 : 3'b101;
						assign node1007 = (inp[2]) ? node1057 : node1008;
							assign node1008 = (inp[1]) ? node1038 : node1009;
								assign node1009 = (inp[8]) ? node1023 : node1010;
									assign node1010 = (inp[11]) ? node1016 : node1011;
										assign node1011 = (inp[9]) ? node1013 : 3'b011;
											assign node1013 = (inp[7]) ? 3'b010 : 3'b110;
										assign node1016 = (inp[5]) ? node1020 : node1017;
											assign node1017 = (inp[9]) ? 3'b001 : 3'b000;
											assign node1020 = (inp[7]) ? 3'b110 : 3'b001;
									assign node1023 = (inp[7]) ? node1031 : node1024;
										assign node1024 = (inp[5]) ? node1028 : node1025;
											assign node1025 = (inp[11]) ? 3'b110 : 3'b000;
											assign node1028 = (inp[11]) ? 3'b011 : 3'b111;
										assign node1031 = (inp[11]) ? node1035 : node1032;
											assign node1032 = (inp[5]) ? 3'b001 : 3'b101;
											assign node1035 = (inp[5]) ? 3'b101 : 3'b001;
								assign node1038 = (inp[5]) ? node1052 : node1039;
									assign node1039 = (inp[9]) ? node1045 : node1040;
										assign node1040 = (inp[8]) ? 3'b011 : node1041;
											assign node1041 = (inp[7]) ? 3'b111 : 3'b101;
										assign node1045 = (inp[11]) ? node1049 : node1046;
											assign node1046 = (inp[7]) ? 3'b101 : 3'b100;
											assign node1049 = (inp[7]) ? 3'b101 : 3'b001;
									assign node1052 = (inp[11]) ? 3'b110 : node1053;
										assign node1053 = (inp[9]) ? 3'b111 : 3'b101;
							assign node1057 = (inp[9]) ? node1081 : node1058;
								assign node1058 = (inp[5]) ? node1068 : node1059;
									assign node1059 = (inp[7]) ? node1065 : node1060;
										assign node1060 = (inp[11]) ? node1062 : 3'b010;
											assign node1062 = (inp[1]) ? 3'b011 : 3'b101;
										assign node1065 = (inp[11]) ? 3'b111 : 3'b101;
									assign node1068 = (inp[7]) ? node1074 : node1069;
										assign node1069 = (inp[1]) ? 3'b101 : node1070;
											assign node1070 = (inp[8]) ? 3'b101 : 3'b111;
										assign node1074 = (inp[11]) ? node1078 : node1075;
											assign node1075 = (inp[8]) ? 3'b011 : 3'b111;
											assign node1078 = (inp[8]) ? 3'b001 : 3'b101;
								assign node1081 = (inp[7]) ? node1085 : node1082;
									assign node1082 = (inp[5]) ? 3'b110 : 3'b001;
									assign node1085 = (inp[5]) ? node1091 : node1086;
										assign node1086 = (inp[11]) ? node1088 : 3'b101;
											assign node1088 = (inp[1]) ? 3'b101 : 3'b001;
										assign node1091 = (inp[11]) ? 3'b001 : node1092;
											assign node1092 = (inp[1]) ? 3'b001 : 3'b001;
		assign node1096 = (inp[4]) ? node1604 : node1097;
			assign node1097 = (inp[9]) ? node1393 : node1098;
				assign node1098 = (inp[6]) ? node1246 : node1099;
					assign node1099 = (inp[0]) ? node1175 : node1100;
						assign node1100 = (inp[1]) ? node1140 : node1101;
							assign node1101 = (inp[7]) ? node1119 : node1102;
								assign node1102 = (inp[5]) ? node1114 : node1103;
									assign node1103 = (inp[10]) ? node1109 : node1104;
										assign node1104 = (inp[11]) ? 3'b100 : node1105;
											assign node1105 = (inp[8]) ? 3'b000 : 3'b000;
										assign node1109 = (inp[11]) ? node1111 : 3'b100;
											assign node1111 = (inp[8]) ? 3'b100 : 3'b000;
									assign node1114 = (inp[10]) ? 3'b000 : node1115;
										assign node1115 = (inp[8]) ? 3'b100 : 3'b000;
								assign node1119 = (inp[8]) ? node1129 : node1120;
									assign node1120 = (inp[10]) ? 3'b100 : node1121;
										assign node1121 = (inp[5]) ? node1125 : node1122;
											assign node1122 = (inp[11]) ? 3'b110 : 3'b100;
											assign node1125 = (inp[11]) ? 3'b100 : 3'b110;
									assign node1129 = (inp[11]) ? node1135 : node1130;
										assign node1130 = (inp[5]) ? node1132 : 3'b000;
											assign node1132 = (inp[10]) ? 3'b000 : 3'b010;
										assign node1135 = (inp[10]) ? 3'b100 : node1136;
											assign node1136 = (inp[5]) ? 3'b100 : 3'b110;
							assign node1140 = (inp[11]) ? node1156 : node1141;
								assign node1141 = (inp[7]) ? node1149 : node1142;
									assign node1142 = (inp[10]) ? node1146 : node1143;
										assign node1143 = (inp[5]) ? 3'b010 : 3'b100;
										assign node1146 = (inp[5]) ? 3'b000 : 3'b010;
									assign node1149 = (inp[5]) ? 3'b110 : node1150;
										assign node1150 = (inp[8]) ? 3'b010 : node1151;
											assign node1151 = (inp[2]) ? 3'b010 : 3'b110;
								assign node1156 = (inp[10]) ? node1166 : node1157;
									assign node1157 = (inp[7]) ? node1161 : node1158;
										assign node1158 = (inp[5]) ? 3'b100 : 3'b010;
										assign node1161 = (inp[5]) ? 3'b000 : node1162;
											assign node1162 = (inp[2]) ? 3'b000 : 3'b100;
									assign node1166 = (inp[7]) ? node1170 : node1167;
										assign node1167 = (inp[5]) ? 3'b000 : 3'b100;
										assign node1170 = (inp[2]) ? node1172 : 3'b000;
											assign node1172 = (inp[5]) ? 3'b100 : 3'b000;
						assign node1175 = (inp[1]) ? node1215 : node1176;
							assign node1176 = (inp[2]) ? node1194 : node1177;
								assign node1177 = (inp[8]) ? node1185 : node1178;
									assign node1178 = (inp[10]) ? node1180 : 3'b010;
										assign node1180 = (inp[11]) ? node1182 : 3'b010;
											assign node1182 = (inp[5]) ? 3'b000 : 3'b100;
									assign node1185 = (inp[7]) ? node1189 : node1186;
										assign node1186 = (inp[11]) ? 3'b110 : 3'b010;
										assign node1189 = (inp[11]) ? node1191 : 3'b110;
											assign node1191 = (inp[10]) ? 3'b110 : 3'b100;
								assign node1194 = (inp[5]) ? node1202 : node1195;
									assign node1195 = (inp[7]) ? node1199 : node1196;
										assign node1196 = (inp[10]) ? 3'b100 : 3'b110;
										assign node1199 = (inp[10]) ? 3'b110 : 3'b100;
									assign node1202 = (inp[11]) ? node1210 : node1203;
										assign node1203 = (inp[10]) ? node1207 : node1204;
											assign node1204 = (inp[8]) ? 3'b000 : 3'b010;
											assign node1207 = (inp[8]) ? 3'b010 : 3'b110;
										assign node1210 = (inp[7]) ? node1212 : 3'b100;
											assign node1212 = (inp[8]) ? 3'b110 : 3'b100;
							assign node1215 = (inp[7]) ? node1225 : node1216;
								assign node1216 = (inp[2]) ? 3'b010 : node1217;
									assign node1217 = (inp[10]) ? node1219 : 3'b110;
										assign node1219 = (inp[5]) ? 3'b100 : node1220;
											assign node1220 = (inp[8]) ? 3'b110 : 3'b010;
								assign node1225 = (inp[10]) ? node1237 : node1226;
									assign node1226 = (inp[11]) ? node1232 : node1227;
										assign node1227 = (inp[8]) ? 3'b011 : node1228;
											assign node1228 = (inp[2]) ? 3'b001 : 3'b101;
										assign node1232 = (inp[5]) ? 3'b110 : node1233;
											assign node1233 = (inp[8]) ? 3'b001 : 3'b101;
									assign node1237 = (inp[11]) ? node1241 : node1238;
										assign node1238 = (inp[2]) ? 3'b101 : 3'b110;
										assign node1241 = (inp[5]) ? node1243 : 3'b110;
											assign node1243 = (inp[8]) ? 3'b110 : 3'b010;
					assign node1246 = (inp[0]) ? node1316 : node1247;
						assign node1247 = (inp[7]) ? node1285 : node1248;
							assign node1248 = (inp[1]) ? node1264 : node1249;
								assign node1249 = (inp[8]) ? node1257 : node1250;
									assign node1250 = (inp[11]) ? node1252 : 3'b100;
										assign node1252 = (inp[5]) ? node1254 : 3'b100;
											assign node1254 = (inp[2]) ? 3'b000 : 3'b000;
									assign node1257 = (inp[5]) ? node1259 : 3'b000;
										assign node1259 = (inp[10]) ? 3'b000 : node1260;
											assign node1260 = (inp[11]) ? 3'b000 : 3'b100;
								assign node1264 = (inp[5]) ? node1278 : node1265;
									assign node1265 = (inp[10]) ? node1271 : node1266;
										assign node1266 = (inp[8]) ? 3'b000 : node1267;
											assign node1267 = (inp[2]) ? 3'b000 : 3'b010;
										assign node1271 = (inp[2]) ? node1275 : node1272;
											assign node1272 = (inp[8]) ? 3'b110 : 3'b010;
											assign node1275 = (inp[11]) ? 3'b110 : 3'b000;
									assign node1278 = (inp[10]) ? 3'b010 : node1279;
										assign node1279 = (inp[11]) ? node1281 : 3'b110;
											assign node1281 = (inp[2]) ? 3'b110 : 3'b010;
							assign node1285 = (inp[10]) ? node1297 : node1286;
								assign node1286 = (inp[1]) ? node1292 : node1287;
									assign node1287 = (inp[5]) ? 3'b110 : node1288;
										assign node1288 = (inp[2]) ? 3'b101 : 3'b110;
									assign node1292 = (inp[11]) ? 3'b001 : node1293;
										assign node1293 = (inp[8]) ? 3'b111 : 3'b101;
								assign node1297 = (inp[5]) ? node1309 : node1298;
									assign node1298 = (inp[11]) ? node1304 : node1299;
										assign node1299 = (inp[1]) ? 3'b011 : node1300;
											assign node1300 = (inp[2]) ? 3'b001 : 3'b011;
										assign node1304 = (inp[2]) ? node1306 : 3'b110;
											assign node1306 = (inp[1]) ? 3'b011 : 3'b110;
									assign node1309 = (inp[11]) ? 3'b010 : node1310;
										assign node1310 = (inp[8]) ? node1312 : 3'b110;
											assign node1312 = (inp[1]) ? 3'b110 : 3'b010;
						assign node1316 = (inp[1]) ? node1352 : node1317;
							assign node1317 = (inp[7]) ? node1337 : node1318;
								assign node1318 = (inp[11]) ? node1328 : node1319;
									assign node1319 = (inp[5]) ? node1325 : node1320;
										assign node1320 = (inp[10]) ? node1322 : 3'b100;
											assign node1322 = (inp[8]) ? 3'b001 : 3'b000;
										assign node1325 = (inp[8]) ? 3'b001 : 3'b110;
									assign node1328 = (inp[10]) ? node1332 : node1329;
										assign node1329 = (inp[5]) ? 3'b110 : 3'b011;
										assign node1332 = (inp[5]) ? node1334 : 3'b110;
											assign node1334 = (inp[8]) ? 3'b010 : 3'b010;
								assign node1337 = (inp[11]) ? node1345 : node1338;
									assign node1338 = (inp[5]) ? node1340 : 3'b101;
										assign node1340 = (inp[10]) ? 3'b001 : node1341;
											assign node1341 = (inp[2]) ? 3'b101 : 3'b001;
									assign node1345 = (inp[5]) ? node1349 : node1346;
										assign node1346 = (inp[10]) ? 3'b001 : 3'b101;
										assign node1349 = (inp[10]) ? 3'b110 : 3'b001;
							assign node1352 = (inp[5]) ? node1372 : node1353;
								assign node1353 = (inp[11]) ? node1363 : node1354;
									assign node1354 = (inp[10]) ? node1360 : node1355;
										assign node1355 = (inp[8]) ? node1357 : 3'b111;
											assign node1357 = (inp[7]) ? 3'b111 : 3'b011;
										assign node1360 = (inp[8]) ? 3'b100 : 3'b111;
									assign node1363 = (inp[10]) ? node1369 : node1364;
										assign node1364 = (inp[7]) ? 3'b011 : node1365;
											assign node1365 = (inp[8]) ? 3'b001 : 3'b101;
										assign node1369 = (inp[7]) ? 3'b101 : 3'b001;
								assign node1372 = (inp[10]) ? node1384 : node1373;
									assign node1373 = (inp[7]) ? node1379 : node1374;
										assign node1374 = (inp[8]) ? node1376 : 3'b001;
											assign node1376 = (inp[2]) ? 3'b101 : 3'b001;
										assign node1379 = (inp[11]) ? 3'b101 : node1380;
											assign node1380 = (inp[8]) ? 3'b011 : 3'b101;
									assign node1384 = (inp[7]) ? node1388 : node1385;
										assign node1385 = (inp[2]) ? 3'b110 : 3'b001;
										assign node1388 = (inp[8]) ? node1390 : 3'b001;
											assign node1390 = (inp[11]) ? 3'b001 : 3'b101;
				assign node1393 = (inp[6]) ? node1465 : node1394;
					assign node1394 = (inp[0]) ? node1410 : node1395;
						assign node1395 = (inp[7]) ? node1397 : 3'b000;
							assign node1397 = (inp[1]) ? node1399 : 3'b000;
								assign node1399 = (inp[10]) ? node1405 : node1400;
									assign node1400 = (inp[5]) ? node1402 : 3'b100;
										assign node1402 = (inp[11]) ? 3'b000 : 3'b100;
									assign node1405 = (inp[5]) ? 3'b000 : node1406;
										assign node1406 = (inp[11]) ? 3'b000 : 3'b010;
						assign node1410 = (inp[10]) ? node1438 : node1411;
							assign node1411 = (inp[5]) ? node1423 : node1412;
								assign node1412 = (inp[7]) ? node1420 : node1413;
									assign node1413 = (inp[8]) ? node1415 : 3'b100;
										assign node1415 = (inp[2]) ? 3'b010 : node1416;
											assign node1416 = (inp[1]) ? 3'b010 : 3'b100;
									assign node1420 = (inp[1]) ? 3'b110 : 3'b010;
								assign node1423 = (inp[1]) ? node1431 : node1424;
									assign node1424 = (inp[8]) ? node1426 : 3'b000;
										assign node1426 = (inp[7]) ? 3'b100 : node1427;
											assign node1427 = (inp[11]) ? 3'b000 : 3'b000;
									assign node1431 = (inp[8]) ? node1433 : 3'b100;
										assign node1433 = (inp[11]) ? node1435 : 3'b010;
											assign node1435 = (inp[7]) ? 3'b100 : 3'b000;
							assign node1438 = (inp[7]) ? node1446 : node1439;
								assign node1439 = (inp[8]) ? node1441 : 3'b000;
									assign node1441 = (inp[1]) ? node1443 : 3'b000;
										assign node1443 = (inp[5]) ? 3'b000 : 3'b100;
								assign node1446 = (inp[5]) ? node1460 : node1447;
									assign node1447 = (inp[8]) ? node1455 : node1448;
										assign node1448 = (inp[1]) ? node1452 : node1449;
											assign node1449 = (inp[11]) ? 3'b000 : 3'b000;
											assign node1452 = (inp[2]) ? 3'b010 : 3'b100;
										assign node1455 = (inp[1]) ? node1457 : 3'b100;
											assign node1457 = (inp[11]) ? 3'b100 : 3'b010;
									assign node1460 = (inp[1]) ? node1462 : 3'b000;
										assign node1462 = (inp[8]) ? 3'b100 : 3'b000;
					assign node1465 = (inp[0]) ? node1531 : node1466;
						assign node1466 = (inp[5]) ? node1502 : node1467;
							assign node1467 = (inp[1]) ? node1483 : node1468;
								assign node1468 = (inp[8]) ? node1478 : node1469;
									assign node1469 = (inp[7]) ? node1471 : 3'b100;
										assign node1471 = (inp[2]) ? node1475 : node1472;
											assign node1472 = (inp[11]) ? 3'b000 : 3'b100;
											assign node1475 = (inp[10]) ? 3'b000 : 3'b010;
									assign node1478 = (inp[7]) ? 3'b100 : node1479;
										assign node1479 = (inp[10]) ? 3'b000 : 3'b100;
								assign node1483 = (inp[11]) ? node1499 : node1484;
									assign node1484 = (inp[8]) ? node1492 : node1485;
										assign node1485 = (inp[10]) ? node1489 : node1486;
											assign node1486 = (inp[2]) ? 3'b100 : 3'b000;
											assign node1489 = (inp[2]) ? 3'b000 : 3'b100;
										assign node1492 = (inp[7]) ? node1496 : node1493;
											assign node1493 = (inp[10]) ? 3'b100 : 3'b110;
											assign node1496 = (inp[10]) ? 3'b010 : 3'b100;
									assign node1499 = (inp[8]) ? 3'b110 : 3'b010;
							assign node1502 = (inp[10]) ? node1522 : node1503;
								assign node1503 = (inp[7]) ? node1513 : node1504;
									assign node1504 = (inp[11]) ? 3'b000 : node1505;
										assign node1505 = (inp[1]) ? node1509 : node1506;
											assign node1506 = (inp[2]) ? 3'b000 : 3'b000;
											assign node1509 = (inp[8]) ? 3'b100 : 3'b000;
									assign node1513 = (inp[1]) ? node1519 : node1514;
										assign node1514 = (inp[8]) ? node1516 : 3'b100;
											assign node1516 = (inp[2]) ? 3'b000 : 3'b100;
										assign node1519 = (inp[11]) ? 3'b100 : 3'b010;
								assign node1522 = (inp[1]) ? node1524 : 3'b000;
									assign node1524 = (inp[8]) ? node1526 : 3'b000;
										assign node1526 = (inp[7]) ? node1528 : 3'b000;
											assign node1528 = (inp[11]) ? 3'b000 : 3'b100;
						assign node1531 = (inp[10]) ? node1573 : node1532;
							assign node1532 = (inp[7]) ? node1550 : node1533;
								assign node1533 = (inp[5]) ? node1543 : node1534;
									assign node1534 = (inp[2]) ? node1538 : node1535;
										assign node1535 = (inp[11]) ? 3'b000 : 3'b010;
										assign node1538 = (inp[8]) ? 3'b110 : node1539;
											assign node1539 = (inp[1]) ? 3'b110 : 3'b010;
									assign node1543 = (inp[2]) ? 3'b010 : node1544;
										assign node1544 = (inp[1]) ? 3'b010 : node1545;
											assign node1545 = (inp[11]) ? 3'b110 : 3'b010;
								assign node1550 = (inp[5]) ? node1560 : node1551;
									assign node1551 = (inp[1]) ? 3'b001 : node1552;
										assign node1552 = (inp[8]) ? node1556 : node1553;
											assign node1553 = (inp[2]) ? 3'b000 : 3'b110;
											assign node1556 = (inp[11]) ? 3'b000 : 3'b001;
									assign node1560 = (inp[1]) ? node1566 : node1561;
										assign node1561 = (inp[8]) ? node1563 : 3'b010;
											assign node1563 = (inp[2]) ? 3'b110 : 3'b010;
										assign node1566 = (inp[11]) ? node1570 : node1567;
											assign node1567 = (inp[2]) ? 3'b001 : 3'b110;
											assign node1570 = (inp[8]) ? 3'b110 : 3'b000;
							assign node1573 = (inp[5]) ? node1589 : node1574;
								assign node1574 = (inp[11]) ? node1578 : node1575;
									assign node1575 = (inp[7]) ? 3'b110 : 3'b010;
									assign node1578 = (inp[1]) ? node1584 : node1579;
										assign node1579 = (inp[7]) ? 3'b010 : node1580;
											assign node1580 = (inp[8]) ? 3'b010 : 3'b100;
										assign node1584 = (inp[7]) ? node1586 : 3'b010;
											assign node1586 = (inp[8]) ? 3'b110 : 3'b010;
								assign node1589 = (inp[11]) ? node1599 : node1590;
									assign node1590 = (inp[7]) ? node1596 : node1591;
										assign node1591 = (inp[8]) ? 3'b100 : node1592;
											assign node1592 = (inp[2]) ? 3'b100 : 3'b000;
										assign node1596 = (inp[2]) ? 3'b110 : 3'b010;
									assign node1599 = (inp[7]) ? 3'b100 : node1600;
										assign node1600 = (inp[1]) ? 3'b100 : 3'b000;
			assign node1604 = (inp[9]) ? node1808 : node1605;
				assign node1605 = (inp[6]) ? node1673 : node1606;
					assign node1606 = (inp[0]) ? node1618 : node1607;
						assign node1607 = (inp[5]) ? 3'b000 : node1608;
							assign node1608 = (inp[8]) ? node1610 : 3'b000;
								assign node1610 = (inp[11]) ? 3'b000 : node1611;
									assign node1611 = (inp[7]) ? node1613 : 3'b000;
										assign node1613 = (inp[1]) ? 3'b100 : 3'b000;
						assign node1618 = (inp[7]) ? node1634 : node1619;
							assign node1619 = (inp[1]) ? node1621 : 3'b000;
								assign node1621 = (inp[11]) ? node1627 : node1622;
									assign node1622 = (inp[5]) ? node1624 : 3'b001;
										assign node1624 = (inp[10]) ? 3'b000 : 3'b100;
									assign node1627 = (inp[5]) ? 3'b000 : node1628;
										assign node1628 = (inp[10]) ? 3'b100 : node1629;
											assign node1629 = (inp[2]) ? 3'b000 : 3'b100;
							assign node1634 = (inp[1]) ? node1650 : node1635;
								assign node1635 = (inp[10]) ? node1643 : node1636;
									assign node1636 = (inp[5]) ? 3'b100 : node1637;
										assign node1637 = (inp[2]) ? node1639 : 3'b100;
											assign node1639 = (inp[8]) ? 3'b001 : 3'b000;
									assign node1643 = (inp[5]) ? 3'b000 : node1644;
										assign node1644 = (inp[11]) ? node1646 : 3'b100;
											assign node1646 = (inp[8]) ? 3'b100 : 3'b000;
								assign node1650 = (inp[8]) ? node1662 : node1651;
									assign node1651 = (inp[2]) ? node1657 : node1652;
										assign node1652 = (inp[5]) ? 3'b100 : node1653;
											assign node1653 = (inp[11]) ? 3'b100 : 3'b110;
										assign node1657 = (inp[5]) ? 3'b000 : node1658;
											assign node1658 = (inp[10]) ? 3'b110 : 3'b000;
									assign node1662 = (inp[11]) ? node1668 : node1663;
										assign node1663 = (inp[10]) ? 3'b010 : node1664;
											assign node1664 = (inp[5]) ? 3'b010 : 3'b000;
										assign node1668 = (inp[10]) ? node1670 : 3'b010;
											assign node1670 = (inp[2]) ? 3'b100 : 3'b000;
					assign node1673 = (inp[0]) ? node1735 : node1674;
						assign node1674 = (inp[10]) ? node1716 : node1675;
							assign node1675 = (inp[7]) ? node1691 : node1676;
								assign node1676 = (inp[5]) ? node1684 : node1677;
									assign node1677 = (inp[1]) ? 3'b000 : node1678;
										assign node1678 = (inp[8]) ? node1680 : 3'b000;
											assign node1680 = (inp[2]) ? 3'b000 : 3'b100;
									assign node1684 = (inp[1]) ? 3'b100 : node1685;
										assign node1685 = (inp[11]) ? 3'b000 : node1686;
											assign node1686 = (inp[2]) ? 3'b100 : 3'b000;
								assign node1691 = (inp[1]) ? node1705 : node1692;
									assign node1692 = (inp[8]) ? node1698 : node1693;
										assign node1693 = (inp[2]) ? node1695 : 3'b100;
											assign node1695 = (inp[5]) ? 3'b100 : 3'b110;
										assign node1698 = (inp[11]) ? node1702 : node1699;
											assign node1699 = (inp[2]) ? 3'b000 : 3'b000;
											assign node1702 = (inp[5]) ? 3'b100 : 3'b110;
									assign node1705 = (inp[11]) ? node1711 : node1706;
										assign node1706 = (inp[2]) ? node1708 : 3'b010;
											assign node1708 = (inp[5]) ? 3'b010 : 3'b110;
										assign node1711 = (inp[8]) ? 3'b010 : node1712;
											assign node1712 = (inp[5]) ? 3'b100 : 3'b010;
							assign node1716 = (inp[5]) ? node1726 : node1717;
								assign node1717 = (inp[7]) ? node1719 : 3'b000;
									assign node1719 = (inp[11]) ? 3'b000 : node1720;
										assign node1720 = (inp[1]) ? 3'b010 : node1721;
											assign node1721 = (inp[8]) ? 3'b010 : 3'b000;
								assign node1726 = (inp[11]) ? 3'b000 : node1727;
									assign node1727 = (inp[1]) ? node1729 : 3'b000;
										assign node1729 = (inp[8]) ? 3'b100 : node1730;
											assign node1730 = (inp[2]) ? 3'b000 : 3'b000;
						assign node1735 = (inp[7]) ? node1769 : node1736;
							assign node1736 = (inp[1]) ? node1754 : node1737;
								assign node1737 = (inp[11]) ? node1745 : node1738;
									assign node1738 = (inp[10]) ? node1742 : node1739;
										assign node1739 = (inp[5]) ? 3'b010 : 3'b000;
										assign node1742 = (inp[8]) ? 3'b010 : 3'b100;
									assign node1745 = (inp[5]) ? node1749 : node1746;
										assign node1746 = (inp[10]) ? 3'b010 : 3'b110;
										assign node1749 = (inp[10]) ? node1751 : 3'b100;
											assign node1751 = (inp[8]) ? 3'b000 : 3'b000;
								assign node1754 = (inp[10]) ? node1762 : node1755;
									assign node1755 = (inp[5]) ? node1757 : 3'b001;
										assign node1757 = (inp[11]) ? 3'b010 : node1758;
											assign node1758 = (inp[2]) ? 3'b110 : 3'b010;
									assign node1762 = (inp[8]) ? 3'b010 : node1763;
										assign node1763 = (inp[5]) ? 3'b100 : node1764;
											assign node1764 = (inp[11]) ? 3'b010 : 3'b110;
							assign node1769 = (inp[10]) ? node1791 : node1770;
								assign node1770 = (inp[5]) ? node1780 : node1771;
									assign node1771 = (inp[1]) ? node1777 : node1772;
										assign node1772 = (inp[8]) ? node1774 : 3'b110;
											assign node1774 = (inp[11]) ? 3'b110 : 3'b001;
										assign node1777 = (inp[8]) ? 3'b001 : 3'b000;
									assign node1780 = (inp[1]) ? node1786 : node1781;
										assign node1781 = (inp[2]) ? node1783 : 3'b010;
											assign node1783 = (inp[11]) ? 3'b010 : 3'b110;
										assign node1786 = (inp[11]) ? 3'b110 : node1787;
											assign node1787 = (inp[2]) ? 3'b000 : 3'b110;
								assign node1791 = (inp[5]) ? node1797 : node1792;
									assign node1792 = (inp[11]) ? node1794 : 3'b110;
										assign node1794 = (inp[1]) ? 3'b110 : 3'b010;
									assign node1797 = (inp[2]) ? node1803 : node1798;
										assign node1798 = (inp[8]) ? node1800 : 3'b100;
											assign node1800 = (inp[11]) ? 3'b000 : 3'b010;
										assign node1803 = (inp[8]) ? node1805 : 3'b010;
											assign node1805 = (inp[11]) ? 3'b010 : 3'b110;
				assign node1808 = (inp[0]) ? node1820 : node1809;
					assign node1809 = (inp[10]) ? 3'b000 : node1810;
						assign node1810 = (inp[5]) ? 3'b000 : node1811;
							assign node1811 = (inp[6]) ? node1813 : 3'b000;
								assign node1813 = (inp[7]) ? node1815 : 3'b000;
									assign node1815 = (inp[1]) ? 3'b100 : 3'b000;
					assign node1820 = (inp[1]) ? node1836 : node1821;
						assign node1821 = (inp[7]) ? node1823 : 3'b000;
							assign node1823 = (inp[5]) ? node1829 : node1824;
								assign node1824 = (inp[10]) ? 3'b000 : node1825;
									assign node1825 = (inp[11]) ? 3'b000 : 3'b010;
								assign node1829 = (inp[6]) ? node1831 : 3'b000;
									assign node1831 = (inp[8]) ? node1833 : 3'b000;
										assign node1833 = (inp[2]) ? 3'b000 : 3'b100;
						assign node1836 = (inp[6]) ? node1846 : node1837;
							assign node1837 = (inp[11]) ? 3'b000 : node1838;
								assign node1838 = (inp[5]) ? 3'b000 : node1839;
									assign node1839 = (inp[7]) ? node1841 : 3'b000;
										assign node1841 = (inp[10]) ? 3'b000 : 3'b100;
							assign node1846 = (inp[5]) ? node1870 : node1847;
								assign node1847 = (inp[7]) ? node1859 : node1848;
									assign node1848 = (inp[10]) ? node1854 : node1849;
										assign node1849 = (inp[2]) ? node1851 : 3'b100;
											assign node1851 = (inp[8]) ? 3'b000 : 3'b100;
										assign node1854 = (inp[8]) ? node1856 : 3'b000;
											assign node1856 = (inp[11]) ? 3'b000 : 3'b100;
									assign node1859 = (inp[10]) ? node1865 : node1860;
										assign node1860 = (inp[8]) ? 3'b010 : node1861;
											assign node1861 = (inp[11]) ? 3'b000 : 3'b010;
										assign node1865 = (inp[11]) ? 3'b100 : node1866;
											assign node1866 = (inp[2]) ? 3'b010 : 3'b100;
								assign node1870 = (inp[10]) ? 3'b000 : node1871;
									assign node1871 = (inp[7]) ? 3'b100 : 3'b000;

endmodule