module dtc_split875_bm59 (
	input  wire [12-1:0] inp,
	output wire [3-1:0] outp
);

	wire [3-1:0] node1;
	wire [3-1:0] node2;
	wire [3-1:0] node3;
	wire [3-1:0] node4;
	wire [3-1:0] node5;
	wire [3-1:0] node6;
	wire [3-1:0] node7;
	wire [3-1:0] node8;
	wire [3-1:0] node9;
	wire [3-1:0] node11;
	wire [3-1:0] node14;
	wire [3-1:0] node17;
	wire [3-1:0] node18;
	wire [3-1:0] node19;
	wire [3-1:0] node20;
	wire [3-1:0] node24;
	wire [3-1:0] node25;
	wire [3-1:0] node29;
	wire [3-1:0] node31;
	wire [3-1:0] node34;
	wire [3-1:0] node35;
	wire [3-1:0] node36;
	wire [3-1:0] node38;
	wire [3-1:0] node42;
	wire [3-1:0] node43;
	wire [3-1:0] node47;
	wire [3-1:0] node48;
	wire [3-1:0] node49;
	wire [3-1:0] node50;
	wire [3-1:0] node52;
	wire [3-1:0] node55;
	wire [3-1:0] node58;
	wire [3-1:0] node59;
	wire [3-1:0] node63;
	wire [3-1:0] node64;
	wire [3-1:0] node65;
	wire [3-1:0] node66;
	wire [3-1:0] node70;
	wire [3-1:0] node71;
	wire [3-1:0] node75;
	wire [3-1:0] node76;
	wire [3-1:0] node80;
	wire [3-1:0] node82;
	wire [3-1:0] node83;
	wire [3-1:0] node84;
	wire [3-1:0] node85;
	wire [3-1:0] node86;
	wire [3-1:0] node88;
	wire [3-1:0] node93;
	wire [3-1:0] node94;
	wire [3-1:0] node95;
	wire [3-1:0] node97;
	wire [3-1:0] node101;
	wire [3-1:0] node102;
	wire [3-1:0] node106;
	wire [3-1:0] node107;
	wire [3-1:0] node108;
	wire [3-1:0] node109;
	wire [3-1:0] node110;
	wire [3-1:0] node114;
	wire [3-1:0] node115;
	wire [3-1:0] node119;
	wire [3-1:0] node120;
	wire [3-1:0] node124;
	wire [3-1:0] node125;
	wire [3-1:0] node126;
	wire [3-1:0] node127;
	wire [3-1:0] node132;
	wire [3-1:0] node134;
	wire [3-1:0] node138;
	wire [3-1:0] node139;
	wire [3-1:0] node140;
	wire [3-1:0] node141;
	wire [3-1:0] node142;
	wire [3-1:0] node143;
	wire [3-1:0] node144;
	wire [3-1:0] node146;
	wire [3-1:0] node147;
	wire [3-1:0] node150;
	wire [3-1:0] node154;
	wire [3-1:0] node155;
	wire [3-1:0] node156;
	wire [3-1:0] node157;
	wire [3-1:0] node161;
	wire [3-1:0] node162;
	wire [3-1:0] node166;
	wire [3-1:0] node167;
	wire [3-1:0] node170;
	wire [3-1:0] node172;
	wire [3-1:0] node175;
	wire [3-1:0] node176;
	wire [3-1:0] node177;
	wire [3-1:0] node178;
	wire [3-1:0] node179;
	wire [3-1:0] node182;
	wire [3-1:0] node185;
	wire [3-1:0] node186;
	wire [3-1:0] node190;
	wire [3-1:0] node191;
	wire [3-1:0] node194;
	wire [3-1:0] node195;
	wire [3-1:0] node199;
	wire [3-1:0] node200;
	wire [3-1:0] node202;
	wire [3-1:0] node205;
	wire [3-1:0] node206;
	wire [3-1:0] node208;
	wire [3-1:0] node212;
	wire [3-1:0] node213;
	wire [3-1:0] node214;
	wire [3-1:0] node215;
	wire [3-1:0] node217;
	wire [3-1:0] node220;
	wire [3-1:0] node221;
	wire [3-1:0] node224;
	wire [3-1:0] node227;
	wire [3-1:0] node228;
	wire [3-1:0] node230;
	wire [3-1:0] node233;
	wire [3-1:0] node234;
	wire [3-1:0] node237;
	wire [3-1:0] node240;
	wire [3-1:0] node241;
	wire [3-1:0] node243;
	wire [3-1:0] node245;
	wire [3-1:0] node248;
	wire [3-1:0] node249;
	wire [3-1:0] node253;
	wire [3-1:0] node254;
	wire [3-1:0] node255;
	wire [3-1:0] node256;
	wire [3-1:0] node257;
	wire [3-1:0] node258;
	wire [3-1:0] node259;
	wire [3-1:0] node263;
	wire [3-1:0] node265;
	wire [3-1:0] node268;
	wire [3-1:0] node269;
	wire [3-1:0] node271;
	wire [3-1:0] node274;
	wire [3-1:0] node276;
	wire [3-1:0] node279;
	wire [3-1:0] node280;
	wire [3-1:0] node282;
	wire [3-1:0] node285;
	wire [3-1:0] node286;
	wire [3-1:0] node290;
	wire [3-1:0] node291;
	wire [3-1:0] node292;
	wire [3-1:0] node295;
	wire [3-1:0] node296;
	wire [3-1:0] node300;
	wire [3-1:0] node301;
	wire [3-1:0] node302;
	wire [3-1:0] node303;
	wire [3-1:0] node307;
	wire [3-1:0] node309;
	wire [3-1:0] node312;
	wire [3-1:0] node314;
	wire [3-1:0] node318;
	wire [3-1:0] node319;
	wire [3-1:0] node320;
	wire [3-1:0] node321;
	wire [3-1:0] node322;
	wire [3-1:0] node323;
	wire [3-1:0] node324;
	wire [3-1:0] node326;
	wire [3-1:0] node329;
	wire [3-1:0] node330;
	wire [3-1:0] node333;
	wire [3-1:0] node336;
	wire [3-1:0] node338;
	wire [3-1:0] node339;
	wire [3-1:0] node342;
	wire [3-1:0] node345;
	wire [3-1:0] node346;
	wire [3-1:0] node347;
	wire [3-1:0] node348;
	wire [3-1:0] node352;
	wire [3-1:0] node353;
	wire [3-1:0] node357;
	wire [3-1:0] node358;
	wire [3-1:0] node359;
	wire [3-1:0] node363;
	wire [3-1:0] node366;
	wire [3-1:0] node367;
	wire [3-1:0] node368;
	wire [3-1:0] node369;
	wire [3-1:0] node373;
	wire [3-1:0] node374;
	wire [3-1:0] node377;
	wire [3-1:0] node378;
	wire [3-1:0] node381;
	wire [3-1:0] node384;
	wire [3-1:0] node385;
	wire [3-1:0] node386;
	wire [3-1:0] node389;
	wire [3-1:0] node392;
	wire [3-1:0] node394;
	wire [3-1:0] node397;
	wire [3-1:0] node398;
	wire [3-1:0] node399;
	wire [3-1:0] node400;
	wire [3-1:0] node401;
	wire [3-1:0] node405;
	wire [3-1:0] node406;
	wire [3-1:0] node410;
	wire [3-1:0] node411;
	wire [3-1:0] node412;
	wire [3-1:0] node413;
	wire [3-1:0] node416;
	wire [3-1:0] node419;
	wire [3-1:0] node420;
	wire [3-1:0] node423;
	wire [3-1:0] node426;
	wire [3-1:0] node427;
	wire [3-1:0] node430;
	wire [3-1:0] node433;
	wire [3-1:0] node434;
	wire [3-1:0] node435;
	wire [3-1:0] node437;
	wire [3-1:0] node440;
	wire [3-1:0] node441;
	wire [3-1:0] node442;
	wire [3-1:0] node445;
	wire [3-1:0] node450;
	wire [3-1:0] node451;
	wire [3-1:0] node452;
	wire [3-1:0] node453;
	wire [3-1:0] node454;
	wire [3-1:0] node455;
	wire [3-1:0] node456;
	wire [3-1:0] node460;
	wire [3-1:0] node462;
	wire [3-1:0] node465;
	wire [3-1:0] node466;
	wire [3-1:0] node470;
	wire [3-1:0] node472;
	wire [3-1:0] node473;
	wire [3-1:0] node475;
	wire [3-1:0] node478;
	wire [3-1:0] node481;
	wire [3-1:0] node482;
	wire [3-1:0] node483;
	wire [3-1:0] node484;
	wire [3-1:0] node488;
	wire [3-1:0] node489;
	wire [3-1:0] node491;
	wire [3-1:0] node496;
	wire [3-1:0] node497;
	wire [3-1:0] node498;
	wire [3-1:0] node499;
	wire [3-1:0] node500;
	wire [3-1:0] node501;
	wire [3-1:0] node505;
	wire [3-1:0] node506;
	wire [3-1:0] node509;
	wire [3-1:0] node512;
	wire [3-1:0] node514;
	wire [3-1:0] node516;
	wire [3-1:0] node521;
	wire [3-1:0] node522;
	wire [3-1:0] node523;
	wire [3-1:0] node524;
	wire [3-1:0] node525;
	wire [3-1:0] node527;
	wire [3-1:0] node528;
	wire [3-1:0] node529;
	wire [3-1:0] node530;
	wire [3-1:0] node533;
	wire [3-1:0] node537;
	wire [3-1:0] node538;
	wire [3-1:0] node540;
	wire [3-1:0] node541;
	wire [3-1:0] node545;
	wire [3-1:0] node546;
	wire [3-1:0] node550;
	wire [3-1:0] node551;
	wire [3-1:0] node552;
	wire [3-1:0] node553;
	wire [3-1:0] node554;
	wire [3-1:0] node558;
	wire [3-1:0] node559;
	wire [3-1:0] node563;
	wire [3-1:0] node564;
	wire [3-1:0] node565;
	wire [3-1:0] node566;
	wire [3-1:0] node570;
	wire [3-1:0] node573;
	wire [3-1:0] node574;
	wire [3-1:0] node575;
	wire [3-1:0] node578;
	wire [3-1:0] node582;
	wire [3-1:0] node583;
	wire [3-1:0] node584;
	wire [3-1:0] node586;
	wire [3-1:0] node589;
	wire [3-1:0] node590;
	wire [3-1:0] node592;
	wire [3-1:0] node595;
	wire [3-1:0] node598;
	wire [3-1:0] node599;
	wire [3-1:0] node601;
	wire [3-1:0] node602;
	wire [3-1:0] node606;
	wire [3-1:0] node607;
	wire [3-1:0] node611;
	wire [3-1:0] node613;
	wire [3-1:0] node615;
	wire [3-1:0] node616;
	wire [3-1:0] node617;
	wire [3-1:0] node618;
	wire [3-1:0] node619;
	wire [3-1:0] node623;
	wire [3-1:0] node625;
	wire [3-1:0] node629;
	wire [3-1:0] node630;
	wire [3-1:0] node632;
	wire [3-1:0] node633;
	wire [3-1:0] node637;
	wire [3-1:0] node639;
	wire [3-1:0] node643;
	wire [3-1:0] node644;
	wire [3-1:0] node645;
	wire [3-1:0] node646;
	wire [3-1:0] node647;
	wire [3-1:0] node648;
	wire [3-1:0] node649;
	wire [3-1:0] node650;
	wire [3-1:0] node653;
	wire [3-1:0] node656;
	wire [3-1:0] node658;
	wire [3-1:0] node661;
	wire [3-1:0] node662;
	wire [3-1:0] node664;
	wire [3-1:0] node667;
	wire [3-1:0] node668;
	wire [3-1:0] node669;
	wire [3-1:0] node672;
	wire [3-1:0] node675;
	wire [3-1:0] node676;
	wire [3-1:0] node679;
	wire [3-1:0] node682;
	wire [3-1:0] node683;
	wire [3-1:0] node684;
	wire [3-1:0] node686;
	wire [3-1:0] node688;
	wire [3-1:0] node692;
	wire [3-1:0] node693;
	wire [3-1:0] node694;
	wire [3-1:0] node696;
	wire [3-1:0] node699;
	wire [3-1:0] node702;
	wire [3-1:0] node704;
	wire [3-1:0] node705;
	wire [3-1:0] node709;
	wire [3-1:0] node710;
	wire [3-1:0] node711;
	wire [3-1:0] node712;
	wire [3-1:0] node715;
	wire [3-1:0] node716;
	wire [3-1:0] node720;
	wire [3-1:0] node721;
	wire [3-1:0] node722;
	wire [3-1:0] node725;
	wire [3-1:0] node728;
	wire [3-1:0] node729;
	wire [3-1:0] node732;
	wire [3-1:0] node735;
	wire [3-1:0] node736;
	wire [3-1:0] node737;
	wire [3-1:0] node740;
	wire [3-1:0] node741;
	wire [3-1:0] node745;
	wire [3-1:0] node746;
	wire [3-1:0] node750;
	wire [3-1:0] node751;
	wire [3-1:0] node752;
	wire [3-1:0] node753;
	wire [3-1:0] node754;
	wire [3-1:0] node755;
	wire [3-1:0] node756;
	wire [3-1:0] node759;
	wire [3-1:0] node762;
	wire [3-1:0] node764;
	wire [3-1:0] node767;
	wire [3-1:0] node768;
	wire [3-1:0] node769;
	wire [3-1:0] node773;
	wire [3-1:0] node776;
	wire [3-1:0] node777;
	wire [3-1:0] node778;
	wire [3-1:0] node780;
	wire [3-1:0] node783;
	wire [3-1:0] node786;
	wire [3-1:0] node787;
	wire [3-1:0] node790;
	wire [3-1:0] node791;
	wire [3-1:0] node795;
	wire [3-1:0] node796;
	wire [3-1:0] node797;
	wire [3-1:0] node798;
	wire [3-1:0] node800;
	wire [3-1:0] node803;
	wire [3-1:0] node804;
	wire [3-1:0] node808;
	wire [3-1:0] node809;
	wire [3-1:0] node810;
	wire [3-1:0] node814;
	wire [3-1:0] node817;
	wire [3-1:0] node819;
	wire [3-1:0] node821;
	wire [3-1:0] node824;
	wire [3-1:0] node825;
	wire [3-1:0] node826;
	wire [3-1:0] node827;
	wire [3-1:0] node828;
	wire [3-1:0] node831;
	wire [3-1:0] node834;
	wire [3-1:0] node836;
	wire [3-1:0] node838;
	wire [3-1:0] node841;
	wire [3-1:0] node842;
	wire [3-1:0] node843;
	wire [3-1:0] node844;
	wire [3-1:0] node847;
	wire [3-1:0] node850;
	wire [3-1:0] node851;
	wire [3-1:0] node854;
	wire [3-1:0] node858;
	wire [3-1:0] node859;
	wire [3-1:0] node860;
	wire [3-1:0] node861;
	wire [3-1:0] node863;
	wire [3-1:0] node866;
	wire [3-1:0] node868;
	wire [3-1:0] node873;
	wire [3-1:0] node874;
	wire [3-1:0] node875;
	wire [3-1:0] node877;
	wire [3-1:0] node878;
	wire [3-1:0] node880;
	wire [3-1:0] node882;
	wire [3-1:0] node883;
	wire [3-1:0] node887;
	wire [3-1:0] node888;
	wire [3-1:0] node890;
	wire [3-1:0] node892;
	wire [3-1:0] node897;
	wire [3-1:0] node898;
	wire [3-1:0] node899;
	wire [3-1:0] node900;
	wire [3-1:0] node901;
	wire [3-1:0] node902;
	wire [3-1:0] node903;
	wire [3-1:0] node906;
	wire [3-1:0] node909;
	wire [3-1:0] node910;
	wire [3-1:0] node913;
	wire [3-1:0] node916;
	wire [3-1:0] node917;
	wire [3-1:0] node919;
	wire [3-1:0] node923;
	wire [3-1:0] node924;
	wire [3-1:0] node925;
	wire [3-1:0] node928;
	wire [3-1:0] node931;
	wire [3-1:0] node932;
	wire [3-1:0] node937;
	wire [3-1:0] node938;
	wire [3-1:0] node939;
	wire [3-1:0] node940;
	wire [3-1:0] node941;
	wire [3-1:0] node945;
	wire [3-1:0] node946;
	wire [3-1:0] node947;
	wire [3-1:0] node952;
	wire [3-1:0] node953;
	wire [3-1:0] node955;
	wire [3-1:0] node956;
	wire [3-1:0] node961;
	wire [3-1:0] node962;
	wire [3-1:0] node963;
	wire [3-1:0] node964;
	wire [3-1:0] node967;
	wire [3-1:0] node969;
	wire [3-1:0] node974;
	wire [3-1:0] node975;
	wire [3-1:0] node976;
	wire [3-1:0] node977;
	wire [3-1:0] node978;
	wire [3-1:0] node979;
	wire [3-1:0] node980;
	wire [3-1:0] node981;
	wire [3-1:0] node983;
	wire [3-1:0] node984;
	wire [3-1:0] node985;
	wire [3-1:0] node990;
	wire [3-1:0] node991;
	wire [3-1:0] node992;
	wire [3-1:0] node996;
	wire [3-1:0] node997;
	wire [3-1:0] node998;
	wire [3-1:0] node1002;
	wire [3-1:0] node1005;
	wire [3-1:0] node1006;
	wire [3-1:0] node1007;
	wire [3-1:0] node1009;
	wire [3-1:0] node1012;
	wire [3-1:0] node1013;
	wire [3-1:0] node1017;
	wire [3-1:0] node1018;
	wire [3-1:0] node1022;
	wire [3-1:0] node1023;
	wire [3-1:0] node1024;
	wire [3-1:0] node1025;
	wire [3-1:0] node1026;
	wire [3-1:0] node1030;
	wire [3-1:0] node1032;
	wire [3-1:0] node1035;
	wire [3-1:0] node1036;
	wire [3-1:0] node1037;
	wire [3-1:0] node1039;
	wire [3-1:0] node1042;
	wire [3-1:0] node1043;
	wire [3-1:0] node1047;
	wire [3-1:0] node1049;
	wire [3-1:0] node1052;
	wire [3-1:0] node1053;
	wire [3-1:0] node1055;
	wire [3-1:0] node1056;
	wire [3-1:0] node1060;
	wire [3-1:0] node1061;
	wire [3-1:0] node1065;
	wire [3-1:0] node1067;
	wire [3-1:0] node1068;
	wire [3-1:0] node1069;
	wire [3-1:0] node1070;
	wire [3-1:0] node1072;
	wire [3-1:0] node1074;
	wire [3-1:0] node1078;
	wire [3-1:0] node1079;
	wire [3-1:0] node1080;
	wire [3-1:0] node1082;
	wire [3-1:0] node1085;
	wire [3-1:0] node1088;
	wire [3-1:0] node1090;
	wire [3-1:0] node1091;
	wire [3-1:0] node1095;
	wire [3-1:0] node1096;
	wire [3-1:0] node1097;
	wire [3-1:0] node1099;
	wire [3-1:0] node1102;
	wire [3-1:0] node1103;
	wire [3-1:0] node1104;
	wire [3-1:0] node1108;
	wire [3-1:0] node1109;
	wire [3-1:0] node1113;
	wire [3-1:0] node1114;
	wire [3-1:0] node1117;
	wire [3-1:0] node1118;
	wire [3-1:0] node1119;
	wire [3-1:0] node1123;
	wire [3-1:0] node1125;
	wire [3-1:0] node1129;
	wire [3-1:0] node1130;
	wire [3-1:0] node1131;
	wire [3-1:0] node1132;
	wire [3-1:0] node1133;
	wire [3-1:0] node1134;
	wire [3-1:0] node1135;
	wire [3-1:0] node1136;
	wire [3-1:0] node1139;
	wire [3-1:0] node1141;
	wire [3-1:0] node1144;
	wire [3-1:0] node1145;
	wire [3-1:0] node1148;
	wire [3-1:0] node1151;
	wire [3-1:0] node1152;
	wire [3-1:0] node1155;
	wire [3-1:0] node1156;
	wire [3-1:0] node1158;
	wire [3-1:0] node1161;
	wire [3-1:0] node1162;
	wire [3-1:0] node1165;
	wire [3-1:0] node1168;
	wire [3-1:0] node1169;
	wire [3-1:0] node1170;
	wire [3-1:0] node1171;
	wire [3-1:0] node1172;
	wire [3-1:0] node1176;
	wire [3-1:0] node1177;
	wire [3-1:0] node1181;
	wire [3-1:0] node1183;
	wire [3-1:0] node1184;
	wire [3-1:0] node1188;
	wire [3-1:0] node1189;
	wire [3-1:0] node1190;
	wire [3-1:0] node1193;
	wire [3-1:0] node1194;
	wire [3-1:0] node1198;
	wire [3-1:0] node1199;
	wire [3-1:0] node1200;
	wire [3-1:0] node1204;
	wire [3-1:0] node1205;
	wire [3-1:0] node1208;
	wire [3-1:0] node1211;
	wire [3-1:0] node1212;
	wire [3-1:0] node1213;
	wire [3-1:0] node1214;
	wire [3-1:0] node1215;
	wire [3-1:0] node1218;
	wire [3-1:0] node1221;
	wire [3-1:0] node1222;
	wire [3-1:0] node1226;
	wire [3-1:0] node1227;
	wire [3-1:0] node1229;
	wire [3-1:0] node1232;
	wire [3-1:0] node1233;
	wire [3-1:0] node1236;
	wire [3-1:0] node1239;
	wire [3-1:0] node1240;
	wire [3-1:0] node1241;
	wire [3-1:0] node1243;
	wire [3-1:0] node1247;
	wire [3-1:0] node1248;
	wire [3-1:0] node1252;
	wire [3-1:0] node1253;
	wire [3-1:0] node1254;
	wire [3-1:0] node1255;
	wire [3-1:0] node1256;
	wire [3-1:0] node1258;
	wire [3-1:0] node1259;
	wire [3-1:0] node1263;
	wire [3-1:0] node1264;
	wire [3-1:0] node1267;
	wire [3-1:0] node1269;
	wire [3-1:0] node1272;
	wire [3-1:0] node1274;
	wire [3-1:0] node1276;
	wire [3-1:0] node1278;
	wire [3-1:0] node1281;
	wire [3-1:0] node1282;
	wire [3-1:0] node1283;
	wire [3-1:0] node1284;
	wire [3-1:0] node1288;
	wire [3-1:0] node1289;
	wire [3-1:0] node1290;
	wire [3-1:0] node1294;
	wire [3-1:0] node1295;
	wire [3-1:0] node1299;
	wire [3-1:0] node1300;
	wire [3-1:0] node1301;
	wire [3-1:0] node1305;
	wire [3-1:0] node1306;
	wire [3-1:0] node1308;
	wire [3-1:0] node1311;
	wire [3-1:0] node1315;
	wire [3-1:0] node1316;
	wire [3-1:0] node1317;
	wire [3-1:0] node1318;
	wire [3-1:0] node1319;
	wire [3-1:0] node1320;
	wire [3-1:0] node1321;
	wire [3-1:0] node1323;
	wire [3-1:0] node1327;
	wire [3-1:0] node1328;
	wire [3-1:0] node1329;
	wire [3-1:0] node1333;
	wire [3-1:0] node1336;
	wire [3-1:0] node1337;
	wire [3-1:0] node1338;
	wire [3-1:0] node1339;
	wire [3-1:0] node1343;
	wire [3-1:0] node1344;
	wire [3-1:0] node1349;
	wire [3-1:0] node1350;
	wire [3-1:0] node1351;
	wire [3-1:0] node1352;
	wire [3-1:0] node1355;
	wire [3-1:0] node1358;
	wire [3-1:0] node1359;
	wire [3-1:0] node1362;
	wire [3-1:0] node1363;
	wire [3-1:0] node1367;
	wire [3-1:0] node1368;
	wire [3-1:0] node1369;
	wire [3-1:0] node1371;
	wire [3-1:0] node1374;
	wire [3-1:0] node1375;
	wire [3-1:0] node1378;
	wire [3-1:0] node1381;
	wire [3-1:0] node1383;
	wire [3-1:0] node1386;
	wire [3-1:0] node1387;
	wire [3-1:0] node1388;
	wire [3-1:0] node1390;
	wire [3-1:0] node1391;
	wire [3-1:0] node1393;
	wire [3-1:0] node1397;
	wire [3-1:0] node1398;
	wire [3-1:0] node1399;
	wire [3-1:0] node1403;
	wire [3-1:0] node1404;
	wire [3-1:0] node1408;
	wire [3-1:0] node1409;
	wire [3-1:0] node1410;
	wire [3-1:0] node1412;
	wire [3-1:0] node1414;
	wire [3-1:0] node1417;
	wire [3-1:0] node1419;
	wire [3-1:0] node1420;
	wire [3-1:0] node1424;
	wire [3-1:0] node1425;
	wire [3-1:0] node1426;
	wire [3-1:0] node1430;
	wire [3-1:0] node1432;
	wire [3-1:0] node1435;
	wire [3-1:0] node1436;
	wire [3-1:0] node1437;
	wire [3-1:0] node1438;
	wire [3-1:0] node1439;
	wire [3-1:0] node1441;
	wire [3-1:0] node1442;
	wire [3-1:0] node1447;
	wire [3-1:0] node1448;
	wire [3-1:0] node1449;
	wire [3-1:0] node1451;
	wire [3-1:0] node1454;
	wire [3-1:0] node1458;
	wire [3-1:0] node1459;
	wire [3-1:0] node1460;
	wire [3-1:0] node1462;
	wire [3-1:0] node1464;
	wire [3-1:0] node1467;
	wire [3-1:0] node1468;
	wire [3-1:0] node1471;
	wire [3-1:0] node1473;
	wire [3-1:0] node1476;
	wire [3-1:0] node1477;
	wire [3-1:0] node1478;
	wire [3-1:0] node1480;
	wire [3-1:0] node1483;
	wire [3-1:0] node1484;
	wire [3-1:0] node1487;
	wire [3-1:0] node1491;
	wire [3-1:0] node1492;
	wire [3-1:0] node1493;
	wire [3-1:0] node1494;
	wire [3-1:0] node1495;
	wire [3-1:0] node1497;
	wire [3-1:0] node1501;
	wire [3-1:0] node1502;
	wire [3-1:0] node1503;
	wire [3-1:0] node1510;
	wire [3-1:0] node1511;
	wire [3-1:0] node1512;
	wire [3-1:0] node1513;
	wire [3-1:0] node1514;
	wire [3-1:0] node1516;
	wire [3-1:0] node1517;
	wire [3-1:0] node1518;
	wire [3-1:0] node1520;
	wire [3-1:0] node1522;
	wire [3-1:0] node1526;
	wire [3-1:0] node1527;
	wire [3-1:0] node1528;
	wire [3-1:0] node1529;
	wire [3-1:0] node1534;
	wire [3-1:0] node1537;
	wire [3-1:0] node1538;
	wire [3-1:0] node1539;
	wire [3-1:0] node1540;
	wire [3-1:0] node1542;
	wire [3-1:0] node1545;
	wire [3-1:0] node1546;
	wire [3-1:0] node1550;
	wire [3-1:0] node1551;
	wire [3-1:0] node1552;
	wire [3-1:0] node1554;
	wire [3-1:0] node1557;
	wire [3-1:0] node1559;
	wire [3-1:0] node1562;
	wire [3-1:0] node1563;
	wire [3-1:0] node1566;
	wire [3-1:0] node1568;
	wire [3-1:0] node1571;
	wire [3-1:0] node1572;
	wire [3-1:0] node1573;
	wire [3-1:0] node1575;
	wire [3-1:0] node1577;
	wire [3-1:0] node1580;
	wire [3-1:0] node1581;
	wire [3-1:0] node1582;
	wire [3-1:0] node1586;
	wire [3-1:0] node1588;
	wire [3-1:0] node1591;
	wire [3-1:0] node1592;
	wire [3-1:0] node1594;
	wire [3-1:0] node1597;
	wire [3-1:0] node1598;
	wire [3-1:0] node1602;
	wire [3-1:0] node1604;
	wire [3-1:0] node1606;
	wire [3-1:0] node1607;
	wire [3-1:0] node1608;
	wire [3-1:0] node1611;
	wire [3-1:0] node1612;
	wire [3-1:0] node1613;
	wire [3-1:0] node1617;
	wire [3-1:0] node1618;
	wire [3-1:0] node1622;
	wire [3-1:0] node1624;
	wire [3-1:0] node1626;
	wire [3-1:0] node1628;
	wire [3-1:0] node1631;
	wire [3-1:0] node1632;
	wire [3-1:0] node1633;
	wire [3-1:0] node1634;
	wire [3-1:0] node1635;
	wire [3-1:0] node1636;
	wire [3-1:0] node1637;
	wire [3-1:0] node1640;
	wire [3-1:0] node1643;
	wire [3-1:0] node1644;
	wire [3-1:0] node1647;
	wire [3-1:0] node1648;
	wire [3-1:0] node1651;
	wire [3-1:0] node1654;
	wire [3-1:0] node1655;
	wire [3-1:0] node1656;
	wire [3-1:0] node1659;
	wire [3-1:0] node1662;
	wire [3-1:0] node1663;
	wire [3-1:0] node1664;
	wire [3-1:0] node1668;
	wire [3-1:0] node1670;
	wire [3-1:0] node1673;
	wire [3-1:0] node1674;
	wire [3-1:0] node1675;
	wire [3-1:0] node1677;
	wire [3-1:0] node1680;
	wire [3-1:0] node1682;
	wire [3-1:0] node1683;
	wire [3-1:0] node1687;
	wire [3-1:0] node1688;
	wire [3-1:0] node1689;
	wire [3-1:0] node1690;
	wire [3-1:0] node1693;
	wire [3-1:0] node1696;
	wire [3-1:0] node1699;
	wire [3-1:0] node1700;
	wire [3-1:0] node1701;
	wire [3-1:0] node1704;
	wire [3-1:0] node1707;
	wire [3-1:0] node1708;
	wire [3-1:0] node1711;
	wire [3-1:0] node1714;
	wire [3-1:0] node1715;
	wire [3-1:0] node1716;
	wire [3-1:0] node1717;
	wire [3-1:0] node1718;
	wire [3-1:0] node1722;
	wire [3-1:0] node1723;
	wire [3-1:0] node1727;
	wire [3-1:0] node1728;
	wire [3-1:0] node1729;
	wire [3-1:0] node1732;
	wire [3-1:0] node1735;
	wire [3-1:0] node1736;
	wire [3-1:0] node1740;
	wire [3-1:0] node1741;
	wire [3-1:0] node1742;
	wire [3-1:0] node1744;
	wire [3-1:0] node1747;
	wire [3-1:0] node1748;
	wire [3-1:0] node1749;
	wire [3-1:0] node1752;
	wire [3-1:0] node1755;
	wire [3-1:0] node1756;
	wire [3-1:0] node1759;
	wire [3-1:0] node1762;
	wire [3-1:0] node1764;
	wire [3-1:0] node1767;
	wire [3-1:0] node1768;
	wire [3-1:0] node1769;
	wire [3-1:0] node1770;
	wire [3-1:0] node1771;
	wire [3-1:0] node1772;
	wire [3-1:0] node1775;
	wire [3-1:0] node1778;
	wire [3-1:0] node1779;
	wire [3-1:0] node1783;
	wire [3-1:0] node1784;
	wire [3-1:0] node1785;
	wire [3-1:0] node1786;
	wire [3-1:0] node1790;
	wire [3-1:0] node1793;
	wire [3-1:0] node1794;
	wire [3-1:0] node1797;
	wire [3-1:0] node1798;
	wire [3-1:0] node1802;
	wire [3-1:0] node1803;
	wire [3-1:0] node1804;
	wire [3-1:0] node1805;
	wire [3-1:0] node1807;
	wire [3-1:0] node1810;
	wire [3-1:0] node1813;
	wire [3-1:0] node1814;
	wire [3-1:0] node1815;
	wire [3-1:0] node1818;
	wire [3-1:0] node1821;
	wire [3-1:0] node1822;
	wire [3-1:0] node1825;
	wire [3-1:0] node1828;
	wire [3-1:0] node1830;
	wire [3-1:0] node1832;
	wire [3-1:0] node1835;
	wire [3-1:0] node1836;
	wire [3-1:0] node1837;
	wire [3-1:0] node1838;
	wire [3-1:0] node1839;
	wire [3-1:0] node1842;
	wire [3-1:0] node1843;
	wire [3-1:0] node1847;
	wire [3-1:0] node1849;
	wire [3-1:0] node1851;
	wire [3-1:0] node1854;
	wire [3-1:0] node1855;
	wire [3-1:0] node1857;
	wire [3-1:0] node1861;
	wire [3-1:0] node1862;
	wire [3-1:0] node1863;
	wire [3-1:0] node1864;
	wire [3-1:0] node1865;
	wire [3-1:0] node1869;
	wire [3-1:0] node1871;
	wire [3-1:0] node1876;
	wire [3-1:0] node1878;
	wire [3-1:0] node1879;
	wire [3-1:0] node1880;
	wire [3-1:0] node1881;
	wire [3-1:0] node1883;
	wire [3-1:0] node1885;
	wire [3-1:0] node1886;
	wire [3-1:0] node1888;
	wire [3-1:0] node1891;
	wire [3-1:0] node1892;
	wire [3-1:0] node1897;
	wire [3-1:0] node1898;
	wire [3-1:0] node1899;
	wire [3-1:0] node1900;
	wire [3-1:0] node1901;
	wire [3-1:0] node1902;
	wire [3-1:0] node1906;
	wire [3-1:0] node1909;
	wire [3-1:0] node1911;
	wire [3-1:0] node1914;
	wire [3-1:0] node1915;
	wire [3-1:0] node1916;
	wire [3-1:0] node1920;
	wire [3-1:0] node1921;
	wire [3-1:0] node1923;
	wire [3-1:0] node1926;
	wire [3-1:0] node1928;
	wire [3-1:0] node1931;
	wire [3-1:0] node1932;
	wire [3-1:0] node1933;
	wire [3-1:0] node1934;
	wire [3-1:0] node1935;
	wire [3-1:0] node1938;
	wire [3-1:0] node1942;
	wire [3-1:0] node1943;
	wire [3-1:0] node1947;
	wire [3-1:0] node1948;
	wire [3-1:0] node1949;
	wire [3-1:0] node1954;
	wire [3-1:0] node1955;
	wire [3-1:0] node1957;
	wire [3-1:0] node1958;
	wire [3-1:0] node1960;
	wire [3-1:0] node1962;

	assign outp = (inp[10]) ? node974 : node1;
		assign node1 = (inp[9]) ? node521 : node2;
			assign node2 = (inp[2]) ? node138 : node3;
				assign node3 = (inp[0]) ? 3'b110 : node4;
					assign node4 = (inp[3]) ? node80 : node5;
						assign node5 = (inp[5]) ? node47 : node6;
							assign node6 = (inp[11]) ? node34 : node7;
								assign node7 = (inp[6]) ? node17 : node8;
									assign node8 = (inp[7]) ? node14 : node9;
										assign node9 = (inp[8]) ? node11 : 3'b000;
											assign node11 = (inp[4]) ? 3'b000 : 3'b100;
										assign node14 = (inp[4]) ? 3'b100 : 3'b000;
									assign node17 = (inp[7]) ? node29 : node18;
										assign node18 = (inp[1]) ? node24 : node19;
											assign node19 = (inp[8]) ? 3'b111 : node20;
												assign node20 = (inp[4]) ? 3'b010 : 3'b111;
											assign node24 = (inp[8]) ? 3'b110 : node25;
												assign node25 = (inp[4]) ? 3'b010 : 3'b110;
										assign node29 = (inp[4]) ? node31 : 3'b010;
											assign node31 = (inp[8]) ? 3'b010 : 3'b110;
								assign node34 = (inp[7]) ? node42 : node35;
									assign node35 = (inp[4]) ? 3'b000 : node36;
										assign node36 = (inp[8]) ? node38 : 3'b000;
											assign node38 = (inp[1]) ? 3'b100 : 3'b111;
									assign node42 = (inp[4]) ? 3'b100 : node43;
										assign node43 = (inp[8]) ? 3'b000 : 3'b100;
							assign node47 = (inp[7]) ? node63 : node48;
								assign node48 = (inp[4]) ? node58 : node49;
									assign node49 = (inp[8]) ? node55 : node50;
										assign node50 = (inp[6]) ? node52 : 3'b010;
											assign node52 = (inp[11]) ? 3'b010 : 3'b000;
										assign node55 = (inp[1]) ? 3'b110 : 3'b111;
									assign node58 = (inp[11]) ? 3'b010 : node59;
										assign node59 = (inp[6]) ? 3'b000 : 3'b010;
								assign node63 = (inp[4]) ? node75 : node64;
									assign node64 = (inp[8]) ? node70 : node65;
										assign node65 = (inp[11]) ? 3'b110 : node66;
											assign node66 = (inp[6]) ? 3'b100 : 3'b110;
										assign node70 = (inp[11]) ? 3'b010 : node71;
											assign node71 = (inp[6]) ? 3'b000 : 3'b010;
									assign node75 = (inp[11]) ? 3'b110 : node76;
										assign node76 = (inp[6]) ? 3'b100 : 3'b110;
						assign node80 = (inp[1]) ? node82 : 3'b111;
							assign node82 = (inp[7]) ? node106 : node83;
								assign node83 = (inp[4]) ? node93 : node84;
									assign node84 = (inp[8]) ? 3'b111 : node85;
										assign node85 = (inp[5]) ? 3'b010 : node86;
											assign node86 = (inp[6]) ? node88 : 3'b000;
												assign node88 = (inp[11]) ? 3'b000 : 3'b111;
									assign node93 = (inp[5]) ? node101 : node94;
										assign node94 = (inp[11]) ? 3'b000 : node95;
											assign node95 = (inp[6]) ? node97 : 3'b000;
												assign node97 = (inp[8]) ? 3'b111 : 3'b010;
										assign node101 = (inp[11]) ? 3'b010 : node102;
											assign node102 = (inp[6]) ? 3'b000 : 3'b010;
								assign node106 = (inp[5]) ? node124 : node107;
									assign node107 = (inp[11]) ? node119 : node108;
										assign node108 = (inp[6]) ? node114 : node109;
											assign node109 = (inp[4]) ? 3'b100 : node110;
												assign node110 = (inp[8]) ? 3'b000 : 3'b100;
											assign node114 = (inp[8]) ? 3'b010 : node115;
												assign node115 = (inp[4]) ? 3'b110 : 3'b010;
										assign node119 = (inp[4]) ? 3'b100 : node120;
											assign node120 = (inp[8]) ? 3'b000 : 3'b100;
									assign node124 = (inp[4]) ? node132 : node125;
										assign node125 = (inp[8]) ? 3'b010 : node126;
											assign node126 = (inp[11]) ? 3'b110 : node127;
												assign node127 = (inp[6]) ? 3'b100 : 3'b110;
										assign node132 = (inp[6]) ? node134 : 3'b110;
											assign node134 = (inp[11]) ? 3'b110 : 3'b100;
				assign node138 = (inp[1]) ? node318 : node139;
					assign node139 = (inp[0]) ? node253 : node140;
						assign node140 = (inp[11]) ? node212 : node141;
							assign node141 = (inp[4]) ? node175 : node142;
								assign node142 = (inp[8]) ? node154 : node143;
									assign node143 = (inp[7]) ? 3'b000 : node144;
										assign node144 = (inp[3]) ? node146 : 3'b000;
											assign node146 = (inp[6]) ? node150 : node147;
												assign node147 = (inp[5]) ? 3'b010 : 3'b000;
												assign node150 = (inp[5]) ? 3'b000 : 3'b110;
									assign node154 = (inp[7]) ? node166 : node155;
										assign node155 = (inp[3]) ? node161 : node156;
											assign node156 = (inp[5]) ? 3'b000 : node157;
												assign node157 = (inp[6]) ? 3'b110 : 3'b100;
											assign node161 = (inp[6]) ? 3'b100 : node162;
												assign node162 = (inp[5]) ? 3'b110 : 3'b100;
										assign node166 = (inp[3]) ? node170 : node167;
											assign node167 = (inp[5]) ? 3'b000 : 3'b100;
											assign node170 = (inp[6]) ? node172 : 3'b000;
												assign node172 = (inp[5]) ? 3'b000 : 3'b010;
								assign node175 = (inp[5]) ? node199 : node176;
									assign node176 = (inp[8]) ? node190 : node177;
										assign node177 = (inp[6]) ? node185 : node178;
											assign node178 = (inp[3]) ? node182 : node179;
												assign node179 = (inp[7]) ? 3'b010 : 3'b100;
												assign node182 = (inp[7]) ? 3'b100 : 3'b000;
											assign node185 = (inp[3]) ? 3'b100 : node186;
												assign node186 = (inp[7]) ? 3'b000 : 3'b100;
										assign node190 = (inp[7]) ? node194 : node191;
											assign node191 = (inp[3]) ? 3'b110 : 3'b000;
											assign node194 = (inp[3]) ? 3'b000 : node195;
												assign node195 = (inp[6]) ? 3'b000 : 3'b010;
									assign node199 = (inp[7]) ? node205 : node200;
										assign node200 = (inp[3]) ? node202 : 3'b100;
											assign node202 = (inp[6]) ? 3'b000 : 3'b010;
										assign node205 = (inp[3]) ? 3'b100 : node206;
											assign node206 = (inp[6]) ? node208 : 3'b100;
												assign node208 = (inp[8]) ? 3'b010 : 3'b110;
							assign node212 = (inp[5]) ? node240 : node213;
								assign node213 = (inp[3]) ? node227 : node214;
									assign node214 = (inp[4]) ? node220 : node215;
										assign node215 = (inp[8]) ? node217 : 3'b010;
											assign node217 = (inp[7]) ? 3'b110 : 3'b100;
										assign node220 = (inp[7]) ? node224 : node221;
											assign node221 = (inp[8]) ? 3'b010 : 3'b110;
											assign node224 = (inp[8]) ? 3'b000 : 3'b100;
									assign node227 = (inp[7]) ? node233 : node228;
										assign node228 = (inp[8]) ? node230 : 3'b000;
											assign node230 = (inp[4]) ? 3'b000 : 3'b100;
										assign node233 = (inp[8]) ? node237 : node234;
											assign node234 = (inp[4]) ? 3'b110 : 3'b010;
											assign node237 = (inp[4]) ? 3'b010 : 3'b000;
								assign node240 = (inp[4]) ? node248 : node241;
									assign node241 = (inp[3]) ? node243 : 3'b010;
										assign node243 = (inp[8]) ? node245 : 3'b010;
											assign node245 = (inp[7]) ? 3'b010 : 3'b110;
									assign node248 = (inp[7]) ? 3'b110 : node249;
										assign node249 = (inp[3]) ? 3'b010 : 3'b110;
						assign node253 = (inp[3]) ? 3'b110 : node254;
							assign node254 = (inp[5]) ? node290 : node255;
								assign node255 = (inp[11]) ? node279 : node256;
									assign node256 = (inp[6]) ? node268 : node257;
										assign node257 = (inp[7]) ? node263 : node258;
											assign node258 = (inp[4]) ? 3'b000 : node259;
												assign node259 = (inp[8]) ? 3'b110 : 3'b000;
											assign node263 = (inp[8]) ? node265 : 3'b100;
												assign node265 = (inp[4]) ? 3'b100 : 3'b000;
										assign node268 = (inp[7]) ? node274 : node269;
											assign node269 = (inp[4]) ? node271 : 3'b110;
												assign node271 = (inp[8]) ? 3'b110 : 3'b010;
											assign node274 = (inp[4]) ? node276 : 3'b010;
												assign node276 = (inp[8]) ? 3'b010 : 3'b110;
									assign node279 = (inp[7]) ? node285 : node280;
										assign node280 = (inp[8]) ? node282 : 3'b000;
											assign node282 = (inp[4]) ? 3'b000 : 3'b110;
										assign node285 = (inp[4]) ? 3'b100 : node286;
											assign node286 = (inp[8]) ? 3'b000 : 3'b100;
								assign node290 = (inp[7]) ? node300 : node291;
									assign node291 = (inp[4]) ? node295 : node292;
										assign node292 = (inp[8]) ? 3'b110 : 3'b010;
										assign node295 = (inp[11]) ? 3'b010 : node296;
											assign node296 = (inp[6]) ? 3'b000 : 3'b010;
									assign node300 = (inp[11]) ? node312 : node301;
										assign node301 = (inp[6]) ? node307 : node302;
											assign node302 = (inp[4]) ? 3'b110 : node303;
												assign node303 = (inp[8]) ? 3'b010 : 3'b110;
											assign node307 = (inp[8]) ? node309 : 3'b100;
												assign node309 = (inp[4]) ? 3'b100 : 3'b000;
										assign node312 = (inp[8]) ? node314 : 3'b110;
											assign node314 = (inp[4]) ? 3'b110 : 3'b010;
					assign node318 = (inp[7]) ? node450 : node319;
						assign node319 = (inp[11]) ? node397 : node320;
							assign node320 = (inp[4]) ? node366 : node321;
								assign node321 = (inp[8]) ? node345 : node322;
									assign node322 = (inp[0]) ? node336 : node323;
										assign node323 = (inp[5]) ? node329 : node324;
											assign node324 = (inp[3]) ? node326 : 3'b010;
												assign node326 = (inp[6]) ? 3'b000 : 3'b010;
											assign node329 = (inp[6]) ? node333 : node330;
												assign node330 = (inp[3]) ? 3'b100 : 3'b110;
												assign node333 = (inp[3]) ? 3'b010 : 3'b110;
										assign node336 = (inp[3]) ? node338 : 3'b000;
											assign node338 = (inp[6]) ? node342 : node339;
												assign node339 = (inp[5]) ? 3'b010 : 3'b000;
												assign node342 = (inp[5]) ? 3'b000 : 3'b110;
									assign node345 = (inp[5]) ? node357 : node346;
										assign node346 = (inp[0]) ? node352 : node347;
											assign node347 = (inp[3]) ? 3'b100 : node348;
												assign node348 = (inp[6]) ? 3'b100 : 3'b110;
											assign node352 = (inp[6]) ? 3'b110 : node353;
												assign node353 = (inp[3]) ? 3'b110 : 3'b100;
										assign node357 = (inp[0]) ? node363 : node358;
											assign node358 = (inp[6]) ? 3'b010 : node359;
												assign node359 = (inp[3]) ? 3'b000 : 3'b010;
											assign node363 = (inp[3]) ? 3'b110 : 3'b000;
								assign node366 = (inp[3]) ? node384 : node367;
									assign node367 = (inp[6]) ? node373 : node368;
										assign node368 = (inp[8]) ? 3'b000 : node369;
											assign node369 = (inp[5]) ? 3'b000 : 3'b100;
										assign node373 = (inp[5]) ? node377 : node374;
											assign node374 = (inp[0]) ? 3'b000 : 3'b010;
											assign node377 = (inp[0]) ? node381 : node378;
												assign node378 = (inp[8]) ? 3'b000 : 3'b100;
												assign node381 = (inp[8]) ? 3'b100 : 3'b010;
									assign node384 = (inp[5]) ? node392 : node385;
										assign node385 = (inp[0]) ? node389 : node386;
											assign node386 = (inp[6]) ? 3'b100 : 3'b110;
											assign node389 = (inp[8]) ? 3'b000 : 3'b010;
										assign node392 = (inp[6]) ? node394 : 3'b010;
											assign node394 = (inp[0]) ? 3'b000 : 3'b010;
							assign node397 = (inp[5]) ? node433 : node398;
								assign node398 = (inp[8]) ? node410 : node399;
									assign node399 = (inp[0]) ? node405 : node400;
										assign node400 = (inp[4]) ? 3'b010 : node401;
											assign node401 = (inp[3]) ? 3'b000 : 3'b010;
										assign node405 = (inp[4]) ? 3'b000 : node406;
											assign node406 = (inp[3]) ? 3'b000 : 3'b010;
									assign node410 = (inp[3]) ? node426 : node411;
										assign node411 = (inp[6]) ? node419 : node412;
											assign node412 = (inp[4]) ? node416 : node413;
												assign node413 = (inp[0]) ? 3'b100 : 3'b010;
												assign node416 = (inp[0]) ? 3'b010 : 3'b100;
											assign node419 = (inp[0]) ? node423 : node420;
												assign node420 = (inp[4]) ? 3'b100 : 3'b010;
												assign node423 = (inp[4]) ? 3'b010 : 3'b100;
										assign node426 = (inp[4]) ? node430 : node427;
											assign node427 = (inp[0]) ? 3'b110 : 3'b000;
											assign node430 = (inp[0]) ? 3'b000 : 3'b010;
								assign node433 = (inp[4]) ? 3'b010 : node434;
									assign node434 = (inp[8]) ? node440 : node435;
										assign node435 = (inp[3]) ? node437 : 3'b010;
											assign node437 = (inp[0]) ? 3'b010 : 3'b110;
										assign node440 = (inp[6]) ? 3'b110 : node441;
											assign node441 = (inp[0]) ? node445 : node442;
												assign node442 = (inp[3]) ? 3'b010 : 3'b110;
												assign node445 = (inp[3]) ? 3'b110 : 3'b010;
						assign node450 = (inp[4]) ? node496 : node451;
							assign node451 = (inp[5]) ? node481 : node452;
								assign node452 = (inp[3]) ? node470 : node453;
									assign node453 = (inp[0]) ? node465 : node454;
										assign node454 = (inp[6]) ? node460 : node455;
											assign node455 = (inp[8]) ? 3'b000 : node456;
												assign node456 = (inp[11]) ? 3'b010 : 3'b000;
											assign node460 = (inp[8]) ? node462 : 3'b010;
												assign node462 = (inp[11]) ? 3'b000 : 3'b010;
										assign node465 = (inp[8]) ? 3'b010 : node466;
											assign node466 = (inp[11]) ? 3'b000 : 3'b010;
									assign node470 = (inp[0]) ? node472 : 3'b000;
										assign node472 = (inp[11]) ? node478 : node473;
											assign node473 = (inp[6]) ? node475 : 3'b000;
												assign node475 = (inp[8]) ? 3'b010 : 3'b000;
											assign node478 = (inp[8]) ? 3'b000 : 3'b010;
								assign node481 = (inp[11]) ? 3'b010 : node482;
									assign node482 = (inp[0]) ? node488 : node483;
										assign node483 = (inp[8]) ? 3'b010 : node484;
											assign node484 = (inp[6]) ? 3'b000 : 3'b010;
										assign node488 = (inp[6]) ? 3'b000 : node489;
											assign node489 = (inp[8]) ? node491 : 3'b000;
												assign node491 = (inp[3]) ? 3'b000 : 3'b010;
							assign node496 = (inp[11]) ? 3'b000 : node497;
								assign node497 = (inp[5]) ? 3'b000 : node498;
									assign node498 = (inp[6]) ? node512 : node499;
										assign node499 = (inp[8]) ? node505 : node500;
											assign node500 = (inp[0]) ? 3'b000 : node501;
												assign node501 = (inp[3]) ? 3'b010 : 3'b000;
											assign node505 = (inp[3]) ? node509 : node506;
												assign node506 = (inp[0]) ? 3'b000 : 3'b010;
												assign node509 = (inp[0]) ? 3'b010 : 3'b000;
										assign node512 = (inp[0]) ? node514 : 3'b000;
											assign node514 = (inp[8]) ? node516 : 3'b000;
												assign node516 = (inp[3]) ? 3'b000 : 3'b010;
			assign node521 = (inp[2]) ? node643 : node522;
				assign node522 = (inp[0]) ? 3'b010 : node523;
					assign node523 = (inp[3]) ? node611 : node524;
						assign node524 = (inp[1]) ? node550 : node525;
							assign node525 = (inp[7]) ? node527 : 3'b011;
								assign node527 = (inp[4]) ? node537 : node528;
									assign node528 = (inp[8]) ? 3'b011 : node529;
										assign node529 = (inp[11]) ? node533 : node530;
											assign node530 = (inp[5]) ? 3'b010 : 3'b011;
											assign node533 = (inp[5]) ? 3'b010 : 3'b000;
									assign node537 = (inp[5]) ? node545 : node538;
										assign node538 = (inp[6]) ? node540 : 3'b000;
											assign node540 = (inp[11]) ? 3'b000 : node541;
												assign node541 = (inp[8]) ? 3'b011 : 3'b010;
										assign node545 = (inp[11]) ? 3'b010 : node546;
											assign node546 = (inp[6]) ? 3'b000 : 3'b010;
							assign node550 = (inp[5]) ? node582 : node551;
								assign node551 = (inp[6]) ? node563 : node552;
									assign node552 = (inp[7]) ? node558 : node553;
										assign node553 = (inp[4]) ? 3'b100 : node554;
											assign node554 = (inp[8]) ? 3'b000 : 3'b100;
										assign node558 = (inp[4]) ? 3'b000 : node559;
											assign node559 = (inp[11]) ? 3'b000 : 3'b100;
									assign node563 = (inp[11]) ? node573 : node564;
										assign node564 = (inp[7]) ? node570 : node565;
											assign node565 = (inp[8]) ? 3'b010 : node566;
												assign node566 = (inp[4]) ? 3'b110 : 3'b010;
											assign node570 = (inp[4]) ? 3'b010 : 3'b110;
										assign node573 = (inp[4]) ? 3'b000 : node574;
											assign node574 = (inp[7]) ? node578 : node575;
												assign node575 = (inp[8]) ? 3'b000 : 3'b100;
												assign node578 = (inp[8]) ? 3'b100 : 3'b000;
								assign node582 = (inp[7]) ? node598 : node583;
									assign node583 = (inp[6]) ? node589 : node584;
										assign node584 = (inp[8]) ? node586 : 3'b110;
											assign node586 = (inp[4]) ? 3'b110 : 3'b010;
										assign node589 = (inp[11]) ? node595 : node590;
											assign node590 = (inp[8]) ? node592 : 3'b100;
												assign node592 = (inp[4]) ? 3'b100 : 3'b000;
											assign node595 = (inp[4]) ? 3'b110 : 3'b010;
									assign node598 = (inp[4]) ? node606 : node599;
										assign node599 = (inp[8]) ? node601 : 3'b010;
											assign node601 = (inp[11]) ? 3'b110 : node602;
												assign node602 = (inp[6]) ? 3'b100 : 3'b110;
										assign node606 = (inp[11]) ? 3'b010 : node607;
											assign node607 = (inp[6]) ? 3'b000 : 3'b010;
						assign node611 = (inp[7]) ? node613 : 3'b011;
							assign node613 = (inp[1]) ? node615 : 3'b011;
								assign node615 = (inp[4]) ? node629 : node616;
									assign node616 = (inp[8]) ? 3'b011 : node617;
										assign node617 = (inp[5]) ? node623 : node618;
											assign node618 = (inp[11]) ? 3'b000 : node619;
												assign node619 = (inp[6]) ? 3'b011 : 3'b000;
											assign node623 = (inp[6]) ? node625 : 3'b010;
												assign node625 = (inp[11]) ? 3'b010 : 3'b000;
									assign node629 = (inp[5]) ? node637 : node630;
										assign node630 = (inp[6]) ? node632 : 3'b000;
											assign node632 = (inp[11]) ? 3'b000 : node633;
												assign node633 = (inp[8]) ? 3'b011 : 3'b010;
										assign node637 = (inp[6]) ? node639 : 3'b010;
											assign node639 = (inp[11]) ? 3'b010 : 3'b000;
				assign node643 = (inp[0]) ? node873 : node644;
					assign node644 = (inp[1]) ? node750 : node645;
						assign node645 = (inp[11]) ? node709 : node646;
							assign node646 = (inp[4]) ? node682 : node647;
								assign node647 = (inp[7]) ? node661 : node648;
									assign node648 = (inp[8]) ? node656 : node649;
										assign node649 = (inp[6]) ? node653 : node650;
											assign node650 = (inp[5]) ? 3'b110 : 3'b100;
											assign node653 = (inp[5]) ? 3'b100 : 3'b010;
										assign node656 = (inp[6]) ? node658 : 3'b010;
											assign node658 = (inp[3]) ? 3'b000 : 3'b010;
									assign node661 = (inp[3]) ? node667 : node662;
										assign node662 = (inp[8]) ? node664 : 3'b100;
											assign node664 = (inp[5]) ? 3'b100 : 3'b000;
										assign node667 = (inp[8]) ? node675 : node668;
											assign node668 = (inp[5]) ? node672 : node669;
												assign node669 = (inp[6]) ? 3'b110 : 3'b000;
												assign node672 = (inp[6]) ? 3'b000 : 3'b010;
											assign node675 = (inp[5]) ? node679 : node676;
												assign node676 = (inp[6]) ? 3'b110 : 3'b100;
												assign node679 = (inp[6]) ? 3'b100 : 3'b110;
								assign node682 = (inp[3]) ? node692 : node683;
									assign node683 = (inp[5]) ? 3'b000 : node684;
										assign node684 = (inp[8]) ? node686 : 3'b000;
											assign node686 = (inp[6]) ? node688 : 3'b100;
												assign node688 = (inp[7]) ? 3'b100 : 3'b010;
									assign node692 = (inp[7]) ? node702 : node693;
										assign node693 = (inp[5]) ? node699 : node694;
											assign node694 = (inp[6]) ? node696 : 3'b100;
												assign node696 = (inp[8]) ? 3'b010 : 3'b110;
											assign node699 = (inp[6]) ? 3'b100 : 3'b110;
										assign node702 = (inp[6]) ? node704 : 3'b000;
											assign node704 = (inp[5]) ? 3'b000 : node705;
												assign node705 = (inp[8]) ? 3'b110 : 3'b000;
							assign node709 = (inp[5]) ? node735 : node710;
								assign node710 = (inp[7]) ? node720 : node711;
									assign node711 = (inp[4]) ? node715 : node712;
										assign node712 = (inp[8]) ? 3'b000 : 3'b100;
										assign node715 = (inp[8]) ? 3'b100 : node716;
											assign node716 = (inp[3]) ? 3'b100 : 3'b010;
									assign node720 = (inp[3]) ? node728 : node721;
										assign node721 = (inp[8]) ? node725 : node722;
											assign node722 = (inp[4]) ? 3'b000 : 3'b110;
											assign node725 = (inp[4]) ? 3'b110 : 3'b010;
										assign node728 = (inp[8]) ? node732 : node729;
											assign node729 = (inp[4]) ? 3'b010 : 3'b000;
											assign node732 = (inp[4]) ? 3'b000 : 3'b100;
								assign node735 = (inp[4]) ? node745 : node736;
									assign node736 = (inp[7]) ? node740 : node737;
										assign node737 = (inp[8]) ? 3'b010 : 3'b110;
										assign node740 = (inp[8]) ? 3'b110 : node741;
											assign node741 = (inp[3]) ? 3'b010 : 3'b110;
									assign node745 = (inp[7]) ? 3'b010 : node746;
										assign node746 = (inp[3]) ? 3'b110 : 3'b010;
						assign node750 = (inp[7]) ? node824 : node751;
							assign node751 = (inp[5]) ? node795 : node752;
								assign node752 = (inp[8]) ? node776 : node753;
									assign node753 = (inp[4]) ? node767 : node754;
										assign node754 = (inp[6]) ? node762 : node755;
											assign node755 = (inp[11]) ? node759 : node756;
												assign node756 = (inp[3]) ? 3'b100 : 3'b110;
												assign node759 = (inp[3]) ? 3'b110 : 3'b100;
											assign node762 = (inp[3]) ? node764 : 3'b100;
												assign node764 = (inp[11]) ? 3'b110 : 3'b100;
										assign node767 = (inp[11]) ? node773 : node768;
											assign node768 = (inp[6]) ? 3'b110 : node769;
												assign node769 = (inp[3]) ? 3'b010 : 3'b000;
											assign node773 = (inp[3]) ? 3'b100 : 3'b000;
									assign node776 = (inp[6]) ? node786 : node777;
										assign node777 = (inp[11]) ? node783 : node778;
											assign node778 = (inp[3]) ? node780 : 3'b010;
												assign node780 = (inp[4]) ? 3'b010 : 3'b000;
											assign node783 = (inp[4]) ? 3'b000 : 3'b010;
										assign node786 = (inp[3]) ? node790 : node787;
											assign node787 = (inp[11]) ? 3'b100 : 3'b000;
											assign node790 = (inp[4]) ? 3'b000 : node791;
												assign node791 = (inp[11]) ? 3'b010 : 3'b000;
								assign node795 = (inp[11]) ? node817 : node796;
									assign node796 = (inp[4]) ? node808 : node797;
										assign node797 = (inp[3]) ? node803 : node798;
											assign node798 = (inp[6]) ? node800 : 3'b100;
												assign node800 = (inp[8]) ? 3'b110 : 3'b010;
											assign node803 = (inp[6]) ? 3'b100 : node804;
												assign node804 = (inp[8]) ? 3'b100 : 3'b000;
										assign node808 = (inp[6]) ? node814 : node809;
											assign node809 = (inp[3]) ? 3'b100 : node810;
												assign node810 = (inp[8]) ? 3'b010 : 3'b000;
											assign node814 = (inp[3]) ? 3'b010 : 3'b000;
									assign node817 = (inp[8]) ? node819 : 3'b010;
										assign node819 = (inp[3]) ? node821 : 3'b010;
											assign node821 = (inp[4]) ? 3'b010 : 3'b110;
							assign node824 = (inp[4]) ? node858 : node825;
								assign node825 = (inp[11]) ? node841 : node826;
									assign node826 = (inp[5]) ? node834 : node827;
										assign node827 = (inp[3]) ? node831 : node828;
											assign node828 = (inp[6]) ? 3'b000 : 3'b010;
											assign node831 = (inp[6]) ? 3'b010 : 3'b000;
										assign node834 = (inp[6]) ? node836 : 3'b000;
											assign node836 = (inp[3]) ? node838 : 3'b000;
												assign node838 = (inp[8]) ? 3'b000 : 3'b010;
									assign node841 = (inp[5]) ? 3'b010 : node842;
										assign node842 = (inp[6]) ? node850 : node843;
											assign node843 = (inp[3]) ? node847 : node844;
												assign node844 = (inp[8]) ? 3'b010 : 3'b000;
												assign node847 = (inp[8]) ? 3'b000 : 3'b010;
											assign node850 = (inp[3]) ? node854 : node851;
												assign node851 = (inp[8]) ? 3'b010 : 3'b000;
												assign node854 = (inp[8]) ? 3'b000 : 3'b010;
								assign node858 = (inp[5]) ? 3'b000 : node859;
									assign node859 = (inp[11]) ? 3'b000 : node860;
										assign node860 = (inp[6]) ? node866 : node861;
											assign node861 = (inp[3]) ? node863 : 3'b000;
												assign node863 = (inp[8]) ? 3'b010 : 3'b000;
											assign node866 = (inp[8]) ? node868 : 3'b010;
												assign node868 = (inp[3]) ? 3'b000 : 3'b010;
					assign node873 = (inp[1]) ? node897 : node874;
						assign node874 = (inp[3]) ? 3'b010 : node875;
							assign node875 = (inp[7]) ? node877 : 3'b010;
								assign node877 = (inp[5]) ? node887 : node878;
									assign node878 = (inp[6]) ? node880 : 3'b000;
										assign node880 = (inp[11]) ? node882 : 3'b010;
											assign node882 = (inp[4]) ? 3'b000 : node883;
												assign node883 = (inp[8]) ? 3'b010 : 3'b000;
									assign node887 = (inp[11]) ? 3'b010 : node888;
										assign node888 = (inp[8]) ? node890 : 3'b000;
											assign node890 = (inp[6]) ? node892 : 3'b010;
												assign node892 = (inp[4]) ? 3'b000 : 3'b010;
						assign node897 = (inp[7]) ? node937 : node898;
							assign node898 = (inp[3]) ? 3'b010 : node899;
								assign node899 = (inp[11]) ? node923 : node900;
									assign node900 = (inp[4]) ? node916 : node901;
										assign node901 = (inp[8]) ? node909 : node902;
											assign node902 = (inp[5]) ? node906 : node903;
												assign node903 = (inp[6]) ? 3'b010 : 3'b100;
												assign node906 = (inp[6]) ? 3'b100 : 3'b110;
											assign node909 = (inp[6]) ? node913 : node910;
												assign node910 = (inp[5]) ? 3'b010 : 3'b000;
												assign node913 = (inp[5]) ? 3'b000 : 3'b010;
										assign node916 = (inp[5]) ? 3'b000 : node917;
											assign node917 = (inp[8]) ? node919 : 3'b000;
												assign node919 = (inp[6]) ? 3'b010 : 3'b100;
									assign node923 = (inp[5]) ? node931 : node924;
										assign node924 = (inp[8]) ? node928 : node925;
											assign node925 = (inp[4]) ? 3'b010 : 3'b100;
											assign node928 = (inp[4]) ? 3'b100 : 3'b000;
										assign node931 = (inp[8]) ? 3'b010 : node932;
											assign node932 = (inp[4]) ? 3'b010 : 3'b110;
							assign node937 = (inp[4]) ? node961 : node938;
								assign node938 = (inp[5]) ? node952 : node939;
									assign node939 = (inp[3]) ? node945 : node940;
										assign node940 = (inp[8]) ? 3'b000 : node941;
											assign node941 = (inp[6]) ? 3'b000 : 3'b010;
										assign node945 = (inp[8]) ? 3'b010 : node946;
											assign node946 = (inp[11]) ? 3'b000 : node947;
												assign node947 = (inp[6]) ? 3'b010 : 3'b000;
									assign node952 = (inp[6]) ? 3'b010 : node953;
										assign node953 = (inp[8]) ? node955 : 3'b010;
											assign node955 = (inp[3]) ? 3'b010 : node956;
												assign node956 = (inp[11]) ? 3'b010 : 3'b000;
								assign node961 = (inp[5]) ? 3'b000 : node962;
									assign node962 = (inp[11]) ? 3'b000 : node963;
										assign node963 = (inp[6]) ? node967 : node964;
											assign node964 = (inp[8]) ? 3'b000 : 3'b010;
											assign node967 = (inp[8]) ? node969 : 3'b000;
												assign node969 = (inp[3]) ? 3'b010 : 3'b000;
		assign node974 = (inp[9]) ? node1510 : node975;
			assign node975 = (inp[2]) ? node1129 : node976;
				assign node976 = (inp[0]) ? 3'b100 : node977;
					assign node977 = (inp[3]) ? node1065 : node978;
						assign node978 = (inp[5]) ? node1022 : node979;
							assign node979 = (inp[7]) ? node1005 : node980;
								assign node980 = (inp[1]) ? node990 : node981;
									assign node981 = (inp[4]) ? node983 : 3'b101;
										assign node983 = (inp[8]) ? 3'b101 : node984;
											assign node984 = (inp[11]) ? 3'b010 : node985;
												assign node985 = (inp[6]) ? 3'b000 : 3'b010;
									assign node990 = (inp[4]) ? node996 : node991;
										assign node991 = (inp[11]) ? 3'b110 : node992;
											assign node992 = (inp[6]) ? 3'b100 : 3'b110;
										assign node996 = (inp[8]) ? node1002 : node997;
											assign node997 = (inp[11]) ? 3'b010 : node998;
												assign node998 = (inp[6]) ? 3'b000 : 3'b010;
											assign node1002 = (inp[11]) ? 3'b110 : 3'b100;
								assign node1005 = (inp[8]) ? node1017 : node1006;
									assign node1006 = (inp[4]) ? node1012 : node1007;
										assign node1007 = (inp[6]) ? node1009 : 3'b010;
											assign node1009 = (inp[11]) ? 3'b010 : 3'b000;
										assign node1012 = (inp[11]) ? 3'b110 : node1013;
											assign node1013 = (inp[6]) ? 3'b100 : 3'b110;
									assign node1017 = (inp[11]) ? 3'b010 : node1018;
										assign node1018 = (inp[6]) ? 3'b000 : 3'b010;
							assign node1022 = (inp[11]) ? node1052 : node1023;
								assign node1023 = (inp[6]) ? node1035 : node1024;
									assign node1024 = (inp[7]) ? node1030 : node1025;
										assign node1025 = (inp[4]) ? 3'b000 : node1026;
											assign node1026 = (inp[8]) ? 3'b101 : 3'b000;
										assign node1030 = (inp[8]) ? node1032 : 3'b100;
											assign node1032 = (inp[4]) ? 3'b100 : 3'b000;
									assign node1035 = (inp[7]) ? node1047 : node1036;
										assign node1036 = (inp[1]) ? node1042 : node1037;
											assign node1037 = (inp[4]) ? node1039 : 3'b101;
												assign node1039 = (inp[8]) ? 3'b101 : 3'b010;
											assign node1042 = (inp[8]) ? 3'b110 : node1043;
												assign node1043 = (inp[4]) ? 3'b010 : 3'b110;
										assign node1047 = (inp[4]) ? node1049 : 3'b010;
											assign node1049 = (inp[8]) ? 3'b010 : 3'b110;
								assign node1052 = (inp[7]) ? node1060 : node1053;
									assign node1053 = (inp[8]) ? node1055 : 3'b000;
										assign node1055 = (inp[4]) ? 3'b000 : node1056;
											assign node1056 = (inp[1]) ? 3'b100 : 3'b101;
									assign node1060 = (inp[4]) ? 3'b100 : node1061;
										assign node1061 = (inp[8]) ? 3'b000 : 3'b100;
						assign node1065 = (inp[1]) ? node1067 : 3'b101;
							assign node1067 = (inp[7]) ? node1095 : node1068;
								assign node1068 = (inp[4]) ? node1078 : node1069;
									assign node1069 = (inp[8]) ? 3'b101 : node1070;
										assign node1070 = (inp[5]) ? node1072 : 3'b101;
											assign node1072 = (inp[6]) ? node1074 : 3'b000;
												assign node1074 = (inp[11]) ? 3'b000 : 3'b101;
									assign node1078 = (inp[8]) ? node1088 : node1079;
										assign node1079 = (inp[5]) ? node1085 : node1080;
											assign node1080 = (inp[6]) ? node1082 : 3'b010;
												assign node1082 = (inp[11]) ? 3'b010 : 3'b000;
											assign node1085 = (inp[11]) ? 3'b000 : 3'b010;
										assign node1088 = (inp[5]) ? node1090 : 3'b101;
											assign node1090 = (inp[11]) ? 3'b000 : node1091;
												assign node1091 = (inp[6]) ? 3'b101 : 3'b000;
								assign node1095 = (inp[4]) ? node1113 : node1096;
									assign node1096 = (inp[5]) ? node1102 : node1097;
										assign node1097 = (inp[6]) ? node1099 : 3'b010;
											assign node1099 = (inp[11]) ? 3'b010 : 3'b000;
										assign node1102 = (inp[8]) ? node1108 : node1103;
											assign node1103 = (inp[11]) ? 3'b100 : node1104;
												assign node1104 = (inp[6]) ? 3'b010 : 3'b100;
											assign node1108 = (inp[11]) ? 3'b000 : node1109;
												assign node1109 = (inp[6]) ? 3'b010 : 3'b000;
									assign node1113 = (inp[6]) ? node1117 : node1114;
										assign node1114 = (inp[5]) ? 3'b100 : 3'b110;
										assign node1117 = (inp[8]) ? node1123 : node1118;
											assign node1118 = (inp[11]) ? 3'b110 : node1119;
												assign node1119 = (inp[5]) ? 3'b110 : 3'b100;
											assign node1123 = (inp[5]) ? node1125 : 3'b010;
												assign node1125 = (inp[11]) ? 3'b100 : 3'b010;
				assign node1129 = (inp[1]) ? node1315 : node1130;
					assign node1130 = (inp[0]) ? node1252 : node1131;
						assign node1131 = (inp[11]) ? node1211 : node1132;
							assign node1132 = (inp[4]) ? node1168 : node1133;
								assign node1133 = (inp[7]) ? node1151 : node1134;
									assign node1134 = (inp[8]) ? node1144 : node1135;
										assign node1135 = (inp[5]) ? node1139 : node1136;
											assign node1136 = (inp[6]) ? 3'b100 : 3'b110;
											assign node1139 = (inp[6]) ? node1141 : 3'b000;
												assign node1141 = (inp[3]) ? 3'b110 : 3'b010;
										assign node1144 = (inp[5]) ? node1148 : node1145;
											assign node1145 = (inp[6]) ? 3'b100 : 3'b110;
											assign node1148 = (inp[6]) ? 3'b110 : 3'b100;
									assign node1151 = (inp[3]) ? node1155 : node1152;
										assign node1152 = (inp[5]) ? 3'b010 : 3'b110;
										assign node1155 = (inp[8]) ? node1161 : node1156;
											assign node1156 = (inp[6]) ? node1158 : 3'b010;
												assign node1158 = (inp[5]) ? 3'b010 : 3'b000;
											assign node1161 = (inp[6]) ? node1165 : node1162;
												assign node1162 = (inp[5]) ? 3'b000 : 3'b010;
												assign node1165 = (inp[5]) ? 3'b010 : 3'b000;
								assign node1168 = (inp[5]) ? node1188 : node1169;
									assign node1169 = (inp[8]) ? node1181 : node1170;
										assign node1170 = (inp[3]) ? node1176 : node1171;
											assign node1171 = (inp[6]) ? 3'b010 : node1172;
												assign node1172 = (inp[7]) ? 3'b000 : 3'b010;
											assign node1176 = (inp[7]) ? 3'b010 : node1177;
												assign node1177 = (inp[6]) ? 3'b000 : 3'b010;
										assign node1181 = (inp[3]) ? node1183 : 3'b010;
											assign node1183 = (inp[7]) ? 3'b010 : node1184;
												assign node1184 = (inp[6]) ? 3'b100 : 3'b110;
									assign node1188 = (inp[8]) ? node1198 : node1189;
										assign node1189 = (inp[7]) ? node1193 : node1190;
											assign node1190 = (inp[6]) ? 3'b110 : 3'b000;
											assign node1193 = (inp[3]) ? 3'b110 : node1194;
												assign node1194 = (inp[6]) ? 3'b100 : 3'b110;
										assign node1198 = (inp[6]) ? node1204 : node1199;
											assign node1199 = (inp[7]) ? 3'b010 : node1200;
												assign node1200 = (inp[3]) ? 3'b000 : 3'b010;
											assign node1204 = (inp[3]) ? node1208 : node1205;
												assign node1205 = (inp[7]) ? 3'b000 : 3'b010;
												assign node1208 = (inp[7]) ? 3'b010 : 3'b110;
							assign node1211 = (inp[5]) ? node1239 : node1212;
								assign node1212 = (inp[7]) ? node1226 : node1213;
									assign node1213 = (inp[3]) ? node1221 : node1214;
										assign node1214 = (inp[8]) ? node1218 : node1215;
											assign node1215 = (inp[4]) ? 3'b100 : 3'b000;
											assign node1218 = (inp[4]) ? 3'b000 : 3'b110;
										assign node1221 = (inp[8]) ? 3'b110 : node1222;
											assign node1222 = (inp[4]) ? 3'b010 : 3'b110;
									assign node1226 = (inp[8]) ? node1232 : node1227;
										assign node1227 = (inp[4]) ? node1229 : 3'b000;
											assign node1229 = (inp[3]) ? 3'b100 : 3'b010;
										assign node1232 = (inp[4]) ? node1236 : node1233;
											assign node1233 = (inp[3]) ? 3'b010 : 3'b100;
											assign node1236 = (inp[3]) ? 3'b000 : 3'b010;
								assign node1239 = (inp[4]) ? node1247 : node1240;
									assign node1240 = (inp[7]) ? 3'b000 : node1241;
										assign node1241 = (inp[3]) ? node1243 : 3'b000;
											assign node1243 = (inp[8]) ? 3'b100 : 3'b000;
									assign node1247 = (inp[7]) ? 3'b100 : node1248;
										assign node1248 = (inp[3]) ? 3'b000 : 3'b100;
						assign node1252 = (inp[3]) ? 3'b100 : node1253;
							assign node1253 = (inp[7]) ? node1281 : node1254;
								assign node1254 = (inp[8]) ? node1272 : node1255;
									assign node1255 = (inp[4]) ? node1263 : node1256;
										assign node1256 = (inp[5]) ? node1258 : 3'b100;
											assign node1258 = (inp[11]) ? 3'b000 : node1259;
												assign node1259 = (inp[6]) ? 3'b100 : 3'b000;
										assign node1263 = (inp[5]) ? node1267 : node1264;
											assign node1264 = (inp[6]) ? 3'b000 : 3'b010;
											assign node1267 = (inp[6]) ? node1269 : 3'b000;
												assign node1269 = (inp[11]) ? 3'b000 : 3'b010;
									assign node1272 = (inp[4]) ? node1274 : 3'b100;
										assign node1274 = (inp[5]) ? node1276 : 3'b100;
											assign node1276 = (inp[6]) ? node1278 : 3'b000;
												assign node1278 = (inp[11]) ? 3'b000 : 3'b100;
								assign node1281 = (inp[5]) ? node1299 : node1282;
									assign node1282 = (inp[6]) ? node1288 : node1283;
										assign node1283 = (inp[8]) ? 3'b010 : node1284;
											assign node1284 = (inp[4]) ? 3'b110 : 3'b010;
										assign node1288 = (inp[11]) ? node1294 : node1289;
											assign node1289 = (inp[8]) ? 3'b000 : node1290;
												assign node1290 = (inp[4]) ? 3'b100 : 3'b000;
											assign node1294 = (inp[8]) ? 3'b010 : node1295;
												assign node1295 = (inp[4]) ? 3'b110 : 3'b010;
									assign node1299 = (inp[6]) ? node1305 : node1300;
										assign node1300 = (inp[4]) ? 3'b100 : node1301;
											assign node1301 = (inp[8]) ? 3'b000 : 3'b100;
										assign node1305 = (inp[11]) ? node1311 : node1306;
											assign node1306 = (inp[4]) ? node1308 : 3'b010;
												assign node1308 = (inp[8]) ? 3'b010 : 3'b110;
											assign node1311 = (inp[8]) ? 3'b000 : 3'b100;
					assign node1315 = (inp[7]) ? node1435 : node1316;
						assign node1316 = (inp[4]) ? node1386 : node1317;
							assign node1317 = (inp[5]) ? node1349 : node1318;
								assign node1318 = (inp[0]) ? node1336 : node1319;
									assign node1319 = (inp[3]) ? node1327 : node1320;
										assign node1320 = (inp[11]) ? 3'b000 : node1321;
											assign node1321 = (inp[8]) ? node1323 : 3'b000;
												assign node1323 = (inp[6]) ? 3'b110 : 3'b100;
										assign node1327 = (inp[8]) ? node1333 : node1328;
											assign node1328 = (inp[6]) ? 3'b110 : node1329;
												assign node1329 = (inp[11]) ? 3'b010 : 3'b000;
											assign node1333 = (inp[11]) ? 3'b100 : 3'b110;
									assign node1336 = (inp[3]) ? 3'b100 : node1337;
										assign node1337 = (inp[8]) ? node1343 : node1338;
											assign node1338 = (inp[11]) ? 3'b000 : node1339;
												assign node1339 = (inp[6]) ? 3'b100 : 3'b110;
											assign node1343 = (inp[11]) ? 3'b110 : node1344;
												assign node1344 = (inp[6]) ? 3'b100 : 3'b110;
								assign node1349 = (inp[11]) ? node1367 : node1350;
									assign node1350 = (inp[0]) ? node1358 : node1351;
										assign node1351 = (inp[3]) ? node1355 : node1352;
											assign node1352 = (inp[8]) ? 3'b000 : 3'b100;
											assign node1355 = (inp[6]) ? 3'b000 : 3'b010;
										assign node1358 = (inp[3]) ? node1362 : node1359;
											assign node1359 = (inp[8]) ? 3'b110 : 3'b010;
											assign node1362 = (inp[6]) ? 3'b100 : node1363;
												assign node1363 = (inp[8]) ? 3'b100 : 3'b000;
									assign node1367 = (inp[0]) ? node1381 : node1368;
										assign node1368 = (inp[6]) ? node1374 : node1369;
											assign node1369 = (inp[8]) ? node1371 : 3'b100;
												assign node1371 = (inp[3]) ? 3'b000 : 3'b100;
											assign node1374 = (inp[8]) ? node1378 : node1375;
												assign node1375 = (inp[3]) ? 3'b100 : 3'b000;
												assign node1378 = (inp[3]) ? 3'b000 : 3'b100;
										assign node1381 = (inp[8]) ? node1383 : 3'b000;
											assign node1383 = (inp[3]) ? 3'b100 : 3'b000;
							assign node1386 = (inp[3]) ? node1408 : node1387;
								assign node1387 = (inp[11]) ? node1397 : node1388;
									assign node1388 = (inp[6]) ? node1390 : 3'b010;
										assign node1390 = (inp[8]) ? 3'b010 : node1391;
											assign node1391 = (inp[0]) ? node1393 : 3'b000;
												assign node1393 = (inp[5]) ? 3'b000 : 3'b010;
									assign node1397 = (inp[8]) ? node1403 : node1398;
										assign node1398 = (inp[5]) ? 3'b000 : node1399;
											assign node1399 = (inp[0]) ? 3'b100 : 3'b000;
										assign node1403 = (inp[0]) ? 3'b000 : node1404;
											assign node1404 = (inp[5]) ? 3'b000 : 3'b010;
								assign node1408 = (inp[8]) ? node1424 : node1409;
									assign node1409 = (inp[0]) ? node1417 : node1410;
										assign node1410 = (inp[5]) ? node1412 : 3'b000;
											assign node1412 = (inp[6]) ? node1414 : 3'b000;
												assign node1414 = (inp[11]) ? 3'b000 : 3'b100;
										assign node1417 = (inp[5]) ? node1419 : 3'b010;
											assign node1419 = (inp[11]) ? 3'b000 : node1420;
												assign node1420 = (inp[6]) ? 3'b010 : 3'b000;
									assign node1424 = (inp[0]) ? node1430 : node1425;
										assign node1425 = (inp[11]) ? 3'b000 : node1426;
											assign node1426 = (inp[5]) ? 3'b000 : 3'b100;
										assign node1430 = (inp[5]) ? node1432 : 3'b100;
											assign node1432 = (inp[6]) ? 3'b100 : 3'b000;
						assign node1435 = (inp[5]) ? node1491 : node1436;
							assign node1436 = (inp[3]) ? node1458 : node1437;
								assign node1437 = (inp[8]) ? node1447 : node1438;
									assign node1438 = (inp[11]) ? 3'b000 : node1439;
										assign node1439 = (inp[0]) ? node1441 : 3'b000;
											assign node1441 = (inp[6]) ? 3'b000 : node1442;
												assign node1442 = (inp[4]) ? 3'b010 : 3'b000;
									assign node1447 = (inp[0]) ? 3'b000 : node1448;
										assign node1448 = (inp[11]) ? node1454 : node1449;
											assign node1449 = (inp[4]) ? node1451 : 3'b000;
												assign node1451 = (inp[6]) ? 3'b010 : 3'b000;
											assign node1454 = (inp[4]) ? 3'b000 : 3'b010;
								assign node1458 = (inp[4]) ? node1476 : node1459;
									assign node1459 = (inp[6]) ? node1467 : node1460;
										assign node1460 = (inp[11]) ? node1462 : 3'b010;
											assign node1462 = (inp[8]) ? node1464 : 3'b010;
												assign node1464 = (inp[0]) ? 3'b010 : 3'b000;
										assign node1467 = (inp[8]) ? node1471 : node1468;
											assign node1468 = (inp[0]) ? 3'b000 : 3'b010;
											assign node1471 = (inp[0]) ? node1473 : 3'b000;
												assign node1473 = (inp[11]) ? 3'b010 : 3'b000;
									assign node1476 = (inp[11]) ? 3'b000 : node1477;
										assign node1477 = (inp[8]) ? node1483 : node1478;
											assign node1478 = (inp[6]) ? node1480 : 3'b000;
												assign node1480 = (inp[0]) ? 3'b000 : 3'b010;
											assign node1483 = (inp[0]) ? node1487 : node1484;
												assign node1484 = (inp[6]) ? 3'b000 : 3'b010;
												assign node1487 = (inp[6]) ? 3'b010 : 3'b000;
							assign node1491 = (inp[4]) ? 3'b000 : node1492;
								assign node1492 = (inp[11]) ? 3'b000 : node1493;
									assign node1493 = (inp[0]) ? node1501 : node1494;
										assign node1494 = (inp[6]) ? 3'b000 : node1495;
											assign node1495 = (inp[8]) ? node1497 : 3'b000;
												assign node1497 = (inp[3]) ? 3'b000 : 3'b010;
										assign node1501 = (inp[3]) ? 3'b010 : node1502;
											assign node1502 = (inp[8]) ? 3'b000 : node1503;
												assign node1503 = (inp[6]) ? 3'b010 : 3'b000;
			assign node1510 = (inp[0]) ? node1876 : node1511;
				assign node1511 = (inp[2]) ? node1631 : node1512;
					assign node1512 = (inp[3]) ? node1602 : node1513;
						assign node1513 = (inp[1]) ? node1537 : node1514;
							assign node1514 = (inp[7]) ? node1516 : 3'b001;
								assign node1516 = (inp[4]) ? node1526 : node1517;
									assign node1517 = (inp[8]) ? 3'b001 : node1518;
										assign node1518 = (inp[5]) ? node1520 : 3'b001;
											assign node1520 = (inp[6]) ? node1522 : 3'b000;
												assign node1522 = (inp[11]) ? 3'b000 : 3'b001;
									assign node1526 = (inp[8]) ? node1534 : node1527;
										assign node1527 = (inp[5]) ? 3'b000 : node1528;
											assign node1528 = (inp[11]) ? 3'b010 : node1529;
												assign node1529 = (inp[6]) ? 3'b000 : 3'b010;
										assign node1534 = (inp[5]) ? 3'b000 : 3'b001;
							assign node1537 = (inp[5]) ? node1571 : node1538;
								assign node1538 = (inp[6]) ? node1550 : node1539;
									assign node1539 = (inp[7]) ? node1545 : node1540;
										assign node1540 = (inp[4]) ? node1542 : 3'b010;
											assign node1542 = (inp[8]) ? 3'b010 : 3'b110;
										assign node1545 = (inp[8]) ? 3'b110 : node1546;
											assign node1546 = (inp[4]) ? 3'b010 : 3'b110;
									assign node1550 = (inp[11]) ? node1562 : node1551;
										assign node1551 = (inp[7]) ? node1557 : node1552;
											assign node1552 = (inp[4]) ? node1554 : 3'b000;
												assign node1554 = (inp[8]) ? 3'b000 : 3'b100;
											assign node1557 = (inp[4]) ? node1559 : 3'b100;
												assign node1559 = (inp[8]) ? 3'b100 : 3'b000;
										assign node1562 = (inp[7]) ? node1566 : node1563;
											assign node1563 = (inp[8]) ? 3'b010 : 3'b110;
											assign node1566 = (inp[4]) ? node1568 : 3'b110;
												assign node1568 = (inp[8]) ? 3'b110 : 3'b010;
								assign node1571 = (inp[11]) ? node1591 : node1572;
									assign node1572 = (inp[6]) ? node1580 : node1573;
										assign node1573 = (inp[7]) ? node1575 : 3'b100;
											assign node1575 = (inp[8]) ? node1577 : 3'b000;
												assign node1577 = (inp[4]) ? 3'b000 : 3'b100;
										assign node1580 = (inp[7]) ? node1586 : node1581;
											assign node1581 = (inp[8]) ? 3'b010 : node1582;
												assign node1582 = (inp[4]) ? 3'b110 : 3'b010;
											assign node1586 = (inp[4]) ? node1588 : 3'b110;
												assign node1588 = (inp[8]) ? 3'b110 : 3'b010;
									assign node1591 = (inp[7]) ? node1597 : node1592;
										assign node1592 = (inp[8]) ? node1594 : 3'b100;
											assign node1594 = (inp[4]) ? 3'b100 : 3'b000;
										assign node1597 = (inp[4]) ? 3'b000 : node1598;
											assign node1598 = (inp[8]) ? 3'b100 : 3'b000;
						assign node1602 = (inp[7]) ? node1604 : 3'b001;
							assign node1604 = (inp[1]) ? node1606 : 3'b001;
								assign node1606 = (inp[8]) ? node1622 : node1607;
									assign node1607 = (inp[4]) ? node1611 : node1608;
										assign node1608 = (inp[5]) ? 3'b000 : 3'b001;
										assign node1611 = (inp[5]) ? node1617 : node1612;
											assign node1612 = (inp[11]) ? 3'b010 : node1613;
												assign node1613 = (inp[6]) ? 3'b000 : 3'b010;
											assign node1617 = (inp[11]) ? 3'b000 : node1618;
												assign node1618 = (inp[6]) ? 3'b010 : 3'b000;
									assign node1622 = (inp[5]) ? node1624 : 3'b001;
										assign node1624 = (inp[4]) ? node1626 : 3'b001;
											assign node1626 = (inp[6]) ? node1628 : 3'b000;
												assign node1628 = (inp[11]) ? 3'b000 : 3'b001;
					assign node1631 = (inp[1]) ? node1767 : node1632;
						assign node1632 = (inp[11]) ? node1714 : node1633;
							assign node1633 = (inp[7]) ? node1673 : node1634;
								assign node1634 = (inp[8]) ? node1654 : node1635;
									assign node1635 = (inp[4]) ? node1643 : node1636;
										assign node1636 = (inp[5]) ? node1640 : node1637;
											assign node1637 = (inp[6]) ? 3'b000 : 3'b010;
											assign node1640 = (inp[6]) ? 3'b010 : 3'b100;
										assign node1643 = (inp[3]) ? node1647 : node1644;
											assign node1644 = (inp[5]) ? 3'b010 : 3'b110;
											assign node1647 = (inp[5]) ? node1651 : node1648;
												assign node1648 = (inp[6]) ? 3'b100 : 3'b110;
												assign node1651 = (inp[6]) ? 3'b110 : 3'b100;
									assign node1654 = (inp[4]) ? node1662 : node1655;
										assign node1655 = (inp[6]) ? node1659 : node1656;
											assign node1656 = (inp[5]) ? 3'b000 : 3'b010;
											assign node1659 = (inp[5]) ? 3'b010 : 3'b000;
										assign node1662 = (inp[3]) ? node1668 : node1663;
											assign node1663 = (inp[5]) ? 3'b100 : node1664;
												assign node1664 = (inp[6]) ? 3'b000 : 3'b010;
											assign node1668 = (inp[6]) ? node1670 : 3'b010;
												assign node1670 = (inp[5]) ? 3'b010 : 3'b000;
								assign node1673 = (inp[3]) ? node1687 : node1674;
									assign node1674 = (inp[4]) ? node1680 : node1675;
										assign node1675 = (inp[5]) ? node1677 : 3'b010;
											assign node1677 = (inp[8]) ? 3'b010 : 3'b110;
										assign node1680 = (inp[5]) ? node1682 : 3'b110;
											assign node1682 = (inp[8]) ? 3'b110 : node1683;
												assign node1683 = (inp[6]) ? 3'b000 : 3'b010;
									assign node1687 = (inp[8]) ? node1699 : node1688;
										assign node1688 = (inp[4]) ? node1696 : node1689;
											assign node1689 = (inp[5]) ? node1693 : node1690;
												assign node1690 = (inp[6]) ? 3'b100 : 3'b110;
												assign node1693 = (inp[6]) ? 3'b110 : 3'b000;
											assign node1696 = (inp[5]) ? 3'b010 : 3'b000;
										assign node1699 = (inp[4]) ? node1707 : node1700;
											assign node1700 = (inp[5]) ? node1704 : node1701;
												assign node1701 = (inp[6]) ? 3'b100 : 3'b110;
												assign node1704 = (inp[6]) ? 3'b110 : 3'b100;
											assign node1707 = (inp[6]) ? node1711 : node1708;
												assign node1708 = (inp[5]) ? 3'b000 : 3'b110;
												assign node1711 = (inp[5]) ? 3'b110 : 3'b100;
							assign node1714 = (inp[5]) ? node1740 : node1715;
								assign node1715 = (inp[7]) ? node1727 : node1716;
									assign node1716 = (inp[3]) ? node1722 : node1717;
										assign node1717 = (inp[8]) ? 3'b010 : node1718;
											assign node1718 = (inp[4]) ? 3'b000 : 3'b010;
										assign node1722 = (inp[8]) ? 3'b010 : node1723;
											assign node1723 = (inp[4]) ? 3'b110 : 3'b010;
									assign node1727 = (inp[3]) ? node1735 : node1728;
										assign node1728 = (inp[4]) ? node1732 : node1729;
											assign node1729 = (inp[8]) ? 3'b000 : 3'b100;
											assign node1732 = (inp[8]) ? 3'b100 : 3'b000;
										assign node1735 = (inp[8]) ? 3'b110 : node1736;
											assign node1736 = (inp[4]) ? 3'b000 : 3'b110;
								assign node1740 = (inp[4]) ? node1762 : node1741;
									assign node1741 = (inp[3]) ? node1747 : node1742;
										assign node1742 = (inp[8]) ? node1744 : 3'b100;
											assign node1744 = (inp[7]) ? 3'b100 : 3'b000;
										assign node1747 = (inp[6]) ? node1755 : node1748;
											assign node1748 = (inp[7]) ? node1752 : node1749;
												assign node1749 = (inp[8]) ? 3'b000 : 3'b100;
												assign node1752 = (inp[8]) ? 3'b100 : 3'b000;
											assign node1755 = (inp[7]) ? node1759 : node1756;
												assign node1756 = (inp[8]) ? 3'b000 : 3'b100;
												assign node1759 = (inp[8]) ? 3'b100 : 3'b000;
									assign node1762 = (inp[3]) ? node1764 : 3'b000;
										assign node1764 = (inp[7]) ? 3'b000 : 3'b100;
						assign node1767 = (inp[7]) ? node1835 : node1768;
							assign node1768 = (inp[5]) ? node1802 : node1769;
								assign node1769 = (inp[8]) ? node1783 : node1770;
									assign node1770 = (inp[4]) ? node1778 : node1771;
										assign node1771 = (inp[11]) ? node1775 : node1772;
											assign node1772 = (inp[3]) ? 3'b010 : 3'b100;
											assign node1775 = (inp[3]) ? 3'b100 : 3'b110;
										assign node1778 = (inp[11]) ? 3'b010 : node1779;
											assign node1779 = (inp[6]) ? 3'b010 : 3'b000;
									assign node1783 = (inp[4]) ? node1793 : node1784;
										assign node1784 = (inp[11]) ? node1790 : node1785;
											assign node1785 = (inp[6]) ? 3'b010 : node1786;
												assign node1786 = (inp[3]) ? 3'b010 : 3'b000;
											assign node1790 = (inp[3]) ? 3'b000 : 3'b010;
										assign node1793 = (inp[3]) ? node1797 : node1794;
											assign node1794 = (inp[11]) ? 3'b100 : 3'b000;
											assign node1797 = (inp[11]) ? 3'b010 : node1798;
												assign node1798 = (inp[6]) ? 3'b110 : 3'b000;
								assign node1802 = (inp[11]) ? node1828 : node1803;
									assign node1803 = (inp[4]) ? node1813 : node1804;
										assign node1804 = (inp[3]) ? node1810 : node1805;
											assign node1805 = (inp[8]) ? node1807 : 3'b000;
												assign node1807 = (inp[6]) ? 3'b100 : 3'b110;
											assign node1810 = (inp[8]) ? 3'b010 : 3'b110;
										assign node1813 = (inp[8]) ? node1821 : node1814;
											assign node1814 = (inp[6]) ? node1818 : node1815;
												assign node1815 = (inp[3]) ? 3'b000 : 3'b100;
												assign node1818 = (inp[3]) ? 3'b000 : 3'b010;
											assign node1821 = (inp[6]) ? node1825 : node1822;
												assign node1822 = (inp[3]) ? 3'b010 : 3'b000;
												assign node1825 = (inp[3]) ? 3'b000 : 3'b010;
									assign node1828 = (inp[3]) ? node1830 : 3'b000;
										assign node1830 = (inp[8]) ? node1832 : 3'b000;
											assign node1832 = (inp[4]) ? 3'b000 : 3'b100;
							assign node1835 = (inp[4]) ? node1861 : node1836;
								assign node1836 = (inp[11]) ? node1854 : node1837;
									assign node1837 = (inp[5]) ? node1847 : node1838;
										assign node1838 = (inp[3]) ? node1842 : node1839;
											assign node1839 = (inp[6]) ? 3'b010 : 3'b000;
											assign node1842 = (inp[6]) ? 3'b000 : node1843;
												assign node1843 = (inp[8]) ? 3'b000 : 3'b010;
										assign node1847 = (inp[6]) ? node1849 : 3'b010;
											assign node1849 = (inp[3]) ? node1851 : 3'b010;
												assign node1851 = (inp[8]) ? 3'b010 : 3'b000;
									assign node1854 = (inp[5]) ? 3'b000 : node1855;
										assign node1855 = (inp[8]) ? node1857 : 3'b000;
											assign node1857 = (inp[6]) ? 3'b010 : 3'b000;
								assign node1861 = (inp[5]) ? 3'b000 : node1862;
									assign node1862 = (inp[11]) ? 3'b000 : node1863;
										assign node1863 = (inp[3]) ? node1869 : node1864;
											assign node1864 = (inp[6]) ? 3'b000 : node1865;
												assign node1865 = (inp[8]) ? 3'b000 : 3'b010;
											assign node1869 = (inp[6]) ? node1871 : 3'b000;
												assign node1871 = (inp[8]) ? 3'b010 : 3'b000;
				assign node1876 = (inp[2]) ? node1878 : 3'b000;
					assign node1878 = (inp[3]) ? node1954 : node1879;
						assign node1879 = (inp[1]) ? node1897 : node1880;
							assign node1880 = (inp[8]) ? 3'b000 : node1881;
								assign node1881 = (inp[7]) ? node1883 : 3'b000;
									assign node1883 = (inp[4]) ? node1885 : 3'b000;
										assign node1885 = (inp[5]) ? node1891 : node1886;
											assign node1886 = (inp[6]) ? node1888 : 3'b010;
												assign node1888 = (inp[11]) ? 3'b010 : 3'b000;
											assign node1891 = (inp[11]) ? 3'b000 : node1892;
												assign node1892 = (inp[6]) ? 3'b010 : 3'b000;
							assign node1897 = (inp[5]) ? node1931 : node1898;
								assign node1898 = (inp[4]) ? node1914 : node1899;
									assign node1899 = (inp[11]) ? node1909 : node1900;
										assign node1900 = (inp[6]) ? node1906 : node1901;
											assign node1901 = (inp[8]) ? 3'b010 : node1902;
												assign node1902 = (inp[7]) ? 3'b000 : 3'b010;
											assign node1906 = (inp[7]) ? 3'b010 : 3'b000;
										assign node1909 = (inp[8]) ? node1911 : 3'b010;
											assign node1911 = (inp[7]) ? 3'b000 : 3'b010;
									assign node1914 = (inp[8]) ? node1920 : node1915;
										assign node1915 = (inp[11]) ? 3'b000 : node1916;
											assign node1916 = (inp[6]) ? 3'b010 : 3'b000;
										assign node1920 = (inp[6]) ? node1926 : node1921;
											assign node1921 = (inp[7]) ? node1923 : 3'b010;
												assign node1923 = (inp[11]) ? 3'b000 : 3'b010;
											assign node1926 = (inp[11]) ? node1928 : 3'b000;
												assign node1928 = (inp[7]) ? 3'b000 : 3'b010;
								assign node1931 = (inp[11]) ? node1947 : node1932;
									assign node1932 = (inp[7]) ? node1942 : node1933;
										assign node1933 = (inp[6]) ? 3'b010 : node1934;
											assign node1934 = (inp[4]) ? node1938 : node1935;
												assign node1935 = (inp[8]) ? 3'b000 : 3'b100;
												assign node1938 = (inp[8]) ? 3'b100 : 3'b010;
										assign node1942 = (inp[6]) ? 3'b000 : node1943;
											assign node1943 = (inp[8]) ? 3'b010 : 3'b000;
									assign node1947 = (inp[8]) ? 3'b000 : node1948;
										assign node1948 = (inp[4]) ? 3'b000 : node1949;
											assign node1949 = (inp[7]) ? 3'b000 : 3'b100;
						assign node1954 = (inp[5]) ? 3'b000 : node1955;
							assign node1955 = (inp[7]) ? node1957 : 3'b000;
								assign node1957 = (inp[11]) ? 3'b000 : node1958;
									assign node1958 = (inp[1]) ? node1960 : 3'b000;
										assign node1960 = (inp[4]) ? node1962 : 3'b000;
											assign node1962 = (inp[8]) ? 3'b000 : 3'b010;

endmodule