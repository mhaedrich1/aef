module dtc_split75_bm61 (
	input  wire [12-1:0] inp,
	output wire [11-1:0] outp
);

	wire [11-1:0] node1;
	wire [11-1:0] node2;
	wire [11-1:0] node3;
	wire [11-1:0] node4;
	wire [11-1:0] node5;
	wire [11-1:0] node6;
	wire [11-1:0] node7;
	wire [11-1:0] node8;
	wire [11-1:0] node9;
	wire [11-1:0] node10;
	wire [11-1:0] node12;
	wire [11-1:0] node15;
	wire [11-1:0] node18;
	wire [11-1:0] node19;
	wire [11-1:0] node22;
	wire [11-1:0] node25;
	wire [11-1:0] node26;
	wire [11-1:0] node27;
	wire [11-1:0] node28;
	wire [11-1:0] node32;
	wire [11-1:0] node35;
	wire [11-1:0] node36;
	wire [11-1:0] node37;
	wire [11-1:0] node40;
	wire [11-1:0] node43;
	wire [11-1:0] node45;
	wire [11-1:0] node48;
	wire [11-1:0] node49;
	wire [11-1:0] node50;
	wire [11-1:0] node51;
	wire [11-1:0] node52;
	wire [11-1:0] node55;
	wire [11-1:0] node58;
	wire [11-1:0] node61;
	wire [11-1:0] node62;
	wire [11-1:0] node64;
	wire [11-1:0] node67;
	wire [11-1:0] node70;
	wire [11-1:0] node71;
	wire [11-1:0] node72;
	wire [11-1:0] node73;
	wire [11-1:0] node77;
	wire [11-1:0] node80;
	wire [11-1:0] node81;
	wire [11-1:0] node82;
	wire [11-1:0] node85;
	wire [11-1:0] node88;
	wire [11-1:0] node90;
	wire [11-1:0] node93;
	wire [11-1:0] node94;
	wire [11-1:0] node95;
	wire [11-1:0] node96;
	wire [11-1:0] node97;
	wire [11-1:0] node98;
	wire [11-1:0] node101;
	wire [11-1:0] node104;
	wire [11-1:0] node105;
	wire [11-1:0] node108;
	wire [11-1:0] node111;
	wire [11-1:0] node112;
	wire [11-1:0] node113;
	wire [11-1:0] node117;
	wire [11-1:0] node118;
	wire [11-1:0] node121;
	wire [11-1:0] node124;
	wire [11-1:0] node125;
	wire [11-1:0] node126;
	wire [11-1:0] node127;
	wire [11-1:0] node131;
	wire [11-1:0] node132;
	wire [11-1:0] node135;
	wire [11-1:0] node138;
	wire [11-1:0] node139;
	wire [11-1:0] node140;
	wire [11-1:0] node143;
	wire [11-1:0] node146;
	wire [11-1:0] node147;
	wire [11-1:0] node150;
	wire [11-1:0] node153;
	wire [11-1:0] node154;
	wire [11-1:0] node155;
	wire [11-1:0] node156;
	wire [11-1:0] node157;
	wire [11-1:0] node160;
	wire [11-1:0] node163;
	wire [11-1:0] node164;
	wire [11-1:0] node167;
	wire [11-1:0] node170;
	wire [11-1:0] node171;
	wire [11-1:0] node172;
	wire [11-1:0] node176;
	wire [11-1:0] node178;
	wire [11-1:0] node181;
	wire [11-1:0] node182;
	wire [11-1:0] node183;
	wire [11-1:0] node184;
	wire [11-1:0] node188;
	wire [11-1:0] node190;
	wire [11-1:0] node193;
	wire [11-1:0] node194;
	wire [11-1:0] node195;
	wire [11-1:0] node198;
	wire [11-1:0] node201;
	wire [11-1:0] node203;
	wire [11-1:0] node206;
	wire [11-1:0] node207;
	wire [11-1:0] node208;
	wire [11-1:0] node209;
	wire [11-1:0] node210;
	wire [11-1:0] node211;
	wire [11-1:0] node214;
	wire [11-1:0] node216;
	wire [11-1:0] node219;
	wire [11-1:0] node220;
	wire [11-1:0] node223;
	wire [11-1:0] node224;
	wire [11-1:0] node228;
	wire [11-1:0] node229;
	wire [11-1:0] node230;
	wire [11-1:0] node231;
	wire [11-1:0] node235;
	wire [11-1:0] node236;
	wire [11-1:0] node239;
	wire [11-1:0] node242;
	wire [11-1:0] node243;
	wire [11-1:0] node244;
	wire [11-1:0] node247;
	wire [11-1:0] node250;
	wire [11-1:0] node251;
	wire [11-1:0] node255;
	wire [11-1:0] node256;
	wire [11-1:0] node257;
	wire [11-1:0] node258;
	wire [11-1:0] node261;
	wire [11-1:0] node264;
	wire [11-1:0] node265;
	wire [11-1:0] node266;
	wire [11-1:0] node269;
	wire [11-1:0] node272;
	wire [11-1:0] node273;
	wire [11-1:0] node277;
	wire [11-1:0] node278;
	wire [11-1:0] node279;
	wire [11-1:0] node280;
	wire [11-1:0] node283;
	wire [11-1:0] node286;
	wire [11-1:0] node288;
	wire [11-1:0] node291;
	wire [11-1:0] node292;
	wire [11-1:0] node295;
	wire [11-1:0] node296;
	wire [11-1:0] node300;
	wire [11-1:0] node301;
	wire [11-1:0] node302;
	wire [11-1:0] node303;
	wire [11-1:0] node304;
	wire [11-1:0] node305;
	wire [11-1:0] node309;
	wire [11-1:0] node310;
	wire [11-1:0] node313;
	wire [11-1:0] node316;
	wire [11-1:0] node317;
	wire [11-1:0] node321;
	wire [11-1:0] node322;
	wire [11-1:0] node323;
	wire [11-1:0] node325;
	wire [11-1:0] node328;
	wire [11-1:0] node331;
	wire [11-1:0] node332;
	wire [11-1:0] node334;
	wire [11-1:0] node337;
	wire [11-1:0] node338;
	wire [11-1:0] node341;
	wire [11-1:0] node344;
	wire [11-1:0] node345;
	wire [11-1:0] node346;
	wire [11-1:0] node347;
	wire [11-1:0] node348;
	wire [11-1:0] node352;
	wire [11-1:0] node353;
	wire [11-1:0] node356;
	wire [11-1:0] node359;
	wire [11-1:0] node360;
	wire [11-1:0] node363;
	wire [11-1:0] node365;
	wire [11-1:0] node368;
	wire [11-1:0] node369;
	wire [11-1:0] node370;
	wire [11-1:0] node372;
	wire [11-1:0] node376;
	wire [11-1:0] node377;
	wire [11-1:0] node378;
	wire [11-1:0] node381;
	wire [11-1:0] node384;
	wire [11-1:0] node387;
	wire [11-1:0] node388;
	wire [11-1:0] node389;
	wire [11-1:0] node390;
	wire [11-1:0] node391;
	wire [11-1:0] node392;
	wire [11-1:0] node393;
	wire [11-1:0] node394;
	wire [11-1:0] node397;
	wire [11-1:0] node400;
	wire [11-1:0] node402;
	wire [11-1:0] node405;
	wire [11-1:0] node406;
	wire [11-1:0] node409;
	wire [11-1:0] node410;
	wire [11-1:0] node414;
	wire [11-1:0] node415;
	wire [11-1:0] node416;
	wire [11-1:0] node417;
	wire [11-1:0] node420;
	wire [11-1:0] node423;
	wire [11-1:0] node424;
	wire [11-1:0] node427;
	wire [11-1:0] node430;
	wire [11-1:0] node431;
	wire [11-1:0] node433;
	wire [11-1:0] node436;
	wire [11-1:0] node437;
	wire [11-1:0] node441;
	wire [11-1:0] node442;
	wire [11-1:0] node443;
	wire [11-1:0] node444;
	wire [11-1:0] node446;
	wire [11-1:0] node449;
	wire [11-1:0] node451;
	wire [11-1:0] node454;
	wire [11-1:0] node455;
	wire [11-1:0] node457;
	wire [11-1:0] node460;
	wire [11-1:0] node461;
	wire [11-1:0] node464;
	wire [11-1:0] node467;
	wire [11-1:0] node468;
	wire [11-1:0] node469;
	wire [11-1:0] node470;
	wire [11-1:0] node473;
	wire [11-1:0] node476;
	wire [11-1:0] node479;
	wire [11-1:0] node480;
	wire [11-1:0] node483;
	wire [11-1:0] node484;
	wire [11-1:0] node487;
	wire [11-1:0] node490;
	wire [11-1:0] node491;
	wire [11-1:0] node492;
	wire [11-1:0] node493;
	wire [11-1:0] node494;
	wire [11-1:0] node495;
	wire [11-1:0] node499;
	wire [11-1:0] node501;
	wire [11-1:0] node504;
	wire [11-1:0] node505;
	wire [11-1:0] node506;
	wire [11-1:0] node510;
	wire [11-1:0] node512;
	wire [11-1:0] node515;
	wire [11-1:0] node516;
	wire [11-1:0] node517;
	wire [11-1:0] node518;
	wire [11-1:0] node521;
	wire [11-1:0] node524;
	wire [11-1:0] node525;
	wire [11-1:0] node529;
	wire [11-1:0] node530;
	wire [11-1:0] node533;
	wire [11-1:0] node534;
	wire [11-1:0] node537;
	wire [11-1:0] node540;
	wire [11-1:0] node541;
	wire [11-1:0] node542;
	wire [11-1:0] node543;
	wire [11-1:0] node544;
	wire [11-1:0] node548;
	wire [11-1:0] node549;
	wire [11-1:0] node552;
	wire [11-1:0] node555;
	wire [11-1:0] node556;
	wire [11-1:0] node558;
	wire [11-1:0] node562;
	wire [11-1:0] node563;
	wire [11-1:0] node564;
	wire [11-1:0] node565;
	wire [11-1:0] node568;
	wire [11-1:0] node572;
	wire [11-1:0] node573;
	wire [11-1:0] node576;
	wire [11-1:0] node578;
	wire [11-1:0] node581;
	wire [11-1:0] node582;
	wire [11-1:0] node583;
	wire [11-1:0] node584;
	wire [11-1:0] node585;
	wire [11-1:0] node586;
	wire [11-1:0] node588;
	wire [11-1:0] node591;
	wire [11-1:0] node594;
	wire [11-1:0] node595;
	wire [11-1:0] node597;
	wire [11-1:0] node600;
	wire [11-1:0] node601;
	wire [11-1:0] node604;
	wire [11-1:0] node607;
	wire [11-1:0] node608;
	wire [11-1:0] node609;
	wire [11-1:0] node610;
	wire [11-1:0] node614;
	wire [11-1:0] node617;
	wire [11-1:0] node618;
	wire [11-1:0] node621;
	wire [11-1:0] node624;
	wire [11-1:0] node625;
	wire [11-1:0] node626;
	wire [11-1:0] node627;
	wire [11-1:0] node630;
	wire [11-1:0] node633;
	wire [11-1:0] node635;
	wire [11-1:0] node637;
	wire [11-1:0] node640;
	wire [11-1:0] node641;
	wire [11-1:0] node642;
	wire [11-1:0] node644;
	wire [11-1:0] node647;
	wire [11-1:0] node649;
	wire [11-1:0] node652;
	wire [11-1:0] node653;
	wire [11-1:0] node654;
	wire [11-1:0] node658;
	wire [11-1:0] node659;
	wire [11-1:0] node663;
	wire [11-1:0] node664;
	wire [11-1:0] node665;
	wire [11-1:0] node666;
	wire [11-1:0] node667;
	wire [11-1:0] node670;
	wire [11-1:0] node673;
	wire [11-1:0] node674;
	wire [11-1:0] node677;
	wire [11-1:0] node678;
	wire [11-1:0] node682;
	wire [11-1:0] node683;
	wire [11-1:0] node684;
	wire [11-1:0] node687;
	wire [11-1:0] node689;
	wire [11-1:0] node692;
	wire [11-1:0] node693;
	wire [11-1:0] node696;
	wire [11-1:0] node697;
	wire [11-1:0] node701;
	wire [11-1:0] node702;
	wire [11-1:0] node703;
	wire [11-1:0] node704;
	wire [11-1:0] node705;
	wire [11-1:0] node709;
	wire [11-1:0] node711;
	wire [11-1:0] node714;
	wire [11-1:0] node715;
	wire [11-1:0] node718;
	wire [11-1:0] node719;
	wire [11-1:0] node722;
	wire [11-1:0] node725;
	wire [11-1:0] node726;
	wire [11-1:0] node727;
	wire [11-1:0] node728;
	wire [11-1:0] node732;
	wire [11-1:0] node733;
	wire [11-1:0] node736;
	wire [11-1:0] node739;
	wire [11-1:0] node741;
	wire [11-1:0] node742;
	wire [11-1:0] node746;
	wire [11-1:0] node747;
	wire [11-1:0] node748;
	wire [11-1:0] node749;
	wire [11-1:0] node750;
	wire [11-1:0] node751;
	wire [11-1:0] node752;
	wire [11-1:0] node753;
	wire [11-1:0] node754;
	wire [11-1:0] node758;
	wire [11-1:0] node761;
	wire [11-1:0] node763;
	wire [11-1:0] node764;
	wire [11-1:0] node768;
	wire [11-1:0] node769;
	wire [11-1:0] node770;
	wire [11-1:0] node771;
	wire [11-1:0] node774;
	wire [11-1:0] node777;
	wire [11-1:0] node778;
	wire [11-1:0] node782;
	wire [11-1:0] node783;
	wire [11-1:0] node784;
	wire [11-1:0] node789;
	wire [11-1:0] node790;
	wire [11-1:0] node791;
	wire [11-1:0] node792;
	wire [11-1:0] node793;
	wire [11-1:0] node797;
	wire [11-1:0] node798;
	wire [11-1:0] node802;
	wire [11-1:0] node803;
	wire [11-1:0] node805;
	wire [11-1:0] node808;
	wire [11-1:0] node809;
	wire [11-1:0] node812;
	wire [11-1:0] node815;
	wire [11-1:0] node816;
	wire [11-1:0] node817;
	wire [11-1:0] node818;
	wire [11-1:0] node821;
	wire [11-1:0] node824;
	wire [11-1:0] node827;
	wire [11-1:0] node828;
	wire [11-1:0] node831;
	wire [11-1:0] node832;
	wire [11-1:0] node835;
	wire [11-1:0] node838;
	wire [11-1:0] node839;
	wire [11-1:0] node840;
	wire [11-1:0] node841;
	wire [11-1:0] node842;
	wire [11-1:0] node843;
	wire [11-1:0] node846;
	wire [11-1:0] node849;
	wire [11-1:0] node850;
	wire [11-1:0] node853;
	wire [11-1:0] node856;
	wire [11-1:0] node857;
	wire [11-1:0] node859;
	wire [11-1:0] node862;
	wire [11-1:0] node864;
	wire [11-1:0] node867;
	wire [11-1:0] node868;
	wire [11-1:0] node869;
	wire [11-1:0] node870;
	wire [11-1:0] node873;
	wire [11-1:0] node876;
	wire [11-1:0] node879;
	wire [11-1:0] node880;
	wire [11-1:0] node881;
	wire [11-1:0] node884;
	wire [11-1:0] node887;
	wire [11-1:0] node888;
	wire [11-1:0] node891;
	wire [11-1:0] node894;
	wire [11-1:0] node895;
	wire [11-1:0] node896;
	wire [11-1:0] node897;
	wire [11-1:0] node900;
	wire [11-1:0] node903;
	wire [11-1:0] node904;
	wire [11-1:0] node905;
	wire [11-1:0] node909;
	wire [11-1:0] node910;
	wire [11-1:0] node913;
	wire [11-1:0] node916;
	wire [11-1:0] node917;
	wire [11-1:0] node918;
	wire [11-1:0] node921;
	wire [11-1:0] node924;
	wire [11-1:0] node925;
	wire [11-1:0] node926;
	wire [11-1:0] node929;
	wire [11-1:0] node932;
	wire [11-1:0] node935;
	wire [11-1:0] node936;
	wire [11-1:0] node937;
	wire [11-1:0] node938;
	wire [11-1:0] node939;
	wire [11-1:0] node940;
	wire [11-1:0] node943;
	wire [11-1:0] node946;
	wire [11-1:0] node947;
	wire [11-1:0] node949;
	wire [11-1:0] node952;
	wire [11-1:0] node954;
	wire [11-1:0] node957;
	wire [11-1:0] node958;
	wire [11-1:0] node959;
	wire [11-1:0] node961;
	wire [11-1:0] node964;
	wire [11-1:0] node965;
	wire [11-1:0] node968;
	wire [11-1:0] node971;
	wire [11-1:0] node972;
	wire [11-1:0] node973;
	wire [11-1:0] node976;
	wire [11-1:0] node979;
	wire [11-1:0] node982;
	wire [11-1:0] node983;
	wire [11-1:0] node984;
	wire [11-1:0] node985;
	wire [11-1:0] node988;
	wire [11-1:0] node990;
	wire [11-1:0] node993;
	wire [11-1:0] node994;
	wire [11-1:0] node995;
	wire [11-1:0] node999;
	wire [11-1:0] node1002;
	wire [11-1:0] node1003;
	wire [11-1:0] node1004;
	wire [11-1:0] node1007;
	wire [11-1:0] node1008;
	wire [11-1:0] node1011;
	wire [11-1:0] node1014;
	wire [11-1:0] node1016;
	wire [11-1:0] node1018;
	wire [11-1:0] node1021;
	wire [11-1:0] node1022;
	wire [11-1:0] node1023;
	wire [11-1:0] node1024;
	wire [11-1:0] node1025;
	wire [11-1:0] node1026;
	wire [11-1:0] node1029;
	wire [11-1:0] node1032;
	wire [11-1:0] node1033;
	wire [11-1:0] node1037;
	wire [11-1:0] node1038;
	wire [11-1:0] node1039;
	wire [11-1:0] node1043;
	wire [11-1:0] node1044;
	wire [11-1:0] node1048;
	wire [11-1:0] node1049;
	wire [11-1:0] node1050;
	wire [11-1:0] node1051;
	wire [11-1:0] node1054;
	wire [11-1:0] node1057;
	wire [11-1:0] node1058;
	wire [11-1:0] node1061;
	wire [11-1:0] node1064;
	wire [11-1:0] node1065;
	wire [11-1:0] node1066;
	wire [11-1:0] node1070;
	wire [11-1:0] node1073;
	wire [11-1:0] node1074;
	wire [11-1:0] node1075;
	wire [11-1:0] node1076;
	wire [11-1:0] node1077;
	wire [11-1:0] node1080;
	wire [11-1:0] node1083;
	wire [11-1:0] node1085;
	wire [11-1:0] node1088;
	wire [11-1:0] node1089;
	wire [11-1:0] node1090;
	wire [11-1:0] node1094;
	wire [11-1:0] node1095;
	wire [11-1:0] node1099;
	wire [11-1:0] node1100;
	wire [11-1:0] node1101;
	wire [11-1:0] node1104;
	wire [11-1:0] node1106;
	wire [11-1:0] node1109;
	wire [11-1:0] node1110;
	wire [11-1:0] node1113;
	wire [11-1:0] node1115;
	wire [11-1:0] node1118;
	wire [11-1:0] node1119;
	wire [11-1:0] node1120;
	wire [11-1:0] node1121;
	wire [11-1:0] node1122;
	wire [11-1:0] node1123;
	wire [11-1:0] node1124;
	wire [11-1:0] node1125;
	wire [11-1:0] node1129;
	wire [11-1:0] node1130;
	wire [11-1:0] node1133;
	wire [11-1:0] node1136;
	wire [11-1:0] node1138;
	wire [11-1:0] node1141;
	wire [11-1:0] node1142;
	wire [11-1:0] node1143;
	wire [11-1:0] node1146;
	wire [11-1:0] node1148;
	wire [11-1:0] node1151;
	wire [11-1:0] node1152;
	wire [11-1:0] node1153;
	wire [11-1:0] node1156;
	wire [11-1:0] node1159;
	wire [11-1:0] node1161;
	wire [11-1:0] node1164;
	wire [11-1:0] node1165;
	wire [11-1:0] node1166;
	wire [11-1:0] node1167;
	wire [11-1:0] node1169;
	wire [11-1:0] node1172;
	wire [11-1:0] node1175;
	wire [11-1:0] node1176;
	wire [11-1:0] node1177;
	wire [11-1:0] node1180;
	wire [11-1:0] node1183;
	wire [11-1:0] node1184;
	wire [11-1:0] node1187;
	wire [11-1:0] node1190;
	wire [11-1:0] node1191;
	wire [11-1:0] node1192;
	wire [11-1:0] node1194;
	wire [11-1:0] node1197;
	wire [11-1:0] node1198;
	wire [11-1:0] node1201;
	wire [11-1:0] node1204;
	wire [11-1:0] node1205;
	wire [11-1:0] node1206;
	wire [11-1:0] node1210;
	wire [11-1:0] node1213;
	wire [11-1:0] node1214;
	wire [11-1:0] node1215;
	wire [11-1:0] node1216;
	wire [11-1:0] node1217;
	wire [11-1:0] node1218;
	wire [11-1:0] node1221;
	wire [11-1:0] node1224;
	wire [11-1:0] node1225;
	wire [11-1:0] node1228;
	wire [11-1:0] node1231;
	wire [11-1:0] node1232;
	wire [11-1:0] node1233;
	wire [11-1:0] node1236;
	wire [11-1:0] node1239;
	wire [11-1:0] node1240;
	wire [11-1:0] node1244;
	wire [11-1:0] node1245;
	wire [11-1:0] node1246;
	wire [11-1:0] node1247;
	wire [11-1:0] node1251;
	wire [11-1:0] node1254;
	wire [11-1:0] node1255;
	wire [11-1:0] node1257;
	wire [11-1:0] node1260;
	wire [11-1:0] node1262;
	wire [11-1:0] node1265;
	wire [11-1:0] node1266;
	wire [11-1:0] node1267;
	wire [11-1:0] node1268;
	wire [11-1:0] node1270;
	wire [11-1:0] node1273;
	wire [11-1:0] node1276;
	wire [11-1:0] node1278;
	wire [11-1:0] node1279;
	wire [11-1:0] node1282;
	wire [11-1:0] node1285;
	wire [11-1:0] node1286;
	wire [11-1:0] node1287;
	wire [11-1:0] node1288;
	wire [11-1:0] node1292;
	wire [11-1:0] node1295;
	wire [11-1:0] node1296;
	wire [11-1:0] node1298;
	wire [11-1:0] node1301;
	wire [11-1:0] node1302;
	wire [11-1:0] node1306;
	wire [11-1:0] node1307;
	wire [11-1:0] node1308;
	wire [11-1:0] node1309;
	wire [11-1:0] node1310;
	wire [11-1:0] node1311;
	wire [11-1:0] node1312;
	wire [11-1:0] node1316;
	wire [11-1:0] node1317;
	wire [11-1:0] node1321;
	wire [11-1:0] node1322;
	wire [11-1:0] node1323;
	wire [11-1:0] node1326;
	wire [11-1:0] node1329;
	wire [11-1:0] node1330;
	wire [11-1:0] node1333;
	wire [11-1:0] node1336;
	wire [11-1:0] node1337;
	wire [11-1:0] node1338;
	wire [11-1:0] node1341;
	wire [11-1:0] node1342;
	wire [11-1:0] node1346;
	wire [11-1:0] node1347;
	wire [11-1:0] node1349;
	wire [11-1:0] node1352;
	wire [11-1:0] node1353;
	wire [11-1:0] node1357;
	wire [11-1:0] node1358;
	wire [11-1:0] node1359;
	wire [11-1:0] node1360;
	wire [11-1:0] node1362;
	wire [11-1:0] node1365;
	wire [11-1:0] node1367;
	wire [11-1:0] node1370;
	wire [11-1:0] node1371;
	wire [11-1:0] node1373;
	wire [11-1:0] node1376;
	wire [11-1:0] node1378;
	wire [11-1:0] node1381;
	wire [11-1:0] node1382;
	wire [11-1:0] node1383;
	wire [11-1:0] node1384;
	wire [11-1:0] node1387;
	wire [11-1:0] node1390;
	wire [11-1:0] node1391;
	wire [11-1:0] node1394;
	wire [11-1:0] node1397;
	wire [11-1:0] node1398;
	wire [11-1:0] node1399;
	wire [11-1:0] node1403;
	wire [11-1:0] node1406;
	wire [11-1:0] node1407;
	wire [11-1:0] node1408;
	wire [11-1:0] node1409;
	wire [11-1:0] node1411;
	wire [11-1:0] node1412;
	wire [11-1:0] node1416;
	wire [11-1:0] node1417;
	wire [11-1:0] node1418;
	wire [11-1:0] node1421;
	wire [11-1:0] node1424;
	wire [11-1:0] node1425;
	wire [11-1:0] node1428;
	wire [11-1:0] node1431;
	wire [11-1:0] node1432;
	wire [11-1:0] node1433;
	wire [11-1:0] node1434;
	wire [11-1:0] node1438;
	wire [11-1:0] node1439;
	wire [11-1:0] node1442;
	wire [11-1:0] node1445;
	wire [11-1:0] node1446;
	wire [11-1:0] node1447;
	wire [11-1:0] node1451;
	wire [11-1:0] node1453;
	wire [11-1:0] node1456;
	wire [11-1:0] node1457;
	wire [11-1:0] node1458;
	wire [11-1:0] node1459;
	wire [11-1:0] node1460;
	wire [11-1:0] node1463;
	wire [11-1:0] node1466;
	wire [11-1:0] node1467;
	wire [11-1:0] node1470;
	wire [11-1:0] node1473;
	wire [11-1:0] node1474;
	wire [11-1:0] node1476;
	wire [11-1:0] node1479;
	wire [11-1:0] node1482;
	wire [11-1:0] node1483;
	wire [11-1:0] node1484;
	wire [11-1:0] node1485;
	wire [11-1:0] node1489;
	wire [11-1:0] node1490;
	wire [11-1:0] node1494;
	wire [11-1:0] node1495;
	wire [11-1:0] node1498;
	wire [11-1:0] node1499;
	wire [11-1:0] node1503;
	wire [11-1:0] node1504;
	wire [11-1:0] node1505;
	wire [11-1:0] node1506;
	wire [11-1:0] node1507;
	wire [11-1:0] node1508;
	wire [11-1:0] node1509;
	wire [11-1:0] node1510;
	wire [11-1:0] node1511;
	wire [11-1:0] node1513;
	wire [11-1:0] node1516;
	wire [11-1:0] node1517;
	wire [11-1:0] node1520;
	wire [11-1:0] node1523;
	wire [11-1:0] node1524;
	wire [11-1:0] node1525;
	wire [11-1:0] node1529;
	wire [11-1:0] node1530;
	wire [11-1:0] node1534;
	wire [11-1:0] node1535;
	wire [11-1:0] node1536;
	wire [11-1:0] node1537;
	wire [11-1:0] node1540;
	wire [11-1:0] node1543;
	wire [11-1:0] node1544;
	wire [11-1:0] node1547;
	wire [11-1:0] node1550;
	wire [11-1:0] node1551;
	wire [11-1:0] node1552;
	wire [11-1:0] node1555;
	wire [11-1:0] node1558;
	wire [11-1:0] node1561;
	wire [11-1:0] node1562;
	wire [11-1:0] node1563;
	wire [11-1:0] node1564;
	wire [11-1:0] node1567;
	wire [11-1:0] node1569;
	wire [11-1:0] node1572;
	wire [11-1:0] node1573;
	wire [11-1:0] node1576;
	wire [11-1:0] node1579;
	wire [11-1:0] node1580;
	wire [11-1:0] node1581;
	wire [11-1:0] node1582;
	wire [11-1:0] node1585;
	wire [11-1:0] node1588;
	wire [11-1:0] node1589;
	wire [11-1:0] node1592;
	wire [11-1:0] node1595;
	wire [11-1:0] node1596;
	wire [11-1:0] node1597;
	wire [11-1:0] node1601;
	wire [11-1:0] node1603;
	wire [11-1:0] node1606;
	wire [11-1:0] node1607;
	wire [11-1:0] node1608;
	wire [11-1:0] node1609;
	wire [11-1:0] node1610;
	wire [11-1:0] node1613;
	wire [11-1:0] node1616;
	wire [11-1:0] node1617;
	wire [11-1:0] node1618;
	wire [11-1:0] node1622;
	wire [11-1:0] node1623;
	wire [11-1:0] node1626;
	wire [11-1:0] node1629;
	wire [11-1:0] node1630;
	wire [11-1:0] node1631;
	wire [11-1:0] node1633;
	wire [11-1:0] node1636;
	wire [11-1:0] node1637;
	wire [11-1:0] node1641;
	wire [11-1:0] node1642;
	wire [11-1:0] node1645;
	wire [11-1:0] node1646;
	wire [11-1:0] node1650;
	wire [11-1:0] node1651;
	wire [11-1:0] node1652;
	wire [11-1:0] node1653;
	wire [11-1:0] node1654;
	wire [11-1:0] node1657;
	wire [11-1:0] node1660;
	wire [11-1:0] node1661;
	wire [11-1:0] node1664;
	wire [11-1:0] node1667;
	wire [11-1:0] node1669;
	wire [11-1:0] node1672;
	wire [11-1:0] node1673;
	wire [11-1:0] node1674;
	wire [11-1:0] node1677;
	wire [11-1:0] node1678;
	wire [11-1:0] node1681;
	wire [11-1:0] node1684;
	wire [11-1:0] node1685;
	wire [11-1:0] node1686;
	wire [11-1:0] node1689;
	wire [11-1:0] node1692;
	wire [11-1:0] node1693;
	wire [11-1:0] node1696;
	wire [11-1:0] node1699;
	wire [11-1:0] node1700;
	wire [11-1:0] node1701;
	wire [11-1:0] node1702;
	wire [11-1:0] node1703;
	wire [11-1:0] node1704;
	wire [11-1:0] node1705;
	wire [11-1:0] node1708;
	wire [11-1:0] node1711;
	wire [11-1:0] node1714;
	wire [11-1:0] node1715;
	wire [11-1:0] node1716;
	wire [11-1:0] node1719;
	wire [11-1:0] node1722;
	wire [11-1:0] node1724;
	wire [11-1:0] node1727;
	wire [11-1:0] node1728;
	wire [11-1:0] node1729;
	wire [11-1:0] node1730;
	wire [11-1:0] node1734;
	wire [11-1:0] node1737;
	wire [11-1:0] node1738;
	wire [11-1:0] node1741;
	wire [11-1:0] node1742;
	wire [11-1:0] node1745;
	wire [11-1:0] node1748;
	wire [11-1:0] node1749;
	wire [11-1:0] node1750;
	wire [11-1:0] node1751;
	wire [11-1:0] node1753;
	wire [11-1:0] node1756;
	wire [11-1:0] node1759;
	wire [11-1:0] node1760;
	wire [11-1:0] node1761;
	wire [11-1:0] node1764;
	wire [11-1:0] node1767;
	wire [11-1:0] node1768;
	wire [11-1:0] node1772;
	wire [11-1:0] node1773;
	wire [11-1:0] node1774;
	wire [11-1:0] node1775;
	wire [11-1:0] node1778;
	wire [11-1:0] node1781;
	wire [11-1:0] node1782;
	wire [11-1:0] node1786;
	wire [11-1:0] node1787;
	wire [11-1:0] node1791;
	wire [11-1:0] node1792;
	wire [11-1:0] node1793;
	wire [11-1:0] node1794;
	wire [11-1:0] node1795;
	wire [11-1:0] node1796;
	wire [11-1:0] node1800;
	wire [11-1:0] node1801;
	wire [11-1:0] node1804;
	wire [11-1:0] node1807;
	wire [11-1:0] node1808;
	wire [11-1:0] node1811;
	wire [11-1:0] node1814;
	wire [11-1:0] node1815;
	wire [11-1:0] node1816;
	wire [11-1:0] node1817;
	wire [11-1:0] node1820;
	wire [11-1:0] node1823;
	wire [11-1:0] node1826;
	wire [11-1:0] node1827;
	wire [11-1:0] node1829;
	wire [11-1:0] node1832;
	wire [11-1:0] node1833;
	wire [11-1:0] node1836;
	wire [11-1:0] node1839;
	wire [11-1:0] node1840;
	wire [11-1:0] node1841;
	wire [11-1:0] node1842;
	wire [11-1:0] node1843;
	wire [11-1:0] node1846;
	wire [11-1:0] node1849;
	wire [11-1:0] node1850;
	wire [11-1:0] node1853;
	wire [11-1:0] node1856;
	wire [11-1:0] node1857;
	wire [11-1:0] node1858;
	wire [11-1:0] node1861;
	wire [11-1:0] node1864;
	wire [11-1:0] node1865;
	wire [11-1:0] node1868;
	wire [11-1:0] node1871;
	wire [11-1:0] node1872;
	wire [11-1:0] node1873;
	wire [11-1:0] node1874;
	wire [11-1:0] node1878;
	wire [11-1:0] node1879;
	wire [11-1:0] node1882;
	wire [11-1:0] node1885;
	wire [11-1:0] node1886;
	wire [11-1:0] node1890;
	wire [11-1:0] node1891;
	wire [11-1:0] node1892;
	wire [11-1:0] node1893;
	wire [11-1:0] node1894;
	wire [11-1:0] node1895;
	wire [11-1:0] node1896;
	wire [11-1:0] node1898;
	wire [11-1:0] node1901;
	wire [11-1:0] node1904;
	wire [11-1:0] node1905;
	wire [11-1:0] node1906;
	wire [11-1:0] node1909;
	wire [11-1:0] node1912;
	wire [11-1:0] node1915;
	wire [11-1:0] node1916;
	wire [11-1:0] node1917;
	wire [11-1:0] node1918;
	wire [11-1:0] node1923;
	wire [11-1:0] node1924;
	wire [11-1:0] node1925;
	wire [11-1:0] node1929;
	wire [11-1:0] node1931;
	wire [11-1:0] node1934;
	wire [11-1:0] node1935;
	wire [11-1:0] node1936;
	wire [11-1:0] node1937;
	wire [11-1:0] node1939;
	wire [11-1:0] node1942;
	wire [11-1:0] node1945;
	wire [11-1:0] node1946;
	wire [11-1:0] node1947;
	wire [11-1:0] node1951;
	wire [11-1:0] node1952;
	wire [11-1:0] node1956;
	wire [11-1:0] node1957;
	wire [11-1:0] node1958;
	wire [11-1:0] node1959;
	wire [11-1:0] node1963;
	wire [11-1:0] node1966;
	wire [11-1:0] node1967;
	wire [11-1:0] node1970;
	wire [11-1:0] node1972;
	wire [11-1:0] node1975;
	wire [11-1:0] node1976;
	wire [11-1:0] node1977;
	wire [11-1:0] node1978;
	wire [11-1:0] node1979;
	wire [11-1:0] node1980;
	wire [11-1:0] node1983;
	wire [11-1:0] node1986;
	wire [11-1:0] node1989;
	wire [11-1:0] node1990;
	wire [11-1:0] node1991;
	wire [11-1:0] node1994;
	wire [11-1:0] node1997;
	wire [11-1:0] node1998;
	wire [11-1:0] node2001;
	wire [11-1:0] node2004;
	wire [11-1:0] node2005;
	wire [11-1:0] node2006;
	wire [11-1:0] node2007;
	wire [11-1:0] node2010;
	wire [11-1:0] node2013;
	wire [11-1:0] node2014;
	wire [11-1:0] node2018;
	wire [11-1:0] node2019;
	wire [11-1:0] node2022;
	wire [11-1:0] node2023;
	wire [11-1:0] node2027;
	wire [11-1:0] node2028;
	wire [11-1:0] node2029;
	wire [11-1:0] node2030;
	wire [11-1:0] node2033;
	wire [11-1:0] node2036;
	wire [11-1:0] node2037;
	wire [11-1:0] node2039;
	wire [11-1:0] node2042;
	wire [11-1:0] node2043;
	wire [11-1:0] node2047;
	wire [11-1:0] node2048;
	wire [11-1:0] node2049;
	wire [11-1:0] node2052;
	wire [11-1:0] node2053;
	wire [11-1:0] node2056;
	wire [11-1:0] node2059;
	wire [11-1:0] node2060;
	wire [11-1:0] node2061;
	wire [11-1:0] node2065;
	wire [11-1:0] node2066;
	wire [11-1:0] node2069;
	wire [11-1:0] node2072;
	wire [11-1:0] node2073;
	wire [11-1:0] node2074;
	wire [11-1:0] node2075;
	wire [11-1:0] node2076;
	wire [11-1:0] node2077;
	wire [11-1:0] node2080;
	wire [11-1:0] node2082;
	wire [11-1:0] node2085;
	wire [11-1:0] node2086;
	wire [11-1:0] node2087;
	wire [11-1:0] node2091;
	wire [11-1:0] node2092;
	wire [11-1:0] node2096;
	wire [11-1:0] node2097;
	wire [11-1:0] node2098;
	wire [11-1:0] node2099;
	wire [11-1:0] node2103;
	wire [11-1:0] node2104;
	wire [11-1:0] node2107;
	wire [11-1:0] node2110;
	wire [11-1:0] node2111;
	wire [11-1:0] node2113;
	wire [11-1:0] node2116;
	wire [11-1:0] node2117;
	wire [11-1:0] node2120;
	wire [11-1:0] node2123;
	wire [11-1:0] node2124;
	wire [11-1:0] node2125;
	wire [11-1:0] node2126;
	wire [11-1:0] node2128;
	wire [11-1:0] node2131;
	wire [11-1:0] node2132;
	wire [11-1:0] node2135;
	wire [11-1:0] node2138;
	wire [11-1:0] node2139;
	wire [11-1:0] node2140;
	wire [11-1:0] node2143;
	wire [11-1:0] node2146;
	wire [11-1:0] node2148;
	wire [11-1:0] node2151;
	wire [11-1:0] node2152;
	wire [11-1:0] node2153;
	wire [11-1:0] node2154;
	wire [11-1:0] node2157;
	wire [11-1:0] node2160;
	wire [11-1:0] node2162;
	wire [11-1:0] node2165;
	wire [11-1:0] node2166;
	wire [11-1:0] node2169;
	wire [11-1:0] node2171;
	wire [11-1:0] node2174;
	wire [11-1:0] node2175;
	wire [11-1:0] node2176;
	wire [11-1:0] node2177;
	wire [11-1:0] node2179;
	wire [11-1:0] node2180;
	wire [11-1:0] node2183;
	wire [11-1:0] node2186;
	wire [11-1:0] node2187;
	wire [11-1:0] node2190;
	wire [11-1:0] node2191;
	wire [11-1:0] node2194;
	wire [11-1:0] node2197;
	wire [11-1:0] node2198;
	wire [11-1:0] node2199;
	wire [11-1:0] node2202;
	wire [11-1:0] node2204;
	wire [11-1:0] node2207;
	wire [11-1:0] node2208;
	wire [11-1:0] node2209;
	wire [11-1:0] node2213;
	wire [11-1:0] node2214;
	wire [11-1:0] node2218;
	wire [11-1:0] node2219;
	wire [11-1:0] node2220;
	wire [11-1:0] node2222;
	wire [11-1:0] node2223;
	wire [11-1:0] node2226;
	wire [11-1:0] node2229;
	wire [11-1:0] node2230;
	wire [11-1:0] node2231;
	wire [11-1:0] node2234;
	wire [11-1:0] node2237;
	wire [11-1:0] node2240;
	wire [11-1:0] node2241;
	wire [11-1:0] node2242;
	wire [11-1:0] node2245;
	wire [11-1:0] node2246;
	wire [11-1:0] node2249;
	wire [11-1:0] node2252;
	wire [11-1:0] node2255;
	wire [11-1:0] node2256;
	wire [11-1:0] node2257;
	wire [11-1:0] node2258;
	wire [11-1:0] node2259;
	wire [11-1:0] node2260;
	wire [11-1:0] node2261;
	wire [11-1:0] node2262;
	wire [11-1:0] node2263;
	wire [11-1:0] node2266;
	wire [11-1:0] node2269;
	wire [11-1:0] node2270;
	wire [11-1:0] node2274;
	wire [11-1:0] node2275;
	wire [11-1:0] node2276;
	wire [11-1:0] node2280;
	wire [11-1:0] node2282;
	wire [11-1:0] node2285;
	wire [11-1:0] node2286;
	wire [11-1:0] node2288;
	wire [11-1:0] node2289;
	wire [11-1:0] node2292;
	wire [11-1:0] node2295;
	wire [11-1:0] node2296;
	wire [11-1:0] node2299;
	wire [11-1:0] node2300;
	wire [11-1:0] node2303;
	wire [11-1:0] node2306;
	wire [11-1:0] node2307;
	wire [11-1:0] node2308;
	wire [11-1:0] node2309;
	wire [11-1:0] node2311;
	wire [11-1:0] node2314;
	wire [11-1:0] node2317;
	wire [11-1:0] node2318;
	wire [11-1:0] node2320;
	wire [11-1:0] node2323;
	wire [11-1:0] node2324;
	wire [11-1:0] node2327;
	wire [11-1:0] node2330;
	wire [11-1:0] node2331;
	wire [11-1:0] node2332;
	wire [11-1:0] node2335;
	wire [11-1:0] node2336;
	wire [11-1:0] node2339;
	wire [11-1:0] node2342;
	wire [11-1:0] node2343;
	wire [11-1:0] node2344;
	wire [11-1:0] node2347;
	wire [11-1:0] node2350;
	wire [11-1:0] node2351;
	wire [11-1:0] node2355;
	wire [11-1:0] node2356;
	wire [11-1:0] node2357;
	wire [11-1:0] node2358;
	wire [11-1:0] node2359;
	wire [11-1:0] node2360;
	wire [11-1:0] node2363;
	wire [11-1:0] node2367;
	wire [11-1:0] node2368;
	wire [11-1:0] node2369;
	wire [11-1:0] node2373;
	wire [11-1:0] node2374;
	wire [11-1:0] node2377;
	wire [11-1:0] node2380;
	wire [11-1:0] node2381;
	wire [11-1:0] node2382;
	wire [11-1:0] node2383;
	wire [11-1:0] node2386;
	wire [11-1:0] node2389;
	wire [11-1:0] node2391;
	wire [11-1:0] node2394;
	wire [11-1:0] node2395;
	wire [11-1:0] node2396;
	wire [11-1:0] node2399;
	wire [11-1:0] node2402;
	wire [11-1:0] node2403;
	wire [11-1:0] node2406;
	wire [11-1:0] node2409;
	wire [11-1:0] node2410;
	wire [11-1:0] node2411;
	wire [11-1:0] node2412;
	wire [11-1:0] node2413;
	wire [11-1:0] node2417;
	wire [11-1:0] node2418;
	wire [11-1:0] node2422;
	wire [11-1:0] node2423;
	wire [11-1:0] node2424;
	wire [11-1:0] node2427;
	wire [11-1:0] node2430;
	wire [11-1:0] node2431;
	wire [11-1:0] node2434;
	wire [11-1:0] node2437;
	wire [11-1:0] node2438;
	wire [11-1:0] node2439;
	wire [11-1:0] node2440;
	wire [11-1:0] node2444;
	wire [11-1:0] node2445;
	wire [11-1:0] node2448;
	wire [11-1:0] node2451;
	wire [11-1:0] node2452;
	wire [11-1:0] node2454;
	wire [11-1:0] node2457;
	wire [11-1:0] node2459;
	wire [11-1:0] node2462;
	wire [11-1:0] node2463;
	wire [11-1:0] node2464;
	wire [11-1:0] node2465;
	wire [11-1:0] node2466;
	wire [11-1:0] node2467;
	wire [11-1:0] node2468;
	wire [11-1:0] node2472;
	wire [11-1:0] node2474;
	wire [11-1:0] node2477;
	wire [11-1:0] node2478;
	wire [11-1:0] node2479;
	wire [11-1:0] node2483;
	wire [11-1:0] node2486;
	wire [11-1:0] node2487;
	wire [11-1:0] node2488;
	wire [11-1:0] node2489;
	wire [11-1:0] node2492;
	wire [11-1:0] node2495;
	wire [11-1:0] node2497;
	wire [11-1:0] node2500;
	wire [11-1:0] node2501;
	wire [11-1:0] node2502;
	wire [11-1:0] node2506;
	wire [11-1:0] node2507;
	wire [11-1:0] node2510;
	wire [11-1:0] node2513;
	wire [11-1:0] node2514;
	wire [11-1:0] node2515;
	wire [11-1:0] node2517;
	wire [11-1:0] node2520;
	wire [11-1:0] node2521;
	wire [11-1:0] node2522;
	wire [11-1:0] node2526;
	wire [11-1:0] node2527;
	wire [11-1:0] node2530;
	wire [11-1:0] node2533;
	wire [11-1:0] node2534;
	wire [11-1:0] node2535;
	wire [11-1:0] node2536;
	wire [11-1:0] node2540;
	wire [11-1:0] node2543;
	wire [11-1:0] node2544;
	wire [11-1:0] node2545;
	wire [11-1:0] node2549;
	wire [11-1:0] node2550;
	wire [11-1:0] node2553;
	wire [11-1:0] node2556;
	wire [11-1:0] node2557;
	wire [11-1:0] node2558;
	wire [11-1:0] node2559;
	wire [11-1:0] node2560;
	wire [11-1:0] node2561;
	wire [11-1:0] node2564;
	wire [11-1:0] node2567;
	wire [11-1:0] node2569;
	wire [11-1:0] node2572;
	wire [11-1:0] node2573;
	wire [11-1:0] node2574;
	wire [11-1:0] node2577;
	wire [11-1:0] node2580;
	wire [11-1:0] node2582;
	wire [11-1:0] node2585;
	wire [11-1:0] node2586;
	wire [11-1:0] node2587;
	wire [11-1:0] node2589;
	wire [11-1:0] node2592;
	wire [11-1:0] node2593;
	wire [11-1:0] node2596;
	wire [11-1:0] node2599;
	wire [11-1:0] node2600;
	wire [11-1:0] node2603;
	wire [11-1:0] node2604;
	wire [11-1:0] node2608;
	wire [11-1:0] node2609;
	wire [11-1:0] node2610;
	wire [11-1:0] node2611;
	wire [11-1:0] node2614;
	wire [11-1:0] node2617;
	wire [11-1:0] node2618;
	wire [11-1:0] node2620;
	wire [11-1:0] node2623;
	wire [11-1:0] node2625;
	wire [11-1:0] node2628;
	wire [11-1:0] node2629;
	wire [11-1:0] node2630;
	wire [11-1:0] node2631;
	wire [11-1:0] node2634;
	wire [11-1:0] node2637;
	wire [11-1:0] node2640;
	wire [11-1:0] node2641;
	wire [11-1:0] node2642;
	wire [11-1:0] node2645;
	wire [11-1:0] node2648;
	wire [11-1:0] node2651;
	wire [11-1:0] node2652;
	wire [11-1:0] node2653;
	wire [11-1:0] node2654;
	wire [11-1:0] node2655;
	wire [11-1:0] node2656;
	wire [11-1:0] node2657;
	wire [11-1:0] node2658;
	wire [11-1:0] node2662;
	wire [11-1:0] node2663;
	wire [11-1:0] node2666;
	wire [11-1:0] node2669;
	wire [11-1:0] node2670;
	wire [11-1:0] node2671;
	wire [11-1:0] node2675;
	wire [11-1:0] node2678;
	wire [11-1:0] node2679;
	wire [11-1:0] node2680;
	wire [11-1:0] node2681;
	wire [11-1:0] node2685;
	wire [11-1:0] node2687;
	wire [11-1:0] node2690;
	wire [11-1:0] node2691;
	wire [11-1:0] node2694;
	wire [11-1:0] node2695;
	wire [11-1:0] node2699;
	wire [11-1:0] node2700;
	wire [11-1:0] node2701;
	wire [11-1:0] node2702;
	wire [11-1:0] node2703;
	wire [11-1:0] node2706;
	wire [11-1:0] node2709;
	wire [11-1:0] node2710;
	wire [11-1:0] node2714;
	wire [11-1:0] node2715;
	wire [11-1:0] node2716;
	wire [11-1:0] node2719;
	wire [11-1:0] node2722;
	wire [11-1:0] node2723;
	wire [11-1:0] node2726;
	wire [11-1:0] node2729;
	wire [11-1:0] node2730;
	wire [11-1:0] node2731;
	wire [11-1:0] node2732;
	wire [11-1:0] node2735;
	wire [11-1:0] node2738;
	wire [11-1:0] node2741;
	wire [11-1:0] node2742;
	wire [11-1:0] node2744;
	wire [11-1:0] node2747;
	wire [11-1:0] node2748;
	wire [11-1:0] node2751;
	wire [11-1:0] node2754;
	wire [11-1:0] node2755;
	wire [11-1:0] node2756;
	wire [11-1:0] node2757;
	wire [11-1:0] node2758;
	wire [11-1:0] node2759;
	wire [11-1:0] node2762;
	wire [11-1:0] node2765;
	wire [11-1:0] node2768;
	wire [11-1:0] node2769;
	wire [11-1:0] node2771;
	wire [11-1:0] node2774;
	wire [11-1:0] node2775;
	wire [11-1:0] node2778;
	wire [11-1:0] node2781;
	wire [11-1:0] node2782;
	wire [11-1:0] node2783;
	wire [11-1:0] node2786;
	wire [11-1:0] node2787;
	wire [11-1:0] node2791;
	wire [11-1:0] node2793;
	wire [11-1:0] node2794;
	wire [11-1:0] node2797;
	wire [11-1:0] node2800;
	wire [11-1:0] node2801;
	wire [11-1:0] node2802;
	wire [11-1:0] node2803;
	wire [11-1:0] node2804;
	wire [11-1:0] node2807;
	wire [11-1:0] node2810;
	wire [11-1:0] node2812;
	wire [11-1:0] node2815;
	wire [11-1:0] node2816;
	wire [11-1:0] node2817;
	wire [11-1:0] node2820;
	wire [11-1:0] node2824;
	wire [11-1:0] node2825;
	wire [11-1:0] node2827;
	wire [11-1:0] node2830;
	wire [11-1:0] node2831;
	wire [11-1:0] node2833;
	wire [11-1:0] node2836;
	wire [11-1:0] node2839;
	wire [11-1:0] node2840;
	wire [11-1:0] node2841;
	wire [11-1:0] node2842;
	wire [11-1:0] node2843;
	wire [11-1:0] node2844;
	wire [11-1:0] node2846;
	wire [11-1:0] node2849;
	wire [11-1:0] node2850;
	wire [11-1:0] node2853;
	wire [11-1:0] node2856;
	wire [11-1:0] node2857;
	wire [11-1:0] node2859;
	wire [11-1:0] node2862;
	wire [11-1:0] node2865;
	wire [11-1:0] node2866;
	wire [11-1:0] node2867;
	wire [11-1:0] node2868;
	wire [11-1:0] node2872;
	wire [11-1:0] node2873;
	wire [11-1:0] node2877;
	wire [11-1:0] node2878;
	wire [11-1:0] node2879;
	wire [11-1:0] node2882;
	wire [11-1:0] node2885;
	wire [11-1:0] node2887;
	wire [11-1:0] node2890;
	wire [11-1:0] node2891;
	wire [11-1:0] node2892;
	wire [11-1:0] node2893;
	wire [11-1:0] node2896;
	wire [11-1:0] node2897;
	wire [11-1:0] node2901;
	wire [11-1:0] node2902;
	wire [11-1:0] node2903;
	wire [11-1:0] node2906;
	wire [11-1:0] node2909;
	wire [11-1:0] node2912;
	wire [11-1:0] node2913;
	wire [11-1:0] node2914;
	wire [11-1:0] node2915;
	wire [11-1:0] node2918;
	wire [11-1:0] node2921;
	wire [11-1:0] node2924;
	wire [11-1:0] node2925;
	wire [11-1:0] node2928;
	wire [11-1:0] node2929;
	wire [11-1:0] node2932;
	wire [11-1:0] node2935;
	wire [11-1:0] node2936;
	wire [11-1:0] node2937;
	wire [11-1:0] node2938;
	wire [11-1:0] node2939;
	wire [11-1:0] node2940;
	wire [11-1:0] node2943;
	wire [11-1:0] node2946;
	wire [11-1:0] node2949;
	wire [11-1:0] node2950;
	wire [11-1:0] node2951;
	wire [11-1:0] node2954;
	wire [11-1:0] node2957;
	wire [11-1:0] node2959;
	wire [11-1:0] node2962;
	wire [11-1:0] node2963;
	wire [11-1:0] node2964;
	wire [11-1:0] node2967;
	wire [11-1:0] node2968;
	wire [11-1:0] node2971;
	wire [11-1:0] node2974;
	wire [11-1:0] node2976;
	wire [11-1:0] node2978;
	wire [11-1:0] node2981;
	wire [11-1:0] node2982;
	wire [11-1:0] node2983;
	wire [11-1:0] node2984;
	wire [11-1:0] node2985;
	wire [11-1:0] node2988;
	wire [11-1:0] node2991;
	wire [11-1:0] node2992;
	wire [11-1:0] node2995;
	wire [11-1:0] node2998;
	wire [11-1:0] node2999;
	wire [11-1:0] node3001;
	wire [11-1:0] node3004;
	wire [11-1:0] node3007;
	wire [11-1:0] node3008;
	wire [11-1:0] node3009;
	wire [11-1:0] node3010;
	wire [11-1:0] node3013;
	wire [11-1:0] node3016;
	wire [11-1:0] node3018;
	wire [11-1:0] node3021;
	wire [11-1:0] node3022;
	wire [11-1:0] node3023;
	wire [11-1:0] node3027;
	wire [11-1:0] node3028;
	wire [11-1:0] node3032;
	wire [11-1:0] node3033;
	wire [11-1:0] node3034;
	wire [11-1:0] node3035;
	wire [11-1:0] node3036;
	wire [11-1:0] node3037;
	wire [11-1:0] node3038;
	wire [11-1:0] node3039;
	wire [11-1:0] node3040;
	wire [11-1:0] node3041;
	wire [11-1:0] node3044;
	wire [11-1:0] node3045;
	wire [11-1:0] node3048;
	wire [11-1:0] node3051;
	wire [11-1:0] node3052;
	wire [11-1:0] node3053;
	wire [11-1:0] node3056;
	wire [11-1:0] node3059;
	wire [11-1:0] node3060;
	wire [11-1:0] node3063;
	wire [11-1:0] node3066;
	wire [11-1:0] node3067;
	wire [11-1:0] node3068;
	wire [11-1:0] node3069;
	wire [11-1:0] node3073;
	wire [11-1:0] node3074;
	wire [11-1:0] node3078;
	wire [11-1:0] node3079;
	wire [11-1:0] node3080;
	wire [11-1:0] node3083;
	wire [11-1:0] node3086;
	wire [11-1:0] node3089;
	wire [11-1:0] node3090;
	wire [11-1:0] node3091;
	wire [11-1:0] node3092;
	wire [11-1:0] node3093;
	wire [11-1:0] node3097;
	wire [11-1:0] node3098;
	wire [11-1:0] node3102;
	wire [11-1:0] node3103;
	wire [11-1:0] node3104;
	wire [11-1:0] node3107;
	wire [11-1:0] node3110;
	wire [11-1:0] node3113;
	wire [11-1:0] node3114;
	wire [11-1:0] node3115;
	wire [11-1:0] node3116;
	wire [11-1:0] node3120;
	wire [11-1:0] node3121;
	wire [11-1:0] node3124;
	wire [11-1:0] node3127;
	wire [11-1:0] node3128;
	wire [11-1:0] node3130;
	wire [11-1:0] node3133;
	wire [11-1:0] node3134;
	wire [11-1:0] node3138;
	wire [11-1:0] node3139;
	wire [11-1:0] node3140;
	wire [11-1:0] node3141;
	wire [11-1:0] node3142;
	wire [11-1:0] node3143;
	wire [11-1:0] node3147;
	wire [11-1:0] node3148;
	wire [11-1:0] node3151;
	wire [11-1:0] node3154;
	wire [11-1:0] node3155;
	wire [11-1:0] node3156;
	wire [11-1:0] node3159;
	wire [11-1:0] node3162;
	wire [11-1:0] node3163;
	wire [11-1:0] node3167;
	wire [11-1:0] node3168;
	wire [11-1:0] node3169;
	wire [11-1:0] node3171;
	wire [11-1:0] node3174;
	wire [11-1:0] node3175;
	wire [11-1:0] node3179;
	wire [11-1:0] node3180;
	wire [11-1:0] node3181;
	wire [11-1:0] node3185;
	wire [11-1:0] node3186;
	wire [11-1:0] node3189;
	wire [11-1:0] node3192;
	wire [11-1:0] node3193;
	wire [11-1:0] node3194;
	wire [11-1:0] node3195;
	wire [11-1:0] node3196;
	wire [11-1:0] node3200;
	wire [11-1:0] node3201;
	wire [11-1:0] node3205;
	wire [11-1:0] node3207;
	wire [11-1:0] node3208;
	wire [11-1:0] node3211;
	wire [11-1:0] node3214;
	wire [11-1:0] node3215;
	wire [11-1:0] node3216;
	wire [11-1:0] node3219;
	wire [11-1:0] node3221;
	wire [11-1:0] node3224;
	wire [11-1:0] node3225;
	wire [11-1:0] node3228;
	wire [11-1:0] node3229;
	wire [11-1:0] node3233;
	wire [11-1:0] node3234;
	wire [11-1:0] node3235;
	wire [11-1:0] node3236;
	wire [11-1:0] node3237;
	wire [11-1:0] node3238;
	wire [11-1:0] node3241;
	wire [11-1:0] node3244;
	wire [11-1:0] node3245;
	wire [11-1:0] node3246;
	wire [11-1:0] node3250;
	wire [11-1:0] node3252;
	wire [11-1:0] node3255;
	wire [11-1:0] node3256;
	wire [11-1:0] node3257;
	wire [11-1:0] node3258;
	wire [11-1:0] node3261;
	wire [11-1:0] node3264;
	wire [11-1:0] node3266;
	wire [11-1:0] node3269;
	wire [11-1:0] node3270;
	wire [11-1:0] node3271;
	wire [11-1:0] node3274;
	wire [11-1:0] node3277;
	wire [11-1:0] node3280;
	wire [11-1:0] node3281;
	wire [11-1:0] node3282;
	wire [11-1:0] node3284;
	wire [11-1:0] node3285;
	wire [11-1:0] node3288;
	wire [11-1:0] node3291;
	wire [11-1:0] node3292;
	wire [11-1:0] node3293;
	wire [11-1:0] node3296;
	wire [11-1:0] node3299;
	wire [11-1:0] node3300;
	wire [11-1:0] node3303;
	wire [11-1:0] node3306;
	wire [11-1:0] node3307;
	wire [11-1:0] node3308;
	wire [11-1:0] node3309;
	wire [11-1:0] node3313;
	wire [11-1:0] node3315;
	wire [11-1:0] node3318;
	wire [11-1:0] node3319;
	wire [11-1:0] node3322;
	wire [11-1:0] node3323;
	wire [11-1:0] node3327;
	wire [11-1:0] node3328;
	wire [11-1:0] node3329;
	wire [11-1:0] node3330;
	wire [11-1:0] node3331;
	wire [11-1:0] node3332;
	wire [11-1:0] node3335;
	wire [11-1:0] node3338;
	wire [11-1:0] node3341;
	wire [11-1:0] node3342;
	wire [11-1:0] node3343;
	wire [11-1:0] node3347;
	wire [11-1:0] node3350;
	wire [11-1:0] node3351;
	wire [11-1:0] node3352;
	wire [11-1:0] node3354;
	wire [11-1:0] node3357;
	wire [11-1:0] node3360;
	wire [11-1:0] node3361;
	wire [11-1:0] node3362;
	wire [11-1:0] node3365;
	wire [11-1:0] node3368;
	wire [11-1:0] node3370;
	wire [11-1:0] node3373;
	wire [11-1:0] node3374;
	wire [11-1:0] node3375;
	wire [11-1:0] node3376;
	wire [11-1:0] node3377;
	wire [11-1:0] node3381;
	wire [11-1:0] node3382;
	wire [11-1:0] node3386;
	wire [11-1:0] node3387;
	wire [11-1:0] node3388;
	wire [11-1:0] node3392;
	wire [11-1:0] node3395;
	wire [11-1:0] node3396;
	wire [11-1:0] node3397;
	wire [11-1:0] node3400;
	wire [11-1:0] node3403;
	wire [11-1:0] node3404;
	wire [11-1:0] node3406;
	wire [11-1:0] node3410;
	wire [11-1:0] node3411;
	wire [11-1:0] node3412;
	wire [11-1:0] node3413;
	wire [11-1:0] node3414;
	wire [11-1:0] node3415;
	wire [11-1:0] node3416;
	wire [11-1:0] node3417;
	wire [11-1:0] node3421;
	wire [11-1:0] node3422;
	wire [11-1:0] node3425;
	wire [11-1:0] node3428;
	wire [11-1:0] node3429;
	wire [11-1:0] node3431;
	wire [11-1:0] node3434;
	wire [11-1:0] node3437;
	wire [11-1:0] node3438;
	wire [11-1:0] node3439;
	wire [11-1:0] node3441;
	wire [11-1:0] node3444;
	wire [11-1:0] node3445;
	wire [11-1:0] node3448;
	wire [11-1:0] node3451;
	wire [11-1:0] node3452;
	wire [11-1:0] node3455;
	wire [11-1:0] node3457;
	wire [11-1:0] node3460;
	wire [11-1:0] node3461;
	wire [11-1:0] node3462;
	wire [11-1:0] node3463;
	wire [11-1:0] node3464;
	wire [11-1:0] node3468;
	wire [11-1:0] node3469;
	wire [11-1:0] node3472;
	wire [11-1:0] node3475;
	wire [11-1:0] node3476;
	wire [11-1:0] node3479;
	wire [11-1:0] node3480;
	wire [11-1:0] node3484;
	wire [11-1:0] node3485;
	wire [11-1:0] node3486;
	wire [11-1:0] node3489;
	wire [11-1:0] node3492;
	wire [11-1:0] node3494;
	wire [11-1:0] node3495;
	wire [11-1:0] node3499;
	wire [11-1:0] node3500;
	wire [11-1:0] node3501;
	wire [11-1:0] node3502;
	wire [11-1:0] node3503;
	wire [11-1:0] node3506;
	wire [11-1:0] node3507;
	wire [11-1:0] node3511;
	wire [11-1:0] node3512;
	wire [11-1:0] node3514;
	wire [11-1:0] node3517;
	wire [11-1:0] node3519;
	wire [11-1:0] node3522;
	wire [11-1:0] node3523;
	wire [11-1:0] node3524;
	wire [11-1:0] node3526;
	wire [11-1:0] node3529;
	wire [11-1:0] node3532;
	wire [11-1:0] node3533;
	wire [11-1:0] node3534;
	wire [11-1:0] node3538;
	wire [11-1:0] node3539;
	wire [11-1:0] node3542;
	wire [11-1:0] node3545;
	wire [11-1:0] node3546;
	wire [11-1:0] node3547;
	wire [11-1:0] node3548;
	wire [11-1:0] node3551;
	wire [11-1:0] node3552;
	wire [11-1:0] node3555;
	wire [11-1:0] node3558;
	wire [11-1:0] node3559;
	wire [11-1:0] node3561;
	wire [11-1:0] node3564;
	wire [11-1:0] node3567;
	wire [11-1:0] node3568;
	wire [11-1:0] node3569;
	wire [11-1:0] node3572;
	wire [11-1:0] node3574;
	wire [11-1:0] node3577;
	wire [11-1:0] node3578;
	wire [11-1:0] node3579;
	wire [11-1:0] node3582;
	wire [11-1:0] node3585;
	wire [11-1:0] node3588;
	wire [11-1:0] node3589;
	wire [11-1:0] node3590;
	wire [11-1:0] node3591;
	wire [11-1:0] node3592;
	wire [11-1:0] node3593;
	wire [11-1:0] node3594;
	wire [11-1:0] node3597;
	wire [11-1:0] node3600;
	wire [11-1:0] node3601;
	wire [11-1:0] node3605;
	wire [11-1:0] node3606;
	wire [11-1:0] node3608;
	wire [11-1:0] node3611;
	wire [11-1:0] node3613;
	wire [11-1:0] node3616;
	wire [11-1:0] node3617;
	wire [11-1:0] node3618;
	wire [11-1:0] node3619;
	wire [11-1:0] node3623;
	wire [11-1:0] node3624;
	wire [11-1:0] node3628;
	wire [11-1:0] node3629;
	wire [11-1:0] node3630;
	wire [11-1:0] node3634;
	wire [11-1:0] node3637;
	wire [11-1:0] node3638;
	wire [11-1:0] node3639;
	wire [11-1:0] node3640;
	wire [11-1:0] node3641;
	wire [11-1:0] node3644;
	wire [11-1:0] node3647;
	wire [11-1:0] node3650;
	wire [11-1:0] node3651;
	wire [11-1:0] node3652;
	wire [11-1:0] node3656;
	wire [11-1:0] node3657;
	wire [11-1:0] node3660;
	wire [11-1:0] node3663;
	wire [11-1:0] node3664;
	wire [11-1:0] node3665;
	wire [11-1:0] node3666;
	wire [11-1:0] node3669;
	wire [11-1:0] node3672;
	wire [11-1:0] node3673;
	wire [11-1:0] node3676;
	wire [11-1:0] node3679;
	wire [11-1:0] node3680;
	wire [11-1:0] node3682;
	wire [11-1:0] node3685;
	wire [11-1:0] node3686;
	wire [11-1:0] node3690;
	wire [11-1:0] node3691;
	wire [11-1:0] node3692;
	wire [11-1:0] node3693;
	wire [11-1:0] node3694;
	wire [11-1:0] node3698;
	wire [11-1:0] node3699;
	wire [11-1:0] node3700;
	wire [11-1:0] node3704;
	wire [11-1:0] node3705;
	wire [11-1:0] node3708;
	wire [11-1:0] node3711;
	wire [11-1:0] node3712;
	wire [11-1:0] node3713;
	wire [11-1:0] node3714;
	wire [11-1:0] node3717;
	wire [11-1:0] node3721;
	wire [11-1:0] node3722;
	wire [11-1:0] node3723;
	wire [11-1:0] node3726;
	wire [11-1:0] node3729;
	wire [11-1:0] node3730;
	wire [11-1:0] node3733;
	wire [11-1:0] node3736;
	wire [11-1:0] node3737;
	wire [11-1:0] node3738;
	wire [11-1:0] node3739;
	wire [11-1:0] node3740;
	wire [11-1:0] node3743;
	wire [11-1:0] node3746;
	wire [11-1:0] node3747;
	wire [11-1:0] node3751;
	wire [11-1:0] node3752;
	wire [11-1:0] node3753;
	wire [11-1:0] node3758;
	wire [11-1:0] node3759;
	wire [11-1:0] node3760;
	wire [11-1:0] node3763;
	wire [11-1:0] node3764;
	wire [11-1:0] node3767;
	wire [11-1:0] node3770;
	wire [11-1:0] node3771;
	wire [11-1:0] node3774;
	wire [11-1:0] node3775;
	wire [11-1:0] node3778;
	wire [11-1:0] node3781;
	wire [11-1:0] node3782;
	wire [11-1:0] node3783;
	wire [11-1:0] node3784;
	wire [11-1:0] node3785;
	wire [11-1:0] node3786;
	wire [11-1:0] node3787;
	wire [11-1:0] node3788;
	wire [11-1:0] node3789;
	wire [11-1:0] node3792;
	wire [11-1:0] node3795;
	wire [11-1:0] node3796;
	wire [11-1:0] node3800;
	wire [11-1:0] node3801;
	wire [11-1:0] node3802;
	wire [11-1:0] node3806;
	wire [11-1:0] node3809;
	wire [11-1:0] node3810;
	wire [11-1:0] node3811;
	wire [11-1:0] node3813;
	wire [11-1:0] node3816;
	wire [11-1:0] node3819;
	wire [11-1:0] node3820;
	wire [11-1:0] node3823;
	wire [11-1:0] node3824;
	wire [11-1:0] node3827;
	wire [11-1:0] node3830;
	wire [11-1:0] node3831;
	wire [11-1:0] node3832;
	wire [11-1:0] node3833;
	wire [11-1:0] node3834;
	wire [11-1:0] node3838;
	wire [11-1:0] node3839;
	wire [11-1:0] node3842;
	wire [11-1:0] node3845;
	wire [11-1:0] node3846;
	wire [11-1:0] node3847;
	wire [11-1:0] node3850;
	wire [11-1:0] node3853;
	wire [11-1:0] node3856;
	wire [11-1:0] node3857;
	wire [11-1:0] node3858;
	wire [11-1:0] node3859;
	wire [11-1:0] node3862;
	wire [11-1:0] node3865;
	wire [11-1:0] node3867;
	wire [11-1:0] node3870;
	wire [11-1:0] node3871;
	wire [11-1:0] node3874;
	wire [11-1:0] node3875;
	wire [11-1:0] node3878;
	wire [11-1:0] node3881;
	wire [11-1:0] node3882;
	wire [11-1:0] node3883;
	wire [11-1:0] node3884;
	wire [11-1:0] node3885;
	wire [11-1:0] node3886;
	wire [11-1:0] node3890;
	wire [11-1:0] node3891;
	wire [11-1:0] node3894;
	wire [11-1:0] node3897;
	wire [11-1:0] node3898;
	wire [11-1:0] node3899;
	wire [11-1:0] node3902;
	wire [11-1:0] node3905;
	wire [11-1:0] node3906;
	wire [11-1:0] node3909;
	wire [11-1:0] node3912;
	wire [11-1:0] node3913;
	wire [11-1:0] node3914;
	wire [11-1:0] node3915;
	wire [11-1:0] node3918;
	wire [11-1:0] node3921;
	wire [11-1:0] node3922;
	wire [11-1:0] node3926;
	wire [11-1:0] node3927;
	wire [11-1:0] node3930;
	wire [11-1:0] node3931;
	wire [11-1:0] node3934;
	wire [11-1:0] node3937;
	wire [11-1:0] node3938;
	wire [11-1:0] node3939;
	wire [11-1:0] node3940;
	wire [11-1:0] node3941;
	wire [11-1:0] node3944;
	wire [11-1:0] node3947;
	wire [11-1:0] node3948;
	wire [11-1:0] node3951;
	wire [11-1:0] node3954;
	wire [11-1:0] node3955;
	wire [11-1:0] node3956;
	wire [11-1:0] node3959;
	wire [11-1:0] node3962;
	wire [11-1:0] node3965;
	wire [11-1:0] node3966;
	wire [11-1:0] node3967;
	wire [11-1:0] node3968;
	wire [11-1:0] node3971;
	wire [11-1:0] node3974;
	wire [11-1:0] node3975;
	wire [11-1:0] node3979;
	wire [11-1:0] node3980;
	wire [11-1:0] node3983;
	wire [11-1:0] node3984;
	wire [11-1:0] node3988;
	wire [11-1:0] node3989;
	wire [11-1:0] node3990;
	wire [11-1:0] node3991;
	wire [11-1:0] node3992;
	wire [11-1:0] node3993;
	wire [11-1:0] node3996;
	wire [11-1:0] node3999;
	wire [11-1:0] node4000;
	wire [11-1:0] node4001;
	wire [11-1:0] node4004;
	wire [11-1:0] node4007;
	wire [11-1:0] node4010;
	wire [11-1:0] node4011;
	wire [11-1:0] node4012;
	wire [11-1:0] node4013;
	wire [11-1:0] node4016;
	wire [11-1:0] node4019;
	wire [11-1:0] node4020;
	wire [11-1:0] node4023;
	wire [11-1:0] node4026;
	wire [11-1:0] node4027;
	wire [11-1:0] node4029;
	wire [11-1:0] node4032;
	wire [11-1:0] node4034;
	wire [11-1:0] node4037;
	wire [11-1:0] node4038;
	wire [11-1:0] node4039;
	wire [11-1:0] node4040;
	wire [11-1:0] node4043;
	wire [11-1:0] node4044;
	wire [11-1:0] node4047;
	wire [11-1:0] node4050;
	wire [11-1:0] node4051;
	wire [11-1:0] node4055;
	wire [11-1:0] node4056;
	wire [11-1:0] node4057;
	wire [11-1:0] node4058;
	wire [11-1:0] node4061;
	wire [11-1:0] node4065;
	wire [11-1:0] node4066;
	wire [11-1:0] node4067;
	wire [11-1:0] node4070;
	wire [11-1:0] node4073;
	wire [11-1:0] node4074;
	wire [11-1:0] node4078;
	wire [11-1:0] node4079;
	wire [11-1:0] node4080;
	wire [11-1:0] node4081;
	wire [11-1:0] node4082;
	wire [11-1:0] node4083;
	wire [11-1:0] node4086;
	wire [11-1:0] node4089;
	wire [11-1:0] node4090;
	wire [11-1:0] node4093;
	wire [11-1:0] node4096;
	wire [11-1:0] node4097;
	wire [11-1:0] node4098;
	wire [11-1:0] node4102;
	wire [11-1:0] node4105;
	wire [11-1:0] node4106;
	wire [11-1:0] node4107;
	wire [11-1:0] node4108;
	wire [11-1:0] node4112;
	wire [11-1:0] node4114;
	wire [11-1:0] node4117;
	wire [11-1:0] node4118;
	wire [11-1:0] node4119;
	wire [11-1:0] node4122;
	wire [11-1:0] node4125;
	wire [11-1:0] node4126;
	wire [11-1:0] node4129;
	wire [11-1:0] node4132;
	wire [11-1:0] node4133;
	wire [11-1:0] node4134;
	wire [11-1:0] node4135;
	wire [11-1:0] node4138;
	wire [11-1:0] node4141;
	wire [11-1:0] node4142;
	wire [11-1:0] node4145;
	wire [11-1:0] node4146;
	wire [11-1:0] node4149;
	wire [11-1:0] node4152;
	wire [11-1:0] node4153;
	wire [11-1:0] node4154;
	wire [11-1:0] node4157;
	wire [11-1:0] node4159;
	wire [11-1:0] node4162;
	wire [11-1:0] node4163;
	wire [11-1:0] node4166;
	wire [11-1:0] node4169;
	wire [11-1:0] node4170;
	wire [11-1:0] node4171;
	wire [11-1:0] node4172;
	wire [11-1:0] node4173;
	wire [11-1:0] node4174;
	wire [11-1:0] node4175;
	wire [11-1:0] node4177;
	wire [11-1:0] node4180;
	wire [11-1:0] node4181;
	wire [11-1:0] node4184;
	wire [11-1:0] node4187;
	wire [11-1:0] node4188;
	wire [11-1:0] node4191;
	wire [11-1:0] node4193;
	wire [11-1:0] node4196;
	wire [11-1:0] node4197;
	wire [11-1:0] node4198;
	wire [11-1:0] node4201;
	wire [11-1:0] node4202;
	wire [11-1:0] node4206;
	wire [11-1:0] node4207;
	wire [11-1:0] node4208;
	wire [11-1:0] node4212;
	wire [11-1:0] node4213;
	wire [11-1:0] node4217;
	wire [11-1:0] node4218;
	wire [11-1:0] node4219;
	wire [11-1:0] node4220;
	wire [11-1:0] node4221;
	wire [11-1:0] node4225;
	wire [11-1:0] node4226;
	wire [11-1:0] node4230;
	wire [11-1:0] node4231;
	wire [11-1:0] node4232;
	wire [11-1:0] node4235;
	wire [11-1:0] node4238;
	wire [11-1:0] node4241;
	wire [11-1:0] node4242;
	wire [11-1:0] node4243;
	wire [11-1:0] node4245;
	wire [11-1:0] node4248;
	wire [11-1:0] node4249;
	wire [11-1:0] node4252;
	wire [11-1:0] node4255;
	wire [11-1:0] node4256;
	wire [11-1:0] node4257;
	wire [11-1:0] node4260;
	wire [11-1:0] node4263;
	wire [11-1:0] node4266;
	wire [11-1:0] node4267;
	wire [11-1:0] node4268;
	wire [11-1:0] node4269;
	wire [11-1:0] node4270;
	wire [11-1:0] node4271;
	wire [11-1:0] node4274;
	wire [11-1:0] node4277;
	wire [11-1:0] node4278;
	wire [11-1:0] node4281;
	wire [11-1:0] node4284;
	wire [11-1:0] node4285;
	wire [11-1:0] node4287;
	wire [11-1:0] node4290;
	wire [11-1:0] node4291;
	wire [11-1:0] node4294;
	wire [11-1:0] node4297;
	wire [11-1:0] node4298;
	wire [11-1:0] node4299;
	wire [11-1:0] node4301;
	wire [11-1:0] node4304;
	wire [11-1:0] node4305;
	wire [11-1:0] node4309;
	wire [11-1:0] node4310;
	wire [11-1:0] node4313;
	wire [11-1:0] node4314;
	wire [11-1:0] node4318;
	wire [11-1:0] node4319;
	wire [11-1:0] node4320;
	wire [11-1:0] node4321;
	wire [11-1:0] node4323;
	wire [11-1:0] node4326;
	wire [11-1:0] node4328;
	wire [11-1:0] node4331;
	wire [11-1:0] node4332;
	wire [11-1:0] node4334;
	wire [11-1:0] node4337;
	wire [11-1:0] node4339;
	wire [11-1:0] node4342;
	wire [11-1:0] node4343;
	wire [11-1:0] node4345;
	wire [11-1:0] node4346;
	wire [11-1:0] node4349;
	wire [11-1:0] node4352;
	wire [11-1:0] node4353;
	wire [11-1:0] node4354;
	wire [11-1:0] node4358;
	wire [11-1:0] node4359;
	wire [11-1:0] node4363;
	wire [11-1:0] node4364;
	wire [11-1:0] node4365;
	wire [11-1:0] node4366;
	wire [11-1:0] node4367;
	wire [11-1:0] node4368;
	wire [11-1:0] node4369;
	wire [11-1:0] node4373;
	wire [11-1:0] node4376;
	wire [11-1:0] node4377;
	wire [11-1:0] node4378;
	wire [11-1:0] node4381;
	wire [11-1:0] node4384;
	wire [11-1:0] node4387;
	wire [11-1:0] node4388;
	wire [11-1:0] node4389;
	wire [11-1:0] node4390;
	wire [11-1:0] node4394;
	wire [11-1:0] node4396;
	wire [11-1:0] node4399;
	wire [11-1:0] node4400;
	wire [11-1:0] node4403;
	wire [11-1:0] node4405;
	wire [11-1:0] node4408;
	wire [11-1:0] node4409;
	wire [11-1:0] node4410;
	wire [11-1:0] node4411;
	wire [11-1:0] node4412;
	wire [11-1:0] node4415;
	wire [11-1:0] node4418;
	wire [11-1:0] node4419;
	wire [11-1:0] node4423;
	wire [11-1:0] node4424;
	wire [11-1:0] node4426;
	wire [11-1:0] node4429;
	wire [11-1:0] node4431;
	wire [11-1:0] node4434;
	wire [11-1:0] node4435;
	wire [11-1:0] node4436;
	wire [11-1:0] node4439;
	wire [11-1:0] node4440;
	wire [11-1:0] node4444;
	wire [11-1:0] node4445;
	wire [11-1:0] node4446;
	wire [11-1:0] node4450;
	wire [11-1:0] node4451;
	wire [11-1:0] node4455;
	wire [11-1:0] node4456;
	wire [11-1:0] node4457;
	wire [11-1:0] node4458;
	wire [11-1:0] node4459;
	wire [11-1:0] node4461;
	wire [11-1:0] node4464;
	wire [11-1:0] node4467;
	wire [11-1:0] node4468;
	wire [11-1:0] node4469;
	wire [11-1:0] node4472;
	wire [11-1:0] node4475;
	wire [11-1:0] node4477;
	wire [11-1:0] node4480;
	wire [11-1:0] node4481;
	wire [11-1:0] node4482;
	wire [11-1:0] node4484;
	wire [11-1:0] node4487;
	wire [11-1:0] node4488;
	wire [11-1:0] node4491;
	wire [11-1:0] node4494;
	wire [11-1:0] node4495;
	wire [11-1:0] node4496;
	wire [11-1:0] node4500;
	wire [11-1:0] node4502;
	wire [11-1:0] node4505;
	wire [11-1:0] node4506;
	wire [11-1:0] node4507;
	wire [11-1:0] node4508;
	wire [11-1:0] node4509;
	wire [11-1:0] node4512;
	wire [11-1:0] node4515;
	wire [11-1:0] node4518;
	wire [11-1:0] node4519;
	wire [11-1:0] node4522;
	wire [11-1:0] node4523;
	wire [11-1:0] node4527;
	wire [11-1:0] node4528;
	wire [11-1:0] node4529;
	wire [11-1:0] node4531;
	wire [11-1:0] node4534;
	wire [11-1:0] node4536;
	wire [11-1:0] node4539;
	wire [11-1:0] node4540;
	wire [11-1:0] node4543;
	wire [11-1:0] node4544;
	wire [11-1:0] node4548;
	wire [11-1:0] node4549;
	wire [11-1:0] node4550;
	wire [11-1:0] node4551;
	wire [11-1:0] node4552;
	wire [11-1:0] node4553;
	wire [11-1:0] node4554;
	wire [11-1:0] node4555;
	wire [11-1:0] node4556;
	wire [11-1:0] node4559;
	wire [11-1:0] node4562;
	wire [11-1:0] node4563;
	wire [11-1:0] node4564;
	wire [11-1:0] node4567;
	wire [11-1:0] node4570;
	wire [11-1:0] node4571;
	wire [11-1:0] node4575;
	wire [11-1:0] node4576;
	wire [11-1:0] node4577;
	wire [11-1:0] node4578;
	wire [11-1:0] node4581;
	wire [11-1:0] node4584;
	wire [11-1:0] node4586;
	wire [11-1:0] node4589;
	wire [11-1:0] node4590;
	wire [11-1:0] node4591;
	wire [11-1:0] node4594;
	wire [11-1:0] node4597;
	wire [11-1:0] node4598;
	wire [11-1:0] node4602;
	wire [11-1:0] node4603;
	wire [11-1:0] node4604;
	wire [11-1:0] node4605;
	wire [11-1:0] node4609;
	wire [11-1:0] node4610;
	wire [11-1:0] node4613;
	wire [11-1:0] node4614;
	wire [11-1:0] node4618;
	wire [11-1:0] node4619;
	wire [11-1:0] node4620;
	wire [11-1:0] node4621;
	wire [11-1:0] node4624;
	wire [11-1:0] node4627;
	wire [11-1:0] node4629;
	wire [11-1:0] node4632;
	wire [11-1:0] node4633;
	wire [11-1:0] node4636;
	wire [11-1:0] node4637;
	wire [11-1:0] node4640;
	wire [11-1:0] node4643;
	wire [11-1:0] node4644;
	wire [11-1:0] node4645;
	wire [11-1:0] node4646;
	wire [11-1:0] node4647;
	wire [11-1:0] node4649;
	wire [11-1:0] node4652;
	wire [11-1:0] node4653;
	wire [11-1:0] node4656;
	wire [11-1:0] node4659;
	wire [11-1:0] node4660;
	wire [11-1:0] node4662;
	wire [11-1:0] node4665;
	wire [11-1:0] node4667;
	wire [11-1:0] node4670;
	wire [11-1:0] node4671;
	wire [11-1:0] node4672;
	wire [11-1:0] node4673;
	wire [11-1:0] node4676;
	wire [11-1:0] node4679;
	wire [11-1:0] node4682;
	wire [11-1:0] node4684;
	wire [11-1:0] node4685;
	wire [11-1:0] node4688;
	wire [11-1:0] node4691;
	wire [11-1:0] node4692;
	wire [11-1:0] node4693;
	wire [11-1:0] node4694;
	wire [11-1:0] node4695;
	wire [11-1:0] node4699;
	wire [11-1:0] node4700;
	wire [11-1:0] node4703;
	wire [11-1:0] node4706;
	wire [11-1:0] node4707;
	wire [11-1:0] node4708;
	wire [11-1:0] node4712;
	wire [11-1:0] node4713;
	wire [11-1:0] node4716;
	wire [11-1:0] node4719;
	wire [11-1:0] node4720;
	wire [11-1:0] node4721;
	wire [11-1:0] node4724;
	wire [11-1:0] node4727;
	wire [11-1:0] node4728;
	wire [11-1:0] node4729;
	wire [11-1:0] node4732;
	wire [11-1:0] node4735;
	wire [11-1:0] node4738;
	wire [11-1:0] node4739;
	wire [11-1:0] node4740;
	wire [11-1:0] node4741;
	wire [11-1:0] node4742;
	wire [11-1:0] node4743;
	wire [11-1:0] node4744;
	wire [11-1:0] node4747;
	wire [11-1:0] node4750;
	wire [11-1:0] node4751;
	wire [11-1:0] node4755;
	wire [11-1:0] node4756;
	wire [11-1:0] node4758;
	wire [11-1:0] node4761;
	wire [11-1:0] node4762;
	wire [11-1:0] node4765;
	wire [11-1:0] node4768;
	wire [11-1:0] node4769;
	wire [11-1:0] node4770;
	wire [11-1:0] node4771;
	wire [11-1:0] node4775;
	wire [11-1:0] node4777;
	wire [11-1:0] node4780;
	wire [11-1:0] node4781;
	wire [11-1:0] node4782;
	wire [11-1:0] node4786;
	wire [11-1:0] node4789;
	wire [11-1:0] node4790;
	wire [11-1:0] node4791;
	wire [11-1:0] node4792;
	wire [11-1:0] node4794;
	wire [11-1:0] node4797;
	wire [11-1:0] node4799;
	wire [11-1:0] node4802;
	wire [11-1:0] node4803;
	wire [11-1:0] node4805;
	wire [11-1:0] node4808;
	wire [11-1:0] node4809;
	wire [11-1:0] node4812;
	wire [11-1:0] node4815;
	wire [11-1:0] node4816;
	wire [11-1:0] node4817;
	wire [11-1:0] node4818;
	wire [11-1:0] node4821;
	wire [11-1:0] node4824;
	wire [11-1:0] node4826;
	wire [11-1:0] node4829;
	wire [11-1:0] node4830;
	wire [11-1:0] node4833;
	wire [11-1:0] node4835;
	wire [11-1:0] node4838;
	wire [11-1:0] node4839;
	wire [11-1:0] node4840;
	wire [11-1:0] node4841;
	wire [11-1:0] node4842;
	wire [11-1:0] node4844;
	wire [11-1:0] node4847;
	wire [11-1:0] node4848;
	wire [11-1:0] node4852;
	wire [11-1:0] node4853;
	wire [11-1:0] node4856;
	wire [11-1:0] node4857;
	wire [11-1:0] node4860;
	wire [11-1:0] node4863;
	wire [11-1:0] node4864;
	wire [11-1:0] node4865;
	wire [11-1:0] node4866;
	wire [11-1:0] node4869;
	wire [11-1:0] node4872;
	wire [11-1:0] node4873;
	wire [11-1:0] node4876;
	wire [11-1:0] node4879;
	wire [11-1:0] node4880;
	wire [11-1:0] node4881;
	wire [11-1:0] node4885;
	wire [11-1:0] node4887;
	wire [11-1:0] node4890;
	wire [11-1:0] node4891;
	wire [11-1:0] node4892;
	wire [11-1:0] node4893;
	wire [11-1:0] node4895;
	wire [11-1:0] node4898;
	wire [11-1:0] node4900;
	wire [11-1:0] node4903;
	wire [11-1:0] node4906;
	wire [11-1:0] node4907;
	wire [11-1:0] node4908;
	wire [11-1:0] node4909;
	wire [11-1:0] node4913;
	wire [11-1:0] node4914;
	wire [11-1:0] node4917;
	wire [11-1:0] node4920;
	wire [11-1:0] node4921;
	wire [11-1:0] node4922;
	wire [11-1:0] node4927;
	wire [11-1:0] node4928;
	wire [11-1:0] node4929;
	wire [11-1:0] node4930;
	wire [11-1:0] node4931;
	wire [11-1:0] node4932;
	wire [11-1:0] node4933;
	wire [11-1:0] node4934;
	wire [11-1:0] node4937;
	wire [11-1:0] node4941;
	wire [11-1:0] node4942;
	wire [11-1:0] node4943;
	wire [11-1:0] node4946;
	wire [11-1:0] node4949;
	wire [11-1:0] node4950;
	wire [11-1:0] node4954;
	wire [11-1:0] node4955;
	wire [11-1:0] node4956;
	wire [11-1:0] node4957;
	wire [11-1:0] node4961;
	wire [11-1:0] node4962;
	wire [11-1:0] node4965;
	wire [11-1:0] node4968;
	wire [11-1:0] node4969;
	wire [11-1:0] node4970;
	wire [11-1:0] node4975;
	wire [11-1:0] node4976;
	wire [11-1:0] node4977;
	wire [11-1:0] node4978;
	wire [11-1:0] node4979;
	wire [11-1:0] node4982;
	wire [11-1:0] node4985;
	wire [11-1:0] node4986;
	wire [11-1:0] node4990;
	wire [11-1:0] node4991;
	wire [11-1:0] node4992;
	wire [11-1:0] node4996;
	wire [11-1:0] node4998;
	wire [11-1:0] node5001;
	wire [11-1:0] node5002;
	wire [11-1:0] node5003;
	wire [11-1:0] node5005;
	wire [11-1:0] node5008;
	wire [11-1:0] node5009;
	wire [11-1:0] node5012;
	wire [11-1:0] node5015;
	wire [11-1:0] node5016;
	wire [11-1:0] node5019;
	wire [11-1:0] node5022;
	wire [11-1:0] node5023;
	wire [11-1:0] node5024;
	wire [11-1:0] node5025;
	wire [11-1:0] node5026;
	wire [11-1:0] node5027;
	wire [11-1:0] node5031;
	wire [11-1:0] node5032;
	wire [11-1:0] node5036;
	wire [11-1:0] node5037;
	wire [11-1:0] node5038;
	wire [11-1:0] node5041;
	wire [11-1:0] node5044;
	wire [11-1:0] node5045;
	wire [11-1:0] node5048;
	wire [11-1:0] node5051;
	wire [11-1:0] node5052;
	wire [11-1:0] node5053;
	wire [11-1:0] node5054;
	wire [11-1:0] node5057;
	wire [11-1:0] node5060;
	wire [11-1:0] node5062;
	wire [11-1:0] node5065;
	wire [11-1:0] node5066;
	wire [11-1:0] node5067;
	wire [11-1:0] node5071;
	wire [11-1:0] node5074;
	wire [11-1:0] node5075;
	wire [11-1:0] node5076;
	wire [11-1:0] node5077;
	wire [11-1:0] node5080;
	wire [11-1:0] node5083;
	wire [11-1:0] node5084;
	wire [11-1:0] node5085;
	wire [11-1:0] node5088;
	wire [11-1:0] node5091;
	wire [11-1:0] node5092;
	wire [11-1:0] node5095;
	wire [11-1:0] node5098;
	wire [11-1:0] node5099;
	wire [11-1:0] node5100;
	wire [11-1:0] node5103;
	wire [11-1:0] node5105;
	wire [11-1:0] node5108;
	wire [11-1:0] node5109;
	wire [11-1:0] node5110;
	wire [11-1:0] node5113;
	wire [11-1:0] node5116;
	wire [11-1:0] node5119;
	wire [11-1:0] node5120;
	wire [11-1:0] node5121;
	wire [11-1:0] node5122;
	wire [11-1:0] node5123;
	wire [11-1:0] node5124;
	wire [11-1:0] node5126;
	wire [11-1:0] node5129;
	wire [11-1:0] node5130;
	wire [11-1:0] node5133;
	wire [11-1:0] node5136;
	wire [11-1:0] node5137;
	wire [11-1:0] node5138;
	wire [11-1:0] node5142;
	wire [11-1:0] node5143;
	wire [11-1:0] node5146;
	wire [11-1:0] node5149;
	wire [11-1:0] node5150;
	wire [11-1:0] node5151;
	wire [11-1:0] node5152;
	wire [11-1:0] node5156;
	wire [11-1:0] node5157;
	wire [11-1:0] node5160;
	wire [11-1:0] node5163;
	wire [11-1:0] node5164;
	wire [11-1:0] node5165;
	wire [11-1:0] node5168;
	wire [11-1:0] node5171;
	wire [11-1:0] node5174;
	wire [11-1:0] node5175;
	wire [11-1:0] node5176;
	wire [11-1:0] node5177;
	wire [11-1:0] node5178;
	wire [11-1:0] node5182;
	wire [11-1:0] node5185;
	wire [11-1:0] node5186;
	wire [11-1:0] node5189;
	wire [11-1:0] node5190;
	wire [11-1:0] node5194;
	wire [11-1:0] node5195;
	wire [11-1:0] node5196;
	wire [11-1:0] node5197;
	wire [11-1:0] node5201;
	wire [11-1:0] node5202;
	wire [11-1:0] node5205;
	wire [11-1:0] node5208;
	wire [11-1:0] node5209;
	wire [11-1:0] node5211;
	wire [11-1:0] node5214;
	wire [11-1:0] node5215;
	wire [11-1:0] node5219;
	wire [11-1:0] node5220;
	wire [11-1:0] node5221;
	wire [11-1:0] node5222;
	wire [11-1:0] node5223;
	wire [11-1:0] node5226;
	wire [11-1:0] node5227;
	wire [11-1:0] node5231;
	wire [11-1:0] node5232;
	wire [11-1:0] node5233;
	wire [11-1:0] node5237;
	wire [11-1:0] node5238;
	wire [11-1:0] node5241;
	wire [11-1:0] node5244;
	wire [11-1:0] node5245;
	wire [11-1:0] node5246;
	wire [11-1:0] node5248;
	wire [11-1:0] node5251;
	wire [11-1:0] node5254;
	wire [11-1:0] node5255;
	wire [11-1:0] node5257;
	wire [11-1:0] node5260;
	wire [11-1:0] node5261;
	wire [11-1:0] node5265;
	wire [11-1:0] node5266;
	wire [11-1:0] node5267;
	wire [11-1:0] node5268;
	wire [11-1:0] node5270;
	wire [11-1:0] node5273;
	wire [11-1:0] node5275;
	wire [11-1:0] node5278;
	wire [11-1:0] node5279;
	wire [11-1:0] node5280;
	wire [11-1:0] node5285;
	wire [11-1:0] node5286;
	wire [11-1:0] node5287;
	wire [11-1:0] node5290;
	wire [11-1:0] node5291;
	wire [11-1:0] node5295;
	wire [11-1:0] node5296;
	wire [11-1:0] node5298;
	wire [11-1:0] node5301;
	wire [11-1:0] node5302;
	wire [11-1:0] node5306;
	wire [11-1:0] node5307;
	wire [11-1:0] node5308;
	wire [11-1:0] node5309;
	wire [11-1:0] node5310;
	wire [11-1:0] node5311;
	wire [11-1:0] node5312;
	wire [11-1:0] node5313;
	wire [11-1:0] node5316;
	wire [11-1:0] node5317;
	wire [11-1:0] node5321;
	wire [11-1:0] node5322;
	wire [11-1:0] node5324;
	wire [11-1:0] node5327;
	wire [11-1:0] node5328;
	wire [11-1:0] node5331;
	wire [11-1:0] node5334;
	wire [11-1:0] node5335;
	wire [11-1:0] node5336;
	wire [11-1:0] node5339;
	wire [11-1:0] node5340;
	wire [11-1:0] node5343;
	wire [11-1:0] node5346;
	wire [11-1:0] node5347;
	wire [11-1:0] node5348;
	wire [11-1:0] node5353;
	wire [11-1:0] node5354;
	wire [11-1:0] node5355;
	wire [11-1:0] node5356;
	wire [11-1:0] node5358;
	wire [11-1:0] node5361;
	wire [11-1:0] node5362;
	wire [11-1:0] node5365;
	wire [11-1:0] node5368;
	wire [11-1:0] node5370;
	wire [11-1:0] node5371;
	wire [11-1:0] node5374;
	wire [11-1:0] node5377;
	wire [11-1:0] node5378;
	wire [11-1:0] node5379;
	wire [11-1:0] node5380;
	wire [11-1:0] node5384;
	wire [11-1:0] node5385;
	wire [11-1:0] node5388;
	wire [11-1:0] node5391;
	wire [11-1:0] node5392;
	wire [11-1:0] node5394;
	wire [11-1:0] node5397;
	wire [11-1:0] node5398;
	wire [11-1:0] node5401;
	wire [11-1:0] node5404;
	wire [11-1:0] node5405;
	wire [11-1:0] node5406;
	wire [11-1:0] node5407;
	wire [11-1:0] node5408;
	wire [11-1:0] node5409;
	wire [11-1:0] node5413;
	wire [11-1:0] node5416;
	wire [11-1:0] node5417;
	wire [11-1:0] node5418;
	wire [11-1:0] node5421;
	wire [11-1:0] node5424;
	wire [11-1:0] node5425;
	wire [11-1:0] node5428;
	wire [11-1:0] node5431;
	wire [11-1:0] node5432;
	wire [11-1:0] node5433;
	wire [11-1:0] node5435;
	wire [11-1:0] node5438;
	wire [11-1:0] node5439;
	wire [11-1:0] node5442;
	wire [11-1:0] node5445;
	wire [11-1:0] node5446;
	wire [11-1:0] node5447;
	wire [11-1:0] node5451;
	wire [11-1:0] node5452;
	wire [11-1:0] node5455;
	wire [11-1:0] node5458;
	wire [11-1:0] node5459;
	wire [11-1:0] node5460;
	wire [11-1:0] node5461;
	wire [11-1:0] node5462;
	wire [11-1:0] node5465;
	wire [11-1:0] node5468;
	wire [11-1:0] node5471;
	wire [11-1:0] node5472;
	wire [11-1:0] node5474;
	wire [11-1:0] node5477;
	wire [11-1:0] node5478;
	wire [11-1:0] node5482;
	wire [11-1:0] node5483;
	wire [11-1:0] node5484;
	wire [11-1:0] node5486;
	wire [11-1:0] node5489;
	wire [11-1:0] node5492;
	wire [11-1:0] node5494;
	wire [11-1:0] node5497;
	wire [11-1:0] node5498;
	wire [11-1:0] node5499;
	wire [11-1:0] node5500;
	wire [11-1:0] node5501;
	wire [11-1:0] node5502;
	wire [11-1:0] node5503;
	wire [11-1:0] node5507;
	wire [11-1:0] node5510;
	wire [11-1:0] node5511;
	wire [11-1:0] node5512;
	wire [11-1:0] node5516;
	wire [11-1:0] node5517;
	wire [11-1:0] node5520;
	wire [11-1:0] node5523;
	wire [11-1:0] node5524;
	wire [11-1:0] node5525;
	wire [11-1:0] node5528;
	wire [11-1:0] node5529;
	wire [11-1:0] node5533;
	wire [11-1:0] node5534;
	wire [11-1:0] node5537;
	wire [11-1:0] node5538;
	wire [11-1:0] node5541;
	wire [11-1:0] node5544;
	wire [11-1:0] node5545;
	wire [11-1:0] node5546;
	wire [11-1:0] node5547;
	wire [11-1:0] node5550;
	wire [11-1:0] node5551;
	wire [11-1:0] node5554;
	wire [11-1:0] node5557;
	wire [11-1:0] node5558;
	wire [11-1:0] node5561;
	wire [11-1:0] node5564;
	wire [11-1:0] node5565;
	wire [11-1:0] node5566;
	wire [11-1:0] node5567;
	wire [11-1:0] node5570;
	wire [11-1:0] node5573;
	wire [11-1:0] node5575;
	wire [11-1:0] node5578;
	wire [11-1:0] node5579;
	wire [11-1:0] node5580;
	wire [11-1:0] node5583;
	wire [11-1:0] node5586;
	wire [11-1:0] node5589;
	wire [11-1:0] node5590;
	wire [11-1:0] node5591;
	wire [11-1:0] node5592;
	wire [11-1:0] node5593;
	wire [11-1:0] node5594;
	wire [11-1:0] node5598;
	wire [11-1:0] node5599;
	wire [11-1:0] node5603;
	wire [11-1:0] node5604;
	wire [11-1:0] node5606;
	wire [11-1:0] node5610;
	wire [11-1:0] node5611;
	wire [11-1:0] node5612;
	wire [11-1:0] node5615;
	wire [11-1:0] node5616;
	wire [11-1:0] node5619;
	wire [11-1:0] node5622;
	wire [11-1:0] node5623;
	wire [11-1:0] node5625;
	wire [11-1:0] node5628;
	wire [11-1:0] node5629;
	wire [11-1:0] node5632;
	wire [11-1:0] node5635;
	wire [11-1:0] node5636;
	wire [11-1:0] node5637;
	wire [11-1:0] node5638;
	wire [11-1:0] node5639;
	wire [11-1:0] node5643;
	wire [11-1:0] node5644;
	wire [11-1:0] node5647;
	wire [11-1:0] node5650;
	wire [11-1:0] node5651;
	wire [11-1:0] node5653;
	wire [11-1:0] node5656;
	wire [11-1:0] node5659;
	wire [11-1:0] node5660;
	wire [11-1:0] node5661;
	wire [11-1:0] node5662;
	wire [11-1:0] node5666;
	wire [11-1:0] node5667;
	wire [11-1:0] node5671;
	wire [11-1:0] node5672;
	wire [11-1:0] node5674;
	wire [11-1:0] node5677;
	wire [11-1:0] node5678;
	wire [11-1:0] node5682;
	wire [11-1:0] node5683;
	wire [11-1:0] node5684;
	wire [11-1:0] node5685;
	wire [11-1:0] node5686;
	wire [11-1:0] node5687;
	wire [11-1:0] node5688;
	wire [11-1:0] node5691;
	wire [11-1:0] node5694;
	wire [11-1:0] node5695;
	wire [11-1:0] node5699;
	wire [11-1:0] node5700;
	wire [11-1:0] node5701;
	wire [11-1:0] node5702;
	wire [11-1:0] node5705;
	wire [11-1:0] node5708;
	wire [11-1:0] node5709;
	wire [11-1:0] node5713;
	wire [11-1:0] node5714;
	wire [11-1:0] node5716;
	wire [11-1:0] node5719;
	wire [11-1:0] node5721;
	wire [11-1:0] node5724;
	wire [11-1:0] node5725;
	wire [11-1:0] node5726;
	wire [11-1:0] node5727;
	wire [11-1:0] node5728;
	wire [11-1:0] node5732;
	wire [11-1:0] node5733;
	wire [11-1:0] node5737;
	wire [11-1:0] node5738;
	wire [11-1:0] node5739;
	wire [11-1:0] node5742;
	wire [11-1:0] node5745;
	wire [11-1:0] node5746;
	wire [11-1:0] node5750;
	wire [11-1:0] node5751;
	wire [11-1:0] node5752;
	wire [11-1:0] node5755;
	wire [11-1:0] node5757;
	wire [11-1:0] node5760;
	wire [11-1:0] node5761;
	wire [11-1:0] node5762;
	wire [11-1:0] node5766;
	wire [11-1:0] node5769;
	wire [11-1:0] node5770;
	wire [11-1:0] node5771;
	wire [11-1:0] node5772;
	wire [11-1:0] node5773;
	wire [11-1:0] node5774;
	wire [11-1:0] node5778;
	wire [11-1:0] node5780;
	wire [11-1:0] node5783;
	wire [11-1:0] node5784;
	wire [11-1:0] node5785;
	wire [11-1:0] node5788;
	wire [11-1:0] node5791;
	wire [11-1:0] node5792;
	wire [11-1:0] node5795;
	wire [11-1:0] node5798;
	wire [11-1:0] node5799;
	wire [11-1:0] node5800;
	wire [11-1:0] node5802;
	wire [11-1:0] node5805;
	wire [11-1:0] node5806;
	wire [11-1:0] node5810;
	wire [11-1:0] node5811;
	wire [11-1:0] node5812;
	wire [11-1:0] node5816;
	wire [11-1:0] node5819;
	wire [11-1:0] node5820;
	wire [11-1:0] node5821;
	wire [11-1:0] node5822;
	wire [11-1:0] node5823;
	wire [11-1:0] node5826;
	wire [11-1:0] node5829;
	wire [11-1:0] node5832;
	wire [11-1:0] node5833;
	wire [11-1:0] node5836;
	wire [11-1:0] node5838;
	wire [11-1:0] node5841;
	wire [11-1:0] node5842;
	wire [11-1:0] node5843;
	wire [11-1:0] node5845;
	wire [11-1:0] node5849;
	wire [11-1:0] node5850;
	wire [11-1:0] node5852;
	wire [11-1:0] node5856;
	wire [11-1:0] node5857;
	wire [11-1:0] node5858;
	wire [11-1:0] node5859;
	wire [11-1:0] node5860;
	wire [11-1:0] node5861;
	wire [11-1:0] node5864;
	wire [11-1:0] node5867;
	wire [11-1:0] node5868;
	wire [11-1:0] node5869;
	wire [11-1:0] node5874;
	wire [11-1:0] node5875;
	wire [11-1:0] node5876;
	wire [11-1:0] node5877;
	wire [11-1:0] node5880;
	wire [11-1:0] node5883;
	wire [11-1:0] node5884;
	wire [11-1:0] node5887;
	wire [11-1:0] node5890;
	wire [11-1:0] node5891;
	wire [11-1:0] node5893;
	wire [11-1:0] node5896;
	wire [11-1:0] node5898;
	wire [11-1:0] node5901;
	wire [11-1:0] node5902;
	wire [11-1:0] node5903;
	wire [11-1:0] node5904;
	wire [11-1:0] node5906;
	wire [11-1:0] node5909;
	wire [11-1:0] node5910;
	wire [11-1:0] node5914;
	wire [11-1:0] node5915;
	wire [11-1:0] node5917;
	wire [11-1:0] node5920;
	wire [11-1:0] node5921;
	wire [11-1:0] node5925;
	wire [11-1:0] node5926;
	wire [11-1:0] node5927;
	wire [11-1:0] node5928;
	wire [11-1:0] node5932;
	wire [11-1:0] node5933;
	wire [11-1:0] node5937;
	wire [11-1:0] node5938;
	wire [11-1:0] node5940;
	wire [11-1:0] node5944;
	wire [11-1:0] node5945;
	wire [11-1:0] node5946;
	wire [11-1:0] node5947;
	wire [11-1:0] node5948;
	wire [11-1:0] node5949;
	wire [11-1:0] node5954;
	wire [11-1:0] node5955;
	wire [11-1:0] node5957;
	wire [11-1:0] node5960;
	wire [11-1:0] node5961;
	wire [11-1:0] node5965;
	wire [11-1:0] node5966;
	wire [11-1:0] node5967;
	wire [11-1:0] node5968;
	wire [11-1:0] node5971;
	wire [11-1:0] node5974;
	wire [11-1:0] node5976;
	wire [11-1:0] node5979;
	wire [11-1:0] node5980;
	wire [11-1:0] node5983;
	wire [11-1:0] node5986;
	wire [11-1:0] node5987;
	wire [11-1:0] node5988;
	wire [11-1:0] node5989;
	wire [11-1:0] node5991;
	wire [11-1:0] node5994;
	wire [11-1:0] node5997;
	wire [11-1:0] node5998;
	wire [11-1:0] node5999;
	wire [11-1:0] node6003;
	wire [11-1:0] node6004;
	wire [11-1:0] node6008;
	wire [11-1:0] node6009;
	wire [11-1:0] node6010;
	wire [11-1:0] node6011;
	wire [11-1:0] node6015;
	wire [11-1:0] node6016;
	wire [11-1:0] node6019;
	wire [11-1:0] node6022;
	wire [11-1:0] node6023;

	assign outp = (inp[1]) ? node3032 : node1;
		assign node1 = (inp[7]) ? node1503 : node2;
			assign node2 = (inp[2]) ? node746 : node3;
				assign node3 = (inp[0]) ? node387 : node4;
					assign node4 = (inp[4]) ? node206 : node5;
						assign node5 = (inp[9]) ? node93 : node6;
							assign node6 = (inp[5]) ? node48 : node7;
								assign node7 = (inp[6]) ? node25 : node8;
									assign node8 = (inp[8]) ? node18 : node9;
										assign node9 = (inp[10]) ? node15 : node10;
											assign node10 = (inp[3]) ? node12 : 11'b01001101011;
												assign node12 = (inp[11]) ? 11'b11001111011 : 11'b11001101011;
											assign node15 = (inp[3]) ? 11'b01000101111 : 11'b11000101011;
										assign node18 = (inp[10]) ? node22 : node19;
											assign node19 = (inp[11]) ? 11'b01000001001 : 11'b01000001010;
											assign node22 = (inp[11]) ? 11'b11111101001 : 11'b11001101011;
									assign node25 = (inp[8]) ? node35 : node26;
										assign node26 = (inp[11]) ? node32 : node27;
											assign node27 = (inp[10]) ? 11'b11000100010 : node28;
												assign node28 = (inp[3]) ? 11'b11011100010 : 11'b01001100010;
											assign node32 = (inp[3]) ? 11'b11000010010 : 11'b01010000010;
										assign node35 = (inp[3]) ? node43 : node36;
											assign node36 = (inp[10]) ? node40 : node37;
												assign node37 = (inp[11]) ? 11'b01011101000 : 11'b01000101010;
												assign node40 = (inp[11]) ? 11'b11110101000 : 11'b11011001010;
											assign node43 = (inp[11]) ? node45 : 11'b01101001100;
												assign node45 = (inp[10]) ? 11'b01010111110 : 11'b11101111000;
								assign node48 = (inp[6]) ? node70 : node49;
									assign node49 = (inp[11]) ? node61 : node50;
										assign node50 = (inp[10]) ? node58 : node51;
											assign node51 = (inp[8]) ? node55 : node52;
												assign node52 = (inp[3]) ? 11'b11001111010 : 11'b01001111010;
												assign node55 = (inp[3]) ? 11'b11000011011 : 11'b01000011011;
											assign node58 = (inp[3]) ? 11'b01111111110 : 11'b11101111010;
										assign node61 = (inp[8]) ? node67 : node62;
											assign node62 = (inp[3]) ? node64 : 11'b11101111000;
												assign node64 = (inp[10]) ? 11'b01010101100 : 11'b11101101000;
											assign node67 = (inp[10]) ? 11'b01001101110 : 11'b11010001010;
									assign node70 = (inp[10]) ? node80 : node71;
										assign node71 = (inp[8]) ? node77 : node72;
											assign node72 = (inp[3]) ? 11'b11011011011 : node73;
												assign node73 = (inp[11]) ? 11'b01011011001 : 11'b01001011011;
											assign node77 = (inp[11]) ? 11'b01010011011 : 11'b01000111011;
										assign node80 = (inp[3]) ? node88 : node81;
											assign node81 = (inp[8]) ? node85 : node82;
												assign node82 = (inp[11]) ? 11'b11110011001 : 11'b11101011001;
												assign node85 = (inp[11]) ? 11'b11001111001 : 11'b11110111001;
											assign node88 = (inp[8]) ? node90 : 11'b01110011101;
												assign node90 = (inp[11]) ? 11'b01011101101 : 11'b01101111101;
							assign node93 = (inp[11]) ? node153 : node94;
								assign node94 = (inp[10]) ? node124 : node95;
									assign node95 = (inp[3]) ? node111 : node96;
										assign node96 = (inp[5]) ? node104 : node97;
											assign node97 = (inp[6]) ? node101 : node98;
												assign node98 = (inp[8]) ? 11'b01010101011 : 11'b01001101011;
												assign node101 = (inp[8]) ? 11'b01010001000 : 11'b01000100000;
											assign node104 = (inp[6]) ? node108 : node105;
												assign node105 = (inp[8]) ? 11'b01010111010 : 11'b01001111010;
												assign node108 = (inp[8]) ? 11'b01001111011 : 11'b01010011001;
										assign node111 = (inp[5]) ? node117 : node112;
											assign node112 = (inp[6]) ? 11'b11011100100 : node113;
												assign node113 = (inp[8]) ? 11'b11111101111 : 11'b11001101111;
											assign node117 = (inp[6]) ? node121 : node118;
												assign node118 = (inp[8]) ? 11'b11000111100 : 11'b11001111110;
												assign node121 = (inp[8]) ? 11'b11010111111 : 11'b11001111111;
									assign node124 = (inp[5]) ? node138 : node125;
										assign node125 = (inp[6]) ? node131 : node126;
											assign node126 = (inp[8]) ? 11'b11011111111 : node127;
												assign node127 = (inp[3]) ? 11'b01000111111 : 11'b11000111111;
											assign node131 = (inp[8]) ? node135 : node132;
												assign node132 = (inp[3]) ? 11'b01010110100 : 11'b11001110100;
												assign node135 = (inp[3]) ? 11'b01111011110 : 11'b11001011110;
										assign node138 = (inp[3]) ? node146 : node139;
											assign node139 = (inp[6]) ? node143 : node140;
												assign node140 = (inp[8]) ? 11'b11000101100 : 11'b11100101110;
												assign node143 = (inp[8]) ? 11'b11010101111 : 11'b11111101111;
											assign node146 = (inp[8]) ? node150 : node147;
												assign node147 = (inp[6]) ? 11'b01000101111 : 11'b01010101110;
												assign node150 = (inp[6]) ? 11'b01100101101 : 11'b01101101100;
								assign node153 = (inp[6]) ? node181 : node154;
									assign node154 = (inp[5]) ? node170 : node155;
										assign node155 = (inp[8]) ? node163 : node156;
											assign node156 = (inp[10]) ? node160 : node157;
												assign node157 = (inp[3]) ? 11'b11101101111 : 11'b01101111011;
												assign node160 = (inp[3]) ? 11'b01010111111 : 11'b11100111111;
											assign node163 = (inp[10]) ? node167 : node164;
												assign node164 = (inp[3]) ? 11'b11100101101 : 11'b01110111001;
												assign node167 = (inp[3]) ? 11'b01101111101 : 11'b11001111101;
										assign node170 = (inp[8]) ? node176 : node171;
											assign node171 = (inp[3]) ? 11'b11011111100 : node172;
												assign node172 = (inp[10]) ? 11'b11111101100 : 11'b01110101000;
											assign node176 = (inp[3]) ? node178 : 11'b01001101010;
												assign node178 = (inp[10]) ? 11'b01111101110 : 11'b11100111110;
									assign node181 = (inp[8]) ? node193 : node182;
										assign node182 = (inp[5]) ? node188 : node183;
											assign node183 = (inp[3]) ? 11'b11100101101 : node184;
												assign node184 = (inp[10]) ? 11'b11110111101 : 11'b01111111001;
											assign node188 = (inp[10]) ? node190 : 11'b11010011111;
												assign node190 = (inp[3]) ? 11'b01010001101 : 11'b11100001101;
										assign node193 = (inp[5]) ? node201 : node194;
											assign node194 = (inp[10]) ? node198 : node195;
												assign node195 = (inp[3]) ? 11'b11111001110 : 11'b01101011010;
												assign node198 = (inp[3]) ? 11'b01100011100 : 11'b11011011100;
											assign node201 = (inp[10]) ? node203 : 11'b11100111111;
												assign node203 = (inp[3]) ? 11'b01111101111 : 11'b11111101111;
						assign node206 = (inp[10]) ? node300 : node207;
							assign node207 = (inp[3]) ? node255 : node208;
								assign node208 = (inp[8]) ? node228 : node209;
									assign node209 = (inp[5]) ? node219 : node210;
										assign node210 = (inp[11]) ? node214 : node211;
											assign node211 = (inp[9]) ? 11'b01101001111 : 11'b01001001111;
											assign node214 = (inp[9]) ? node216 : 11'b01011101111;
												assign node216 = (inp[6]) ? 11'b01001011101 : 11'b01011011111;
										assign node219 = (inp[11]) ? node223 : node220;
											assign node220 = (inp[9]) ? 11'b01111011110 : 11'b01011011110;
											assign node223 = (inp[9]) ? 11'b01011101110 : node224;
												assign node224 = (inp[6]) ? 11'b01001111100 : 11'b01000111100;
									assign node228 = (inp[5]) ? node242 : node229;
										assign node229 = (inp[6]) ? node235 : node230;
											assign node230 = (inp[9]) ? 11'b01000011111 : node231;
												assign node231 = (inp[11]) ? 11'b01110101101 : 11'b01100101111;
											assign node235 = (inp[9]) ? node239 : node236;
												assign node236 = (inp[11]) ? 11'b01110001100 : 11'b01100001110;
												assign node239 = (inp[11]) ? 11'b01010011100 : 11'b01111101100;
										assign node242 = (inp[9]) ? node250 : node243;
											assign node243 = (inp[6]) ? node247 : node244;
												assign node244 = (inp[11]) ? 11'b01101111100 : 11'b01111111100;
												assign node247 = (inp[11]) ? 11'b01101111101 : 11'b01111011101;
											assign node250 = (inp[6]) ? 11'b01101001111 : node251;
												assign node251 = (inp[11]) ? 11'b01101001100 : 11'b01101011100;
								assign node255 = (inp[9]) ? node277 : node256;
									assign node256 = (inp[5]) ? node264 : node257;
										assign node257 = (inp[11]) ? node261 : node258;
											assign node258 = (inp[6]) ? 11'b11000001100 : 11'b11001001111;
											assign node261 = (inp[8]) ? 11'b11010101101 : 11'b11100101111;
										assign node264 = (inp[11]) ? node272 : node265;
											assign node265 = (inp[6]) ? node269 : node266;
												assign node266 = (inp[8]) ? 11'b11010111100 : 11'b11111011110;
												assign node269 = (inp[8]) ? 11'b11011011101 : 11'b11100111101;
											assign node272 = (inp[6]) ? 11'b11111111100 : node273;
												assign node273 = (inp[8]) ? 11'b11101111100 : 11'b11101011100;
									assign node277 = (inp[5]) ? node291 : node278;
										assign node278 = (inp[6]) ? node286 : node279;
											assign node279 = (inp[8]) ? node283 : node280;
												assign node280 = (inp[11]) ? 11'b11011011011 : 11'b11101011011;
												assign node283 = (inp[11]) ? 11'b11010011011 : 11'b11011011011;
											assign node286 = (inp[8]) ? node288 : 11'b11011011001;
												assign node288 = (inp[11]) ? 11'b11000011000 : 11'b11010111010;
										assign node291 = (inp[8]) ? node295 : node292;
											assign node292 = (inp[6]) ? 11'b11010101011 : 11'b11001001000;
											assign node295 = (inp[6]) ? 11'b11101001001 : node296;
												assign node296 = (inp[11]) ? 11'b11101001000 : 11'b11110001000;
							assign node300 = (inp[3]) ? node344 : node301;
								assign node301 = (inp[9]) ? node321 : node302;
									assign node302 = (inp[5]) ? node316 : node303;
										assign node303 = (inp[8]) ? node309 : node304;
											assign node304 = (inp[11]) ? 11'b11110111111 : node305;
												assign node305 = (inp[6]) ? 11'b11001010110 : 11'b11000011111;
											assign node309 = (inp[6]) ? node313 : node310;
												assign node310 = (inp[11]) ? 11'b11111011101 : 11'b11101011111;
												assign node313 = (inp[11]) ? 11'b11101011110 : 11'b11110011100;
										assign node316 = (inp[8]) ? 11'b11110101101 : node317;
											assign node317 = (inp[6]) ? 11'b11010101110 : 11'b11010001110;
									assign node321 = (inp[5]) ? node331 : node322;
										assign node322 = (inp[6]) ? node328 : node323;
											assign node323 = (inp[11]) ? node325 : 11'b11100001011;
												assign node325 = (inp[8]) ? 11'b11111011011 : 11'b11110011011;
											assign node328 = (inp[8]) ? 11'b11000101010 : 11'b11101000000;
										assign node331 = (inp[8]) ? node337 : node332;
											assign node332 = (inp[11]) ? node334 : 11'b11001011000;
												assign node334 = (inp[6]) ? 11'b11001101000 : 11'b11011001000;
											assign node337 = (inp[11]) ? node341 : node338;
												assign node338 = (inp[6]) ? 11'b11101011001 : 11'b11110011000;
												assign node341 = (inp[6]) ? 11'b11110001001 : 11'b11110001000;
								assign node344 = (inp[5]) ? node368 : node345;
									assign node345 = (inp[6]) ? node359 : node346;
										assign node346 = (inp[8]) ? node352 : node347;
											assign node347 = (inp[11]) ? 11'b01110011011 : node348;
												assign node348 = (inp[9]) ? 11'b01100011011 : 11'b01100001011;
											assign node352 = (inp[9]) ? node356 : node353;
												assign node353 = (inp[11]) ? 11'b01101011011 : 11'b01010001011;
												assign node356 = (inp[11]) ? 11'b01111011011 : 11'b01101011001;
										assign node359 = (inp[8]) ? node363 : node360;
											assign node360 = (inp[9]) ? 11'b01111010000 : 11'b01110000010;
											assign node363 = (inp[9]) ? node365 : 11'b01110011010;
												assign node365 = (inp[11]) ? 11'b01111111011 : 11'b01111111010;
									assign node368 = (inp[6]) ? node376 : node369;
										assign node369 = (inp[11]) ? 11'b01110101000 : node370;
											assign node370 = (inp[9]) ? node372 : 11'b01001011000;
												assign node372 = (inp[8]) ? 11'b01101001010 : 11'b01100001000;
										assign node376 = (inp[9]) ? node384 : node377;
											assign node377 = (inp[11]) ? node381 : node378;
												assign node378 = (inp[8]) ? 11'b01000011011 : 11'b01011111001;
												assign node381 = (inp[8]) ? 11'b01111001011 : 11'b01100101010;
											assign node384 = (inp[8]) ? 11'b01110001001 : 11'b01111001011;
					assign node387 = (inp[3]) ? node581 : node388;
						assign node388 = (inp[4]) ? node490 : node389;
							assign node389 = (inp[11]) ? node441 : node390;
								assign node390 = (inp[8]) ? node414 : node391;
									assign node391 = (inp[6]) ? node405 : node392;
										assign node392 = (inp[10]) ? node400 : node393;
											assign node393 = (inp[5]) ? node397 : node394;
												assign node394 = (inp[9]) ? 11'b01001101101 : 11'b01001101001;
												assign node397 = (inp[9]) ? 11'b01001101100 : 11'b01001101000;
											assign node400 = (inp[5]) ? node402 : 11'b01000111001;
												assign node402 = (inp[9]) ? 11'b01100111000 : 11'b01100101100;
										assign node405 = (inp[5]) ? node409 : node406;
											assign node406 = (inp[10]) ? 11'b01010100100 : 11'b01011100000;
											assign node409 = (inp[10]) ? 11'b01110001111 : node410;
												assign node410 = (inp[9]) ? 11'b01011101111 : 11'b01011001001;
									assign node414 = (inp[10]) ? node430 : node415;
										assign node415 = (inp[9]) ? node423 : node416;
											assign node416 = (inp[6]) ? node420 : node417;
												assign node417 = (inp[5]) ? 11'b01100001001 : 11'b01100001000;
												assign node420 = (inp[5]) ? 11'b01110101001 : 11'b01110101000;
											assign node423 = (inp[6]) ? node427 : node424;
												assign node424 = (inp[5]) ? 11'b01110101100 : 11'b01110101101;
												assign node427 = (inp[5]) ? 11'b01101101101 : 11'b01100001110;
										assign node430 = (inp[9]) ? node436 : node431;
											assign node431 = (inp[5]) ? node433 : 11'b01111001100;
												assign node433 = (inp[6]) ? 11'b01001101111 : 11'b01011101100;
											assign node436 = (inp[5]) ? 11'b01010111001 : node437;
												assign node437 = (inp[6]) ? 11'b01101011000 : 11'b01111111001;
								assign node441 = (inp[10]) ? node467 : node442;
									assign node442 = (inp[9]) ? node454 : node443;
										assign node443 = (inp[6]) ? node449 : node444;
											assign node444 = (inp[5]) ? node446 : 11'b01100011011;
												assign node446 = (inp[8]) ? 11'b01101011000 : 11'b01001111010;
											assign node449 = (inp[5]) ? node451 : 11'b01111111010;
												assign node451 = (inp[8]) ? 11'b01110011001 : 11'b01010011011;
										assign node454 = (inp[8]) ? node460 : node455;
											assign node455 = (inp[6]) ? node457 : 11'b01111111110;
												assign node457 = (inp[5]) ? 11'b01101011101 : 11'b01110111111;
											assign node460 = (inp[6]) ? node464 : node461;
												assign node461 = (inp[5]) ? 11'b01001111100 : 11'b01000111111;
												assign node464 = (inp[5]) ? 11'b01010111111 : 11'b01011011100;
									assign node467 = (inp[9]) ? node479 : node468;
										assign node468 = (inp[8]) ? node476 : node469;
											assign node469 = (inp[5]) ? node473 : node470;
												assign node470 = (inp[6]) ? 11'b01011111101 : 11'b01000111101;
												assign node473 = (inp[6]) ? 11'b01000011101 : 11'b01010111110;
											assign node476 = (inp[6]) ? 11'b01100111100 : 11'b01111111111;
										assign node479 = (inp[6]) ? node483 : node480;
											assign node480 = (inp[5]) ? 11'b01110101010 : 11'b01010101001;
											assign node483 = (inp[8]) ? node487 : node484;
												assign node484 = (inp[5]) ? 11'b01100001011 : 11'b01000101001;
												assign node487 = (inp[5]) ? 11'b01001101001 : 11'b01110001010;
							assign node490 = (inp[5]) ? node540 : node491;
								assign node491 = (inp[6]) ? node515 : node492;
									assign node492 = (inp[11]) ? node504 : node493;
										assign node493 = (inp[9]) ? node499 : node494;
											assign node494 = (inp[10]) ? 11'b01101011101 : node495;
												assign node495 = (inp[8]) ? 11'b01100101001 : 11'b01001001001;
											assign node499 = (inp[10]) ? node501 : 11'b01010011101;
												assign node501 = (inp[8]) ? 11'b01001011011 : 11'b01100011001;
										assign node504 = (inp[9]) ? node510 : node505;
											assign node505 = (inp[10]) ? 11'b01001001101 : node506;
												assign node506 = (inp[8]) ? 11'b01110111011 : 11'b01011011001;
											assign node510 = (inp[10]) ? node512 : 11'b01100001101;
												assign node512 = (inp[8]) ? 11'b01011001001 : 11'b01110001001;
									assign node515 = (inp[11]) ? node529 : node516;
										assign node516 = (inp[8]) ? node524 : node517;
											assign node517 = (inp[9]) ? node521 : node518;
												assign node518 = (inp[10]) ? 11'b01011010100 : 11'b01010100000;
												assign node521 = (inp[10]) ? 11'b01111010010 : 11'b01110010110;
											assign node524 = (inp[9]) ? 11'b01001111100 : node525;
												assign node525 = (inp[10]) ? 11'b01111111110 : 11'b01110001000;
										assign node529 = (inp[10]) ? node533 : node530;
											assign node530 = (inp[9]) ? 11'b01110001110 : 11'b01100011000;
											assign node533 = (inp[8]) ? node537 : node534;
												assign node534 = (inp[9]) ? 11'b01100001001 : 11'b01100101111;
												assign node537 = (inp[9]) ? 11'b01001101001 : 11'b01011001100;
								assign node540 = (inp[6]) ? node562 : node541;
									assign node541 = (inp[8]) ? node555 : node542;
										assign node542 = (inp[10]) ? node548 : node543;
											assign node543 = (inp[9]) ? 11'b01111001110 : node544;
												assign node544 = (inp[11]) ? 11'b01101011010 : 11'b01111001000;
											assign node548 = (inp[11]) ? node552 : node549;
												assign node549 = (inp[9]) ? 11'b01100011010 : 11'b01010011100;
												assign node552 = (inp[9]) ? 11'b01110001010 : 11'b01100001110;
										assign node555 = (inp[10]) ? 11'b01101011110 : node556;
											assign node556 = (inp[11]) ? node558 : 11'b01010101010;
												assign node558 = (inp[9]) ? 11'b01001001110 : 11'b01001111010;
									assign node562 = (inp[8]) ? node572 : node563;
										assign node563 = (inp[11]) ? 11'b01111111010 : node564;
											assign node564 = (inp[10]) ? node568 : node565;
												assign node565 = (inp[9]) ? 11'b01100111101 : 11'b01100101011;
												assign node568 = (inp[9]) ? 11'b01111011001 : 11'b01001111111;
										assign node572 = (inp[9]) ? node576 : node573;
											assign node573 = (inp[10]) ? 11'b01000101101 : 11'b01010111011;
											assign node576 = (inp[10]) ? node578 : 11'b01001011111;
												assign node578 = (inp[11]) ? 11'b01000001011 : 11'b01010011011;
						assign node581 = (inp[10]) ? node663 : node582;
							assign node582 = (inp[4]) ? node624 : node583;
								assign node583 = (inp[9]) ? node607 : node584;
									assign node584 = (inp[5]) ? node594 : node585;
										assign node585 = (inp[11]) ? node591 : node586;
											assign node586 = (inp[6]) ? node588 : 11'b01001101001;
												assign node588 = (inp[8]) ? 11'b01001001000 : 11'b01001100000;
											assign node591 = (inp[8]) ? 11'b01010101010 : 11'b01000000000;
										assign node594 = (inp[6]) ? node600 : node595;
											assign node595 = (inp[8]) ? node597 : 11'b01101101000;
												assign node597 = (inp[11]) ? 11'b01110001000 : 11'b01100001001;
											assign node600 = (inp[8]) ? node604 : node601;
												assign node601 = (inp[11]) ? 11'b01100001011 : 11'b01101001011;
												assign node604 = (inp[11]) ? 11'b01111101001 : 11'b01100101011;
									assign node607 = (inp[5]) ? node617 : node608;
										assign node608 = (inp[6]) ? node614 : node609;
											assign node609 = (inp[11]) ? 11'b01101111011 : node610;
												assign node610 = (inp[8]) ? 11'b01011111001 : 11'b01001111001;
											assign node614 = (inp[11]) ? 11'b01101011010 : 11'b01011011010;
										assign node617 = (inp[11]) ? node621 : node618;
											assign node618 = (inp[8]) ? 11'b01100111001 : 11'b01101111001;
											assign node621 = (inp[8]) ? 11'b01010111000 : 11'b01010011001;
								assign node624 = (inp[9]) ? node640 : node625;
									assign node625 = (inp[8]) ? node633 : node626;
										assign node626 = (inp[5]) ? node630 : node627;
											assign node627 = (inp[6]) ? 11'b01001010000 : 11'b01111011001;
											assign node630 = (inp[6]) ? 11'b01111111011 : 11'b01001011010;
										assign node633 = (inp[5]) ? node635 : 11'b01000011010;
											assign node635 = (inp[6]) ? node637 : 11'b01110111010;
												assign node637 = (inp[11]) ? 11'b01010111011 : 11'b01110011011;
									assign node640 = (inp[5]) ? node652 : node641;
										assign node641 = (inp[6]) ? node647 : node642;
											assign node642 = (inp[8]) ? node644 : 11'b01111001001;
												assign node644 = (inp[11]) ? 11'b01110001001 : 11'b01111001001;
											assign node647 = (inp[8]) ? node649 : 11'b01101000010;
												assign node649 = (inp[11]) ? 11'b01111101011 : 11'b01110101000;
										assign node652 = (inp[6]) ? node658 : node653;
											assign node653 = (inp[8]) ? 11'b01010001010 : node654;
												assign node654 = (inp[11]) ? 11'b01011001010 : 11'b01001001010;
											assign node658 = (inp[8]) ? 11'b01011001011 : node659;
												assign node659 = (inp[11]) ? 11'b01011101010 : 11'b01000101001;
							assign node663 = (inp[4]) ? node701 : node664;
								assign node664 = (inp[11]) ? node682 : node665;
									assign node665 = (inp[6]) ? node673 : node666;
										assign node666 = (inp[5]) ? node670 : node667;
											assign node667 = (inp[9]) ? 11'b01000101001 : 11'b01010101001;
											assign node670 = (inp[9]) ? 11'b01010101000 : 11'b01000101000;
										assign node673 = (inp[5]) ? node677 : node674;
											assign node674 = (inp[9]) ? 11'b01000100000 : 11'b01000100010;
											assign node677 = (inp[8]) ? 11'b01011001011 : node678;
												assign node678 = (inp[9]) ? 11'b01010101001 : 11'b01000001011;
									assign node682 = (inp[9]) ? node692 : node683;
										assign node683 = (inp[6]) ? node687 : node684;
											assign node684 = (inp[8]) ? 11'b01110101011 : 11'b01110101010;
											assign node687 = (inp[8]) ? node689 : 11'b01111001001;
												assign node689 = (inp[5]) ? 11'b01100101011 : 11'b01110101000;
										assign node692 = (inp[5]) ? node696 : node693;
											assign node693 = (inp[8]) ? 11'b01010001010 : 11'b01011101001;
											assign node696 = (inp[6]) ? 11'b01001101011 : node697;
												assign node697 = (inp[8]) ? 11'b01001101010 : 11'b01000101010;
								assign node701 = (inp[9]) ? node725 : node702;
									assign node702 = (inp[11]) ? node714 : node703;
										assign node703 = (inp[8]) ? node709 : node704;
											assign node704 = (inp[6]) ? 11'b01100000010 : node705;
												assign node705 = (inp[5]) ? 11'b01110001000 : 11'b01100001001;
											assign node709 = (inp[5]) ? node711 : 11'b01111101010;
												assign node711 = (inp[6]) ? 11'b01100001001 : 11'b01101001010;
										assign node714 = (inp[8]) ? node718 : node715;
											assign node715 = (inp[5]) ? 11'b01010001010 : 11'b01011001011;
											assign node718 = (inp[6]) ? node722 : node719;
												assign node719 = (inp[5]) ? 11'b01001001010 : 11'b01001001001;
												assign node722 = (inp[5]) ? 11'b01001001001 : 11'b01000001010;
									assign node725 = (inp[11]) ? node739 : node726;
										assign node726 = (inp[6]) ? node732 : node727;
											assign node727 = (inp[5]) ? 11'b01001001000 : node728;
												assign node728 = (inp[8]) ? 11'b01000001011 : 11'b01000001001;
											assign node732 = (inp[5]) ? node736 : node733;
												assign node733 = (inp[8]) ? 11'b01001101010 : 11'b01001000000;
												assign node736 = (inp[8]) ? 11'b01000001001 : 11'b01001001011;
										assign node739 = (inp[6]) ? node741 : 11'b01000001000;
											assign node741 = (inp[8]) ? 11'b01000001001 : node742;
												assign node742 = (inp[5]) ? 11'b01000101000 : 11'b01000001001;
				assign node746 = (inp[0]) ? node1118 : node747;
					assign node747 = (inp[8]) ? node935 : node748;
						assign node748 = (inp[6]) ? node838 : node749;
							assign node749 = (inp[4]) ? node789 : node750;
								assign node750 = (inp[5]) ? node768 : node751;
									assign node751 = (inp[9]) ? node761 : node752;
										assign node752 = (inp[11]) ? node758 : node753;
											assign node753 = (inp[10]) ? 11'b11110001010 : node754;
												assign node754 = (inp[3]) ? 11'b11101001010 : 11'b01101001010;
											assign node758 = (inp[10]) ? 11'b11111000011 : 11'b01100000011;
										assign node761 = (inp[3]) ? node763 : 11'b01010010011;
											assign node763 = (inp[10]) ? 11'b01101110101 : node764;
												assign node764 = (inp[11]) ? 11'b11011100111 : 11'b11101100111;
									assign node768 = (inp[11]) ? node782 : node769;
										assign node769 = (inp[10]) ? node777 : node770;
											assign node770 = (inp[3]) ? node774 : node771;
												assign node771 = (inp[9]) ? 11'b01101010001 : 11'b01100010011;
												assign node774 = (inp[9]) ? 11'b11110010101 : 11'b11100010011;
											assign node777 = (inp[9]) ? 11'b11000000101 : node778;
												assign node778 = (inp[3]) ? 11'b01001010101 : 11'b11011010011;
										assign node782 = (inp[10]) ? 11'b11010000110 : node783;
											assign node783 = (inp[3]) ? 11'b11011000000 : node784;
												assign node784 = (inp[9]) ? 11'b01011000000 : 11'b01101010000;
								assign node789 = (inp[5]) ? node815 : node790;
									assign node790 = (inp[9]) ? node802 : node791;
										assign node791 = (inp[3]) ? node797 : node792;
											assign node792 = (inp[10]) ? 11'b11111110101 : node793;
												assign node793 = (inp[11]) ? 11'b01110100101 : 11'b01100100101;
											assign node797 = (inp[10]) ? 11'b01000100001 : node798;
												assign node798 = (inp[11]) ? 11'b11000100101 : 11'b11101100101;
										assign node802 = (inp[10]) ? node808 : node803;
											assign node803 = (inp[11]) ? node805 : 11'b11011010001;
												assign node805 = (inp[3]) ? 11'b11100110011 : 11'b01110110101;
											assign node808 = (inp[3]) ? node812 : node809;
												assign node809 = (inp[11]) ? 11'b11011010011 : 11'b11011000001;
												assign node812 = (inp[11]) ? 11'b01011010011 : 11'b01000010011;
									assign node815 = (inp[3]) ? node827 : node816;
										assign node816 = (inp[10]) ? node824 : node817;
											assign node817 = (inp[11]) ? node821 : node818;
												assign node818 = (inp[9]) ? 11'b01001110110 : 11'b01111110100;
												assign node821 = (inp[9]) ? 11'b01110100100 : 11'b01101110110;
											assign node824 = (inp[11]) ? 11'b11101100000 : 11'b11110110010;
										assign node827 = (inp[10]) ? node831 : node828;
											assign node828 = (inp[11]) ? 11'b11001100000 : 11'b11100100010;
											assign node831 = (inp[11]) ? node835 : node832;
												assign node832 = (inp[9]) ? 11'b01000100000 : 11'b01111110010;
												assign node835 = (inp[9]) ? 11'b01010100000 : 11'b01000100000;
							assign node838 = (inp[5]) ? node894 : node839;
								assign node839 = (inp[4]) ? node867 : node840;
									assign node840 = (inp[10]) ? node856 : node841;
										assign node841 = (inp[3]) ? node849 : node842;
											assign node842 = (inp[11]) ? node846 : node843;
												assign node843 = (inp[9]) ? 11'b01100001001 : 11'b01101001011;
												assign node846 = (inp[9]) ? 11'b01011011000 : 11'b01111001010;
											assign node849 = (inp[9]) ? node853 : node850;
												assign node850 = (inp[11]) ? 11'b11100011010 : 11'b11101001011;
												assign node853 = (inp[11]) ? 11'b11011001110 : 11'b11101101110;
										assign node856 = (inp[11]) ? node862 : node857;
											assign node857 = (inp[9]) ? node859 : 11'b11110001011;
												assign node859 = (inp[3]) ? 11'b01110111110 : 11'b11111111110;
											assign node862 = (inp[3]) ? node864 : 11'b11100001000;
												assign node864 = (inp[9]) ? 11'b01100011100 : 11'b01110011100;
									assign node867 = (inp[10]) ? node879 : node868;
										assign node868 = (inp[3]) ? node876 : node869;
											assign node869 = (inp[9]) ? node873 : node870;
												assign node870 = (inp[11]) ? 11'b01110001100 : 11'b01100101100;
												assign node873 = (inp[11]) ? 11'b01100111100 : 11'b01010101110;
											assign node876 = (inp[9]) ? 11'b11110111000 : 11'b11100101100;
										assign node879 = (inp[3]) ? node887 : node880;
											assign node880 = (inp[9]) ? node884 : node881;
												assign node881 = (inp[11]) ? 11'b11011111110 : 11'b11111111100;
												assign node884 = (inp[11]) ? 11'b11011111000 : 11'b11000101000;
											assign node887 = (inp[9]) ? node891 : node888;
												assign node888 = (inp[11]) ? 11'b01000111010 : 11'b01011101010;
												assign node891 = (inp[11]) ? 11'b01011111010 : 11'b01011011000;
								assign node894 = (inp[11]) ? node916 : node895;
									assign node895 = (inp[4]) ? node903 : node896;
										assign node896 = (inp[3]) ? node900 : node897;
											assign node897 = (inp[9]) ? 11'b01111011010 : 11'b01100111010;
											assign node900 = (inp[10]) ? 11'b01100001100 : 11'b11100011110;
										assign node903 = (inp[9]) ? node909 : node904;
											assign node904 = (inp[10]) ? 11'b01100011000 : node905;
												assign node905 = (inp[3]) ? 11'b11011011110 : 11'b01111011100;
											assign node909 = (inp[10]) ? node913 : node910;
												assign node910 = (inp[3]) ? 11'b11101100011 : 11'b01000011100;
												assign node913 = (inp[3]) ? 11'b01010100011 : 11'b11111110011;
									assign node916 = (inp[4]) ? node924 : node917;
										assign node917 = (inp[3]) ? node921 : node918;
											assign node918 = (inp[9]) ? 11'b01001100001 : 11'b11001110011;
											assign node921 = (inp[9]) ? 11'b11110110101 : 11'b11010100001;
										assign node924 = (inp[9]) ? node932 : node925;
											assign node925 = (inp[10]) ? node929 : node926;
												assign node926 = (inp[3]) ? 11'b11001010101 : 11'b01101010111;
												assign node929 = (inp[3]) ? 11'b01000000011 : 11'b11100000101;
											assign node932 = (inp[10]) ? 11'b01010000001 : 11'b11011000011;
						assign node935 = (inp[5]) ? node1021 : node936;
							assign node936 = (inp[10]) ? node982 : node937;
								assign node937 = (inp[3]) ? node957 : node938;
									assign node938 = (inp[4]) ? node946 : node939;
										assign node939 = (inp[9]) ? node943 : node940;
											assign node940 = (inp[6]) ? 11'b01110000001 : 11'b01101100001;
											assign node943 = (inp[11]) ? 11'b01001010011 : 11'b01110000010;
										assign node946 = (inp[11]) ? node952 : node947;
											assign node947 = (inp[6]) ? node949 : 11'b01000000100;
												assign node949 = (inp[9]) ? 11'b01001000101 : 11'b01011100101;
											assign node952 = (inp[6]) ? node954 : 11'b01011000111;
												assign node954 = (inp[9]) ? 11'b01111110110 : 11'b01001100100;
									assign node957 = (inp[4]) ? node971 : node958;
										assign node958 = (inp[9]) ? node964 : node959;
											assign node959 = (inp[11]) ? node961 : 11'b11011000010;
												assign node961 = (inp[6]) ? 11'b11011010001 : 11'b11010110001;
											assign node964 = (inp[6]) ? node968 : node965;
												assign node965 = (inp[11]) ? 11'b11010000111 : 11'b11000000100;
												assign node968 = (inp[11]) ? 11'b11000000101 : 11'b11010100111;
										assign node971 = (inp[9]) ? node979 : node972;
											assign node972 = (inp[6]) ? node976 : node973;
												assign node973 = (inp[11]) ? 11'b11101000101 : 11'b11110000100;
												assign node976 = (inp[11]) ? 11'b11110100100 : 11'b11100100111;
											assign node979 = (inp[11]) ? 11'b11111110000 : 11'b11111010001;
								assign node982 = (inp[3]) ? node1002 : node983;
									assign node983 = (inp[4]) ? node993 : node984;
										assign node984 = (inp[9]) ? node988 : node985;
											assign node985 = (inp[6]) ? 11'b11011000011 : 11'b11111000010;
											assign node988 = (inp[11]) ? node990 : 11'b11101010100;
												assign node990 = (inp[6]) ? 11'b11101110110 : 11'b11110010111;
										assign node993 = (inp[11]) ? node999 : node994;
											assign node994 = (inp[9]) ? 11'b11111100011 : node995;
												assign node995 = (inp[6]) ? 11'b11000110111 : 11'b11001110111;
											assign node999 = (inp[9]) ? 11'b11010110000 : 11'b11010110100;
									assign node1002 = (inp[4]) ? node1014 : node1003;
										assign node1003 = (inp[9]) ? node1007 : node1004;
											assign node1004 = (inp[6]) ? 11'b01100010111 : 11'b01111010101;
											assign node1007 = (inp[11]) ? node1011 : node1008;
												assign node1008 = (inp[6]) ? 11'b01011110101 : 11'b01011010100;
												assign node1011 = (inp[6]) ? 11'b01001110110 : 11'b01001010111;
										assign node1014 = (inp[11]) ? node1016 : 11'b01001110001;
											assign node1016 = (inp[6]) ? node1018 : 11'b01010110011;
												assign node1018 = (inp[9]) ? 11'b01010110010 : 11'b01011110010;
							assign node1021 = (inp[11]) ? node1073 : node1022;
								assign node1022 = (inp[6]) ? node1048 : node1023;
									assign node1023 = (inp[9]) ? node1037 : node1024;
										assign node1024 = (inp[4]) ? node1032 : node1025;
											assign node1025 = (inp[10]) ? node1029 : node1026;
												assign node1026 = (inp[3]) ? 11'b11111110011 : 11'b01101110011;
												assign node1029 = (inp[3]) ? 11'b01010110101 : 11'b11001110001;
											assign node1032 = (inp[3]) ? 11'b01101010001 : node1033;
												assign node1033 = (inp[10]) ? 11'b11111000111 : 11'b01010010111;
										assign node1037 = (inp[3]) ? node1043 : node1038;
											assign node1038 = (inp[4]) ? 11'b11011110000 : node1039;
												assign node1039 = (inp[10]) ? 11'b11111000101 : 11'b01110110001;
											assign node1043 = (inp[10]) ? 11'b01000000111 : node1044;
												assign node1044 = (inp[4]) ? 11'b11000000001 : 11'b11101010101;
									assign node1048 = (inp[4]) ? node1064 : node1049;
										assign node1049 = (inp[10]) ? node1057 : node1050;
											assign node1050 = (inp[3]) ? node1054 : node1051;
												assign node1051 = (inp[9]) ? 11'b01100010010 : 11'b01101010010;
												assign node1054 = (inp[9]) ? 11'b11100010100 : 11'b11101010000;
											assign node1057 = (inp[3]) ? node1061 : node1058;
												assign node1058 = (inp[9]) ? 11'b11101000100 : 11'b11001010000;
												assign node1061 = (inp[9]) ? 11'b01001000110 : 11'b01000010110;
										assign node1064 = (inp[10]) ? node1070 : node1065;
											assign node1065 = (inp[9]) ? 11'b11010100010 : node1066;
												assign node1066 = (inp[3]) ? 11'b11110010110 : 11'b01000010110;
											assign node1070 = (inp[3]) ? 11'b01111110000 : 11'b11110000100;
								assign node1073 = (inp[4]) ? node1099 : node1074;
									assign node1074 = (inp[9]) ? node1088 : node1075;
										assign node1075 = (inp[3]) ? node1083 : node1076;
											assign node1076 = (inp[10]) ? node1080 : node1077;
												assign node1077 = (inp[6]) ? 11'b01111110010 : 11'b01100110010;
												assign node1080 = (inp[6]) ? 11'b11111110000 : 11'b11101110010;
											assign node1083 = (inp[10]) ? node1085 : 11'b11111100010;
												assign node1085 = (inp[6]) ? 11'b01110100100 : 11'b01111100110;
										assign node1088 = (inp[10]) ? node1094 : node1089;
											assign node1089 = (inp[3]) ? 11'b11010110100 : node1090;
												assign node1090 = (inp[6]) ? 11'b01110100010 : 11'b01101100000;
											assign node1094 = (inp[3]) ? 11'b01011000100 : node1095;
												assign node1095 = (inp[6]) ? 11'b11011000100 : 11'b11000100100;
									assign node1099 = (inp[9]) ? node1109 : node1100;
										assign node1100 = (inp[10]) ? node1104 : node1101;
											assign node1101 = (inp[3]) ? 11'b11010010110 : 11'b01001010110;
											assign node1104 = (inp[3]) ? node1106 : 11'b11010000100;
												assign node1106 = (inp[6]) ? 11'b01011000000 : 11'b01011000010;
										assign node1109 = (inp[6]) ? node1113 : node1110;
											assign node1110 = (inp[3]) ? 11'b11011000000 : 11'b11000000000;
											assign node1113 = (inp[10]) ? node1115 : 11'b11010000010;
												assign node1115 = (inp[3]) ? 11'b01010000000 : 11'b11010000000;
					assign node1118 = (inp[3]) ? node1306 : node1119;
						assign node1119 = (inp[8]) ? node1213 : node1120;
							assign node1120 = (inp[6]) ? node1164 : node1121;
								assign node1121 = (inp[5]) ? node1141 : node1122;
									assign node1122 = (inp[4]) ? node1136 : node1123;
										assign node1123 = (inp[9]) ? node1129 : node1124;
											assign node1124 = (inp[11]) ? 11'b01010010001 : node1125;
												assign node1125 = (inp[10]) ? 11'b01010001100 : 11'b01001001000;
											assign node1129 = (inp[10]) ? node1133 : node1130;
												assign node1130 = (inp[11]) ? 11'b01110010101 : 11'b01001100101;
												assign node1133 = (inp[11]) ? 11'b01001100011 : 11'b01010110001;
										assign node1136 = (inp[9]) ? node1138 : 11'b01010110011;
											assign node1138 = (inp[10]) ? 11'b01110010011 : 11'b01101010111;
									assign node1141 = (inp[4]) ? node1151 : node1142;
										assign node1142 = (inp[10]) ? node1146 : node1143;
											assign node1143 = (inp[11]) ? 11'b01111010110 : 11'b01010000111;
											assign node1146 = (inp[9]) ? node1148 : 11'b01111000101;
												assign node1148 = (inp[11]) ? 11'b01110000000 : 11'b01101110010;
										assign node1151 = (inp[10]) ? node1159 : node1152;
											assign node1152 = (inp[9]) ? node1156 : node1153;
												assign node1153 = (inp[11]) ? 11'b01101110000 : 11'b01110100010;
												assign node1156 = (inp[11]) ? 11'b01111100110 : 11'b01101110100;
											assign node1159 = (inp[9]) ? node1161 : 11'b01010110100;
												assign node1161 = (inp[11]) ? 11'b01110100010 : 11'b01110110000;
								assign node1164 = (inp[5]) ? node1190 : node1165;
									assign node1165 = (inp[4]) ? node1175 : node1166;
										assign node1166 = (inp[9]) ? node1172 : node1167;
											assign node1167 = (inp[10]) ? node1169 : 11'b01011001001;
												assign node1169 = (inp[11]) ? 11'b01010011110 : 11'b01000001111;
											assign node1172 = (inp[11]) ? 11'b01010001000 : 11'b01001111000;
										assign node1175 = (inp[10]) ? node1183 : node1176;
											assign node1176 = (inp[9]) ? node1180 : node1177;
												assign node1177 = (inp[11]) ? 11'b01001111010 : 11'b01010101010;
												assign node1180 = (inp[11]) ? 11'b01010101110 : 11'b01110111100;
											assign node1183 = (inp[9]) ? node1187 : node1184;
												assign node1184 = (inp[11]) ? 11'b01111101100 : 11'b01001111100;
												assign node1187 = (inp[11]) ? 11'b01101101000 : 11'b01101011010;
									assign node1190 = (inp[11]) ? node1204 : node1191;
										assign node1191 = (inp[9]) ? node1197 : node1192;
											assign node1192 = (inp[10]) ? node1194 : 11'b01101001000;
												assign node1194 = (inp[4]) ? 11'b01000011110 : 11'b01101001110;
											assign node1197 = (inp[4]) ? node1201 : node1198;
												assign node1198 = (inp[10]) ? 11'b01110011010 : 11'b01001001100;
												assign node1201 = (inp[10]) ? 11'b01101110001 : 11'b01111110111;
										assign node1204 = (inp[4]) ? node1210 : node1205;
											assign node1205 = (inp[10]) ? 11'b01100100001 : node1206;
												assign node1206 = (inp[9]) ? 11'b01100110111 : 11'b01000110011;
											assign node1210 = (inp[9]) ? 11'b01101000101 : 11'b01110000111;
							assign node1213 = (inp[5]) ? node1265 : node1214;
								assign node1214 = (inp[9]) ? node1244 : node1215;
									assign node1215 = (inp[10]) ? node1231 : node1216;
										assign node1216 = (inp[11]) ? node1224 : node1217;
											assign node1217 = (inp[6]) ? node1221 : node1218;
												assign node1218 = (inp[4]) ? 11'b01100000010 : 11'b01100100000;
												assign node1221 = (inp[4]) ? 11'b01110100011 : 11'b01110000001;
											assign node1224 = (inp[6]) ? node1228 : node1225;
												assign node1225 = (inp[4]) ? 11'b01111010001 : 11'b01110110011;
												assign node1228 = (inp[4]) ? 11'b01100110010 : 11'b01101010011;
										assign node1231 = (inp[11]) ? node1239 : node1232;
											assign node1232 = (inp[4]) ? node1236 : node1233;
												assign node1233 = (inp[6]) ? 11'b01111100111 : 11'b01101000100;
												assign node1236 = (inp[6]) ? 11'b01110110101 : 11'b01101110101;
											assign node1239 = (inp[4]) ? 11'b01010000111 : node1240;
												assign node1240 = (inp[6]) ? 11'b01111010101 : 11'b01101010111;
									assign node1244 = (inp[10]) ? node1254 : node1245;
										assign node1245 = (inp[6]) ? node1251 : node1246;
											assign node1246 = (inp[4]) ? 11'b01111100111 : node1247;
												assign node1247 = (inp[11]) ? 11'b01001010101 : 11'b01110000100;
											assign node1251 = (inp[4]) ? 11'b01011010111 : 11'b01010010111;
										assign node1254 = (inp[11]) ? node1260 : node1255;
											assign node1255 = (inp[4]) ? node1257 : 11'b01111010010;
												assign node1257 = (inp[6]) ? 11'b01000010001 : 11'b01011110001;
											assign node1260 = (inp[6]) ? node1262 : 11'b01100000001;
												assign node1262 = (inp[4]) ? 11'b01000100000 : 11'b01111100000;
								assign node1265 = (inp[6]) ? node1285 : node1266;
									assign node1266 = (inp[11]) ? node1276 : node1267;
										assign node1267 = (inp[4]) ? node1273 : node1268;
											assign node1268 = (inp[9]) ? node1270 : 11'b01000100111;
												assign node1270 = (inp[10]) ? 11'b01001010001 : 11'b01101000111;
											assign node1273 = (inp[9]) ? 11'b01010010111 : 11'b01111010101;
										assign node1276 = (inp[4]) ? node1278 : 11'b01110110000;
											assign node1278 = (inp[9]) ? node1282 : node1279;
												assign node1279 = (inp[10]) ? 11'b01010000100 : 11'b01011010000;
												assign node1282 = (inp[10]) ? 11'b01010000010 : 11'b01011000110;
									assign node1285 = (inp[10]) ? node1295 : node1286;
										assign node1286 = (inp[9]) ? node1292 : node1287;
											assign node1287 = (inp[11]) ? 11'b01101110000 : node1288;
												assign node1288 = (inp[4]) ? 11'b01010000000 : 11'b01111000000;
											assign node1292 = (inp[11]) ? 11'b01001000100 : 11'b01001110100;
										assign node1295 = (inp[9]) ? node1301 : node1296;
											assign node1296 = (inp[4]) ? node1298 : 11'b01100110110;
												assign node1298 = (inp[11]) ? 11'b01001000110 : 11'b01101110110;
											assign node1301 = (inp[4]) ? 11'b01000110010 : node1302;
												assign node1302 = (inp[11]) ? 11'b01001000010 : 11'b01011010010;
						assign node1306 = (inp[10]) ? node1406 : node1307;
							assign node1307 = (inp[5]) ? node1357 : node1308;
								assign node1308 = (inp[4]) ? node1336 : node1309;
									assign node1309 = (inp[9]) ? node1321 : node1310;
										assign node1310 = (inp[8]) ? node1316 : node1311;
											assign node1311 = (inp[11]) ? 11'b01010001000 : node1312;
												assign node1312 = (inp[6]) ? 11'b01011001001 : 11'b01011001000;
											assign node1316 = (inp[11]) ? 11'b01000100011 : node1317;
												assign node1317 = (inp[6]) ? 11'b01011100001 : 11'b01011000000;
										assign node1321 = (inp[11]) ? node1329 : node1322;
											assign node1322 = (inp[8]) ? node1326 : node1323;
												assign node1323 = (inp[6]) ? 11'b01011111000 : 11'b01011110001;
												assign node1326 = (inp[6]) ? 11'b01000110001 : 11'b01001010010;
											assign node1329 = (inp[6]) ? node1333 : node1330;
												assign node1330 = (inp[8]) ? 11'b01110010001 : 11'b01111110001;
												assign node1333 = (inp[8]) ? 11'b01111110010 : 11'b01111011000;
									assign node1336 = (inp[9]) ? node1346 : node1337;
										assign node1337 = (inp[11]) ? node1341 : node1338;
											assign node1338 = (inp[6]) ? 11'b01010110001 : 11'b01011110011;
											assign node1341 = (inp[8]) ? 11'b01100110010 : node1342;
												assign node1342 = (inp[6]) ? 11'b01101111000 : 11'b01101110011;
										assign node1346 = (inp[8]) ? node1352 : node1347;
											assign node1347 = (inp[6]) ? node1349 : 11'b01111000011;
												assign node1349 = (inp[11]) ? 11'b01101101010 : 11'b01110101010;
											assign node1352 = (inp[6]) ? 11'b01101000001 : node1353;
												assign node1353 = (inp[11]) ? 11'b01101100001 : 11'b01100100001;
								assign node1357 = (inp[11]) ? node1381 : node1358;
									assign node1358 = (inp[8]) ? node1370 : node1359;
										assign node1359 = (inp[4]) ? node1365 : node1360;
											assign node1360 = (inp[6]) ? node1362 : 11'b01110000001;
												assign node1362 = (inp[9]) ? 11'b01110011000 : 11'b01110101010;
											assign node1365 = (inp[9]) ? node1367 : 11'b01100110000;
												assign node1367 = (inp[6]) ? 11'b01011100001 : 11'b01010100000;
										assign node1370 = (inp[4]) ? node1376 : node1371;
											assign node1371 = (inp[6]) ? node1373 : 11'b01111010011;
												assign node1373 = (inp[9]) ? 11'b01111010010 : 11'b01111000010;
											assign node1376 = (inp[6]) ? node1378 : 11'b01101010001;
												assign node1378 = (inp[9]) ? 11'b01000100010 : 11'b01100010010;
									assign node1381 = (inp[8]) ? node1397 : node1382;
										assign node1382 = (inp[9]) ? node1390 : node1383;
											assign node1383 = (inp[4]) ? node1387 : node1384;
												assign node1384 = (inp[6]) ? 11'b01111100011 : 11'b01110000010;
												assign node1387 = (inp[6]) ? 11'b01010010011 : 11'b01011110000;
											assign node1390 = (inp[6]) ? node1394 : node1391;
												assign node1391 = (inp[4]) ? 11'b01001100010 : 11'b01001010000;
												assign node1394 = (inp[4]) ? 11'b01001000011 : 11'b01000110011;
										assign node1397 = (inp[4]) ? node1403 : node1398;
											assign node1398 = (inp[9]) ? 11'b01000110010 : node1399;
												assign node1399 = (inp[6]) ? 11'b01101100010 : 11'b01100100000;
											assign node1403 = (inp[9]) ? 11'b01000000010 : 11'b01000010010;
							assign node1406 = (inp[9]) ? node1456 : node1407;
								assign node1407 = (inp[6]) ? node1431 : node1408;
									assign node1408 = (inp[5]) ? node1416 : node1409;
										assign node1409 = (inp[8]) ? node1411 : 11'b01010100011;
											assign node1411 = (inp[11]) ? 11'b01111000011 : node1412;
												assign node1412 = (inp[4]) ? 11'b01111100001 : 11'b01010000000;
										assign node1416 = (inp[11]) ? node1424 : node1417;
											assign node1417 = (inp[4]) ? node1421 : node1418;
												assign node1418 = (inp[8]) ? 11'b01010100011 : 11'b01001000011;
												assign node1421 = (inp[8]) ? 11'b01100000011 : 11'b01111100000;
											assign node1424 = (inp[4]) ? node1428 : node1425;
												assign node1425 = (inp[8]) ? 11'b01101100010 : 11'b01111000010;
												assign node1428 = (inp[8]) ? 11'b01001000010 : 11'b01010100010;
									assign node1431 = (inp[8]) ? node1445 : node1432;
										assign node1432 = (inp[5]) ? node1438 : node1433;
											assign node1433 = (inp[4]) ? 11'b01101101000 : node1434;
												assign node1434 = (inp[11]) ? 11'b01101001010 : 11'b01000001011;
											assign node1438 = (inp[11]) ? node1442 : node1439;
												assign node1439 = (inp[4]) ? 11'b01110001010 : 11'b01001001000;
												assign node1442 = (inp[4]) ? 11'b01010000001 : 11'b01111100001;
										assign node1445 = (inp[5]) ? node1451 : node1446;
											assign node1446 = (inp[11]) ? 11'b01110000001 : node1447;
												assign node1447 = (inp[4]) ? 11'b01111000011 : 11'b01010100011;
											assign node1451 = (inp[4]) ? node1453 : 11'b01100100000;
												assign node1453 = (inp[11]) ? 11'b01001000000 : 11'b01101100000;
								assign node1456 = (inp[4]) ? node1482 : node1457;
									assign node1457 = (inp[5]) ? node1473 : node1458;
										assign node1458 = (inp[11]) ? node1466 : node1459;
											assign node1459 = (inp[6]) ? node1463 : node1460;
												assign node1460 = (inp[8]) ? 11'b01000000010 : 11'b01000100011;
												assign node1463 = (inp[8]) ? 11'b01001100011 : 11'b01000101010;
											assign node1466 = (inp[8]) ? node1470 : node1467;
												assign node1467 = (inp[6]) ? 11'b01010001010 : 11'b01010100011;
												assign node1470 = (inp[6]) ? 11'b01011100000 : 11'b01011000001;
										assign node1473 = (inp[11]) ? node1479 : node1474;
											assign node1474 = (inp[6]) ? node1476 : 11'b01010000001;
												assign node1476 = (inp[8]) ? 11'b01011000000 : 11'b01011001010;
											assign node1479 = (inp[8]) ? 11'b01001000000 : 11'b01001000001;
									assign node1482 = (inp[5]) ? node1494 : node1483;
										assign node1483 = (inp[6]) ? node1489 : node1484;
											assign node1484 = (inp[8]) ? 11'b01001100011 : node1485;
												assign node1485 = (inp[11]) ? 11'b01001000001 : 11'b01000000001;
											assign node1489 = (inp[8]) ? 11'b01000100000 : node1490;
												assign node1490 = (inp[11]) ? 11'b01001101000 : 11'b01001001000;
										assign node1494 = (inp[11]) ? node1498 : node1495;
											assign node1495 = (inp[8]) ? 11'b01000100000 : 11'b01001000010;
											assign node1498 = (inp[8]) ? 11'b01000000000 : node1499;
												assign node1499 = (inp[6]) ? 11'b01000000001 : 11'b01000100000;
			assign node1503 = (inp[6]) ? node2255 : node1504;
				assign node1504 = (inp[2]) ? node1890 : node1505;
					assign node1505 = (inp[8]) ? node1699 : node1506;
						assign node1506 = (inp[5]) ? node1606 : node1507;
							assign node1507 = (inp[0]) ? node1561 : node1508;
								assign node1508 = (inp[10]) ? node1534 : node1509;
									assign node1509 = (inp[3]) ? node1523 : node1510;
										assign node1510 = (inp[4]) ? node1516 : node1511;
											assign node1511 = (inp[11]) ? node1513 : 11'b01010100011;
												assign node1513 = (inp[9]) ? 11'b01110010011 : 11'b01011000011;
											assign node1516 = (inp[11]) ? node1520 : node1517;
												assign node1517 = (inp[9]) ? 11'b01111000111 : 11'b01010100111;
												assign node1520 = (inp[9]) ? 11'b01001110111 : 11'b01000100111;
										assign node1523 = (inp[4]) ? node1529 : node1524;
											assign node1524 = (inp[11]) ? 11'b11111100111 : node1525;
												assign node1525 = (inp[9]) ? 11'b11011100111 : 11'b11011100011;
											assign node1529 = (inp[9]) ? 11'b11110010011 : node1530;
												assign node1530 = (inp[11]) ? 11'b11100100101 : 11'b11010100111;
									assign node1534 = (inp[4]) ? node1550 : node1535;
										assign node1535 = (inp[3]) ? node1543 : node1536;
											assign node1536 = (inp[9]) ? node1540 : node1537;
												assign node1537 = (inp[11]) ? 11'b11011000001 : 11'b11011100001;
												assign node1540 = (inp[11]) ? 11'b11111110101 : 11'b11011110101;
											assign node1543 = (inp[9]) ? node1547 : node1544;
												assign node1544 = (inp[11]) ? 11'b01010010101 : 11'b01010100101;
												assign node1547 = (inp[11]) ? 11'b01001110111 : 11'b01011110101;
										assign node1550 = (inp[11]) ? node1558 : node1551;
											assign node1551 = (inp[3]) ? node1555 : node1552;
												assign node1552 = (inp[9]) ? 11'b11110000001 : 11'b11010110101;
												assign node1555 = (inp[9]) ? 11'b01110010001 : 11'b01111000001;
											assign node1558 = (inp[3]) ? 11'b01100110011 : 11'b11100110001;
								assign node1561 = (inp[11]) ? node1579 : node1562;
									assign node1562 = (inp[4]) ? node1572 : node1563;
										assign node1563 = (inp[10]) ? node1567 : node1564;
											assign node1564 = (inp[9]) ? 11'b01000100101 : 11'b01001100001;
											assign node1567 = (inp[9]) ? node1569 : 11'b01000100111;
												assign node1569 = (inp[3]) ? 11'b01001100001 : 11'b01001110011;
										assign node1572 = (inp[3]) ? node1576 : node1573;
											assign node1573 = (inp[9]) ? 11'b01100010011 : 11'b01001010111;
											assign node1576 = (inp[10]) ? 11'b01000000001 : 11'b01000110011;
									assign node1579 = (inp[4]) ? node1595 : node1580;
										assign node1580 = (inp[9]) ? node1588 : node1581;
											assign node1581 = (inp[3]) ? node1585 : node1582;
												assign node1582 = (inp[10]) ? 11'b01000010111 : 11'b01001010001;
												assign node1585 = (inp[10]) ? 11'b01100000001 : 11'b01001000011;
											assign node1588 = (inp[10]) ? node1592 : node1589;
												assign node1589 = (inp[3]) ? 11'b01101110011 : 11'b01100010101;
												assign node1592 = (inp[3]) ? 11'b01011100001 : 11'b01011100011;
										assign node1595 = (inp[9]) ? node1601 : node1596;
											assign node1596 = (inp[10]) ? 11'b01111100111 : node1597;
												assign node1597 = (inp[3]) ? 11'b01110110011 : 11'b01010110001;
											assign node1601 = (inp[10]) ? node1603 : 11'b01011100101;
												assign node1603 = (inp[3]) ? 11'b01000100001 : 11'b01110100011;
							assign node1606 = (inp[11]) ? node1650 : node1607;
								assign node1607 = (inp[4]) ? node1629 : node1608;
									assign node1608 = (inp[0]) ? node1616 : node1609;
										assign node1609 = (inp[9]) ? node1613 : node1610;
											assign node1610 = (inp[10]) ? 11'b11111010001 : 11'b01011010011;
											assign node1613 = (inp[10]) ? 11'b01001000111 : 11'b11010010101;
										assign node1616 = (inp[10]) ? node1622 : node1617;
											assign node1617 = (inp[3]) ? 11'b01101010011 : node1618;
												assign node1618 = (inp[9]) ? 11'b01000000111 : 11'b01001000011;
											assign node1622 = (inp[3]) ? node1626 : node1623;
												assign node1623 = (inp[9]) ? 11'b01101010001 : 11'b01101000101;
												assign node1626 = (inp[9]) ? 11'b01011000001 : 11'b01000000001;
									assign node1629 = (inp[9]) ? node1641 : node1630;
										assign node1630 = (inp[0]) ? node1636 : node1631;
											assign node1631 = (inp[10]) ? node1633 : 11'b11100010101;
												assign node1633 = (inp[3]) ? 11'b01001110010 : 11'b11000000111;
											assign node1636 = (inp[10]) ? 11'b01111100000 : node1637;
												assign node1637 = (inp[3]) ? 11'b01110010011 : 11'b01110000011;
										assign node1641 = (inp[3]) ? node1645 : node1642;
											assign node1642 = (inp[10]) ? 11'b01100110000 : 11'b01101110100;
											assign node1645 = (inp[10]) ? 11'b01110100010 : node1646;
												assign node1646 = (inp[0]) ? 11'b01001100000 : 11'b11011100000;
								assign node1650 = (inp[4]) ? node1672 : node1651;
									assign node1651 = (inp[10]) ? node1667 : node1652;
										assign node1652 = (inp[9]) ? node1660 : node1653;
											assign node1653 = (inp[3]) ? node1657 : node1654;
												assign node1654 = (inp[0]) ? 11'b01001110010 : 11'b01010110000;
												assign node1657 = (inp[0]) ? 11'b01101100000 : 11'b11111100000;
											assign node1660 = (inp[3]) ? node1664 : node1661;
												assign node1661 = (inp[0]) ? 11'b01110110110 : 11'b01100100000;
												assign node1664 = (inp[0]) ? 11'b01010110000 : 11'b11000110110;
										assign node1667 = (inp[9]) ? node1669 : 11'b01011110100;
											assign node1669 = (inp[3]) ? 11'b01011000100 : 11'b01111000000;
									assign node1672 = (inp[9]) ? node1684 : node1673;
										assign node1673 = (inp[10]) ? node1677 : node1674;
											assign node1674 = (inp[3]) ? 11'b11110010110 : 11'b01011010100;
											assign node1677 = (inp[3]) ? node1681 : node1678;
												assign node1678 = (inp[0]) ? 11'b01100000110 : 11'b11010000110;
												assign node1681 = (inp[0]) ? 11'b01011000010 : 11'b01110000000;
										assign node1684 = (inp[10]) ? node1692 : node1685;
											assign node1685 = (inp[0]) ? node1689 : node1686;
												assign node1686 = (inp[3]) ? 11'b11101000010 : 11'b01001000110;
												assign node1689 = (inp[3]) ? 11'b01011000000 : 11'b01111000100;
											assign node1692 = (inp[3]) ? node1696 : node1693;
												assign node1693 = (inp[0]) ? 11'b01110000010 : 11'b11001000000;
												assign node1696 = (inp[0]) ? 11'b01000000000 : 11'b01100000000;
						assign node1699 = (inp[5]) ? node1791 : node1700;
							assign node1700 = (inp[11]) ? node1748 : node1701;
								assign node1701 = (inp[4]) ? node1727 : node1702;
									assign node1702 = (inp[10]) ? node1714 : node1703;
										assign node1703 = (inp[9]) ? node1711 : node1704;
											assign node1704 = (inp[3]) ? node1708 : node1705;
												assign node1705 = (inp[0]) ? 11'b01100000000 : 11'b01010000010;
												assign node1708 = (inp[0]) ? 11'b01001100010 : 11'b11111100010;
											assign node1711 = (inp[0]) ? 11'b01110100100 : 11'b11100100100;
										assign node1714 = (inp[9]) ? node1722 : node1715;
											assign node1715 = (inp[0]) ? node1719 : node1716;
												assign node1716 = (inp[3]) ? 11'b01111100100 : 11'b11011100000;
												assign node1719 = (inp[3]) ? 11'b01011100000 : 11'b01101100110;
											assign node1722 = (inp[0]) ? node1724 : 11'b01101110110;
												assign node1724 = (inp[3]) ? 11'b01001100000 : 11'b01111110010;
									assign node1727 = (inp[9]) ? node1737 : node1728;
										assign node1728 = (inp[3]) ? node1734 : node1729;
											assign node1729 = (inp[10]) ? 11'b01100110100 : node1730;
												assign node1730 = (inp[0]) ? 11'b01101100010 : 11'b01111100110;
											assign node1734 = (inp[0]) ? 11'b01000110010 : 11'b01000100010;
										assign node1737 = (inp[10]) ? node1741 : node1738;
											assign node1738 = (inp[3]) ? 11'b11001010000 : 11'b01011010110;
											assign node1741 = (inp[0]) ? node1745 : node1742;
												assign node1742 = (inp[3]) ? 11'b01110010010 : 11'b11011000010;
												assign node1745 = (inp[3]) ? 11'b01000000010 : 11'b01001010000;
								assign node1748 = (inp[4]) ? node1772 : node1749;
									assign node1749 = (inp[0]) ? node1759 : node1750;
										assign node1750 = (inp[10]) ? node1756 : node1751;
											assign node1751 = (inp[3]) ? node1753 : 11'b01101010000;
												assign node1753 = (inp[9]) ? 11'b11110000110 : 11'b11110010000;
											assign node1756 = (inp[3]) ? 11'b01110010100 : 11'b11010010110;
										assign node1759 = (inp[10]) ? node1767 : node1760;
											assign node1760 = (inp[9]) ? node1764 : node1761;
												assign node1761 = (inp[3]) ? 11'b01010000000 : 11'b01100010010;
												assign node1764 = (inp[3]) ? 11'b01100010000 : 11'b01001010100;
											assign node1767 = (inp[9]) ? 11'b00011101011 : node1768;
												assign node1768 = (inp[3]) ? 11'b01111000010 : 11'b01111010100;
									assign node1772 = (inp[0]) ? node1786 : node1773;
										assign node1773 = (inp[10]) ? node1781 : node1774;
											assign node1774 = (inp[9]) ? node1778 : node1775;
												assign node1775 = (inp[3]) ? 11'b10001101111 : 11'b00101101111;
												assign node1778 = (inp[3]) ? 11'b10000111001 : 11'b00010111111;
											assign node1781 = (inp[3]) ? 11'b00101111011 : node1782;
												assign node1782 = (inp[9]) ? 11'b10101111001 : 11'b10101111101;
										assign node1786 = (inp[10]) ? 11'b00000101001 : node1787;
											assign node1787 = (inp[9]) ? 11'b00100101101 : 11'b00111111001;
							assign node1791 = (inp[0]) ? node1839 : node1792;
								assign node1792 = (inp[4]) ? node1814 : node1793;
									assign node1793 = (inp[9]) ? node1807 : node1794;
										assign node1794 = (inp[11]) ? node1800 : node1795;
											assign node1795 = (inp[10]) ? 11'b10110111001 : node1796;
												assign node1796 = (inp[3]) ? 11'b10010111001 : 11'b00010111011;
											assign node1800 = (inp[3]) ? node1804 : node1801;
												assign node1801 = (inp[10]) ? 11'b10000111001 : 11'b00011111011;
												assign node1804 = (inp[10]) ? 11'b00010101111 : 11'b10001101001;
										assign node1807 = (inp[10]) ? node1811 : node1808;
											assign node1808 = (inp[11]) ? 11'b10111111101 : 11'b10011011101;
											assign node1811 = (inp[11]) ? 11'b00100101111 : 11'b00110001111;
									assign node1814 = (inp[9]) ? node1826 : node1815;
										assign node1815 = (inp[11]) ? node1823 : node1816;
											assign node1816 = (inp[10]) ? node1820 : node1817;
												assign node1817 = (inp[3]) ? 11'b10001011111 : 11'b00100011101;
												assign node1820 = (inp[3]) ? 11'b00011011001 : 11'b10011001111;
											assign node1823 = (inp[3]) ? 11'b00101001001 : 11'b10101001111;
										assign node1826 = (inp[10]) ? node1832 : node1827;
											assign node1827 = (inp[3]) ? node1829 : 11'b00111001101;
												assign node1829 = (inp[11]) ? 11'b10110001011 : 11'b10100001011;
											assign node1832 = (inp[3]) ? node1836 : node1833;
												assign node1833 = (inp[11]) ? 11'b10100001001 : 11'b10100011001;
												assign node1836 = (inp[11]) ? 11'b00100001001 : 11'b00111101001;
								assign node1839 = (inp[3]) ? node1871 : node1840;
									assign node1840 = (inp[4]) ? node1856 : node1841;
										assign node1841 = (inp[10]) ? node1849 : node1842;
											assign node1842 = (inp[11]) ? node1846 : node1843;
												assign node1843 = (inp[9]) ? 11'b00111001111 : 11'b00100101011;
												assign node1846 = (inp[9]) ? 11'b00001111111 : 11'b00101111001;
											assign node1849 = (inp[9]) ? node1853 : node1850;
												assign node1850 = (inp[11]) ? 11'b00110111111 : 11'b00010101101;
												assign node1853 = (inp[11]) ? 11'b00011101001 : 11'b00000011001;
										assign node1856 = (inp[11]) ? node1864 : node1857;
											assign node1857 = (inp[10]) ? node1861 : node1858;
												assign node1858 = (inp[9]) ? 11'b00010011101 : 11'b00011001011;
												assign node1861 = (inp[9]) ? 11'b00001111011 : 11'b00101011111;
											assign node1864 = (inp[10]) ? node1868 : node1865;
												assign node1865 = (inp[9]) ? 11'b00001001101 : 11'b00000111011;
												assign node1868 = (inp[9]) ? 11'b00010001011 : 11'b00011001101;
									assign node1871 = (inp[11]) ? node1885 : node1872;
										assign node1872 = (inp[10]) ? node1878 : node1873;
											assign node1873 = (inp[4]) ? 11'b00111011001 : node1874;
												assign node1874 = (inp[9]) ? 11'b00101011001 : 11'b00100101011;
											assign node1878 = (inp[4]) ? node1882 : node1879;
												assign node1879 = (inp[9]) ? 11'b00010001011 : 11'b00011001001;
												assign node1882 = (inp[9]) ? 11'b00001101001 : 11'b00100001011;
										assign node1885 = (inp[10]) ? 11'b00100101001 : node1886;
											assign node1886 = (inp[9]) ? 11'b00010001001 : 11'b00010111001;
					assign node1890 = (inp[0]) ? node2072 : node1891;
						assign node1891 = (inp[8]) ? node1975 : node1892;
							assign node1892 = (inp[10]) ? node1934 : node1893;
								assign node1893 = (inp[3]) ? node1915 : node1894;
									assign node1894 = (inp[4]) ? node1904 : node1895;
										assign node1895 = (inp[11]) ? node1901 : node1896;
											assign node1896 = (inp[5]) ? node1898 : 11'b00111001011;
												assign node1898 = (inp[9]) ? 11'b00111111000 : 11'b00110111010;
											assign node1901 = (inp[9]) ? 11'b00000001010 : 11'b00110101010;
										assign node1904 = (inp[11]) ? node1912 : node1905;
											assign node1905 = (inp[5]) ? node1909 : node1906;
												assign node1906 = (inp[9]) ? 11'b00011101100 : 11'b00111101100;
												assign node1909 = (inp[9]) ? 11'b00010011110 : 11'b00100111110;
											assign node1912 = (inp[5]) ? 11'b00101101101 : 11'b00100011110;
									assign node1915 = (inp[4]) ? node1923 : node1916;
										assign node1916 = (inp[11]) ? 11'b10100111000 : node1917;
											assign node1917 = (inp[5]) ? 11'b10110111000 : node1918;
												assign node1918 = (inp[9]) ? 11'b10110001101 : 11'b10111001011;
										assign node1923 = (inp[9]) ? node1929 : node1924;
											assign node1924 = (inp[5]) ? 11'b10011011110 : node1925;
												assign node1925 = (inp[11]) ? 11'b10011001110 : 11'b10110101100;
											assign node1929 = (inp[5]) ? node1931 : 11'b10001111010;
												assign node1931 = (inp[11]) ? 11'b10011101011 : 11'b10110001000;
								assign node1934 = (inp[3]) ? node1956 : node1935;
									assign node1935 = (inp[11]) ? node1945 : node1936;
										assign node1936 = (inp[5]) ? node1942 : node1937;
											assign node1937 = (inp[9]) ? node1939 : 11'b10100111110;
												assign node1939 = (inp[4]) ? 11'b10001101000 : 11'b10101111110;
											assign node1942 = (inp[4]) ? 11'b10100011010 : 11'b10000111010;
										assign node1945 = (inp[9]) ? node1951 : node1946;
											assign node1946 = (inp[4]) ? 11'b10100101111 : node1947;
												assign node1947 = (inp[5]) ? 11'b10010011010 : 11'b10101001000;
											assign node1951 = (inp[5]) ? 11'b10001101101 : node1952;
												assign node1952 = (inp[4]) ? 11'b10001111000 : 11'b10010011110;
									assign node1956 = (inp[4]) ? node1966 : node1957;
										assign node1957 = (inp[5]) ? node1963 : node1958;
											assign node1958 = (inp[9]) ? 11'b00101111110 : node1959;
												assign node1959 = (inp[11]) ? 11'b00111011110 : 11'b00100001111;
											assign node1963 = (inp[9]) ? 11'b00110101100 : 11'b00011111110;
										assign node1966 = (inp[11]) ? node1970 : node1967;
											assign node1967 = (inp[9]) ? 11'b00011001010 : 11'b00101011010;
											assign node1970 = (inp[5]) ? node1972 : 11'b00001111010;
												assign node1972 = (inp[9]) ? 11'b00000101001 : 11'b00011101011;
							assign node1975 = (inp[5]) ? node2027 : node1976;
								assign node1976 = (inp[11]) ? node2004 : node1977;
									assign node1977 = (inp[10]) ? node1989 : node1978;
										assign node1978 = (inp[3]) ? node1986 : node1979;
											assign node1979 = (inp[4]) ? node1983 : node1980;
												assign node1980 = (inp[9]) ? 11'b00101001001 : 11'b00110101011;
												assign node1983 = (inp[9]) ? 11'b00000001111 : 11'b00011001101;
											assign node1986 = (inp[9]) ? 11'b10010001101 : 11'b10101001111;
										assign node1989 = (inp[3]) ? node1997 : node1990;
											assign node1990 = (inp[9]) ? node1994 : node1991;
												assign node1991 = (inp[4]) ? 11'b10011011101 : 11'b10101001001;
												assign node1994 = (inp[4]) ? 11'b10101101011 : 11'b10110011111;
											assign node1997 = (inp[4]) ? node2001 : node1998;
												assign node1998 = (inp[9]) ? 11'b00000011101 : 11'b00011001111;
												assign node2001 = (inp[9]) ? 11'b00011111011 : 11'b00110001001;
									assign node2004 = (inp[4]) ? node2018 : node2005;
										assign node2005 = (inp[3]) ? node2013 : node2006;
											assign node2006 = (inp[10]) ? node2010 : node2007;
												assign node2007 = (inp[9]) ? 11'b00011111011 : 11'b00111101001;
												assign node2010 = (inp[9]) ? 11'b10101111101 : 11'b10010101011;
											assign node2013 = (inp[10]) ? 11'b00100111101 : node2014;
												assign node2014 = (inp[9]) ? 11'b10001101101 : 11'b10000111011;
										assign node2018 = (inp[10]) ? node2022 : node2019;
											assign node2019 = (inp[9]) ? 11'b00111011101 : 11'b10110101101;
											assign node2022 = (inp[9]) ? 11'b10010011001 : node2023;
												assign node2023 = (inp[3]) ? 11'b00011011001 : 11'b10001011111;
								assign node2027 = (inp[4]) ? node2047 : node2028;
									assign node2028 = (inp[9]) ? node2036 : node2029;
										assign node2029 = (inp[11]) ? node2033 : node2030;
											assign node2030 = (inp[3]) ? 11'b00001011101 : 11'b00111011011;
											assign node2033 = (inp[10]) ? 11'b10110111000 : 11'b00110111010;
										assign node2036 = (inp[10]) ? node2042 : node2037;
											assign node2037 = (inp[3]) ? node2039 : 11'b00111001000;
												assign node2039 = (inp[11]) ? 11'b10001011110 : 11'b10110011111;
											assign node2042 = (inp[3]) ? 11'b00011101100 : node2043;
												assign node2043 = (inp[11]) ? 11'b10010001110 : 11'b10100001101;
									assign node2047 = (inp[11]) ? node2059 : node2048;
										assign node2048 = (inp[9]) ? node2052 : node2049;
											assign node2049 = (inp[10]) ? 11'b10100101110 : 11'b10111111100;
											assign node2052 = (inp[3]) ? node2056 : node2053;
												assign node2053 = (inp[10]) ? 11'b10001111000 : 11'b00000111100;
												assign node2056 = (inp[10]) ? 11'b00011101000 : 11'b10011101010;
										assign node2059 = (inp[3]) ? node2065 : node2060;
											assign node2060 = (inp[10]) ? 11'b10011001100 : node2061;
												assign node2061 = (inp[9]) ? 11'b00011001100 : 11'b00010011110;
											assign node2065 = (inp[10]) ? node2069 : node2066;
												assign node2066 = (inp[9]) ? 11'b10000001010 : 11'b10000011100;
												assign node2069 = (inp[9]) ? 11'b00000001000 : 11'b00001001010;
						assign node2072 = (inp[3]) ? node2174 : node2073;
							assign node2073 = (inp[8]) ? node2123 : node2074;
								assign node2074 = (inp[5]) ? node2096 : node2075;
									assign node2075 = (inp[11]) ? node2085 : node2076;
										assign node2076 = (inp[10]) ? node2080 : node2077;
											assign node2077 = (inp[4]) ? 11'b00000101010 : 11'b00001001001;
											assign node2080 = (inp[9]) ? node2082 : 11'b00010111100;
												assign node2082 = (inp[4]) ? 11'b00110111010 : 11'b00011111000;
										assign node2085 = (inp[9]) ? node2091 : node2086;
											assign node2086 = (inp[10]) ? 11'b00001011100 : node2087;
												assign node2087 = (inp[4]) ? 11'b00011011010 : 11'b00010111000;
											assign node2091 = (inp[10]) ? 11'b00000001000 : node2092;
												assign node2092 = (inp[4]) ? 11'b00000001100 : 11'b00110011110;
									assign node2096 = (inp[9]) ? node2110 : node2097;
										assign node2097 = (inp[10]) ? node2103 : node2098;
											assign node2098 = (inp[4]) ? 11'b00100111011 : node2099;
												assign node2099 = (inp[11]) ? 11'b00011011010 : 11'b00000101010;
											assign node2103 = (inp[11]) ? node2107 : node2104;
												assign node2104 = (inp[4]) ? 11'b00011011110 : 11'b00110101100;
												assign node2107 = (inp[4]) ? 11'b00100101101 : 11'b00000011110;
										assign node2110 = (inp[10]) ? node2116 : node2111;
											assign node2111 = (inp[11]) ? node2113 : 11'b00011101110;
												assign node2113 = (inp[4]) ? 11'b00111101111 : 11'b00110011100;
											assign node2116 = (inp[11]) ? node2120 : node2117;
												assign node2117 = (inp[4]) ? 11'b00110011000 : 11'b00100111010;
												assign node2120 = (inp[4]) ? 11'b00110101011 : 11'b00111101011;
								assign node2123 = (inp[5]) ? node2151 : node2124;
									assign node2124 = (inp[4]) ? node2138 : node2125;
										assign node2125 = (inp[11]) ? node2131 : node2126;
											assign node2126 = (inp[9]) ? node2128 : 11'b00101001101;
												assign node2128 = (inp[10]) ? 11'b00110011001 : 11'b00110001111;
											assign node2131 = (inp[9]) ? node2135 : node2132;
												assign node2132 = (inp[10]) ? 11'b00100111111 : 11'b00110111011;
												assign node2135 = (inp[10]) ? 11'b00101101001 : 11'b00001111101;
										assign node2138 = (inp[10]) ? node2146 : node2139;
											assign node2139 = (inp[9]) ? node2143 : node2140;
												assign node2140 = (inp[11]) ? 11'b00110111011 : 11'b00101001001;
												assign node2143 = (inp[11]) ? 11'b00111001101 : 11'b00000011111;
											assign node2146 = (inp[11]) ? node2148 : 11'b00011111001;
												assign node2148 = (inp[9]) ? 11'b00010001011 : 11'b00011001101;
									assign node2151 = (inp[11]) ? node2165 : node2152;
										assign node2152 = (inp[4]) ? node2160 : node2153;
											assign node2153 = (inp[10]) ? node2157 : node2154;
												assign node2154 = (inp[9]) ? 11'b00100001101 : 11'b00101001011;
												assign node2157 = (inp[9]) ? 11'b00001111010 : 11'b00001001101;
											assign node2160 = (inp[9]) ? node2162 : 11'b00001101010;
												assign node2162 = (inp[10]) ? 11'b00011111010 : 11'b00011111110;
										assign node2165 = (inp[9]) ? node2169 : node2166;
											assign node2166 = (inp[4]) ? 11'b00010011000 : 11'b00110111100;
											assign node2169 = (inp[4]) ? node2171 : 11'b00011011110;
												assign node2171 = (inp[10]) ? 11'b00010001010 : 11'b00010001110;
							assign node2174 = (inp[8]) ? node2218 : node2175;
								assign node2175 = (inp[10]) ? node2197 : node2176;
									assign node2176 = (inp[11]) ? node2186 : node2177;
										assign node2177 = (inp[9]) ? node2179 : 11'b00110101010;
											assign node2179 = (inp[4]) ? node2183 : node2180;
												assign node2180 = (inp[5]) ? 11'b00111111000 : 11'b00011111010;
												assign node2183 = (inp[5]) ? 11'b00010001010 : 11'b00111101000;
										assign node2186 = (inp[5]) ? node2190 : node2187;
											assign node2187 = (inp[9]) ? 11'b00110011010 : 11'b00011001010;
											assign node2190 = (inp[9]) ? node2194 : node2191;
												assign node2191 = (inp[4]) ? 11'b00010111011 : 11'b00111001000;
												assign node2194 = (inp[4]) ? 11'b00001101001 : 11'b00001111011;
									assign node2197 = (inp[9]) ? node2207 : node2198;
										assign node2198 = (inp[11]) ? node2202 : node2199;
											assign node2199 = (inp[4]) ? 11'b00111001000 : 11'b00001101010;
											assign node2202 = (inp[4]) ? node2204 : 11'b00110001010;
												assign node2204 = (inp[5]) ? 11'b00011101011 : 11'b00010001010;
										assign node2207 = (inp[4]) ? node2213 : node2208;
											assign node2208 = (inp[11]) ? 11'b00011001010 : node2209;
												assign node2209 = (inp[5]) ? 11'b00010101010 : 11'b00001101010;
											assign node2213 = (inp[5]) ? 11'b00001001010 : node2214;
												assign node2214 = (inp[11]) ? 11'b00001101000 : 11'b00000101000;
								assign node2218 = (inp[5]) ? node2240 : node2219;
									assign node2219 = (inp[10]) ? node2229 : node2220;
										assign node2220 = (inp[11]) ? node2222 : 11'b00000011001;
											assign node2222 = (inp[9]) ? node2226 : node2223;
												assign node2223 = (inp[4]) ? 11'b00100111001 : 11'b00000101001;
												assign node2226 = (inp[4]) ? 11'b00100001011 : 11'b00111111011;
										assign node2229 = (inp[9]) ? node2237 : node2230;
											assign node2230 = (inp[11]) ? node2234 : node2231;
												assign node2231 = (inp[4]) ? 11'b00110001001 : 11'b00011001001;
												assign node2234 = (inp[4]) ? 11'b00001001011 : 11'b00111101011;
											assign node2237 = (inp[11]) ? 11'b00000001001 : 11'b00001101011;
									assign node2240 = (inp[9]) ? node2252 : node2241;
										assign node2241 = (inp[11]) ? node2245 : node2242;
											assign node2242 = (inp[10]) ? 11'b00100101010 : 11'b00111001011;
											assign node2245 = (inp[4]) ? node2249 : node2246;
												assign node2246 = (inp[10]) ? 11'b00101001010 : 11'b00100101010;
												assign node2249 = (inp[10]) ? 11'b00001001010 : 11'b00001011010;
										assign node2252 = (inp[10]) ? 11'b00000001000 : 11'b00001011000;
				assign node2255 = (inp[8]) ? node2651 : node2256;
					assign node2256 = (inp[5]) ? node2462 : node2257;
						assign node2257 = (inp[2]) ? node2355 : node2258;
							assign node2258 = (inp[4]) ? node2306 : node2259;
								assign node2259 = (inp[11]) ? node2285 : node2260;
									assign node2260 = (inp[3]) ? node2274 : node2261;
										assign node2261 = (inp[10]) ? node2269 : node2262;
											assign node2262 = (inp[9]) ? node2266 : node2263;
												assign node2263 = (inp[0]) ? 11'b00011101000 : 11'b00011101010;
												assign node2266 = (inp[0]) ? 11'b00010101110 : 11'b00010101000;
											assign node2269 = (inp[9]) ? 11'b10011111110 : node2270;
												assign node2270 = (inp[0]) ? 11'b00011101100 : 11'b10011101000;
										assign node2274 = (inp[0]) ? node2280 : node2275;
											assign node2275 = (inp[10]) ? 11'b00001111100 : node2276;
												assign node2276 = (inp[9]) ? 11'b10000101110 : 11'b10001101000;
											assign node2280 = (inp[9]) ? node2282 : 11'b00000101010;
												assign node2282 = (inp[10]) ? 11'b00001101000 : 11'b00000111000;
									assign node2285 = (inp[0]) ? node2295 : node2286;
										assign node2286 = (inp[3]) ? node2288 : 11'b10000001010;
											assign node2288 = (inp[10]) ? node2292 : node2289;
												assign node2289 = (inp[9]) ? 11'b10111001110 : 11'b10010011000;
												assign node2292 = (inp[9]) ? 11'b00010011100 : 11'b00011011110;
										assign node2295 = (inp[3]) ? node2299 : node2296;
											assign node2296 = (inp[10]) ? 11'b00010011100 : 11'b00010011000;
											assign node2299 = (inp[9]) ? node2303 : node2300;
												assign node2300 = (inp[10]) ? 11'b00101001010 : 11'b00000001010;
												assign node2303 = (inp[10]) ? 11'b00010001000 : 11'b00101011000;
								assign node2306 = (inp[11]) ? node2330 : node2307;
									assign node2307 = (inp[9]) ? node2317 : node2308;
										assign node2308 = (inp[3]) ? node2314 : node2309;
											assign node2309 = (inp[10]) ? node2311 : 11'b00011101110;
												assign node2311 = (inp[0]) ? 11'b00010111100 : 11'b10010111100;
											assign node2314 = (inp[10]) ? 11'b00100101010 : 11'b10001101100;
										assign node2317 = (inp[3]) ? node2323 : node2318;
											assign node2318 = (inp[0]) ? node2320 : 11'b10111001010;
												assign node2320 = (inp[10]) ? 11'b00111011010 : 11'b00111011110;
											assign node2323 = (inp[0]) ? node2327 : node2324;
												assign node2324 = (inp[10]) ? 11'b00101011000 : 11'b10101011010;
												assign node2327 = (inp[10]) ? 11'b00001001000 : 11'b00101001000;
									assign node2330 = (inp[0]) ? node2342 : node2331;
										assign node2331 = (inp[10]) ? node2335 : node2332;
											assign node2332 = (inp[9]) ? 11'b10000110011 : 11'b10110001100;
											assign node2335 = (inp[9]) ? node2339 : node2336;
												assign node2336 = (inp[3]) ? 11'b00111110011 : 11'b10101110111;
												assign node2339 = (inp[3]) ? 11'b00100110011 : 11'b10110110001;
										assign node2342 = (inp[3]) ? node2350 : node2343;
											assign node2343 = (inp[10]) ? node2347 : node2344;
												assign node2344 = (inp[9]) ? 11'b00001100101 : 11'b00000011010;
												assign node2347 = (inp[9]) ? 11'b00100100011 : 11'b00101100101;
											assign node2350 = (inp[9]) ? 11'b00110100001 : node2351;
												assign node2351 = (inp[10]) ? 11'b00011100011 : 11'b00111110011;
							assign node2355 = (inp[0]) ? node2409 : node2356;
								assign node2356 = (inp[4]) ? node2380 : node2357;
									assign node2357 = (inp[10]) ? node2367 : node2358;
										assign node2358 = (inp[11]) ? 11'b00101100011 : node2359;
											assign node2359 = (inp[9]) ? node2363 : node2360;
												assign node2360 = (inp[3]) ? 11'b10111000000 : 11'b00111000010;
												assign node2363 = (inp[3]) ? 11'b10110000110 : 11'b00110000000;
										assign node2367 = (inp[3]) ? node2373 : node2368;
											assign node2368 = (inp[11]) ? 11'b10011010101 : node2369;
												assign node2369 = (inp[9]) ? 11'b10100010100 : 11'b10101000010;
											assign node2373 = (inp[9]) ? node2377 : node2374;
												assign node2374 = (inp[11]) ? 11'b00100110101 : 11'b00101000100;
												assign node2377 = (inp[11]) ? 11'b00111010111 : 11'b00101110111;
									assign node2380 = (inp[11]) ? node2394 : node2381;
										assign node2381 = (inp[9]) ? node2389 : node2382;
											assign node2382 = (inp[3]) ? node2386 : node2383;
												assign node2383 = (inp[10]) ? 11'b10101110101 : 11'b00111100101;
												assign node2386 = (inp[10]) ? 11'b00000100011 : 11'b10111100111;
											assign node2389 = (inp[3]) ? node2391 : 11'b00000100101;
												assign node2391 = (inp[10]) ? 11'b00001110001 : 11'b10010110001;
										assign node2394 = (inp[3]) ? node2402 : node2395;
											assign node2395 = (inp[10]) ? node2399 : node2396;
												assign node2396 = (inp[9]) ? 11'b00110010101 : 11'b00101000101;
												assign node2399 = (inp[9]) ? 11'b10001010001 : 11'b10000010101;
											assign node2402 = (inp[9]) ? node2406 : node2403;
												assign node2403 = (inp[10]) ? 11'b00010010011 : 11'b10000000111;
												assign node2406 = (inp[10]) ? 11'b00001010011 : 11'b10101010011;
								assign node2409 = (inp[11]) ? node2437 : node2410;
									assign node2410 = (inp[4]) ? node2422 : node2411;
										assign node2411 = (inp[3]) ? node2417 : node2412;
											assign node2412 = (inp[9]) ? 11'b00000010000 : node2413;
												assign node2413 = (inp[10]) ? 11'b00001000100 : 11'b00011000000;
											assign node2417 = (inp[9]) ? 11'b00001100011 : node2418;
												assign node2418 = (inp[10]) ? 11'b00000000010 : 11'b00011000010;
										assign node2422 = (inp[3]) ? node2430 : node2423;
											assign node2423 = (inp[9]) ? node2427 : node2424;
												assign node2424 = (inp[10]) ? 11'b00000110111 : 11'b00011100011;
												assign node2427 = (inp[10]) ? 11'b00101110011 : 11'b00110110111;
											assign node2430 = (inp[10]) ? node2434 : node2431;
												assign node2431 = (inp[9]) ? 11'b00110100001 : 11'b00011110001;
												assign node2434 = (inp[9]) ? 11'b00001100001 : 11'b00100100001;
									assign node2437 = (inp[10]) ? node2451 : node2438;
										assign node2438 = (inp[3]) ? node2444 : node2439;
											assign node2439 = (inp[9]) ? 11'b00100110101 : node2440;
												assign node2440 = (inp[4]) ? 11'b00001010001 : 11'b00001110011;
											assign node2444 = (inp[4]) ? node2448 : node2445;
												assign node2445 = (inp[9]) ? 11'b00111010011 : 11'b00010100011;
												assign node2448 = (inp[9]) ? 11'b00101000001 : 11'b00100010011;
										assign node2451 = (inp[9]) ? node2457 : node2452;
											assign node2452 = (inp[4]) ? node2454 : 11'b00100100011;
												assign node2454 = (inp[3]) ? 11'b00010000001 : 11'b00110000111;
											assign node2457 = (inp[4]) ? node2459 : 11'b00011000001;
												assign node2459 = (inp[3]) ? 11'b00001000001 : 11'b00101000011;
						assign node2462 = (inp[0]) ? node2556 : node2463;
							assign node2463 = (inp[11]) ? node2513 : node2464;
								assign node2464 = (inp[10]) ? node2486 : node2465;
									assign node2465 = (inp[3]) ? node2477 : node2466;
										assign node2466 = (inp[4]) ? node2472 : node2467;
											assign node2467 = (inp[2]) ? 11'b00110010011 : node2468;
												assign node2468 = (inp[9]) ? 11'b00000110011 : 11'b00011110011;
											assign node2472 = (inp[2]) ? node2474 : 11'b00110010111;
												assign node2474 = (inp[9]) ? 11'b00011110101 : 11'b00100110111;
										assign node2477 = (inp[9]) ? node2483 : node2478;
											assign node2478 = (inp[4]) ? 11'b10000110101 : node2479;
												assign node2479 = (inp[2]) ? 11'b10110010001 : 11'b10001110001;
											assign node2483 = (inp[2]) ? 11'b10111110101 : 11'b10010110111;
									assign node2486 = (inp[3]) ? node2500 : node2487;
										assign node2487 = (inp[9]) ? node2495 : node2488;
											assign node2488 = (inp[4]) ? node2492 : node2489;
												assign node2489 = (inp[2]) ? 11'b10010010011 : 11'b10111110011;
												assign node2492 = (inp[2]) ? 11'b10100100111 : 11'b10010000111;
											assign node2495 = (inp[4]) ? node2497 : 11'b10100100101;
												assign node2497 = (inp[2]) ? 11'b10101110001 : 11'b10011010001;
										assign node2500 = (inp[4]) ? node2506 : node2501;
											assign node2501 = (inp[9]) ? 11'b00111100101 : node2502;
												assign node2502 = (inp[2]) ? 11'b00000010101 : 11'b00101110101;
											assign node2506 = (inp[2]) ? node2510 : node2507;
												assign node2507 = (inp[9]) ? 11'b00101000011 : 11'b00000010001;
												assign node2510 = (inp[9]) ? 11'b00000100011 : 11'b00111110011;
								assign node2513 = (inp[9]) ? node2533 : node2514;
									assign node2514 = (inp[3]) ? node2520 : node2515;
										assign node2515 = (inp[10]) ? node2517 : 11'b00001010001;
											assign node2517 = (inp[2]) ? 11'b10010110001 : 11'b10100010001;
										assign node2520 = (inp[10]) ? node2526 : node2521;
											assign node2521 = (inp[4]) ? 11'b10100110111 : node2522;
												assign node2522 = (inp[2]) ? 11'b10000100011 : 11'b10110000011;
											assign node2526 = (inp[4]) ? node2530 : node2527;
												assign node2527 = (inp[2]) ? 11'b00111000111 : 11'b00010000101;
												assign node2530 = (inp[2]) ? 11'b00011000001 : 11'b00111100011;
									assign node2533 = (inp[2]) ? node2543 : node2534;
										assign node2534 = (inp[4]) ? node2540 : node2535;
											assign node2535 = (inp[3]) ? 11'b00001100101 : node2536;
												assign node2536 = (inp[10]) ? 11'b10111100111 : 11'b00101100011;
											assign node2540 = (inp[10]) ? 11'b00100100001 : 11'b10111100001;
										assign node2543 = (inp[10]) ? node2549 : node2544;
											assign node2544 = (inp[3]) ? 11'b10101010111 : node2545;
												assign node2545 = (inp[4]) ? 11'b00101000111 : 11'b00011000001;
											assign node2549 = (inp[4]) ? node2553 : node2550;
												assign node2550 = (inp[3]) ? 11'b00100000111 : 11'b10001000101;
												assign node2553 = (inp[3]) ? 11'b00000000001 : 11'b10100000011;
							assign node2556 = (inp[3]) ? node2608 : node2557;
								assign node2557 = (inp[9]) ? node2585 : node2558;
									assign node2558 = (inp[10]) ? node2572 : node2559;
										assign node2559 = (inp[4]) ? node2567 : node2560;
											assign node2560 = (inp[11]) ? node2564 : node2561;
												assign node2561 = (inp[2]) ? 11'b00010000011 : 11'b00011100011;
												assign node2564 = (inp[2]) ? 11'b00000110001 : 11'b00010010011;
											assign node2567 = (inp[11]) ? node2569 : 11'b00100100001;
												assign node2569 = (inp[2]) ? 11'b00110010011 : 11'b00110110001;
										assign node2572 = (inp[11]) ? node2580 : node2573;
											assign node2573 = (inp[4]) ? node2577 : node2574;
												assign node2574 = (inp[2]) ? 11'b00100000111 : 11'b00111100101;
												assign node2577 = (inp[2]) ? 11'b00000110101 : 11'b00000010111;
											assign node2580 = (inp[4]) ? node2582 : 11'b00011010111;
												assign node2582 = (inp[2]) ? 11'b00111000111 : 11'b00111100111;
									assign node2585 = (inp[10]) ? node2599 : node2586;
										assign node2586 = (inp[11]) ? node2592 : node2587;
											assign node2587 = (inp[4]) ? node2589 : 11'b00001100111;
												assign node2589 = (inp[2]) ? 11'b00111110101 : 11'b00100010101;
											assign node2592 = (inp[2]) ? node2596 : node2593;
												assign node2593 = (inp[4]) ? 11'b00101100111 : 11'b00101110111;
												assign node2596 = (inp[4]) ? 11'b00101000111 : 11'b00101010111;
										assign node2599 = (inp[11]) ? node2603 : node2600;
											assign node2600 = (inp[2]) ? 11'b00111110001 : 11'b00111010001;
											assign node2603 = (inp[2]) ? 11'b00100000011 : node2604;
												assign node2604 = (inp[4]) ? 11'b00100100011 : 11'b00101100001;
								assign node2608 = (inp[10]) ? node2628 : node2609;
									assign node2609 = (inp[11]) ? node2617 : node2610;
										assign node2610 = (inp[2]) ? node2614 : node2611;
											assign node2611 = (inp[4]) ? 11'b00111010001 : 11'b00101100001;
											assign node2614 = (inp[4]) ? 11'b00100110011 : 11'b00110000001;
										assign node2617 = (inp[2]) ? node2623 : node2618;
											assign node2618 = (inp[9]) ? node2620 : 11'b00000110011;
												assign node2620 = (inp[4]) ? 11'b00011100001 : 11'b00011110011;
											assign node2623 = (inp[9]) ? node2625 : 11'b00010010001;
												assign node2625 = (inp[4]) ? 11'b00001000001 : 11'b00001010001;
									assign node2628 = (inp[11]) ? node2640 : node2629;
										assign node2629 = (inp[4]) ? node2637 : node2630;
											assign node2630 = (inp[9]) ? node2634 : node2631;
												assign node2631 = (inp[2]) ? 11'b00000000001 : 11'b00000100011;
												assign node2634 = (inp[2]) ? 11'b00010100011 : 11'b00011000001;
											assign node2637 = (inp[9]) ? 11'b00000100011 : 11'b00110000011;
										assign node2640 = (inp[9]) ? node2648 : node2641;
											assign node2641 = (inp[4]) ? node2645 : node2642;
												assign node2642 = (inp[2]) ? 11'b00111000001 : 11'b00110000001;
												assign node2645 = (inp[2]) ? 11'b00011000001 : 11'b00011100001;
											assign node2648 = (inp[2]) ? 11'b00000000001 : 11'b00000100001;
					assign node2651 = (inp[0]) ? node2839 : node2652;
						assign node2652 = (inp[11]) ? node2754 : node2653;
							assign node2653 = (inp[2]) ? node2699 : node2654;
								assign node2654 = (inp[5]) ? node2678 : node2655;
									assign node2655 = (inp[10]) ? node2669 : node2656;
										assign node2656 = (inp[3]) ? node2662 : node2657;
											assign node2657 = (inp[4]) ? 11'b00111000111 : node2658;
												assign node2658 = (inp[9]) ? 11'b00001000001 : 11'b00010100011;
											assign node2662 = (inp[4]) ? node2666 : node2663;
												assign node2663 = (inp[9]) ? 11'b10110000111 : 11'b10100100001;
												assign node2666 = (inp[9]) ? 11'b10000010001 : 11'b10011000101;
										assign node2669 = (inp[9]) ? node2675 : node2670;
											assign node2670 = (inp[3]) ? 11'b00011000001 : node2671;
												assign node2671 = (inp[4]) ? 11'b10101010111 : 11'b10001000011;
											assign node2675 = (inp[4]) ? 11'b00101110010 : 11'b00100010111;
									assign node2678 = (inp[9]) ? node2690 : node2679;
										assign node2679 = (inp[3]) ? node2685 : node2680;
											assign node2680 = (inp[4]) ? 11'b00100010100 : node2681;
												assign node2681 = (inp[10]) ? 11'b10100010010 : 11'b00010010010;
											assign node2685 = (inp[4]) ? node2687 : 11'b00110010100;
												assign node2687 = (inp[10]) ? 11'b00011110010 : 11'b10000010110;
										assign node2690 = (inp[4]) ? node2694 : node2691;
											assign node2691 = (inp[10]) ? 11'b10001000110 : 11'b00011010010;
											assign node2694 = (inp[10]) ? 11'b10110110010 : node2695;
												assign node2695 = (inp[3]) ? 11'b10111100000 : 11'b00101110100;
								assign node2699 = (inp[9]) ? node2729 : node2700;
									assign node2700 = (inp[5]) ? node2714 : node2701;
										assign node2701 = (inp[10]) ? node2709 : node2702;
											assign node2702 = (inp[4]) ? node2706 : node2703;
												assign node2703 = (inp[3]) ? 11'b10010000001 : 11'b00110000011;
												assign node2706 = (inp[3]) ? 11'b10111100110 : 11'b00000100110;
											assign node2709 = (inp[4]) ? 11'b10011110100 : node2710;
												assign node2710 = (inp[3]) ? 11'b00011100100 : 11'b10111100010;
										assign node2714 = (inp[3]) ? node2722 : node2715;
											assign node2715 = (inp[10]) ? node2719 : node2716;
												assign node2716 = (inp[4]) ? 11'b00011110110 : 11'b00111110010;
												assign node2719 = (inp[4]) ? 11'b10101100110 : 11'b10011110010;
											assign node2722 = (inp[10]) ? node2726 : node2723;
												assign node2723 = (inp[4]) ? 11'b10101110100 : 11'b10111110000;
												assign node2726 = (inp[4]) ? 11'b00101110000 : 11'b00011110100;
									assign node2729 = (inp[4]) ? node2741 : node2730;
										assign node2730 = (inp[3]) ? node2738 : node2731;
											assign node2731 = (inp[10]) ? node2735 : node2732;
												assign node2732 = (inp[5]) ? 11'b00110110010 : 11'b00101100010;
												assign node2735 = (inp[5]) ? 11'b10110100110 : 11'b10100110110;
											assign node2738 = (inp[10]) ? 11'b00000110100 : 11'b10110110100;
										assign node2741 = (inp[3]) ? node2747 : node2742;
											assign node2742 = (inp[5]) ? node2744 : 11'b00011100100;
												assign node2744 = (inp[10]) ? 11'b10000110010 : 11'b00000110110;
											assign node2747 = (inp[5]) ? node2751 : node2748;
												assign node2748 = (inp[10]) ? 11'b00000110010 : 11'b10100110010;
												assign node2751 = (inp[10]) ? 11'b00000100000 : 11'b10000100000;
							assign node2754 = (inp[2]) ? node2800 : node2755;
								assign node2755 = (inp[5]) ? node2781 : node2756;
									assign node2756 = (inp[9]) ? node2768 : node2757;
										assign node2757 = (inp[10]) ? node2765 : node2758;
											assign node2758 = (inp[3]) ? node2762 : node2759;
												assign node2759 = (inp[4]) ? 11'b00101100110 : 11'b00001100000;
												assign node2762 = (inp[4]) ? 11'b10001100100 : 11'b10111110010;
											assign node2765 = (inp[3]) ? 11'b00100110010 : 11'b10110110100;
										assign node2768 = (inp[4]) ? node2774 : node2769;
											assign node2769 = (inp[10]) ? node2771 : 11'b00110110010;
												assign node2771 = (inp[3]) ? 11'b00111110100 : 11'b10001110110;
											assign node2774 = (inp[10]) ? node2778 : node2775;
												assign node2775 = (inp[3]) ? 11'b10011010010 : 11'b00000110100;
												assign node2778 = (inp[3]) ? 11'b00101010010 : 11'b10101010000;
									assign node2781 = (inp[10]) ? node2791 : node2782;
										assign node2782 = (inp[4]) ? node2786 : node2783;
											assign node2783 = (inp[3]) ? 11'b10110110110 : 11'b00001100010;
											assign node2786 = (inp[3]) ? 11'b10110000000 : node2787;
												assign node2787 = (inp[9]) ? 11'b00110000110 : 11'b00110110100;
										assign node2791 = (inp[4]) ? node2793 : 11'b00100100110;
											assign node2793 = (inp[9]) ? node2797 : node2794;
												assign node2794 = (inp[3]) ? 11'b00101000010 : 11'b10101000100;
												assign node2797 = (inp[3]) ? 11'b00100000000 : 11'b10100000010;
								assign node2800 = (inp[9]) ? node2824 : node2801;
									assign node2801 = (inp[4]) ? node2815 : node2802;
										assign node2802 = (inp[10]) ? node2810 : node2803;
											assign node2803 = (inp[3]) ? node2807 : node2804;
												assign node2804 = (inp[5]) ? 11'b00101010010 : 11'b00100100000;
												assign node2807 = (inp[5]) ? 11'b10101000000 : 11'b10001010010;
											assign node2810 = (inp[3]) ? node2812 : 11'b10001000000;
												assign node2812 = (inp[5]) ? 11'b00101000100 : 11'b00111010110;
										assign node2815 = (inp[3]) ? 11'b00001000000 : node2816;
											assign node2816 = (inp[10]) ? node2820 : node2817;
												assign node2817 = (inp[5]) ? 11'b00001010110 : 11'b00010000100;
												assign node2820 = (inp[5]) ? 11'b10001000110 : 11'b10001010100;
									assign node2824 = (inp[4]) ? node2830 : node2825;
										assign node2825 = (inp[5]) ? node2827 : 11'b00010010110;
											assign node2827 = (inp[10]) ? 11'b00000000100 : 11'b10000010100;
										assign node2830 = (inp[5]) ? node2836 : node2831;
											assign node2831 = (inp[10]) ? node2833 : 11'b10100010010;
												assign node2833 = (inp[3]) ? 11'b00000010010 : 11'b10000010000;
											assign node2836 = (inp[10]) ? 11'b10000000010 : 11'b00000000110;
						assign node2839 = (inp[9]) ? node2935 : node2840;
							assign node2840 = (inp[10]) ? node2890 : node2841;
								assign node2841 = (inp[11]) ? node2865 : node2842;
									assign node2842 = (inp[2]) ? node2856 : node2843;
										assign node2843 = (inp[5]) ? node2849 : node2844;
											assign node2844 = (inp[3]) ? node2846 : 11'b00110100001;
												assign node2846 = (inp[4]) ? 11'b00001010001 : 11'b00001000011;
											assign node2849 = (inp[3]) ? node2853 : node2850;
												assign node2850 = (inp[4]) ? 11'b00000000000 : 11'b00110000010;
												assign node2853 = (inp[4]) ? 11'b00110010000 : 11'b00100000000;
										assign node2856 = (inp[3]) ? node2862 : node2857;
											assign node2857 = (inp[5]) ? node2859 : 11'b00110100000;
												assign node2859 = (inp[4]) ? 11'b00011100010 : 11'b00111100010;
											assign node2862 = (inp[5]) ? 11'b00101110000 : 11'b00011110010;
									assign node2865 = (inp[2]) ? node2877 : node2866;
										assign node2866 = (inp[3]) ? node2872 : node2867;
											assign node2867 = (inp[4]) ? 11'b00101110000 : node2868;
												assign node2868 = (inp[5]) ? 11'b00110110000 : 11'b00111110010;
											assign node2872 = (inp[5]) ? 11'b00011010000 : node2873;
												assign node2873 = (inp[4]) ? 11'b00110110010 : 11'b00011100000;
										assign node2877 = (inp[3]) ? node2885 : node2878;
											assign node2878 = (inp[4]) ? node2882 : node2879;
												assign node2879 = (inp[5]) ? 11'b00101010010 : 11'b00100110000;
												assign node2882 = (inp[5]) ? 11'b00001010010 : 11'b00101010010;
											assign node2885 = (inp[5]) ? node2887 : 11'b00001000010;
												assign node2887 = (inp[4]) ? 11'b00001010000 : 11'b00101000000;
								assign node2890 = (inp[3]) ? node2912 : node2891;
									assign node2891 = (inp[5]) ? node2901 : node2892;
										assign node2892 = (inp[2]) ? node2896 : node2893;
											assign node2893 = (inp[11]) ? 11'b00010100100 : 11'b00111000101;
											assign node2896 = (inp[11]) ? 11'b00111010110 : node2897;
												assign node2897 = (inp[4]) ? 11'b00111110100 : 11'b00111100100;
										assign node2901 = (inp[11]) ? node2909 : node2902;
											assign node2902 = (inp[4]) ? node2906 : node2903;
												assign node2903 = (inp[2]) ? 11'b00011100110 : 11'b00000000110;
												assign node2906 = (inp[2]) ? 11'b00101110110 : 11'b00111110110;
											assign node2909 = (inp[4]) ? 11'b00001000110 : 11'b00101110100;
									assign node2912 = (inp[5]) ? node2924 : node2913;
										assign node2913 = (inp[11]) ? node2921 : node2914;
											assign node2914 = (inp[2]) ? node2918 : node2915;
												assign node2915 = (inp[4]) ? 11'b00110000011 : 11'b00011000011;
												assign node2918 = (inp[4]) ? 11'b00111100010 : 11'b00011100010;
											assign node2921 = (inp[2]) ? 11'b00111000000 : 11'b00110100000;
										assign node2924 = (inp[2]) ? node2928 : node2925;
											assign node2925 = (inp[4]) ? 11'b00101100000 : 11'b00101100010;
											assign node2928 = (inp[11]) ? node2932 : node2929;
												assign node2929 = (inp[4]) ? 11'b00101100000 : 11'b00011100000;
												assign node2932 = (inp[4]) ? 11'b00001000000 : 11'b00101000000;
							assign node2935 = (inp[10]) ? node2981 : node2936;
								assign node2936 = (inp[3]) ? node2962 : node2937;
									assign node2937 = (inp[11]) ? node2949 : node2938;
										assign node2938 = (inp[4]) ? node2946 : node2939;
											assign node2939 = (inp[2]) ? node2943 : node2940;
												assign node2940 = (inp[5]) ? 11'b00101000100 : 11'b00101000101;
												assign node2943 = (inp[5]) ? 11'b00110100110 : 11'b00101100100;
											assign node2946 = (inp[5]) ? 11'b00001110110 : 11'b00000010101;
										assign node2949 = (inp[4]) ? node2957 : node2950;
											assign node2950 = (inp[2]) ? node2954 : node2951;
												assign node2951 = (inp[5]) ? 11'b00011110100 : 11'b00010110110;
												assign node2954 = (inp[5]) ? 11'b00000010110 : 11'b00010010110;
											assign node2957 = (inp[5]) ? node2959 : 11'b00111000110;
												assign node2959 = (inp[2]) ? 11'b00000000110 : 11'b00010000110;
									assign node2962 = (inp[4]) ? node2974 : node2963;
										assign node2963 = (inp[5]) ? node2967 : node2964;
											assign node2964 = (inp[2]) ? 11'b00000110010 : 11'b00100110000;
											assign node2967 = (inp[11]) ? node2971 : node2968;
												assign node2968 = (inp[2]) ? 11'b00110110000 : 11'b00101010010;
												assign node2971 = (inp[2]) ? 11'b00000010000 : 11'b00010110010;
										assign node2974 = (inp[5]) ? node2976 : 11'b00111000000;
											assign node2976 = (inp[2]) ? node2978 : 11'b00010000000;
												assign node2978 = (inp[11]) ? 11'b00000000000 : 11'b00000100000;
								assign node2981 = (inp[11]) ? node3007 : node2982;
									assign node2982 = (inp[3]) ? node2998 : node2983;
										assign node2983 = (inp[2]) ? node2991 : node2984;
											assign node2984 = (inp[5]) ? node2988 : node2985;
												assign node2985 = (inp[4]) ? 11'b00010010001 : 11'b00100010011;
												assign node2988 = (inp[4]) ? 11'b00010110010 : 11'b00011010000;
											assign node2991 = (inp[5]) ? node2995 : node2992;
												assign node2992 = (inp[4]) ? 11'b00000110000 : 11'b00100110000;
												assign node2995 = (inp[4]) ? 11'b00000110010 : 11'b00010110010;
										assign node2998 = (inp[4]) ? node3004 : node2999;
											assign node2999 = (inp[5]) ? node3001 : 11'b00000000001;
												assign node3001 = (inp[2]) ? 11'b00010100000 : 11'b00010000010;
											assign node3004 = (inp[2]) ? 11'b00000100010 : 11'b00001100010;
									assign node3007 = (inp[4]) ? node3021 : node3008;
										assign node3008 = (inp[5]) ? node3016 : node3009;
											assign node3009 = (inp[2]) ? node3013 : node3010;
												assign node3010 = (inp[3]) ? 11'b00011100010 : 11'b00111100000;
												assign node3013 = (inp[3]) ? 11'b00010000000 : 11'b00110000010;
											assign node3016 = (inp[2]) ? node3018 : 11'b00000100000;
												assign node3018 = (inp[3]) ? 11'b00000000000 : 11'b00000000010;
										assign node3021 = (inp[3]) ? node3027 : node3022;
											assign node3022 = (inp[2]) ? 11'b00000000010 : node3023;
												assign node3023 = (inp[5]) ? 11'b00000000010 : 11'b00001000010;
											assign node3027 = (inp[5]) ? 11'b00000000000 : node3028;
												assign node3028 = (inp[2]) ? 11'b00000000000 : 11'b00001000000;
		assign node3032 = (inp[7]) ? node4548 : node3033;
			assign node3033 = (inp[6]) ? node3781 : node3034;
				assign node3034 = (inp[8]) ? node3410 : node3035;
					assign node3035 = (inp[0]) ? node3233 : node3036;
						assign node3036 = (inp[9]) ? node3138 : node3037;
							assign node3037 = (inp[4]) ? node3089 : node3038;
								assign node3038 = (inp[2]) ? node3066 : node3039;
									assign node3039 = (inp[11]) ? node3051 : node3040;
										assign node3040 = (inp[5]) ? node3044 : node3041;
											assign node3041 = (inp[10]) ? 11'b10001101011 : 11'b00001101011;
											assign node3044 = (inp[3]) ? node3048 : node3045;
												assign node3045 = (inp[10]) ? 11'b10101111001 : 11'b00000011001;
												assign node3048 = (inp[10]) ? 11'b00101111111 : 11'b10001111011;
										assign node3051 = (inp[10]) ? node3059 : node3052;
											assign node3052 = (inp[3]) ? node3056 : node3053;
												assign node3053 = (inp[5]) ? 11'b00000111001 : 11'b00001001011;
												assign node3056 = (inp[5]) ? 11'b10101001011 : 11'b10001011001;
											assign node3059 = (inp[3]) ? node3063 : node3060;
												assign node3060 = (inp[5]) ? 11'b10101011001 : 11'b10001001011;
												assign node3063 = (inp[5]) ? 11'b00011001111 : 11'b00001011101;
									assign node3066 = (inp[11]) ? node3078 : node3067;
										assign node3067 = (inp[5]) ? node3073 : node3068;
											assign node3068 = (inp[3]) ? 11'b10101001000 : node3069;
												assign node3069 = (inp[10]) ? 11'b10111001010 : 11'b00101001010;
											assign node3073 = (inp[3]) ? 11'b00000011111 : node3074;
												assign node3074 = (inp[10]) ? 11'b10010011001 : 11'b00101011001;
										assign node3078 = (inp[5]) ? node3086 : node3079;
											assign node3079 = (inp[3]) ? node3083 : node3080;
												assign node3080 = (inp[10]) ? 11'b10111101011 : 11'b00100101011;
												assign node3083 = (inp[10]) ? 11'b00101111111 : 11'b10110111001;
											assign node3086 = (inp[10]) ? 11'b10001111011 : 11'b10011101011;
								assign node3089 = (inp[5]) ? node3113 : node3090;
									assign node3090 = (inp[2]) ? node3102 : node3091;
										assign node3091 = (inp[11]) ? node3097 : node3092;
											assign node3092 = (inp[10]) ? 11'b00101101001 : node3093;
												assign node3093 = (inp[3]) ? 11'b10001101101 : 11'b00001101111;
											assign node3097 = (inp[10]) ? 11'b10111011111 : node3098;
												assign node3098 = (inp[3]) ? 11'b10111001101 : 11'b00011001111;
										assign node3102 = (inp[10]) ? node3110 : node3103;
											assign node3103 = (inp[3]) ? node3107 : node3104;
												assign node3104 = (inp[11]) ? 11'b00110101101 : 11'b00100001100;
												assign node3107 = (inp[11]) ? 11'b10000101101 : 11'b10101101111;
											assign node3110 = (inp[11]) ? 11'b10000111111 : 11'b10111111101;
									assign node3113 = (inp[10]) ? node3127 : node3114;
										assign node3114 = (inp[3]) ? node3120 : node3115;
											assign node3115 = (inp[2]) ? 11'b00111011111 : node3116;
												assign node3116 = (inp[11]) ? 11'b00000011111 : 11'b00010111101;
											assign node3120 = (inp[2]) ? node3124 : node3121;
												assign node3121 = (inp[11]) ? 11'b10100011101 : 11'b10111111111;
												assign node3124 = (inp[11]) ? 11'b10011111111 : 11'b10001011101;
										assign node3127 = (inp[3]) ? node3133 : node3128;
											assign node3128 = (inp[11]) ? node3130 : 11'b10100001111;
												assign node3130 = (inp[2]) ? 11'b10111101101 : 11'b10001001111;
											assign node3133 = (inp[11]) ? 11'b00101001001 : node3134;
												assign node3134 = (inp[2]) ? 11'b00110011001 : 11'b00011111011;
							assign node3138 = (inp[4]) ? node3192 : node3139;
								assign node3139 = (inp[10]) ? node3167 : node3140;
									assign node3140 = (inp[3]) ? node3154 : node3141;
										assign node3141 = (inp[11]) ? node3147 : node3142;
											assign node3142 = (inp[2]) ? 11'b00100011001 : node3143;
												assign node3143 = (inp[5]) ? 11'b00001111001 : 11'b00000101011;
											assign node3147 = (inp[2]) ? node3151 : node3148;
												assign node3148 = (inp[5]) ? 11'b00111001001 : 11'b00100011011;
												assign node3151 = (inp[5]) ? 11'b00010101011 : 11'b00011111001;
										assign node3154 = (inp[5]) ? node3162 : node3155;
											assign node3155 = (inp[2]) ? node3159 : node3156;
												assign node3156 = (inp[11]) ? 11'b10100001101 : 11'b10000101101;
												assign node3159 = (inp[11]) ? 11'b10011101111 : 11'b10100001110;
											assign node3162 = (inp[11]) ? 11'b10100111101 : node3163;
												assign node3163 = (inp[2]) ? 11'b10111011111 : 11'b10000111111;
									assign node3167 = (inp[5]) ? node3179 : node3168;
										assign node3168 = (inp[3]) ? node3174 : node3169;
											assign node3169 = (inp[11]) ? node3171 : 11'b10110011100;
												assign node3171 = (inp[2]) ? 11'b10001111101 : 11'b10100011111;
											assign node3174 = (inp[2]) ? 11'b00110011110 : node3175;
												assign node3175 = (inp[11]) ? 11'b00010011101 : 11'b00000111101;
										assign node3179 = (inp[3]) ? node3185 : node3180;
											assign node3180 = (inp[2]) ? 11'b10010101111 : node3181;
												assign node3181 = (inp[11]) ? 11'b10110001101 : 11'b10100101101;
											assign node3185 = (inp[2]) ? node3189 : node3186;
												assign node3186 = (inp[11]) ? 11'b00000001101 : 11'b00010101111;
												assign node3189 = (inp[11]) ? 11'b00110101101 : 11'b00101001101;
								assign node3192 = (inp[10]) ? node3214 : node3193;
									assign node3193 = (inp[3]) ? node3205 : node3194;
										assign node3194 = (inp[11]) ? node3200 : node3195;
											assign node3195 = (inp[5]) ? 11'b00000011101 : node3196;
												assign node3196 = (inp[2]) ? 11'b00001101111 : 11'b00100101111;
											assign node3200 = (inp[2]) ? 11'b00111101101 : node3201;
												assign node3201 = (inp[5]) ? 11'b00011001111 : 11'b00010011111;
										assign node3205 = (inp[5]) ? node3207 : 11'b10011111001;
											assign node3207 = (inp[11]) ? node3211 : node3208;
												assign node3208 = (inp[2]) ? 11'b10100001011 : 11'b10000101011;
												assign node3211 = (inp[2]) ? 11'b10001101001 : 11'b10111001001;
									assign node3214 = (inp[3]) ? node3224 : node3215;
										assign node3215 = (inp[2]) ? node3219 : node3216;
											assign node3216 = (inp[5]) ? 11'b10010001011 : 11'b10110011011;
											assign node3219 = (inp[5]) ? node3221 : 11'b10010101011;
												assign node3221 = (inp[11]) ? 11'b10100101011 : 11'b10110011001;
										assign node3224 = (inp[11]) ? node3228 : node3225;
											assign node3225 = (inp[2]) ? 11'b00001101011 : 11'b00100101011;
											assign node3228 = (inp[2]) ? 11'b00010101001 : node3229;
												assign node3229 = (inp[5]) ? 11'b00110001001 : 11'b00110011001;
						assign node3233 = (inp[3]) ? node3327 : node3234;
							assign node3234 = (inp[5]) ? node3280 : node3235;
								assign node3235 = (inp[2]) ? node3255 : node3236;
									assign node3236 = (inp[11]) ? node3244 : node3237;
										assign node3237 = (inp[9]) ? node3241 : node3238;
											assign node3238 = (inp[10]) ? 11'b00001101111 : 11'b00001101011;
											assign node3241 = (inp[10]) ? 11'b00000111011 : 11'b00000101111;
										assign node3244 = (inp[4]) ? node3250 : node3245;
											assign node3245 = (inp[10]) ? 11'b00010001011 : node3246;
												assign node3246 = (inp[9]) ? 11'b00100011111 : 11'b00001011011;
											assign node3250 = (inp[9]) ? node3252 : 11'b00111001111;
												assign node3252 = (inp[10]) ? 11'b00110001011 : 11'b00010001111;
									assign node3255 = (inp[11]) ? node3269 : node3256;
										assign node3256 = (inp[4]) ? node3264 : node3257;
											assign node3257 = (inp[10]) ? node3261 : node3258;
												assign node3258 = (inp[9]) ? 11'b00000001110 : 11'b00001001010;
												assign node3261 = (inp[9]) ? 11'b00010011010 : 11'b00011001110;
											assign node3264 = (inp[10]) ? node3266 : 11'b00000001000;
												assign node3266 = (inp[9]) ? 11'b00110111001 : 11'b00011111101;
										assign node3269 = (inp[10]) ? node3277 : node3270;
											assign node3270 = (inp[9]) ? node3274 : node3271;
												assign node3271 = (inp[4]) ? 11'b00010111001 : 11'b00010111011;
												assign node3274 = (inp[4]) ? 11'b00001001111 : 11'b00111111111;
											assign node3277 = (inp[9]) ? 11'b00001101001 : 11'b00100101101;
								assign node3280 = (inp[11]) ? node3306 : node3281;
									assign node3281 = (inp[2]) ? node3291 : node3282;
										assign node3282 = (inp[9]) ? node3284 : 11'b00011111111;
											assign node3284 = (inp[10]) ? node3288 : node3285;
												assign node3285 = (inp[4]) ? 11'b00110111111 : 11'b00000101111;
												assign node3288 = (inp[4]) ? 11'b00100111001 : 11'b00100111011;
										assign node3291 = (inp[9]) ? node3299 : node3292;
											assign node3292 = (inp[10]) ? node3296 : node3293;
												assign node3293 = (inp[4]) ? 11'b00111001001 : 11'b00000001011;
												assign node3296 = (inp[4]) ? 11'b00010011111 : 11'b00110001111;
											assign node3299 = (inp[10]) ? node3303 : node3300;
												assign node3300 = (inp[4]) ? 11'b00100011111 : 11'b00010001101;
												assign node3303 = (inp[4]) ? 11'b00111111011 : 11'b00101011001;
									assign node3306 = (inp[4]) ? node3318 : node3307;
										assign node3307 = (inp[9]) ? node3313 : node3308;
											assign node3308 = (inp[10]) ? 11'b00011011101 : node3309;
												assign node3309 = (inp[2]) ? 11'b00011111001 : 11'b00000111001;
											assign node3313 = (inp[10]) ? node3315 : 11'b00110111101;
												assign node3315 = (inp[2]) ? 11'b00110101011 : 11'b00110001001;
										assign node3318 = (inp[9]) ? node3322 : node3319;
											assign node3319 = (inp[2]) ? 11'b00101101101 : 11'b00101001101;
											assign node3322 = (inp[10]) ? 11'b00110101001 : node3323;
												assign node3323 = (inp[2]) ? 11'b00111101101 : 11'b00111001101;
							assign node3327 = (inp[9]) ? node3373 : node3328;
								assign node3328 = (inp[2]) ? node3350 : node3329;
									assign node3329 = (inp[11]) ? node3341 : node3330;
										assign node3330 = (inp[5]) ? node3338 : node3331;
											assign node3331 = (inp[10]) ? node3335 : node3332;
												assign node3332 = (inp[4]) ? 11'b00001111001 : 11'b00001101001;
												assign node3335 = (inp[4]) ? 11'b00101101001 : 11'b00001101001;
											assign node3338 = (inp[4]) ? 11'b00111101001 : 11'b00101101001;
										assign node3341 = (inp[5]) ? node3347 : node3342;
											assign node3342 = (inp[4]) ? 11'b00011001001 : node3343;
												assign node3343 = (inp[10]) ? 11'b00101001001 : 11'b00001001001;
											assign node3347 = (inp[4]) ? 11'b00001011011 : 11'b00111001011;
									assign node3350 = (inp[4]) ? node3360 : node3351;
										assign node3351 = (inp[11]) ? node3357 : node3352;
											assign node3352 = (inp[5]) ? node3354 : 11'b00001001000;
												assign node3354 = (inp[10]) ? 11'b00000001011 : 11'b00110001001;
											assign node3357 = (inp[10]) ? 11'b00110101011 : 11'b00010101001;
										assign node3360 = (inp[10]) ? node3368 : node3361;
											assign node3361 = (inp[5]) ? node3365 : node3362;
												assign node3362 = (inp[11]) ? 11'b00100111011 : 11'b00011111011;
												assign node3365 = (inp[11]) ? 11'b00011111001 : 11'b00101011001;
											assign node3368 = (inp[11]) ? node3370 : 11'b00101101011;
												assign node3370 = (inp[5]) ? 11'b00011101011 : 11'b00011001011;
								assign node3373 = (inp[10]) ? node3395 : node3374;
									assign node3374 = (inp[4]) ? node3386 : node3375;
										assign node3375 = (inp[2]) ? node3381 : node3376;
											assign node3376 = (inp[11]) ? 11'b00010011011 : node3377;
												assign node3377 = (inp[5]) ? 11'b00100111001 : 11'b00000111001;
											assign node3381 = (inp[11]) ? 11'b00111111001 : node3382;
												assign node3382 = (inp[5]) ? 11'b00111011011 : 11'b00010011000;
										assign node3386 = (inp[5]) ? node3392 : node3387;
											assign node3387 = (inp[11]) ? 11'b00110001001 : node3388;
												assign node3388 = (inp[2]) ? 11'b00110101011 : 11'b00100101001;
											assign node3392 = (inp[2]) ? 11'b00000101011 : 11'b00010001011;
									assign node3395 = (inp[4]) ? node3403 : node3396;
										assign node3396 = (inp[5]) ? node3400 : node3397;
											assign node3397 = (inp[11]) ? 11'b00010101011 : 11'b00000001010;
											assign node3400 = (inp[11]) ? 11'b00000101001 : 11'b00010101001;
										assign node3403 = (inp[5]) ? 11'b00001101011 : node3404;
											assign node3404 = (inp[11]) ? node3406 : 11'b00000101001;
												assign node3406 = (inp[2]) ? 11'b00001001001 : 11'b00000001001;
					assign node3410 = (inp[0]) ? node3588 : node3411;
						assign node3411 = (inp[11]) ? node3499 : node3412;
							assign node3412 = (inp[5]) ? node3460 : node3413;
								assign node3413 = (inp[2]) ? node3437 : node3414;
									assign node3414 = (inp[9]) ? node3428 : node3415;
										assign node3415 = (inp[10]) ? node3421 : node3416;
											assign node3416 = (inp[4]) ? 11'b10000101110 : node3417;
												assign node3417 = (inp[3]) ? 11'b10100001001 : 11'b00000001011;
											assign node3421 = (inp[3]) ? node3425 : node3422;
												assign node3422 = (inp[4]) ? 11'b10100111100 : 11'b10001101010;
												assign node3425 = (inp[4]) ? 11'b00011101010 : 11'b00101101100;
										assign node3428 = (inp[10]) ? node3434 : node3429;
											assign node3429 = (inp[3]) ? node3431 : 11'b00011101010;
												assign node3431 = (inp[4]) ? 11'b10011111010 : 11'b10111101100;
											assign node3434 = (inp[3]) ? 11'b00100111010 : 11'b10010111110;
									assign node3437 = (inp[9]) ? node3451 : node3438;
										assign node3438 = (inp[10]) ? node3444 : node3439;
											assign node3439 = (inp[3]) ? node3441 : 11'b00100101011;
												assign node3441 = (inp[4]) ? 11'b10110001101 : 11'b10010101001;
											assign node3444 = (inp[3]) ? node3448 : node3445;
												assign node3445 = (inp[4]) ? 11'b10000011111 : 11'b10111001011;
												assign node3448 = (inp[4]) ? 11'b00100001001 : 11'b00001001111;
										assign node3451 = (inp[3]) ? node3455 : node3452;
											assign node3452 = (inp[10]) ? 11'b10111001001 : 11'b00011001111;
											assign node3455 = (inp[4]) ? node3457 : 11'b10001001111;
												assign node3457 = (inp[10]) ? 11'b00001011011 : 11'b10101011011;
								assign node3460 = (inp[9]) ? node3484 : node3461;
									assign node3461 = (inp[3]) ? node3475 : node3462;
										assign node3462 = (inp[4]) ? node3468 : node3463;
											assign node3463 = (inp[2]) ? 11'b10001111000 : node3464;
												assign node3464 = (inp[10]) ? 11'b10100011000 : 11'b00001011000;
											assign node3468 = (inp[10]) ? node3472 : node3469;
												assign node3469 = (inp[2]) ? 11'b00010111110 : 11'b00111111100;
												assign node3472 = (inp[2]) ? 11'b10110101100 : 11'b10000101110;
										assign node3475 = (inp[10]) ? node3479 : node3476;
											assign node3476 = (inp[4]) ? 11'b10010111110 : 11'b10111111010;
											assign node3479 = (inp[4]) ? 11'b00101011010 : node3480;
												assign node3480 = (inp[2]) ? 11'b00011111110 : 11'b00110011110;
									assign node3484 = (inp[4]) ? node3492 : node3485;
										assign node3485 = (inp[10]) ? node3489 : node3486;
											assign node3486 = (inp[3]) ? 11'b10001111110 : 11'b00010011000;
											assign node3489 = (inp[3]) ? 11'b00000101100 : 11'b10110101110;
										assign node3492 = (inp[3]) ? node3494 : 11'b10111111010;
											assign node3494 = (inp[2]) ? 11'b10001001000 : node3495;
												assign node3495 = (inp[10]) ? 11'b00101101000 : 11'b10110101000;
							assign node3499 = (inp[5]) ? node3545 : node3500;
								assign node3500 = (inp[2]) ? node3522 : node3501;
									assign node3501 = (inp[9]) ? node3511 : node3502;
										assign node3502 = (inp[4]) ? node3506 : node3503;
											assign node3503 = (inp[10]) ? 11'b10110101000 : 11'b00000101000;
											assign node3506 = (inp[10]) ? 11'b00100011000 : node3507;
												assign node3507 = (inp[3]) ? 11'b10010001100 : 11'b00110001110;
										assign node3511 = (inp[4]) ? node3517 : node3512;
											assign node3512 = (inp[3]) ? node3514 : 11'b00111011000;
												assign node3514 = (inp[10]) ? 11'b00101011100 : 11'b10101001100;
											assign node3517 = (inp[3]) ? node3519 : 11'b00001011110;
												assign node3519 = (inp[10]) ? 11'b00111011000 : 11'b10011011000;
									assign node3522 = (inp[4]) ? node3532 : node3523;
										assign node3523 = (inp[10]) ? node3529 : node3524;
											assign node3524 = (inp[3]) ? node3526 : 11'b00000011011;
												assign node3526 = (inp[9]) ? 11'b10010001101 : 11'b10010011011;
											assign node3529 = (inp[9]) ? 11'b00001111110 : 11'b10000001011;
										assign node3532 = (inp[9]) ? node3538 : node3533;
											assign node3533 = (inp[10]) ? 11'b00001111000 : node3534;
												assign node3534 = (inp[3]) ? 11'b10101101110 : 11'b00011101100;
											assign node3538 = (inp[3]) ? node3542 : node3539;
												assign node3539 = (inp[10]) ? 11'b10000111010 : 11'b00100111110;
												assign node3542 = (inp[10]) ? 11'b00010111000 : 11'b10110111000;
								assign node3545 = (inp[3]) ? node3567 : node3546;
									assign node3546 = (inp[10]) ? node3558 : node3547;
										assign node3547 = (inp[9]) ? node3551 : node3548;
											assign node3548 = (inp[4]) ? 11'b00001011110 : 11'b00100011010;
											assign node3551 = (inp[4]) ? node3555 : node3552;
												assign node3552 = (inp[2]) ? 11'b00100001000 : 11'b00000101000;
												assign node3555 = (inp[2]) ? 11'b00000001100 : 11'b00100001110;
										assign node3558 = (inp[9]) ? node3564 : node3559;
											assign node3559 = (inp[4]) ? node3561 : 11'b10100011000;
												assign node3561 = (inp[2]) ? 11'b10001001100 : 11'b10111001100;
											assign node3564 = (inp[4]) ? 11'b10000001010 : 11'b10001001110;
									assign node3567 = (inp[10]) ? node3577 : node3568;
										assign node3568 = (inp[2]) ? node3572 : node3569;
											assign node3569 = (inp[4]) ? 11'b10100001000 : 11'b10100111110;
											assign node3572 = (inp[9]) ? node3574 : 11'b10011011100;
												assign node3574 = (inp[4]) ? 11'b10010001010 : 11'b10011011110;
										assign node3577 = (inp[9]) ? node3585 : node3578;
											assign node3578 = (inp[4]) ? node3582 : node3579;
												assign node3579 = (inp[2]) ? 11'b00110001110 : 11'b00000101110;
												assign node3582 = (inp[2]) ? 11'b00010001010 : 11'b00110001010;
											assign node3585 = (inp[2]) ? 11'b00011001100 : 11'b00111001110;
						assign node3588 = (inp[3]) ? node3690 : node3589;
							assign node3589 = (inp[4]) ? node3637 : node3590;
								assign node3590 = (inp[5]) ? node3616 : node3591;
									assign node3591 = (inp[11]) ? node3605 : node3592;
										assign node3592 = (inp[9]) ? node3600 : node3593;
											assign node3593 = (inp[10]) ? node3597 : node3594;
												assign node3594 = (inp[2]) ? 11'b00100101011 : 11'b00100001011;
												assign node3597 = (inp[2]) ? 11'b00101001111 : 11'b00101101110;
											assign node3600 = (inp[2]) ? 11'b00111011001 : node3601;
												assign node3601 = (inp[10]) ? 11'b00110111010 : 11'b00111101110;
										assign node3605 = (inp[9]) ? node3611 : node3606;
											assign node3606 = (inp[2]) ? node3608 : 11'b00110111100;
												assign node3608 = (inp[10]) ? 11'b00100011101 : 11'b00111011001;
											assign node3611 = (inp[10]) ? node3613 : 11'b00001011100;
												assign node3613 = (inp[2]) ? 11'b00101101010 : 11'b00101001000;
									assign node3616 = (inp[11]) ? node3628 : node3617;
										assign node3617 = (inp[2]) ? node3623 : node3618;
											assign node3618 = (inp[9]) ? 11'b00001111000 : node3619;
												assign node3619 = (inp[10]) ? 11'b00010001110 : 11'b00100001010;
											assign node3623 = (inp[10]) ? 11'b00001101100 : node3624;
												assign node3624 = (inp[9]) ? 11'b00101101100 : 11'b00101101010;
										assign node3628 = (inp[2]) ? node3634 : node3629;
											assign node3629 = (inp[10]) ? 11'b00011001010 : node3630;
												assign node3630 = (inp[9]) ? 11'b00000111110 : 11'b00101111010;
											assign node3634 = (inp[10]) ? 11'b00110011110 : 11'b00110011010;
								assign node3637 = (inp[11]) ? node3663 : node3638;
									assign node3638 = (inp[9]) ? node3650 : node3639;
										assign node3639 = (inp[10]) ? node3647 : node3640;
											assign node3640 = (inp[5]) ? node3644 : node3641;
												assign node3641 = (inp[2]) ? 11'b00100001001 : 11'b00100101010;
												assign node3644 = (inp[2]) ? 11'b00000101010 : 11'b00011101000;
											assign node3647 = (inp[5]) ? 11'b00100111100 : 11'b00101111110;
										assign node3650 = (inp[2]) ? node3656 : node3651;
											assign node3651 = (inp[10]) ? 11'b00001111000 : node3652;
												assign node3652 = (inp[5]) ? 11'b00010111100 : 11'b00011111110;
											assign node3656 = (inp[5]) ? node3660 : node3657;
												assign node3657 = (inp[10]) ? 11'b00011011011 : 11'b00001011111;
												assign node3660 = (inp[10]) ? 11'b00011011000 : 11'b00011011100;
									assign node3663 = (inp[5]) ? node3679 : node3664;
										assign node3664 = (inp[2]) ? node3672 : node3665;
											assign node3665 = (inp[9]) ? node3669 : node3666;
												assign node3666 = (inp[10]) ? 11'b00000001110 : 11'b00110011000;
												assign node3669 = (inp[10]) ? 11'b00011001010 : 11'b00101001110;
											assign node3672 = (inp[9]) ? node3676 : node3673;
												assign node3673 = (inp[10]) ? 11'b00011101100 : 11'b00111111010;
												assign node3676 = (inp[10]) ? 11'b00010101010 : 11'b00110101100;
										assign node3679 = (inp[9]) ? node3685 : node3680;
											assign node3680 = (inp[10]) ? node3682 : 11'b00011011010;
												assign node3682 = (inp[2]) ? 11'b00010001110 : 11'b00011001100;
											assign node3685 = (inp[10]) ? 11'b00010001000 : node3686;
												assign node3686 = (inp[2]) ? 11'b00010001100 : 11'b00000001100;
							assign node3690 = (inp[10]) ? node3736 : node3691;
								assign node3691 = (inp[2]) ? node3711 : node3692;
									assign node3692 = (inp[11]) ? node3698 : node3693;
										assign node3693 = (inp[9]) ? 11'b00111101000 : node3694;
											assign node3694 = (inp[5]) ? 11'b00110111010 : 11'b00000111000;
										assign node3698 = (inp[4]) ? node3704 : node3699;
											assign node3699 = (inp[9]) ? 11'b00101011010 : node3700;
												assign node3700 = (inp[5]) ? 11'b00111101000 : 11'b00010101010;
											assign node3704 = (inp[5]) ? node3708 : node3705;
												assign node3705 = (inp[9]) ? 11'b00111001000 : 11'b00110011010;
												assign node3708 = (inp[9]) ? 11'b00010001010 : 11'b00011011010;
									assign node3711 = (inp[5]) ? node3721 : node3712;
										assign node3712 = (inp[11]) ? 11'b00100101000 : node3713;
											assign node3713 = (inp[9]) ? node3717 : node3714;
												assign node3714 = (inp[4]) ? 11'b00010011011 : 11'b00010101001;
												assign node3717 = (inp[4]) ? 11'b00101001001 : 11'b00001011011;
										assign node3721 = (inp[9]) ? node3729 : node3722;
											assign node3722 = (inp[4]) ? node3726 : node3723;
												assign node3723 = (inp[11]) ? 11'b00100001000 : 11'b00111101000;
												assign node3726 = (inp[11]) ? 11'b00001011000 : 11'b00100111000;
											assign node3729 = (inp[4]) ? node3733 : node3730;
												assign node3730 = (inp[11]) ? 11'b00001011010 : 11'b00110111010;
												assign node3733 = (inp[11]) ? 11'b00000001010 : 11'b00001001010;
								assign node3736 = (inp[9]) ? node3758 : node3737;
									assign node3737 = (inp[2]) ? node3751 : node3738;
										assign node3738 = (inp[5]) ? node3746 : node3739;
											assign node3739 = (inp[11]) ? node3743 : node3740;
												assign node3740 = (inp[4]) ? 11'b00111101000 : 11'b00011101000;
												assign node3743 = (inp[4]) ? 11'b00000001000 : 11'b00111001010;
											assign node3746 = (inp[4]) ? 11'b00100101010 : node3747;
												assign node3747 = (inp[11]) ? 11'b00100101000 : 11'b00010001000;
										assign node3751 = (inp[5]) ? 11'b00101001010 : node3752;
											assign node3752 = (inp[11]) ? 11'b00110001011 : node3753;
												assign node3753 = (inp[4]) ? 11'b00110001001 : 11'b00011001001;
									assign node3758 = (inp[11]) ? node3770 : node3759;
										assign node3759 = (inp[5]) ? node3763 : node3760;
											assign node3760 = (inp[2]) ? 11'b00000001011 : 11'b00000101010;
											assign node3763 = (inp[4]) ? node3767 : node3764;
												assign node3764 = (inp[2]) ? 11'b00010101000 : 11'b00011101010;
												assign node3767 = (inp[2]) ? 11'b00001001000 : 11'b00001101000;
										assign node3770 = (inp[4]) ? node3774 : node3771;
											assign node3771 = (inp[2]) ? 11'b00001001000 : 11'b00001001010;
											assign node3774 = (inp[2]) ? node3778 : node3775;
												assign node3775 = (inp[5]) ? 11'b00000001000 : 11'b00001001000;
												assign node3778 = (inp[5]) ? 11'b00000001000 : 11'b00000101000;
				assign node3781 = (inp[2]) ? node4169 : node3782;
					assign node3782 = (inp[8]) ? node3988 : node3783;
						assign node3783 = (inp[5]) ? node3881 : node3784;
							assign node3784 = (inp[11]) ? node3830 : node3785;
								assign node3785 = (inp[4]) ? node3809 : node3786;
									assign node3786 = (inp[9]) ? node3800 : node3787;
										assign node3787 = (inp[10]) ? node3795 : node3788;
											assign node3788 = (inp[3]) ? node3792 : node3789;
												assign node3789 = (inp[0]) ? 11'b00011101010 : 11'b00001101010;
												assign node3792 = (inp[0]) ? 11'b00001101000 : 11'b10011101000;
											assign node3795 = (inp[0]) ? 11'b00011101110 : node3796;
												assign node3796 = (inp[3]) ? 11'b00011101110 : 11'b10001101000;
										assign node3800 = (inp[0]) ? node3806 : node3801;
											assign node3801 = (inp[10]) ? 11'b10000111110 : node3802;
												assign node3802 = (inp[3]) ? 11'b10010101110 : 11'b00001101000;
											assign node3806 = (inp[3]) ? 11'b00000101000 : 11'b00010111000;
									assign node3809 = (inp[3]) ? node3819 : node3810;
										assign node3810 = (inp[0]) ? node3816 : node3811;
											assign node3811 = (inp[9]) ? node3813 : 11'b00000101110;
												assign node3813 = (inp[10]) ? 11'b10101101010 : 11'b00101101100;
											assign node3816 = (inp[10]) ? 11'b00011111110 : 11'b00111111100;
										assign node3819 = (inp[0]) ? node3823 : node3820;
											assign node3820 = (inp[9]) ? 11'b10111111010 : 11'b00111101010;
											assign node3823 = (inp[9]) ? node3827 : node3824;
												assign node3824 = (inp[10]) ? 11'b00101101010 : 11'b00000111000;
												assign node3827 = (inp[10]) ? 11'b00001101000 : 11'b00101101010;
								assign node3830 = (inp[0]) ? node3856 : node3831;
									assign node3831 = (inp[4]) ? node3845 : node3832;
										assign node3832 = (inp[9]) ? node3838 : node3833;
											assign node3833 = (inp[3]) ? 11'b10000111010 : node3834;
												assign node3834 = (inp[10]) ? 11'b10010101000 : 11'b00010101010;
											assign node3838 = (inp[10]) ? node3842 : node3839;
												assign node3839 = (inp[3]) ? 11'b10100101100 : 11'b00110111000;
												assign node3842 = (inp[3]) ? 11'b00001011100 : 11'b10111011110;
										assign node3845 = (inp[9]) ? node3853 : node3846;
											assign node3846 = (inp[3]) ? node3850 : node3847;
												assign node3847 = (inp[10]) ? 11'b10111011100 : 11'b00011001110;
												assign node3850 = (inp[10]) ? 11'b00100011010 : 11'b10101001110;
											assign node3853 = (inp[3]) ? 11'b10010011000 : 11'b10100011010;
									assign node3856 = (inp[4]) ? node3870 : node3857;
										assign node3857 = (inp[9]) ? node3865 : node3858;
											assign node3858 = (inp[3]) ? node3862 : node3859;
												assign node3859 = (inp[10]) ? 11'b00010111110 : 11'b00010111010;
												assign node3862 = (inp[10]) ? 11'b00100101010 : 11'b00000101000;
											assign node3865 = (inp[10]) ? node3867 : 11'b00101011010;
												assign node3867 = (inp[3]) ? 11'b00011001000 : 11'b00001001010;
										assign node3870 = (inp[9]) ? node3874 : node3871;
											assign node3871 = (inp[3]) ? 11'b00111011000 : 11'b00101001100;
											assign node3874 = (inp[10]) ? node3878 : node3875;
												assign node3875 = (inp[3]) ? 11'b00110001010 : 11'b00000001100;
												assign node3878 = (inp[3]) ? 11'b00000001000 : 11'b00100001010;
							assign node3881 = (inp[11]) ? node3937 : node3882;
								assign node3882 = (inp[4]) ? node3912 : node3883;
									assign node3883 = (inp[0]) ? node3897 : node3884;
										assign node3884 = (inp[3]) ? node3890 : node3885;
											assign node3885 = (inp[9]) ? 11'b00011011010 : node3886;
												assign node3886 = (inp[10]) ? 11'b10101011000 : 11'b00000011000;
											assign node3890 = (inp[10]) ? node3894 : node3891;
												assign node3891 = (inp[9]) ? 11'b10001011100 : 11'b10011011010;
												assign node3894 = (inp[9]) ? 11'b00000001110 : 11'b00111011110;
										assign node3897 = (inp[3]) ? node3905 : node3898;
											assign node3898 = (inp[10]) ? node3902 : node3899;
												assign node3899 = (inp[9]) ? 11'b00011001100 : 11'b00011001010;
												assign node3902 = (inp[9]) ? 11'b00110011010 : 11'b00111001100;
											assign node3905 = (inp[10]) ? node3909 : node3906;
												assign node3906 = (inp[9]) ? 11'b00101011000 : 11'b00101001010;
												assign node3909 = (inp[9]) ? 11'b00010001000 : 11'b00001001010;
									assign node3912 = (inp[9]) ? node3926 : node3913;
										assign node3913 = (inp[0]) ? node3921 : node3914;
											assign node3914 = (inp[3]) ? node3918 : node3915;
												assign node3915 = (inp[10]) ? 11'b10000001110 : 11'b00010011100;
												assign node3918 = (inp[10]) ? 11'b00010011000 : 11'b10100011110;
											assign node3921 = (inp[3]) ? 11'b00111100011 : node3922;
												assign node3922 = (inp[10]) ? 11'b00000011100 : 11'b00100001000;
										assign node3926 = (inp[3]) ? node3930 : node3927;
											assign node3927 = (inp[10]) ? 11'b00111110011 : 11'b00101110111;
											assign node3930 = (inp[10]) ? node3934 : node3931;
												assign node3931 = (inp[0]) ? 11'b00001100001 : 11'b10011100001;
												assign node3934 = (inp[0]) ? 11'b00001100011 : 11'b00111100011;
								assign node3937 = (inp[9]) ? node3965 : node3938;
									assign node3938 = (inp[10]) ? node3954 : node3939;
										assign node3939 = (inp[3]) ? node3947 : node3940;
											assign node3940 = (inp[0]) ? node3944 : node3941;
												assign node3941 = (inp[4]) ? 11'b00001110111 : 11'b00011110001;
												assign node3944 = (inp[4]) ? 11'b00111110001 : 11'b00011110001;
											assign node3947 = (inp[0]) ? node3951 : node3948;
												assign node3948 = (inp[4]) ? 11'b10111110101 : 11'b10101100001;
												assign node3951 = (inp[4]) ? 11'b00001110001 : 11'b00100100011;
										assign node3954 = (inp[3]) ? node3962 : node3955;
											assign node3955 = (inp[4]) ? node3959 : node3956;
												assign node3956 = (inp[0]) ? 11'b00000110111 : 11'b10110110011;
												assign node3959 = (inp[0]) ? 11'b00111100111 : 11'b10011100111;
											assign node3962 = (inp[4]) ? 11'b00011100001 : 11'b00110100001;
									assign node3965 = (inp[3]) ? node3979 : node3966;
										assign node3966 = (inp[10]) ? node3974 : node3967;
											assign node3967 = (inp[4]) ? node3971 : node3968;
												assign node3968 = (inp[0]) ? 11'b00100110111 : 11'b00110100011;
												assign node3971 = (inp[0]) ? 11'b00101100101 : 11'b00011100101;
											assign node3974 = (inp[4]) ? 11'b10000100011 : node3975;
												assign node3975 = (inp[0]) ? 11'b00100100001 : 11'b10100100101;
										assign node3979 = (inp[0]) ? node3983 : node3980;
											assign node3980 = (inp[10]) ? 11'b00110100001 : 11'b10100100011;
											assign node3983 = (inp[10]) ? 11'b00001100011 : node3984;
												assign node3984 = (inp[4]) ? 11'b00010100011 : 11'b00010110001;
						assign node3988 = (inp[0]) ? node4078 : node3989;
							assign node3989 = (inp[11]) ? node4037 : node3990;
								assign node3990 = (inp[5]) ? node4010 : node3991;
									assign node3991 = (inp[9]) ? node3999 : node3992;
										assign node3992 = (inp[4]) ? node3996 : node3993;
											assign node3993 = (inp[10]) ? 11'b10010100001 : 11'b00000100011;
											assign node3996 = (inp[10]) ? 11'b00000000001 : 11'b00101000101;
										assign node3999 = (inp[10]) ? node4007 : node4000;
											assign node4000 = (inp[4]) ? node4004 : node4001;
												assign node4001 = (inp[3]) ? 11'b10101000101 : 11'b00011000001;
												assign node4004 = (inp[3]) ? 11'b10010010001 : 11'b00110000111;
											assign node4007 = (inp[4]) ? 11'b00111010011 : 11'b00111010101;
									assign node4010 = (inp[9]) ? node4026 : node4011;
										assign node4011 = (inp[4]) ? node4019 : node4012;
											assign node4012 = (inp[10]) ? node4016 : node4013;
												assign node4013 = (inp[3]) ? 11'b10000110011 : 11'b00001110001;
												assign node4016 = (inp[3]) ? 11'b00100110101 : 11'b10110110001;
											assign node4019 = (inp[10]) ? node4023 : node4020;
												assign node4020 = (inp[3]) ? 11'b10011110101 : 11'b00111110101;
												assign node4023 = (inp[3]) ? 11'b00001110011 : 11'b10001100111;
										assign node4026 = (inp[4]) ? node4032 : node4027;
											assign node4027 = (inp[10]) ? node4029 : 11'b10010110101;
												assign node4029 = (inp[3]) ? 11'b00101100111 : 11'b10010100101;
											assign node4032 = (inp[3]) ? node4034 : 11'b10100110011;
												assign node4034 = (inp[10]) ? 11'b00110100001 : 11'b10100100011;
								assign node4037 = (inp[10]) ? node4055 : node4038;
									assign node4038 = (inp[3]) ? node4050 : node4039;
										assign node4039 = (inp[4]) ? node4043 : node4040;
											assign node4040 = (inp[5]) ? 11'b00011000011 : 11'b00101010001;
											assign node4043 = (inp[5]) ? node4047 : node4044;
												assign node4044 = (inp[9]) ? 11'b00011110101 : 11'b00110000111;
												assign node4047 = (inp[9]) ? 11'b00100000101 : 11'b00101010101;
										assign node4050 = (inp[5]) ? 11'b10101010101 : node4051;
											assign node4051 = (inp[9]) ? 11'b10110000111 : 11'b10101010001;
									assign node4055 = (inp[3]) ? node4065 : node4056;
										assign node4056 = (inp[4]) ? 11'b10110000111 : node4057;
											assign node4057 = (inp[9]) ? node4061 : node4058;
												assign node4058 = (inp[5]) ? 11'b10000110001 : 11'b10111000011;
												assign node4061 = (inp[5]) ? 11'b10111000111 : 11'b10010010101;
										assign node4065 = (inp[4]) ? node4073 : node4066;
											assign node4066 = (inp[5]) ? node4070 : node4067;
												assign node4067 = (inp[9]) ? 11'b00100010101 : 11'b00011010101;
												assign node4070 = (inp[9]) ? 11'b00111000111 : 11'b00011000111;
											assign node4073 = (inp[5]) ? 11'b00110000001 : node4074;
												assign node4074 = (inp[9]) ? 11'b00111110001 : 11'b00111110011;
							assign node4078 = (inp[3]) ? node4132 : node4079;
								assign node4079 = (inp[5]) ? node4105 : node4080;
									assign node4080 = (inp[9]) ? node4096 : node4081;
										assign node4081 = (inp[10]) ? node4089 : node4082;
											assign node4082 = (inp[11]) ? node4086 : node4083;
												assign node4083 = (inp[4]) ? 11'b00110000011 : 11'b00110100011;
												assign node4086 = (inp[4]) ? 11'b00100010011 : 11'b00111010001;
											assign node4089 = (inp[4]) ? node4093 : node4090;
												assign node4090 = (inp[11]) ? 11'b00101010111 : 11'b00111000111;
												assign node4093 = (inp[11]) ? 11'b00011100111 : 11'b00110010101;
										assign node4096 = (inp[11]) ? node4102 : node4097;
											assign node4097 = (inp[4]) ? 11'b00000010111 : node4098;
												assign node4098 = (inp[10]) ? 11'b00101010011 : 11'b00101000101;
											assign node4102 = (inp[10]) ? 11'b00110000001 : 11'b00010010111;
									assign node4105 = (inp[11]) ? node4117 : node4106;
										assign node4106 = (inp[4]) ? node4112 : node4107;
											assign node4107 = (inp[10]) ? 11'b00000100101 : node4108;
												assign node4108 = (inp[9]) ? 11'b00100100111 : 11'b00110100011;
											assign node4112 = (inp[9]) ? node4114 : 11'b00111110111;
												assign node4114 = (inp[10]) ? 11'b00010110001 : 11'b00001110101;
										assign node4117 = (inp[10]) ? node4125 : node4118;
											assign node4118 = (inp[9]) ? node4122 : node4119;
												assign node4119 = (inp[4]) ? 11'b00011010001 : 11'b00110110011;
												assign node4122 = (inp[4]) ? 11'b00010000111 : 11'b00011010101;
											assign node4125 = (inp[9]) ? node4129 : node4126;
												assign node4126 = (inp[4]) ? 11'b00000000111 : 11'b00100110101;
												assign node4129 = (inp[4]) ? 11'b00000000001 : 11'b00001000011;
								assign node4132 = (inp[10]) ? node4152 : node4133;
									assign node4133 = (inp[11]) ? node4141 : node4134;
										assign node4134 = (inp[5]) ? node4138 : node4135;
											assign node4135 = (inp[9]) ? 11'b00011010011 : 11'b00000100001;
											assign node4138 = (inp[9]) ? 11'b00100110001 : 11'b00111110011;
										assign node4141 = (inp[5]) ? node4145 : node4142;
											assign node4142 = (inp[9]) ? 11'b00111100011 : 11'b00011000011;
											assign node4145 = (inp[4]) ? node4149 : node4146;
												assign node4146 = (inp[9]) ? 11'b00011010001 : 11'b00110100001;
												assign node4149 = (inp[9]) ? 11'b00010000011 : 11'b00010010011;
									assign node4152 = (inp[4]) ? node4162 : node4153;
										assign node4153 = (inp[9]) ? node4157 : node4154;
											assign node4154 = (inp[11]) ? 11'b00111000001 : 11'b00011000011;
											assign node4157 = (inp[11]) ? node4159 : 11'b00001000001;
												assign node4159 = (inp[5]) ? 11'b00001000011 : 11'b00010000011;
										assign node4162 = (inp[5]) ? node4166 : node4163;
											assign node4163 = (inp[11]) ? 11'b00001100001 : 11'b00001000011;
											assign node4166 = (inp[11]) ? 11'b00000000001 : 11'b00000100001;
					assign node4169 = (inp[5]) ? node4363 : node4170;
						assign node4170 = (inp[11]) ? node4266 : node4171;
							assign node4171 = (inp[8]) ? node4217 : node4172;
								assign node4172 = (inp[0]) ? node4196 : node4173;
									assign node4173 = (inp[4]) ? node4187 : node4174;
										assign node4174 = (inp[10]) ? node4180 : node4175;
											assign node4175 = (inp[3]) ? node4177 : 11'b00101000011;
												assign node4177 = (inp[9]) ? 11'b10101000101 : 11'b10101000011;
											assign node4180 = (inp[9]) ? node4184 : node4181;
												assign node4181 = (inp[3]) ? 11'b00111000111 : 11'b10111000001;
												assign node4184 = (inp[3]) ? 11'b00110010111 : 11'b10110010111;
										assign node4187 = (inp[9]) ? node4191 : node4188;
											assign node4188 = (inp[10]) ? 11'b10110010111 : 11'b00100000101;
											assign node4191 = (inp[3]) ? node4193 : 11'b10001100010;
												assign node4193 = (inp[10]) ? 11'b00011110000 : 11'b10001110010;
									assign node4196 = (inp[10]) ? node4206 : node4197;
										assign node4197 = (inp[9]) ? node4201 : node4198;
											assign node4198 = (inp[4]) ? 11'b00010000001 : 11'b00011000011;
											assign node4201 = (inp[4]) ? 11'b00111110110 : node4202;
												assign node4202 = (inp[3]) ? 11'b00011010001 : 11'b00011000101;
										assign node4206 = (inp[3]) ? node4212 : node4207;
											assign node4207 = (inp[9]) ? 11'b00000010011 : node4208;
												assign node4208 = (inp[4]) ? 11'b00000010111 : 11'b00001000101;
											assign node4212 = (inp[4]) ? 11'b00001100000 : node4213;
												assign node4213 = (inp[9]) ? 11'b00000000011 : 11'b00001000011;
								assign node4217 = (inp[9]) ? node4241 : node4218;
									assign node4218 = (inp[4]) ? node4230 : node4219;
										assign node4219 = (inp[3]) ? node4225 : node4220;
											assign node4220 = (inp[10]) ? 11'b10100000000 : node4221;
												assign node4221 = (inp[0]) ? 11'b00110000010 : 11'b00100000010;
											assign node4225 = (inp[0]) ? 11'b00010000000 : node4226;
												assign node4226 = (inp[10]) ? 11'b00000000100 : 11'b10000000010;
										assign node4230 = (inp[0]) ? node4238 : node4231;
											assign node4231 = (inp[3]) ? node4235 : node4232;
												assign node4232 = (inp[10]) ? 11'b10001110100 : 11'b00011100110;
												assign node4235 = (inp[10]) ? 11'b00100100010 : 11'b10101100100;
											assign node4238 = (inp[10]) ? 11'b00110100010 : 11'b00011110000;
									assign node4241 = (inp[4]) ? node4255 : node4242;
										assign node4242 = (inp[0]) ? node4248 : node4243;
											assign node4243 = (inp[10]) ? node4245 : 11'b00111100010;
												assign node4245 = (inp[3]) ? 11'b00011110110 : 11'b10111110100;
											assign node4248 = (inp[3]) ? node4252 : node4249;
												assign node4249 = (inp[10]) ? 11'b00101110000 : 11'b00101100110;
												assign node4252 = (inp[10]) ? 11'b00001100010 : 11'b00001110000;
										assign node4255 = (inp[10]) ? node4263 : node4256;
											assign node4256 = (inp[3]) ? node4260 : node4257;
												assign node4257 = (inp[0]) ? 11'b00010110100 : 11'b00000100110;
												assign node4260 = (inp[0]) ? 11'b00100100000 : 11'b10110110000;
											assign node4263 = (inp[3]) ? 11'b00000100010 : 11'b00000110010;
							assign node4266 = (inp[0]) ? node4318 : node4267;
								assign node4267 = (inp[10]) ? node4297 : node4268;
									assign node4268 = (inp[3]) ? node4284 : node4269;
										assign node4269 = (inp[4]) ? node4277 : node4270;
											assign node4270 = (inp[9]) ? node4274 : node4271;
												assign node4271 = (inp[8]) ? 11'b00110100000 : 11'b00111100010;
												assign node4274 = (inp[8]) ? 11'b00001110000 : 11'b00010110010;
											assign node4277 = (inp[9]) ? node4281 : node4278;
												assign node4278 = (inp[8]) ? 11'b00001100100 : 11'b00110100100;
												assign node4281 = (inp[8]) ? 11'b00110110100 : 11'b00101110100;
										assign node4284 = (inp[4]) ? node4290 : node4285;
											assign node4285 = (inp[9]) ? node4287 : 11'b10101110010;
												assign node4287 = (inp[8]) ? 11'b10001100100 : 11'b10010100100;
											assign node4290 = (inp[9]) ? node4294 : node4291;
												assign node4291 = (inp[8]) ? 11'b10110100110 : 11'b10010100100;
												assign node4294 = (inp[8]) ? 11'b10110110010 : 11'b10111110010;
									assign node4297 = (inp[4]) ? node4309 : node4298;
										assign node4298 = (inp[3]) ? node4304 : node4299;
											assign node4299 = (inp[9]) ? node4301 : 11'b10011100010;
												assign node4301 = (inp[8]) ? 11'b10101110110 : 11'b10000110100;
											assign node4304 = (inp[8]) ? 11'b00101110110 : node4305;
												assign node4305 = (inp[9]) ? 11'b00100110110 : 11'b00110110110;
										assign node4309 = (inp[3]) ? node4313 : node4310;
											assign node4310 = (inp[9]) ? 11'b10011110010 : 11'b10011110110;
											assign node4313 = (inp[8]) ? 11'b00010110000 : node4314;
												assign node4314 = (inp[9]) ? 11'b00011110000 : 11'b00001110010;
								assign node4318 = (inp[10]) ? node4342 : node4319;
									assign node4319 = (inp[9]) ? node4331 : node4320;
										assign node4320 = (inp[4]) ? node4326 : node4321;
											assign node4321 = (inp[3]) ? node4323 : 11'b00100110000;
												assign node4323 = (inp[8]) ? 11'b00000100000 : 11'b00011100000;
											assign node4326 = (inp[3]) ? node4328 : 11'b00101110000;
												assign node4328 = (inp[8]) ? 11'b00100110010 : 11'b00100110000;
										assign node4331 = (inp[4]) ? node4337 : node4332;
											assign node4332 = (inp[3]) ? node4334 : 11'b00100110110;
												assign node4334 = (inp[8]) ? 11'b00111110010 : 11'b00110110000;
											assign node4337 = (inp[3]) ? node4339 : 11'b00100100100;
												assign node4339 = (inp[8]) ? 11'b00100100010 : 11'b00101100010;
									assign node4342 = (inp[3]) ? node4352 : node4343;
										assign node4343 = (inp[4]) ? node4345 : 11'b00011110100;
											assign node4345 = (inp[8]) ? node4349 : node4346;
												assign node4346 = (inp[9]) ? 11'b00101100010 : 11'b00111100110;
												assign node4349 = (inp[9]) ? 11'b00000100010 : 11'b00000100110;
										assign node4352 = (inp[8]) ? node4358 : node4353;
											assign node4353 = (inp[4]) ? 11'b00011100000 : node4354;
												assign node4354 = (inp[9]) ? 11'b00010100010 : 11'b00100100010;
											assign node4358 = (inp[4]) ? 11'b00000100000 : node4359;
												assign node4359 = (inp[9]) ? 11'b00011100000 : 11'b00111100000;
						assign node4363 = (inp[0]) ? node4455 : node4364;
							assign node4364 = (inp[11]) ? node4408 : node4365;
								assign node4365 = (inp[4]) ? node4387 : node4366;
									assign node4366 = (inp[8]) ? node4376 : node4367;
										assign node4367 = (inp[10]) ? node4373 : node4368;
											assign node4368 = (inp[3]) ? 11'b10100110110 : node4369;
												assign node4369 = (inp[9]) ? 11'b00110110010 : 11'b00101110000;
											assign node4373 = (inp[3]) ? 11'b00010110100 : 11'b10000110010;
										assign node4376 = (inp[10]) ? node4384 : node4377;
											assign node4377 = (inp[3]) ? node4381 : node4378;
												assign node4378 = (inp[9]) ? 11'b00101010000 : 11'b00100110000;
												assign node4381 = (inp[9]) ? 11'b10101010110 : 11'b10101010010;
											assign node4384 = (inp[9]) ? 11'b00001000100 : 11'b00001010100;
									assign node4387 = (inp[8]) ? node4399 : node4388;
										assign node4388 = (inp[3]) ? node4394 : node4389;
											assign node4389 = (inp[10]) ? 11'b10110010010 : node4390;
												assign node4390 = (inp[9]) ? 11'b00001010110 : 11'b00111010110;
											assign node4394 = (inp[10]) ? node4396 : 11'b10101000000;
												assign node4396 = (inp[9]) ? 11'b00010000010 : 11'b00101010010;
										assign node4399 = (inp[10]) ? node4403 : node4400;
											assign node4400 = (inp[3]) ? 11'b10010000010 : 11'b00010010110;
											assign node4403 = (inp[3]) ? node4405 : 11'b10010010000;
												assign node4405 = (inp[9]) ? 11'b00010000000 : 11'b00110010000;
								assign node4408 = (inp[4]) ? node4434 : node4409;
									assign node4409 = (inp[9]) ? node4423 : node4410;
										assign node4410 = (inp[8]) ? node4418 : node4411;
											assign node4411 = (inp[10]) ? node4415 : node4412;
												assign node4412 = (inp[3]) ? 11'b10010000000 : 11'b00110010000;
												assign node4415 = (inp[3]) ? 11'b00100000110 : 11'b10000010010;
											assign node4418 = (inp[10]) ? 11'b10111010000 : node4419;
												assign node4419 = (inp[3]) ? 11'b10111000010 : 11'b00111010010;
										assign node4423 = (inp[10]) ? node4429 : node4424;
											assign node4424 = (inp[3]) ? node4426 : 11'b00111000010;
												assign node4426 = (inp[8]) ? 11'b10011010110 : 11'b10111010110;
											assign node4429 = (inp[3]) ? node4431 : 11'b10011000100;
												assign node4431 = (inp[8]) ? 11'b00011000100 : 11'b00111000100;
									assign node4434 = (inp[9]) ? node4444 : node4435;
										assign node4435 = (inp[8]) ? node4439 : node4436;
											assign node4436 = (inp[10]) ? 11'b10101000110 : 11'b00101010100;
											assign node4439 = (inp[10]) ? 11'b10010000100 : node4440;
												assign node4440 = (inp[3]) ? 11'b10010010110 : 11'b00010010110;
										assign node4444 = (inp[10]) ? node4450 : node4445;
											assign node4445 = (inp[3]) ? 11'b10010000010 : node4446;
												assign node4446 = (inp[8]) ? 11'b00010000110 : 11'b00110000110;
											assign node4450 = (inp[3]) ? 11'b00010000000 : node4451;
												assign node4451 = (inp[8]) ? 11'b10010000000 : 11'b10110000000;
							assign node4455 = (inp[3]) ? node4505 : node4456;
								assign node4456 = (inp[10]) ? node4480 : node4457;
									assign node4457 = (inp[9]) ? node4467 : node4458;
										assign node4458 = (inp[11]) ? node4464 : node4459;
											assign node4459 = (inp[8]) ? node4461 : 11'b00101000010;
												assign node4461 = (inp[4]) ? 11'b00010000010 : 11'b00111000010;
											assign node4464 = (inp[8]) ? 11'b00101010010 : 11'b00111010010;
										assign node4467 = (inp[11]) ? node4475 : node4468;
											assign node4468 = (inp[4]) ? node4472 : node4469;
												assign node4469 = (inp[8]) ? 11'b00111000110 : 11'b00000100110;
												assign node4472 = (inp[8]) ? 11'b00000010110 : 11'b00111010100;
											assign node4475 = (inp[4]) ? node4477 : 11'b00100010100;
												assign node4477 = (inp[8]) ? 11'b00000000110 : 11'b00100000110;
									assign node4480 = (inp[9]) ? node4494 : node4481;
										assign node4481 = (inp[8]) ? node4487 : node4482;
											assign node4482 = (inp[11]) ? node4484 : 11'b00100100100;
												assign node4484 = (inp[4]) ? 11'b00111000100 : 11'b00010010110;
											assign node4487 = (inp[4]) ? node4491 : node4488;
												assign node4488 = (inp[11]) ? 11'b00101010100 : 11'b00011000100;
												assign node4491 = (inp[11]) ? 11'b00000000100 : 11'b00100010100;
										assign node4494 = (inp[8]) ? node4500 : node4495;
											assign node4495 = (inp[11]) ? 11'b00101000010 : node4496;
												assign node4496 = (inp[4]) ? 11'b00100010010 : 11'b00110110000;
											assign node4500 = (inp[4]) ? node4502 : 11'b00011010000;
												assign node4502 = (inp[11]) ? 11'b00000000000 : 11'b00000010000;
								assign node4505 = (inp[10]) ? node4527 : node4506;
									assign node4506 = (inp[4]) ? node4518 : node4507;
										assign node4507 = (inp[9]) ? node4515 : node4508;
											assign node4508 = (inp[8]) ? node4512 : node4509;
												assign node4509 = (inp[11]) ? 11'b00110000010 : 11'b00110100010;
												assign node4512 = (inp[11]) ? 11'b00101000010 : 11'b00111000010;
											assign node4515 = (inp[11]) ? 11'b00001010010 : 11'b00110110000;
										assign node4518 = (inp[9]) ? node4522 : node4519;
											assign node4519 = (inp[11]) ? 11'b00000010010 : 11'b00100010010;
											assign node4522 = (inp[8]) ? 11'b00000000010 : node4523;
												assign node4523 = (inp[11]) ? 11'b00000000010 : 11'b00011000000;
									assign node4527 = (inp[9]) ? node4539 : node4528;
										assign node4528 = (inp[8]) ? node4534 : node4529;
											assign node4529 = (inp[4]) ? node4531 : 11'b00110000000;
												assign node4531 = (inp[11]) ? 11'b00011000000 : 11'b00111000010;
											assign node4534 = (inp[11]) ? node4536 : 11'b00011000000;
												assign node4536 = (inp[4]) ? 11'b00000000000 : 11'b00101000000;
										assign node4539 = (inp[4]) ? node4543 : node4540;
											assign node4540 = (inp[11]) ? 11'b00001000000 : 11'b00011000010;
											assign node4543 = (inp[8]) ? 11'b00000000000 : node4544;
												assign node4544 = (inp[11]) ? 11'b00000000000 : 11'b00000000010;
			assign node4548 = (inp[6]) ? node5306 : node4549;
				assign node4549 = (inp[2]) ? node4927 : node4550;
					assign node4550 = (inp[5]) ? node4738 : node4551;
						assign node4551 = (inp[0]) ? node4643 : node4552;
							assign node4552 = (inp[10]) ? node4602 : node4553;
								assign node4553 = (inp[3]) ? node4575 : node4554;
									assign node4554 = (inp[4]) ? node4562 : node4555;
										assign node4555 = (inp[8]) ? node4559 : node4556;
											assign node4556 = (inp[9]) ? 11'b00111110011 : 11'b00011100011;
											assign node4559 = (inp[9]) ? 11'b00000000001 : 11'b00010100001;
										assign node4562 = (inp[11]) ? node4570 : node4563;
											assign node4563 = (inp[8]) ? node4567 : node4564;
												assign node4564 = (inp[9]) ? 11'b00110100111 : 11'b00010100111;
												assign node4567 = (inp[9]) ? 11'b00101100101 : 11'b00111100101;
											assign node4570 = (inp[8]) ? 11'b00011110111 : node4571;
												assign node4571 = (inp[9]) ? 11'b00000110101 : 11'b00001100101;
									assign node4575 = (inp[4]) ? node4589 : node4576;
										assign node4576 = (inp[8]) ? node4584 : node4577;
											assign node4577 = (inp[9]) ? node4581 : node4578;
												assign node4578 = (inp[11]) ? 11'b10011110011 : 11'b10011100011;
												assign node4581 = (inp[11]) ? 11'b10111100111 : 11'b10011100111;
											assign node4584 = (inp[11]) ? node4586 : 11'b10110000011;
												assign node4586 = (inp[9]) ? 11'b10110100101 : 11'b10110110001;
										assign node4589 = (inp[9]) ? node4597 : node4590;
											assign node4590 = (inp[8]) ? node4594 : node4591;
												assign node4591 = (inp[11]) ? 11'b10100100111 : 11'b10010100111;
												assign node4594 = (inp[11]) ? 11'b10001100111 : 11'b10011100111;
											assign node4597 = (inp[8]) ? 11'b10001110001 : node4598;
												assign node4598 = (inp[11]) ? 11'b10000110011 : 11'b10110110011;
								assign node4602 = (inp[3]) ? node4618 : node4603;
									assign node4603 = (inp[4]) ? node4609 : node4604;
										assign node4604 = (inp[8]) ? 11'b10100100001 : node4605;
											assign node4605 = (inp[9]) ? 11'b10011110101 : 11'b10011100001;
										assign node4609 = (inp[8]) ? node4613 : node4610;
											assign node4610 = (inp[11]) ? 11'b10100110111 : 11'b10010110101;
											assign node4613 = (inp[9]) ? 11'b10101110011 : node4614;
												assign node4614 = (inp[11]) ? 11'b10101110101 : 11'b10111110111;
									assign node4618 = (inp[4]) ? node4632 : node4619;
										assign node4619 = (inp[8]) ? node4627 : node4620;
											assign node4620 = (inp[9]) ? node4624 : node4621;
												assign node4621 = (inp[11]) ? 11'b00011110101 : 11'b00011100101;
												assign node4624 = (inp[11]) ? 11'b00001110101 : 11'b00011110101;
											assign node4627 = (inp[11]) ? node4629 : 11'b00110000101;
												assign node4629 = (inp[9]) ? 11'b00111110111 : 11'b00000110111;
										assign node4632 = (inp[9]) ? node4636 : node4633;
											assign node4633 = (inp[8]) ? 11'b00001100011 : 11'b00110100001;
											assign node4636 = (inp[11]) ? node4640 : node4637;
												assign node4637 = (inp[8]) ? 11'b00110110011 : 11'b00110110001;
												assign node4640 = (inp[8]) ? 11'b00101110001 : 11'b00100110001;
							assign node4643 = (inp[10]) ? node4691 : node4644;
								assign node4644 = (inp[9]) ? node4670 : node4645;
									assign node4645 = (inp[11]) ? node4659 : node4646;
										assign node4646 = (inp[3]) ? node4652 : node4647;
											assign node4647 = (inp[8]) ? node4649 : 11'b00000100011;
												assign node4649 = (inp[4]) ? 11'b00101100001 : 11'b00100000011;
											assign node4652 = (inp[4]) ? node4656 : node4653;
												assign node4653 = (inp[8]) ? 11'b00000000011 : 11'b00001100011;
												assign node4656 = (inp[8]) ? 11'b00001110011 : 11'b00000110011;
										assign node4659 = (inp[4]) ? node4665 : node4660;
											assign node4660 = (inp[8]) ? node4662 : 11'b00001110011;
												assign node4662 = (inp[3]) ? 11'b00010100001 : 11'b00100110001;
											assign node4665 = (inp[8]) ? node4667 : 11'b00110110011;
												assign node4667 = (inp[3]) ? 11'b00111110001 : 11'b00111110011;
									assign node4670 = (inp[3]) ? node4682 : node4671;
										assign node4671 = (inp[8]) ? node4679 : node4672;
											assign node4672 = (inp[4]) ? node4676 : node4673;
												assign node4673 = (inp[11]) ? 11'b00101110111 : 11'b00001100111;
												assign node4676 = (inp[11]) ? 11'b00010100111 : 11'b00100110111;
											assign node4679 = (inp[11]) ? 11'b00000110111 : 11'b00011110101;
										assign node4682 = (inp[4]) ? node4684 : 11'b00011110011;
											assign node4684 = (inp[11]) ? node4688 : node4685;
												assign node4685 = (inp[8]) ? 11'b00110100011 : 11'b00100100011;
												assign node4688 = (inp[8]) ? 11'b00111100011 : 11'b00110100011;
								assign node4691 = (inp[3]) ? node4719 : node4692;
									assign node4692 = (inp[9]) ? node4706 : node4693;
										assign node4693 = (inp[8]) ? node4699 : node4694;
											assign node4694 = (inp[4]) ? 11'b00110100101 : node4695;
												assign node4695 = (inp[11]) ? 11'b00001110101 : 11'b00001100101;
											assign node4699 = (inp[4]) ? node4703 : node4700;
												assign node4700 = (inp[11]) ? 11'b00110110111 : 11'b00100000101;
												assign node4703 = (inp[11]) ? 11'b00001100101 : 11'b00101110111;
										assign node4706 = (inp[11]) ? node4712 : node4707;
											assign node4707 = (inp[4]) ? 11'b00000110011 : node4708;
												assign node4708 = (inp[8]) ? 11'b00111110001 : 11'b00001110001;
											assign node4712 = (inp[8]) ? node4716 : node4713;
												assign node4713 = (inp[4]) ? 11'b00110100001 : 11'b00011100001;
												assign node4716 = (inp[4]) ? 11'b00011100001 : 11'b00100100001;
									assign node4719 = (inp[8]) ? node4727 : node4720;
										assign node4720 = (inp[4]) ? node4724 : node4721;
											assign node4721 = (inp[11]) ? 11'b00101100001 : 11'b00001100001;
											assign node4724 = (inp[9]) ? 11'b00000100001 : 11'b00100100001;
										assign node4727 = (inp[4]) ? node4735 : node4728;
											assign node4728 = (inp[9]) ? node4732 : node4729;
												assign node4729 = (inp[11]) ? 11'b00110100011 : 11'b00010000001;
												assign node4732 = (inp[11]) ? 11'b00011100011 : 11'b00001100001;
											assign node4735 = (inp[11]) ? 11'b00001100001 : 11'b00000100011;
						assign node4738 = (inp[0]) ? node4838 : node4739;
							assign node4739 = (inp[11]) ? node4789 : node4740;
								assign node4740 = (inp[8]) ? node4768 : node4741;
									assign node4741 = (inp[10]) ? node4755 : node4742;
										assign node4742 = (inp[4]) ? node4750 : node4743;
											assign node4743 = (inp[3]) ? node4747 : node4744;
												assign node4744 = (inp[9]) ? 11'b00011010001 : 11'b00010110001;
												assign node4747 = (inp[9]) ? 11'b10011010111 : 11'b10011010011;
											assign node4750 = (inp[3]) ? 11'b10101010101 : node4751;
												assign node4751 = (inp[9]) ? 11'b00100010101 : 11'b00001010101;
										assign node4755 = (inp[4]) ? node4761 : node4756;
											assign node4756 = (inp[9]) ? node4758 : 11'b00111010101;
												assign node4758 = (inp[3]) ? 11'b00001000111 : 11'b10111000111;
											assign node4761 = (inp[9]) ? node4765 : node4762;
												assign node4762 = (inp[3]) ? 11'b00000010011 : 11'b10000000111;
												assign node4765 = (inp[3]) ? 11'b00110000011 : 11'b10010010011;
									assign node4768 = (inp[4]) ? node4780 : node4769;
										assign node4769 = (inp[10]) ? node4775 : node4770;
											assign node4770 = (inp[3]) ? 11'b10010110011 : node4771;
												assign node4771 = (inp[9]) ? 11'b00000110001 : 11'b00011110001;
											assign node4775 = (inp[3]) ? node4777 : 11'b10010100111;
												assign node4777 = (inp[9]) ? 11'b00110100111 : 11'b00100110111;
										assign node4780 = (inp[9]) ? node4786 : node4781;
											assign node4781 = (inp[3]) ? 11'b00011010011 : node4782;
												assign node4782 = (inp[10]) ? 11'b10010100101 : 11'b00100110111;
											assign node4786 = (inp[10]) ? 11'b10101010001 : 11'b10101000011;
								assign node4789 = (inp[9]) ? node4815 : node4790;
									assign node4790 = (inp[10]) ? node4802 : node4791;
										assign node4791 = (inp[3]) ? node4797 : node4792;
											assign node4792 = (inp[4]) ? node4794 : 11'b00011010011;
												assign node4794 = (inp[8]) ? 11'b00110010101 : 11'b00011010111;
											assign node4797 = (inp[4]) ? node4799 : 11'b10110000001;
												assign node4799 = (inp[8]) ? 11'b10110010101 : 11'b10111010101;
										assign node4802 = (inp[3]) ? node4808 : node4803;
											assign node4803 = (inp[4]) ? node4805 : 11'b10001010011;
												assign node4805 = (inp[8]) ? 11'b10100000101 : 11'b10011000101;
											assign node4808 = (inp[4]) ? node4812 : node4809;
												assign node4809 = (inp[8]) ? 11'b00011000101 : 11'b00001000111;
												assign node4812 = (inp[8]) ? 11'b00100000011 : 11'b00110000011;
									assign node4815 = (inp[10]) ? node4829 : node4816;
										assign node4816 = (inp[3]) ? node4824 : node4817;
											assign node4817 = (inp[4]) ? node4821 : node4818;
												assign node4818 = (inp[8]) ? 11'b00011000001 : 11'b00101000011;
												assign node4821 = (inp[8]) ? 11'b00110000111 : 11'b00000000111;
											assign node4824 = (inp[4]) ? node4826 : 11'b10110010111;
												assign node4826 = (inp[8]) ? 11'b10110000001 : 11'b10100000011;
										assign node4829 = (inp[4]) ? node4833 : node4830;
											assign node4830 = (inp[3]) ? 11'b00100000111 : 11'b10100000111;
											assign node4833 = (inp[8]) ? node4835 : 11'b10000000001;
												assign node4835 = (inp[3]) ? 11'b00100000001 : 11'b10100000001;
							assign node4838 = (inp[11]) ? node4890 : node4839;
								assign node4839 = (inp[8]) ? node4863 : node4840;
									assign node4840 = (inp[4]) ? node4852 : node4841;
										assign node4841 = (inp[9]) ? node4847 : node4842;
											assign node4842 = (inp[10]) ? node4844 : 11'b00000100001;
												assign node4844 = (inp[3]) ? 11'b00001000001 : 11'b00101000111;
											assign node4847 = (inp[3]) ? 11'b00101010011 : node4848;
												assign node4848 = (inp[10]) ? 11'b00101010011 : 11'b00001000101;
										assign node4852 = (inp[9]) ? node4856 : node4853;
											assign node4853 = (inp[10]) ? 11'b00110000001 : 11'b00111000001;
											assign node4856 = (inp[3]) ? node4860 : node4857;
												assign node4857 = (inp[10]) ? 11'b00100010011 : 11'b00110010101;
												assign node4860 = (inp[10]) ? 11'b00000000011 : 11'b00000000001;
									assign node4863 = (inp[4]) ? node4879 : node4864;
										assign node4864 = (inp[10]) ? node4872 : node4865;
											assign node4865 = (inp[9]) ? node4869 : node4866;
												assign node4866 = (inp[3]) ? 11'b00100100011 : 11'b00101100001;
												assign node4869 = (inp[3]) ? 11'b00100110001 : 11'b00110100101;
											assign node4872 = (inp[9]) ? node4876 : node4873;
												assign node4873 = (inp[3]) ? 11'b00010100001 : 11'b00010100111;
												assign node4876 = (inp[3]) ? 11'b00010100011 : 11'b00000110011;
										assign node4879 = (inp[9]) ? node4885 : node4880;
											assign node4880 = (inp[10]) ? 11'b00100110101 : node4881;
												assign node4881 = (inp[3]) ? 11'b00110110001 : 11'b00010100001;
											assign node4885 = (inp[10]) ? node4887 : 11'b00011000001;
												assign node4887 = (inp[3]) ? 11'b00001000001 : 11'b00001010001;
								assign node4890 = (inp[4]) ? node4906 : node4891;
									assign node4891 = (inp[10]) ? node4903 : node4892;
										assign node4892 = (inp[3]) ? node4898 : node4893;
											assign node4893 = (inp[8]) ? node4895 : 11'b00000010001;
												assign node4895 = (inp[9]) ? 11'b00001010101 : 11'b00101010011;
											assign node4898 = (inp[9]) ? node4900 : 11'b00111000011;
												assign node4900 = (inp[8]) ? 11'b00010010011 : 11'b00011010001;
										assign node4903 = (inp[9]) ? 11'b00111000011 : 11'b00011010111;
									assign node4906 = (inp[9]) ? node4920 : node4907;
										assign node4907 = (inp[10]) ? node4913 : node4908;
											assign node4908 = (inp[8]) ? 11'b00010010001 : node4909;
												assign node4909 = (inp[3]) ? 11'b00001010001 : 11'b00101010011;
											assign node4913 = (inp[3]) ? node4917 : node4914;
												assign node4914 = (inp[8]) ? 11'b00010000111 : 11'b00101000101;
												assign node4917 = (inp[8]) ? 11'b00000000011 : 11'b00010000011;
										assign node4920 = (inp[8]) ? 11'b00010000001 : node4921;
											assign node4921 = (inp[3]) ? 11'b00010000001 : node4922;
												assign node4922 = (inp[10]) ? 11'b00110000001 : 11'b00110000111;
					assign node4927 = (inp[8]) ? node5119 : node4928;
						assign node4928 = (inp[5]) ? node5022 : node4929;
							assign node4929 = (inp[11]) ? node4975 : node4930;
								assign node4930 = (inp[0]) ? node4954 : node4931;
									assign node4931 = (inp[10]) ? node4941 : node4932;
										assign node4932 = (inp[9]) ? 11'b00010000111 : node4933;
											assign node4933 = (inp[4]) ? node4937 : node4934;
												assign node4934 = (inp[3]) ? 11'b10111000011 : 11'b00111000011;
												assign node4937 = (inp[3]) ? 11'b10111000101 : 11'b00111000101;
										assign node4941 = (inp[4]) ? node4949 : node4942;
											assign node4942 = (inp[3]) ? node4946 : node4943;
												assign node4943 = (inp[9]) ? 11'b10101010111 : 11'b10101000011;
												assign node4946 = (inp[9]) ? 11'b00101010111 : 11'b00101000101;
											assign node4949 = (inp[3]) ? 11'b00010000011 : node4950;
												assign node4950 = (inp[9]) ? 11'b10000000001 : 11'b10101010101;
									assign node4954 = (inp[4]) ? node4968 : node4955;
										assign node4955 = (inp[3]) ? node4961 : node4956;
											assign node4956 = (inp[10]) ? 11'b00011000101 : node4957;
												assign node4957 = (inp[9]) ? 11'b00001000101 : 11'b00001000011;
											assign node4961 = (inp[10]) ? node4965 : node4962;
												assign node4962 = (inp[9]) ? 11'b00011010011 : 11'b00011000011;
												assign node4965 = (inp[9]) ? 11'b00001000011 : 11'b00001000001;
										assign node4968 = (inp[3]) ? 11'b00000000001 : node4969;
											assign node4969 = (inp[10]) ? 11'b00010010111 : node4970;
												assign node4970 = (inp[9]) ? 11'b00100010111 : 11'b00001000001;
								assign node4975 = (inp[4]) ? node5001 : node4976;
									assign node4976 = (inp[9]) ? node4990 : node4977;
										assign node4977 = (inp[0]) ? node4985 : node4978;
											assign node4978 = (inp[3]) ? node4982 : node4979;
												assign node4979 = (inp[10]) ? 11'b10100000011 : 11'b00110000011;
												assign node4982 = (inp[10]) ? 11'b00110010101 : 11'b10100010011;
											assign node4985 = (inp[10]) ? 11'b00000010111 : node4986;
												assign node4986 = (inp[3]) ? 11'b00010000011 : 11'b00010010011;
										assign node4990 = (inp[10]) ? node4996 : node4991;
											assign node4991 = (inp[0]) ? 11'b00110010101 : node4992;
												assign node4992 = (inp[3]) ? 11'b10000000101 : 11'b00000010001;
											assign node4996 = (inp[0]) ? node4998 : 11'b10011110110;
												assign node4998 = (inp[3]) ? 11'b00011100010 : 11'b00001100010;
									assign node5001 = (inp[0]) ? node5015 : node5002;
										assign node5002 = (inp[9]) ? node5008 : node5003;
											assign node5003 = (inp[10]) ? node5005 : 11'b10011100100;
												assign node5005 = (inp[3]) ? 11'b00001110000 : 11'b10011110100;
											assign node5008 = (inp[10]) ? node5012 : node5009;
												assign node5009 = (inp[3]) ? 11'b10111110010 : 11'b00101110110;
												assign node5012 = (inp[3]) ? 11'b00001110000 : 11'b10001110010;
										assign node5015 = (inp[9]) ? node5019 : node5016;
											assign node5016 = (inp[3]) ? 11'b00101110000 : 11'b00011110000;
											assign node5019 = (inp[10]) ? 11'b00111100000 : 11'b00101100010;
							assign node5022 = (inp[0]) ? node5074 : node5023;
								assign node5023 = (inp[11]) ? node5051 : node5024;
									assign node5024 = (inp[10]) ? node5036 : node5025;
										assign node5025 = (inp[3]) ? node5031 : node5026;
											assign node5026 = (inp[4]) ? 11'b00100110110 : node5027;
												assign node5027 = (inp[9]) ? 11'b00110110000 : 11'b00111110000;
											assign node5031 = (inp[9]) ? 11'b10100110100 : node5032;
												assign node5032 = (inp[4]) ? 11'b10010110110 : 11'b10110110010;
										assign node5036 = (inp[3]) ? node5044 : node5037;
											assign node5037 = (inp[4]) ? node5041 : node5038;
												assign node5038 = (inp[9]) ? 11'b10010100100 : 11'b10000110010;
												assign node5041 = (inp[9]) ? 11'b10101110010 : 11'b10110100100;
											assign node5044 = (inp[4]) ? node5048 : node5045;
												assign node5045 = (inp[9]) ? 11'b00110100110 : 11'b00010110110;
												assign node5048 = (inp[9]) ? 11'b00011100010 : 11'b00100110000;
									assign node5051 = (inp[4]) ? node5065 : node5052;
										assign node5052 = (inp[9]) ? node5060 : node5053;
											assign node5053 = (inp[3]) ? node5057 : node5054;
												assign node5054 = (inp[10]) ? 11'b10011110000 : 11'b00111110000;
												assign node5057 = (inp[10]) ? 11'b00111100110 : 11'b10001100000;
											assign node5060 = (inp[10]) ? node5062 : 11'b10111110110;
												assign node5062 = (inp[3]) ? 11'b00101100100 : 11'b10001100110;
										assign node5065 = (inp[9]) ? node5071 : node5066;
											assign node5066 = (inp[10]) ? 11'b00010100010 : node5067;
												assign node5067 = (inp[3]) ? 11'b10001110100 : 11'b00111110100;
											assign node5071 = (inp[3]) ? 11'b10010100000 : 11'b10110100000;
								assign node5074 = (inp[3]) ? node5098 : node5075;
									assign node5075 = (inp[9]) ? node5083 : node5076;
										assign node5076 = (inp[11]) ? node5080 : node5077;
											assign node5077 = (inp[10]) ? 11'b00110100110 : 11'b00110100010;
											assign node5080 = (inp[4]) ? 11'b00100100110 : 11'b00001110100;
										assign node5083 = (inp[10]) ? node5091 : node5084;
											assign node5084 = (inp[11]) ? node5088 : node5085;
												assign node5085 = (inp[4]) ? 11'b00100110100 : 11'b00010100100;
												assign node5088 = (inp[4]) ? 11'b00110100100 : 11'b00111110110;
											assign node5091 = (inp[11]) ? node5095 : node5092;
												assign node5092 = (inp[4]) ? 11'b00111110010 : 11'b00100110000;
												assign node5095 = (inp[4]) ? 11'b00110100000 : 11'b00111100000;
									assign node5098 = (inp[9]) ? node5108 : node5099;
										assign node5099 = (inp[4]) ? node5103 : node5100;
											assign node5100 = (inp[11]) ? 11'b00111100010 : 11'b00110100010;
											assign node5103 = (inp[11]) ? node5105 : 11'b00100110010;
												assign node5105 = (inp[10]) ? 11'b00010100010 : 11'b00010110010;
										assign node5108 = (inp[11]) ? node5116 : node5109;
											assign node5109 = (inp[4]) ? node5113 : node5110;
												assign node5110 = (inp[10]) ? 11'b00010100010 : 11'b00110110000;
												assign node5113 = (inp[10]) ? 11'b00001100010 : 11'b00011100010;
											assign node5116 = (inp[4]) ? 11'b00000100000 : 11'b00001100000;
						assign node5119 = (inp[11]) ? node5219 : node5120;
							assign node5120 = (inp[4]) ? node5174 : node5121;
								assign node5121 = (inp[5]) ? node5149 : node5122;
									assign node5122 = (inp[10]) ? node5136 : node5123;
										assign node5123 = (inp[3]) ? node5129 : node5124;
											assign node5124 = (inp[9]) ? node5126 : 11'b00100100010;
												assign node5126 = (inp[0]) ? 11'b00110100100 : 11'b00100100000;
											assign node5129 = (inp[0]) ? node5133 : node5130;
												assign node5130 = (inp[9]) ? 11'b10010100100 : 11'b10000100010;
												assign node5133 = (inp[9]) ? 11'b00000110000 : 11'b00010100010;
										assign node5136 = (inp[9]) ? node5142 : node5137;
											assign node5137 = (inp[3]) ? 11'b00010100100 : node5138;
												assign node5138 = (inp[0]) ? 11'b00100100110 : 11'b10100100010;
											assign node5142 = (inp[3]) ? node5146 : node5143;
												assign node5143 = (inp[0]) ? 11'b00111010010 : 11'b10111010110;
												assign node5146 = (inp[0]) ? 11'b00001000010 : 11'b00001010110;
									assign node5149 = (inp[10]) ? node5163 : node5150;
										assign node5150 = (inp[0]) ? node5156 : node5151;
											assign node5151 = (inp[9]) ? 11'b00101010010 : node5152;
												assign node5152 = (inp[3]) ? 11'b10100010000 : 11'b00110010000;
											assign node5156 = (inp[3]) ? node5160 : node5157;
												assign node5157 = (inp[9]) ? 11'b00101000110 : 11'b00100000000;
												assign node5160 = (inp[9]) ? 11'b00111010000 : 11'b00111000010;
										assign node5163 = (inp[9]) ? node5171 : node5164;
											assign node5164 = (inp[0]) ? node5168 : node5165;
												assign node5165 = (inp[3]) ? 11'b00001010110 : 11'b10011010010;
												assign node5168 = (inp[3]) ? 11'b00011000010 : 11'b00001000110;
											assign node5171 = (inp[0]) ? 11'b00011000000 : 11'b10101000100;
								assign node5174 = (inp[3]) ? node5194 : node5175;
									assign node5175 = (inp[0]) ? node5185 : node5176;
										assign node5176 = (inp[10]) ? node5182 : node5177;
											assign node5177 = (inp[5]) ? 11'b00001010110 : node5178;
												assign node5178 = (inp[9]) ? 11'b00001000100 : 11'b00011000110;
											assign node5182 = (inp[9]) ? 11'b10101000010 : 11'b10101000110;
										assign node5185 = (inp[9]) ? node5189 : node5186;
											assign node5186 = (inp[10]) ? 11'b00101010100 : 11'b00101000010;
											assign node5189 = (inp[10]) ? 11'b00011010010 : node5190;
												assign node5190 = (inp[5]) ? 11'b00011010100 : 11'b00001010100;
									assign node5194 = (inp[0]) ? node5208 : node5195;
										assign node5195 = (inp[10]) ? node5201 : node5196;
											assign node5196 = (inp[5]) ? 11'b10011000000 : node5197;
												assign node5197 = (inp[9]) ? 11'b10111010010 : 11'b10101000110;
											assign node5201 = (inp[9]) ? node5205 : node5202;
												assign node5202 = (inp[5]) ? 11'b00111010010 : 11'b00111000000;
												assign node5205 = (inp[5]) ? 11'b00011000000 : 11'b00011010010;
										assign node5208 = (inp[9]) ? node5214 : node5209;
											assign node5209 = (inp[5]) ? node5211 : 11'b00011010000;
												assign node5211 = (inp[10]) ? 11'b00101000010 : 11'b00101010010;
											assign node5214 = (inp[5]) ? 11'b00001000000 : node5215;
												assign node5215 = (inp[10]) ? 11'b00001000010 : 11'b00101000010;
							assign node5219 = (inp[3]) ? node5265 : node5220;
								assign node5220 = (inp[9]) ? node5244 : node5221;
									assign node5221 = (inp[5]) ? node5231 : node5222;
										assign node5222 = (inp[0]) ? node5226 : node5223;
											assign node5223 = (inp[10]) ? 11'b10011000000 : 11'b00111000000;
											assign node5226 = (inp[10]) ? 11'b00101010100 : node5227;
												assign node5227 = (inp[4]) ? 11'b00110010000 : 11'b00111010000;
										assign node5231 = (inp[4]) ? node5237 : node5232;
											assign node5232 = (inp[0]) ? 11'b00110010110 : node5233;
												assign node5233 = (inp[10]) ? 11'b10110010010 : 11'b00110010010;
											assign node5237 = (inp[10]) ? node5241 : node5238;
												assign node5238 = (inp[0]) ? 11'b00010010010 : 11'b00010010110;
												assign node5241 = (inp[0]) ? 11'b00010000110 : 11'b10010000110;
									assign node5244 = (inp[10]) ? node5254 : node5245;
										assign node5245 = (inp[5]) ? node5251 : node5246;
											assign node5246 = (inp[4]) ? node5248 : 11'b00000010110;
												assign node5248 = (inp[0]) ? 11'b00110000110 : 11'b00110010110;
											assign node5251 = (inp[4]) ? 11'b00010000100 : 11'b00110000000;
										assign node5254 = (inp[0]) ? node5260 : node5255;
											assign node5255 = (inp[5]) ? node5257 : 11'b10010010000;
												assign node5257 = (inp[4]) ? 11'b10010000000 : 11'b10010000100;
											assign node5260 = (inp[4]) ? 11'b00010000000 : node5261;
												assign node5261 = (inp[5]) ? 11'b00010000000 : 11'b00100000010;
								assign node5265 = (inp[5]) ? node5285 : node5266;
									assign node5266 = (inp[0]) ? node5278 : node5267;
										assign node5267 = (inp[10]) ? node5273 : node5268;
											assign node5268 = (inp[9]) ? node5270 : 11'b10001010000;
												assign node5270 = (inp[4]) ? 11'b10100010010 : 11'b10000000110;
											assign node5273 = (inp[9]) ? node5275 : 11'b00101010100;
												assign node5275 = (inp[4]) ? 11'b00000010000 : 11'b00010010100;
										assign node5278 = (inp[4]) ? 11'b00100010000 : node5279;
											assign node5279 = (inp[9]) ? 11'b00110010010 : node5280;
												assign node5280 = (inp[10]) ? 11'b00110000010 : 11'b00001000000;
									assign node5285 = (inp[9]) ? node5295 : node5286;
										assign node5286 = (inp[10]) ? node5290 : node5287;
											assign node5287 = (inp[0]) ? 11'b00000010010 : 11'b10000010110;
											assign node5290 = (inp[4]) ? 11'b00000000010 : node5291;
												assign node5291 = (inp[0]) ? 11'b00100000010 : 11'b00100000110;
										assign node5295 = (inp[4]) ? node5301 : node5296;
											assign node5296 = (inp[10]) ? node5298 : 11'b00000010000;
												assign node5298 = (inp[0]) ? 11'b00000000000 : 11'b00000000100;
											assign node5301 = (inp[0]) ? 11'b00000000000 : node5302;
												assign node5302 = (inp[10]) ? 11'b00000000000 : 11'b10000000000;
				assign node5306 = (inp[2]) ? node5682 : node5307;
					assign node5307 = (inp[8]) ? node5497 : node5308;
						assign node5308 = (inp[11]) ? node5404 : node5309;
							assign node5309 = (inp[3]) ? node5353 : node5310;
								assign node5310 = (inp[10]) ? node5334 : node5311;
									assign node5311 = (inp[4]) ? node5321 : node5312;
										assign node5312 = (inp[9]) ? node5316 : node5313;
											assign node5313 = (inp[5]) ? 11'b00010100000 : 11'b00011100010;
											assign node5316 = (inp[5]) ? 11'b00011100110 : node5317;
												assign node5317 = (inp[0]) ? 11'b00011100100 : 11'b00011100000;
										assign node5321 = (inp[9]) ? node5327 : node5322;
											assign node5322 = (inp[0]) ? node5324 : 11'b00001110100;
												assign node5324 = (inp[5]) ? 11'b00101100000 : 11'b00011100010;
											assign node5327 = (inp[5]) ? node5331 : node5328;
												assign node5328 = (inp[0]) ? 11'b00111110100 : 11'b00111100100;
												assign node5331 = (inp[0]) ? 11'b00101110110 : 11'b00111110110;
									assign node5334 = (inp[0]) ? node5346 : node5335;
										assign node5335 = (inp[5]) ? node5339 : node5336;
											assign node5336 = (inp[9]) ? 11'b10011110100 : 11'b10011100010;
											assign node5339 = (inp[4]) ? node5343 : node5340;
												assign node5340 = (inp[9]) ? 11'b10101100110 : 11'b10111110010;
												assign node5343 = (inp[9]) ? 11'b10011110010 : 11'b10011100100;
										assign node5346 = (inp[9]) ? 11'b00111110000 : node5347;
											assign node5347 = (inp[4]) ? 11'b00011110110 : node5348;
												assign node5348 = (inp[5]) ? 11'b00111100110 : 11'b00011100110;
								assign node5353 = (inp[0]) ? node5377 : node5354;
									assign node5354 = (inp[10]) ? node5368 : node5355;
										assign node5355 = (inp[5]) ? node5361 : node5356;
											assign node5356 = (inp[9]) ? node5358 : 11'b10001100110;
												assign node5358 = (inp[4]) ? 11'b10101110000 : 11'b10001100100;
											assign node5361 = (inp[9]) ? node5365 : node5362;
												assign node5362 = (inp[4]) ? 11'b10111110100 : 11'b10000110000;
												assign node5365 = (inp[4]) ? 11'b10001100010 : 11'b10011110110;
										assign node5368 = (inp[4]) ? node5370 : 11'b00101110110;
											assign node5370 = (inp[9]) ? node5374 : node5371;
												assign node5371 = (inp[5]) ? 11'b00001110000 : 11'b00101100010;
												assign node5374 = (inp[5]) ? 11'b00101100010 : 11'b00101110000;
									assign node5377 = (inp[10]) ? node5391 : node5378;
										assign node5378 = (inp[5]) ? node5384 : node5379;
											assign node5379 = (inp[9]) ? 11'b00001110000 : node5380;
												assign node5380 = (inp[4]) ? 11'b00001110010 : 11'b00001100010;
											assign node5384 = (inp[9]) ? node5388 : node5385;
												assign node5385 = (inp[4]) ? 11'b00111110000 : 11'b00100100000;
												assign node5388 = (inp[4]) ? 11'b00001100010 : 11'b00101110010;
										assign node5391 = (inp[9]) ? node5397 : node5392;
											assign node5392 = (inp[4]) ? node5394 : 11'b00001100010;
												assign node5394 = (inp[5]) ? 11'b00111100010 : 11'b00101100010;
											assign node5397 = (inp[4]) ? node5401 : node5398;
												assign node5398 = (inp[5]) ? 11'b00011100000 : 11'b00001100000;
												assign node5401 = (inp[5]) ? 11'b00001100010 : 11'b00001100000;
							assign node5404 = (inp[0]) ? node5458 : node5405;
								assign node5405 = (inp[5]) ? node5431 : node5406;
									assign node5406 = (inp[3]) ? node5416 : node5407;
										assign node5407 = (inp[9]) ? node5413 : node5408;
											assign node5408 = (inp[10]) ? 11'b10000100010 : node5409;
												assign node5409 = (inp[4]) ? 11'b00000100100 : 11'b00001100000;
											assign node5413 = (inp[4]) ? 11'b10110110000 : 11'b00100110010;
										assign node5416 = (inp[10]) ? node5424 : node5417;
											assign node5417 = (inp[4]) ? node5421 : node5418;
												assign node5418 = (inp[9]) ? 11'b10110100100 : 11'b10010110010;
												assign node5421 = (inp[9]) ? 11'b10000110010 : 11'b10110100110;
											assign node5424 = (inp[4]) ? node5428 : node5425;
												assign node5425 = (inp[9]) ? 11'b00010110100 : 11'b00010110110;
												assign node5428 = (inp[9]) ? 11'b00100110000 : 11'b00110110010;
									assign node5431 = (inp[4]) ? node5445 : node5432;
										assign node5432 = (inp[9]) ? node5438 : node5433;
											assign node5433 = (inp[3]) ? node5435 : 11'b10101110000;
												assign node5435 = (inp[10]) ? 11'b00011100100 : 11'b10111100000;
											assign node5438 = (inp[10]) ? node5442 : node5439;
												assign node5439 = (inp[3]) ? 11'b10001110100 : 11'b00101100000;
												assign node5442 = (inp[3]) ? 11'b00000100110 : 11'b10110100110;
										assign node5445 = (inp[3]) ? node5451 : node5446;
											assign node5446 = (inp[10]) ? 11'b10010100000 : node5447;
												assign node5447 = (inp[9]) ? 11'b00000100100 : 11'b00010110110;
											assign node5451 = (inp[10]) ? node5455 : node5452;
												assign node5452 = (inp[9]) ? 11'b10110100000 : 11'b10100110110;
												assign node5455 = (inp[9]) ? 11'b00100100000 : 11'b00110100000;
								assign node5458 = (inp[10]) ? node5482 : node5459;
									assign node5459 = (inp[9]) ? node5471 : node5460;
										assign node5460 = (inp[3]) ? node5468 : node5461;
											assign node5461 = (inp[4]) ? node5465 : node5462;
												assign node5462 = (inp[5]) ? 11'b00011110000 : 11'b00010110010;
												assign node5465 = (inp[5]) ? 11'b00110110010 : 11'b00000110000;
											assign node5468 = (inp[4]) ? 11'b00000110010 : 11'b00000100010;
										assign node5471 = (inp[3]) ? node5477 : node5472;
											assign node5472 = (inp[5]) ? node5474 : 11'b00000100110;
												assign node5474 = (inp[4]) ? 11'b00100100100 : 11'b00101110100;
											assign node5477 = (inp[5]) ? 11'b00010110010 : node5478;
												assign node5478 = (inp[4]) ? 11'b00110100000 : 11'b00100110000;
									assign node5482 = (inp[9]) ? node5492 : node5483;
										assign node5483 = (inp[5]) ? node5489 : node5484;
											assign node5484 = (inp[3]) ? node5486 : 11'b00100100110;
												assign node5486 = (inp[4]) ? 11'b00010100010 : 11'b00100100010;
											assign node5489 = (inp[3]) ? 11'b00111100000 : 11'b00110100100;
										assign node5492 = (inp[3]) ? node5494 : 11'b00100100000;
											assign node5494 = (inp[4]) ? 11'b00000100000 : 11'b00000100010;
						assign node5497 = (inp[5]) ? node5589 : node5498;
							assign node5498 = (inp[11]) ? node5544 : node5499;
								assign node5499 = (inp[4]) ? node5523 : node5500;
									assign node5500 = (inp[9]) ? node5510 : node5501;
										assign node5501 = (inp[0]) ? node5507 : node5502;
											assign node5502 = (inp[3]) ? 11'b10100100010 : node5503;
												assign node5503 = (inp[10]) ? 11'b10000100010 : 11'b00010100010;
											assign node5507 = (inp[10]) ? 11'b00010100010 : 11'b00000100010;
										assign node5510 = (inp[0]) ? node5516 : node5511;
											assign node5511 = (inp[3]) ? 11'b10110100100 : node5512;
												assign node5512 = (inp[10]) ? 11'b10010110100 : 11'b00000100010;
											assign node5516 = (inp[3]) ? node5520 : node5517;
												assign node5517 = (inp[10]) ? 11'b00100110000 : 11'b00100100110;
												assign node5520 = (inp[10]) ? 11'b00000100000 : 11'b00010110000;
									assign node5523 = (inp[9]) ? node5533 : node5524;
										assign node5524 = (inp[3]) ? node5528 : node5525;
											assign node5525 = (inp[10]) ? 11'b10100110100 : 11'b00110100000;
											assign node5528 = (inp[10]) ? 11'b00011000010 : node5529;
												assign node5529 = (inp[0]) ? 11'b00000110000 : 11'b10010100100;
										assign node5533 = (inp[10]) ? node5537 : node5534;
											assign node5534 = (inp[0]) ? 11'b00111000010 : 11'b00101000110;
											assign node5537 = (inp[3]) ? node5541 : node5538;
												assign node5538 = (inp[0]) ? 11'b00011010010 : 11'b10011000010;
												assign node5541 = (inp[0]) ? 11'b00001000010 : 11'b00101010010;
								assign node5544 = (inp[0]) ? node5564 : node5545;
									assign node5545 = (inp[3]) ? node5557 : node5546;
										assign node5546 = (inp[10]) ? node5550 : node5547;
											assign node5547 = (inp[4]) ? 11'b00001010110 : 11'b00001000010;
											assign node5550 = (inp[4]) ? node5554 : node5551;
												assign node5551 = (inp[9]) ? 11'b10001010100 : 11'b10101000000;
												assign node5554 = (inp[9]) ? 11'b10101010000 : 11'b10111010110;
										assign node5557 = (inp[10]) ? node5561 : node5558;
											assign node5558 = (inp[4]) ? 11'b10011010000 : 11'b10111010000;
											assign node5561 = (inp[9]) ? 11'b00101010000 : 11'b00001010100;
									assign node5564 = (inp[10]) ? node5578 : node5565;
										assign node5565 = (inp[9]) ? node5573 : node5566;
											assign node5566 = (inp[4]) ? node5570 : node5567;
												assign node5567 = (inp[3]) ? 11'b00011000000 : 11'b00111010000;
												assign node5570 = (inp[3]) ? 11'b00111010010 : 11'b00101010010;
											assign node5573 = (inp[4]) ? node5575 : 11'b00101010000;
												assign node5575 = (inp[3]) ? 11'b00111000000 : 11'b00111000100;
										assign node5578 = (inp[4]) ? node5586 : node5579;
											assign node5579 = (inp[9]) ? node5583 : node5580;
												assign node5580 = (inp[3]) ? 11'b00111000000 : 11'b00101010100;
												assign node5583 = (inp[3]) ? 11'b00011000010 : 11'b00111000010;
											assign node5586 = (inp[3]) ? 11'b00001000010 : 11'b00001000000;
							assign node5589 = (inp[4]) ? node5635 : node5590;
								assign node5590 = (inp[11]) ? node5610 : node5591;
									assign node5591 = (inp[9]) ? node5603 : node5592;
										assign node5592 = (inp[0]) ? node5598 : node5593;
											assign node5593 = (inp[3]) ? 11'b00110010110 : node5594;
												assign node5594 = (inp[10]) ? 11'b10101010000 : 11'b00011010000;
											assign node5598 = (inp[10]) ? 11'b00001000100 : node5599;
												assign node5599 = (inp[3]) ? 11'b00101000000 : 11'b00111000000;
										assign node5603 = (inp[10]) ? 11'b00010000010 : node5604;
											assign node5604 = (inp[3]) ? node5606 : 11'b00010010010;
												assign node5606 = (inp[0]) ? 11'b00100010010 : 11'b10000010110;
									assign node5610 = (inp[10]) ? node5622 : node5611;
										assign node5611 = (inp[0]) ? node5615 : node5612;
											assign node5612 = (inp[3]) ? 11'b10010000010 : 11'b00000000010;
											assign node5615 = (inp[9]) ? node5619 : node5616;
												assign node5616 = (inp[3]) ? 11'b00110000010 : 11'b00110010010;
												assign node5619 = (inp[3]) ? 11'b00010010010 : 11'b00010010110;
										assign node5622 = (inp[3]) ? node5628 : node5623;
											assign node5623 = (inp[0]) ? node5625 : 11'b10010010010;
												assign node5625 = (inp[9]) ? 11'b00000000010 : 11'b00100010110;
											assign node5628 = (inp[0]) ? node5632 : node5629;
												assign node5629 = (inp[9]) ? 11'b00100000110 : 11'b00000000110;
												assign node5632 = (inp[9]) ? 11'b00000000010 : 11'b00100000010;
								assign node5635 = (inp[0]) ? node5659 : node5636;
									assign node5636 = (inp[9]) ? node5650 : node5637;
										assign node5637 = (inp[10]) ? node5643 : node5638;
											assign node5638 = (inp[11]) ? 11'b00110010100 : node5639;
												assign node5639 = (inp[3]) ? 11'b10000010110 : 11'b00100010110;
											assign node5643 = (inp[3]) ? node5647 : node5644;
												assign node5644 = (inp[11]) ? 11'b10100000100 : 11'b10010000100;
												assign node5647 = (inp[11]) ? 11'b00100000000 : 11'b00010010000;
										assign node5650 = (inp[3]) ? node5656 : node5651;
											assign node5651 = (inp[10]) ? node5653 : 11'b00100010100;
												assign node5653 = (inp[11]) ? 11'b10100000000 : 11'b10110010000;
											assign node5656 = (inp[10]) ? 11'b00100000000 : 11'b10110000000;
									assign node5659 = (inp[10]) ? node5671 : node5660;
										assign node5660 = (inp[9]) ? node5666 : node5661;
											assign node5661 = (inp[11]) ? 11'b00010010000 : node5662;
												assign node5662 = (inp[3]) ? 11'b00110010000 : 11'b00000000010;
											assign node5666 = (inp[3]) ? 11'b00010000000 : node5667;
												assign node5667 = (inp[11]) ? 11'b00010000100 : 11'b00000010100;
										assign node5671 = (inp[3]) ? node5677 : node5672;
											assign node5672 = (inp[11]) ? node5674 : 11'b00010010000;
												assign node5674 = (inp[9]) ? 11'b00000000000 : 11'b00000000100;
											assign node5677 = (inp[11]) ? 11'b00000000000 : node5678;
												assign node5678 = (inp[9]) ? 11'b00000000000 : 11'b00100000000;
					assign node5682 = (inp[8]) ? node5856 : node5683;
						assign node5683 = (inp[5]) ? node5769 : node5684;
							assign node5684 = (inp[4]) ? node5724 : node5685;
								assign node5685 = (inp[0]) ? node5699 : node5686;
									assign node5686 = (inp[10]) ? node5694 : node5687;
										assign node5687 = (inp[3]) ? node5691 : node5688;
											assign node5688 = (inp[11]) ? 11'b00101000000 : 11'b00111000010;
											assign node5691 = (inp[11]) ? 11'b10111010010 : 11'b10111000010;
										assign node5694 = (inp[9]) ? 11'b00111010110 : node5695;
											assign node5695 = (inp[11]) ? 11'b00101010110 : 11'b00101000110;
									assign node5699 = (inp[3]) ? node5713 : node5700;
										assign node5700 = (inp[11]) ? node5708 : node5701;
											assign node5701 = (inp[10]) ? node5705 : node5702;
												assign node5702 = (inp[9]) ? 11'b00011000110 : 11'b00011000010;
												assign node5705 = (inp[9]) ? 11'b00001010010 : 11'b00001000110;
											assign node5708 = (inp[9]) ? 11'b00101010110 : node5709;
												assign node5709 = (inp[10]) ? 11'b00011010110 : 11'b00001010000;
										assign node5713 = (inp[10]) ? node5719 : node5714;
											assign node5714 = (inp[9]) ? node5716 : 11'b00011000010;
												assign node5716 = (inp[11]) ? 11'b00111010010 : 11'b00011010010;
											assign node5719 = (inp[11]) ? node5721 : 11'b00001000010;
												assign node5721 = (inp[9]) ? 11'b00011000010 : 11'b00101000010;
								assign node5724 = (inp[10]) ? node5750 : node5725;
									assign node5725 = (inp[11]) ? node5737 : node5726;
										assign node5726 = (inp[0]) ? node5732 : node5727;
											assign node5727 = (inp[9]) ? 11'b10011010000 : node5728;
												assign node5728 = (inp[3]) ? 11'b10111000100 : 11'b00111000100;
											assign node5732 = (inp[9]) ? 11'b00111000000 : node5733;
												assign node5733 = (inp[3]) ? 11'b00011010000 : 11'b00011000000;
										assign node5737 = (inp[9]) ? node5745 : node5738;
											assign node5738 = (inp[0]) ? node5742 : node5739;
												assign node5739 = (inp[3]) ? 11'b10001000110 : 11'b00101000110;
												assign node5742 = (inp[3]) ? 11'b00101010010 : 11'b00001010010;
											assign node5745 = (inp[3]) ? 11'b10101010000 : node5746;
												assign node5746 = (inp[0]) ? 11'b00011000100 : 11'b00111010100;
									assign node5750 = (inp[3]) ? node5760 : node5751;
										assign node5751 = (inp[0]) ? node5755 : node5752;
											assign node5752 = (inp[11]) ? 11'b10001010000 : 11'b10101010100;
											assign node5755 = (inp[9]) ? node5757 : 11'b00001010100;
												assign node5757 = (inp[11]) ? 11'b00101000000 : 11'b00101010000;
										assign node5760 = (inp[0]) ? node5766 : node5761;
											assign node5761 = (inp[11]) ? 11'b00011010000 : node5762;
												assign node5762 = (inp[9]) ? 11'b00001010000 : 11'b00001000000;
											assign node5766 = (inp[9]) ? 11'b00001000000 : 11'b00011000000;
							assign node5769 = (inp[11]) ? node5819 : node5770;
								assign node5770 = (inp[4]) ? node5798 : node5771;
									assign node5771 = (inp[9]) ? node5783 : node5772;
										assign node5772 = (inp[0]) ? node5778 : node5773;
											assign node5773 = (inp[3]) ? 11'b00001010100 : node5774;
												assign node5774 = (inp[10]) ? 11'b10011010000 : 11'b00111010000;
											assign node5778 = (inp[3]) ? node5780 : 11'b00101000100;
												assign node5780 = (inp[10]) ? 11'b00001000000 : 11'b00111000000;
										assign node5783 = (inp[10]) ? node5791 : node5784;
											assign node5784 = (inp[3]) ? node5788 : node5785;
												assign node5785 = (inp[0]) ? 11'b00001000100 : 11'b00101010000;
												assign node5788 = (inp[0]) ? 11'b00110010010 : 11'b10110010110;
											assign node5791 = (inp[0]) ? node5795 : node5792;
												assign node5792 = (inp[3]) ? 11'b00110000110 : 11'b10010000110;
												assign node5795 = (inp[3]) ? 11'b00010000010 : 11'b00110010010;
									assign node5798 = (inp[0]) ? node5810 : node5799;
										assign node5799 = (inp[10]) ? node5805 : node5800;
											assign node5800 = (inp[3]) ? node5802 : 11'b00010010110;
												assign node5802 = (inp[9]) ? 11'b10110000010 : 11'b10000010110;
											assign node5805 = (inp[3]) ? 11'b00110010010 : node5806;
												assign node5806 = (inp[9]) ? 11'b10100010010 : 11'b10100000110;
										assign node5810 = (inp[9]) ? node5816 : node5811;
											assign node5811 = (inp[10]) ? 11'b00110000010 : node5812;
												assign node5812 = (inp[3]) ? 11'b00100010010 : 11'b00100000010;
											assign node5816 = (inp[10]) ? 11'b00000000010 : 11'b00010000010;
								assign node5819 = (inp[9]) ? node5841 : node5820;
									assign node5820 = (inp[3]) ? node5832 : node5821;
										assign node5821 = (inp[10]) ? node5829 : node5822;
											assign node5822 = (inp[4]) ? node5826 : node5823;
												assign node5823 = (inp[0]) ? 11'b00000010010 : 11'b00100010010;
												assign node5826 = (inp[0]) ? 11'b00110010000 : 11'b00110010100;
											assign node5829 = (inp[0]) ? 11'b00010010100 : 11'b10010010000;
										assign node5832 = (inp[0]) ? node5836 : node5833;
											assign node5833 = (inp[10]) ? 11'b00110000100 : 11'b10000000010;
											assign node5836 = (inp[4]) ? node5838 : 11'b00110000000;
												assign node5838 = (inp[10]) ? 11'b00010000000 : 11'b00010010000;
									assign node5841 = (inp[4]) ? node5849 : node5842;
										assign node5842 = (inp[10]) ? 11'b00100000100 : node5843;
											assign node5843 = (inp[0]) ? node5845 : 11'b10100010100;
												assign node5845 = (inp[3]) ? 11'b00000010000 : 11'b00100010100;
										assign node5849 = (inp[3]) ? 11'b00000000000 : node5850;
											assign node5850 = (inp[10]) ? node5852 : 11'b00100000100;
												assign node5852 = (inp[0]) ? 11'b00100000000 : 11'b10100000000;
						assign node5856 = (inp[5]) ? node5944 : node5857;
							assign node5857 = (inp[11]) ? node5901 : node5858;
								assign node5858 = (inp[9]) ? node5874 : node5859;
									assign node5859 = (inp[4]) ? node5867 : node5860;
										assign node5860 = (inp[3]) ? node5864 : node5861;
											assign node5861 = (inp[0]) ? 11'b00110000110 : 11'b00110000010;
											assign node5864 = (inp[10]) ? 11'b00010000010 : 11'b10010000010;
										assign node5867 = (inp[0]) ? 11'b00010010010 : node5868;
											assign node5868 = (inp[3]) ? 11'b10110000110 : node5869;
												assign node5869 = (inp[10]) ? 11'b10010010110 : 11'b00000000110;
									assign node5874 = (inp[0]) ? node5890 : node5875;
										assign node5875 = (inp[3]) ? node5883 : node5876;
											assign node5876 = (inp[10]) ? node5880 : node5877;
												assign node5877 = (inp[4]) ? 11'b00010000110 : 11'b00100000010;
												assign node5880 = (inp[4]) ? 11'b10100000010 : 11'b10100010110;
											assign node5883 = (inp[4]) ? node5887 : node5884;
												assign node5884 = (inp[10]) ? 11'b00000010110 : 11'b10000000110;
												assign node5887 = (inp[10]) ? 11'b00000010010 : 11'b10100010010;
										assign node5890 = (inp[3]) ? node5896 : node5891;
											assign node5891 = (inp[10]) ? node5893 : 11'b00010010110;
												assign node5893 = (inp[4]) ? 11'b00000010010 : 11'b00100010010;
											assign node5896 = (inp[4]) ? node5898 : 11'b00000010010;
												assign node5898 = (inp[10]) ? 11'b00000000010 : 11'b00100000010;
								assign node5901 = (inp[4]) ? node5925 : node5902;
									assign node5902 = (inp[10]) ? node5914 : node5903;
										assign node5903 = (inp[9]) ? node5909 : node5904;
											assign node5904 = (inp[3]) ? node5906 : 11'b00100000010;
												assign node5906 = (inp[0]) ? 11'b00000000010 : 11'b10000010010;
											assign node5909 = (inp[3]) ? 11'b00110010000 : node5910;
												assign node5910 = (inp[0]) ? 11'b00010010100 : 11'b00010010000;
										assign node5914 = (inp[0]) ? node5920 : node5915;
											assign node5915 = (inp[3]) ? node5917 : 11'b10110010100;
												assign node5917 = (inp[9]) ? 11'b00010010100 : 11'b00110010100;
											assign node5920 = (inp[9]) ? 11'b00110000000 : node5921;
												assign node5921 = (inp[3]) ? 11'b00110000000 : 11'b00110010100;
									assign node5925 = (inp[0]) ? node5937 : node5926;
										assign node5926 = (inp[9]) ? node5932 : node5927;
											assign node5927 = (inp[10]) ? 11'b10000010100 : node5928;
												assign node5928 = (inp[3]) ? 11'b10100000100 : 11'b00010000100;
											assign node5932 = (inp[10]) ? 11'b10000010000 : node5933;
												assign node5933 = (inp[3]) ? 11'b10100010000 : 11'b00100010100;
										assign node5937 = (inp[10]) ? 11'b00000000000 : node5938;
											assign node5938 = (inp[3]) ? node5940 : 11'b00100000100;
												assign node5940 = (inp[9]) ? 11'b00100000000 : 11'b00100010000;
							assign node5944 = (inp[11]) ? node5986 : node5945;
								assign node5945 = (inp[4]) ? node5965 : node5946;
									assign node5946 = (inp[0]) ? node5954 : node5947;
										assign node5947 = (inp[9]) ? 11'b10110000100 : node5948;
											assign node5948 = (inp[10]) ? 11'b10010010000 : node5949;
												assign node5949 = (inp[3]) ? 11'b10110010000 : 11'b00110010000;
										assign node5954 = (inp[10]) ? node5960 : node5955;
											assign node5955 = (inp[3]) ? node5957 : 11'b00110000100;
												assign node5957 = (inp[9]) ? 11'b00110010000 : 11'b00110000000;
											assign node5960 = (inp[9]) ? 11'b00010010000 : node5961;
												assign node5961 = (inp[3]) ? 11'b00010000000 : 11'b00010000100;
									assign node5965 = (inp[9]) ? node5979 : node5966;
										assign node5966 = (inp[3]) ? node5974 : node5967;
											assign node5967 = (inp[10]) ? node5971 : node5968;
												assign node5968 = (inp[0]) ? 11'b00010000000 : 11'b00010010100;
												assign node5971 = (inp[0]) ? 11'b00100010100 : 11'b10100000100;
											assign node5974 = (inp[10]) ? node5976 : 11'b00100010000;
												assign node5976 = (inp[0]) ? 11'b00100000000 : 11'b00100010000;
										assign node5979 = (inp[0]) ? node5983 : node5980;
											assign node5980 = (inp[10]) ? 11'b10000010000 : 11'b10000000000;
											assign node5983 = (inp[3]) ? 11'b00000000000 : 11'b00000010000;
								assign node5986 = (inp[4]) ? node6008 : node5987;
									assign node5987 = (inp[9]) ? node5997 : node5988;
										assign node5988 = (inp[10]) ? node5994 : node5989;
											assign node5989 = (inp[3]) ? node5991 : 11'b00100010000;
												assign node5991 = (inp[0]) ? 11'b00100000000 : 11'b10100000000;
											assign node5994 = (inp[0]) ? 11'b00100010100 : 11'b00100000100;
										assign node5997 = (inp[0]) ? node6003 : node5998;
											assign node5998 = (inp[3]) ? 11'b10000010100 : node5999;
												assign node5999 = (inp[10]) ? 11'b10000000100 : 11'b00100000000;
											assign node6003 = (inp[10]) ? 11'b00000000000 : node6004;
												assign node6004 = (inp[3]) ? 11'b00000010000 : 11'b00000010100;
									assign node6008 = (inp[3]) ? node6022 : node6009;
										assign node6009 = (inp[10]) ? node6015 : node6010;
											assign node6010 = (inp[9]) ? 11'b00000000100 : node6011;
												assign node6011 = (inp[0]) ? 11'b00000010000 : 11'b00000010100;
											assign node6015 = (inp[9]) ? node6019 : node6016;
												assign node6016 = (inp[0]) ? 11'b00000000100 : 11'b10000000100;
												assign node6019 = (inp[0]) ? 11'b00000000000 : 11'b10000000000;
										assign node6022 = (inp[10]) ? 11'b00000000000 : node6023;
											assign node6023 = (inp[9]) ? 11'b00000000000 : 11'b00000010000;

endmodule