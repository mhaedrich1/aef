module dtc_split66_bm21 (
	input  wire [10-1:0] inp,
	output wire [10-1:0] outp
);

	wire [10-1:0] node1;
	wire [10-1:0] node2;
	wire [10-1:0] node3;
	wire [10-1:0] node4;
	wire [10-1:0] node5;
	wire [10-1:0] node8;
	wire [10-1:0] node11;
	wire [10-1:0] node12;
	wire [10-1:0] node15;
	wire [10-1:0] node18;
	wire [10-1:0] node19;
	wire [10-1:0] node20;
	wire [10-1:0] node23;
	wire [10-1:0] node26;
	wire [10-1:0] node27;
	wire [10-1:0] node30;
	wire [10-1:0] node33;
	wire [10-1:0] node34;
	wire [10-1:0] node35;
	wire [10-1:0] node36;
	wire [10-1:0] node39;
	wire [10-1:0] node42;
	wire [10-1:0] node43;
	wire [10-1:0] node46;
	wire [10-1:0] node49;
	wire [10-1:0] node50;
	wire [10-1:0] node51;
	wire [10-1:0] node54;
	wire [10-1:0] node57;
	wire [10-1:0] node58;
	wire [10-1:0] node61;
	wire [10-1:0] node64;
	wire [10-1:0] node65;
	wire [10-1:0] node66;
	wire [10-1:0] node67;
	wire [10-1:0] node68;
	wire [10-1:0] node71;
	wire [10-1:0] node74;
	wire [10-1:0] node75;
	wire [10-1:0] node78;
	wire [10-1:0] node81;
	wire [10-1:0] node82;
	wire [10-1:0] node83;
	wire [10-1:0] node86;
	wire [10-1:0] node89;
	wire [10-1:0] node90;
	wire [10-1:0] node93;
	wire [10-1:0] node96;
	wire [10-1:0] node97;
	wire [10-1:0] node98;
	wire [10-1:0] node99;
	wire [10-1:0] node102;
	wire [10-1:0] node105;
	wire [10-1:0] node106;
	wire [10-1:0] node109;
	wire [10-1:0] node112;
	wire [10-1:0] node113;
	wire [10-1:0] node114;
	wire [10-1:0] node117;
	wire [10-1:0] node120;
	wire [10-1:0] node121;
	wire [10-1:0] node124;

	assign outp = (inp[2]) ? node64 : node1;
		assign node1 = (inp[9]) ? node33 : node2;
			assign node2 = (inp[8]) ? node18 : node3;
				assign node3 = (inp[5]) ? node11 : node4;
					assign node4 = (inp[7]) ? node8 : node5;
						assign node5 = (inp[4]) ? 10'b0001111111 : 10'b0011111111;
						assign node8 = (inp[1]) ? 10'b0000111111 : 10'b0001111111;
					assign node11 = (inp[3]) ? node15 : node12;
						assign node12 = (inp[4]) ? 10'b0000111111 : 10'b0001111111;
						assign node15 = (inp[1]) ? 10'b0000011111 : 10'b0000111111;
				assign node18 = (inp[4]) ? node26 : node19;
					assign node19 = (inp[5]) ? node23 : node20;
						assign node20 = (inp[3]) ? 10'b0000111111 : 10'b0001111111;
						assign node23 = (inp[7]) ? 10'b0000011111 : 10'b0000111111;
					assign node26 = (inp[7]) ? node30 : node27;
						assign node27 = (inp[5]) ? 10'b0000011111 : 10'b0000111111;
						assign node30 = (inp[1]) ? 10'b0000001111 : 10'b0000011111;
			assign node33 = (inp[0]) ? node49 : node34;
				assign node34 = (inp[1]) ? node42 : node35;
					assign node35 = (inp[7]) ? node39 : node36;
						assign node36 = (inp[6]) ? 10'b0000111111 : 10'b0001111111;
						assign node39 = (inp[6]) ? 10'b0000011111 : 10'b0000111111;
					assign node42 = (inp[8]) ? node46 : node43;
						assign node43 = (inp[5]) ? 10'b0000011111 : 10'b0000111111;
						assign node46 = (inp[7]) ? 10'b0000001111 : 10'b0000011111;
				assign node49 = (inp[7]) ? node57 : node50;
					assign node50 = (inp[3]) ? node54 : node51;
						assign node51 = (inp[1]) ? 10'b0000011111 : 10'b0000111111;
						assign node54 = (inp[8]) ? 10'b0000001111 : 10'b0000011111;
					assign node57 = (inp[8]) ? node61 : node58;
						assign node58 = (inp[6]) ? 10'b0000001111 : 10'b0000011111;
						assign node61 = (inp[5]) ? 10'b0000000111 : 10'b0000001111;
		assign node64 = (inp[8]) ? node96 : node65;
			assign node65 = (inp[6]) ? node81 : node66;
				assign node66 = (inp[0]) ? node74 : node67;
					assign node67 = (inp[4]) ? node71 : node68;
						assign node68 = (inp[3]) ? 10'b0000111111 : 10'b0001111111;
						assign node71 = (inp[9]) ? 10'b0000011111 : 10'b0000111111;
					assign node74 = (inp[1]) ? node78 : node75;
						assign node75 = (inp[5]) ? 10'b0000011111 : 10'b0000111111;
						assign node78 = (inp[5]) ? 10'b0000001111 : 10'b0000011111;
				assign node81 = (inp[9]) ? node89 : node82;
					assign node82 = (inp[7]) ? node86 : node83;
						assign node83 = (inp[3]) ? 10'b0000011111 : 10'b0000111111;
						assign node86 = (inp[5]) ? 10'b0000001111 : 10'b0000011111;
					assign node89 = (inp[3]) ? node93 : node90;
						assign node90 = (inp[4]) ? 10'b0000001111 : 10'b0000011111;
						assign node93 = (inp[5]) ? 10'b0000000111 : 10'b0000001111;
			assign node96 = (inp[1]) ? node112 : node97;
				assign node97 = (inp[7]) ? node105 : node98;
					assign node98 = (inp[4]) ? node102 : node99;
						assign node99 = (inp[9]) ? 10'b0000011111 : 10'b0000111111;
						assign node102 = (inp[9]) ? 10'b0000001111 : 10'b0000011111;
					assign node105 = (inp[6]) ? node109 : node106;
						assign node106 = (inp[9]) ? 10'b0000001111 : 10'b0000011111;
						assign node109 = (inp[0]) ? 10'b0000000111 : 10'b0000001111;
				assign node112 = (inp[5]) ? node120 : node113;
					assign node113 = (inp[7]) ? node117 : node114;
						assign node114 = (inp[4]) ? 10'b0000001111 : 10'b0000011111;
						assign node117 = (inp[6]) ? 10'b0000000111 : 10'b0000001111;
					assign node120 = (inp[7]) ? node124 : node121;
						assign node121 = (inp[9]) ? 10'b0000000111 : 10'b0000001111;
						assign node124 = (inp[0]) ? 10'b0000000011 : 10'b0000000111;

endmodule