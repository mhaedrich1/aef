module dtc_split05_bm65 (
	input  wire [16-1:0] inp,
	output wire [4-1:0] outp
);

	wire [4-1:0] node1;
	wire [4-1:0] node2;
	wire [4-1:0] node3;
	wire [4-1:0] node4;
	wire [4-1:0] node5;
	wire [4-1:0] node6;
	wire [4-1:0] node7;
	wire [4-1:0] node8;
	wire [4-1:0] node9;
	wire [4-1:0] node10;
	wire [4-1:0] node14;
	wire [4-1:0] node16;
	wire [4-1:0] node18;
	wire [4-1:0] node21;
	wire [4-1:0] node22;
	wire [4-1:0] node23;
	wire [4-1:0] node25;
	wire [4-1:0] node28;
	wire [4-1:0] node29;
	wire [4-1:0] node33;
	wire [4-1:0] node34;
	wire [4-1:0] node36;
	wire [4-1:0] node39;
	wire [4-1:0] node42;
	wire [4-1:0] node43;
	wire [4-1:0] node44;
	wire [4-1:0] node45;
	wire [4-1:0] node48;
	wire [4-1:0] node49;
	wire [4-1:0] node53;
	wire [4-1:0] node54;
	wire [4-1:0] node57;
	wire [4-1:0] node58;
	wire [4-1:0] node62;
	wire [4-1:0] node63;
	wire [4-1:0] node66;
	wire [4-1:0] node67;
	wire [4-1:0] node69;
	wire [4-1:0] node73;
	wire [4-1:0] node75;
	wire [4-1:0] node76;
	wire [4-1:0] node77;
	wire [4-1:0] node80;
	wire [4-1:0] node81;
	wire [4-1:0] node85;
	wire [4-1:0] node86;
	wire [4-1:0] node88;
	wire [4-1:0] node91;
	wire [4-1:0] node95;
	wire [4-1:0] node96;
	wire [4-1:0] node97;
	wire [4-1:0] node98;
	wire [4-1:0] node99;
	wire [4-1:0] node100;
	wire [4-1:0] node101;
	wire [4-1:0] node103;
	wire [4-1:0] node106;
	wire [4-1:0] node107;
	wire [4-1:0] node111;
	wire [4-1:0] node112;
	wire [4-1:0] node113;
	wire [4-1:0] node117;
	wire [4-1:0] node120;
	wire [4-1:0] node121;
	wire [4-1:0] node123;
	wire [4-1:0] node126;
	wire [4-1:0] node127;
	wire [4-1:0] node128;
	wire [4-1:0] node132;
	wire [4-1:0] node133;
	wire [4-1:0] node136;
	wire [4-1:0] node139;
	wire [4-1:0] node140;
	wire [4-1:0] node141;
	wire [4-1:0] node143;
	wire [4-1:0] node145;
	wire [4-1:0] node148;
	wire [4-1:0] node149;
	wire [4-1:0] node153;
	wire [4-1:0] node154;
	wire [4-1:0] node156;
	wire [4-1:0] node157;
	wire [4-1:0] node161;
	wire [4-1:0] node162;
	wire [4-1:0] node163;
	wire [4-1:0] node166;
	wire [4-1:0] node170;
	wire [4-1:0] node171;
	wire [4-1:0] node172;
	wire [4-1:0] node173;
	wire [4-1:0] node175;
	wire [4-1:0] node177;
	wire [4-1:0] node180;
	wire [4-1:0] node182;
	wire [4-1:0] node185;
	wire [4-1:0] node186;
	wire [4-1:0] node187;
	wire [4-1:0] node188;
	wire [4-1:0] node192;
	wire [4-1:0] node193;
	wire [4-1:0] node197;
	wire [4-1:0] node198;
	wire [4-1:0] node200;
	wire [4-1:0] node205;
	wire [4-1:0] node206;
	wire [4-1:0] node207;
	wire [4-1:0] node208;
	wire [4-1:0] node209;
	wire [4-1:0] node210;
	wire [4-1:0] node214;
	wire [4-1:0] node215;
	wire [4-1:0] node217;
	wire [4-1:0] node220;
	wire [4-1:0] node223;
	wire [4-1:0] node224;
	wire [4-1:0] node225;
	wire [4-1:0] node227;
	wire [4-1:0] node231;
	wire [4-1:0] node232;
	wire [4-1:0] node234;
	wire [4-1:0] node238;
	wire [4-1:0] node239;
	wire [4-1:0] node240;
	wire [4-1:0] node242;
	wire [4-1:0] node245;
	wire [4-1:0] node247;
	wire [4-1:0] node250;
	wire [4-1:0] node251;
	wire [4-1:0] node253;
	wire [4-1:0] node256;
	wire [4-1:0] node259;
	wire [4-1:0] node260;
	wire [4-1:0] node261;
	wire [4-1:0] node262;
	wire [4-1:0] node263;
	wire [4-1:0] node264;
	wire [4-1:0] node268;
	wire [4-1:0] node269;
	wire [4-1:0] node273;
	wire [4-1:0] node274;
	wire [4-1:0] node277;
	wire [4-1:0] node279;
	wire [4-1:0] node282;
	wire [4-1:0] node283;
	wire [4-1:0] node285;
	wire [4-1:0] node288;
	wire [4-1:0] node289;
	wire [4-1:0] node290;
	wire [4-1:0] node295;
	wire [4-1:0] node296;
	wire [4-1:0] node297;
	wire [4-1:0] node298;
	wire [4-1:0] node301;
	wire [4-1:0] node303;
	wire [4-1:0] node306;
	wire [4-1:0] node307;
	wire [4-1:0] node311;
	wire [4-1:0] node312;
	wire [4-1:0] node314;
	wire [4-1:0] node317;
	wire [4-1:0] node318;
	wire [4-1:0] node322;
	wire [4-1:0] node323;
	wire [4-1:0] node324;
	wire [4-1:0] node325;
	wire [4-1:0] node326;
	wire [4-1:0] node328;
	wire [4-1:0] node329;
	wire [4-1:0] node330;
	wire [4-1:0] node333;
	wire [4-1:0] node336;
	wire [4-1:0] node337;
	wire [4-1:0] node340;
	wire [4-1:0] node342;
	wire [4-1:0] node345;
	wire [4-1:0] node346;
	wire [4-1:0] node347;
	wire [4-1:0] node348;
	wire [4-1:0] node350;
	wire [4-1:0] node353;
	wire [4-1:0] node355;
	wire [4-1:0] node358;
	wire [4-1:0] node360;
	wire [4-1:0] node361;
	wire [4-1:0] node364;
	wire [4-1:0] node367;
	wire [4-1:0] node368;
	wire [4-1:0] node369;
	wire [4-1:0] node372;
	wire [4-1:0] node375;
	wire [4-1:0] node376;
	wire [4-1:0] node378;
	wire [4-1:0] node381;
	wire [4-1:0] node383;
	wire [4-1:0] node386;
	wire [4-1:0] node388;
	wire [4-1:0] node390;
	wire [4-1:0] node391;
	wire [4-1:0] node392;
	wire [4-1:0] node393;
	wire [4-1:0] node396;
	wire [4-1:0] node400;
	wire [4-1:0] node401;
	wire [4-1:0] node402;
	wire [4-1:0] node406;
	wire [4-1:0] node410;
	wire [4-1:0] node411;
	wire [4-1:0] node412;
	wire [4-1:0] node413;
	wire [4-1:0] node414;
	wire [4-1:0] node415;
	wire [4-1:0] node416;
	wire [4-1:0] node417;
	wire [4-1:0] node420;
	wire [4-1:0] node424;
	wire [4-1:0] node425;
	wire [4-1:0] node426;
	wire [4-1:0] node430;
	wire [4-1:0] node433;
	wire [4-1:0] node434;
	wire [4-1:0] node436;
	wire [4-1:0] node439;
	wire [4-1:0] node440;
	wire [4-1:0] node442;
	wire [4-1:0] node445;
	wire [4-1:0] node448;
	wire [4-1:0] node449;
	wire [4-1:0] node450;
	wire [4-1:0] node452;
	wire [4-1:0] node454;
	wire [4-1:0] node457;
	wire [4-1:0] node459;
	wire [4-1:0] node462;
	wire [4-1:0] node463;
	wire [4-1:0] node465;
	wire [4-1:0] node468;
	wire [4-1:0] node470;
	wire [4-1:0] node473;
	wire [4-1:0] node474;
	wire [4-1:0] node475;
	wire [4-1:0] node476;
	wire [4-1:0] node479;
	wire [4-1:0] node480;
	wire [4-1:0] node482;
	wire [4-1:0] node485;
	wire [4-1:0] node487;
	wire [4-1:0] node490;
	wire [4-1:0] node491;
	wire [4-1:0] node492;
	wire [4-1:0] node493;
	wire [4-1:0] node497;
	wire [4-1:0] node499;
	wire [4-1:0] node502;
	wire [4-1:0] node503;
	wire [4-1:0] node504;
	wire [4-1:0] node508;
	wire [4-1:0] node511;
	wire [4-1:0] node512;
	wire [4-1:0] node513;
	wire [4-1:0] node514;
	wire [4-1:0] node515;
	wire [4-1:0] node518;
	wire [4-1:0] node521;
	wire [4-1:0] node524;
	wire [4-1:0] node525;
	wire [4-1:0] node526;
	wire [4-1:0] node530;
	wire [4-1:0] node531;
	wire [4-1:0] node534;
	wire [4-1:0] node537;
	wire [4-1:0] node538;
	wire [4-1:0] node539;
	wire [4-1:0] node543;
	wire [4-1:0] node545;
	wire [4-1:0] node548;
	wire [4-1:0] node549;
	wire [4-1:0] node551;
	wire [4-1:0] node552;
	wire [4-1:0] node553;
	wire [4-1:0] node557;
	wire [4-1:0] node558;
	wire [4-1:0] node559;
	wire [4-1:0] node561;
	wire [4-1:0] node564;
	wire [4-1:0] node565;
	wire [4-1:0] node568;
	wire [4-1:0] node572;
	wire [4-1:0] node573;
	wire [4-1:0] node574;
	wire [4-1:0] node575;
	wire [4-1:0] node576;
	wire [4-1:0] node577;
	wire [4-1:0] node580;
	wire [4-1:0] node583;
	wire [4-1:0] node585;
	wire [4-1:0] node589;
	wire [4-1:0] node590;
	wire [4-1:0] node591;
	wire [4-1:0] node593;
	wire [4-1:0] node596;
	wire [4-1:0] node599;
	wire [4-1:0] node600;
	wire [4-1:0] node601;
	wire [4-1:0] node606;
	wire [4-1:0] node608;
	wire [4-1:0] node609;
	wire [4-1:0] node610;
	wire [4-1:0] node612;
	wire [4-1:0] node616;
	wire [4-1:0] node618;
	wire [4-1:0] node619;
	wire [4-1:0] node623;
	wire [4-1:0] node624;
	wire [4-1:0] node625;
	wire [4-1:0] node626;
	wire [4-1:0] node627;
	wire [4-1:0] node628;
	wire [4-1:0] node629;
	wire [4-1:0] node630;
	wire [4-1:0] node631;
	wire [4-1:0] node635;
	wire [4-1:0] node638;
	wire [4-1:0] node639;
	wire [4-1:0] node640;
	wire [4-1:0] node644;
	wire [4-1:0] node645;
	wire [4-1:0] node646;
	wire [4-1:0] node650;
	wire [4-1:0] node654;
	wire [4-1:0] node655;
	wire [4-1:0] node656;
	wire [4-1:0] node657;
	wire [4-1:0] node658;
	wire [4-1:0] node663;
	wire [4-1:0] node664;
	wire [4-1:0] node666;
	wire [4-1:0] node669;
	wire [4-1:0] node670;
	wire [4-1:0] node672;
	wire [4-1:0] node675;
	wire [4-1:0] node676;
	wire [4-1:0] node680;
	wire [4-1:0] node681;
	wire [4-1:0] node682;
	wire [4-1:0] node683;
	wire [4-1:0] node684;
	wire [4-1:0] node688;
	wire [4-1:0] node689;
	wire [4-1:0] node693;
	wire [4-1:0] node694;
	wire [4-1:0] node697;
	wire [4-1:0] node698;
	wire [4-1:0] node701;
	wire [4-1:0] node704;
	wire [4-1:0] node705;
	wire [4-1:0] node706;
	wire [4-1:0] node709;
	wire [4-1:0] node712;
	wire [4-1:0] node713;
	wire [4-1:0] node716;
	wire [4-1:0] node720;
	wire [4-1:0] node721;
	wire [4-1:0] node722;
	wire [4-1:0] node723;
	wire [4-1:0] node724;
	wire [4-1:0] node725;
	wire [4-1:0] node727;
	wire [4-1:0] node729;
	wire [4-1:0] node732;
	wire [4-1:0] node733;
	wire [4-1:0] node736;
	wire [4-1:0] node737;
	wire [4-1:0] node741;
	wire [4-1:0] node742;
	wire [4-1:0] node743;
	wire [4-1:0] node747;
	wire [4-1:0] node748;
	wire [4-1:0] node750;
	wire [4-1:0] node753;
	wire [4-1:0] node756;
	wire [4-1:0] node757;
	wire [4-1:0] node758;
	wire [4-1:0] node759;
	wire [4-1:0] node760;
	wire [4-1:0] node765;
	wire [4-1:0] node766;
	wire [4-1:0] node770;
	wire [4-1:0] node771;
	wire [4-1:0] node772;
	wire [4-1:0] node775;
	wire [4-1:0] node777;
	wire [4-1:0] node780;
	wire [4-1:0] node781;
	wire [4-1:0] node784;
	wire [4-1:0] node787;
	wire [4-1:0] node788;
	wire [4-1:0] node789;
	wire [4-1:0] node790;
	wire [4-1:0] node791;
	wire [4-1:0] node795;
	wire [4-1:0] node797;
	wire [4-1:0] node798;
	wire [4-1:0] node802;
	wire [4-1:0] node803;
	wire [4-1:0] node806;
	wire [4-1:0] node810;
	wire [4-1:0] node811;
	wire [4-1:0] node812;
	wire [4-1:0] node813;
	wire [4-1:0] node814;
	wire [4-1:0] node816;
	wire [4-1:0] node819;
	wire [4-1:0] node820;
	wire [4-1:0] node822;
	wire [4-1:0] node826;
	wire [4-1:0] node827;
	wire [4-1:0] node828;
	wire [4-1:0] node830;
	wire [4-1:0] node834;
	wire [4-1:0] node836;
	wire [4-1:0] node839;
	wire [4-1:0] node840;
	wire [4-1:0] node841;
	wire [4-1:0] node842;
	wire [4-1:0] node843;
	wire [4-1:0] node846;
	wire [4-1:0] node849;
	wire [4-1:0] node850;
	wire [4-1:0] node853;
	wire [4-1:0] node856;
	wire [4-1:0] node857;
	wire [4-1:0] node861;
	wire [4-1:0] node862;
	wire [4-1:0] node863;
	wire [4-1:0] node865;
	wire [4-1:0] node870;
	wire [4-1:0] node871;
	wire [4-1:0] node872;
	wire [4-1:0] node873;
	wire [4-1:0] node874;
	wire [4-1:0] node875;
	wire [4-1:0] node878;
	wire [4-1:0] node881;
	wire [4-1:0] node882;
	wire [4-1:0] node887;
	wire [4-1:0] node888;
	wire [4-1:0] node889;
	wire [4-1:0] node891;
	wire [4-1:0] node894;
	wire [4-1:0] node896;
	wire [4-1:0] node899;
	wire [4-1:0] node900;
	wire [4-1:0] node901;
	wire [4-1:0] node905;
	wire [4-1:0] node908;
	wire [4-1:0] node909;
	wire [4-1:0] node910;
	wire [4-1:0] node911;
	wire [4-1:0] node912;
	wire [4-1:0] node915;
	wire [4-1:0] node918;
	wire [4-1:0] node921;
	wire [4-1:0] node922;
	wire [4-1:0] node923;
	wire [4-1:0] node927;
	wire [4-1:0] node930;
	wire [4-1:0] node931;
	wire [4-1:0] node935;
	wire [4-1:0] node936;
	wire [4-1:0] node937;
	wire [4-1:0] node938;
	wire [4-1:0] node940;
	wire [4-1:0] node942;
	wire [4-1:0] node943;
	wire [4-1:0] node944;
	wire [4-1:0] node946;
	wire [4-1:0] node949;
	wire [4-1:0] node951;
	wire [4-1:0] node955;
	wire [4-1:0] node956;
	wire [4-1:0] node957;
	wire [4-1:0] node958;
	wire [4-1:0] node959;
	wire [4-1:0] node963;
	wire [4-1:0] node966;
	wire [4-1:0] node967;
	wire [4-1:0] node970;
	wire [4-1:0] node971;
	wire [4-1:0] node973;
	wire [4-1:0] node976;
	wire [4-1:0] node977;
	wire [4-1:0] node980;
	wire [4-1:0] node983;
	wire [4-1:0] node985;
	wire [4-1:0] node986;
	wire [4-1:0] node989;
	wire [4-1:0] node991;
	wire [4-1:0] node994;
	wire [4-1:0] node995;
	wire [4-1:0] node996;
	wire [4-1:0] node997;
	wire [4-1:0] node998;
	wire [4-1:0] node999;
	wire [4-1:0] node1000;
	wire [4-1:0] node1003;
	wire [4-1:0] node1006;
	wire [4-1:0] node1009;
	wire [4-1:0] node1010;
	wire [4-1:0] node1013;
	wire [4-1:0] node1014;
	wire [4-1:0] node1018;
	wire [4-1:0] node1019;
	wire [4-1:0] node1020;
	wire [4-1:0] node1023;
	wire [4-1:0] node1026;
	wire [4-1:0] node1027;
	wire [4-1:0] node1028;
	wire [4-1:0] node1031;
	wire [4-1:0] node1035;
	wire [4-1:0] node1036;
	wire [4-1:0] node1037;
	wire [4-1:0] node1038;
	wire [4-1:0] node1041;
	wire [4-1:0] node1044;
	wire [4-1:0] node1046;
	wire [4-1:0] node1047;
	wire [4-1:0] node1051;
	wire [4-1:0] node1052;
	wire [4-1:0] node1053;
	wire [4-1:0] node1056;
	wire [4-1:0] node1057;
	wire [4-1:0] node1061;
	wire [4-1:0] node1063;
	wire [4-1:0] node1065;
	wire [4-1:0] node1068;
	wire [4-1:0] node1069;
	wire [4-1:0] node1070;
	wire [4-1:0] node1071;
	wire [4-1:0] node1074;
	wire [4-1:0] node1075;
	wire [4-1:0] node1077;
	wire [4-1:0] node1080;
	wire [4-1:0] node1083;
	wire [4-1:0] node1084;
	wire [4-1:0] node1085;
	wire [4-1:0] node1086;
	wire [4-1:0] node1091;
	wire [4-1:0] node1092;
	wire [4-1:0] node1096;
	wire [4-1:0] node1097;
	wire [4-1:0] node1098;
	wire [4-1:0] node1101;
	wire [4-1:0] node1103;
	wire [4-1:0] node1106;
	wire [4-1:0] node1107;
	wire [4-1:0] node1108;
	wire [4-1:0] node1110;
	wire [4-1:0] node1113;
	wire [4-1:0] node1116;
	wire [4-1:0] node1119;
	wire [4-1:0] node1121;
	wire [4-1:0] node1122;
	wire [4-1:0] node1123;
	wire [4-1:0] node1125;
	wire [4-1:0] node1126;
	wire [4-1:0] node1127;
	wire [4-1:0] node1130;
	wire [4-1:0] node1133;
	wire [4-1:0] node1135;
	wire [4-1:0] node1138;
	wire [4-1:0] node1139;
	wire [4-1:0] node1140;
	wire [4-1:0] node1141;
	wire [4-1:0] node1142;
	wire [4-1:0] node1146;
	wire [4-1:0] node1148;
	wire [4-1:0] node1151;
	wire [4-1:0] node1153;
	wire [4-1:0] node1156;
	wire [4-1:0] node1157;
	wire [4-1:0] node1158;
	wire [4-1:0] node1161;
	wire [4-1:0] node1164;
	wire [4-1:0] node1165;
	wire [4-1:0] node1166;
	wire [4-1:0] node1170;
	wire [4-1:0] node1174;
	wire [4-1:0] node1175;
	wire [4-1:0] node1176;
	wire [4-1:0] node1177;
	wire [4-1:0] node1178;
	wire [4-1:0] node1179;
	wire [4-1:0] node1180;
	wire [4-1:0] node1181;
	wire [4-1:0] node1182;
	wire [4-1:0] node1183;
	wire [4-1:0] node1186;
	wire [4-1:0] node1189;
	wire [4-1:0] node1192;
	wire [4-1:0] node1193;
	wire [4-1:0] node1194;
	wire [4-1:0] node1195;
	wire [4-1:0] node1199;
	wire [4-1:0] node1201;
	wire [4-1:0] node1206;
	wire [4-1:0] node1207;
	wire [4-1:0] node1208;
	wire [4-1:0] node1209;
	wire [4-1:0] node1210;
	wire [4-1:0] node1212;
	wire [4-1:0] node1215;
	wire [4-1:0] node1218;
	wire [4-1:0] node1220;
	wire [4-1:0] node1222;
	wire [4-1:0] node1225;
	wire [4-1:0] node1226;
	wire [4-1:0] node1229;
	wire [4-1:0] node1231;
	wire [4-1:0] node1233;
	wire [4-1:0] node1236;
	wire [4-1:0] node1237;
	wire [4-1:0] node1238;
	wire [4-1:0] node1240;
	wire [4-1:0] node1243;
	wire [4-1:0] node1244;
	wire [4-1:0] node1247;
	wire [4-1:0] node1250;
	wire [4-1:0] node1251;
	wire [4-1:0] node1252;
	wire [4-1:0] node1254;
	wire [4-1:0] node1257;
	wire [4-1:0] node1259;
	wire [4-1:0] node1262;
	wire [4-1:0] node1263;
	wire [4-1:0] node1266;
	wire [4-1:0] node1268;
	wire [4-1:0] node1272;
	wire [4-1:0] node1273;
	wire [4-1:0] node1274;
	wire [4-1:0] node1275;
	wire [4-1:0] node1276;
	wire [4-1:0] node1277;
	wire [4-1:0] node1278;
	wire [4-1:0] node1279;
	wire [4-1:0] node1282;
	wire [4-1:0] node1285;
	wire [4-1:0] node1287;
	wire [4-1:0] node1290;
	wire [4-1:0] node1293;
	wire [4-1:0] node1294;
	wire [4-1:0] node1295;
	wire [4-1:0] node1296;
	wire [4-1:0] node1300;
	wire [4-1:0] node1302;
	wire [4-1:0] node1305;
	wire [4-1:0] node1306;
	wire [4-1:0] node1307;
	wire [4-1:0] node1310;
	wire [4-1:0] node1314;
	wire [4-1:0] node1315;
	wire [4-1:0] node1316;
	wire [4-1:0] node1317;
	wire [4-1:0] node1319;
	wire [4-1:0] node1322;
	wire [4-1:0] node1325;
	wire [4-1:0] node1328;
	wire [4-1:0] node1329;
	wire [4-1:0] node1331;
	wire [4-1:0] node1333;
	wire [4-1:0] node1336;
	wire [4-1:0] node1338;
	wire [4-1:0] node1340;
	wire [4-1:0] node1343;
	wire [4-1:0] node1345;
	wire [4-1:0] node1346;
	wire [4-1:0] node1347;
	wire [4-1:0] node1349;
	wire [4-1:0] node1352;
	wire [4-1:0] node1354;
	wire [4-1:0] node1355;
	wire [4-1:0] node1358;
	wire [4-1:0] node1361;
	wire [4-1:0] node1362;
	wire [4-1:0] node1363;
	wire [4-1:0] node1367;
	wire [4-1:0] node1369;
	wire [4-1:0] node1371;
	wire [4-1:0] node1375;
	wire [4-1:0] node1376;
	wire [4-1:0] node1377;
	wire [4-1:0] node1378;
	wire [4-1:0] node1379;
	wire [4-1:0] node1380;
	wire [4-1:0] node1381;
	wire [4-1:0] node1382;
	wire [4-1:0] node1384;
	wire [4-1:0] node1387;
	wire [4-1:0] node1389;
	wire [4-1:0] node1392;
	wire [4-1:0] node1393;
	wire [4-1:0] node1394;
	wire [4-1:0] node1398;
	wire [4-1:0] node1399;
	wire [4-1:0] node1402;
	wire [4-1:0] node1405;
	wire [4-1:0] node1406;
	wire [4-1:0] node1407;
	wire [4-1:0] node1410;
	wire [4-1:0] node1413;
	wire [4-1:0] node1414;
	wire [4-1:0] node1416;
	wire [4-1:0] node1419;
	wire [4-1:0] node1421;
	wire [4-1:0] node1424;
	wire [4-1:0] node1425;
	wire [4-1:0] node1426;
	wire [4-1:0] node1427;
	wire [4-1:0] node1429;
	wire [4-1:0] node1432;
	wire [4-1:0] node1433;
	wire [4-1:0] node1436;
	wire [4-1:0] node1439;
	wire [4-1:0] node1440;
	wire [4-1:0] node1442;
	wire [4-1:0] node1445;
	wire [4-1:0] node1446;
	wire [4-1:0] node1450;
	wire [4-1:0] node1451;
	wire [4-1:0] node1452;
	wire [4-1:0] node1453;
	wire [4-1:0] node1458;
	wire [4-1:0] node1460;
	wire [4-1:0] node1463;
	wire [4-1:0] node1464;
	wire [4-1:0] node1465;
	wire [4-1:0] node1466;
	wire [4-1:0] node1467;
	wire [4-1:0] node1468;
	wire [4-1:0] node1472;
	wire [4-1:0] node1473;
	wire [4-1:0] node1477;
	wire [4-1:0] node1479;
	wire [4-1:0] node1482;
	wire [4-1:0] node1483;
	wire [4-1:0] node1484;
	wire [4-1:0] node1485;
	wire [4-1:0] node1489;
	wire [4-1:0] node1492;
	wire [4-1:0] node1493;
	wire [4-1:0] node1497;
	wire [4-1:0] node1498;
	wire [4-1:0] node1499;
	wire [4-1:0] node1502;
	wire [4-1:0] node1504;
	wire [4-1:0] node1505;
	wire [4-1:0] node1508;
	wire [4-1:0] node1511;
	wire [4-1:0] node1512;
	wire [4-1:0] node1514;
	wire [4-1:0] node1515;
	wire [4-1:0] node1519;
	wire [4-1:0] node1521;
	wire [4-1:0] node1522;
	wire [4-1:0] node1526;
	wire [4-1:0] node1527;
	wire [4-1:0] node1528;
	wire [4-1:0] node1529;
	wire [4-1:0] node1530;
	wire [4-1:0] node1531;
	wire [4-1:0] node1532;
	wire [4-1:0] node1537;
	wire [4-1:0] node1538;
	wire [4-1:0] node1542;
	wire [4-1:0] node1543;
	wire [4-1:0] node1544;
	wire [4-1:0] node1547;
	wire [4-1:0] node1550;
	wire [4-1:0] node1552;
	wire [4-1:0] node1553;
	wire [4-1:0] node1556;
	wire [4-1:0] node1559;
	wire [4-1:0] node1560;
	wire [4-1:0] node1561;
	wire [4-1:0] node1562;
	wire [4-1:0] node1563;
	wire [4-1:0] node1567;
	wire [4-1:0] node1570;
	wire [4-1:0] node1572;
	wire [4-1:0] node1575;
	wire [4-1:0] node1576;
	wire [4-1:0] node1578;
	wire [4-1:0] node1579;
	wire [4-1:0] node1583;
	wire [4-1:0] node1584;
	wire [4-1:0] node1585;
	wire [4-1:0] node1589;
	wire [4-1:0] node1592;
	wire [4-1:0] node1595;
	wire [4-1:0] node1596;
	wire [4-1:0] node1597;
	wire [4-1:0] node1598;
	wire [4-1:0] node1599;
	wire [4-1:0] node1600;
	wire [4-1:0] node1601;
	wire [4-1:0] node1602;
	wire [4-1:0] node1606;
	wire [4-1:0] node1608;
	wire [4-1:0] node1611;
	wire [4-1:0] node1612;
	wire [4-1:0] node1613;
	wire [4-1:0] node1618;
	wire [4-1:0] node1619;
	wire [4-1:0] node1621;
	wire [4-1:0] node1623;
	wire [4-1:0] node1626;
	wire [4-1:0] node1627;
	wire [4-1:0] node1630;
	wire [4-1:0] node1633;
	wire [4-1:0] node1634;
	wire [4-1:0] node1635;
	wire [4-1:0] node1636;
	wire [4-1:0] node1639;
	wire [4-1:0] node1642;
	wire [4-1:0] node1643;
	wire [4-1:0] node1644;
	wire [4-1:0] node1648;
	wire [4-1:0] node1651;
	wire [4-1:0] node1652;
	wire [4-1:0] node1654;
	wire [4-1:0] node1657;
	wire [4-1:0] node1658;
	wire [4-1:0] node1660;
	wire [4-1:0] node1664;
	wire [4-1:0] node1665;
	wire [4-1:0] node1666;
	wire [4-1:0] node1667;
	wire [4-1:0] node1670;
	wire [4-1:0] node1672;
	wire [4-1:0] node1674;
	wire [4-1:0] node1677;
	wire [4-1:0] node1678;
	wire [4-1:0] node1679;
	wire [4-1:0] node1680;
	wire [4-1:0] node1685;
	wire [4-1:0] node1686;
	wire [4-1:0] node1687;
	wire [4-1:0] node1691;
	wire [4-1:0] node1694;
	wire [4-1:0] node1695;
	wire [4-1:0] node1696;
	wire [4-1:0] node1697;
	wire [4-1:0] node1698;
	wire [4-1:0] node1702;
	wire [4-1:0] node1704;
	wire [4-1:0] node1708;
	wire [4-1:0] node1709;
	wire [4-1:0] node1711;
	wire [4-1:0] node1714;
	wire [4-1:0] node1715;
	wire [4-1:0] node1717;
	wire [4-1:0] node1720;
	wire [4-1:0] node1721;
	wire [4-1:0] node1725;
	wire [4-1:0] node1726;
	wire [4-1:0] node1727;
	wire [4-1:0] node1728;
	wire [4-1:0] node1729;
	wire [4-1:0] node1731;
	wire [4-1:0] node1734;
	wire [4-1:0] node1735;
	wire [4-1:0] node1738;
	wire [4-1:0] node1739;
	wire [4-1:0] node1743;
	wire [4-1:0] node1744;
	wire [4-1:0] node1746;
	wire [4-1:0] node1747;
	wire [4-1:0] node1751;
	wire [4-1:0] node1754;
	wire [4-1:0] node1755;
	wire [4-1:0] node1757;
	wire [4-1:0] node1758;
	wire [4-1:0] node1759;
	wire [4-1:0] node1763;
	wire [4-1:0] node1765;
	wire [4-1:0] node1768;
	wire [4-1:0] node1769;
	wire [4-1:0] node1772;
	wire [4-1:0] node1773;
	wire [4-1:0] node1777;
	wire [4-1:0] node1778;
	wire [4-1:0] node1779;
	wire [4-1:0] node1780;
	wire [4-1:0] node1781;
	wire [4-1:0] node1784;
	wire [4-1:0] node1787;
	wire [4-1:0] node1790;
	wire [4-1:0] node1791;
	wire [4-1:0] node1792;
	wire [4-1:0] node1794;
	wire [4-1:0] node1797;
	wire [4-1:0] node1798;
	wire [4-1:0] node1802;
	wire [4-1:0] node1803;
	wire [4-1:0] node1804;
	wire [4-1:0] node1809;
	wire [4-1:0] node1811;
	wire [4-1:0] node1812;
	wire [4-1:0] node1813;
	wire [4-1:0] node1817;
	wire [4-1:0] node1818;
	wire [4-1:0] node1822;
	wire [4-1:0] node1823;
	wire [4-1:0] node1824;
	wire [4-1:0] node1825;
	wire [4-1:0] node1826;
	wire [4-1:0] node1828;
	wire [4-1:0] node1829;
	wire [4-1:0] node1830;
	wire [4-1:0] node1831;
	wire [4-1:0] node1832;
	wire [4-1:0] node1839;
	wire [4-1:0] node1840;
	wire [4-1:0] node1841;
	wire [4-1:0] node1842;
	wire [4-1:0] node1843;
	wire [4-1:0] node1844;
	wire [4-1:0] node1847;
	wire [4-1:0] node1850;
	wire [4-1:0] node1853;
	wire [4-1:0] node1854;
	wire [4-1:0] node1857;
	wire [4-1:0] node1860;
	wire [4-1:0] node1861;
	wire [4-1:0] node1862;
	wire [4-1:0] node1863;
	wire [4-1:0] node1868;
	wire [4-1:0] node1869;
	wire [4-1:0] node1873;
	wire [4-1:0] node1875;
	wire [4-1:0] node1876;
	wire [4-1:0] node1877;
	wire [4-1:0] node1880;
	wire [4-1:0] node1883;
	wire [4-1:0] node1885;
	wire [4-1:0] node1887;
	wire [4-1:0] node1891;
	wire [4-1:0] node1892;
	wire [4-1:0] node1893;
	wire [4-1:0] node1894;
	wire [4-1:0] node1895;
	wire [4-1:0] node1896;
	wire [4-1:0] node1898;
	wire [4-1:0] node1899;
	wire [4-1:0] node1902;
	wire [4-1:0] node1905;
	wire [4-1:0] node1906;
	wire [4-1:0] node1908;
	wire [4-1:0] node1911;
	wire [4-1:0] node1912;
	wire [4-1:0] node1915;
	wire [4-1:0] node1918;
	wire [4-1:0] node1919;
	wire [4-1:0] node1920;
	wire [4-1:0] node1922;
	wire [4-1:0] node1925;
	wire [4-1:0] node1928;
	wire [4-1:0] node1929;
	wire [4-1:0] node1931;
	wire [4-1:0] node1934;
	wire [4-1:0] node1935;
	wire [4-1:0] node1938;
	wire [4-1:0] node1941;
	wire [4-1:0] node1942;
	wire [4-1:0] node1943;
	wire [4-1:0] node1944;
	wire [4-1:0] node1947;
	wire [4-1:0] node1948;
	wire [4-1:0] node1951;
	wire [4-1:0] node1954;
	wire [4-1:0] node1956;
	wire [4-1:0] node1959;
	wire [4-1:0] node1960;
	wire [4-1:0] node1962;
	wire [4-1:0] node1963;
	wire [4-1:0] node1966;
	wire [4-1:0] node1969;
	wire [4-1:0] node1970;
	wire [4-1:0] node1974;
	wire [4-1:0] node1975;
	wire [4-1:0] node1976;
	wire [4-1:0] node1977;
	wire [4-1:0] node1978;
	wire [4-1:0] node1981;
	wire [4-1:0] node1982;
	wire [4-1:0] node1985;
	wire [4-1:0] node1988;
	wire [4-1:0] node1989;
	wire [4-1:0] node1990;
	wire [4-1:0] node1995;
	wire [4-1:0] node1996;
	wire [4-1:0] node1998;
	wire [4-1:0] node1999;
	wire [4-1:0] node2004;
	wire [4-1:0] node2005;
	wire [4-1:0] node2006;
	wire [4-1:0] node2009;
	wire [4-1:0] node2012;
	wire [4-1:0] node2013;
	wire [4-1:0] node2016;
	wire [4-1:0] node2017;
	wire [4-1:0] node2018;
	wire [4-1:0] node2023;
	wire [4-1:0] node2024;
	wire [4-1:0] node2026;
	wire [4-1:0] node2027;
	wire [4-1:0] node2028;
	wire [4-1:0] node2030;
	wire [4-1:0] node2033;
	wire [4-1:0] node2034;
	wire [4-1:0] node2036;
	wire [4-1:0] node2041;
	wire [4-1:0] node2042;
	wire [4-1:0] node2043;
	wire [4-1:0] node2044;
	wire [4-1:0] node2045;
	wire [4-1:0] node2046;
	wire [4-1:0] node2049;
	wire [4-1:0] node2052;
	wire [4-1:0] node2055;
	wire [4-1:0] node2056;
	wire [4-1:0] node2057;
	wire [4-1:0] node2060;
	wire [4-1:0] node2063;
	wire [4-1:0] node2066;
	wire [4-1:0] node2067;
	wire [4-1:0] node2068;
	wire [4-1:0] node2072;
	wire [4-1:0] node2073;
	wire [4-1:0] node2076;
	wire [4-1:0] node2079;
	wire [4-1:0] node2081;
	wire [4-1:0] node2082;
	wire [4-1:0] node2083;
	wire [4-1:0] node2084;
	wire [4-1:0] node2089;
	wire [4-1:0] node2091;
	wire [4-1:0] node2094;
	wire [4-1:0] node2095;
	wire [4-1:0] node2096;
	wire [4-1:0] node2097;
	wire [4-1:0] node2098;
	wire [4-1:0] node2100;
	wire [4-1:0] node2101;
	wire [4-1:0] node2103;
	wire [4-1:0] node2107;
	wire [4-1:0] node2108;
	wire [4-1:0] node2109;
	wire [4-1:0] node2110;
	wire [4-1:0] node2113;
	wire [4-1:0] node2114;
	wire [4-1:0] node2118;
	wire [4-1:0] node2119;
	wire [4-1:0] node2120;
	wire [4-1:0] node2123;
	wire [4-1:0] node2126;
	wire [4-1:0] node2127;
	wire [4-1:0] node2131;
	wire [4-1:0] node2132;
	wire [4-1:0] node2134;
	wire [4-1:0] node2136;
	wire [4-1:0] node2139;
	wire [4-1:0] node2140;
	wire [4-1:0] node2143;
	wire [4-1:0] node2146;
	wire [4-1:0] node2148;
	wire [4-1:0] node2149;
	wire [4-1:0] node2151;
	wire [4-1:0] node2153;
	wire [4-1:0] node2157;
	wire [4-1:0] node2158;
	wire [4-1:0] node2159;
	wire [4-1:0] node2160;
	wire [4-1:0] node2161;
	wire [4-1:0] node2163;
	wire [4-1:0] node2166;
	wire [4-1:0] node2167;
	wire [4-1:0] node2169;
	wire [4-1:0] node2172;
	wire [4-1:0] node2173;
	wire [4-1:0] node2176;
	wire [4-1:0] node2179;
	wire [4-1:0] node2180;
	wire [4-1:0] node2183;
	wire [4-1:0] node2184;
	wire [4-1:0] node2186;
	wire [4-1:0] node2189;
	wire [4-1:0] node2192;
	wire [4-1:0] node2193;
	wire [4-1:0] node2194;
	wire [4-1:0] node2195;
	wire [4-1:0] node2197;
	wire [4-1:0] node2201;
	wire [4-1:0] node2204;
	wire [4-1:0] node2205;
	wire [4-1:0] node2208;
	wire [4-1:0] node2209;
	wire [4-1:0] node2211;
	wire [4-1:0] node2215;
	wire [4-1:0] node2216;
	wire [4-1:0] node2217;
	wire [4-1:0] node2218;
	wire [4-1:0] node2219;
	wire [4-1:0] node2223;
	wire [4-1:0] node2224;
	wire [4-1:0] node2227;
	wire [4-1:0] node2230;
	wire [4-1:0] node2231;
	wire [4-1:0] node2233;
	wire [4-1:0] node2234;
	wire [4-1:0] node2238;
	wire [4-1:0] node2241;
	wire [4-1:0] node2242;
	wire [4-1:0] node2243;
	wire [4-1:0] node2244;
	wire [4-1:0] node2247;
	wire [4-1:0] node2248;
	wire [4-1:0] node2251;
	wire [4-1:0] node2255;
	wire [4-1:0] node2256;
	wire [4-1:0] node2260;
	wire [4-1:0] node2262;
	wire [4-1:0] node2263;
	wire [4-1:0] node2264;
	wire [4-1:0] node2265;
	wire [4-1:0] node2267;
	wire [4-1:0] node2269;
	wire [4-1:0] node2273;
	wire [4-1:0] node2274;
	wire [4-1:0] node2275;
	wire [4-1:0] node2276;
	wire [4-1:0] node2279;
	wire [4-1:0] node2282;
	wire [4-1:0] node2283;
	wire [4-1:0] node2287;
	wire [4-1:0] node2288;
	wire [4-1:0] node2289;
	wire [4-1:0] node2290;
	wire [4-1:0] node2294;
	wire [4-1:0] node2296;
	wire [4-1:0] node2299;
	wire [4-1:0] node2300;
	wire [4-1:0] node2303;
	wire [4-1:0] node2304;
	wire [4-1:0] node2308;
	wire [4-1:0] node2309;
	wire [4-1:0] node2311;
	wire [4-1:0] node2312;

	assign outp = (inp[8]) ? node1174 : node1;
		assign node1 = (inp[9]) ? node623 : node2;
			assign node2 = (inp[15]) ? node322 : node3;
				assign node3 = (inp[6]) ? node95 : node4;
					assign node4 = (inp[0]) ? 4'b1101 : node5;
						assign node5 = (inp[2]) ? node73 : node6;
							assign node6 = (inp[3]) ? node42 : node7;
								assign node7 = (inp[4]) ? node21 : node8;
									assign node8 = (inp[7]) ? node14 : node9;
										assign node9 = (inp[13]) ? 4'b1001 : node10;
											assign node10 = (inp[5]) ? 4'b0000 : 4'b0001;
										assign node14 = (inp[5]) ? node16 : 4'b1111;
											assign node16 = (inp[12]) ? node18 : 4'b0100;
												assign node18 = (inp[11]) ? 4'b0100 : 4'b1100;
									assign node21 = (inp[10]) ? node33 : node22;
										assign node22 = (inp[11]) ? node28 : node23;
											assign node23 = (inp[7]) ? node25 : 4'b1001;
												assign node25 = (inp[14]) ? 4'b1101 : 4'b1001;
											assign node28 = (inp[13]) ? 4'b1001 : node29;
												assign node29 = (inp[1]) ? 4'b0001 : 4'b0000;
										assign node33 = (inp[13]) ? node39 : node34;
											assign node34 = (inp[7]) ? node36 : 4'b0000;
												assign node36 = (inp[5]) ? 4'b0001 : 4'b0000;
											assign node39 = (inp[1]) ? 4'b1001 : 4'b0001;
								assign node42 = (inp[1]) ? node62 : node43;
									assign node43 = (inp[14]) ? node53 : node44;
										assign node44 = (inp[4]) ? node48 : node45;
											assign node45 = (inp[11]) ? 4'b1000 : 4'b1100;
											assign node48 = (inp[10]) ? 4'b0100 : node49;
												assign node49 = (inp[11]) ? 4'b1100 : 4'b0100;
										assign node53 = (inp[13]) ? node57 : node54;
											assign node54 = (inp[12]) ? 4'b1001 : 4'b0000;
											assign node57 = (inp[5]) ? 4'b0101 : node58;
												assign node58 = (inp[11]) ? 4'b1100 : 4'b1101;
									assign node62 = (inp[13]) ? node66 : node63;
										assign node63 = (inp[5]) ? 4'b0001 : 4'b0101;
										assign node66 = (inp[4]) ? 4'b1101 : node67;
											assign node67 = (inp[7]) ? node69 : 4'b1101;
												assign node69 = (inp[14]) ? 4'b0001 : 4'b1001;
							assign node73 = (inp[5]) ? node75 : 4'b1111;
								assign node75 = (inp[4]) ? node85 : node76;
									assign node76 = (inp[3]) ? node80 : node77;
										assign node77 = (inp[7]) ? 4'b1111 : 4'b1001;
										assign node80 = (inp[7]) ? 4'b1001 : node81;
											assign node81 = (inp[13]) ? 4'b1101 : 4'b0101;
									assign node85 = (inp[10]) ? node91 : node86;
										assign node86 = (inp[13]) ? node88 : 4'b1001;
											assign node88 = (inp[12]) ? 4'b0001 : 4'b1001;
										assign node91 = (inp[13]) ? 4'b1000 : 4'b0000;
					assign node95 = (inp[5]) ? node205 : node96;
						assign node96 = (inp[0]) ? node170 : node97;
							assign node97 = (inp[11]) ? node139 : node98;
								assign node98 = (inp[14]) ? node120 : node99;
									assign node99 = (inp[4]) ? node111 : node100;
										assign node100 = (inp[1]) ? node106 : node101;
											assign node101 = (inp[3]) ? node103 : 4'b0000;
												assign node103 = (inp[12]) ? 4'b0001 : 4'b0000;
											assign node106 = (inp[3]) ? 4'b0001 : node107;
												assign node107 = (inp[7]) ? 4'b0101 : 4'b0001;
										assign node111 = (inp[7]) ? node117 : node112;
											assign node112 = (inp[2]) ? 4'b1001 : node113;
												assign node113 = (inp[13]) ? 4'b1100 : 4'b1000;
											assign node117 = (inp[12]) ? 4'b0100 : 4'b0000;
									assign node120 = (inp[4]) ? node126 : node121;
										assign node121 = (inp[13]) ? node123 : 4'b1101;
											assign node123 = (inp[7]) ? 4'b0000 : 4'b1000;
										assign node126 = (inp[7]) ? node132 : node127;
											assign node127 = (inp[1]) ? 4'b1101 : node128;
												assign node128 = (inp[2]) ? 4'b1100 : 4'b0100;
											assign node132 = (inp[12]) ? node136 : node133;
												assign node133 = (inp[13]) ? 4'b0100 : 4'b0000;
												assign node136 = (inp[3]) ? 4'b1000 : 4'b0100;
								assign node139 = (inp[4]) ? node153 : node140;
									assign node140 = (inp[1]) ? node148 : node141;
										assign node141 = (inp[3]) ? node143 : 4'b1100;
											assign node143 = (inp[7]) ? node145 : 4'b1001;
												assign node145 = (inp[12]) ? 4'b0101 : 4'b1101;
										assign node148 = (inp[3]) ? 4'b0001 : node149;
											assign node149 = (inp[10]) ? 4'b1001 : 4'b0001;
									assign node153 = (inp[7]) ? node161 : node154;
										assign node154 = (inp[12]) ? node156 : 4'b0101;
											assign node156 = (inp[10]) ? 4'b0101 : node157;
												assign node157 = (inp[13]) ? 4'b0100 : 4'b1001;
										assign node161 = (inp[10]) ? 4'b1101 : node162;
											assign node162 = (inp[12]) ? node166 : node163;
												assign node163 = (inp[3]) ? 4'b0001 : 4'b0101;
												assign node166 = (inp[3]) ? 4'b1000 : 4'b1001;
							assign node170 = (inp[2]) ? 4'b1101 : node171;
								assign node171 = (inp[3]) ? node185 : node172;
									assign node172 = (inp[12]) ? node180 : node173;
										assign node173 = (inp[10]) ? node175 : 4'b0000;
											assign node175 = (inp[11]) ? node177 : 4'b0001;
												assign node177 = (inp[7]) ? 4'b1101 : 4'b0001;
										assign node180 = (inp[1]) ? node182 : 4'b1101;
											assign node182 = (inp[11]) ? 4'b0001 : 4'b0000;
									assign node185 = (inp[13]) ? node197 : node186;
										assign node186 = (inp[4]) ? node192 : node187;
											assign node187 = (inp[14]) ? 4'b1001 : node188;
												assign node188 = (inp[7]) ? 4'b0000 : 4'b1000;
											assign node192 = (inp[1]) ? 4'b0101 : node193;
												assign node193 = (inp[14]) ? 4'b1100 : 4'b0100;
										assign node197 = (inp[12]) ? 4'b0101 : node198;
											assign node198 = (inp[4]) ? node200 : 4'b1100;
												assign node200 = (inp[14]) ? 4'b1100 : 4'b1101;
						assign node205 = (inp[3]) ? node259 : node206;
							assign node206 = (inp[4]) ? node238 : node207;
								assign node207 = (inp[2]) ? node223 : node208;
									assign node208 = (inp[7]) ? node214 : node209;
										assign node209 = (inp[12]) ? 4'b0001 : node210;
											assign node210 = (inp[1]) ? 4'b1001 : 4'b0001;
										assign node214 = (inp[13]) ? node220 : node215;
											assign node215 = (inp[14]) ? node217 : 4'b0101;
												assign node217 = (inp[12]) ? 4'b0100 : 4'b0101;
											assign node220 = (inp[1]) ? 4'b1001 : 4'b0101;
									assign node223 = (inp[11]) ? node231 : node224;
										assign node224 = (inp[0]) ? 4'b1101 : node225;
											assign node225 = (inp[13]) ? node227 : 4'b1100;
												assign node227 = (inp[7]) ? 4'b1000 : 4'b1100;
										assign node231 = (inp[10]) ? 4'b1101 : node232;
											assign node232 = (inp[7]) ? node234 : 4'b0000;
												assign node234 = (inp[0]) ? 4'b1101 : 4'b0101;
								assign node238 = (inp[1]) ? node250 : node239;
									assign node239 = (inp[14]) ? node245 : node240;
										assign node240 = (inp[7]) ? node242 : 4'b0000;
											assign node242 = (inp[13]) ? 4'b0000 : 4'b1000;
										assign node245 = (inp[13]) ? node247 : 4'b0101;
											assign node247 = (inp[2]) ? 4'b0001 : 4'b1000;
									assign node250 = (inp[0]) ? node256 : node251;
										assign node251 = (inp[13]) ? node253 : 4'b1000;
											assign node253 = (inp[10]) ? 4'b1001 : 4'b0001;
										assign node256 = (inp[10]) ? 4'b0001 : 4'b0101;
							assign node259 = (inp[1]) ? node295 : node260;
								assign node260 = (inp[4]) ? node282 : node261;
									assign node261 = (inp[2]) ? node273 : node262;
										assign node262 = (inp[13]) ? node268 : node263;
											assign node263 = (inp[10]) ? 4'b0000 : node264;
												assign node264 = (inp[11]) ? 4'b1001 : 4'b0001;
											assign node268 = (inp[12]) ? 4'b0000 : node269;
												assign node269 = (inp[7]) ? 4'b0000 : 4'b0001;
										assign node273 = (inp[13]) ? node277 : node274;
											assign node274 = (inp[0]) ? 4'b0000 : 4'b1000;
											assign node277 = (inp[14]) ? node279 : 4'b0001;
												assign node279 = (inp[12]) ? 4'b0000 : 4'b1000;
									assign node282 = (inp[12]) ? node288 : node283;
										assign node283 = (inp[11]) ? node285 : 4'b0000;
											assign node285 = (inp[7]) ? 4'b1000 : 4'b0000;
										assign node288 = (inp[11]) ? 4'b0000 : node289;
											assign node289 = (inp[7]) ? 4'b0001 : node290;
												assign node290 = (inp[14]) ? 4'b0001 : 4'b0000;
								assign node295 = (inp[11]) ? node311 : node296;
									assign node296 = (inp[14]) ? node306 : node297;
										assign node297 = (inp[4]) ? node301 : node298;
											assign node298 = (inp[7]) ? 4'b1001 : 4'b0001;
											assign node301 = (inp[12]) ? node303 : 4'b0001;
												assign node303 = (inp[10]) ? 4'b0000 : 4'b0000;
										assign node306 = (inp[0]) ? 4'b0000 : node307;
											assign node307 = (inp[12]) ? 4'b0000 : 4'b1000;
									assign node311 = (inp[13]) ? node317 : node312;
										assign node312 = (inp[4]) ? node314 : 4'b0001;
											assign node314 = (inp[10]) ? 4'b0001 : 4'b1001;
										assign node317 = (inp[10]) ? 4'b1001 : node318;
											assign node318 = (inp[0]) ? 4'b0001 : 4'b1001;
				assign node322 = (inp[6]) ? node410 : node323;
					assign node323 = (inp[0]) ? 4'b1001 : node324;
						assign node324 = (inp[2]) ? node386 : node325;
							assign node325 = (inp[5]) ? node345 : node326;
								assign node326 = (inp[3]) ? node328 : 4'b1011;
									assign node328 = (inp[4]) ? node336 : node329;
										assign node329 = (inp[14]) ? node333 : node330;
											assign node330 = (inp[12]) ? 4'b1011 : 4'b1001;
											assign node333 = (inp[1]) ? 4'b1000 : 4'b0001;
										assign node336 = (inp[12]) ? node340 : node337;
											assign node337 = (inp[13]) ? 4'b1001 : 4'b0001;
											assign node340 = (inp[14]) ? node342 : 4'b0000;
												assign node342 = (inp[11]) ? 4'b0000 : 4'b0001;
								assign node345 = (inp[3]) ? node367 : node346;
									assign node346 = (inp[7]) ? node358 : node347;
										assign node347 = (inp[12]) ? node353 : node348;
											assign node348 = (inp[13]) ? node350 : 4'b0100;
												assign node350 = (inp[11]) ? 4'b1101 : 4'b1100;
											assign node353 = (inp[14]) ? node355 : 4'b0100;
												assign node355 = (inp[11]) ? 4'b0101 : 4'b0100;
										assign node358 = (inp[4]) ? node360 : 4'b1001;
											assign node360 = (inp[13]) ? node364 : node361;
												assign node361 = (inp[1]) ? 4'b1001 : 4'b1000;
												assign node364 = (inp[12]) ? 4'b1101 : 4'b1100;
									assign node367 = (inp[4]) ? node375 : node368;
										assign node368 = (inp[10]) ? node372 : node369;
											assign node369 = (inp[7]) ? 4'b1100 : 4'b1101;
											assign node372 = (inp[12]) ? 4'b1000 : 4'b1001;
										assign node375 = (inp[1]) ? node381 : node376;
											assign node376 = (inp[13]) ? node378 : 4'b0000;
												assign node378 = (inp[10]) ? 4'b1001 : 4'b0001;
											assign node381 = (inp[10]) ? node383 : 4'b1001;
												assign node383 = (inp[13]) ? 4'b1001 : 4'b0001;
							assign node386 = (inp[3]) ? node388 : 4'b1011;
								assign node388 = (inp[5]) ? node390 : 4'b1011;
									assign node390 = (inp[4]) ? node400 : node391;
										assign node391 = (inp[7]) ? 4'b1011 : node392;
											assign node392 = (inp[11]) ? node396 : node393;
												assign node393 = (inp[13]) ? 4'b1001 : 4'b1011;
												assign node396 = (inp[1]) ? 4'b1001 : 4'b0000;
										assign node400 = (inp[11]) ? node406 : node401;
											assign node401 = (inp[7]) ? 4'b0001 : node402;
												assign node402 = (inp[14]) ? 4'b0000 : 4'b0001;
											assign node406 = (inp[14]) ? 4'b1000 : 4'b0000;
					assign node410 = (inp[0]) ? node548 : node411;
						assign node411 = (inp[1]) ? node473 : node412;
							assign node412 = (inp[4]) ? node448 : node413;
								assign node413 = (inp[12]) ? node433 : node414;
									assign node414 = (inp[5]) ? node424 : node415;
										assign node415 = (inp[10]) ? 4'b1100 : node416;
											assign node416 = (inp[3]) ? node420 : node417;
												assign node417 = (inp[11]) ? 4'b0100 : 4'b0000;
												assign node420 = (inp[7]) ? 4'b0100 : 4'b1101;
										assign node424 = (inp[7]) ? node430 : node425;
											assign node425 = (inp[3]) ? 4'b0001 : node426;
												assign node426 = (inp[14]) ? 4'b0100 : 4'b0101;
											assign node430 = (inp[13]) ? 4'b1101 : 4'b1001;
									assign node433 = (inp[7]) ? node439 : node434;
										assign node434 = (inp[3]) ? node436 : 4'b0101;
											assign node436 = (inp[5]) ? 4'b0000 : 4'b0001;
										assign node439 = (inp[3]) ? node445 : node440;
											assign node440 = (inp[14]) ? node442 : 4'b1000;
												assign node442 = (inp[5]) ? 4'b0000 : 4'b0001;
											assign node445 = (inp[14]) ? 4'b1100 : 4'b0100;
								assign node448 = (inp[11]) ? node462 : node449;
									assign node449 = (inp[5]) ? node457 : node450;
										assign node450 = (inp[2]) ? node452 : 4'b0000;
											assign node452 = (inp[7]) ? node454 : 4'b1000;
												assign node454 = (inp[13]) ? 4'b0100 : 4'b0000;
										assign node457 = (inp[14]) ? node459 : 4'b0001;
											assign node459 = (inp[12]) ? 4'b0001 : 4'b0000;
									assign node462 = (inp[13]) ? node468 : node463;
										assign node463 = (inp[12]) ? node465 : 4'b0001;
											assign node465 = (inp[7]) ? 4'b0101 : 4'b1101;
										assign node468 = (inp[7]) ? node470 : 4'b1000;
											assign node470 = (inp[5]) ? 4'b0000 : 4'b0001;
							assign node473 = (inp[3]) ? node511 : node474;
								assign node474 = (inp[13]) ? node490 : node475;
									assign node475 = (inp[7]) ? node479 : node476;
										assign node476 = (inp[10]) ? 4'b0101 : 4'b0001;
										assign node479 = (inp[2]) ? node485 : node480;
											assign node480 = (inp[14]) ? node482 : 4'b0101;
												assign node482 = (inp[5]) ? 4'b0001 : 4'b1000;
											assign node485 = (inp[11]) ? node487 : 4'b1001;
												assign node487 = (inp[4]) ? 4'b1001 : 4'b0001;
									assign node490 = (inp[2]) ? node502 : node491;
										assign node491 = (inp[14]) ? node497 : node492;
											assign node492 = (inp[4]) ? 4'b1000 : node493;
												assign node493 = (inp[7]) ? 4'b0101 : 4'b1101;
											assign node497 = (inp[12]) ? node499 : 4'b1001;
												assign node499 = (inp[5]) ? 4'b0001 : 4'b0000;
										assign node502 = (inp[12]) ? node508 : node503;
											assign node503 = (inp[14]) ? 4'b1101 : node504;
												assign node504 = (inp[10]) ? 4'b1001 : 4'b1101;
											assign node508 = (inp[11]) ? 4'b1101 : 4'b0101;
								assign node511 = (inp[11]) ? node537 : node512;
									assign node512 = (inp[5]) ? node524 : node513;
										assign node513 = (inp[12]) ? node521 : node514;
											assign node514 = (inp[7]) ? node518 : node515;
												assign node515 = (inp[13]) ? 4'b1001 : 4'b1000;
												assign node518 = (inp[13]) ? 4'b1101 : 4'b0100;
											assign node521 = (inp[10]) ? 4'b0001 : 4'b0000;
										assign node524 = (inp[12]) ? node530 : node525;
											assign node525 = (inp[4]) ? 4'b0001 : node526;
												assign node526 = (inp[2]) ? 4'b1000 : 4'b0000;
											assign node530 = (inp[2]) ? node534 : node531;
												assign node531 = (inp[4]) ? 4'b0000 : 4'b1000;
												assign node534 = (inp[10]) ? 4'b1001 : 4'b1000;
									assign node537 = (inp[10]) ? node543 : node538;
										assign node538 = (inp[7]) ? 4'b0001 : node539;
											assign node539 = (inp[5]) ? 4'b0001 : 4'b0101;
										assign node543 = (inp[4]) ? node545 : 4'b1001;
											assign node545 = (inp[5]) ? 4'b0000 : 4'b1001;
						assign node548 = (inp[5]) ? node572 : node549;
							assign node549 = (inp[3]) ? node551 : 4'b1001;
								assign node551 = (inp[4]) ? node557 : node552;
									assign node552 = (inp[12]) ? 4'b1001 : node553;
										assign node553 = (inp[7]) ? 4'b1001 : 4'b1000;
									assign node557 = (inp[2]) ? 4'b1001 : node558;
										assign node558 = (inp[13]) ? node564 : node559;
											assign node559 = (inp[10]) ? node561 : 4'b1001;
												assign node561 = (inp[1]) ? 4'b0001 : 4'b0000;
											assign node564 = (inp[14]) ? node568 : node565;
												assign node565 = (inp[1]) ? 4'b1001 : 4'b1000;
												assign node568 = (inp[1]) ? 4'b1000 : 4'b0001;
							assign node572 = (inp[2]) ? node606 : node573;
								assign node573 = (inp[12]) ? node589 : node574;
									assign node574 = (inp[14]) ? 4'b0001 : node575;
										assign node575 = (inp[13]) ? node583 : node576;
											assign node576 = (inp[3]) ? node580 : node577;
												assign node577 = (inp[1]) ? 4'b0101 : 4'b0100;
												assign node580 = (inp[1]) ? 4'b0001 : 4'b0000;
											assign node583 = (inp[7]) ? node585 : 4'b1101;
												assign node585 = (inp[4]) ? 4'b1000 : 4'b1001;
									assign node589 = (inp[1]) ? node599 : node590;
										assign node590 = (inp[11]) ? node596 : node591;
											assign node591 = (inp[13]) ? node593 : 4'b1000;
												assign node593 = (inp[14]) ? 4'b0000 : 4'b0000;
											assign node596 = (inp[3]) ? 4'b0000 : 4'b1000;
										assign node599 = (inp[7]) ? 4'b1001 : node600;
											assign node600 = (inp[13]) ? 4'b1000 : node601;
												assign node601 = (inp[14]) ? 4'b0001 : 4'b0000;
								assign node606 = (inp[3]) ? node608 : 4'b1001;
									assign node608 = (inp[7]) ? node616 : node609;
										assign node609 = (inp[1]) ? 4'b0001 : node610;
											assign node610 = (inp[11]) ? node612 : 4'b0000;
												assign node612 = (inp[12]) ? 4'b1000 : 4'b0000;
										assign node616 = (inp[4]) ? node618 : 4'b1001;
											assign node618 = (inp[14]) ? 4'b1001 : node619;
												assign node619 = (inp[1]) ? 4'b0001 : 4'b0000;
			assign node623 = (inp[15]) ? node935 : node624;
				assign node624 = (inp[6]) ? node720 : node625;
					assign node625 = (inp[0]) ? 4'b0101 : node626;
						assign node626 = (inp[5]) ? node654 : node627;
							assign node627 = (inp[2]) ? 4'b0111 : node628;
								assign node628 = (inp[4]) ? node638 : node629;
									assign node629 = (inp[3]) ? node635 : node630;
										assign node630 = (inp[14]) ? 4'b0111 : node631;
											assign node631 = (inp[10]) ? 4'b0000 : 4'b0111;
										assign node635 = (inp[1]) ? 4'b1000 : 4'b0101;
									assign node638 = (inp[1]) ? node644 : node639;
										assign node639 = (inp[12]) ? 4'b0111 : node640;
											assign node640 = (inp[11]) ? 4'b0100 : 4'b0000;
										assign node644 = (inp[14]) ? node650 : node645;
											assign node645 = (inp[3]) ? 4'b1001 : node646;
												assign node646 = (inp[13]) ? 4'b0001 : 4'b0111;
											assign node650 = (inp[12]) ? 4'b0000 : 4'b1000;
							assign node654 = (inp[3]) ? node680 : node655;
								assign node655 = (inp[13]) ? node663 : node656;
									assign node656 = (inp[2]) ? 4'b0111 : node657;
										assign node657 = (inp[12]) ? 4'b0100 : node658;
											assign node658 = (inp[7]) ? 4'b1100 : 4'b1101;
									assign node663 = (inp[14]) ? node669 : node664;
										assign node664 = (inp[1]) ? node666 : 4'b0000;
											assign node666 = (inp[11]) ? 4'b1101 : 4'b0001;
										assign node669 = (inp[1]) ? node675 : node670;
											assign node670 = (inp[12]) ? node672 : 4'b0111;
												assign node672 = (inp[2]) ? 4'b0000 : 4'b1100;
											assign node675 = (inp[10]) ? 4'b0000 : node676;
												assign node676 = (inp[4]) ? 4'b0000 : 4'b0100;
								assign node680 = (inp[4]) ? node704 : node681;
									assign node681 = (inp[7]) ? node693 : node682;
										assign node682 = (inp[13]) ? node688 : node683;
											assign node683 = (inp[14]) ? 4'b0001 : node684;
												assign node684 = (inp[1]) ? 4'b0001 : 4'b1000;
											assign node688 = (inp[10]) ? 4'b0100 : node689;
												assign node689 = (inp[11]) ? 4'b0101 : 4'b1000;
										assign node693 = (inp[12]) ? node697 : node694;
											assign node694 = (inp[13]) ? 4'b0000 : 4'b1000;
											assign node697 = (inp[1]) ? node701 : node698;
												assign node698 = (inp[14]) ? 4'b1001 : 4'b1000;
												assign node701 = (inp[13]) ? 4'b0001 : 4'b1001;
									assign node704 = (inp[10]) ? node712 : node705;
										assign node705 = (inp[7]) ? node709 : node706;
											assign node706 = (inp[14]) ? 4'b1101 : 4'b1100;
											assign node709 = (inp[1]) ? 4'b1001 : 4'b1000;
										assign node712 = (inp[13]) ? node716 : node713;
											assign node713 = (inp[1]) ? 4'b1101 : 4'b1100;
											assign node716 = (inp[7]) ? 4'b0100 : 4'b0101;
					assign node720 = (inp[5]) ? node810 : node721;
						assign node721 = (inp[0]) ? node787 : node722;
							assign node722 = (inp[11]) ? node756 : node723;
								assign node723 = (inp[3]) ? node741 : node724;
									assign node724 = (inp[4]) ? node732 : node725;
										assign node725 = (inp[13]) ? node727 : 4'b0101;
											assign node727 = (inp[7]) ? node729 : 4'b0000;
												assign node729 = (inp[10]) ? 4'b0000 : 4'b0100;
										assign node732 = (inp[2]) ? node736 : node733;
											assign node733 = (inp[12]) ? 4'b0000 : 4'b0100;
											assign node736 = (inp[13]) ? 4'b1101 : node737;
												assign node737 = (inp[14]) ? 4'b0100 : 4'b1100;
									assign node741 = (inp[7]) ? node747 : node742;
										assign node742 = (inp[2]) ? 4'b0100 : node743;
											assign node743 = (inp[12]) ? 4'b0001 : 4'b1101;
										assign node747 = (inp[10]) ? node753 : node748;
											assign node748 = (inp[2]) ? node750 : 4'b1100;
												assign node750 = (inp[12]) ? 4'b0001 : 4'b1001;
											assign node753 = (inp[14]) ? 4'b1000 : 4'b0000;
								assign node756 = (inp[12]) ? node770 : node757;
									assign node757 = (inp[10]) ? node765 : node758;
										assign node758 = (inp[4]) ? 4'b1001 : node759;
											assign node759 = (inp[2]) ? 4'b1001 : node760;
												assign node760 = (inp[13]) ? 4'b1001 : 4'b1101;
										assign node765 = (inp[7]) ? 4'b0101 : node766;
											assign node766 = (inp[4]) ? 4'b1001 : 4'b0001;
									assign node770 = (inp[10]) ? node780 : node771;
										assign node771 = (inp[2]) ? node775 : node772;
											assign node772 = (inp[4]) ? 4'b0001 : 4'b0101;
											assign node775 = (inp[13]) ? node777 : 4'b0000;
												assign node777 = (inp[14]) ? 4'b0101 : 4'b1000;
										assign node780 = (inp[2]) ? node784 : node781;
											assign node781 = (inp[13]) ? 4'b1000 : 4'b1001;
											assign node784 = (inp[3]) ? 4'b0101 : 4'b1101;
							assign node787 = (inp[2]) ? 4'b0101 : node788;
								assign node788 = (inp[3]) ? node802 : node789;
									assign node789 = (inp[13]) ? node795 : node790;
										assign node790 = (inp[7]) ? 4'b0101 : node791;
											assign node791 = (inp[4]) ? 4'b1000 : 4'b0101;
										assign node795 = (inp[10]) ? node797 : 4'b0101;
											assign node797 = (inp[7]) ? 4'b0001 : node798;
												assign node798 = (inp[12]) ? 4'b0001 : 4'b0000;
									assign node802 = (inp[7]) ? node806 : node803;
										assign node803 = (inp[4]) ? 4'b0100 : 4'b1001;
										assign node806 = (inp[12]) ? 4'b1001 : 4'b1000;
						assign node810 = (inp[3]) ? node870 : node811;
							assign node811 = (inp[4]) ? node839 : node812;
								assign node812 = (inp[0]) ? node826 : node813;
									assign node813 = (inp[10]) ? node819 : node814;
										assign node814 = (inp[11]) ? node816 : 4'b1100;
											assign node816 = (inp[1]) ? 4'b1101 : 4'b1001;
										assign node819 = (inp[14]) ? 4'b0001 : node820;
											assign node820 = (inp[7]) ? node822 : 4'b1101;
												assign node822 = (inp[12]) ? 4'b0100 : 4'b0101;
									assign node826 = (inp[2]) ? node834 : node827;
										assign node827 = (inp[13]) ? 4'b0001 : node828;
											assign node828 = (inp[1]) ? node830 : 4'b1100;
												assign node830 = (inp[14]) ? 4'b0000 : 4'b1101;
										assign node834 = (inp[11]) ? node836 : 4'b0101;
											assign node836 = (inp[12]) ? 4'b0101 : 4'b0000;
								assign node839 = (inp[11]) ? node861 : node840;
									assign node840 = (inp[14]) ? node856 : node841;
										assign node841 = (inp[2]) ? node849 : node842;
											assign node842 = (inp[7]) ? node846 : node843;
												assign node843 = (inp[12]) ? 4'b0000 : 4'b0100;
												assign node846 = (inp[12]) ? 4'b1000 : 4'b0000;
											assign node849 = (inp[13]) ? node853 : node850;
												assign node850 = (inp[0]) ? 4'b1000 : 4'b0001;
												assign node853 = (inp[1]) ? 4'b0001 : 4'b0000;
										assign node856 = (inp[0]) ? 4'b0101 : node857;
											assign node857 = (inp[1]) ? 4'b1000 : 4'b1001;
									assign node861 = (inp[1]) ? 4'b0001 : node862;
										assign node862 = (inp[10]) ? 4'b0101 : node863;
											assign node863 = (inp[13]) ? node865 : 4'b1000;
												assign node865 = (inp[2]) ? 4'b0000 : 4'b0001;
							assign node870 = (inp[4]) ? node908 : node871;
								assign node871 = (inp[10]) ? node887 : node872;
									assign node872 = (inp[12]) ? 4'b1000 : node873;
										assign node873 = (inp[0]) ? node881 : node874;
											assign node874 = (inp[2]) ? node878 : node875;
												assign node875 = (inp[14]) ? 4'b1000 : 4'b1001;
												assign node878 = (inp[7]) ? 4'b0001 : 4'b1001;
											assign node881 = (inp[14]) ? 4'b0001 : node882;
												assign node882 = (inp[2]) ? 4'b1000 : 4'b0000;
									assign node887 = (inp[0]) ? node899 : node888;
										assign node888 = (inp[13]) ? node894 : node889;
											assign node889 = (inp[7]) ? node891 : 4'b0000;
												assign node891 = (inp[12]) ? 4'b1000 : 4'b1001;
											assign node894 = (inp[12]) ? node896 : 4'b0001;
												assign node896 = (inp[2]) ? 4'b0000 : 4'b0000;
										assign node899 = (inp[11]) ? node905 : node900;
											assign node900 = (inp[14]) ? 4'b0000 : node901;
												assign node901 = (inp[1]) ? 4'b1000 : 4'b1000;
											assign node905 = (inp[1]) ? 4'b0001 : 4'b1001;
								assign node908 = (inp[13]) ? node930 : node909;
									assign node909 = (inp[2]) ? node921 : node910;
										assign node910 = (inp[11]) ? node918 : node911;
											assign node911 = (inp[0]) ? node915 : node912;
												assign node912 = (inp[7]) ? 4'b1001 : 4'b0000;
												assign node915 = (inp[14]) ? 4'b1000 : 4'b1001;
											assign node918 = (inp[0]) ? 4'b0000 : 4'b0001;
										assign node921 = (inp[1]) ? node927 : node922;
											assign node922 = (inp[11]) ? 4'b1000 : node923;
												assign node923 = (inp[10]) ? 4'b0001 : 4'b0000;
											assign node927 = (inp[7]) ? 4'b0001 : 4'b0000;
									assign node930 = (inp[10]) ? 4'b0000 : node931;
										assign node931 = (inp[1]) ? 4'b0001 : 4'b0000;
				assign node935 = (inp[0]) ? node1119 : node936;
					assign node936 = (inp[6]) ? node994 : node937;
						assign node937 = (inp[5]) ? node955 : node938;
							assign node938 = (inp[3]) ? node940 : 4'b0011;
								assign node940 = (inp[4]) ? node942 : 4'b0011;
									assign node942 = (inp[2]) ? 4'b0011 : node943;
										assign node943 = (inp[7]) ? node949 : node944;
											assign node944 = (inp[12]) ? node946 : 4'b1001;
												assign node946 = (inp[10]) ? 4'b1000 : 4'b0000;
											assign node949 = (inp[13]) ? node951 : 4'b0011;
												assign node951 = (inp[12]) ? 4'b0000 : 4'b0001;
							assign node955 = (inp[2]) ? node983 : node956;
								assign node956 = (inp[10]) ? node966 : node957;
									assign node957 = (inp[12]) ? node963 : node958;
										assign node958 = (inp[7]) ? 4'b1001 : node959;
											assign node959 = (inp[3]) ? 4'b1101 : 4'b0101;
										assign node963 = (inp[13]) ? 4'b1100 : 4'b0100;
									assign node966 = (inp[13]) ? node970 : node967;
										assign node967 = (inp[3]) ? 4'b1101 : 4'b1000;
										assign node970 = (inp[3]) ? node976 : node971;
											assign node971 = (inp[11]) ? node973 : 4'b0100;
												assign node973 = (inp[12]) ? 4'b0100 : 4'b0000;
											assign node976 = (inp[1]) ? node980 : node977;
												assign node977 = (inp[11]) ? 4'b0000 : 4'b0000;
												assign node980 = (inp[7]) ? 4'b0101 : 4'b0000;
								assign node983 = (inp[3]) ? node985 : 4'b0011;
									assign node985 = (inp[7]) ? node989 : node986;
										assign node986 = (inp[1]) ? 4'b0011 : 4'b0000;
										assign node989 = (inp[4]) ? node991 : 4'b0011;
											assign node991 = (inp[13]) ? 4'b0000 : 4'b0011;
						assign node994 = (inp[1]) ? node1068 : node995;
							assign node995 = (inp[5]) ? node1035 : node996;
								assign node996 = (inp[11]) ? node1018 : node997;
									assign node997 = (inp[14]) ? node1009 : node998;
										assign node998 = (inp[10]) ? node1006 : node999;
											assign node999 = (inp[4]) ? node1003 : node1000;
												assign node1000 = (inp[13]) ? 4'b1000 : 4'b0000;
												assign node1003 = (inp[7]) ? 4'b0000 : 4'b0100;
											assign node1006 = (inp[4]) ? 4'b1000 : 4'b0000;
										assign node1009 = (inp[13]) ? node1013 : node1010;
											assign node1010 = (inp[3]) ? 4'b0101 : 4'b0001;
											assign node1013 = (inp[3]) ? 4'b1101 : node1014;
												assign node1014 = (inp[4]) ? 4'b1000 : 4'b1001;
									assign node1018 = (inp[10]) ? node1026 : node1019;
										assign node1019 = (inp[7]) ? node1023 : node1020;
											assign node1020 = (inp[2]) ? 4'b0000 : 4'b0100;
											assign node1023 = (inp[12]) ? 4'b0100 : 4'b1100;
										assign node1026 = (inp[2]) ? 4'b1100 : node1027;
											assign node1027 = (inp[3]) ? node1031 : node1028;
												assign node1028 = (inp[13]) ? 4'b0100 : 4'b1000;
												assign node1031 = (inp[12]) ? 4'b1001 : 4'b0001;
								assign node1035 = (inp[2]) ? node1051 : node1036;
									assign node1036 = (inp[14]) ? node1044 : node1037;
										assign node1037 = (inp[11]) ? node1041 : node1038;
											assign node1038 = (inp[10]) ? 4'b0000 : 4'b0001;
											assign node1041 = (inp[4]) ? 4'b1001 : 4'b1000;
										assign node1044 = (inp[13]) ? node1046 : 4'b0000;
											assign node1046 = (inp[4]) ? 4'b0000 : node1047;
												assign node1047 = (inp[10]) ? 4'b1100 : 4'b0100;
									assign node1051 = (inp[10]) ? node1061 : node1052;
										assign node1052 = (inp[3]) ? node1056 : node1053;
											assign node1053 = (inp[11]) ? 4'b1001 : 4'b1000;
											assign node1056 = (inp[7]) ? 4'b0001 : node1057;
												assign node1057 = (inp[12]) ? 4'b1001 : 4'b0000;
										assign node1061 = (inp[4]) ? node1063 : 4'b0001;
											assign node1063 = (inp[7]) ? node1065 : 4'b1000;
												assign node1065 = (inp[11]) ? 4'b0000 : 4'b0001;
							assign node1068 = (inp[11]) ? node1096 : node1069;
								assign node1069 = (inp[13]) ? node1083 : node1070;
									assign node1070 = (inp[14]) ? node1074 : node1071;
										assign node1071 = (inp[7]) ? 4'b1000 : 4'b1001;
										assign node1074 = (inp[5]) ? node1080 : node1075;
											assign node1075 = (inp[4]) ? node1077 : 4'b0100;
												assign node1077 = (inp[10]) ? 4'b0000 : 4'b1100;
											assign node1080 = (inp[10]) ? 4'b0001 : 4'b1001;
									assign node1083 = (inp[3]) ? node1091 : node1084;
										assign node1084 = (inp[4]) ? 4'b1001 : node1085;
											assign node1085 = (inp[12]) ? 4'b0100 : node1086;
												assign node1086 = (inp[2]) ? 4'b0100 : 4'b0001;
										assign node1091 = (inp[10]) ? 4'b0000 : node1092;
											assign node1092 = (inp[4]) ? 4'b0001 : 4'b1000;
								assign node1096 = (inp[10]) ? node1106 : node1097;
									assign node1097 = (inp[2]) ? node1101 : node1098;
										assign node1098 = (inp[5]) ? 4'b0101 : 4'b1101;
										assign node1101 = (inp[4]) ? node1103 : 4'b1001;
											assign node1103 = (inp[13]) ? 4'b0101 : 4'b0001;
									assign node1106 = (inp[3]) ? node1116 : node1107;
										assign node1107 = (inp[12]) ? node1113 : node1108;
											assign node1108 = (inp[4]) ? node1110 : 4'b0101;
												assign node1110 = (inp[13]) ? 4'b0101 : 4'b1001;
											assign node1113 = (inp[13]) ? 4'b0001 : 4'b1001;
										assign node1116 = (inp[7]) ? 4'b0000 : 4'b0001;
					assign node1119 = (inp[6]) ? node1121 : 4'b0001;
						assign node1121 = (inp[2]) ? 4'b0001 : node1122;
							assign node1122 = (inp[5]) ? node1138 : node1123;
								assign node1123 = (inp[3]) ? node1125 : 4'b0001;
									assign node1125 = (inp[7]) ? node1133 : node1126;
										assign node1126 = (inp[4]) ? node1130 : node1127;
											assign node1127 = (inp[10]) ? 4'b0000 : 4'b0001;
											assign node1130 = (inp[11]) ? 4'b0000 : 4'b1000;
										assign node1133 = (inp[11]) ? node1135 : 4'b0001;
											assign node1135 = (inp[13]) ? 4'b0000 : 4'b0001;
								assign node1138 = (inp[1]) ? node1156 : node1139;
									assign node1139 = (inp[14]) ? node1151 : node1140;
										assign node1140 = (inp[13]) ? node1146 : node1141;
											assign node1141 = (inp[12]) ? 4'b0000 : node1142;
												assign node1142 = (inp[4]) ? 4'b0000 : 4'b1001;
											assign node1146 = (inp[7]) ? node1148 : 4'b0100;
												assign node1148 = (inp[4]) ? 4'b0001 : 4'b0000;
										assign node1151 = (inp[12]) ? node1153 : 4'b1000;
											assign node1153 = (inp[11]) ? 4'b0000 : 4'b1000;
									assign node1156 = (inp[11]) ? node1164 : node1157;
										assign node1157 = (inp[10]) ? node1161 : node1158;
											assign node1158 = (inp[12]) ? 4'b0000 : 4'b1000;
											assign node1161 = (inp[13]) ? 4'b0100 : 4'b0001;
										assign node1164 = (inp[13]) ? node1170 : node1165;
											assign node1165 = (inp[10]) ? 4'b1001 : node1166;
												assign node1166 = (inp[4]) ? 4'b1001 : 4'b0001;
											assign node1170 = (inp[12]) ? 4'b0001 : 4'b0101;
		assign node1174 = (inp[15]) ? node1822 : node1175;
			assign node1175 = (inp[6]) ? node1375 : node1176;
				assign node1176 = (inp[9]) ? node1272 : node1177;
					assign node1177 = (inp[0]) ? 4'b1100 : node1178;
						assign node1178 = (inp[5]) ? node1206 : node1179;
							assign node1179 = (inp[2]) ? 4'b1110 : node1180;
								assign node1180 = (inp[3]) ? node1192 : node1181;
									assign node1181 = (inp[14]) ? node1189 : node1182;
										assign node1182 = (inp[1]) ? node1186 : node1183;
											assign node1183 = (inp[4]) ? 4'b1001 : 4'b0001;
											assign node1186 = (inp[13]) ? 4'b1000 : 4'b0000;
										assign node1189 = (inp[12]) ? 4'b1110 : 4'b1000;
									assign node1192 = (inp[1]) ? 4'b0100 : node1193;
										assign node1193 = (inp[13]) ? node1199 : node1194;
											assign node1194 = (inp[14]) ? 4'b1100 : node1195;
												assign node1195 = (inp[12]) ? 4'b1001 : 4'b0001;
											assign node1199 = (inp[7]) ? node1201 : 4'b0101;
												assign node1201 = (inp[10]) ? 4'b0000 : 4'b0100;
							assign node1206 = (inp[3]) ? node1236 : node1207;
								assign node1207 = (inp[7]) ? node1225 : node1208;
									assign node1208 = (inp[1]) ? node1218 : node1209;
										assign node1209 = (inp[13]) ? node1215 : node1210;
											assign node1210 = (inp[4]) ? node1212 : 4'b1101;
												assign node1212 = (inp[11]) ? 4'b1001 : 4'b1000;
											assign node1215 = (inp[14]) ? 4'b0001 : 4'b1001;
										assign node1218 = (inp[4]) ? node1220 : 4'b0000;
											assign node1220 = (inp[12]) ? node1222 : 4'b0001;
												assign node1222 = (inp[10]) ? 4'b1000 : 4'b1000;
									assign node1225 = (inp[4]) ? node1229 : node1226;
										assign node1226 = (inp[2]) ? 4'b1110 : 4'b0100;
										assign node1229 = (inp[10]) ? node1231 : 4'b1101;
											assign node1231 = (inp[13]) ? node1233 : 4'b0000;
												assign node1233 = (inp[1]) ? 4'b1000 : 4'b1000;
								assign node1236 = (inp[1]) ? node1250 : node1237;
									assign node1237 = (inp[13]) ? node1243 : node1238;
										assign node1238 = (inp[12]) ? node1240 : 4'b0101;
											assign node1240 = (inp[2]) ? 4'b1001 : 4'b1101;
										assign node1243 = (inp[14]) ? node1247 : node1244;
											assign node1244 = (inp[7]) ? 4'b0001 : 4'b0101;
											assign node1247 = (inp[11]) ? 4'b0101 : 4'b0100;
									assign node1250 = (inp[4]) ? node1262 : node1251;
										assign node1251 = (inp[7]) ? node1257 : node1252;
											assign node1252 = (inp[10]) ? node1254 : 4'b1001;
												assign node1254 = (inp[13]) ? 4'b1101 : 4'b0100;
											assign node1257 = (inp[2]) ? node1259 : 4'b0001;
												assign node1259 = (inp[14]) ? 4'b1000 : 4'b0000;
										assign node1262 = (inp[14]) ? node1266 : node1263;
											assign node1263 = (inp[13]) ? 4'b1100 : 4'b0100;
											assign node1266 = (inp[11]) ? node1268 : 4'b1101;
												assign node1268 = (inp[2]) ? 4'b0100 : 4'b1100;
					assign node1272 = (inp[0]) ? 4'b0100 : node1273;
						assign node1273 = (inp[2]) ? node1343 : node1274;
							assign node1274 = (inp[1]) ? node1314 : node1275;
								assign node1275 = (inp[14]) ? node1293 : node1276;
									assign node1276 = (inp[13]) ? node1290 : node1277;
										assign node1277 = (inp[12]) ? node1285 : node1278;
											assign node1278 = (inp[4]) ? node1282 : node1279;
												assign node1279 = (inp[10]) ? 4'b1101 : 4'b0101;
												assign node1282 = (inp[11]) ? 4'b0001 : 4'b1001;
											assign node1285 = (inp[11]) ? node1287 : 4'b0101;
												assign node1287 = (inp[5]) ? 4'b0001 : 4'b0101;
										assign node1290 = (inp[12]) ? 4'b1101 : 4'b0101;
									assign node1293 = (inp[11]) ? node1305 : node1294;
										assign node1294 = (inp[4]) ? node1300 : node1295;
											assign node1295 = (inp[7]) ? 4'b0110 : node1296;
												assign node1296 = (inp[3]) ? 4'b0000 : 4'b0000;
											assign node1300 = (inp[7]) ? node1302 : 4'b1100;
												assign node1302 = (inp[5]) ? 4'b1100 : 4'b0110;
										assign node1305 = (inp[13]) ? 4'b1001 : node1306;
											assign node1306 = (inp[12]) ? node1310 : node1307;
												assign node1307 = (inp[3]) ? 4'b1101 : 4'b1001;
												assign node1310 = (inp[5]) ? 4'b0101 : 4'b0110;
								assign node1314 = (inp[13]) ? node1328 : node1315;
									assign node1315 = (inp[3]) ? node1325 : node1316;
										assign node1316 = (inp[5]) ? node1322 : node1317;
											assign node1317 = (inp[11]) ? node1319 : 4'b0110;
												assign node1319 = (inp[7]) ? 4'b0110 : 4'b1000;
											assign node1322 = (inp[4]) ? 4'b0100 : 4'b1100;
										assign node1325 = (inp[10]) ? 4'b1000 : 4'b0001;
									assign node1328 = (inp[12]) ? node1336 : node1329;
										assign node1329 = (inp[11]) ? node1331 : 4'b0000;
											assign node1331 = (inp[14]) ? node1333 : 4'b0100;
												assign node1333 = (inp[10]) ? 4'b0100 : 4'b0000;
										assign node1336 = (inp[14]) ? node1338 : 4'b0000;
											assign node1338 = (inp[5]) ? node1340 : 4'b1001;
												assign node1340 = (inp[4]) ? 4'b1001 : 4'b1101;
							assign node1343 = (inp[5]) ? node1345 : 4'b0110;
								assign node1345 = (inp[14]) ? node1361 : node1346;
									assign node1346 = (inp[1]) ? node1352 : node1347;
										assign node1347 = (inp[3]) ? node1349 : 4'b1001;
											assign node1349 = (inp[13]) ? 4'b0101 : 4'b0001;
										assign node1352 = (inp[13]) ? node1354 : 4'b1000;
											assign node1354 = (inp[10]) ? node1358 : node1355;
												assign node1355 = (inp[12]) ? 4'b1000 : 4'b0000;
												assign node1358 = (inp[3]) ? 4'b0100 : 4'b0000;
									assign node1361 = (inp[3]) ? node1367 : node1362;
										assign node1362 = (inp[1]) ? 4'b0110 : node1363;
											assign node1363 = (inp[11]) ? 4'b0001 : 4'b0110;
										assign node1367 = (inp[13]) ? node1369 : 4'b0001;
											assign node1369 = (inp[1]) ? node1371 : 4'b1000;
												assign node1371 = (inp[10]) ? 4'b0100 : 4'b0000;
				assign node1375 = (inp[5]) ? node1595 : node1376;
					assign node1376 = (inp[0]) ? node1526 : node1377;
						assign node1377 = (inp[11]) ? node1463 : node1378;
							assign node1378 = (inp[3]) ? node1424 : node1379;
								assign node1379 = (inp[4]) ? node1405 : node1380;
									assign node1380 = (inp[7]) ? node1392 : node1381;
										assign node1381 = (inp[2]) ? node1387 : node1382;
											assign node1382 = (inp[13]) ? node1384 : 4'b0001;
												assign node1384 = (inp[1]) ? 4'b0001 : 4'b1001;
											assign node1387 = (inp[1]) ? node1389 : 4'b0000;
												assign node1389 = (inp[14]) ? 4'b1101 : 4'b1100;
										assign node1392 = (inp[9]) ? node1398 : node1393;
											assign node1393 = (inp[13]) ? 4'b0101 : node1394;
												assign node1394 = (inp[12]) ? 4'b1100 : 4'b1101;
											assign node1398 = (inp[2]) ? node1402 : node1399;
												assign node1399 = (inp[1]) ? 4'b1100 : 4'b0100;
												assign node1402 = (inp[10]) ? 4'b1101 : 4'b0100;
									assign node1405 = (inp[9]) ? node1413 : node1406;
										assign node1406 = (inp[10]) ? node1410 : node1407;
											assign node1407 = (inp[14]) ? 4'b1101 : 4'b1001;
											assign node1410 = (inp[2]) ? 4'b0000 : 4'b0101;
										assign node1413 = (inp[10]) ? node1419 : node1414;
											assign node1414 = (inp[13]) ? node1416 : 4'b0001;
												assign node1416 = (inp[12]) ? 4'b0101 : 4'b1101;
											assign node1419 = (inp[14]) ? node1421 : 4'b1001;
												assign node1421 = (inp[12]) ? 4'b1001 : 4'b0001;
								assign node1424 = (inp[13]) ? node1450 : node1425;
									assign node1425 = (inp[4]) ? node1439 : node1426;
										assign node1426 = (inp[7]) ? node1432 : node1427;
											assign node1427 = (inp[12]) ? node1429 : 4'b0001;
												assign node1429 = (inp[10]) ? 4'b0001 : 4'b1001;
											assign node1432 = (inp[14]) ? node1436 : node1433;
												assign node1433 = (inp[1]) ? 4'b0000 : 4'b0001;
												assign node1436 = (inp[10]) ? 4'b0000 : 4'b1000;
										assign node1439 = (inp[9]) ? node1445 : node1440;
											assign node1440 = (inp[1]) ? node1442 : 4'b1001;
												assign node1442 = (inp[7]) ? 4'b0001 : 4'b1001;
											assign node1445 = (inp[12]) ? 4'b0000 : node1446;
												assign node1446 = (inp[2]) ? 4'b0001 : 4'b1001;
									assign node1450 = (inp[12]) ? node1458 : node1451;
										assign node1451 = (inp[2]) ? 4'b0101 : node1452;
											assign node1452 = (inp[14]) ? 4'b0100 : node1453;
												assign node1453 = (inp[10]) ? 4'b0000 : 4'b0001;
										assign node1458 = (inp[4]) ? node1460 : 4'b1101;
											assign node1460 = (inp[9]) ? 4'b0001 : 4'b0101;
							assign node1463 = (inp[12]) ? node1497 : node1464;
								assign node1464 = (inp[14]) ? node1482 : node1465;
									assign node1465 = (inp[1]) ? node1477 : node1466;
										assign node1466 = (inp[13]) ? node1472 : node1467;
											assign node1467 = (inp[3]) ? 4'b0001 : node1468;
												assign node1468 = (inp[9]) ? 4'b0101 : 4'b1101;
											assign node1472 = (inp[4]) ? 4'b1101 : node1473;
												assign node1473 = (inp[2]) ? 4'b1000 : 4'b0000;
										assign node1477 = (inp[9]) ? node1479 : 4'b1100;
											assign node1479 = (inp[13]) ? 4'b0000 : 4'b1000;
									assign node1482 = (inp[4]) ? node1492 : node1483;
										assign node1483 = (inp[7]) ? node1489 : node1484;
											assign node1484 = (inp[1]) ? 4'b0000 : node1485;
												assign node1485 = (inp[10]) ? 4'b0000 : 4'b0000;
											assign node1489 = (inp[13]) ? 4'b0000 : 4'b1001;
										assign node1492 = (inp[13]) ? 4'b0100 : node1493;
											assign node1493 = (inp[9]) ? 4'b0000 : 4'b1000;
								assign node1497 = (inp[9]) ? node1511 : node1498;
									assign node1498 = (inp[1]) ? node1502 : node1499;
										assign node1499 = (inp[10]) ? 4'b1001 : 4'b1000;
										assign node1502 = (inp[2]) ? node1504 : 4'b0000;
											assign node1504 = (inp[3]) ? node1508 : node1505;
												assign node1505 = (inp[4]) ? 4'b0000 : 4'b0100;
												assign node1508 = (inp[4]) ? 4'b0100 : 4'b0000;
									assign node1511 = (inp[4]) ? node1519 : node1512;
										assign node1512 = (inp[3]) ? node1514 : 4'b0100;
											assign node1514 = (inp[10]) ? 4'b1100 : node1515;
												assign node1515 = (inp[1]) ? 4'b1100 : 4'b0100;
										assign node1519 = (inp[14]) ? node1521 : 4'b1000;
											assign node1521 = (inp[1]) ? 4'b0100 : node1522;
												assign node1522 = (inp[7]) ? 4'b0000 : 4'b1100;
						assign node1526 = (inp[2]) ? node1592 : node1527;
							assign node1527 = (inp[1]) ? node1559 : node1528;
								assign node1528 = (inp[3]) ? node1542 : node1529;
									assign node1529 = (inp[9]) ? node1537 : node1530;
										assign node1530 = (inp[13]) ? 4'b0001 : node1531;
											assign node1531 = (inp[7]) ? 4'b1100 : node1532;
												assign node1532 = (inp[4]) ? 4'b1000 : 4'b1100;
										assign node1537 = (inp[11]) ? 4'b0100 : node1538;
											assign node1538 = (inp[4]) ? 4'b0001 : 4'b0100;
									assign node1542 = (inp[11]) ? node1550 : node1543;
										assign node1543 = (inp[14]) ? node1547 : node1544;
											assign node1544 = (inp[4]) ? 4'b1101 : 4'b1001;
											assign node1547 = (inp[10]) ? 4'b0100 : 4'b1100;
										assign node1550 = (inp[7]) ? node1552 : 4'b1001;
											assign node1552 = (inp[14]) ? node1556 : node1553;
												assign node1553 = (inp[12]) ? 4'b1001 : 4'b0001;
												assign node1556 = (inp[12]) ? 4'b0001 : 4'b1001;
								assign node1559 = (inp[11]) ? node1575 : node1560;
									assign node1560 = (inp[14]) ? node1570 : node1561;
										assign node1561 = (inp[9]) ? node1567 : node1562;
											assign node1562 = (inp[4]) ? 4'b1100 : node1563;
												assign node1563 = (inp[13]) ? 4'b1000 : 4'b0000;
											assign node1567 = (inp[12]) ? 4'b0000 : 4'b1000;
										assign node1570 = (inp[12]) ? node1572 : 4'b0100;
											assign node1572 = (inp[9]) ? 4'b1001 : 4'b0101;
									assign node1575 = (inp[14]) ? node1583 : node1576;
										assign node1576 = (inp[10]) ? node1578 : 4'b0000;
											assign node1578 = (inp[3]) ? 4'b0100 : node1579;
												assign node1579 = (inp[9]) ? 4'b0100 : 4'b0000;
										assign node1583 = (inp[7]) ? node1589 : node1584;
											assign node1584 = (inp[12]) ? 4'b0100 : node1585;
												assign node1585 = (inp[4]) ? 4'b0100 : 4'b1100;
											assign node1589 = (inp[12]) ? 4'b1100 : 4'b0000;
							assign node1592 = (inp[9]) ? 4'b0100 : 4'b1100;
					assign node1595 = (inp[3]) ? node1725 : node1596;
						assign node1596 = (inp[11]) ? node1664 : node1597;
							assign node1597 = (inp[7]) ? node1633 : node1598;
								assign node1598 = (inp[9]) ? node1618 : node1599;
									assign node1599 = (inp[10]) ? node1611 : node1600;
										assign node1600 = (inp[0]) ? node1606 : node1601;
											assign node1601 = (inp[2]) ? 4'b1100 : node1602;
												assign node1602 = (inp[1]) ? 4'b1000 : 4'b1000;
											assign node1606 = (inp[2]) ? node1608 : 4'b1000;
												assign node1608 = (inp[13]) ? 4'b0001 : 4'b1001;
										assign node1611 = (inp[14]) ? 4'b0001 : node1612;
											assign node1612 = (inp[13]) ? 4'b1000 : node1613;
												assign node1613 = (inp[2]) ? 4'b1001 : 4'b0001;
									assign node1618 = (inp[14]) ? node1626 : node1619;
										assign node1619 = (inp[4]) ? node1621 : 4'b0000;
											assign node1621 = (inp[12]) ? node1623 : 4'b0001;
												assign node1623 = (inp[2]) ? 4'b0000 : 4'b0001;
										assign node1626 = (inp[12]) ? node1630 : node1627;
											assign node1627 = (inp[13]) ? 4'b0100 : 4'b0000;
											assign node1630 = (inp[4]) ? 4'b0001 : 4'b0101;
								assign node1633 = (inp[12]) ? node1651 : node1634;
									assign node1634 = (inp[0]) ? node1642 : node1635;
										assign node1635 = (inp[13]) ? node1639 : node1636;
											assign node1636 = (inp[10]) ? 4'b0000 : 4'b0100;
											assign node1639 = (inp[2]) ? 4'b1001 : 4'b1000;
										assign node1642 = (inp[1]) ? node1648 : node1643;
											assign node1643 = (inp[13]) ? 4'b1100 : node1644;
												assign node1644 = (inp[9]) ? 4'b1001 : 4'b1101;
											assign node1648 = (inp[9]) ? 4'b0100 : 4'b1100;
									assign node1651 = (inp[4]) ? node1657 : node1652;
										assign node1652 = (inp[9]) ? node1654 : 4'b1101;
											assign node1654 = (inp[14]) ? 4'b1101 : 4'b0101;
										assign node1657 = (inp[14]) ? 4'b1001 : node1658;
											assign node1658 = (inp[10]) ? node1660 : 4'b1100;
												assign node1660 = (inp[2]) ? 4'b0000 : 4'b0001;
							assign node1664 = (inp[1]) ? node1694 : node1665;
								assign node1665 = (inp[4]) ? node1677 : node1666;
									assign node1666 = (inp[13]) ? node1670 : node1667;
										assign node1667 = (inp[14]) ? 4'b0100 : 4'b1100;
										assign node1670 = (inp[10]) ? node1672 : 4'b0100;
											assign node1672 = (inp[2]) ? node1674 : 4'b1000;
												assign node1674 = (inp[14]) ? 4'b1001 : 4'b0001;
									assign node1677 = (inp[0]) ? node1685 : node1678;
										assign node1678 = (inp[9]) ? 4'b1000 : node1679;
											assign node1679 = (inp[12]) ? 4'b0001 : node1680;
												assign node1680 = (inp[10]) ? 4'b0000 : 4'b0000;
										assign node1685 = (inp[2]) ? node1691 : node1686;
											assign node1686 = (inp[7]) ? 4'b1000 : node1687;
												assign node1687 = (inp[12]) ? 4'b0100 : 4'b1100;
											assign node1691 = (inp[7]) ? 4'b0001 : 4'b1001;
								assign node1694 = (inp[9]) ? node1708 : node1695;
									assign node1695 = (inp[7]) ? 4'b1100 : node1696;
										assign node1696 = (inp[13]) ? node1702 : node1697;
											assign node1697 = (inp[0]) ? 4'b0000 : node1698;
												assign node1698 = (inp[10]) ? 4'b0000 : 4'b1000;
											assign node1702 = (inp[12]) ? node1704 : 4'b1000;
												assign node1704 = (inp[4]) ? 4'b1000 : 4'b1100;
									assign node1708 = (inp[10]) ? node1714 : node1709;
										assign node1709 = (inp[4]) ? node1711 : 4'b1000;
											assign node1711 = (inp[14]) ? 4'b1000 : 4'b0000;
										assign node1714 = (inp[2]) ? node1720 : node1715;
											assign node1715 = (inp[0]) ? node1717 : 4'b0000;
												assign node1717 = (inp[14]) ? 4'b0100 : 4'b0000;
											assign node1720 = (inp[7]) ? 4'b0100 : node1721;
												assign node1721 = (inp[0]) ? 4'b0100 : 4'b1000;
						assign node1725 = (inp[11]) ? node1777 : node1726;
							assign node1726 = (inp[4]) ? node1754 : node1727;
								assign node1727 = (inp[2]) ? node1743 : node1728;
									assign node1728 = (inp[1]) ? node1734 : node1729;
										assign node1729 = (inp[14]) ? node1731 : 4'b1001;
											assign node1731 = (inp[10]) ? 4'b0000 : 4'b0001;
										assign node1734 = (inp[12]) ? node1738 : node1735;
											assign node1735 = (inp[14]) ? 4'b1000 : 4'b0000;
											assign node1738 = (inp[9]) ? 4'b0001 : node1739;
												assign node1739 = (inp[14]) ? 4'b0000 : 4'b0000;
									assign node1743 = (inp[9]) ? node1751 : node1744;
										assign node1744 = (inp[0]) ? node1746 : 4'b1001;
											assign node1746 = (inp[10]) ? 4'b0001 : node1747;
												assign node1747 = (inp[7]) ? 4'b0001 : 4'b1001;
										assign node1751 = (inp[12]) ? 4'b0000 : 4'b0001;
								assign node1754 = (inp[7]) ? node1768 : node1755;
									assign node1755 = (inp[1]) ? node1757 : 4'b0000;
										assign node1757 = (inp[0]) ? node1763 : node1758;
											assign node1758 = (inp[12]) ? 4'b0000 : node1759;
												assign node1759 = (inp[2]) ? 4'b0000 : 4'b0001;
											assign node1763 = (inp[13]) ? node1765 : 4'b0001;
												assign node1765 = (inp[2]) ? 4'b0001 : 4'b0000;
									assign node1768 = (inp[10]) ? node1772 : node1769;
										assign node1769 = (inp[12]) ? 4'b1000 : 4'b1001;
										assign node1772 = (inp[14]) ? 4'b0000 : node1773;
											assign node1773 = (inp[13]) ? 4'b0000 : 4'b1000;
							assign node1777 = (inp[13]) ? node1809 : node1778;
								assign node1778 = (inp[1]) ? node1790 : node1779;
									assign node1779 = (inp[10]) ? node1787 : node1780;
										assign node1780 = (inp[9]) ? node1784 : node1781;
											assign node1781 = (inp[14]) ? 4'b1000 : 4'b0000;
											assign node1784 = (inp[4]) ? 4'b0001 : 4'b1001;
										assign node1787 = (inp[0]) ? 4'b0001 : 4'b1001;
									assign node1790 = (inp[10]) ? node1802 : node1791;
										assign node1791 = (inp[12]) ? node1797 : node1792;
											assign node1792 = (inp[4]) ? node1794 : 4'b0000;
												assign node1794 = (inp[2]) ? 4'b1000 : 4'b0000;
											assign node1797 = (inp[0]) ? 4'b1000 : node1798;
												assign node1798 = (inp[2]) ? 4'b0000 : 4'b1000;
										assign node1802 = (inp[2]) ? 4'b0000 : node1803;
											assign node1803 = (inp[4]) ? 4'b0000 : node1804;
												assign node1804 = (inp[9]) ? 4'b0000 : 4'b1000;
								assign node1809 = (inp[12]) ? node1811 : 4'b0000;
									assign node1811 = (inp[4]) ? node1817 : node1812;
										assign node1812 = (inp[0]) ? 4'b0000 : node1813;
											assign node1813 = (inp[9]) ? 4'b0001 : 4'b1001;
										assign node1817 = (inp[7]) ? 4'b0000 : node1818;
											assign node1818 = (inp[1]) ? 4'b0000 : 4'b0001;
			assign node1822 = (inp[9]) ? node2094 : node1823;
				assign node1823 = (inp[6]) ? node1891 : node1824;
					assign node1824 = (inp[0]) ? 4'b1000 : node1825;
						assign node1825 = (inp[5]) ? node1839 : node1826;
							assign node1826 = (inp[3]) ? node1828 : 4'b1010;
								assign node1828 = (inp[2]) ? 4'b1010 : node1829;
									assign node1829 = (inp[7]) ? 4'b1010 : node1830;
										assign node1830 = (inp[1]) ? 4'b0000 : node1831;
											assign node1831 = (inp[11]) ? 4'b1010 : node1832;
												assign node1832 = (inp[13]) ? 4'b0000 : 4'b1000;
							assign node1839 = (inp[2]) ? node1873 : node1840;
								assign node1840 = (inp[1]) ? node1860 : node1841;
									assign node1841 = (inp[11]) ? node1853 : node1842;
										assign node1842 = (inp[14]) ? node1850 : node1843;
											assign node1843 = (inp[13]) ? node1847 : node1844;
												assign node1844 = (inp[10]) ? 4'b0101 : 4'b1001;
												assign node1847 = (inp[7]) ? 4'b0001 : 4'b0001;
											assign node1850 = (inp[12]) ? 4'b0000 : 4'b1000;
										assign node1853 = (inp[10]) ? node1857 : node1854;
											assign node1854 = (inp[3]) ? 4'b1101 : 4'b1001;
											assign node1857 = (inp[7]) ? 4'b0101 : 4'b1101;
									assign node1860 = (inp[11]) ? node1868 : node1861;
										assign node1861 = (inp[14]) ? 4'b1101 : node1862;
											assign node1862 = (inp[4]) ? 4'b1100 : node1863;
												assign node1863 = (inp[3]) ? 4'b1100 : 4'b0100;
										assign node1868 = (inp[3]) ? 4'b0000 : node1869;
											assign node1869 = (inp[14]) ? 4'b1100 : 4'b1000;
								assign node1873 = (inp[3]) ? node1875 : 4'b1010;
									assign node1875 = (inp[1]) ? node1883 : node1876;
										assign node1876 = (inp[12]) ? node1880 : node1877;
											assign node1877 = (inp[10]) ? 4'b1001 : 4'b0001;
											assign node1880 = (inp[7]) ? 4'b0001 : 4'b0000;
										assign node1883 = (inp[7]) ? node1885 : 4'b0000;
											assign node1885 = (inp[4]) ? node1887 : 4'b1010;
												assign node1887 = (inp[14]) ? 4'b0000 : 4'b0000;
					assign node1891 = (inp[0]) ? node2023 : node1892;
						assign node1892 = (inp[5]) ? node1974 : node1893;
							assign node1893 = (inp[11]) ? node1941 : node1894;
								assign node1894 = (inp[13]) ? node1918 : node1895;
									assign node1895 = (inp[4]) ? node1905 : node1896;
										assign node1896 = (inp[7]) ? node1898 : 4'b0100;
											assign node1898 = (inp[3]) ? node1902 : node1899;
												assign node1899 = (inp[1]) ? 4'b0000 : 4'b1001;
												assign node1902 = (inp[1]) ? 4'b0101 : 4'b0001;
										assign node1905 = (inp[2]) ? node1911 : node1906;
											assign node1906 = (inp[10]) ? node1908 : 4'b1101;
												assign node1908 = (inp[14]) ? 4'b1000 : 4'b1001;
											assign node1911 = (inp[10]) ? node1915 : node1912;
												assign node1912 = (inp[7]) ? 4'b1101 : 4'b1000;
												assign node1915 = (inp[1]) ? 4'b0100 : 4'b0101;
									assign node1918 = (inp[12]) ? node1928 : node1919;
										assign node1919 = (inp[14]) ? node1925 : node1920;
											assign node1920 = (inp[2]) ? node1922 : 4'b1001;
												assign node1922 = (inp[1]) ? 4'b0001 : 4'b1001;
											assign node1925 = (inp[2]) ? 4'b1001 : 4'b1000;
										assign node1928 = (inp[2]) ? node1934 : node1929;
											assign node1929 = (inp[10]) ? node1931 : 4'b1001;
												assign node1931 = (inp[3]) ? 4'b0101 : 4'b0001;
											assign node1934 = (inp[4]) ? node1938 : node1935;
												assign node1935 = (inp[3]) ? 4'b0101 : 4'b0000;
												assign node1938 = (inp[3]) ? 4'b0001 : 4'b0101;
								assign node1941 = (inp[1]) ? node1959 : node1942;
									assign node1942 = (inp[3]) ? node1954 : node1943;
										assign node1943 = (inp[2]) ? node1947 : node1944;
											assign node1944 = (inp[4]) ? 4'b0000 : 4'b0101;
											assign node1947 = (inp[7]) ? node1951 : node1948;
												assign node1948 = (inp[13]) ? 4'b0101 : 4'b0101;
												assign node1951 = (inp[13]) ? 4'b0001 : 4'b1001;
										assign node1954 = (inp[7]) ? node1956 : 4'b0001;
											assign node1956 = (inp[2]) ? 4'b1101 : 4'b1100;
									assign node1959 = (inp[10]) ? node1969 : node1960;
										assign node1960 = (inp[14]) ? node1962 : 4'b0000;
											assign node1962 = (inp[2]) ? node1966 : node1963;
												assign node1963 = (inp[13]) ? 4'b0000 : 4'b0100;
												assign node1966 = (inp[12]) ? 4'b1100 : 4'b0000;
										assign node1969 = (inp[3]) ? 4'b1000 : node1970;
											assign node1970 = (inp[2]) ? 4'b1100 : 4'b1000;
							assign node1974 = (inp[3]) ? node2004 : node1975;
								assign node1975 = (inp[4]) ? node1995 : node1976;
									assign node1976 = (inp[2]) ? node1988 : node1977;
										assign node1977 = (inp[1]) ? node1981 : node1978;
											assign node1978 = (inp[11]) ? 4'b1001 : 4'b1000;
											assign node1981 = (inp[11]) ? node1985 : node1982;
												assign node1982 = (inp[12]) ? 4'b1100 : 4'b0101;
												assign node1985 = (inp[14]) ? 4'b0100 : 4'b1000;
										assign node1988 = (inp[11]) ? 4'b0100 : node1989;
											assign node1989 = (inp[13]) ? 4'b0101 : node1990;
												assign node1990 = (inp[1]) ? 4'b0001 : 4'b0101;
									assign node1995 = (inp[13]) ? 4'b1000 : node1996;
										assign node1996 = (inp[1]) ? node1998 : 4'b0100;
											assign node1998 = (inp[10]) ? 4'b0000 : node1999;
												assign node1999 = (inp[2]) ? 4'b1000 : 4'b0000;
								assign node2004 = (inp[14]) ? node2012 : node2005;
									assign node2005 = (inp[10]) ? node2009 : node2006;
										assign node2006 = (inp[1]) ? 4'b1001 : 4'b0001;
										assign node2009 = (inp[11]) ? 4'b1000 : 4'b0000;
									assign node2012 = (inp[4]) ? node2016 : node2013;
										assign node2013 = (inp[2]) ? 4'b1000 : 4'b0000;
										assign node2016 = (inp[1]) ? 4'b0000 : node2017;
											assign node2017 = (inp[12]) ? 4'b0000 : node2018;
												assign node2018 = (inp[7]) ? 4'b0000 : 4'b0001;
						assign node2023 = (inp[5]) ? node2041 : node2024;
							assign node2024 = (inp[3]) ? node2026 : 4'b1000;
								assign node2026 = (inp[2]) ? 4'b1000 : node2027;
									assign node2027 = (inp[7]) ? node2033 : node2028;
										assign node2028 = (inp[11]) ? node2030 : 4'b0001;
											assign node2030 = (inp[4]) ? 4'b1001 : 4'b1000;
										assign node2033 = (inp[13]) ? 4'b1000 : node2034;
											assign node2034 = (inp[10]) ? node2036 : 4'b1000;
												assign node2036 = (inp[11]) ? 4'b0001 : 4'b0000;
							assign node2041 = (inp[2]) ? node2079 : node2042;
								assign node2042 = (inp[3]) ? node2066 : node2043;
									assign node2043 = (inp[7]) ? node2055 : node2044;
										assign node2044 = (inp[4]) ? node2052 : node2045;
											assign node2045 = (inp[12]) ? node2049 : node2046;
												assign node2046 = (inp[11]) ? 4'b0100 : 4'b0101;
												assign node2049 = (inp[1]) ? 4'b1000 : 4'b0101;
											assign node2052 = (inp[1]) ? 4'b1000 : 4'b1100;
										assign node2055 = (inp[1]) ? node2063 : node2056;
											assign node2056 = (inp[11]) ? node2060 : node2057;
												assign node2057 = (inp[12]) ? 4'b1001 : 4'b1000;
												assign node2060 = (inp[12]) ? 4'b0001 : 4'b1001;
											assign node2063 = (inp[14]) ? 4'b0001 : 4'b0000;
									assign node2066 = (inp[1]) ? node2072 : node2067;
										assign node2067 = (inp[7]) ? 4'b0000 : node2068;
											assign node2068 = (inp[14]) ? 4'b0001 : 4'b0000;
										assign node2072 = (inp[12]) ? node2076 : node2073;
											assign node2073 = (inp[7]) ? 4'b1001 : 4'b0001;
											assign node2076 = (inp[14]) ? 4'b0000 : 4'b0001;
								assign node2079 = (inp[3]) ? node2081 : 4'b1000;
									assign node2081 = (inp[7]) ? node2089 : node2082;
										assign node2082 = (inp[4]) ? 4'b0000 : node2083;
											assign node2083 = (inp[10]) ? 4'b0000 : node2084;
												assign node2084 = (inp[14]) ? 4'b0000 : 4'b1000;
										assign node2089 = (inp[4]) ? node2091 : 4'b1000;
											assign node2091 = (inp[14]) ? 4'b1000 : 4'b0001;
				assign node2094 = (inp[0]) ? node2260 : node2095;
					assign node2095 = (inp[6]) ? node2157 : node2096;
						assign node2096 = (inp[2]) ? node2146 : node2097;
							assign node2097 = (inp[5]) ? node2107 : node2098;
								assign node2098 = (inp[3]) ? node2100 : 4'b0010;
									assign node2100 = (inp[4]) ? 4'b0001 : node2101;
										assign node2101 = (inp[12]) ? node2103 : 4'b0010;
											assign node2103 = (inp[14]) ? 4'b0000 : 4'b0010;
								assign node2107 = (inp[1]) ? node2131 : node2108;
									assign node2108 = (inp[13]) ? node2118 : node2109;
										assign node2109 = (inp[3]) ? node2113 : node2110;
											assign node2110 = (inp[10]) ? 4'b1001 : 4'b0001;
											assign node2113 = (inp[12]) ? 4'b0001 : node2114;
												assign node2114 = (inp[14]) ? 4'b0100 : 4'b0101;
										assign node2118 = (inp[11]) ? node2126 : node2119;
											assign node2119 = (inp[14]) ? node2123 : node2120;
												assign node2120 = (inp[3]) ? 4'b1101 : 4'b1001;
												assign node2123 = (inp[10]) ? 4'b1000 : 4'b1100;
											assign node2126 = (inp[10]) ? 4'b0101 : node2127;
												assign node2127 = (inp[12]) ? 4'b1101 : 4'b1001;
									assign node2131 = (inp[10]) ? node2139 : node2132;
										assign node2132 = (inp[3]) ? node2134 : 4'b0000;
											assign node2134 = (inp[11]) ? node2136 : 4'b1100;
												assign node2136 = (inp[7]) ? 4'b0100 : 4'b0000;
										assign node2139 = (inp[13]) ? node2143 : node2140;
											assign node2140 = (inp[3]) ? 4'b1001 : 4'b1000;
											assign node2143 = (inp[7]) ? 4'b0001 : 4'b0100;
							assign node2146 = (inp[3]) ? node2148 : 4'b0010;
								assign node2148 = (inp[7]) ? 4'b0010 : node2149;
									assign node2149 = (inp[4]) ? node2151 : 4'b0010;
										assign node2151 = (inp[5]) ? node2153 : 4'b0010;
											assign node2153 = (inp[11]) ? 4'b1001 : 4'b0000;
						assign node2157 = (inp[11]) ? node2215 : node2158;
							assign node2158 = (inp[5]) ? node2192 : node2159;
								assign node2159 = (inp[3]) ? node2179 : node2160;
									assign node2160 = (inp[7]) ? node2166 : node2161;
										assign node2161 = (inp[4]) ? node2163 : 4'b1001;
											assign node2163 = (inp[10]) ? 4'b0100 : 4'b0101;
										assign node2166 = (inp[2]) ? node2172 : node2167;
											assign node2167 = (inp[4]) ? node2169 : 4'b0000;
												assign node2169 = (inp[10]) ? 4'b0001 : 4'b0001;
											assign node2172 = (inp[4]) ? node2176 : node2173;
												assign node2173 = (inp[13]) ? 4'b1001 : 4'b0001;
												assign node2176 = (inp[14]) ? 4'b0000 : 4'b1000;
									assign node2179 = (inp[4]) ? node2183 : node2180;
										assign node2180 = (inp[14]) ? 4'b1100 : 4'b1101;
										assign node2183 = (inp[7]) ? node2189 : node2184;
											assign node2184 = (inp[13]) ? node2186 : 4'b0001;
												assign node2186 = (inp[1]) ? 4'b1001 : 4'b0001;
											assign node2189 = (inp[14]) ? 4'b1101 : 4'b0101;
								assign node2192 = (inp[1]) ? node2204 : node2193;
									assign node2193 = (inp[10]) ? node2201 : node2194;
										assign node2194 = (inp[4]) ? 4'b0001 : node2195;
											assign node2195 = (inp[14]) ? node2197 : 4'b0000;
												assign node2197 = (inp[2]) ? 4'b0101 : 4'b1000;
										assign node2201 = (inp[3]) ? 4'b0000 : 4'b1000;
									assign node2204 = (inp[3]) ? node2208 : node2205;
										assign node2205 = (inp[2]) ? 4'b1001 : 4'b0001;
										assign node2208 = (inp[13]) ? 4'b1000 : node2209;
											assign node2209 = (inp[14]) ? node2211 : 4'b0001;
												assign node2211 = (inp[4]) ? 4'b0000 : 4'b0001;
							assign node2215 = (inp[13]) ? node2241 : node2216;
								assign node2216 = (inp[1]) ? node2230 : node2217;
									assign node2217 = (inp[5]) ? node2223 : node2218;
										assign node2218 = (inp[7]) ? 4'b0101 : node2219;
											assign node2219 = (inp[10]) ? 4'b1001 : 4'b0001;
										assign node2223 = (inp[10]) ? node2227 : node2224;
											assign node2224 = (inp[2]) ? 4'b1100 : 4'b1000;
											assign node2227 = (inp[4]) ? 4'b0001 : 4'b0100;
									assign node2230 = (inp[10]) ? node2238 : node2231;
										assign node2231 = (inp[4]) ? node2233 : 4'b0100;
											assign node2233 = (inp[7]) ? 4'b0000 : node2234;
												assign node2234 = (inp[3]) ? 4'b0000 : 4'b0100;
										assign node2238 = (inp[4]) ? 4'b1100 : 4'b1000;
								assign node2241 = (inp[10]) ? node2255 : node2242;
									assign node2242 = (inp[2]) ? 4'b1000 : node2243;
										assign node2243 = (inp[3]) ? node2247 : node2244;
											assign node2244 = (inp[7]) ? 4'b0000 : 4'b0101;
											assign node2247 = (inp[12]) ? node2251 : node2248;
												assign node2248 = (inp[5]) ? 4'b0000 : 4'b1000;
												assign node2251 = (inp[4]) ? 4'b0000 : 4'b1100;
									assign node2255 = (inp[3]) ? 4'b0000 : node2256;
										assign node2256 = (inp[12]) ? 4'b0000 : 4'b1000;
					assign node2260 = (inp[6]) ? node2262 : 4'b0000;
						assign node2262 = (inp[2]) ? node2308 : node2263;
							assign node2263 = (inp[5]) ? node2273 : node2264;
								assign node2264 = (inp[7]) ? 4'b0000 : node2265;
									assign node2265 = (inp[14]) ? node2267 : 4'b0000;
										assign node2267 = (inp[4]) ? node2269 : 4'b0001;
											assign node2269 = (inp[1]) ? 4'b0000 : 4'b1000;
								assign node2273 = (inp[1]) ? node2287 : node2274;
									assign node2274 = (inp[4]) ? node2282 : node2275;
										assign node2275 = (inp[7]) ? node2279 : node2276;
											assign node2276 = (inp[13]) ? 4'b0101 : 4'b0001;
											assign node2279 = (inp[14]) ? 4'b1001 : 4'b0001;
										assign node2282 = (inp[12]) ? 4'b1001 : node2283;
											assign node2283 = (inp[3]) ? 4'b1000 : 4'b1100;
									assign node2287 = (inp[14]) ? node2299 : node2288;
										assign node2288 = (inp[4]) ? node2294 : node2289;
											assign node2289 = (inp[10]) ? 4'b1000 : node2290;
												assign node2290 = (inp[11]) ? 4'b0000 : 4'b1000;
											assign node2294 = (inp[13]) ? node2296 : 4'b1100;
												assign node2296 = (inp[11]) ? 4'b0000 : 4'b0100;
										assign node2299 = (inp[11]) ? node2303 : node2300;
											assign node2300 = (inp[3]) ? 4'b0001 : 4'b1001;
											assign node2303 = (inp[4]) ? 4'b0000 : node2304;
												assign node2304 = (inp[7]) ? 4'b0000 : 4'b1000;
							assign node2308 = (inp[10]) ? 4'b0000 : node2309;
								assign node2309 = (inp[5]) ? node2311 : 4'b0000;
									assign node2311 = (inp[7]) ? 4'b0000 : node2312;
										assign node2312 = (inp[3]) ? 4'b0001 : 4'b0000;

endmodule