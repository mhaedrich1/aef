module dtc_split75_bm37 (
	input  wire [8-1:0] inp,
	output wire [63-1:0] outp
);

	wire [63-1:0] node1;
	wire [63-1:0] node2;
	wire [63-1:0] node3;
	wire [63-1:0] node4;
	wire [63-1:0] node5;
	wire [63-1:0] node7;
	wire [63-1:0] node10;
	wire [63-1:0] node12;
	wire [63-1:0] node14;
	wire [63-1:0] node17;
	wire [63-1:0] node18;
	wire [63-1:0] node19;
	wire [63-1:0] node20;
	wire [63-1:0] node24;
	wire [63-1:0] node27;
	wire [63-1:0] node28;
	wire [63-1:0] node29;
	wire [63-1:0] node33;
	wire [63-1:0] node35;
	wire [63-1:0] node38;
	wire [63-1:0] node39;
	wire [63-1:0] node40;
	wire [63-1:0] node42;
	wire [63-1:0] node46;
	wire [63-1:0] node47;
	wire [63-1:0] node48;
	wire [63-1:0] node49;
	wire [63-1:0] node52;
	wire [63-1:0] node56;
	wire [63-1:0] node57;
	wire [63-1:0] node58;
	wire [63-1:0] node62;
	wire [63-1:0] node63;
	wire [63-1:0] node67;
	wire [63-1:0] node68;
	wire [63-1:0] node69;
	wire [63-1:0] node70;
	wire [63-1:0] node72;
	wire [63-1:0] node76;
	wire [63-1:0] node77;
	wire [63-1:0] node79;
	wire [63-1:0] node81;
	wire [63-1:0] node84;
	wire [63-1:0] node86;
	wire [63-1:0] node88;
	wire [63-1:0] node91;
	wire [63-1:0] node92;
	wire [63-1:0] node93;
	wire [63-1:0] node94;
	wire [63-1:0] node97;
	wire [63-1:0] node99;
	wire [63-1:0] node102;
	wire [63-1:0] node104;
	wire [63-1:0] node106;
	wire [63-1:0] node109;
	wire [63-1:0] node110;
	wire [63-1:0] node112;
	wire [63-1:0] node115;
	wire [63-1:0] node116;
	wire [63-1:0] node117;
	wire [63-1:0] node121;
	wire [63-1:0] node124;
	wire [63-1:0] node125;
	wire [63-1:0] node126;
	wire [63-1:0] node127;
	wire [63-1:0] node129;
	wire [63-1:0] node131;
	wire [63-1:0] node134;
	wire [63-1:0] node135;
	wire [63-1:0] node137;
	wire [63-1:0] node140;
	wire [63-1:0] node143;
	wire [63-1:0] node144;
	wire [63-1:0] node145;
	wire [63-1:0] node148;
	wire [63-1:0] node150;
	wire [63-1:0] node153;
	wire [63-1:0] node154;
	wire [63-1:0] node156;
	wire [63-1:0] node158;
	wire [63-1:0] node161;
	wire [63-1:0] node163;
	wire [63-1:0] node165;
	wire [63-1:0] node168;
	wire [63-1:0] node169;
	wire [63-1:0] node170;
	wire [63-1:0] node171;
	wire [63-1:0] node172;
	wire [63-1:0] node174;
	wire [63-1:0] node177;
	wire [63-1:0] node178;
	wire [63-1:0] node182;
	wire [63-1:0] node183;
	wire [63-1:0] node185;
	wire [63-1:0] node188;
	wire [63-1:0] node189;
	wire [63-1:0] node192;
	wire [63-1:0] node195;
	wire [63-1:0] node196;
	wire [63-1:0] node197;
	wire [63-1:0] node201;
	wire [63-1:0] node203;
	wire [63-1:0] node206;
	wire [63-1:0] node207;
	wire [63-1:0] node209;
	wire [63-1:0] node211;
	wire [63-1:0] node214;
	wire [63-1:0] node215;
	wire [63-1:0] node216;
	wire [63-1:0] node218;
	wire [63-1:0] node221;
	wire [63-1:0] node224;
	wire [63-1:0] node225;
	wire [63-1:0] node227;
	wire [63-1:0] node230;
	wire [63-1:0] node231;
	wire [63-1:0] node234;

	assign outp = (inp[7]) ? node124 : node1;
		assign node1 = (inp[6]) ? node67 : node2;
			assign node2 = (inp[1]) ? node38 : node3;
				assign node3 = (inp[2]) ? node17 : node4;
					assign node4 = (inp[3]) ? node10 : node5;
						assign node5 = (inp[5]) ? node7 : 63'b100111101001100000110001101110110010010101001100001101001010101;
							assign node7 = (inp[0]) ? 63'b100111101001100000110001101110110010010101001101001101001010101 : 63'b100111101001100000110001101110110010010101001100001101001010101;
						assign node10 = (inp[0]) ? node12 : 63'b100110101001100000110001101110110011010101001100000101001010101;
							assign node12 = (inp[5]) ? node14 : 63'b100110101001100000110001101110110011010101001100000101001010101;
								assign node14 = (inp[4]) ? 63'b100110101001100000110001101110110011010101001101000101001010101 : 63'b100110101001100000110001101110110011010101001100000101001010101;
					assign node17 = (inp[4]) ? node27 : node18;
						assign node18 = (inp[0]) ? node24 : node19;
							assign node19 = (inp[5]) ? 63'b100111101001100100110001101110110011010101001100101101001010101 : node20;
								assign node20 = (inp[3]) ? 63'b100111101001100000110001101110110011010101001100101101001010111 : 63'b100110100001100000110001101110110001010101000100001101001010101;
							assign node24 = (inp[5]) ? 63'b100111101001000000110001101110110011000110001100101001001010101 : 63'b100111101001100000110001101110110011010101001100101101001010101;
						assign node27 = (inp[0]) ? node33 : node28;
							assign node28 = (inp[3]) ? 63'b100111001001100000110001101110110011010101001100100101001000101 : node29;
								assign node29 = (inp[5]) ? 63'b100101101001110000110001101110110011010101001100101101001010101 : 63'b100111101001100000110001101110110011010101001100101101001010101;
							assign node33 = (inp[3]) ? node35 : 63'b100111101001100000110001101110110010010101011100001101001010101;
								assign node35 = (inp[5]) ? 63'b100110101001100000110001101110110011010101011101000101001010101 : 63'b100110101001100000110001101110110011010101011100000101001010101;
				assign node38 = (inp[2]) ? node46 : node39;
					assign node39 = (inp[3]) ? 63'b100001101001100000010001101110010010010101001100101101000010101 : node40;
						assign node40 = (inp[5]) ? node42 : 63'b100111101001100000010001101110010010010101001100101101000000101;
							assign node42 = (inp[4]) ? 63'b100111101001100000010001101110010010010101001101101101000000101 : 63'b100111101001100000010001101110010010010101001100101101000000101;
					assign node46 = (inp[3]) ? node56 : node47;
						assign node47 = (inp[0]) ? 63'b100111101001100000110001101110010010010101011100101101000000101 : node48;
							assign node48 = (inp[5]) ? node52 : node49;
								assign node49 = (inp[4]) ? 63'b110111100001000000110001101100110011010101001100111101001010101 : 63'b101110100001100000110001101110110011010101001100101101001010100;
								assign node52 = (inp[4]) ? 63'b100111101001100000110001101110110011010101001100101101001010101 : 63'b100111101001100100110001101110110011010101001100101101001010101;
						assign node56 = (inp[0]) ? node62 : node57;
							assign node57 = (inp[4]) ? 63'b100001101001100000110001101110110011010101001100101101001010101 : node58;
								assign node58 = (inp[5]) ? 63'b100001101001100100110001101110110011010101001100101101001010101 : 63'b100001111001100000110001101110110010010101001100101101001010100;
							assign node62 = (inp[4]) ? 63'b100001101001100000110001101110010010010101011101101101000010101 : node63;
								assign node63 = (inp[5]) ? 63'b100001101001000000110001101110110011010100001100101101001110101 : 63'b100001101001100000110001101110110011010101001100101101001010101;
			assign node67 = (inp[2]) ? node91 : node68;
				assign node68 = (inp[3]) ? node76 : node69;
					assign node69 = (inp[1]) ? 63'b100110101001100000110001101110110011010101000100001101001010001 : node70;
						assign node70 = (inp[0]) ? node72 : 63'b100110101001100000110001101110110001010101000100101101001010000;
							assign node72 = (inp[4]) ? 63'b100110101001100000110001101110110001010101000101101101001010000 : 63'b100110101001100000110001101110110001010101000100101101001010000;
					assign node76 = (inp[1]) ? node84 : node77;
						assign node77 = (inp[4]) ? node79 : 63'b100110101001100000110001101110110011010001001100001101001010101;
							assign node79 = (inp[5]) ? node81 : 63'b100110101001100000110001101110110011010001001100001101001010101;
								assign node81 = (inp[0]) ? 63'b100110101001100000110001101110110011010001001101001101001010101 : 63'b100110101001100000110001101110110011010001001100001101001010101;
						assign node84 = (inp[5]) ? node86 : 63'b100110101001100000110001101110100011010101001100100101001010100;
							assign node86 = (inp[0]) ? node88 : 63'b100110101001100000110001101110100011010101001100100101001010100;
								assign node88 = (inp[4]) ? 63'b100110101001100000110001101110100011010101001101100101001010100 : 63'b100110101001100000110001101110100011010101001100100101001010100;
				assign node91 = (inp[0]) ? node109 : node92;
					assign node92 = (inp[5]) ? node102 : node93;
						assign node93 = (inp[4]) ? node97 : node94;
							assign node94 = (inp[3]) ? 63'b100111101001100000110011101110110011010101001100001101001010101 : 63'b100111101001100000111001101110110011010001001100100101001010100;
							assign node97 = (inp[3]) ? node99 : 63'b100111101001100000110001101110110011010101001100101101001010101;
								assign node99 = (inp[1]) ? 63'b100111001001100000110001101110100011010101001100100101001000101 : 63'b100111001001100000110001101110110011010001001100101101001000101;
						assign node102 = (inp[4]) ? node104 : 63'b100111101001100100110001101110110011010101001100101101001010101;
							assign node104 = (inp[1]) ? node106 : 63'b100101101001110000110001101110110011010101001100101101001010101;
								assign node106 = (inp[3]) ? 63'b100111101001100000110101101110110011010101001100101101001010101 : 63'b100111101001100001110001101110110011010101001100101101001010101;
					assign node109 = (inp[4]) ? node115 : node110;
						assign node110 = (inp[5]) ? node112 : 63'b100111101001100000110001101110110011010101001100101101001010101;
							assign node112 = (inp[1]) ? 63'b100111101001000000110001101110110011010100001100101101001110101 : 63'b100111101001000000110001101110110011000110001100101001001010101;
						assign node115 = (inp[3]) ? node121 : node116;
							assign node116 = (inp[1]) ? 63'b100110101001100000110001101110110011010101010101001101001010001 : node117;
								assign node117 = (inp[5]) ? 63'b100110101001100000110001101110110001010101010101101101001010000 : 63'b100110101001100000110001101110110001010101010100101101001010000;
							assign node121 = (inp[1]) ? 63'b100110101001100000110001101110100011010101011101100101001010100 : 63'b100110101001100000110001101110110011010001011101001101001010101;
		assign node124 = (inp[2]) ? node168 : node125;
			assign node125 = (inp[3]) ? node143 : node126;
				assign node126 = (inp[1]) ? node134 : node127;
					assign node127 = (inp[6]) ? node129 : 63'b100111101001100000110001101110110011010101001000101101001000101;
						assign node129 = (inp[4]) ? node131 : 63'b100111101000000000110001100000110011010101001100101100001010101;
							assign node131 = (inp[5]) ? 63'b100111101001000000110001101000110111010101001101101100001010101 : 63'b100111101001000000110001101000110111010101001100101100001010101;
					assign node134 = (inp[6]) ? node140 : node135;
						assign node135 = (inp[5]) ? node137 : 63'b100111101001100000110001101110110011010101001100101101000010101;
							assign node137 = (inp[0]) ? 63'b100111101001100000110001101110110011010101001101101101000010101 : 63'b100111101001100000110001101110110011010101001100101101000010101;
						assign node140 = (inp[0]) ? 63'b100111101001100000110001001110110011010101001101101101000010101 : 63'b100111101001100000110001001110110011010101001100101101000010101;
				assign node143 = (inp[6]) ? node153 : node144;
					assign node144 = (inp[4]) ? node148 : node145;
						assign node145 = (inp[1]) ? 63'b100111101000000000110001100000110011010101001100101100001010101 : 63'b100001101000000000110001100000110011010101001100101100001010101;
						assign node148 = (inp[5]) ? node150 : 63'b000111101001001000110001101010110011000101001100101101001010101;
							assign node150 = (inp[0]) ? 63'b000111101001001000110001101010110011000101001101101101001010101 : 63'b000111101001001000110001101010110011000101001100101101001010101;
					assign node153 = (inp[1]) ? node161 : node154;
						assign node154 = (inp[4]) ? node156 : 63'b100111101011100000100001101110110010010101001100101101000010101;
							assign node156 = (inp[5]) ? node158 : 63'b100111101001100000100001101110110010010101001100101101000010101;
								assign node158 = (inp[0]) ? 63'b100111101001100000100001101110110010010101001101101101000010101 : 63'b100111101001100000100001101110110010010101001100101101000010101;
						assign node161 = (inp[4]) ? node163 : 63'b100111101000000000110000100100110011010101101100101101001010101;
							assign node163 = (inp[5]) ? node165 : 63'b100111101001000000110000100100110011010101101100101101001010101;
								assign node165 = (inp[0]) ? 63'b100111101001000000110000100100110011010101101101101101001010101 : 63'b100111101001000000110000100100110011010101101100101101001010101;
			assign node168 = (inp[0]) ? node206 : node169;
				assign node169 = (inp[5]) ? node195 : node170;
					assign node170 = (inp[6]) ? node182 : node171;
						assign node171 = (inp[4]) ? node177 : node172;
							assign node172 = (inp[1]) ? node174 : 63'b100001101001100000110001111110110011010101001100101101001010101;
								assign node174 = (inp[3]) ? 63'b100111101001100000110001101110110011010101001100001101001010101 : 63'b100111101001100000110001101110110011010101001110101101001010101;
							assign node177 = (inp[3]) ? 63'b100111101001000000110001101110110011100100001100101001001010101 : node178;
								assign node178 = (inp[1]) ? 63'b100111100001000000110001101100110011010101001100111101001010101 : 63'b100111100001000000110001101110110011011100001100101101001010101;
						assign node182 = (inp[4]) ? node188 : node183;
							assign node183 = (inp[1]) ? node185 : 63'b100111101001100000010001101110110011010101001100000101001010101;
								assign node185 = (inp[3]) ? 63'b100111101001100000010001101110110011010101001100001101001010101 : 63'b100111101001100000110001101110110011010001001100101101001010100;
							assign node188 = (inp[3]) ? node192 : node189;
								assign node189 = (inp[1]) ? 63'b100111101001100010110001101110110011010101001100101101001000101 : 63'b100111101001100000110001101110110011010101001100101101001010101;
								assign node192 = (inp[1]) ? 63'b100111001001100000110001101110110011010101000100101101001000001 : 63'b100111001001100000110001101110110001010101000100101101001000001;
					assign node195 = (inp[4]) ? node201 : node196;
						assign node196 = (inp[1]) ? 63'b100111101001100100110001101110110011010101001100101101001010101 : node197;
							assign node197 = (inp[3]) ? 63'b100001101001100100110001101110110011010101001100101101001010101 : 63'b100111101001100100110001101110110011010101001100101101001010101;
						assign node201 = (inp[1]) ? node203 : 63'b100101101001110000110001101110110011010101001100101101001010101;
							assign node203 = (inp[6]) ? 63'b000111101001100000110001101110110011000101001100101101001010101 : 63'b100111101001100000110001101110110011010101001100101101001010101;
				assign node206 = (inp[4]) ? node214 : node207;
					assign node207 = (inp[5]) ? node209 : 63'b100111101001100000110001101110110011010101001100101101001010101;
						assign node209 = (inp[3]) ? node211 : 63'b100111101001000000110001101110110011000110001100101001001010101;
							assign node211 = (inp[6]) ? 63'b100111101011000000110001101110110011000110001100101001001010101 : 63'b100001101001000000110001101110110011000110001100101001001010101;
					assign node214 = (inp[6]) ? node224 : node215;
						assign node215 = (inp[3]) ? node221 : node216;
							assign node216 = (inp[1]) ? node218 : 63'b100111101001100000110001101110110011010101011000101101001000101;
								assign node218 = (inp[5]) ? 63'b100111101001100000110001101110110011010101011101101101000010101 : 63'b100111101001100000110001101110110011010101011100101101000010101;
							assign node221 = (inp[1]) ? 63'b100111101000000000110000101100110011010101011100101101001011101 : 63'b100111101000000000110001101001110011010101011100101100001010101;
						assign node224 = (inp[1]) ? node230 : node225;
							assign node225 = (inp[3]) ? node227 : 63'b100111101001100000110001001110111010010101011100101101000010101;
								assign node227 = (inp[5]) ? 63'b100111101001100000100001101110110010010101011101101101000010101 : 63'b100111101001100000100001101110110010010101011100101101000010101;
							assign node230 = (inp[3]) ? node234 : node231;
								assign node231 = (inp[5]) ? 63'b100111101001100000110001001110110011010101011101101101000010101 : 63'b100111101001100000110001001110110011010101011100101101000010101;
								assign node234 = (inp[5]) ? 63'b100111101001100000110001101110110011010101011101101101001010101 : 63'b100111101101100000110001101110110011010101011100101101001010101;

endmodule