module dtc_split66_bm59 (
	input  wire [12-1:0] inp,
	output wire [3-1:0] outp
);

	wire [3-1:0] node1;
	wire [3-1:0] node2;
	wire [3-1:0] node3;
	wire [3-1:0] node4;
	wire [3-1:0] node5;
	wire [3-1:0] node6;
	wire [3-1:0] node7;
	wire [3-1:0] node8;
	wire [3-1:0] node10;
	wire [3-1:0] node11;
	wire [3-1:0] node15;
	wire [3-1:0] node17;
	wire [3-1:0] node20;
	wire [3-1:0] node21;
	wire [3-1:0] node23;
	wire [3-1:0] node24;
	wire [3-1:0] node27;
	wire [3-1:0] node30;
	wire [3-1:0] node32;
	wire [3-1:0] node33;
	wire [3-1:0] node37;
	wire [3-1:0] node38;
	wire [3-1:0] node39;
	wire [3-1:0] node41;
	wire [3-1:0] node42;
	wire [3-1:0] node46;
	wire [3-1:0] node48;
	wire [3-1:0] node51;
	wire [3-1:0] node52;
	wire [3-1:0] node53;
	wire [3-1:0] node55;
	wire [3-1:0] node58;
	wire [3-1:0] node61;
	wire [3-1:0] node62;
	wire [3-1:0] node65;
	wire [3-1:0] node66;
	wire [3-1:0] node70;
	wire [3-1:0] node72;
	wire [3-1:0] node73;
	wire [3-1:0] node74;
	wire [3-1:0] node75;
	wire [3-1:0] node77;
	wire [3-1:0] node79;
	wire [3-1:0] node82;
	wire [3-1:0] node83;
	wire [3-1:0] node84;
	wire [3-1:0] node89;
	wire [3-1:0] node90;
	wire [3-1:0] node91;
	wire [3-1:0] node95;
	wire [3-1:0] node97;
	wire [3-1:0] node100;
	wire [3-1:0] node101;
	wire [3-1:0] node102;
	wire [3-1:0] node106;
	wire [3-1:0] node108;
	wire [3-1:0] node112;
	wire [3-1:0] node113;
	wire [3-1:0] node114;
	wire [3-1:0] node115;
	wire [3-1:0] node116;
	wire [3-1:0] node117;
	wire [3-1:0] node119;
	wire [3-1:0] node120;
	wire [3-1:0] node122;
	wire [3-1:0] node126;
	wire [3-1:0] node127;
	wire [3-1:0] node130;
	wire [3-1:0] node131;
	wire [3-1:0] node135;
	wire [3-1:0] node136;
	wire [3-1:0] node137;
	wire [3-1:0] node140;
	wire [3-1:0] node141;
	wire [3-1:0] node143;
	wire [3-1:0] node147;
	wire [3-1:0] node148;
	wire [3-1:0] node149;
	wire [3-1:0] node152;
	wire [3-1:0] node153;
	wire [3-1:0] node157;
	wire [3-1:0] node159;
	wire [3-1:0] node162;
	wire [3-1:0] node163;
	wire [3-1:0] node164;
	wire [3-1:0] node165;
	wire [3-1:0] node167;
	wire [3-1:0] node170;
	wire [3-1:0] node171;
	wire [3-1:0] node174;
	wire [3-1:0] node177;
	wire [3-1:0] node178;
	wire [3-1:0] node180;
	wire [3-1:0] node183;
	wire [3-1:0] node184;
	wire [3-1:0] node187;
	wire [3-1:0] node190;
	wire [3-1:0] node191;
	wire [3-1:0] node192;
	wire [3-1:0] node194;
	wire [3-1:0] node198;
	wire [3-1:0] node200;
	wire [3-1:0] node203;
	wire [3-1:0] node204;
	wire [3-1:0] node205;
	wire [3-1:0] node206;
	wire [3-1:0] node207;
	wire [3-1:0] node208;
	wire [3-1:0] node212;
	wire [3-1:0] node215;
	wire [3-1:0] node217;
	wire [3-1:0] node218;
	wire [3-1:0] node220;
	wire [3-1:0] node224;
	wire [3-1:0] node225;
	wire [3-1:0] node226;
	wire [3-1:0] node228;
	wire [3-1:0] node229;
	wire [3-1:0] node233;
	wire [3-1:0] node234;
	wire [3-1:0] node237;
	wire [3-1:0] node240;
	wire [3-1:0] node241;
	wire [3-1:0] node243;
	wire [3-1:0] node246;
	wire [3-1:0] node248;
	wire [3-1:0] node252;
	wire [3-1:0] node253;
	wire [3-1:0] node254;
	wire [3-1:0] node255;
	wire [3-1:0] node256;
	wire [3-1:0] node257;
	wire [3-1:0] node259;
	wire [3-1:0] node260;
	wire [3-1:0] node264;
	wire [3-1:0] node265;
	wire [3-1:0] node269;
	wire [3-1:0] node270;
	wire [3-1:0] node271;
	wire [3-1:0] node272;
	wire [3-1:0] node278;
	wire [3-1:0] node279;
	wire [3-1:0] node281;
	wire [3-1:0] node282;
	wire [3-1:0] node284;
	wire [3-1:0] node287;
	wire [3-1:0] node289;
	wire [3-1:0] node292;
	wire [3-1:0] node293;
	wire [3-1:0] node297;
	wire [3-1:0] node298;
	wire [3-1:0] node299;
	wire [3-1:0] node300;
	wire [3-1:0] node301;
	wire [3-1:0] node305;
	wire [3-1:0] node306;
	wire [3-1:0] node310;
	wire [3-1:0] node311;
	wire [3-1:0] node312;
	wire [3-1:0] node313;
	wire [3-1:0] node316;
	wire [3-1:0] node319;
	wire [3-1:0] node321;
	wire [3-1:0] node324;
	wire [3-1:0] node325;
	wire [3-1:0] node327;
	wire [3-1:0] node331;
	wire [3-1:0] node332;
	wire [3-1:0] node333;
	wire [3-1:0] node335;
	wire [3-1:0] node338;
	wire [3-1:0] node341;
	wire [3-1:0] node342;
	wire [3-1:0] node344;
	wire [3-1:0] node345;
	wire [3-1:0] node350;
	wire [3-1:0] node351;
	wire [3-1:0] node352;
	wire [3-1:0] node353;
	wire [3-1:0] node354;
	wire [3-1:0] node355;
	wire [3-1:0] node359;
	wire [3-1:0] node360;
	wire [3-1:0] node362;
	wire [3-1:0] node365;
	wire [3-1:0] node366;
	wire [3-1:0] node369;
	wire [3-1:0] node372;
	wire [3-1:0] node374;
	wire [3-1:0] node376;
	wire [3-1:0] node379;
	wire [3-1:0] node380;
	wire [3-1:0] node382;
	wire [3-1:0] node383;
	wire [3-1:0] node384;
	wire [3-1:0] node390;
	wire [3-1:0] node391;
	wire [3-1:0] node392;
	wire [3-1:0] node393;
	wire [3-1:0] node394;
	wire [3-1:0] node396;
	wire [3-1:0] node399;
	wire [3-1:0] node401;
	wire [3-1:0] node404;
	wire [3-1:0] node406;
	wire [3-1:0] node407;
	wire [3-1:0] node410;
	wire [3-1:0] node415;
	wire [3-1:0] node416;
	wire [3-1:0] node417;
	wire [3-1:0] node418;
	wire [3-1:0] node420;
	wire [3-1:0] node421;
	wire [3-1:0] node422;
	wire [3-1:0] node423;
	wire [3-1:0] node427;
	wire [3-1:0] node428;
	wire [3-1:0] node431;
	wire [3-1:0] node433;
	wire [3-1:0] node437;
	wire [3-1:0] node438;
	wire [3-1:0] node439;
	wire [3-1:0] node440;
	wire [3-1:0] node441;
	wire [3-1:0] node443;
	wire [3-1:0] node445;
	wire [3-1:0] node448;
	wire [3-1:0] node449;
	wire [3-1:0] node450;
	wire [3-1:0] node455;
	wire [3-1:0] node456;
	wire [3-1:0] node459;
	wire [3-1:0] node460;
	wire [3-1:0] node464;
	wire [3-1:0] node465;
	wire [3-1:0] node466;
	wire [3-1:0] node467;
	wire [3-1:0] node469;
	wire [3-1:0] node473;
	wire [3-1:0] node474;
	wire [3-1:0] node478;
	wire [3-1:0] node479;
	wire [3-1:0] node482;
	wire [3-1:0] node484;
	wire [3-1:0] node487;
	wire [3-1:0] node489;
	wire [3-1:0] node490;
	wire [3-1:0] node492;
	wire [3-1:0] node493;
	wire [3-1:0] node497;
	wire [3-1:0] node499;
	wire [3-1:0] node500;
	wire [3-1:0] node504;
	wire [3-1:0] node505;
	wire [3-1:0] node506;
	wire [3-1:0] node507;
	wire [3-1:0] node508;
	wire [3-1:0] node510;
	wire [3-1:0] node511;
	wire [3-1:0] node512;
	wire [3-1:0] node515;
	wire [3-1:0] node518;
	wire [3-1:0] node521;
	wire [3-1:0] node522;
	wire [3-1:0] node523;
	wire [3-1:0] node525;
	wire [3-1:0] node528;
	wire [3-1:0] node530;
	wire [3-1:0] node533;
	wire [3-1:0] node534;
	wire [3-1:0] node537;
	wire [3-1:0] node538;
	wire [3-1:0] node542;
	wire [3-1:0] node543;
	wire [3-1:0] node544;
	wire [3-1:0] node546;
	wire [3-1:0] node547;
	wire [3-1:0] node550;
	wire [3-1:0] node553;
	wire [3-1:0] node554;
	wire [3-1:0] node557;
	wire [3-1:0] node560;
	wire [3-1:0] node561;
	wire [3-1:0] node563;
	wire [3-1:0] node566;
	wire [3-1:0] node569;
	wire [3-1:0] node570;
	wire [3-1:0] node571;
	wire [3-1:0] node572;
	wire [3-1:0] node573;
	wire [3-1:0] node574;
	wire [3-1:0] node578;
	wire [3-1:0] node581;
	wire [3-1:0] node582;
	wire [3-1:0] node583;
	wire [3-1:0] node588;
	wire [3-1:0] node589;
	wire [3-1:0] node591;
	wire [3-1:0] node594;
	wire [3-1:0] node597;
	wire [3-1:0] node598;
	wire [3-1:0] node599;
	wire [3-1:0] node600;
	wire [3-1:0] node605;
	wire [3-1:0] node606;
	wire [3-1:0] node607;
	wire [3-1:0] node611;
	wire [3-1:0] node614;
	wire [3-1:0] node615;
	wire [3-1:0] node616;
	wire [3-1:0] node617;
	wire [3-1:0] node618;
	wire [3-1:0] node619;
	wire [3-1:0] node623;
	wire [3-1:0] node624;
	wire [3-1:0] node625;
	wire [3-1:0] node629;
	wire [3-1:0] node632;
	wire [3-1:0] node633;
	wire [3-1:0] node634;
	wire [3-1:0] node639;
	wire [3-1:0] node640;
	wire [3-1:0] node641;
	wire [3-1:0] node642;
	wire [3-1:0] node645;
	wire [3-1:0] node648;
	wire [3-1:0] node650;
	wire [3-1:0] node654;
	wire [3-1:0] node655;
	wire [3-1:0] node656;
	wire [3-1:0] node657;
	wire [3-1:0] node658;
	wire [3-1:0] node661;
	wire [3-1:0] node664;
	wire [3-1:0] node665;
	wire [3-1:0] node668;
	wire [3-1:0] node671;
	wire [3-1:0] node672;
	wire [3-1:0] node673;
	wire [3-1:0] node674;
	wire [3-1:0] node677;
	wire [3-1:0] node680;
	wire [3-1:0] node682;
	wire [3-1:0] node686;
	wire [3-1:0] node687;
	wire [3-1:0] node688;
	wire [3-1:0] node689;
	wire [3-1:0] node694;
	wire [3-1:0] node697;
	wire [3-1:0] node699;
	wire [3-1:0] node700;
	wire [3-1:0] node702;
	wire [3-1:0] node703;
	wire [3-1:0] node704;
	wire [3-1:0] node705;
	wire [3-1:0] node706;
	wire [3-1:0] node710;
	wire [3-1:0] node711;
	wire [3-1:0] node715;
	wire [3-1:0] node717;
	wire [3-1:0] node718;
	wire [3-1:0] node720;
	wire [3-1:0] node723;
	wire [3-1:0] node727;
	wire [3-1:0] node728;
	wire [3-1:0] node729;
	wire [3-1:0] node730;
	wire [3-1:0] node731;
	wire [3-1:0] node732;
	wire [3-1:0] node734;
	wire [3-1:0] node737;
	wire [3-1:0] node739;
	wire [3-1:0] node742;
	wire [3-1:0] node745;
	wire [3-1:0] node746;
	wire [3-1:0] node747;
	wire [3-1:0] node750;
	wire [3-1:0] node753;
	wire [3-1:0] node754;
	wire [3-1:0] node755;
	wire [3-1:0] node760;
	wire [3-1:0] node761;
	wire [3-1:0] node762;
	wire [3-1:0] node763;
	wire [3-1:0] node768;
	wire [3-1:0] node769;
	wire [3-1:0] node770;
	wire [3-1:0] node775;
	wire [3-1:0] node777;
	wire [3-1:0] node778;
	wire [3-1:0] node779;
	wire [3-1:0] node780;
	wire [3-1:0] node785;
	wire [3-1:0] node787;
	wire [3-1:0] node788;
	wire [3-1:0] node792;
	wire [3-1:0] node793;
	wire [3-1:0] node794;
	wire [3-1:0] node795;
	wire [3-1:0] node796;
	wire [3-1:0] node797;
	wire [3-1:0] node798;
	wire [3-1:0] node799;
	wire [3-1:0] node801;
	wire [3-1:0] node802;
	wire [3-1:0] node803;
	wire [3-1:0] node808;
	wire [3-1:0] node809;
	wire [3-1:0] node811;
	wire [3-1:0] node813;
	wire [3-1:0] node816;
	wire [3-1:0] node819;
	wire [3-1:0] node820;
	wire [3-1:0] node821;
	wire [3-1:0] node822;
	wire [3-1:0] node823;
	wire [3-1:0] node829;
	wire [3-1:0] node830;
	wire [3-1:0] node831;
	wire [3-1:0] node834;
	wire [3-1:0] node835;
	wire [3-1:0] node839;
	wire [3-1:0] node840;
	wire [3-1:0] node842;
	wire [3-1:0] node847;
	wire [3-1:0] node848;
	wire [3-1:0] node849;
	wire [3-1:0] node850;
	wire [3-1:0] node851;
	wire [3-1:0] node853;
	wire [3-1:0] node854;
	wire [3-1:0] node858;
	wire [3-1:0] node859;
	wire [3-1:0] node863;
	wire [3-1:0] node864;
	wire [3-1:0] node868;
	wire [3-1:0] node869;
	wire [3-1:0] node870;
	wire [3-1:0] node874;
	wire [3-1:0] node875;
	wire [3-1:0] node876;
	wire [3-1:0] node880;
	wire [3-1:0] node883;
	wire [3-1:0] node884;
	wire [3-1:0] node885;
	wire [3-1:0] node886;
	wire [3-1:0] node890;
	wire [3-1:0] node891;
	wire [3-1:0] node895;
	wire [3-1:0] node896;
	wire [3-1:0] node897;
	wire [3-1:0] node899;
	wire [3-1:0] node902;
	wire [3-1:0] node904;
	wire [3-1:0] node907;
	wire [3-1:0] node908;
	wire [3-1:0] node911;
	wire [3-1:0] node915;
	wire [3-1:0] node916;
	wire [3-1:0] node917;
	wire [3-1:0] node918;
	wire [3-1:0] node919;
	wire [3-1:0] node920;
	wire [3-1:0] node921;
	wire [3-1:0] node922;
	wire [3-1:0] node923;
	wire [3-1:0] node927;
	wire [3-1:0] node930;
	wire [3-1:0] node932;
	wire [3-1:0] node935;
	wire [3-1:0] node936;
	wire [3-1:0] node937;
	wire [3-1:0] node941;
	wire [3-1:0] node943;
	wire [3-1:0] node945;
	wire [3-1:0] node948;
	wire [3-1:0] node949;
	wire [3-1:0] node950;
	wire [3-1:0] node952;
	wire [3-1:0] node955;
	wire [3-1:0] node956;
	wire [3-1:0] node959;
	wire [3-1:0] node960;
	wire [3-1:0] node963;
	wire [3-1:0] node966;
	wire [3-1:0] node967;
	wire [3-1:0] node969;
	wire [3-1:0] node972;
	wire [3-1:0] node975;
	wire [3-1:0] node976;
	wire [3-1:0] node977;
	wire [3-1:0] node978;
	wire [3-1:0] node980;
	wire [3-1:0] node983;
	wire [3-1:0] node986;
	wire [3-1:0] node987;
	wire [3-1:0] node988;
	wire [3-1:0] node992;
	wire [3-1:0] node995;
	wire [3-1:0] node996;
	wire [3-1:0] node997;
	wire [3-1:0] node999;
	wire [3-1:0] node1003;
	wire [3-1:0] node1005;
	wire [3-1:0] node1008;
	wire [3-1:0] node1009;
	wire [3-1:0] node1010;
	wire [3-1:0] node1011;
	wire [3-1:0] node1012;
	wire [3-1:0] node1015;
	wire [3-1:0] node1019;
	wire [3-1:0] node1021;
	wire [3-1:0] node1022;
	wire [3-1:0] node1023;
	wire [3-1:0] node1026;
	wire [3-1:0] node1029;
	wire [3-1:0] node1031;
	wire [3-1:0] node1035;
	wire [3-1:0] node1036;
	wire [3-1:0] node1037;
	wire [3-1:0] node1038;
	wire [3-1:0] node1039;
	wire [3-1:0] node1040;
	wire [3-1:0] node1042;
	wire [3-1:0] node1044;
	wire [3-1:0] node1047;
	wire [3-1:0] node1048;
	wire [3-1:0] node1052;
	wire [3-1:0] node1054;
	wire [3-1:0] node1055;
	wire [3-1:0] node1059;
	wire [3-1:0] node1060;
	wire [3-1:0] node1061;
	wire [3-1:0] node1062;
	wire [3-1:0] node1065;
	wire [3-1:0] node1067;
	wire [3-1:0] node1070;
	wire [3-1:0] node1071;
	wire [3-1:0] node1073;
	wire [3-1:0] node1077;
	wire [3-1:0] node1078;
	wire [3-1:0] node1080;
	wire [3-1:0] node1083;
	wire [3-1:0] node1084;
	wire [3-1:0] node1087;
	wire [3-1:0] node1090;
	wire [3-1:0] node1091;
	wire [3-1:0] node1092;
	wire [3-1:0] node1094;
	wire [3-1:0] node1095;
	wire [3-1:0] node1099;
	wire [3-1:0] node1100;
	wire [3-1:0] node1103;
	wire [3-1:0] node1105;
	wire [3-1:0] node1107;
	wire [3-1:0] node1110;
	wire [3-1:0] node1111;
	wire [3-1:0] node1112;
	wire [3-1:0] node1114;
	wire [3-1:0] node1117;
	wire [3-1:0] node1118;
	wire [3-1:0] node1123;
	wire [3-1:0] node1124;
	wire [3-1:0] node1125;
	wire [3-1:0] node1126;
	wire [3-1:0] node1128;
	wire [3-1:0] node1129;
	wire [3-1:0] node1131;
	wire [3-1:0] node1134;
	wire [3-1:0] node1137;
	wire [3-1:0] node1139;
	wire [3-1:0] node1140;
	wire [3-1:0] node1144;
	wire [3-1:0] node1145;
	wire [3-1:0] node1146;
	wire [3-1:0] node1147;
	wire [3-1:0] node1149;
	wire [3-1:0] node1153;
	wire [3-1:0] node1155;
	wire [3-1:0] node1157;
	wire [3-1:0] node1161;
	wire [3-1:0] node1162;
	wire [3-1:0] node1163;
	wire [3-1:0] node1165;
	wire [3-1:0] node1166;
	wire [3-1:0] node1167;
	wire [3-1:0] node1174;
	wire [3-1:0] node1175;
	wire [3-1:0] node1176;
	wire [3-1:0] node1177;
	wire [3-1:0] node1178;
	wire [3-1:0] node1180;
	wire [3-1:0] node1181;
	wire [3-1:0] node1182;
	wire [3-1:0] node1183;
	wire [3-1:0] node1188;
	wire [3-1:0] node1190;
	wire [3-1:0] node1192;
	wire [3-1:0] node1195;
	wire [3-1:0] node1196;
	wire [3-1:0] node1197;
	wire [3-1:0] node1198;
	wire [3-1:0] node1200;
	wire [3-1:0] node1203;
	wire [3-1:0] node1205;
	wire [3-1:0] node1208;
	wire [3-1:0] node1209;
	wire [3-1:0] node1210;
	wire [3-1:0] node1215;
	wire [3-1:0] node1216;
	wire [3-1:0] node1217;
	wire [3-1:0] node1219;
	wire [3-1:0] node1222;
	wire [3-1:0] node1224;
	wire [3-1:0] node1227;
	wire [3-1:0] node1228;
	wire [3-1:0] node1229;
	wire [3-1:0] node1234;
	wire [3-1:0] node1236;
	wire [3-1:0] node1238;
	wire [3-1:0] node1239;
	wire [3-1:0] node1240;
	wire [3-1:0] node1242;
	wire [3-1:0] node1246;
	wire [3-1:0] node1247;
	wire [3-1:0] node1249;
	wire [3-1:0] node1252;
	wire [3-1:0] node1254;
	wire [3-1:0] node1256;
	wire [3-1:0] node1259;
	wire [3-1:0] node1260;
	wire [3-1:0] node1261;
	wire [3-1:0] node1262;
	wire [3-1:0] node1263;
	wire [3-1:0] node1264;
	wire [3-1:0] node1265;
	wire [3-1:0] node1268;
	wire [3-1:0] node1271;
	wire [3-1:0] node1272;
	wire [3-1:0] node1273;
	wire [3-1:0] node1278;
	wire [3-1:0] node1279;
	wire [3-1:0] node1280;
	wire [3-1:0] node1284;
	wire [3-1:0] node1285;
	wire [3-1:0] node1287;
	wire [3-1:0] node1290;
	wire [3-1:0] node1292;
	wire [3-1:0] node1295;
	wire [3-1:0] node1296;
	wire [3-1:0] node1297;
	wire [3-1:0] node1298;
	wire [3-1:0] node1301;
	wire [3-1:0] node1302;
	wire [3-1:0] node1306;
	wire [3-1:0] node1307;
	wire [3-1:0] node1309;
	wire [3-1:0] node1312;
	wire [3-1:0] node1315;
	wire [3-1:0] node1316;
	wire [3-1:0] node1317;
	wire [3-1:0] node1318;
	wire [3-1:0] node1321;
	wire [3-1:0] node1325;
	wire [3-1:0] node1328;
	wire [3-1:0] node1329;
	wire [3-1:0] node1330;
	wire [3-1:0] node1331;
	wire [3-1:0] node1332;
	wire [3-1:0] node1334;
	wire [3-1:0] node1337;
	wire [3-1:0] node1339;
	wire [3-1:0] node1343;
	wire [3-1:0] node1344;
	wire [3-1:0] node1346;
	wire [3-1:0] node1349;
	wire [3-1:0] node1352;
	wire [3-1:0] node1353;
	wire [3-1:0] node1354;
	wire [3-1:0] node1355;
	wire [3-1:0] node1358;
	wire [3-1:0] node1361;
	wire [3-1:0] node1362;
	wire [3-1:0] node1363;
	wire [3-1:0] node1366;
	wire [3-1:0] node1369;
	wire [3-1:0] node1372;
	wire [3-1:0] node1374;
	wire [3-1:0] node1377;
	wire [3-1:0] node1378;
	wire [3-1:0] node1379;
	wire [3-1:0] node1380;
	wire [3-1:0] node1381;
	wire [3-1:0] node1382;
	wire [3-1:0] node1386;
	wire [3-1:0] node1387;
	wire [3-1:0] node1391;
	wire [3-1:0] node1392;
	wire [3-1:0] node1393;
	wire [3-1:0] node1397;
	wire [3-1:0] node1398;
	wire [3-1:0] node1401;
	wire [3-1:0] node1404;
	wire [3-1:0] node1405;
	wire [3-1:0] node1406;
	wire [3-1:0] node1407;
	wire [3-1:0] node1410;
	wire [3-1:0] node1414;
	wire [3-1:0] node1416;
	wire [3-1:0] node1418;
	wire [3-1:0] node1421;
	wire [3-1:0] node1422;
	wire [3-1:0] node1423;
	wire [3-1:0] node1424;
	wire [3-1:0] node1426;
	wire [3-1:0] node1429;
	wire [3-1:0] node1432;
	wire [3-1:0] node1433;
	wire [3-1:0] node1437;
	wire [3-1:0] node1439;
	wire [3-1:0] node1441;
	wire [3-1:0] node1442;
	wire [3-1:0] node1446;
	wire [3-1:0] node1447;
	wire [3-1:0] node1449;
	wire [3-1:0] node1450;
	wire [3-1:0] node1452;
	wire [3-1:0] node1453;
	wire [3-1:0] node1455;
	wire [3-1:0] node1457;
	wire [3-1:0] node1459;
	wire [3-1:0] node1463;
	wire [3-1:0] node1464;
	wire [3-1:0] node1465;
	wire [3-1:0] node1466;
	wire [3-1:0] node1467;
	wire [3-1:0] node1470;
	wire [3-1:0] node1471;
	wire [3-1:0] node1476;
	wire [3-1:0] node1477;
	wire [3-1:0] node1480;
	wire [3-1:0] node1482;
	wire [3-1:0] node1483;
	wire [3-1:0] node1487;
	wire [3-1:0] node1488;
	wire [3-1:0] node1489;
	wire [3-1:0] node1490;
	wire [3-1:0] node1492;
	wire [3-1:0] node1496;
	wire [3-1:0] node1497;
	wire [3-1:0] node1498;
	wire [3-1:0] node1503;
	wire [3-1:0] node1504;
	wire [3-1:0] node1505;

	assign outp = (inp[10]) ? node792 : node1;
		assign node1 = (inp[9]) ? node415 : node2;
			assign node2 = (inp[2]) ? node112 : node3;
				assign node3 = (inp[0]) ? 3'b110 : node4;
					assign node4 = (inp[3]) ? node70 : node5;
						assign node5 = (inp[7]) ? node37 : node6;
							assign node6 = (inp[8]) ? node20 : node7;
								assign node7 = (inp[5]) ? node15 : node8;
									assign node8 = (inp[6]) ? node10 : 3'b000;
										assign node10 = (inp[11]) ? 3'b000 : node11;
											assign node11 = (inp[4]) ? 3'b010 : 3'b110;
									assign node15 = (inp[6]) ? node17 : 3'b010;
										assign node17 = (inp[11]) ? 3'b010 : 3'b000;
								assign node20 = (inp[4]) ? node30 : node21;
									assign node21 = (inp[1]) ? node23 : 3'b111;
										assign node23 = (inp[5]) ? node27 : node24;
											assign node24 = (inp[6]) ? 3'b110 : 3'b100;
											assign node27 = (inp[11]) ? 3'b110 : 3'b100;
									assign node30 = (inp[5]) ? node32 : 3'b000;
										assign node32 = (inp[11]) ? 3'b010 : node33;
											assign node33 = (inp[6]) ? 3'b000 : 3'b010;
							assign node37 = (inp[8]) ? node51 : node38;
								assign node38 = (inp[5]) ? node46 : node39;
									assign node39 = (inp[6]) ? node41 : 3'b100;
										assign node41 = (inp[11]) ? 3'b100 : node42;
											assign node42 = (inp[1]) ? 3'b110 : 3'b010;
									assign node46 = (inp[6]) ? node48 : 3'b110;
										assign node48 = (inp[11]) ? 3'b110 : 3'b100;
								assign node51 = (inp[4]) ? node61 : node52;
									assign node52 = (inp[5]) ? node58 : node53;
										assign node53 = (inp[6]) ? node55 : 3'b000;
											assign node55 = (inp[11]) ? 3'b000 : 3'b010;
										assign node58 = (inp[6]) ? 3'b000 : 3'b010;
									assign node61 = (inp[6]) ? node65 : node62;
										assign node62 = (inp[5]) ? 3'b110 : 3'b100;
										assign node65 = (inp[5]) ? 3'b100 : node66;
											assign node66 = (inp[11]) ? 3'b100 : 3'b010;
						assign node70 = (inp[1]) ? node72 : 3'b111;
							assign node72 = (inp[5]) ? node100 : node73;
								assign node73 = (inp[11]) ? node89 : node74;
									assign node74 = (inp[6]) ? node82 : node75;
										assign node75 = (inp[7]) ? node77 : 3'b000;
											assign node77 = (inp[8]) ? node79 : 3'b100;
												assign node79 = (inp[4]) ? 3'b100 : 3'b000;
										assign node82 = (inp[7]) ? 3'b010 : node83;
											assign node83 = (inp[8]) ? 3'b111 : node84;
												assign node84 = (inp[4]) ? 3'b010 : 3'b111;
									assign node89 = (inp[7]) ? node95 : node90;
										assign node90 = (inp[4]) ? 3'b000 : node91;
											assign node91 = (inp[6]) ? 3'b000 : 3'b111;
										assign node95 = (inp[8]) ? node97 : 3'b100;
											assign node97 = (inp[4]) ? 3'b100 : 3'b000;
								assign node100 = (inp[7]) ? node106 : node101;
									assign node101 = (inp[8]) ? 3'b111 : node102;
										assign node102 = (inp[6]) ? 3'b000 : 3'b010;
									assign node106 = (inp[8]) ? node108 : 3'b110;
										assign node108 = (inp[4]) ? 3'b100 : 3'b010;
				assign node112 = (inp[1]) ? node252 : node113;
					assign node113 = (inp[0]) ? node203 : node114;
						assign node114 = (inp[11]) ? node162 : node115;
							assign node115 = (inp[4]) ? node135 : node116;
								assign node116 = (inp[8]) ? node126 : node117;
									assign node117 = (inp[3]) ? node119 : 3'b000;
										assign node119 = (inp[7]) ? 3'b000 : node120;
											assign node120 = (inp[5]) ? node122 : 3'b000;
												assign node122 = (inp[6]) ? 3'b000 : 3'b010;
									assign node126 = (inp[7]) ? node130 : node127;
										assign node127 = (inp[6]) ? 3'b000 : 3'b110;
										assign node130 = (inp[3]) ? 3'b000 : node131;
											assign node131 = (inp[5]) ? 3'b000 : 3'b100;
								assign node135 = (inp[8]) ? node147 : node136;
									assign node136 = (inp[3]) ? node140 : node137;
										assign node137 = (inp[7]) ? 3'b000 : 3'b100;
										assign node140 = (inp[7]) ? 3'b100 : node141;
											assign node141 = (inp[6]) ? node143 : 3'b000;
												assign node143 = (inp[5]) ? 3'b000 : 3'b010;
									assign node147 = (inp[5]) ? node157 : node148;
										assign node148 = (inp[7]) ? node152 : node149;
											assign node149 = (inp[3]) ? 3'b110 : 3'b000;
											assign node152 = (inp[6]) ? 3'b000 : node153;
												assign node153 = (inp[3]) ? 3'b000 : 3'b010;
										assign node157 = (inp[7]) ? node159 : 3'b100;
											assign node159 = (inp[3]) ? 3'b100 : 3'b010;
							assign node162 = (inp[5]) ? node190 : node163;
								assign node163 = (inp[3]) ? node177 : node164;
									assign node164 = (inp[4]) ? node170 : node165;
										assign node165 = (inp[8]) ? node167 : 3'b010;
											assign node167 = (inp[7]) ? 3'b110 : 3'b100;
										assign node170 = (inp[8]) ? node174 : node171;
											assign node171 = (inp[7]) ? 3'b100 : 3'b110;
											assign node174 = (inp[7]) ? 3'b000 : 3'b010;
									assign node177 = (inp[7]) ? node183 : node178;
										assign node178 = (inp[8]) ? node180 : 3'b000;
											assign node180 = (inp[4]) ? 3'b000 : 3'b100;
										assign node183 = (inp[8]) ? node187 : node184;
											assign node184 = (inp[4]) ? 3'b110 : 3'b010;
											assign node187 = (inp[4]) ? 3'b010 : 3'b000;
								assign node190 = (inp[4]) ? node198 : node191;
									assign node191 = (inp[7]) ? 3'b010 : node192;
										assign node192 = (inp[3]) ? node194 : 3'b010;
											assign node194 = (inp[8]) ? 3'b110 : 3'b010;
									assign node198 = (inp[3]) ? node200 : 3'b110;
										assign node200 = (inp[7]) ? 3'b110 : 3'b010;
						assign node203 = (inp[3]) ? 3'b110 : node204;
							assign node204 = (inp[5]) ? node224 : node205;
								assign node205 = (inp[6]) ? node215 : node206;
									assign node206 = (inp[7]) ? node212 : node207;
										assign node207 = (inp[4]) ? 3'b000 : node208;
											assign node208 = (inp[8]) ? 3'b110 : 3'b000;
										assign node212 = (inp[8]) ? 3'b000 : 3'b100;
									assign node215 = (inp[11]) ? node217 : 3'b010;
										assign node217 = (inp[7]) ? 3'b100 : node218;
											assign node218 = (inp[8]) ? node220 : 3'b000;
												assign node220 = (inp[4]) ? 3'b000 : 3'b110;
								assign node224 = (inp[11]) ? node240 : node225;
									assign node225 = (inp[6]) ? node233 : node226;
										assign node226 = (inp[8]) ? node228 : 3'b010;
											assign node228 = (inp[4]) ? 3'b110 : node229;
												assign node229 = (inp[7]) ? 3'b010 : 3'b110;
										assign node233 = (inp[8]) ? node237 : node234;
											assign node234 = (inp[7]) ? 3'b100 : 3'b000;
											assign node237 = (inp[7]) ? 3'b000 : 3'b110;
									assign node240 = (inp[7]) ? node246 : node241;
										assign node241 = (inp[8]) ? node243 : 3'b010;
											assign node243 = (inp[4]) ? 3'b010 : 3'b110;
										assign node246 = (inp[8]) ? node248 : 3'b110;
											assign node248 = (inp[4]) ? 3'b110 : 3'b010;
					assign node252 = (inp[7]) ? node350 : node253;
						assign node253 = (inp[8]) ? node297 : node254;
							assign node254 = (inp[0]) ? node278 : node255;
								assign node255 = (inp[5]) ? node269 : node256;
									assign node256 = (inp[4]) ? node264 : node257;
										assign node257 = (inp[3]) ? node259 : 3'b010;
											assign node259 = (inp[11]) ? 3'b000 : node260;
												assign node260 = (inp[6]) ? 3'b000 : 3'b010;
										assign node264 = (inp[11]) ? 3'b010 : node265;
											assign node265 = (inp[3]) ? 3'b010 : 3'b100;
									assign node269 = (inp[6]) ? 3'b010 : node270;
										assign node270 = (inp[4]) ? 3'b010 : node271;
											assign node271 = (inp[3]) ? 3'b110 : node272;
												assign node272 = (inp[11]) ? 3'b010 : 3'b110;
								assign node278 = (inp[11]) ? node292 : node279;
									assign node279 = (inp[4]) ? node281 : 3'b000;
										assign node281 = (inp[3]) ? node287 : node282;
											assign node282 = (inp[5]) ? node284 : 3'b100;
												assign node284 = (inp[6]) ? 3'b010 : 3'b000;
											assign node287 = (inp[6]) ? node289 : 3'b010;
												assign node289 = (inp[5]) ? 3'b000 : 3'b010;
									assign node292 = (inp[5]) ? 3'b010 : node293;
										assign node293 = (inp[4]) ? 3'b000 : 3'b010;
							assign node297 = (inp[5]) ? node331 : node298;
								assign node298 = (inp[4]) ? node310 : node299;
									assign node299 = (inp[0]) ? node305 : node300;
										assign node300 = (inp[6]) ? 3'b100 : node301;
											assign node301 = (inp[3]) ? 3'b000 : 3'b010;
										assign node305 = (inp[3]) ? 3'b110 : node306;
											assign node306 = (inp[6]) ? 3'b110 : 3'b100;
									assign node310 = (inp[6]) ? node324 : node311;
										assign node311 = (inp[0]) ? node319 : node312;
											assign node312 = (inp[3]) ? node316 : node313;
												assign node313 = (inp[11]) ? 3'b100 : 3'b000;
												assign node316 = (inp[11]) ? 3'b010 : 3'b110;
											assign node319 = (inp[11]) ? node321 : 3'b000;
												assign node321 = (inp[3]) ? 3'b000 : 3'b010;
										assign node324 = (inp[3]) ? 3'b110 : node325;
											assign node325 = (inp[11]) ? node327 : 3'b010;
												assign node327 = (inp[0]) ? 3'b010 : 3'b100;
								assign node331 = (inp[4]) ? node341 : node332;
									assign node332 = (inp[0]) ? node338 : node333;
										assign node333 = (inp[11]) ? node335 : 3'b010;
											assign node335 = (inp[3]) ? 3'b010 : 3'b110;
										assign node338 = (inp[3]) ? 3'b110 : 3'b010;
									assign node341 = (inp[11]) ? 3'b010 : node342;
										assign node342 = (inp[6]) ? node344 : 3'b010;
											assign node344 = (inp[0]) ? 3'b000 : node345;
												assign node345 = (inp[3]) ? 3'b010 : 3'b000;
						assign node350 = (inp[4]) ? node390 : node351;
							assign node351 = (inp[5]) ? node379 : node352;
								assign node352 = (inp[3]) ? node372 : node353;
									assign node353 = (inp[11]) ? node359 : node354;
										assign node354 = (inp[8]) ? 3'b010 : node355;
											assign node355 = (inp[0]) ? 3'b010 : 3'b000;
										assign node359 = (inp[6]) ? node365 : node360;
											assign node360 = (inp[8]) ? node362 : 3'b010;
												assign node362 = (inp[0]) ? 3'b010 : 3'b000;
											assign node365 = (inp[0]) ? node369 : node366;
												assign node366 = (inp[8]) ? 3'b000 : 3'b010;
												assign node369 = (inp[8]) ? 3'b010 : 3'b000;
									assign node372 = (inp[0]) ? node374 : 3'b000;
										assign node374 = (inp[8]) ? node376 : 3'b000;
											assign node376 = (inp[6]) ? 3'b010 : 3'b000;
								assign node379 = (inp[11]) ? 3'b010 : node380;
									assign node380 = (inp[0]) ? node382 : 3'b010;
										assign node382 = (inp[6]) ? 3'b000 : node383;
											assign node383 = (inp[3]) ? 3'b000 : node384;
												assign node384 = (inp[8]) ? 3'b010 : 3'b000;
							assign node390 = (inp[5]) ? 3'b000 : node391;
								assign node391 = (inp[11]) ? 3'b000 : node392;
									assign node392 = (inp[6]) ? node404 : node393;
										assign node393 = (inp[0]) ? node399 : node394;
											assign node394 = (inp[8]) ? node396 : 3'b010;
												assign node396 = (inp[3]) ? 3'b000 : 3'b010;
											assign node399 = (inp[3]) ? node401 : 3'b000;
												assign node401 = (inp[8]) ? 3'b010 : 3'b000;
										assign node404 = (inp[0]) ? node406 : 3'b000;
											assign node406 = (inp[3]) ? node410 : node407;
												assign node407 = (inp[8]) ? 3'b010 : 3'b000;
												assign node410 = (inp[8]) ? 3'b000 : 3'b010;
			assign node415 = (inp[0]) ? node697 : node416;
				assign node416 = (inp[2]) ? node504 : node417;
					assign node417 = (inp[1]) ? node437 : node418;
						assign node418 = (inp[7]) ? node420 : 3'b011;
							assign node420 = (inp[3]) ? 3'b011 : node421;
								assign node421 = (inp[4]) ? node427 : node422;
									assign node422 = (inp[8]) ? 3'b011 : node423;
										assign node423 = (inp[11]) ? 3'b010 : 3'b000;
									assign node427 = (inp[5]) ? node431 : node428;
										assign node428 = (inp[11]) ? 3'b000 : 3'b010;
										assign node431 = (inp[6]) ? node433 : 3'b010;
											assign node433 = (inp[11]) ? 3'b010 : 3'b000;
						assign node437 = (inp[3]) ? node487 : node438;
							assign node438 = (inp[5]) ? node464 : node439;
								assign node439 = (inp[11]) ? node455 : node440;
									assign node440 = (inp[6]) ? node448 : node441;
										assign node441 = (inp[7]) ? node443 : 3'b100;
											assign node443 = (inp[8]) ? node445 : 3'b000;
												assign node445 = (inp[4]) ? 3'b000 : 3'b100;
										assign node448 = (inp[8]) ? 3'b110 : node449;
											assign node449 = (inp[7]) ? 3'b010 : node450;
												assign node450 = (inp[4]) ? 3'b110 : 3'b010;
									assign node455 = (inp[7]) ? node459 : node456;
										assign node456 = (inp[4]) ? 3'b100 : 3'b000;
										assign node459 = (inp[4]) ? 3'b000 : node460;
											assign node460 = (inp[8]) ? 3'b100 : 3'b000;
								assign node464 = (inp[7]) ? node478 : node465;
									assign node465 = (inp[4]) ? node473 : node466;
										assign node466 = (inp[8]) ? 3'b010 : node467;
											assign node467 = (inp[6]) ? node469 : 3'b110;
												assign node469 = (inp[11]) ? 3'b110 : 3'b100;
										assign node473 = (inp[11]) ? 3'b110 : node474;
											assign node474 = (inp[6]) ? 3'b100 : 3'b110;
									assign node478 = (inp[4]) ? node482 : node479;
										assign node479 = (inp[8]) ? 3'b110 : 3'b010;
										assign node482 = (inp[6]) ? node484 : 3'b010;
											assign node484 = (inp[11]) ? 3'b010 : 3'b000;
							assign node487 = (inp[7]) ? node489 : 3'b011;
								assign node489 = (inp[8]) ? node497 : node490;
									assign node490 = (inp[5]) ? node492 : 3'b000;
										assign node492 = (inp[11]) ? 3'b010 : node493;
											assign node493 = (inp[4]) ? 3'b010 : 3'b000;
									assign node497 = (inp[4]) ? node499 : 3'b011;
										assign node499 = (inp[6]) ? 3'b000 : node500;
											assign node500 = (inp[5]) ? 3'b010 : 3'b000;
					assign node504 = (inp[7]) ? node614 : node505;
						assign node505 = (inp[5]) ? node569 : node506;
							assign node506 = (inp[8]) ? node542 : node507;
								assign node507 = (inp[6]) ? node521 : node508;
									assign node508 = (inp[1]) ? node510 : 3'b100;
										assign node510 = (inp[4]) ? node518 : node511;
											assign node511 = (inp[11]) ? node515 : node512;
												assign node512 = (inp[3]) ? 3'b100 : 3'b110;
												assign node515 = (inp[3]) ? 3'b110 : 3'b100;
											assign node518 = (inp[3]) ? 3'b100 : 3'b000;
									assign node521 = (inp[11]) ? node533 : node522;
										assign node522 = (inp[1]) ? node528 : node523;
											assign node523 = (inp[4]) ? node525 : 3'b010;
												assign node525 = (inp[3]) ? 3'b110 : 3'b000;
											assign node528 = (inp[3]) ? node530 : 3'b110;
												assign node530 = (inp[4]) ? 3'b000 : 3'b100;
										assign node533 = (inp[3]) ? node537 : node534;
											assign node534 = (inp[4]) ? 3'b010 : 3'b100;
											assign node537 = (inp[4]) ? 3'b100 : node538;
												assign node538 = (inp[1]) ? 3'b110 : 3'b100;
								assign node542 = (inp[4]) ? node560 : node543;
									assign node543 = (inp[6]) ? node553 : node544;
										assign node544 = (inp[1]) ? node546 : 3'b000;
											assign node546 = (inp[11]) ? node550 : node547;
												assign node547 = (inp[3]) ? 3'b000 : 3'b010;
												assign node550 = (inp[3]) ? 3'b010 : 3'b100;
										assign node553 = (inp[1]) ? node557 : node554;
											assign node554 = (inp[11]) ? 3'b000 : 3'b010;
											assign node557 = (inp[11]) ? 3'b010 : 3'b000;
									assign node560 = (inp[1]) ? node566 : node561;
										assign node561 = (inp[6]) ? node563 : 3'b100;
											assign node563 = (inp[11]) ? 3'b100 : 3'b010;
										assign node566 = (inp[11]) ? 3'b000 : 3'b010;
							assign node569 = (inp[11]) ? node597 : node570;
								assign node570 = (inp[6]) ? node588 : node571;
									assign node571 = (inp[3]) ? node581 : node572;
										assign node572 = (inp[4]) ? node578 : node573;
											assign node573 = (inp[1]) ? 3'b010 : node574;
												assign node574 = (inp[8]) ? 3'b010 : 3'b110;
											assign node578 = (inp[8]) ? 3'b010 : 3'b000;
										assign node581 = (inp[1]) ? 3'b100 : node582;
											assign node582 = (inp[4]) ? 3'b110 : node583;
												assign node583 = (inp[8]) ? 3'b010 : 3'b110;
									assign node588 = (inp[4]) ? node594 : node589;
										assign node589 = (inp[8]) ? node591 : 3'b100;
											assign node591 = (inp[1]) ? 3'b110 : 3'b000;
										assign node594 = (inp[3]) ? 3'b100 : 3'b000;
								assign node597 = (inp[3]) ? node605 : node598;
									assign node598 = (inp[1]) ? 3'b010 : node599;
										assign node599 = (inp[4]) ? 3'b010 : node600;
											assign node600 = (inp[8]) ? 3'b010 : 3'b110;
									assign node605 = (inp[1]) ? node611 : node606;
										assign node606 = (inp[4]) ? 3'b110 : node607;
											assign node607 = (inp[8]) ? 3'b010 : 3'b110;
										assign node611 = (inp[4]) ? 3'b010 : 3'b110;
						assign node614 = (inp[11]) ? node654 : node615;
							assign node615 = (inp[1]) ? node639 : node616;
								assign node616 = (inp[4]) ? node632 : node617;
									assign node617 = (inp[3]) ? node623 : node618;
										assign node618 = (inp[5]) ? 3'b100 : node619;
											assign node619 = (inp[8]) ? 3'b000 : 3'b100;
										assign node623 = (inp[8]) ? node629 : node624;
											assign node624 = (inp[6]) ? 3'b110 : node625;
												assign node625 = (inp[5]) ? 3'b010 : 3'b000;
											assign node629 = (inp[5]) ? 3'b110 : 3'b100;
									assign node632 = (inp[3]) ? 3'b000 : node633;
										assign node633 = (inp[5]) ? 3'b000 : node634;
											assign node634 = (inp[8]) ? 3'b100 : 3'b000;
								assign node639 = (inp[5]) ? 3'b000 : node640;
									assign node640 = (inp[4]) ? node648 : node641;
										assign node641 = (inp[3]) ? node645 : node642;
											assign node642 = (inp[6]) ? 3'b000 : 3'b010;
											assign node645 = (inp[6]) ? 3'b010 : 3'b000;
										assign node648 = (inp[6]) ? node650 : 3'b000;
											assign node650 = (inp[3]) ? 3'b010 : 3'b000;
							assign node654 = (inp[5]) ? node686 : node655;
								assign node655 = (inp[1]) ? node671 : node656;
									assign node656 = (inp[3]) ? node664 : node657;
										assign node657 = (inp[4]) ? node661 : node658;
											assign node658 = (inp[8]) ? 3'b010 : 3'b110;
											assign node661 = (inp[8]) ? 3'b110 : 3'b000;
										assign node664 = (inp[8]) ? node668 : node665;
											assign node665 = (inp[4]) ? 3'b010 : 3'b000;
											assign node668 = (inp[4]) ? 3'b000 : 3'b100;
									assign node671 = (inp[4]) ? 3'b000 : node672;
										assign node672 = (inp[6]) ? node680 : node673;
											assign node673 = (inp[3]) ? node677 : node674;
												assign node674 = (inp[8]) ? 3'b010 : 3'b000;
												assign node677 = (inp[8]) ? 3'b000 : 3'b010;
											assign node680 = (inp[8]) ? node682 : 3'b010;
												assign node682 = (inp[3]) ? 3'b000 : 3'b010;
								assign node686 = (inp[4]) ? node694 : node687;
									assign node687 = (inp[1]) ? 3'b010 : node688;
										assign node688 = (inp[8]) ? 3'b110 : node689;
											assign node689 = (inp[3]) ? 3'b010 : 3'b110;
									assign node694 = (inp[1]) ? 3'b000 : 3'b010;
				assign node697 = (inp[2]) ? node699 : 3'b010;
					assign node699 = (inp[1]) ? node727 : node700;
						assign node700 = (inp[7]) ? node702 : 3'b010;
							assign node702 = (inp[3]) ? 3'b010 : node703;
								assign node703 = (inp[8]) ? node715 : node704;
									assign node704 = (inp[5]) ? node710 : node705;
										assign node705 = (inp[11]) ? 3'b000 : node706;
											assign node706 = (inp[6]) ? 3'b010 : 3'b000;
										assign node710 = (inp[11]) ? 3'b010 : node711;
											assign node711 = (inp[6]) ? 3'b000 : 3'b010;
									assign node715 = (inp[4]) ? node717 : 3'b010;
										assign node717 = (inp[11]) ? node723 : node718;
											assign node718 = (inp[6]) ? node720 : 3'b010;
												assign node720 = (inp[5]) ? 3'b000 : 3'b010;
											assign node723 = (inp[5]) ? 3'b010 : 3'b000;
						assign node727 = (inp[3]) ? node775 : node728;
							assign node728 = (inp[7]) ? node760 : node729;
								assign node729 = (inp[8]) ? node745 : node730;
									assign node730 = (inp[4]) ? node742 : node731;
										assign node731 = (inp[5]) ? node737 : node732;
											assign node732 = (inp[6]) ? node734 : 3'b100;
												assign node734 = (inp[11]) ? 3'b100 : 3'b010;
											assign node737 = (inp[6]) ? node739 : 3'b110;
												assign node739 = (inp[11]) ? 3'b110 : 3'b100;
										assign node742 = (inp[11]) ? 3'b010 : 3'b000;
									assign node745 = (inp[5]) ? node753 : node746;
										assign node746 = (inp[11]) ? node750 : node747;
											assign node747 = (inp[6]) ? 3'b010 : 3'b000;
											assign node750 = (inp[4]) ? 3'b100 : 3'b000;
										assign node753 = (inp[11]) ? 3'b010 : node754;
											assign node754 = (inp[4]) ? 3'b000 : node755;
												assign node755 = (inp[6]) ? 3'b000 : 3'b010;
								assign node760 = (inp[4]) ? node768 : node761;
									assign node761 = (inp[5]) ? 3'b010 : node762;
										assign node762 = (inp[11]) ? 3'b000 : node763;
											assign node763 = (inp[8]) ? 3'b000 : 3'b010;
									assign node768 = (inp[6]) ? 3'b000 : node769;
										assign node769 = (inp[8]) ? 3'b000 : node770;
											assign node770 = (inp[5]) ? 3'b000 : 3'b010;
							assign node775 = (inp[7]) ? node777 : 3'b010;
								assign node777 = (inp[4]) ? node785 : node778;
									assign node778 = (inp[5]) ? 3'b010 : node779;
										assign node779 = (inp[11]) ? 3'b000 : node780;
											assign node780 = (inp[6]) ? 3'b010 : 3'b000;
									assign node785 = (inp[8]) ? node787 : 3'b000;
										assign node787 = (inp[5]) ? 3'b000 : node788;
											assign node788 = (inp[11]) ? 3'b000 : 3'b010;
		assign node792 = (inp[9]) ? node1174 : node793;
			assign node793 = (inp[2]) ? node915 : node794;
				assign node794 = (inp[0]) ? 3'b100 : node795;
					assign node795 = (inp[1]) ? node847 : node796;
						assign node796 = (inp[3]) ? 3'b101 : node797;
							assign node797 = (inp[7]) ? node819 : node798;
								assign node798 = (inp[4]) ? node808 : node799;
									assign node799 = (inp[5]) ? node801 : 3'b101;
										assign node801 = (inp[8]) ? 3'b101 : node802;
											assign node802 = (inp[11]) ? 3'b000 : node803;
												assign node803 = (inp[6]) ? 3'b101 : 3'b000;
									assign node808 = (inp[8]) ? node816 : node809;
										assign node809 = (inp[5]) ? node811 : 3'b010;
											assign node811 = (inp[6]) ? node813 : 3'b000;
												assign node813 = (inp[11]) ? 3'b000 : 3'b010;
										assign node816 = (inp[5]) ? 3'b000 : 3'b101;
								assign node819 = (inp[4]) ? node829 : node820;
									assign node820 = (inp[8]) ? 3'b000 : node821;
										assign node821 = (inp[11]) ? 3'b010 : node822;
											assign node822 = (inp[5]) ? 3'b010 : node823;
												assign node823 = (inp[6]) ? 3'b000 : 3'b010;
									assign node829 = (inp[8]) ? node839 : node830;
										assign node830 = (inp[5]) ? node834 : node831;
											assign node831 = (inp[11]) ? 3'b110 : 3'b100;
											assign node834 = (inp[11]) ? 3'b100 : node835;
												assign node835 = (inp[6]) ? 3'b110 : 3'b100;
										assign node839 = (inp[11]) ? 3'b100 : node840;
											assign node840 = (inp[5]) ? node842 : 3'b010;
												assign node842 = (inp[6]) ? 3'b010 : 3'b100;
						assign node847 = (inp[5]) ? node883 : node848;
							assign node848 = (inp[7]) ? node868 : node849;
								assign node849 = (inp[3]) ? node863 : node850;
									assign node850 = (inp[11]) ? node858 : node851;
										assign node851 = (inp[6]) ? node853 : 3'b110;
											assign node853 = (inp[8]) ? 3'b100 : node854;
												assign node854 = (inp[4]) ? 3'b000 : 3'b100;
										assign node858 = (inp[8]) ? 3'b110 : node859;
											assign node859 = (inp[4]) ? 3'b010 : 3'b110;
									assign node863 = (inp[8]) ? 3'b101 : node864;
										assign node864 = (inp[4]) ? 3'b010 : 3'b101;
								assign node868 = (inp[4]) ? node874 : node869;
									assign node869 = (inp[11]) ? 3'b010 : node870;
										assign node870 = (inp[6]) ? 3'b000 : 3'b010;
									assign node874 = (inp[8]) ? node880 : node875;
										assign node875 = (inp[3]) ? 3'b110 : node876;
											assign node876 = (inp[11]) ? 3'b110 : 3'b100;
										assign node880 = (inp[6]) ? 3'b000 : 3'b010;
							assign node883 = (inp[6]) ? node895 : node884;
								assign node884 = (inp[7]) ? node890 : node885;
									assign node885 = (inp[4]) ? 3'b000 : node886;
										assign node886 = (inp[8]) ? 3'b101 : 3'b000;
									assign node890 = (inp[4]) ? 3'b100 : node891;
										assign node891 = (inp[8]) ? 3'b000 : 3'b100;
								assign node895 = (inp[11]) ? node907 : node896;
									assign node896 = (inp[7]) ? node902 : node897;
										assign node897 = (inp[8]) ? node899 : 3'b010;
											assign node899 = (inp[3]) ? 3'b101 : 3'b110;
										assign node902 = (inp[4]) ? node904 : 3'b010;
											assign node904 = (inp[8]) ? 3'b010 : 3'b110;
									assign node907 = (inp[7]) ? node911 : node908;
										assign node908 = (inp[8]) ? 3'b100 : 3'b000;
										assign node911 = (inp[4]) ? 3'b100 : 3'b000;
				assign node915 = (inp[1]) ? node1035 : node916;
					assign node916 = (inp[0]) ? node1008 : node917;
						assign node917 = (inp[11]) ? node975 : node918;
							assign node918 = (inp[7]) ? node948 : node919;
								assign node919 = (inp[8]) ? node935 : node920;
									assign node920 = (inp[3]) ? node930 : node921;
										assign node921 = (inp[4]) ? node927 : node922;
											assign node922 = (inp[5]) ? 3'b010 : node923;
												assign node923 = (inp[6]) ? 3'b100 : 3'b110;
											assign node927 = (inp[5]) ? 3'b110 : 3'b010;
										assign node930 = (inp[6]) ? node932 : 3'b000;
											assign node932 = (inp[4]) ? 3'b010 : 3'b110;
									assign node935 = (inp[4]) ? node941 : node936;
										assign node936 = (inp[6]) ? 3'b100 : node937;
											assign node937 = (inp[5]) ? 3'b100 : 3'b110;
										assign node941 = (inp[3]) ? node943 : 3'b010;
											assign node943 = (inp[6]) ? node945 : 3'b110;
												assign node945 = (inp[5]) ? 3'b110 : 3'b100;
								assign node948 = (inp[3]) ? node966 : node949;
									assign node949 = (inp[4]) ? node955 : node950;
										assign node950 = (inp[5]) ? node952 : 3'b110;
											assign node952 = (inp[8]) ? 3'b110 : 3'b010;
										assign node955 = (inp[8]) ? node959 : node956;
											assign node956 = (inp[5]) ? 3'b100 : 3'b010;
											assign node959 = (inp[5]) ? node963 : node960;
												assign node960 = (inp[6]) ? 3'b010 : 3'b000;
												assign node963 = (inp[6]) ? 3'b000 : 3'b010;
									assign node966 = (inp[8]) ? node972 : node967;
										assign node967 = (inp[4]) ? node969 : 3'b010;
											assign node969 = (inp[5]) ? 3'b110 : 3'b010;
										assign node972 = (inp[4]) ? 3'b010 : 3'b000;
							assign node975 = (inp[5]) ? node995 : node976;
								assign node976 = (inp[3]) ? node986 : node977;
									assign node977 = (inp[7]) ? node983 : node978;
										assign node978 = (inp[6]) ? node980 : 3'b000;
											assign node980 = (inp[4]) ? 3'b100 : 3'b000;
										assign node983 = (inp[4]) ? 3'b010 : 3'b000;
									assign node986 = (inp[7]) ? node992 : node987;
										assign node987 = (inp[8]) ? 3'b110 : node988;
											assign node988 = (inp[4]) ? 3'b010 : 3'b110;
										assign node992 = (inp[6]) ? 3'b100 : 3'b000;
								assign node995 = (inp[4]) ? node1003 : node996;
									assign node996 = (inp[7]) ? 3'b000 : node997;
										assign node997 = (inp[8]) ? node999 : 3'b000;
											assign node999 = (inp[3]) ? 3'b100 : 3'b000;
									assign node1003 = (inp[3]) ? node1005 : 3'b100;
										assign node1005 = (inp[7]) ? 3'b100 : 3'b000;
						assign node1008 = (inp[3]) ? 3'b100 : node1009;
							assign node1009 = (inp[7]) ? node1019 : node1010;
								assign node1010 = (inp[8]) ? 3'b100 : node1011;
									assign node1011 = (inp[4]) ? node1015 : node1012;
										assign node1012 = (inp[5]) ? 3'b000 : 3'b100;
										assign node1015 = (inp[5]) ? 3'b000 : 3'b010;
								assign node1019 = (inp[5]) ? node1021 : 3'b010;
									assign node1021 = (inp[11]) ? node1029 : node1022;
										assign node1022 = (inp[6]) ? node1026 : node1023;
											assign node1023 = (inp[8]) ? 3'b000 : 3'b100;
											assign node1026 = (inp[4]) ? 3'b110 : 3'b010;
										assign node1029 = (inp[8]) ? node1031 : 3'b100;
											assign node1031 = (inp[4]) ? 3'b100 : 3'b000;
					assign node1035 = (inp[7]) ? node1123 : node1036;
						assign node1036 = (inp[4]) ? node1090 : node1037;
							assign node1037 = (inp[5]) ? node1059 : node1038;
								assign node1038 = (inp[8]) ? node1052 : node1039;
									assign node1039 = (inp[0]) ? node1047 : node1040;
										assign node1040 = (inp[3]) ? node1042 : 3'b000;
											assign node1042 = (inp[6]) ? node1044 : 3'b000;
												assign node1044 = (inp[11]) ? 3'b010 : 3'b110;
										assign node1047 = (inp[3]) ? 3'b100 : node1048;
											assign node1048 = (inp[11]) ? 3'b000 : 3'b100;
									assign node1052 = (inp[3]) ? node1054 : 3'b110;
										assign node1054 = (inp[0]) ? 3'b100 : node1055;
											assign node1055 = (inp[11]) ? 3'b100 : 3'b110;
								assign node1059 = (inp[11]) ? node1077 : node1060;
									assign node1060 = (inp[0]) ? node1070 : node1061;
										assign node1061 = (inp[8]) ? node1065 : node1062;
											assign node1062 = (inp[3]) ? 3'b000 : 3'b100;
											assign node1065 = (inp[3]) ? node1067 : 3'b000;
												assign node1067 = (inp[6]) ? 3'b000 : 3'b010;
										assign node1070 = (inp[8]) ? 3'b100 : node1071;
											assign node1071 = (inp[3]) ? node1073 : 3'b010;
												assign node1073 = (inp[6]) ? 3'b100 : 3'b000;
									assign node1077 = (inp[8]) ? node1083 : node1078;
										assign node1078 = (inp[3]) ? node1080 : 3'b000;
											assign node1080 = (inp[0]) ? 3'b000 : 3'b100;
										assign node1083 = (inp[3]) ? node1087 : node1084;
											assign node1084 = (inp[0]) ? 3'b000 : 3'b100;
											assign node1087 = (inp[0]) ? 3'b100 : 3'b000;
							assign node1090 = (inp[11]) ? node1110 : node1091;
								assign node1091 = (inp[3]) ? node1099 : node1092;
									assign node1092 = (inp[6]) ? node1094 : 3'b010;
										assign node1094 = (inp[5]) ? 3'b010 : node1095;
											assign node1095 = (inp[0]) ? 3'b010 : 3'b000;
									assign node1099 = (inp[5]) ? node1103 : node1100;
										assign node1100 = (inp[6]) ? 3'b010 : 3'b100;
										assign node1103 = (inp[6]) ? node1105 : 3'b000;
											assign node1105 = (inp[8]) ? node1107 : 3'b100;
												assign node1107 = (inp[0]) ? 3'b100 : 3'b000;
								assign node1110 = (inp[5]) ? 3'b000 : node1111;
									assign node1111 = (inp[0]) ? node1117 : node1112;
										assign node1112 = (inp[8]) ? node1114 : 3'b000;
											assign node1114 = (inp[3]) ? 3'b000 : 3'b010;
										assign node1117 = (inp[8]) ? 3'b100 : node1118;
											assign node1118 = (inp[3]) ? 3'b010 : 3'b100;
						assign node1123 = (inp[5]) ? node1161 : node1124;
							assign node1124 = (inp[4]) ? node1144 : node1125;
								assign node1125 = (inp[3]) ? node1137 : node1126;
									assign node1126 = (inp[8]) ? node1128 : 3'b000;
										assign node1128 = (inp[11]) ? node1134 : node1129;
											assign node1129 = (inp[0]) ? node1131 : 3'b000;
												assign node1131 = (inp[6]) ? 3'b010 : 3'b000;
											assign node1134 = (inp[0]) ? 3'b000 : 3'b010;
									assign node1137 = (inp[6]) ? node1139 : 3'b010;
										assign node1139 = (inp[0]) ? 3'b000 : node1140;
											assign node1140 = (inp[8]) ? 3'b000 : 3'b010;
								assign node1144 = (inp[11]) ? 3'b000 : node1145;
									assign node1145 = (inp[8]) ? node1153 : node1146;
										assign node1146 = (inp[6]) ? 3'b000 : node1147;
											assign node1147 = (inp[0]) ? node1149 : 3'b000;
												assign node1149 = (inp[3]) ? 3'b000 : 3'b010;
										assign node1153 = (inp[6]) ? node1155 : 3'b000;
											assign node1155 = (inp[3]) ? node1157 : 3'b010;
												assign node1157 = (inp[0]) ? 3'b010 : 3'b000;
							assign node1161 = (inp[11]) ? 3'b000 : node1162;
								assign node1162 = (inp[4]) ? 3'b000 : node1163;
									assign node1163 = (inp[0]) ? node1165 : 3'b000;
										assign node1165 = (inp[3]) ? 3'b010 : node1166;
											assign node1166 = (inp[8]) ? 3'b000 : node1167;
												assign node1167 = (inp[6]) ? 3'b010 : 3'b000;
			assign node1174 = (inp[0]) ? node1446 : node1175;
				assign node1175 = (inp[2]) ? node1259 : node1176;
					assign node1176 = (inp[3]) ? node1234 : node1177;
						assign node1177 = (inp[1]) ? node1195 : node1178;
							assign node1178 = (inp[7]) ? node1180 : 3'b001;
								assign node1180 = (inp[8]) ? node1188 : node1181;
									assign node1181 = (inp[5]) ? 3'b000 : node1182;
										assign node1182 = (inp[11]) ? 3'b010 : node1183;
											assign node1183 = (inp[4]) ? 3'b000 : 3'b001;
									assign node1188 = (inp[4]) ? node1190 : 3'b001;
										assign node1190 = (inp[5]) ? node1192 : 3'b001;
											assign node1192 = (inp[11]) ? 3'b000 : 3'b001;
							assign node1195 = (inp[5]) ? node1215 : node1196;
								assign node1196 = (inp[7]) ? node1208 : node1197;
									assign node1197 = (inp[8]) ? node1203 : node1198;
										assign node1198 = (inp[4]) ? node1200 : 3'b010;
											assign node1200 = (inp[6]) ? 3'b100 : 3'b110;
										assign node1203 = (inp[6]) ? node1205 : 3'b010;
											assign node1205 = (inp[11]) ? 3'b010 : 3'b000;
									assign node1208 = (inp[11]) ? 3'b110 : node1209;
										assign node1209 = (inp[6]) ? 3'b100 : node1210;
											assign node1210 = (inp[8]) ? 3'b110 : 3'b010;
								assign node1215 = (inp[11]) ? node1227 : node1216;
									assign node1216 = (inp[6]) ? node1222 : node1217;
										assign node1217 = (inp[7]) ? node1219 : 3'b100;
											assign node1219 = (inp[8]) ? 3'b100 : 3'b000;
										assign node1222 = (inp[7]) ? node1224 : 3'b010;
											assign node1224 = (inp[8]) ? 3'b110 : 3'b010;
									assign node1227 = (inp[7]) ? 3'b000 : node1228;
										assign node1228 = (inp[4]) ? 3'b100 : node1229;
											assign node1229 = (inp[8]) ? 3'b000 : 3'b100;
						assign node1234 = (inp[7]) ? node1236 : 3'b001;
							assign node1236 = (inp[1]) ? node1238 : 3'b001;
								assign node1238 = (inp[4]) ? node1246 : node1239;
									assign node1239 = (inp[8]) ? 3'b001 : node1240;
										assign node1240 = (inp[5]) ? node1242 : 3'b001;
											assign node1242 = (inp[11]) ? 3'b000 : 3'b001;
									assign node1246 = (inp[8]) ? node1252 : node1247;
										assign node1247 = (inp[11]) ? node1249 : 3'b010;
											assign node1249 = (inp[5]) ? 3'b000 : 3'b010;
										assign node1252 = (inp[5]) ? node1254 : 3'b001;
											assign node1254 = (inp[6]) ? node1256 : 3'b000;
												assign node1256 = (inp[11]) ? 3'b000 : 3'b001;
					assign node1259 = (inp[11]) ? node1377 : node1260;
						assign node1260 = (inp[1]) ? node1328 : node1261;
							assign node1261 = (inp[3]) ? node1295 : node1262;
								assign node1262 = (inp[7]) ? node1278 : node1263;
									assign node1263 = (inp[4]) ? node1271 : node1264;
										assign node1264 = (inp[5]) ? node1268 : node1265;
											assign node1265 = (inp[6]) ? 3'b000 : 3'b010;
											assign node1268 = (inp[6]) ? 3'b010 : 3'b000;
										assign node1271 = (inp[5]) ? 3'b010 : node1272;
											assign node1272 = (inp[8]) ? 3'b010 : node1273;
												assign node1273 = (inp[6]) ? 3'b100 : 3'b110;
									assign node1278 = (inp[6]) ? node1284 : node1279;
										assign node1279 = (inp[8]) ? 3'b010 : node1280;
											assign node1280 = (inp[4]) ? 3'b010 : 3'b110;
										assign node1284 = (inp[4]) ? node1290 : node1285;
											assign node1285 = (inp[5]) ? node1287 : 3'b010;
												assign node1287 = (inp[8]) ? 3'b010 : 3'b110;
											assign node1290 = (inp[5]) ? node1292 : 3'b110;
												assign node1292 = (inp[8]) ? 3'b110 : 3'b000;
								assign node1295 = (inp[6]) ? node1315 : node1296;
									assign node1296 = (inp[5]) ? node1306 : node1297;
										assign node1297 = (inp[7]) ? node1301 : node1298;
											assign node1298 = (inp[8]) ? 3'b010 : 3'b110;
											assign node1301 = (inp[8]) ? 3'b110 : node1302;
												assign node1302 = (inp[4]) ? 3'b010 : 3'b110;
										assign node1306 = (inp[7]) ? node1312 : node1307;
											assign node1307 = (inp[8]) ? node1309 : 3'b100;
												assign node1309 = (inp[4]) ? 3'b100 : 3'b000;
											assign node1312 = (inp[4]) ? 3'b010 : 3'b000;
									assign node1315 = (inp[5]) ? node1325 : node1316;
										assign node1316 = (inp[8]) ? 3'b100 : node1317;
											assign node1317 = (inp[7]) ? node1321 : node1318;
												assign node1318 = (inp[4]) ? 3'b100 : 3'b000;
												assign node1321 = (inp[4]) ? 3'b000 : 3'b100;
										assign node1325 = (inp[7]) ? 3'b110 : 3'b010;
							assign node1328 = (inp[4]) ? node1352 : node1329;
								assign node1329 = (inp[3]) ? node1343 : node1330;
									assign node1330 = (inp[7]) ? 3'b010 : node1331;
										assign node1331 = (inp[8]) ? node1337 : node1332;
											assign node1332 = (inp[6]) ? node1334 : 3'b100;
												assign node1334 = (inp[5]) ? 3'b000 : 3'b010;
											assign node1337 = (inp[5]) ? node1339 : 3'b000;
												assign node1339 = (inp[6]) ? 3'b100 : 3'b110;
									assign node1343 = (inp[7]) ? node1349 : node1344;
										assign node1344 = (inp[5]) ? node1346 : 3'b010;
											assign node1346 = (inp[8]) ? 3'b010 : 3'b110;
										assign node1349 = (inp[8]) ? 3'b000 : 3'b010;
								assign node1352 = (inp[7]) ? node1372 : node1353;
									assign node1353 = (inp[6]) ? node1361 : node1354;
										assign node1354 = (inp[8]) ? node1358 : node1355;
											assign node1355 = (inp[3]) ? 3'b000 : 3'b100;
											assign node1358 = (inp[3]) ? 3'b010 : 3'b000;
										assign node1361 = (inp[5]) ? node1369 : node1362;
											assign node1362 = (inp[3]) ? node1366 : node1363;
												assign node1363 = (inp[8]) ? 3'b000 : 3'b100;
												assign node1366 = (inp[8]) ? 3'b110 : 3'b010;
											assign node1369 = (inp[3]) ? 3'b000 : 3'b010;
									assign node1372 = (inp[3]) ? node1374 : 3'b000;
										assign node1374 = (inp[5]) ? 3'b000 : 3'b010;
						assign node1377 = (inp[5]) ? node1421 : node1378;
							assign node1378 = (inp[7]) ? node1404 : node1379;
								assign node1379 = (inp[1]) ? node1391 : node1380;
									assign node1380 = (inp[3]) ? node1386 : node1381;
										assign node1381 = (inp[8]) ? 3'b010 : node1382;
											assign node1382 = (inp[4]) ? 3'b000 : 3'b010;
										assign node1386 = (inp[8]) ? 3'b010 : node1387;
											assign node1387 = (inp[4]) ? 3'b110 : 3'b010;
									assign node1391 = (inp[8]) ? node1397 : node1392;
										assign node1392 = (inp[4]) ? 3'b010 : node1393;
											assign node1393 = (inp[3]) ? 3'b100 : 3'b110;
										assign node1397 = (inp[4]) ? node1401 : node1398;
											assign node1398 = (inp[3]) ? 3'b000 : 3'b010;
											assign node1401 = (inp[3]) ? 3'b010 : 3'b100;
								assign node1404 = (inp[3]) ? node1414 : node1405;
									assign node1405 = (inp[1]) ? 3'b000 : node1406;
										assign node1406 = (inp[8]) ? node1410 : node1407;
											assign node1407 = (inp[4]) ? 3'b000 : 3'b100;
											assign node1410 = (inp[4]) ? 3'b100 : 3'b000;
									assign node1414 = (inp[1]) ? node1416 : 3'b110;
										assign node1416 = (inp[8]) ? node1418 : 3'b000;
											assign node1418 = (inp[4]) ? 3'b000 : 3'b010;
							assign node1421 = (inp[1]) ? node1437 : node1422;
								assign node1422 = (inp[4]) ? node1432 : node1423;
									assign node1423 = (inp[8]) ? node1429 : node1424;
										assign node1424 = (inp[7]) ? node1426 : 3'b100;
											assign node1426 = (inp[3]) ? 3'b000 : 3'b100;
										assign node1429 = (inp[7]) ? 3'b100 : 3'b000;
									assign node1432 = (inp[7]) ? 3'b000 : node1433;
										assign node1433 = (inp[3]) ? 3'b100 : 3'b000;
								assign node1437 = (inp[8]) ? node1439 : 3'b000;
									assign node1439 = (inp[3]) ? node1441 : 3'b000;
										assign node1441 = (inp[7]) ? 3'b000 : node1442;
											assign node1442 = (inp[4]) ? 3'b000 : 3'b100;
				assign node1446 = (inp[3]) ? 3'b000 : node1447;
					assign node1447 = (inp[2]) ? node1449 : 3'b000;
						assign node1449 = (inp[1]) ? node1463 : node1450;
							assign node1450 = (inp[4]) ? node1452 : 3'b000;
								assign node1452 = (inp[8]) ? 3'b000 : node1453;
									assign node1453 = (inp[7]) ? node1455 : 3'b000;
										assign node1455 = (inp[5]) ? node1457 : 3'b010;
											assign node1457 = (inp[6]) ? node1459 : 3'b000;
												assign node1459 = (inp[11]) ? 3'b000 : 3'b010;
							assign node1463 = (inp[5]) ? node1487 : node1464;
								assign node1464 = (inp[4]) ? node1476 : node1465;
									assign node1465 = (inp[11]) ? 3'b010 : node1466;
										assign node1466 = (inp[7]) ? node1470 : node1467;
											assign node1467 = (inp[6]) ? 3'b000 : 3'b010;
											assign node1470 = (inp[6]) ? 3'b010 : node1471;
												assign node1471 = (inp[8]) ? 3'b010 : 3'b000;
									assign node1476 = (inp[8]) ? node1480 : node1477;
										assign node1477 = (inp[11]) ? 3'b000 : 3'b100;
										assign node1480 = (inp[7]) ? node1482 : 3'b010;
											assign node1482 = (inp[6]) ? 3'b000 : node1483;
												assign node1483 = (inp[11]) ? 3'b000 : 3'b010;
								assign node1487 = (inp[11]) ? node1503 : node1488;
									assign node1488 = (inp[7]) ? node1496 : node1489;
										assign node1489 = (inp[6]) ? 3'b010 : node1490;
											assign node1490 = (inp[8]) ? node1492 : 3'b010;
												assign node1492 = (inp[4]) ? 3'b100 : 3'b000;
										assign node1496 = (inp[6]) ? 3'b000 : node1497;
											assign node1497 = (inp[4]) ? 3'b000 : node1498;
												assign node1498 = (inp[8]) ? 3'b010 : 3'b000;
									assign node1503 = (inp[4]) ? 3'b000 : node1504;
										assign node1504 = (inp[8]) ? 3'b000 : node1505;
											assign node1505 = (inp[7]) ? 3'b000 : 3'b100;

endmodule