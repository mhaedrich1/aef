module dtc_split33_bm55 (
	input  wire [8-1:0] inp,
	output wire [7-1:0] outp
);

	wire [7-1:0] node1;
	wire [7-1:0] node2;
	wire [7-1:0] node3;
	wire [7-1:0] node4;
	wire [7-1:0] node5;
	wire [7-1:0] node6;
	wire [7-1:0] node11;
	wire [7-1:0] node12;
	wire [7-1:0] node14;
	wire [7-1:0] node18;
	wire [7-1:0] node19;
	wire [7-1:0] node20;
	wire [7-1:0] node21;
	wire [7-1:0] node22;
	wire [7-1:0] node25;
	wire [7-1:0] node29;
	wire [7-1:0] node32;
	wire [7-1:0] node34;
	wire [7-1:0] node36;
	wire [7-1:0] node39;
	wire [7-1:0] node40;
	wire [7-1:0] node41;
	wire [7-1:0] node43;
	wire [7-1:0] node46;
	wire [7-1:0] node47;
	wire [7-1:0] node48;
	wire [7-1:0] node51;
	wire [7-1:0] node54;
	wire [7-1:0] node55;
	wire [7-1:0] node57;
	wire [7-1:0] node61;
	wire [7-1:0] node62;
	wire [7-1:0] node63;
	wire [7-1:0] node66;
	wire [7-1:0] node67;
	wire [7-1:0] node69;
	wire [7-1:0] node73;
	wire [7-1:0] node75;
	wire [7-1:0] node77;
	wire [7-1:0] node80;
	wire [7-1:0] node81;
	wire [7-1:0] node82;
	wire [7-1:0] node83;
	wire [7-1:0] node84;
	wire [7-1:0] node85;
	wire [7-1:0] node89;
	wire [7-1:0] node91;
	wire [7-1:0] node94;
	wire [7-1:0] node95;
	wire [7-1:0] node96;
	wire [7-1:0] node98;
	wire [7-1:0] node102;
	wire [7-1:0] node105;
	wire [7-1:0] node106;
	wire [7-1:0] node107;
	wire [7-1:0] node109;
	wire [7-1:0] node112;
	wire [7-1:0] node113;
	wire [7-1:0] node117;
	wire [7-1:0] node119;
	wire [7-1:0] node120;
	wire [7-1:0] node123;
	wire [7-1:0] node126;
	wire [7-1:0] node127;
	wire [7-1:0] node128;
	wire [7-1:0] node129;
	wire [7-1:0] node132;
	wire [7-1:0] node135;
	wire [7-1:0] node136;
	wire [7-1:0] node139;
	wire [7-1:0] node140;
	wire [7-1:0] node144;
	wire [7-1:0] node145;
	wire [7-1:0] node146;
	wire [7-1:0] node149;
	wire [7-1:0] node152;
	wire [7-1:0] node153;

	assign outp = (inp[2]) ? node80 : node1;
		assign node1 = (inp[6]) ? node39 : node2;
			assign node2 = (inp[4]) ? node18 : node3;
				assign node3 = (inp[3]) ? node11 : node4;
					assign node4 = (inp[1]) ? 7'b1100100 : node5;
						assign node5 = (inp[0]) ? 7'b1110111 : node6;
							assign node6 = (inp[7]) ? 7'b0110111 : 7'b0110101;
					assign node11 = (inp[5]) ? 7'b0100100 : node12;
						assign node12 = (inp[7]) ? node14 : 7'b1111110;
							assign node14 = (inp[1]) ? 7'b1111101 : 7'b1111100;
				assign node18 = (inp[3]) ? node32 : node19;
					assign node19 = (inp[5]) ? node29 : node20;
						assign node20 = (inp[0]) ? 7'b0101110 : node21;
							assign node21 = (inp[1]) ? node25 : node22;
								assign node22 = (inp[7]) ? 7'b0011111 : 7'b0011101;
								assign node25 = (inp[7]) ? 7'b1000111 : 7'b0001100;
						assign node29 = (inp[7]) ? 7'b1000101 : 7'b1100100;
					assign node32 = (inp[7]) ? node34 : 7'b1010100;
						assign node34 = (inp[1]) ? node36 : 7'b1000101;
							assign node36 = (inp[5]) ? 7'b0000100 : 7'b1000100;
			assign node39 = (inp[0]) ? node61 : node40;
				assign node40 = (inp[7]) ? node46 : node41;
					assign node41 = (inp[3]) ? node43 : 7'b0001100;
						assign node43 = (inp[5]) ? 7'b1101000 : 7'b0101011;
					assign node46 = (inp[3]) ? node54 : node47;
						assign node47 = (inp[4]) ? node51 : node48;
							assign node48 = (inp[1]) ? 7'b1110001 : 7'b1010111;
							assign node51 = (inp[1]) ? 7'b0110011 : 7'b1101010;
						assign node54 = (inp[5]) ? 7'b0000100 : node55;
							assign node55 = (inp[4]) ? node57 : 7'b0111001;
								assign node57 = (inp[1]) ? 7'b0100000 : 7'b1110001;
				assign node61 = (inp[3]) ? node73 : node62;
					assign node62 = (inp[1]) ? node66 : node63;
						assign node63 = (inp[5]) ? 7'b1010001 : 7'b1110000;
						assign node66 = (inp[4]) ? 7'b0011000 : node67;
							assign node67 = (inp[5]) ? node69 : 7'b1011010;
								assign node69 = (inp[7]) ? 7'b1000000 : 7'b1011000;
					assign node73 = (inp[1]) ? node75 : 7'b0000001;
						assign node75 = (inp[4]) ? node77 : 7'b0011000;
							assign node77 = (inp[7]) ? 7'b0000000 : 7'b0010000;
		assign node80 = (inp[0]) ? node126 : node81;
			assign node81 = (inp[6]) ? node105 : node82;
				assign node82 = (inp[1]) ? node94 : node83;
					assign node83 = (inp[7]) ? node89 : node84;
						assign node84 = (inp[4]) ? 7'b1101011 : node85;
							assign node85 = (inp[5]) ? 7'b0111001 : 7'b0110011;
						assign node89 = (inp[5]) ? node91 : 7'b0110001;
							assign node91 = (inp[4]) ? 7'b1100001 : 7'b0100001;
					assign node94 = (inp[4]) ? node102 : node95;
						assign node95 = (inp[7]) ? 7'b0101010 : node96;
							assign node96 = (inp[3]) ? node98 : 7'b0110000;
								assign node98 = (inp[5]) ? 7'b1110000 : 7'b1111010;
						assign node102 = (inp[7]) ? 7'b1100000 : 7'b1101001;
				assign node105 = (inp[4]) ? node117 : node106;
					assign node106 = (inp[3]) ? node112 : node107;
						assign node107 = (inp[1]) ? node109 : 7'b1010001;
							assign node109 = (inp[5]) ? 7'b0011001 : 7'b1011011;
						assign node112 = (inp[7]) ? 7'b0000001 : node113;
							assign node113 = (inp[1]) ? 7'b1000001 : 7'b1000011;
					assign node117 = (inp[3]) ? node119 : 7'b0000001;
						assign node119 = (inp[1]) ? node123 : node120;
							assign node120 = (inp[7]) ? 7'b1010000 : 7'b1011000;
							assign node123 = (inp[7]) ? 7'b0000000 : 7'b1000010;
			assign node126 = (inp[5]) ? node144 : node127;
				assign node127 = (inp[6]) ? node135 : node128;
					assign node128 = (inp[7]) ? node132 : node129;
						assign node129 = (inp[4]) ? 7'b1001010 : 7'b0100010;
						assign node132 = (inp[4]) ? 7'b1000000 : 7'b1001001;
					assign node135 = (inp[4]) ? node139 : node136;
						assign node136 = (inp[1]) ? 7'b0010000 : 7'b0011000;
						assign node139 = (inp[1]) ? 7'b0000010 : node140;
							assign node140 = (inp[7]) ? 7'b0000000 : 7'b1001000;
				assign node144 = (inp[3]) ? node152 : node145;
					assign node145 = (inp[6]) ? node149 : node146;
						assign node146 = (inp[1]) ? 7'b0010000 : 7'b1010000;
						assign node149 = (inp[7]) ? 7'b1000000 : 7'b1001000;
					assign node152 = (inp[7]) ? 7'b0010001 : node153;
						assign node153 = (inp[1]) ? 7'b0000000 : 7'b0001000;

endmodule