module dtc_split5_bm49 (
	input  wire [7-1:0] inp,
	output wire [10-1:0] outp
);

	wire [10-1:0] node1;
	wire [10-1:0] node2;
	wire [10-1:0] node3;
	wire [10-1:0] node4;
	wire [10-1:0] node6;
	wire [10-1:0] node9;
	wire [10-1:0] node10;
	wire [10-1:0] node14;
	wire [10-1:0] node15;
	wire [10-1:0] node17;
	wire [10-1:0] node20;
	wire [10-1:0] node21;
	wire [10-1:0] node23;
	wire [10-1:0] node26;
	wire [10-1:0] node29;
	wire [10-1:0] node30;
	wire [10-1:0] node31;
	wire [10-1:0] node32;
	wire [10-1:0] node33;
	wire [10-1:0] node36;
	wire [10-1:0] node39;
	wire [10-1:0] node41;
	wire [10-1:0] node44;
	wire [10-1:0] node46;
	wire [10-1:0] node49;
	wire [10-1:0] node50;
	wire [10-1:0] node51;
	wire [10-1:0] node54;
	wire [10-1:0] node57;
	wire [10-1:0] node58;
	wire [10-1:0] node61;
	wire [10-1:0] node64;
	wire [10-1:0] node65;
	wire [10-1:0] node66;
	wire [10-1:0] node67;
	wire [10-1:0] node70;
	wire [10-1:0] node71;
	wire [10-1:0] node74;
	wire [10-1:0] node75;
	wire [10-1:0] node78;
	wire [10-1:0] node81;
	wire [10-1:0] node82;
	wire [10-1:0] node83;
	wire [10-1:0] node86;
	wire [10-1:0] node89;
	wire [10-1:0] node90;
	wire [10-1:0] node93;
	wire [10-1:0] node96;
	wire [10-1:0] node97;
	wire [10-1:0] node98;
	wire [10-1:0] node99;
	wire [10-1:0] node103;
	wire [10-1:0] node104;
	wire [10-1:0] node105;
	wire [10-1:0] node110;
	wire [10-1:0] node111;
	wire [10-1:0] node112;
	wire [10-1:0] node113;
	wire [10-1:0] node116;
	wire [10-1:0] node119;
	wire [10-1:0] node122;
	wire [10-1:0] node124;

	assign outp = (inp[3]) ? node64 : node1;
		assign node1 = (inp[1]) ? node29 : node2;
			assign node2 = (inp[0]) ? node14 : node3;
				assign node3 = (inp[4]) ? node9 : node4;
					assign node4 = (inp[6]) ? node6 : 10'b1101000010;
						assign node6 = (inp[2]) ? 10'b1000011110 : 10'b1100001111;
					assign node9 = (inp[6]) ? 10'b1000010000 : node10;
						assign node10 = (inp[2]) ? 10'b1001000000 : 10'b1001010001;
				assign node14 = (inp[2]) ? node20 : node15;
					assign node15 = (inp[5]) ? node17 : 10'b0001000011;
						assign node17 = (inp[6]) ? 10'b0000010011 : 10'b0100001011;
					assign node20 = (inp[4]) ? node26 : node21;
						assign node21 = (inp[6]) ? node23 : 10'b0101000000;
							assign node23 = (inp[5]) ? 10'b0100010000 : 10'b0000011100;
						assign node26 = (inp[6]) ? 10'b0100000110 : 10'b0100011110;
			assign node29 = (inp[0]) ? node49 : node30;
				assign node30 = (inp[2]) ? node44 : node31;
					assign node31 = (inp[6]) ? node39 : node32;
						assign node32 = (inp[4]) ? node36 : node33;
							assign node33 = (inp[5]) ? 10'b0000110110 : 10'b0101110010;
							assign node36 = (inp[5]) ? 10'b0100111000 : 10'b0001110000;
						assign node39 = (inp[5]) ? node41 : 10'b0000101100;
							assign node41 = (inp[4]) ? 10'b0100100000 : 10'b0000101010;
					assign node44 = (inp[6]) ? node46 : 10'b0000100101;
						assign node46 = (inp[5]) ? 10'b0100110001 : 10'b0000111101;
				assign node49 = (inp[4]) ? node57 : node50;
					assign node50 = (inp[2]) ? node54 : node51;
						assign node51 = (inp[6]) ? 10'b1100110011 : 10'b1101100011;
						assign node54 = (inp[6]) ? 10'b1100100010 : 10'b1100111010;
					assign node57 = (inp[5]) ? node61 : node58;
						assign node58 = (inp[6]) ? 10'b1100100100 : 10'b1100111100;
						assign node61 = (inp[6]) ? 10'b1000100000 : 10'b1000111000;
		assign node64 = (inp[1]) ? node96 : node65;
			assign node65 = (inp[2]) ? node81 : node66;
				assign node66 = (inp[6]) ? node70 : node67;
					assign node67 = (inp[0]) ? 10'b0111110000 : 10'b1111110010;
					assign node70 = (inp[0]) ? node74 : node71;
						assign node71 = (inp[5]) ? 10'b1110100000 : 10'b1010101100;
						assign node74 = (inp[4]) ? node78 : node75;
							assign node75 = (inp[5]) ? 10'b0010101000 : 10'b0110101100;
							assign node78 = (inp[5]) ? 10'b0010110010 : 10'b0110110110;
				assign node81 = (inp[0]) ? node89 : node82;
					assign node82 = (inp[6]) ? node86 : node83;
						assign node83 = (inp[5]) ? 10'b1010111011 : 10'b1110111111;
						assign node86 = (inp[4]) ? 10'b1010100011 : 10'b1110110001;
					assign node89 = (inp[6]) ? node93 : node90;
						assign node90 = (inp[4]) ? 10'b0010111001 : 10'b0011110011;
						assign node93 = (inp[5]) ? 10'b0110100011 : 10'b0010101111;
			assign node96 = (inp[0]) ? node110 : node97;
				assign node97 = (inp[4]) ? node103 : node98;
					assign node98 = (inp[6]) ? 10'b1110001101 : node99;
						assign node99 = (inp[2]) ? 10'b1111000000 : 10'b1111010001;
					assign node103 = (inp[2]) ? 10'b1010000010 : node104;
						assign node104 = (inp[6]) ? 10'b1110010111 : node105;
							assign node105 = (inp[5]) ? 10'b1110001011 : 10'b1011000011;
				assign node110 = (inp[4]) ? node122 : node111;
					assign node111 = (inp[6]) ? node119 : node112;
						assign node112 = (inp[2]) ? node116 : node113;
							assign node113 = (inp[5]) ? 10'b0010000111 : 10'b0111000011;
							assign node116 = (inp[5]) ? 10'b0110011010 : 10'b0011010010;
						assign node119 = (inp[2]) ? 10'b0010001110 : 10'b0010011111;
					assign node122 = (inp[6]) ? node124 : 10'b0110001001;
						assign node124 = (inp[2]) ? 10'b0110000100 : 10'b0110010101;

endmodule