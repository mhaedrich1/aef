module dtc_split25_bm22 (
	input  wire [11-1:0] inp,
	output wire [11-1:0] outp
);

	wire [11-1:0] node1;
	wire [11-1:0] node2;
	wire [11-1:0] node3;
	wire [11-1:0] node4;
	wire [11-1:0] node5;
	wire [11-1:0] node6;
	wire [11-1:0] node7;
	wire [11-1:0] node11;
	wire [11-1:0] node12;
	wire [11-1:0] node14;
	wire [11-1:0] node15;
	wire [11-1:0] node16;
	wire [11-1:0] node21;
	wire [11-1:0] node22;
	wire [11-1:0] node26;
	wire [11-1:0] node27;
	wire [11-1:0] node28;
	wire [11-1:0] node29;
	wire [11-1:0] node32;
	wire [11-1:0] node34;
	wire [11-1:0] node38;
	wire [11-1:0] node39;
	wire [11-1:0] node40;
	wire [11-1:0] node44;
	wire [11-1:0] node46;
	wire [11-1:0] node49;
	wire [11-1:0] node50;
	wire [11-1:0] node51;
	wire [11-1:0] node53;
	wire [11-1:0] node55;
	wire [11-1:0] node58;
	wire [11-1:0] node60;
	wire [11-1:0] node61;
	wire [11-1:0] node62;
	wire [11-1:0] node67;
	wire [11-1:0] node68;
	wire [11-1:0] node69;
	wire [11-1:0] node71;
	wire [11-1:0] node74;
	wire [11-1:0] node75;
	wire [11-1:0] node79;
	wire [11-1:0] node81;
	wire [11-1:0] node82;
	wire [11-1:0] node85;
	wire [11-1:0] node88;
	wire [11-1:0] node89;
	wire [11-1:0] node90;
	wire [11-1:0] node91;
	wire [11-1:0] node92;
	wire [11-1:0] node94;
	wire [11-1:0] node98;
	wire [11-1:0] node99;
	wire [11-1:0] node100;
	wire [11-1:0] node103;
	wire [11-1:0] node105;
	wire [11-1:0] node108;
	wire [11-1:0] node109;
	wire [11-1:0] node111;
	wire [11-1:0] node115;
	wire [11-1:0] node116;
	wire [11-1:0] node117;
	wire [11-1:0] node120;
	wire [11-1:0] node121;
	wire [11-1:0] node125;
	wire [11-1:0] node127;
	wire [11-1:0] node130;
	wire [11-1:0] node131;
	wire [11-1:0] node132;
	wire [11-1:0] node134;
	wire [11-1:0] node135;
	wire [11-1:0] node136;
	wire [11-1:0] node138;
	wire [11-1:0] node142;
	wire [11-1:0] node144;
	wire [11-1:0] node147;
	wire [11-1:0] node148;
	wire [11-1:0] node149;
	wire [11-1:0] node153;
	wire [11-1:0] node154;
	wire [11-1:0] node158;
	wire [11-1:0] node159;
	wire [11-1:0] node160;
	wire [11-1:0] node161;
	wire [11-1:0] node162;
	wire [11-1:0] node166;
	wire [11-1:0] node169;
	wire [11-1:0] node172;
	wire [11-1:0] node174;
	wire [11-1:0] node175;
	wire [11-1:0] node179;
	wire [11-1:0] node180;
	wire [11-1:0] node181;
	wire [11-1:0] node182;
	wire [11-1:0] node183;
	wire [11-1:0] node184;
	wire [11-1:0] node187;
	wire [11-1:0] node188;
	wire [11-1:0] node192;
	wire [11-1:0] node193;
	wire [11-1:0] node194;
	wire [11-1:0] node196;
	wire [11-1:0] node199;
	wire [11-1:0] node202;
	wire [11-1:0] node203;
	wire [11-1:0] node205;
	wire [11-1:0] node208;
	wire [11-1:0] node211;
	wire [11-1:0] node212;
	wire [11-1:0] node213;
	wire [11-1:0] node214;
	wire [11-1:0] node217;
	wire [11-1:0] node219;
	wire [11-1:0] node222;
	wire [11-1:0] node223;
	wire [11-1:0] node226;
	wire [11-1:0] node229;
	wire [11-1:0] node230;
	wire [11-1:0] node232;
	wire [11-1:0] node235;
	wire [11-1:0] node236;
	wire [11-1:0] node239;
	wire [11-1:0] node240;
	wire [11-1:0] node242;
	wire [11-1:0] node246;
	wire [11-1:0] node247;
	wire [11-1:0] node248;
	wire [11-1:0] node249;
	wire [11-1:0] node253;
	wire [11-1:0] node254;
	wire [11-1:0] node255;
	wire [11-1:0] node258;
	wire [11-1:0] node260;
	wire [11-1:0] node263;
	wire [11-1:0] node266;
	wire [11-1:0] node267;
	wire [11-1:0] node268;
	wire [11-1:0] node269;
	wire [11-1:0] node272;
	wire [11-1:0] node275;
	wire [11-1:0] node277;
	wire [11-1:0] node280;
	wire [11-1:0] node281;
	wire [11-1:0] node285;
	wire [11-1:0] node286;
	wire [11-1:0] node287;
	wire [11-1:0] node288;
	wire [11-1:0] node289;
	wire [11-1:0] node292;
	wire [11-1:0] node293;
	wire [11-1:0] node295;
	wire [11-1:0] node299;
	wire [11-1:0] node300;
	wire [11-1:0] node303;
	wire [11-1:0] node304;
	wire [11-1:0] node308;
	wire [11-1:0] node309;
	wire [11-1:0] node310;
	wire [11-1:0] node311;
	wire [11-1:0] node313;
	wire [11-1:0] node316;
	wire [11-1:0] node318;
	wire [11-1:0] node321;
	wire [11-1:0] node322;
	wire [11-1:0] node326;
	wire [11-1:0] node327;
	wire [11-1:0] node328;
	wire [11-1:0] node332;
	wire [11-1:0] node333;
	wire [11-1:0] node334;
	wire [11-1:0] node336;
	wire [11-1:0] node341;
	wire [11-1:0] node342;
	wire [11-1:0] node343;
	wire [11-1:0] node344;
	wire [11-1:0] node347;
	wire [11-1:0] node348;
	wire [11-1:0] node352;
	wire [11-1:0] node353;
	wire [11-1:0] node355;
	wire [11-1:0] node358;
	wire [11-1:0] node359;
	wire [11-1:0] node363;
	wire [11-1:0] node364;
	wire [11-1:0] node365;
	wire [11-1:0] node368;
	wire [11-1:0] node370;
	wire [11-1:0] node371;
	wire [11-1:0] node373;
	wire [11-1:0] node377;
	wire [11-1:0] node378;
	wire [11-1:0] node382;
	wire [11-1:0] node383;
	wire [11-1:0] node384;
	wire [11-1:0] node385;
	wire [11-1:0] node386;
	wire [11-1:0] node387;
	wire [11-1:0] node388;
	wire [11-1:0] node390;
	wire [11-1:0] node393;
	wire [11-1:0] node394;
	wire [11-1:0] node395;
	wire [11-1:0] node397;
	wire [11-1:0] node402;
	wire [11-1:0] node403;
	wire [11-1:0] node404;
	wire [11-1:0] node408;
	wire [11-1:0] node409;
	wire [11-1:0] node413;
	wire [11-1:0] node414;
	wire [11-1:0] node415;
	wire [11-1:0] node416;
	wire [11-1:0] node417;
	wire [11-1:0] node421;
	wire [11-1:0] node423;
	wire [11-1:0] node425;
	wire [11-1:0] node429;
	wire [11-1:0] node431;
	wire [11-1:0] node432;
	wire [11-1:0] node436;
	wire [11-1:0] node437;
	wire [11-1:0] node438;
	wire [11-1:0] node439;
	wire [11-1:0] node440;
	wire [11-1:0] node443;
	wire [11-1:0] node444;
	wire [11-1:0] node446;
	wire [11-1:0] node450;
	wire [11-1:0] node451;
	wire [11-1:0] node455;
	wire [11-1:0] node456;
	wire [11-1:0] node458;
	wire [11-1:0] node459;
	wire [11-1:0] node463;
	wire [11-1:0] node464;
	wire [11-1:0] node468;
	wire [11-1:0] node469;
	wire [11-1:0] node470;
	wire [11-1:0] node472;
	wire [11-1:0] node473;
	wire [11-1:0] node477;
	wire [11-1:0] node480;
	wire [11-1:0] node483;
	wire [11-1:0] node484;
	wire [11-1:0] node485;
	wire [11-1:0] node486;
	wire [11-1:0] node487;
	wire [11-1:0] node488;
	wire [11-1:0] node489;
	wire [11-1:0] node491;
	wire [11-1:0] node495;
	wire [11-1:0] node496;
	wire [11-1:0] node498;
	wire [11-1:0] node502;
	wire [11-1:0] node505;
	wire [11-1:0] node506;
	wire [11-1:0] node508;
	wire [11-1:0] node512;
	wire [11-1:0] node513;
	wire [11-1:0] node514;
	wire [11-1:0] node517;
	wire [11-1:0] node518;
	wire [11-1:0] node521;
	wire [11-1:0] node524;
	wire [11-1:0] node525;
	wire [11-1:0] node527;
	wire [11-1:0] node530;
	wire [11-1:0] node532;
	wire [11-1:0] node535;
	wire [11-1:0] node536;
	wire [11-1:0] node537;
	wire [11-1:0] node538;
	wire [11-1:0] node542;
	wire [11-1:0] node543;
	wire [11-1:0] node545;
	wire [11-1:0] node547;
	wire [11-1:0] node548;
	wire [11-1:0] node552;
	wire [11-1:0] node553;
	wire [11-1:0] node554;
	wire [11-1:0] node559;
	wire [11-1:0] node560;
	wire [11-1:0] node562;
	wire [11-1:0] node564;
	wire [11-1:0] node567;
	wire [11-1:0] node568;
	wire [11-1:0] node570;
	wire [11-1:0] node573;
	wire [11-1:0] node575;
	wire [11-1:0] node576;
	wire [11-1:0] node578;
	wire [11-1:0] node582;
	wire [11-1:0] node583;
	wire [11-1:0] node584;
	wire [11-1:0] node585;
	wire [11-1:0] node586;
	wire [11-1:0] node587;
	wire [11-1:0] node588;
	wire [11-1:0] node589;
	wire [11-1:0] node593;
	wire [11-1:0] node597;
	wire [11-1:0] node598;
	wire [11-1:0] node599;
	wire [11-1:0] node604;
	wire [11-1:0] node605;
	wire [11-1:0] node606;
	wire [11-1:0] node609;
	wire [11-1:0] node610;
	wire [11-1:0] node614;
	wire [11-1:0] node615;
	wire [11-1:0] node616;
	wire [11-1:0] node619;
	wire [11-1:0] node621;
	wire [11-1:0] node622;
	wire [11-1:0] node626;
	wire [11-1:0] node629;
	wire [11-1:0] node630;
	wire [11-1:0] node631;
	wire [11-1:0] node632;
	wire [11-1:0] node634;
	wire [11-1:0] node638;
	wire [11-1:0] node640;
	wire [11-1:0] node641;
	wire [11-1:0] node643;
	wire [11-1:0] node647;
	wire [11-1:0] node648;
	wire [11-1:0] node649;
	wire [11-1:0] node652;
	wire [11-1:0] node653;
	wire [11-1:0] node656;
	wire [11-1:0] node658;
	wire [11-1:0] node661;
	wire [11-1:0] node662;
	wire [11-1:0] node663;
	wire [11-1:0] node666;
	wire [11-1:0] node669;
	wire [11-1:0] node671;
	wire [11-1:0] node672;
	wire [11-1:0] node676;
	wire [11-1:0] node677;
	wire [11-1:0] node678;
	wire [11-1:0] node679;
	wire [11-1:0] node680;
	wire [11-1:0] node682;
	wire [11-1:0] node684;
	wire [11-1:0] node687;
	wire [11-1:0] node689;
	wire [11-1:0] node692;
	wire [11-1:0] node693;
	wire [11-1:0] node696;
	wire [11-1:0] node698;
	wire [11-1:0] node700;
	wire [11-1:0] node703;
	wire [11-1:0] node704;
	wire [11-1:0] node707;
	wire [11-1:0] node708;
	wire [11-1:0] node709;
	wire [11-1:0] node713;
	wire [11-1:0] node714;
	wire [11-1:0] node715;
	wire [11-1:0] node720;
	wire [11-1:0] node721;
	wire [11-1:0] node722;
	wire [11-1:0] node723;
	wire [11-1:0] node724;
	wire [11-1:0] node725;
	wire [11-1:0] node730;
	wire [11-1:0] node731;
	wire [11-1:0] node735;
	wire [11-1:0] node736;
	wire [11-1:0] node737;
	wire [11-1:0] node741;
	wire [11-1:0] node744;
	wire [11-1:0] node745;
	wire [11-1:0] node746;
	wire [11-1:0] node747;
	wire [11-1:0] node751;
	wire [11-1:0] node754;
	wire [11-1:0] node755;
	wire [11-1:0] node757;
	wire [11-1:0] node759;
	wire [11-1:0] node762;
	wire [11-1:0] node763;
	wire [11-1:0] node765;
	wire [11-1:0] node768;
	wire [11-1:0] node769;

	assign outp = (inp[5]) ? node382 : node1;
		assign node1 = (inp[1]) ? node179 : node2;
			assign node2 = (inp[8]) ? node88 : node3;
				assign node3 = (inp[6]) ? node49 : node4;
					assign node4 = (inp[10]) ? node26 : node5;
						assign node5 = (inp[0]) ? node11 : node6;
							assign node6 = (inp[9]) ? 11'b00111111111 : node7;
								assign node7 = (inp[2]) ? 11'b00111111111 : 11'b01111111111;
							assign node11 = (inp[4]) ? node21 : node12;
								assign node12 = (inp[3]) ? node14 : 11'b00111111111;
									assign node14 = (inp[7]) ? 11'b00011111111 : node15;
										assign node15 = (inp[2]) ? 11'b00011111111 : node16;
											assign node16 = (inp[9]) ? 11'b00011111111 : 11'b00111111111;
								assign node21 = (inp[9]) ? 11'b00000111111 : node22;
									assign node22 = (inp[3]) ? 11'b00001111111 : 11'b00011111111;
						assign node26 = (inp[9]) ? node38 : node27;
							assign node27 = (inp[2]) ? 11'b00001111111 : node28;
								assign node28 = (inp[4]) ? node32 : node29;
									assign node29 = (inp[7]) ? 11'b00011111111 : 11'b00111111111;
									assign node32 = (inp[3]) ? node34 : 11'b00011111111;
										assign node34 = (inp[7]) ? 11'b00001111111 : 11'b00011111111;
							assign node38 = (inp[3]) ? node44 : node39;
								assign node39 = (inp[7]) ? 11'b00001111111 : node40;
									assign node40 = (inp[4]) ? 11'b00001111111 : 11'b00011111111;
								assign node44 = (inp[2]) ? node46 : 11'b00001111111;
									assign node46 = (inp[7]) ? 11'b00000011111 : 11'b00000111111;
					assign node49 = (inp[3]) ? node67 : node50;
						assign node50 = (inp[10]) ? node58 : node51;
							assign node51 = (inp[4]) ? node53 : 11'b00111111111;
								assign node53 = (inp[7]) ? node55 : 11'b00011111111;
									assign node55 = (inp[2]) ? 11'b00001111111 : 11'b00011111111;
							assign node58 = (inp[0]) ? node60 : 11'b00001111111;
								assign node60 = (inp[7]) ? 11'b00001111111 : node61;
									assign node61 = (inp[9]) ? 11'b00001111111 : node62;
										assign node62 = (inp[4]) ? 11'b00001111111 : 11'b00011111111;
						assign node67 = (inp[4]) ? node79 : node68;
							assign node68 = (inp[2]) ? node74 : node69;
								assign node69 = (inp[9]) ? node71 : 11'b00001111111;
									assign node71 = (inp[10]) ? 11'b00000011111 : 11'b00001111111;
								assign node74 = (inp[7]) ? 11'b00000111111 : node75;
									assign node75 = (inp[10]) ? 11'b00000111111 : 11'b00001111111;
							assign node79 = (inp[9]) ? node81 : 11'b00000111111;
								assign node81 = (inp[10]) ? node85 : node82;
									assign node82 = (inp[2]) ? 11'b00000011111 : 11'b00000111111;
									assign node85 = (inp[0]) ? 11'b00000001111 : 11'b00000011111;
				assign node88 = (inp[0]) ? node130 : node89;
					assign node89 = (inp[9]) ? node115 : node90;
						assign node90 = (inp[7]) ? node98 : node91;
							assign node91 = (inp[4]) ? 11'b00001111111 : node92;
								assign node92 = (inp[6]) ? node94 : 11'b00111111111;
									assign node94 = (inp[3]) ? 11'b00000111111 : 11'b00011111111;
							assign node98 = (inp[2]) ? node108 : node99;
								assign node99 = (inp[3]) ? node103 : node100;
									assign node100 = (inp[6]) ? 11'b00001111111 : 11'b00011111111;
									assign node103 = (inp[6]) ? node105 : 11'b00001111111;
										assign node105 = (inp[4]) ? 11'b00000111111 : 11'b00001111111;
								assign node108 = (inp[6]) ? 11'b00000111111 : node109;
									assign node109 = (inp[10]) ? node111 : 11'b00001111111;
										assign node111 = (inp[4]) ? 11'b00000111111 : 11'b00001111111;
						assign node115 = (inp[7]) ? node125 : node116;
							assign node116 = (inp[3]) ? node120 : node117;
								assign node117 = (inp[10]) ? 11'b00001111111 : 11'b00000111111;
								assign node120 = (inp[4]) ? 11'b00000011111 : node121;
									assign node121 = (inp[2]) ? 11'b00000111111 : 11'b00001111111;
							assign node125 = (inp[4]) ? node127 : 11'b00000111111;
								assign node127 = (inp[3]) ? 11'b00000001111 : 11'b00000011111;
					assign node130 = (inp[10]) ? node158 : node131;
						assign node131 = (inp[6]) ? node147 : node132;
							assign node132 = (inp[9]) ? node134 : 11'b00001111111;
								assign node134 = (inp[3]) ? node142 : node135;
									assign node135 = (inp[4]) ? 11'b00000111111 : node136;
										assign node136 = (inp[7]) ? node138 : 11'b00001111111;
											assign node138 = (inp[2]) ? 11'b00000111111 : 11'b00001111111;
									assign node142 = (inp[4]) ? node144 : 11'b00000111111;
										assign node144 = (inp[7]) ? 11'b00000011111 : 11'b00000111111;
							assign node147 = (inp[2]) ? node153 : node148;
								assign node148 = (inp[7]) ? 11'b00000111111 : node149;
									assign node149 = (inp[3]) ? 11'b00000111111 : 11'b00001111111;
								assign node153 = (inp[9]) ? 11'b00000011111 : node154;
									assign node154 = (inp[3]) ? 11'b00000011111 : 11'b00000111111;
						assign node158 = (inp[3]) ? node172 : node159;
							assign node159 = (inp[2]) ? node169 : node160;
								assign node160 = (inp[4]) ? node166 : node161;
									assign node161 = (inp[9]) ? 11'b00000111111 : node162;
										assign node162 = (inp[6]) ? 11'b00001111111 : 11'b00011111111;
									assign node166 = (inp[9]) ? 11'b00000011111 : 11'b00000111111;
								assign node169 = (inp[9]) ? 11'b00000001111 : 11'b00000011111;
							assign node172 = (inp[4]) ? node174 : 11'b00000011111;
								assign node174 = (inp[9]) ? 11'b00000001111 : node175;
									assign node175 = (inp[6]) ? 11'b00000001111 : 11'b00000011111;
			assign node179 = (inp[3]) ? node285 : node180;
				assign node180 = (inp[9]) ? node246 : node181;
					assign node181 = (inp[2]) ? node211 : node182;
						assign node182 = (inp[7]) ? node192 : node183;
							assign node183 = (inp[10]) ? node187 : node184;
								assign node184 = (inp[8]) ? 11'b00111111111 : 11'b00011111111;
								assign node187 = (inp[4]) ? 11'b00001111111 : node188;
									assign node188 = (inp[0]) ? 11'b00001111111 : 11'b00011111111;
							assign node192 = (inp[6]) ? node202 : node193;
								assign node193 = (inp[0]) ? node199 : node194;
									assign node194 = (inp[4]) ? node196 : 11'b00011111111;
										assign node196 = (inp[8]) ? 11'b00001111111 : 11'b00011111111;
									assign node199 = (inp[10]) ? 11'b00000111111 : 11'b00001111111;
								assign node202 = (inp[4]) ? node208 : node203;
									assign node203 = (inp[8]) ? node205 : 11'b00001111111;
										assign node205 = (inp[10]) ? 11'b00000111111 : 11'b00001111111;
									assign node208 = (inp[10]) ? 11'b00000011111 : 11'b00000111111;
						assign node211 = (inp[0]) ? node229 : node212;
							assign node212 = (inp[4]) ? node222 : node213;
								assign node213 = (inp[7]) ? node217 : node214;
									assign node214 = (inp[6]) ? 11'b00001111111 : 11'b00011111111;
									assign node217 = (inp[10]) ? node219 : 11'b00001111111;
										assign node219 = (inp[8]) ? 11'b00000111111 : 11'b00001111111;
								assign node222 = (inp[6]) ? node226 : node223;
									assign node223 = (inp[8]) ? 11'b00000111111 : 11'b00001111111;
									assign node226 = (inp[10]) ? 11'b00000011111 : 11'b00000111111;
							assign node229 = (inp[10]) ? node235 : node230;
								assign node230 = (inp[4]) ? node232 : 11'b00001111111;
									assign node232 = (inp[7]) ? 11'b00000011111 : 11'b00000111111;
								assign node235 = (inp[4]) ? node239 : node236;
									assign node236 = (inp[8]) ? 11'b00000011111 : 11'b00000111111;
									assign node239 = (inp[7]) ? 11'b00000001111 : node240;
										assign node240 = (inp[8]) ? node242 : 11'b00000011111;
											assign node242 = (inp[6]) ? 11'b00000001111 : 11'b00000011111;
					assign node246 = (inp[6]) ? node266 : node247;
						assign node247 = (inp[8]) ? node253 : node248;
							assign node248 = (inp[0]) ? 11'b00000111111 : node249;
								assign node249 = (inp[4]) ? 11'b00000111111 : 11'b00001111111;
							assign node253 = (inp[2]) ? node263 : node254;
								assign node254 = (inp[4]) ? node258 : node255;
									assign node255 = (inp[7]) ? 11'b00000111111 : 11'b00001111111;
									assign node258 = (inp[10]) ? node260 : 11'b00000111111;
										assign node260 = (inp[7]) ? 11'b00000011111 : 11'b00000111111;
								assign node263 = (inp[10]) ? 11'b00000001111 : 11'b00000011111;
						assign node266 = (inp[2]) ? node280 : node267;
							assign node267 = (inp[8]) ? node275 : node268;
								assign node268 = (inp[7]) ? node272 : node269;
									assign node269 = (inp[0]) ? 11'b00001111111 : 11'b00000111111;
									assign node272 = (inp[4]) ? 11'b00000011111 : 11'b00000111111;
								assign node275 = (inp[10]) ? node277 : 11'b00000011111;
									assign node277 = (inp[4]) ? 11'b00000001111 : 11'b00000011111;
							assign node280 = (inp[4]) ? 11'b00000001111 : node281;
								assign node281 = (inp[0]) ? 11'b00000001111 : 11'b00000011111;
				assign node285 = (inp[4]) ? node341 : node286;
					assign node286 = (inp[0]) ? node308 : node287;
						assign node287 = (inp[10]) ? node299 : node288;
							assign node288 = (inp[6]) ? node292 : node289;
								assign node289 = (inp[7]) ? 11'b00000111111 : 11'b00011111111;
								assign node292 = (inp[2]) ? 11'b00000111111 : node293;
									assign node293 = (inp[7]) ? node295 : 11'b00001111111;
										assign node295 = (inp[9]) ? 11'b00000111111 : 11'b00001111111;
							assign node299 = (inp[8]) ? node303 : node300;
								assign node300 = (inp[2]) ? 11'b00000111111 : 11'b00001111111;
								assign node303 = (inp[2]) ? 11'b00000001111 : node304;
									assign node304 = (inp[7]) ? 11'b00000011111 : 11'b00000111111;
						assign node308 = (inp[6]) ? node326 : node309;
							assign node309 = (inp[10]) ? node321 : node310;
								assign node310 = (inp[2]) ? node316 : node311;
									assign node311 = (inp[9]) ? node313 : 11'b00011111111;
										assign node313 = (inp[8]) ? 11'b00000111111 : 11'b00001111111;
									assign node316 = (inp[8]) ? node318 : 11'b00000111111;
										assign node318 = (inp[9]) ? 11'b00000011111 : 11'b00000111111;
								assign node321 = (inp[7]) ? 11'b00000001111 : node322;
									assign node322 = (inp[9]) ? 11'b00000011111 : 11'b00000111111;
							assign node326 = (inp[8]) ? node332 : node327;
								assign node327 = (inp[9]) ? 11'b00000011111 : node328;
									assign node328 = (inp[7]) ? 11'b00000011111 : 11'b00000111111;
								assign node332 = (inp[7]) ? 11'b00000000011 : node333;
									assign node333 = (inp[2]) ? 11'b00000001111 : node334;
										assign node334 = (inp[9]) ? node336 : 11'b00000011111;
											assign node336 = (inp[10]) ? 11'b00000001111 : 11'b00000011111;
					assign node341 = (inp[2]) ? node363 : node342;
						assign node342 = (inp[10]) ? node352 : node343;
							assign node343 = (inp[7]) ? node347 : node344;
								assign node344 = (inp[6]) ? 11'b00000111111 : 11'b00011111111;
								assign node347 = (inp[9]) ? 11'b00000011111 : node348;
									assign node348 = (inp[8]) ? 11'b00000011111 : 11'b00000111111;
							assign node352 = (inp[8]) ? node358 : node353;
								assign node353 = (inp[9]) ? node355 : 11'b00000011111;
									assign node355 = (inp[0]) ? 11'b00000001111 : 11'b00000011111;
								assign node358 = (inp[7]) ? 11'b00000001111 : node359;
									assign node359 = (inp[9]) ? 11'b00000001111 : 11'b00000011111;
						assign node363 = (inp[10]) ? node377 : node364;
							assign node364 = (inp[7]) ? node368 : node365;
								assign node365 = (inp[8]) ? 11'b00000001111 : 11'b00000011111;
								assign node368 = (inp[9]) ? node370 : 11'b00000001111;
									assign node370 = (inp[6]) ? 11'b00000000111 : node371;
										assign node371 = (inp[0]) ? node373 : 11'b00000001111;
											assign node373 = (inp[8]) ? 11'b00000000111 : 11'b00000001111;
							assign node377 = (inp[7]) ? 11'b00000000011 : node378;
								assign node378 = (inp[9]) ? 11'b00000000111 : 11'b00000001111;
		assign node382 = (inp[0]) ? node582 : node383;
			assign node383 = (inp[9]) ? node483 : node384;
				assign node384 = (inp[4]) ? node436 : node385;
					assign node385 = (inp[1]) ? node413 : node386;
						assign node386 = (inp[7]) ? node402 : node387;
							assign node387 = (inp[10]) ? node393 : node388;
								assign node388 = (inp[6]) ? node390 : 11'b00111111111;
									assign node390 = (inp[2]) ? 11'b00000111111 : 11'b00011111111;
								assign node393 = (inp[3]) ? 11'b00001111111 : node394;
									assign node394 = (inp[8]) ? 11'b00001111111 : node395;
										assign node395 = (inp[2]) ? node397 : 11'b00011111111;
											assign node397 = (inp[6]) ? 11'b00001111111 : 11'b00011111111;
							assign node402 = (inp[10]) ? node408 : node403;
								assign node403 = (inp[2]) ? 11'b00001111111 : node404;
									assign node404 = (inp[8]) ? 11'b00001111111 : 11'b00011111111;
								assign node408 = (inp[2]) ? 11'b00000111111 : node409;
									assign node409 = (inp[8]) ? 11'b00000111111 : 11'b00001111111;
						assign node413 = (inp[2]) ? node429 : node414;
							assign node414 = (inp[10]) ? 11'b00000111111 : node415;
								assign node415 = (inp[7]) ? node421 : node416;
									assign node416 = (inp[6]) ? 11'b00001111111 : node417;
										assign node417 = (inp[8]) ? 11'b00011111111 : 11'b00111111111;
									assign node421 = (inp[8]) ? node423 : 11'b00001111111;
										assign node423 = (inp[3]) ? node425 : 11'b00000111111;
											assign node425 = (inp[6]) ? 11'b00000011111 : 11'b00000111111;
							assign node429 = (inp[3]) ? node431 : 11'b00000111111;
								assign node431 = (inp[8]) ? 11'b00000011111 : node432;
									assign node432 = (inp[6]) ? 11'b00000001111 : 11'b00000011111;
					assign node436 = (inp[1]) ? node468 : node437;
						assign node437 = (inp[6]) ? node455 : node438;
							assign node438 = (inp[7]) ? node450 : node439;
								assign node439 = (inp[10]) ? node443 : node440;
									assign node440 = (inp[3]) ? 11'b00001111111 : 11'b00111111111;
									assign node443 = (inp[3]) ? 11'b00000111111 : node444;
										assign node444 = (inp[8]) ? node446 : 11'b00001111111;
											assign node446 = (inp[2]) ? 11'b00000111111 : 11'b00001111111;
								assign node450 = (inp[8]) ? 11'b00000011111 : node451;
									assign node451 = (inp[10]) ? 11'b00000111111 : 11'b00001111111;
							assign node455 = (inp[8]) ? node463 : node456;
								assign node456 = (inp[7]) ? node458 : 11'b00000111111;
									assign node458 = (inp[10]) ? 11'b00000011111 : node459;
										assign node459 = (inp[3]) ? 11'b00000011111 : 11'b00000111111;
								assign node463 = (inp[2]) ? 11'b00000011111 : node464;
									assign node464 = (inp[10]) ? 11'b00000011111 : 11'b00000111111;
						assign node468 = (inp[6]) ? node480 : node469;
							assign node469 = (inp[7]) ? node477 : node470;
								assign node470 = (inp[3]) ? node472 : 11'b00000111111;
									assign node472 = (inp[2]) ? 11'b00000011111 : node473;
										assign node473 = (inp[8]) ? 11'b00000011111 : 11'b00000111111;
								assign node477 = (inp[10]) ? 11'b00000001111 : 11'b00000011111;
							assign node480 = (inp[2]) ? 11'b00000000111 : 11'b00000001111;
				assign node483 = (inp[10]) ? node535 : node484;
					assign node484 = (inp[4]) ? node512 : node485;
						assign node485 = (inp[1]) ? node505 : node486;
							assign node486 = (inp[2]) ? node502 : node487;
								assign node487 = (inp[7]) ? node495 : node488;
									assign node488 = (inp[3]) ? 11'b00001111111 : node489;
										assign node489 = (inp[6]) ? node491 : 11'b00011111111;
											assign node491 = (inp[8]) ? 11'b00001111111 : 11'b00011111111;
									assign node495 = (inp[8]) ? 11'b00000111111 : node496;
										assign node496 = (inp[3]) ? node498 : 11'b00001111111;
											assign node498 = (inp[6]) ? 11'b00000111111 : 11'b00001111111;
								assign node502 = (inp[8]) ? 11'b00000011111 : 11'b00001111111;
							assign node505 = (inp[3]) ? 11'b00000011111 : node506;
								assign node506 = (inp[6]) ? node508 : 11'b00000111111;
									assign node508 = (inp[7]) ? 11'b00000111111 : 11'b00000011111;
						assign node512 = (inp[2]) ? node524 : node513;
							assign node513 = (inp[8]) ? node517 : node514;
								assign node514 = (inp[7]) ? 11'b00000111111 : 11'b00001111111;
								assign node517 = (inp[6]) ? node521 : node518;
									assign node518 = (inp[3]) ? 11'b00000011111 : 11'b00000111111;
									assign node521 = (inp[3]) ? 11'b00000001111 : 11'b00000011111;
							assign node524 = (inp[6]) ? node530 : node525;
								assign node525 = (inp[1]) ? node527 : 11'b00000111111;
									assign node527 = (inp[7]) ? 11'b00000001111 : 11'b00000011111;
								assign node530 = (inp[7]) ? node532 : 11'b00000001111;
									assign node532 = (inp[3]) ? 11'b00000000111 : 11'b00000001111;
					assign node535 = (inp[6]) ? node559 : node536;
						assign node536 = (inp[2]) ? node542 : node537;
							assign node537 = (inp[1]) ? 11'b00000011111 : node538;
								assign node538 = (inp[4]) ? 11'b00000111111 : 11'b00011111111;
							assign node542 = (inp[3]) ? node552 : node543;
								assign node543 = (inp[8]) ? node545 : 11'b00000111111;
									assign node545 = (inp[1]) ? node547 : 11'b00000011111;
										assign node547 = (inp[4]) ? 11'b00000001111 : node548;
											assign node548 = (inp[7]) ? 11'b00000001111 : 11'b00000011111;
								assign node552 = (inp[4]) ? 11'b00000000111 : node553;
									assign node553 = (inp[8]) ? 11'b00000001111 : node554;
										assign node554 = (inp[1]) ? 11'b00000001111 : 11'b00000011111;
						assign node559 = (inp[8]) ? node567 : node560;
							assign node560 = (inp[3]) ? node562 : 11'b00000011111;
								assign node562 = (inp[2]) ? node564 : 11'b00000011111;
									assign node564 = (inp[1]) ? 11'b00000000011 : 11'b00000001111;
							assign node567 = (inp[4]) ? node573 : node568;
								assign node568 = (inp[7]) ? node570 : 11'b00000011111;
									assign node570 = (inp[2]) ? 11'b00000000111 : 11'b00000011111;
								assign node573 = (inp[7]) ? node575 : 11'b00000000111;
									assign node575 = (inp[2]) ? 11'b00000000011 : node576;
										assign node576 = (inp[3]) ? node578 : 11'b00000000111;
											assign node578 = (inp[1]) ? 11'b00000000011 : 11'b00000000111;
			assign node582 = (inp[2]) ? node676 : node583;
				assign node583 = (inp[10]) ? node629 : node584;
					assign node584 = (inp[7]) ? node604 : node585;
						assign node585 = (inp[1]) ? node597 : node586;
							assign node586 = (inp[6]) ? 11'b00000111111 : node587;
								assign node587 = (inp[4]) ? node593 : node588;
									assign node588 = (inp[8]) ? 11'b00011111111 : node589;
										assign node589 = (inp[3]) ? 11'b00011111111 : 11'b00111111111;
									assign node593 = (inp[8]) ? 11'b00000111111 : 11'b00001111111;
							assign node597 = (inp[4]) ? 11'b00000011111 : node598;
								assign node598 = (inp[3]) ? 11'b00000111111 : node599;
									assign node599 = (inp[8]) ? 11'b00000111111 : 11'b00001111111;
						assign node604 = (inp[6]) ? node614 : node605;
							assign node605 = (inp[9]) ? node609 : node606;
								assign node606 = (inp[8]) ? 11'b00001111111 : 11'b00000111111;
								assign node609 = (inp[1]) ? 11'b00000011111 : node610;
									assign node610 = (inp[3]) ? 11'b00000011111 : 11'b00000111111;
							assign node614 = (inp[4]) ? node626 : node615;
								assign node615 = (inp[1]) ? node619 : node616;
									assign node616 = (inp[3]) ? 11'b00000011111 : 11'b00000111111;
									assign node619 = (inp[8]) ? node621 : 11'b00000011111;
										assign node621 = (inp[3]) ? 11'b00000001111 : node622;
											assign node622 = (inp[9]) ? 11'b00000001111 : 11'b00000011111;
								assign node626 = (inp[3]) ? 11'b00000000111 : 11'b00000001111;
					assign node629 = (inp[1]) ? node647 : node630;
						assign node630 = (inp[7]) ? node638 : node631;
							assign node631 = (inp[6]) ? 11'b00000011111 : node632;
								assign node632 = (inp[9]) ? node634 : 11'b00000111111;
									assign node634 = (inp[3]) ? 11'b00000011111 : 11'b00000111111;
							assign node638 = (inp[3]) ? node640 : 11'b00000011111;
								assign node640 = (inp[9]) ? 11'b00000000111 : node641;
									assign node641 = (inp[6]) ? node643 : 11'b00000011111;
										assign node643 = (inp[8]) ? 11'b00000001111 : 11'b00000011111;
						assign node647 = (inp[8]) ? node661 : node648;
							assign node648 = (inp[7]) ? node652 : node649;
								assign node649 = (inp[3]) ? 11'b00000011111 : 11'b00000111111;
								assign node652 = (inp[3]) ? node656 : node653;
									assign node653 = (inp[9]) ? 11'b00000000111 : 11'b00000011111;
									assign node656 = (inp[4]) ? node658 : 11'b00000001111;
										assign node658 = (inp[6]) ? 11'b00000000111 : 11'b00000001111;
							assign node661 = (inp[4]) ? node669 : node662;
								assign node662 = (inp[7]) ? node666 : node663;
									assign node663 = (inp[3]) ? 11'b00000001111 : 11'b00000011111;
									assign node666 = (inp[6]) ? 11'b00000000111 : 11'b00000001111;
								assign node669 = (inp[3]) ? node671 : 11'b00000001111;
									assign node671 = (inp[7]) ? 11'b00000000011 : node672;
										assign node672 = (inp[6]) ? 11'b00000000011 : 11'b00000000111;
				assign node676 = (inp[3]) ? node720 : node677;
					assign node677 = (inp[6]) ? node703 : node678;
						assign node678 = (inp[8]) ? node692 : node679;
							assign node679 = (inp[4]) ? node687 : node680;
								assign node680 = (inp[10]) ? node682 : 11'b00001111111;
									assign node682 = (inp[1]) ? node684 : 11'b00000111111;
										assign node684 = (inp[9]) ? 11'b00000011111 : 11'b00000111111;
								assign node687 = (inp[1]) ? node689 : 11'b00000011111;
									assign node689 = (inp[10]) ? 11'b00000001111 : 11'b00000011111;
							assign node692 = (inp[10]) ? node696 : node693;
								assign node693 = (inp[4]) ? 11'b00000111111 : 11'b00000011111;
								assign node696 = (inp[1]) ? node698 : 11'b00000001111;
									assign node698 = (inp[9]) ? node700 : 11'b00000000111;
										assign node700 = (inp[4]) ? 11'b00000000011 : 11'b00000000111;
						assign node703 = (inp[9]) ? node707 : node704;
							assign node704 = (inp[10]) ? 11'b00000001111 : 11'b00000011111;
							assign node707 = (inp[8]) ? node713 : node708;
								assign node708 = (inp[4]) ? 11'b00000001111 : node709;
									assign node709 = (inp[7]) ? 11'b00000000111 : 11'b00000001111;
								assign node713 = (inp[10]) ? 11'b00000000011 : node714;
									assign node714 = (inp[1]) ? 11'b00000000111 : node715;
										assign node715 = (inp[7]) ? 11'b00000000111 : 11'b00000001111;
					assign node720 = (inp[10]) ? node744 : node721;
						assign node721 = (inp[1]) ? node735 : node722;
							assign node722 = (inp[8]) ? node730 : node723;
								assign node723 = (inp[6]) ? 11'b00000011111 : node724;
									assign node724 = (inp[7]) ? 11'b00000011111 : node725;
										assign node725 = (inp[9]) ? 11'b00000011111 : 11'b00000111111;
								assign node730 = (inp[6]) ? 11'b00000000111 : node731;
									assign node731 = (inp[4]) ? 11'b00000001111 : 11'b00000011111;
							assign node735 = (inp[4]) ? node741 : node736;
								assign node736 = (inp[8]) ? 11'b00000000111 : node737;
									assign node737 = (inp[9]) ? 11'b00000000111 : 11'b00000001111;
								assign node741 = (inp[6]) ? 11'b00000000011 : 11'b00000000111;
						assign node744 = (inp[4]) ? node754 : node745;
							assign node745 = (inp[6]) ? node751 : node746;
								assign node746 = (inp[8]) ? 11'b00000000111 : node747;
									assign node747 = (inp[7]) ? 11'b00000001111 : 11'b00000011111;
								assign node751 = (inp[1]) ? 11'b00000000011 : 11'b00000000111;
							assign node754 = (inp[8]) ? node762 : node755;
								assign node755 = (inp[6]) ? node757 : 11'b00000000111;
									assign node757 = (inp[9]) ? node759 : 11'b00000000111;
										assign node759 = (inp[1]) ? 11'b00000000001 : 11'b00000000011;
								assign node762 = (inp[1]) ? node768 : node763;
									assign node763 = (inp[7]) ? node765 : 11'b00000000011;
										assign node765 = (inp[9]) ? 11'b00000000001 : 11'b00000000011;
									assign node768 = (inp[7]) ? 11'b00000000001 : node769;
										assign node769 = (inp[6]) ? 11'b00000000001 : 11'b00000000011;

endmodule