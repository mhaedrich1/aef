module dtc_split5_bm7 (
	input  wire [12-1:0] inp,
	output wire [1-1:0] outp
);

	wire [1-1:0] node1;
	wire [1-1:0] node2;
	wire [1-1:0] node3;
	wire [1-1:0] node4;
	wire [1-1:0] node5;
	wire [1-1:0] node6;
	wire [1-1:0] node7;
	wire [1-1:0] node9;
	wire [1-1:0] node11;
	wire [1-1:0] node14;
	wire [1-1:0] node15;
	wire [1-1:0] node16;
	wire [1-1:0] node19;
	wire [1-1:0] node20;
	wire [1-1:0] node24;
	wire [1-1:0] node26;
	wire [1-1:0] node29;
	wire [1-1:0] node30;
	wire [1-1:0] node31;
	wire [1-1:0] node33;
	wire [1-1:0] node35;
	wire [1-1:0] node38;
	wire [1-1:0] node39;
	wire [1-1:0] node41;
	wire [1-1:0] node44;
	wire [1-1:0] node46;
	wire [1-1:0] node49;
	wire [1-1:0] node51;
	wire [1-1:0] node53;
	wire [1-1:0] node55;
	wire [1-1:0] node58;
	wire [1-1:0] node59;
	wire [1-1:0] node60;
	wire [1-1:0] node61;
	wire [1-1:0] node62;
	wire [1-1:0] node64;
	wire [1-1:0] node67;
	wire [1-1:0] node68;
	wire [1-1:0] node72;
	wire [1-1:0] node74;
	wire [1-1:0] node75;
	wire [1-1:0] node78;
	wire [1-1:0] node81;
	wire [1-1:0] node82;
	wire [1-1:0] node83;
	wire [1-1:0] node84;
	wire [1-1:0] node88;
	wire [1-1:0] node89;
	wire [1-1:0] node93;
	wire [1-1:0] node95;
	wire [1-1:0] node96;
	wire [1-1:0] node100;
	wire [1-1:0] node101;
	wire [1-1:0] node102;
	wire [1-1:0] node103;
	wire [1-1:0] node104;
	wire [1-1:0] node108;
	wire [1-1:0] node111;
	wire [1-1:0] node113;
	wire [1-1:0] node114;
	wire [1-1:0] node118;
	wire [1-1:0] node119;
	wire [1-1:0] node120;
	wire [1-1:0] node124;
	wire [1-1:0] node125;
	wire [1-1:0] node126;
	wire [1-1:0] node130;
	wire [1-1:0] node131;
	wire [1-1:0] node135;
	wire [1-1:0] node136;
	wire [1-1:0] node137;
	wire [1-1:0] node138;
	wire [1-1:0] node139;
	wire [1-1:0] node140;
	wire [1-1:0] node141;
	wire [1-1:0] node145;
	wire [1-1:0] node147;
	wire [1-1:0] node150;
	wire [1-1:0] node152;
	wire [1-1:0] node153;
	wire [1-1:0] node156;
	wire [1-1:0] node159;
	wire [1-1:0] node160;
	wire [1-1:0] node161;
	wire [1-1:0] node165;
	wire [1-1:0] node167;
	wire [1-1:0] node170;
	wire [1-1:0] node171;
	wire [1-1:0] node172;
	wire [1-1:0] node174;
	wire [1-1:0] node177;
	wire [1-1:0] node178;
	wire [1-1:0] node182;
	wire [1-1:0] node183;
	wire [1-1:0] node185;
	wire [1-1:0] node186;
	wire [1-1:0] node189;
	wire [1-1:0] node192;
	wire [1-1:0] node193;
	wire [1-1:0] node194;
	wire [1-1:0] node199;
	wire [1-1:0] node200;
	wire [1-1:0] node201;
	wire [1-1:0] node202;
	wire [1-1:0] node203;
	wire [1-1:0] node204;
	wire [1-1:0] node208;
	wire [1-1:0] node210;
	wire [1-1:0] node213;
	wire [1-1:0] node214;
	wire [1-1:0] node215;
	wire [1-1:0] node218;
	wire [1-1:0] node221;
	wire [1-1:0] node223;
	wire [1-1:0] node226;
	wire [1-1:0] node227;
	wire [1-1:0] node229;
	wire [1-1:0] node231;
	wire [1-1:0] node234;
	wire [1-1:0] node235;
	wire [1-1:0] node236;
	wire [1-1:0] node239;
	wire [1-1:0] node243;
	wire [1-1:0] node244;
	wire [1-1:0] node245;
	wire [1-1:0] node246;
	wire [1-1:0] node249;
	wire [1-1:0] node252;
	wire [1-1:0] node254;
	wire [1-1:0] node256;
	wire [1-1:0] node259;
	wire [1-1:0] node260;
	wire [1-1:0] node262;
	wire [1-1:0] node266;
	wire [1-1:0] node267;
	wire [1-1:0] node268;
	wire [1-1:0] node269;
	wire [1-1:0] node270;
	wire [1-1:0] node271;
	wire [1-1:0] node275;
	wire [1-1:0] node276;
	wire [1-1:0] node278;
	wire [1-1:0] node280;
	wire [1-1:0] node283;
	wire [1-1:0] node284;
	wire [1-1:0] node286;
	wire [1-1:0] node289;
	wire [1-1:0] node291;
	wire [1-1:0] node294;
	wire [1-1:0] node295;
	wire [1-1:0] node296;
	wire [1-1:0] node297;
	wire [1-1:0] node300;
	wire [1-1:0] node303;
	wire [1-1:0] node304;
	wire [1-1:0] node307;
	wire [1-1:0] node309;
	wire [1-1:0] node312;
	wire [1-1:0] node313;
	wire [1-1:0] node314;
	wire [1-1:0] node318;
	wire [1-1:0] node319;
	wire [1-1:0] node320;
	wire [1-1:0] node324;
	wire [1-1:0] node327;
	wire [1-1:0] node328;
	wire [1-1:0] node329;
	wire [1-1:0] node330;
	wire [1-1:0] node332;
	wire [1-1:0] node336;
	wire [1-1:0] node337;
	wire [1-1:0] node338;
	wire [1-1:0] node339;
	wire [1-1:0] node344;
	wire [1-1:0] node345;
	wire [1-1:0] node346;
	wire [1-1:0] node350;
	wire [1-1:0] node351;
	wire [1-1:0] node355;
	wire [1-1:0] node356;
	wire [1-1:0] node357;
	wire [1-1:0] node360;
	wire [1-1:0] node362;
	wire [1-1:0] node363;
	wire [1-1:0] node367;
	wire [1-1:0] node368;
	wire [1-1:0] node369;
	wire [1-1:0] node371;
	wire [1-1:0] node374;
	wire [1-1:0] node377;
	wire [1-1:0] node378;
	wire [1-1:0] node382;
	wire [1-1:0] node383;
	wire [1-1:0] node384;
	wire [1-1:0] node385;
	wire [1-1:0] node387;
	wire [1-1:0] node388;
	wire [1-1:0] node389;
	wire [1-1:0] node393;
	wire [1-1:0] node394;
	wire [1-1:0] node398;
	wire [1-1:0] node399;
	wire [1-1:0] node401;
	wire [1-1:0] node404;
	wire [1-1:0] node406;
	wire [1-1:0] node408;
	wire [1-1:0] node411;
	wire [1-1:0] node412;
	wire [1-1:0] node413;
	wire [1-1:0] node414;
	wire [1-1:0] node418;
	wire [1-1:0] node420;
	wire [1-1:0] node421;
	wire [1-1:0] node425;
	wire [1-1:0] node426;
	wire [1-1:0] node428;
	wire [1-1:0] node432;
	wire [1-1:0] node433;
	wire [1-1:0] node434;
	wire [1-1:0] node435;
	wire [1-1:0] node436;
	wire [1-1:0] node437;
	wire [1-1:0] node440;
	wire [1-1:0] node444;
	wire [1-1:0] node445;
	wire [1-1:0] node448;
	wire [1-1:0] node451;
	wire [1-1:0] node452;
	wire [1-1:0] node453;
	wire [1-1:0] node454;
	wire [1-1:0] node458;
	wire [1-1:0] node460;
	wire [1-1:0] node463;
	wire [1-1:0] node464;
	wire [1-1:0] node468;
	wire [1-1:0] node469;
	wire [1-1:0] node470;
	wire [1-1:0] node471;
	wire [1-1:0] node473;
	wire [1-1:0] node476;
	wire [1-1:0] node478;
	wire [1-1:0] node481;
	wire [1-1:0] node482;
	wire [1-1:0] node485;
	wire [1-1:0] node486;
	wire [1-1:0] node491;
	wire [1-1:0] node492;
	wire [1-1:0] node493;
	wire [1-1:0] node494;
	wire [1-1:0] node495;
	wire [1-1:0] node496;
	wire [1-1:0] node497;
	wire [1-1:0] node498;
	wire [1-1:0] node501;
	wire [1-1:0] node502;
	wire [1-1:0] node506;
	wire [1-1:0] node508;
	wire [1-1:0] node511;
	wire [1-1:0] node512;
	wire [1-1:0] node513;
	wire [1-1:0] node517;
	wire [1-1:0] node518;
	wire [1-1:0] node519;
	wire [1-1:0] node523;
	wire [1-1:0] node524;
	wire [1-1:0] node527;
	wire [1-1:0] node530;
	wire [1-1:0] node531;
	wire [1-1:0] node532;
	wire [1-1:0] node533;
	wire [1-1:0] node535;
	wire [1-1:0] node538;
	wire [1-1:0] node539;
	wire [1-1:0] node542;
	wire [1-1:0] node545;
	wire [1-1:0] node546;
	wire [1-1:0] node547;
	wire [1-1:0] node550;
	wire [1-1:0] node554;
	wire [1-1:0] node556;
	wire [1-1:0] node557;
	wire [1-1:0] node558;
	wire [1-1:0] node562;
	wire [1-1:0] node563;
	wire [1-1:0] node567;
	wire [1-1:0] node568;
	wire [1-1:0] node569;
	wire [1-1:0] node570;
	wire [1-1:0] node572;
	wire [1-1:0] node573;
	wire [1-1:0] node576;
	wire [1-1:0] node579;
	wire [1-1:0] node580;
	wire [1-1:0] node582;
	wire [1-1:0] node586;
	wire [1-1:0] node587;
	wire [1-1:0] node588;
	wire [1-1:0] node590;
	wire [1-1:0] node594;
	wire [1-1:0] node596;
	wire [1-1:0] node597;
	wire [1-1:0] node601;
	wire [1-1:0] node602;
	wire [1-1:0] node603;
	wire [1-1:0] node605;
	wire [1-1:0] node606;
	wire [1-1:0] node609;
	wire [1-1:0] node612;
	wire [1-1:0] node614;
	wire [1-1:0] node615;
	wire [1-1:0] node618;
	wire [1-1:0] node621;
	wire [1-1:0] node622;
	wire [1-1:0] node624;
	wire [1-1:0] node625;
	wire [1-1:0] node628;
	wire [1-1:0] node631;
	wire [1-1:0] node632;
	wire [1-1:0] node634;
	wire [1-1:0] node638;
	wire [1-1:0] node639;
	wire [1-1:0] node640;
	wire [1-1:0] node641;
	wire [1-1:0] node642;
	wire [1-1:0] node644;
	wire [1-1:0] node647;
	wire [1-1:0] node648;
	wire [1-1:0] node649;
	wire [1-1:0] node653;
	wire [1-1:0] node654;
	wire [1-1:0] node658;
	wire [1-1:0] node659;
	wire [1-1:0] node660;
	wire [1-1:0] node663;
	wire [1-1:0] node665;
	wire [1-1:0] node669;
	wire [1-1:0] node670;
	wire [1-1:0] node671;
	wire [1-1:0] node673;
	wire [1-1:0] node675;
	wire [1-1:0] node678;
	wire [1-1:0] node679;
	wire [1-1:0] node680;
	wire [1-1:0] node685;
	wire [1-1:0] node686;
	wire [1-1:0] node687;
	wire [1-1:0] node689;
	wire [1-1:0] node693;
	wire [1-1:0] node695;
	wire [1-1:0] node696;
	wire [1-1:0] node700;
	wire [1-1:0] node701;
	wire [1-1:0] node702;
	wire [1-1:0] node703;
	wire [1-1:0] node704;
	wire [1-1:0] node705;
	wire [1-1:0] node710;
	wire [1-1:0] node712;
	wire [1-1:0] node715;
	wire [1-1:0] node716;
	wire [1-1:0] node717;
	wire [1-1:0] node719;
	wire [1-1:0] node722;
	wire [1-1:0] node725;
	wire [1-1:0] node726;
	wire [1-1:0] node727;
	wire [1-1:0] node730;
	wire [1-1:0] node733;
	wire [1-1:0] node735;
	wire [1-1:0] node738;
	wire [1-1:0] node739;
	wire [1-1:0] node741;
	wire [1-1:0] node742;
	wire [1-1:0] node745;
	wire [1-1:0] node747;
	wire [1-1:0] node750;
	wire [1-1:0] node751;
	wire [1-1:0] node753;
	wire [1-1:0] node756;
	wire [1-1:0] node757;
	wire [1-1:0] node759;
	wire [1-1:0] node763;
	wire [1-1:0] node764;
	wire [1-1:0] node765;
	wire [1-1:0] node766;
	wire [1-1:0] node767;
	wire [1-1:0] node768;
	wire [1-1:0] node769;
	wire [1-1:0] node771;
	wire [1-1:0] node774;
	wire [1-1:0] node775;
	wire [1-1:0] node780;
	wire [1-1:0] node781;
	wire [1-1:0] node783;
	wire [1-1:0] node784;
	wire [1-1:0] node787;
	wire [1-1:0] node790;
	wire [1-1:0] node792;
	wire [1-1:0] node793;
	wire [1-1:0] node797;
	wire [1-1:0] node798;
	wire [1-1:0] node799;
	wire [1-1:0] node801;
	wire [1-1:0] node804;
	wire [1-1:0] node807;
	wire [1-1:0] node808;
	wire [1-1:0] node809;
	wire [1-1:0] node814;
	wire [1-1:0] node815;
	wire [1-1:0] node816;
	wire [1-1:0] node817;
	wire [1-1:0] node818;
	wire [1-1:0] node821;
	wire [1-1:0] node823;
	wire [1-1:0] node826;
	wire [1-1:0] node827;
	wire [1-1:0] node830;
	wire [1-1:0] node832;
	wire [1-1:0] node835;
	wire [1-1:0] node836;
	wire [1-1:0] node837;
	wire [1-1:0] node839;
	wire [1-1:0] node842;
	wire [1-1:0] node845;
	wire [1-1:0] node846;
	wire [1-1:0] node847;
	wire [1-1:0] node852;
	wire [1-1:0] node853;
	wire [1-1:0] node855;
	wire [1-1:0] node856;
	wire [1-1:0] node860;
	wire [1-1:0] node861;
	wire [1-1:0] node863;
	wire [1-1:0] node864;
	wire [1-1:0] node867;
	wire [1-1:0] node870;
	wire [1-1:0] node871;
	wire [1-1:0] node874;
	wire [1-1:0] node877;
	wire [1-1:0] node878;
	wire [1-1:0] node879;
	wire [1-1:0] node880;
	wire [1-1:0] node881;
	wire [1-1:0] node882;
	wire [1-1:0] node884;
	wire [1-1:0] node888;
	wire [1-1:0] node890;
	wire [1-1:0] node893;
	wire [1-1:0] node894;
	wire [1-1:0] node896;
	wire [1-1:0] node897;
	wire [1-1:0] node900;
	wire [1-1:0] node903;
	wire [1-1:0] node905;
	wire [1-1:0] node906;
	wire [1-1:0] node910;
	wire [1-1:0] node911;
	wire [1-1:0] node912;
	wire [1-1:0] node913;
	wire [1-1:0] node916;
	wire [1-1:0] node917;
	wire [1-1:0] node921;
	wire [1-1:0] node922;
	wire [1-1:0] node926;
	wire [1-1:0] node927;
	wire [1-1:0] node928;
	wire [1-1:0] node930;
	wire [1-1:0] node934;
	wire [1-1:0] node936;
	wire [1-1:0] node937;
	wire [1-1:0] node941;
	wire [1-1:0] node942;
	wire [1-1:0] node943;
	wire [1-1:0] node944;
	wire [1-1:0] node945;
	wire [1-1:0] node947;
	wire [1-1:0] node950;
	wire [1-1:0] node952;
	wire [1-1:0] node955;
	wire [1-1:0] node957;
	wire [1-1:0] node959;
	wire [1-1:0] node962;
	wire [1-1:0] node963;
	wire [1-1:0] node964;
	wire [1-1:0] node965;
	wire [1-1:0] node969;
	wire [1-1:0] node970;
	wire [1-1:0] node973;
	wire [1-1:0] node976;
	wire [1-1:0] node977;
	wire [1-1:0] node978;
	wire [1-1:0] node982;
	wire [1-1:0] node985;
	wire [1-1:0] node986;
	wire [1-1:0] node988;
	wire [1-1:0] node990;
	wire [1-1:0] node992;
	wire [1-1:0] node995;
	wire [1-1:0] node996;
	wire [1-1:0] node997;
	wire [1-1:0] node998;
	wire [1-1:0] node1001;
	wire [1-1:0] node1004;
	wire [1-1:0] node1005;
	wire [1-1:0] node1009;
	wire [1-1:0] node1011;
	wire [1-1:0] node1013;
	wire [1-1:0] node1016;
	wire [1-1:0] node1017;
	wire [1-1:0] node1018;
	wire [1-1:0] node1019;
	wire [1-1:0] node1020;
	wire [1-1:0] node1021;
	wire [1-1:0] node1022;
	wire [1-1:0] node1023;
	wire [1-1:0] node1025;
	wire [1-1:0] node1027;
	wire [1-1:0] node1031;
	wire [1-1:0] node1032;
	wire [1-1:0] node1033;
	wire [1-1:0] node1034;
	wire [1-1:0] node1037;
	wire [1-1:0] node1042;
	wire [1-1:0] node1043;
	wire [1-1:0] node1044;
	wire [1-1:0] node1045;
	wire [1-1:0] node1049;
	wire [1-1:0] node1051;
	wire [1-1:0] node1054;
	wire [1-1:0] node1055;
	wire [1-1:0] node1056;
	wire [1-1:0] node1057;
	wire [1-1:0] node1061;
	wire [1-1:0] node1064;
	wire [1-1:0] node1066;
	wire [1-1:0] node1067;
	wire [1-1:0] node1071;
	wire [1-1:0] node1072;
	wire [1-1:0] node1073;
	wire [1-1:0] node1075;
	wire [1-1:0] node1076;
	wire [1-1:0] node1077;
	wire [1-1:0] node1081;
	wire [1-1:0] node1082;
	wire [1-1:0] node1085;
	wire [1-1:0] node1088;
	wire [1-1:0] node1089;
	wire [1-1:0] node1090;
	wire [1-1:0] node1092;
	wire [1-1:0] node1096;
	wire [1-1:0] node1097;
	wire [1-1:0] node1098;
	wire [1-1:0] node1103;
	wire [1-1:0] node1104;
	wire [1-1:0] node1105;
	wire [1-1:0] node1107;
	wire [1-1:0] node1108;
	wire [1-1:0] node1111;
	wire [1-1:0] node1114;
	wire [1-1:0] node1115;
	wire [1-1:0] node1118;
	wire [1-1:0] node1121;
	wire [1-1:0] node1122;
	wire [1-1:0] node1123;
	wire [1-1:0] node1126;
	wire [1-1:0] node1127;
	wire [1-1:0] node1131;
	wire [1-1:0] node1132;
	wire [1-1:0] node1136;
	wire [1-1:0] node1137;
	wire [1-1:0] node1138;
	wire [1-1:0] node1139;
	wire [1-1:0] node1141;
	wire [1-1:0] node1142;
	wire [1-1:0] node1146;
	wire [1-1:0] node1147;
	wire [1-1:0] node1148;
	wire [1-1:0] node1152;
	wire [1-1:0] node1154;
	wire [1-1:0] node1157;
	wire [1-1:0] node1159;
	wire [1-1:0] node1160;
	wire [1-1:0] node1164;
	wire [1-1:0] node1165;
	wire [1-1:0] node1166;
	wire [1-1:0] node1167;
	wire [1-1:0] node1169;
	wire [1-1:0] node1172;
	wire [1-1:0] node1173;
	wire [1-1:0] node1174;
	wire [1-1:0] node1177;
	wire [1-1:0] node1181;
	wire [1-1:0] node1183;
	wire [1-1:0] node1184;
	wire [1-1:0] node1185;
	wire [1-1:0] node1190;
	wire [1-1:0] node1191;
	wire [1-1:0] node1192;
	wire [1-1:0] node1193;
	wire [1-1:0] node1194;
	wire [1-1:0] node1198;
	wire [1-1:0] node1201;
	wire [1-1:0] node1203;
	wire [1-1:0] node1206;
	wire [1-1:0] node1207;
	wire [1-1:0] node1208;
	wire [1-1:0] node1209;
	wire [1-1:0] node1213;
	wire [1-1:0] node1214;
	wire [1-1:0] node1217;
	wire [1-1:0] node1220;
	wire [1-1:0] node1222;
	wire [1-1:0] node1225;
	wire [1-1:0] node1226;
	wire [1-1:0] node1227;
	wire [1-1:0] node1228;
	wire [1-1:0] node1229;
	wire [1-1:0] node1230;
	wire [1-1:0] node1231;
	wire [1-1:0] node1232;
	wire [1-1:0] node1236;
	wire [1-1:0] node1237;
	wire [1-1:0] node1241;
	wire [1-1:0] node1242;
	wire [1-1:0] node1243;
	wire [1-1:0] node1248;
	wire [1-1:0] node1249;
	wire [1-1:0] node1250;
	wire [1-1:0] node1251;
	wire [1-1:0] node1256;
	wire [1-1:0] node1257;
	wire [1-1:0] node1261;
	wire [1-1:0] node1262;
	wire [1-1:0] node1263;
	wire [1-1:0] node1265;
	wire [1-1:0] node1267;
	wire [1-1:0] node1271;
	wire [1-1:0] node1273;
	wire [1-1:0] node1276;
	wire [1-1:0] node1277;
	wire [1-1:0] node1278;
	wire [1-1:0] node1279;
	wire [1-1:0] node1280;
	wire [1-1:0] node1281;
	wire [1-1:0] node1285;
	wire [1-1:0] node1286;
	wire [1-1:0] node1290;
	wire [1-1:0] node1292;
	wire [1-1:0] node1293;
	wire [1-1:0] node1297;
	wire [1-1:0] node1298;
	wire [1-1:0] node1299;
	wire [1-1:0] node1301;
	wire [1-1:0] node1305;
	wire [1-1:0] node1306;
	wire [1-1:0] node1307;
	wire [1-1:0] node1310;
	wire [1-1:0] node1314;
	wire [1-1:0] node1315;
	wire [1-1:0] node1316;
	wire [1-1:0] node1317;
	wire [1-1:0] node1318;
	wire [1-1:0] node1321;
	wire [1-1:0] node1325;
	wire [1-1:0] node1326;
	wire [1-1:0] node1328;
	wire [1-1:0] node1331;
	wire [1-1:0] node1332;
	wire [1-1:0] node1336;
	wire [1-1:0] node1338;
	wire [1-1:0] node1339;
	wire [1-1:0] node1343;
	wire [1-1:0] node1344;
	wire [1-1:0] node1345;
	wire [1-1:0] node1346;
	wire [1-1:0] node1347;
	wire [1-1:0] node1349;
	wire [1-1:0] node1352;
	wire [1-1:0] node1353;
	wire [1-1:0] node1354;
	wire [1-1:0] node1358;
	wire [1-1:0] node1359;
	wire [1-1:0] node1362;
	wire [1-1:0] node1365;
	wire [1-1:0] node1366;
	wire [1-1:0] node1367;
	wire [1-1:0] node1369;
	wire [1-1:0] node1372;
	wire [1-1:0] node1373;
	wire [1-1:0] node1377;
	wire [1-1:0] node1379;
	wire [1-1:0] node1381;
	wire [1-1:0] node1384;
	wire [1-1:0] node1385;
	wire [1-1:0] node1386;
	wire [1-1:0] node1388;
	wire [1-1:0] node1389;
	wire [1-1:0] node1394;
	wire [1-1:0] node1396;
	wire [1-1:0] node1397;
	wire [1-1:0] node1399;
	wire [1-1:0] node1402;
	wire [1-1:0] node1403;
	wire [1-1:0] node1407;
	wire [1-1:0] node1408;
	wire [1-1:0] node1409;
	wire [1-1:0] node1410;
	wire [1-1:0] node1411;
	wire [1-1:0] node1412;
	wire [1-1:0] node1416;
	wire [1-1:0] node1417;
	wire [1-1:0] node1420;
	wire [1-1:0] node1423;
	wire [1-1:0] node1425;
	wire [1-1:0] node1427;
	wire [1-1:0] node1430;
	wire [1-1:0] node1431;
	wire [1-1:0] node1432;
	wire [1-1:0] node1433;
	wire [1-1:0] node1437;
	wire [1-1:0] node1439;
	wire [1-1:0] node1442;
	wire [1-1:0] node1444;
	wire [1-1:0] node1446;
	wire [1-1:0] node1449;
	wire [1-1:0] node1450;
	wire [1-1:0] node1451;
	wire [1-1:0] node1452;
	wire [1-1:0] node1453;
	wire [1-1:0] node1457;
	wire [1-1:0] node1458;
	wire [1-1:0] node1462;
	wire [1-1:0] node1463;
	wire [1-1:0] node1466;
	wire [1-1:0] node1468;
	wire [1-1:0] node1471;
	wire [1-1:0] node1472;
	wire [1-1:0] node1473;
	wire [1-1:0] node1474;
	wire [1-1:0] node1479;
	wire [1-1:0] node1480;
	wire [1-1:0] node1483;
	wire [1-1:0] node1486;
	wire [1-1:0] node1487;
	wire [1-1:0] node1488;
	wire [1-1:0] node1489;
	wire [1-1:0] node1490;
	wire [1-1:0] node1491;
	wire [1-1:0] node1492;
	wire [1-1:0] node1494;
	wire [1-1:0] node1496;
	wire [1-1:0] node1499;
	wire [1-1:0] node1501;
	wire [1-1:0] node1502;
	wire [1-1:0] node1505;
	wire [1-1:0] node1508;
	wire [1-1:0] node1510;
	wire [1-1:0] node1511;
	wire [1-1:0] node1513;
	wire [1-1:0] node1516;
	wire [1-1:0] node1519;
	wire [1-1:0] node1520;
	wire [1-1:0] node1521;
	wire [1-1:0] node1522;
	wire [1-1:0] node1523;
	wire [1-1:0] node1527;
	wire [1-1:0] node1528;
	wire [1-1:0] node1532;
	wire [1-1:0] node1534;
	wire [1-1:0] node1537;
	wire [1-1:0] node1538;
	wire [1-1:0] node1539;
	wire [1-1:0] node1543;
	wire [1-1:0] node1544;
	wire [1-1:0] node1546;
	wire [1-1:0] node1550;
	wire [1-1:0] node1551;
	wire [1-1:0] node1552;
	wire [1-1:0] node1553;
	wire [1-1:0] node1555;
	wire [1-1:0] node1558;
	wire [1-1:0] node1559;
	wire [1-1:0] node1560;
	wire [1-1:0] node1563;
	wire [1-1:0] node1566;
	wire [1-1:0] node1567;
	wire [1-1:0] node1570;
	wire [1-1:0] node1573;
	wire [1-1:0] node1574;
	wire [1-1:0] node1577;
	wire [1-1:0] node1579;
	wire [1-1:0] node1581;
	wire [1-1:0] node1584;
	wire [1-1:0] node1585;
	wire [1-1:0] node1586;
	wire [1-1:0] node1587;
	wire [1-1:0] node1592;
	wire [1-1:0] node1593;
	wire [1-1:0] node1595;
	wire [1-1:0] node1598;
	wire [1-1:0] node1600;
	wire [1-1:0] node1601;
	wire [1-1:0] node1604;
	wire [1-1:0] node1607;
	wire [1-1:0] node1608;
	wire [1-1:0] node1609;
	wire [1-1:0] node1610;
	wire [1-1:0] node1611;
	wire [1-1:0] node1612;
	wire [1-1:0] node1614;
	wire [1-1:0] node1617;
	wire [1-1:0] node1619;
	wire [1-1:0] node1623;
	wire [1-1:0] node1624;
	wire [1-1:0] node1625;
	wire [1-1:0] node1627;
	wire [1-1:0] node1630;
	wire [1-1:0] node1632;
	wire [1-1:0] node1635;
	wire [1-1:0] node1636;
	wire [1-1:0] node1639;
	wire [1-1:0] node1640;
	wire [1-1:0] node1644;
	wire [1-1:0] node1645;
	wire [1-1:0] node1646;
	wire [1-1:0] node1647;
	wire [1-1:0] node1648;
	wire [1-1:0] node1651;
	wire [1-1:0] node1655;
	wire [1-1:0] node1656;
	wire [1-1:0] node1657;
	wire [1-1:0] node1661;
	wire [1-1:0] node1664;
	wire [1-1:0] node1666;
	wire [1-1:0] node1669;
	wire [1-1:0] node1670;
	wire [1-1:0] node1671;
	wire [1-1:0] node1672;
	wire [1-1:0] node1673;
	wire [1-1:0] node1677;
	wire [1-1:0] node1678;
	wire [1-1:0] node1681;
	wire [1-1:0] node1682;
	wire [1-1:0] node1686;
	wire [1-1:0] node1687;
	wire [1-1:0] node1689;
	wire [1-1:0] node1690;
	wire [1-1:0] node1694;
	wire [1-1:0] node1696;
	wire [1-1:0] node1697;
	wire [1-1:0] node1701;
	wire [1-1:0] node1702;
	wire [1-1:0] node1703;
	wire [1-1:0] node1704;
	wire [1-1:0] node1705;
	wire [1-1:0] node1708;
	wire [1-1:0] node1712;
	wire [1-1:0] node1713;
	wire [1-1:0] node1714;
	wire [1-1:0] node1717;
	wire [1-1:0] node1721;
	wire [1-1:0] node1722;
	wire [1-1:0] node1724;
	wire [1-1:0] node1726;
	wire [1-1:0] node1729;
	wire [1-1:0] node1730;
	wire [1-1:0] node1731;
	wire [1-1:0] node1736;
	wire [1-1:0] node1737;
	wire [1-1:0] node1738;
	wire [1-1:0] node1739;
	wire [1-1:0] node1740;
	wire [1-1:0] node1741;
	wire [1-1:0] node1743;
	wire [1-1:0] node1746;
	wire [1-1:0] node1748;
	wire [1-1:0] node1750;
	wire [1-1:0] node1753;
	wire [1-1:0] node1754;
	wire [1-1:0] node1755;
	wire [1-1:0] node1757;
	wire [1-1:0] node1761;
	wire [1-1:0] node1762;
	wire [1-1:0] node1764;
	wire [1-1:0] node1767;
	wire [1-1:0] node1769;
	wire [1-1:0] node1772;
	wire [1-1:0] node1773;
	wire [1-1:0] node1774;
	wire [1-1:0] node1775;
	wire [1-1:0] node1777;
	wire [1-1:0] node1780;
	wire [1-1:0] node1783;
	wire [1-1:0] node1784;
	wire [1-1:0] node1788;
	wire [1-1:0] node1789;
	wire [1-1:0] node1790;
	wire [1-1:0] node1791;
	wire [1-1:0] node1796;
	wire [1-1:0] node1797;
	wire [1-1:0] node1799;
	wire [1-1:0] node1803;
	wire [1-1:0] node1804;
	wire [1-1:0] node1805;
	wire [1-1:0] node1806;
	wire [1-1:0] node1807;
	wire [1-1:0] node1809;
	wire [1-1:0] node1813;
	wire [1-1:0] node1814;
	wire [1-1:0] node1815;
	wire [1-1:0] node1819;
	wire [1-1:0] node1820;
	wire [1-1:0] node1823;
	wire [1-1:0] node1826;
	wire [1-1:0] node1827;
	wire [1-1:0] node1828;
	wire [1-1:0] node1830;
	wire [1-1:0] node1833;
	wire [1-1:0] node1834;
	wire [1-1:0] node1838;
	wire [1-1:0] node1839;
	wire [1-1:0] node1841;
	wire [1-1:0] node1844;
	wire [1-1:0] node1846;
	wire [1-1:0] node1849;
	wire [1-1:0] node1850;
	wire [1-1:0] node1851;
	wire [1-1:0] node1852;
	wire [1-1:0] node1853;
	wire [1-1:0] node1856;
	wire [1-1:0] node1861;
	wire [1-1:0] node1862;
	wire [1-1:0] node1863;
	wire [1-1:0] node1865;
	wire [1-1:0] node1869;
	wire [1-1:0] node1870;
	wire [1-1:0] node1872;
	wire [1-1:0] node1876;
	wire [1-1:0] node1877;
	wire [1-1:0] node1878;
	wire [1-1:0] node1879;
	wire [1-1:0] node1880;
	wire [1-1:0] node1881;
	wire [1-1:0] node1882;
	wire [1-1:0] node1886;
	wire [1-1:0] node1890;
	wire [1-1:0] node1891;
	wire [1-1:0] node1892;
	wire [1-1:0] node1893;
	wire [1-1:0] node1896;
	wire [1-1:0] node1900;
	wire [1-1:0] node1903;
	wire [1-1:0] node1904;
	wire [1-1:0] node1905;
	wire [1-1:0] node1907;
	wire [1-1:0] node1909;
	wire [1-1:0] node1912;
	wire [1-1:0] node1913;
	wire [1-1:0] node1915;
	wire [1-1:0] node1919;
	wire [1-1:0] node1920;
	wire [1-1:0] node1921;
	wire [1-1:0] node1922;
	wire [1-1:0] node1927;
	wire [1-1:0] node1929;
	wire [1-1:0] node1931;
	wire [1-1:0] node1934;
	wire [1-1:0] node1935;
	wire [1-1:0] node1936;
	wire [1-1:0] node1937;
	wire [1-1:0] node1939;
	wire [1-1:0] node1942;
	wire [1-1:0] node1944;
	wire [1-1:0] node1945;
	wire [1-1:0] node1949;
	wire [1-1:0] node1951;
	wire [1-1:0] node1953;
	wire [1-1:0] node1955;
	wire [1-1:0] node1958;
	wire [1-1:0] node1959;
	wire [1-1:0] node1960;
	wire [1-1:0] node1961;
	wire [1-1:0] node1963;
	wire [1-1:0] node1967;
	wire [1-1:0] node1968;
	wire [1-1:0] node1971;
	wire [1-1:0] node1974;
	wire [1-1:0] node1975;
	wire [1-1:0] node1977;
	wire [1-1:0] node1980;
	wire [1-1:0] node1981;
	wire [1-1:0] node1982;
	wire [1-1:0] node1985;
	wire [1-1:0] node1988;
	wire [1-1:0] node1990;

	assign outp = (inp[9]) ? node1016 : node1;
		assign node1 = (inp[3]) ? node491 : node2;
			assign node2 = (inp[8]) ? node266 : node3;
				assign node3 = (inp[11]) ? node135 : node4;
					assign node4 = (inp[5]) ? node58 : node5;
						assign node5 = (inp[0]) ? node29 : node6;
							assign node6 = (inp[7]) ? node14 : node7;
								assign node7 = (inp[6]) ? node9 : 1'b0;
									assign node9 = (inp[10]) ? node11 : 1'b0;
										assign node11 = (inp[2]) ? 1'b1 : 1'b0;
								assign node14 = (inp[2]) ? node24 : node15;
									assign node15 = (inp[6]) ? node19 : node16;
										assign node16 = (inp[10]) ? 1'b0 : 1'b1;
										assign node19 = (inp[10]) ? 1'b1 : node20;
											assign node20 = (inp[1]) ? 1'b0 : 1'b0;
									assign node24 = (inp[10]) ? node26 : 1'b0;
										assign node26 = (inp[1]) ? 1'b1 : 1'b0;
							assign node29 = (inp[7]) ? node49 : node30;
								assign node30 = (inp[1]) ? node38 : node31;
									assign node31 = (inp[10]) ? node33 : 1'b1;
										assign node33 = (inp[6]) ? node35 : 1'b1;
											assign node35 = (inp[4]) ? 1'b0 : 1'b1;
									assign node38 = (inp[4]) ? node44 : node39;
										assign node39 = (inp[6]) ? node41 : 1'b1;
											assign node41 = (inp[10]) ? 1'b1 : 1'b0;
										assign node44 = (inp[6]) ? node46 : 1'b0;
											assign node46 = (inp[2]) ? 1'b0 : 1'b0;
								assign node49 = (inp[4]) ? node51 : 1'b0;
									assign node51 = (inp[10]) ? node53 : 1'b0;
										assign node53 = (inp[1]) ? node55 : 1'b1;
											assign node55 = (inp[6]) ? 1'b0 : 1'b0;
						assign node58 = (inp[1]) ? node100 : node59;
							assign node59 = (inp[6]) ? node81 : node60;
								assign node60 = (inp[2]) ? node72 : node61;
									assign node61 = (inp[0]) ? node67 : node62;
										assign node62 = (inp[7]) ? node64 : 1'b1;
											assign node64 = (inp[10]) ? 1'b0 : 1'b1;
										assign node67 = (inp[10]) ? 1'b0 : node68;
											assign node68 = (inp[7]) ? 1'b1 : 1'b0;
									assign node72 = (inp[7]) ? node74 : 1'b0;
										assign node74 = (inp[4]) ? node78 : node75;
											assign node75 = (inp[10]) ? 1'b0 : 1'b1;
											assign node78 = (inp[10]) ? 1'b1 : 1'b0;
								assign node81 = (inp[4]) ? node93 : node82;
									assign node82 = (inp[2]) ? node88 : node83;
										assign node83 = (inp[7]) ? 1'b0 : node84;
											assign node84 = (inp[10]) ? 1'b0 : 1'b1;
										assign node88 = (inp[10]) ? 1'b1 : node89;
											assign node89 = (inp[7]) ? 1'b0 : 1'b0;
									assign node93 = (inp[10]) ? node95 : 1'b1;
										assign node95 = (inp[7]) ? 1'b1 : node96;
											assign node96 = (inp[0]) ? 1'b0 : 1'b1;
							assign node100 = (inp[10]) ? node118 : node101;
								assign node101 = (inp[7]) ? node111 : node102;
									assign node102 = (inp[6]) ? node108 : node103;
										assign node103 = (inp[4]) ? 1'b1 : node104;
											assign node104 = (inp[0]) ? 1'b1 : 1'b0;
										assign node108 = (inp[0]) ? 1'b0 : 1'b1;
									assign node111 = (inp[0]) ? node113 : 1'b1;
										assign node113 = (inp[2]) ? 1'b1 : node114;
											assign node114 = (inp[4]) ? 1'b0 : 1'b1;
								assign node118 = (inp[7]) ? node124 : node119;
									assign node119 = (inp[0]) ? 1'b1 : node120;
										assign node120 = (inp[4]) ? 1'b1 : 1'b0;
									assign node124 = (inp[6]) ? node130 : node125;
										assign node125 = (inp[0]) ? 1'b0 : node126;
											assign node126 = (inp[4]) ? 1'b0 : 1'b1;
										assign node130 = (inp[4]) ? 1'b1 : node131;
											assign node131 = (inp[0]) ? 1'b0 : 1'b1;
					assign node135 = (inp[7]) ? node199 : node136;
						assign node136 = (inp[2]) ? node170 : node137;
							assign node137 = (inp[6]) ? node159 : node138;
								assign node138 = (inp[4]) ? node150 : node139;
									assign node139 = (inp[1]) ? node145 : node140;
										assign node140 = (inp[5]) ? 1'b1 : node141;
											assign node141 = (inp[10]) ? 1'b1 : 1'b0;
										assign node145 = (inp[0]) ? node147 : 1'b0;
											assign node147 = (inp[10]) ? 1'b1 : 1'b0;
									assign node150 = (inp[10]) ? node152 : 1'b1;
										assign node152 = (inp[0]) ? node156 : node153;
											assign node153 = (inp[5]) ? 1'b1 : 1'b0;
											assign node156 = (inp[1]) ? 1'b1 : 1'b0;
								assign node159 = (inp[4]) ? node165 : node160;
									assign node160 = (inp[1]) ? 1'b0 : node161;
										assign node161 = (inp[5]) ? 1'b0 : 1'b1;
									assign node165 = (inp[0]) ? node167 : 1'b1;
										assign node167 = (inp[5]) ? 1'b0 : 1'b1;
							assign node170 = (inp[10]) ? node182 : node171;
								assign node171 = (inp[4]) ? node177 : node172;
									assign node172 = (inp[0]) ? node174 : 1'b0;
										assign node174 = (inp[6]) ? 1'b1 : 1'b0;
									assign node177 = (inp[6]) ? 1'b0 : node178;
										assign node178 = (inp[0]) ? 1'b0 : 1'b1;
								assign node182 = (inp[6]) ? node192 : node183;
									assign node183 = (inp[0]) ? node185 : 1'b0;
										assign node185 = (inp[1]) ? node189 : node186;
											assign node186 = (inp[5]) ? 1'b0 : 1'b1;
											assign node189 = (inp[5]) ? 1'b1 : 1'b0;
									assign node192 = (inp[4]) ? 1'b1 : node193;
										assign node193 = (inp[1]) ? 1'b1 : node194;
											assign node194 = (inp[5]) ? 1'b0 : 1'b0;
						assign node199 = (inp[1]) ? node243 : node200;
							assign node200 = (inp[10]) ? node226 : node201;
								assign node201 = (inp[4]) ? node213 : node202;
									assign node202 = (inp[6]) ? node208 : node203;
										assign node203 = (inp[0]) ? 1'b0 : node204;
											assign node204 = (inp[5]) ? 1'b0 : 1'b0;
										assign node208 = (inp[2]) ? node210 : 1'b0;
											assign node210 = (inp[5]) ? 1'b0 : 1'b0;
									assign node213 = (inp[0]) ? node221 : node214;
										assign node214 = (inp[6]) ? node218 : node215;
											assign node215 = (inp[5]) ? 1'b1 : 1'b0;
											assign node218 = (inp[5]) ? 1'b0 : 1'b0;
										assign node221 = (inp[2]) ? node223 : 1'b0;
											assign node223 = (inp[5]) ? 1'b0 : 1'b0;
								assign node226 = (inp[0]) ? node234 : node227;
									assign node227 = (inp[2]) ? node229 : 1'b0;
										assign node229 = (inp[5]) ? node231 : 1'b1;
											assign node231 = (inp[4]) ? 1'b0 : 1'b1;
									assign node234 = (inp[4]) ? 1'b1 : node235;
										assign node235 = (inp[6]) ? node239 : node236;
											assign node236 = (inp[5]) ? 1'b1 : 1'b0;
											assign node239 = (inp[2]) ? 1'b0 : 1'b1;
							assign node243 = (inp[5]) ? node259 : node244;
								assign node244 = (inp[2]) ? node252 : node245;
									assign node245 = (inp[4]) ? node249 : node246;
										assign node246 = (inp[6]) ? 1'b1 : 1'b0;
										assign node249 = (inp[6]) ? 1'b0 : 1'b1;
									assign node252 = (inp[4]) ? node254 : 1'b0;
										assign node254 = (inp[0]) ? node256 : 1'b0;
											assign node256 = (inp[6]) ? 1'b1 : 1'b0;
								assign node259 = (inp[6]) ? 1'b0 : node260;
									assign node260 = (inp[10]) ? node262 : 1'b0;
										assign node262 = (inp[2]) ? 1'b1 : 1'b0;
				assign node266 = (inp[5]) ? node382 : node267;
					assign node267 = (inp[7]) ? node327 : node268;
						assign node268 = (inp[2]) ? node294 : node269;
							assign node269 = (inp[0]) ? node275 : node270;
								assign node270 = (inp[11]) ? 1'b0 : node271;
									assign node271 = (inp[4]) ? 1'b0 : 1'b1;
								assign node275 = (inp[1]) ? node283 : node276;
									assign node276 = (inp[10]) ? node278 : 1'b0;
										assign node278 = (inp[6]) ? node280 : 1'b0;
											assign node280 = (inp[4]) ? 1'b1 : 1'b0;
									assign node283 = (inp[4]) ? node289 : node284;
										assign node284 = (inp[11]) ? node286 : 1'b0;
											assign node286 = (inp[10]) ? 1'b1 : 1'b0;
										assign node289 = (inp[11]) ? node291 : 1'b1;
											assign node291 = (inp[10]) ? 1'b0 : 1'b1;
							assign node294 = (inp[1]) ? node312 : node295;
								assign node295 = (inp[6]) ? node303 : node296;
									assign node296 = (inp[0]) ? node300 : node297;
										assign node297 = (inp[11]) ? 1'b0 : 1'b1;
										assign node300 = (inp[11]) ? 1'b1 : 1'b0;
									assign node303 = (inp[0]) ? node307 : node304;
										assign node304 = (inp[11]) ? 1'b1 : 1'b0;
										assign node307 = (inp[10]) ? node309 : 1'b1;
											assign node309 = (inp[11]) ? 1'b0 : 1'b1;
								assign node312 = (inp[10]) ? node318 : node313;
									assign node313 = (inp[11]) ? 1'b0 : node314;
										assign node314 = (inp[4]) ? 1'b1 : 1'b0;
									assign node318 = (inp[11]) ? node324 : node319;
										assign node319 = (inp[0]) ? 1'b0 : node320;
											assign node320 = (inp[4]) ? 1'b0 : 1'b1;
										assign node324 = (inp[6]) ? 1'b1 : 1'b0;
						assign node327 = (inp[2]) ? node355 : node328;
							assign node328 = (inp[4]) ? node336 : node329;
								assign node329 = (inp[0]) ? 1'b0 : node330;
									assign node330 = (inp[6]) ? node332 : 1'b1;
										assign node332 = (inp[1]) ? 1'b0 : 1'b1;
								assign node336 = (inp[10]) ? node344 : node337;
									assign node337 = (inp[6]) ? 1'b1 : node338;
										assign node338 = (inp[1]) ? 1'b1 : node339;
											assign node339 = (inp[0]) ? 1'b0 : 1'b1;
									assign node344 = (inp[11]) ? node350 : node345;
										assign node345 = (inp[6]) ? 1'b0 : node346;
											assign node346 = (inp[1]) ? 1'b0 : 1'b0;
										assign node350 = (inp[6]) ? 1'b1 : node351;
											assign node351 = (inp[1]) ? 1'b0 : 1'b0;
							assign node355 = (inp[1]) ? node367 : node356;
								assign node356 = (inp[11]) ? node360 : node357;
									assign node357 = (inp[10]) ? 1'b1 : 1'b0;
									assign node360 = (inp[6]) ? node362 : 1'b0;
										assign node362 = (inp[0]) ? 1'b0 : node363;
											assign node363 = (inp[4]) ? 1'b0 : 1'b1;
								assign node367 = (inp[6]) ? node377 : node368;
									assign node368 = (inp[0]) ? node374 : node369;
										assign node369 = (inp[10]) ? node371 : 1'b0;
											assign node371 = (inp[11]) ? 1'b0 : 1'b1;
										assign node374 = (inp[4]) ? 1'b0 : 1'b1;
									assign node377 = (inp[11]) ? 1'b1 : node378;
										assign node378 = (inp[10]) ? 1'b0 : 1'b1;
					assign node382 = (inp[10]) ? node432 : node383;
						assign node383 = (inp[6]) ? node411 : node384;
							assign node384 = (inp[2]) ? node398 : node385;
								assign node385 = (inp[7]) ? node387 : 1'b1;
									assign node387 = (inp[11]) ? node393 : node388;
										assign node388 = (inp[4]) ? 1'b1 : node389;
											assign node389 = (inp[0]) ? 1'b0 : 1'b1;
										assign node393 = (inp[1]) ? 1'b0 : node394;
											assign node394 = (inp[0]) ? 1'b1 : 1'b0;
								assign node398 = (inp[7]) ? node404 : node399;
									assign node399 = (inp[1]) ? node401 : 1'b0;
										assign node401 = (inp[11]) ? 1'b0 : 1'b1;
									assign node404 = (inp[4]) ? node406 : 1'b1;
										assign node406 = (inp[0]) ? node408 : 1'b1;
											assign node408 = (inp[1]) ? 1'b0 : 1'b0;
							assign node411 = (inp[7]) ? node425 : node412;
								assign node412 = (inp[11]) ? node418 : node413;
									assign node413 = (inp[4]) ? 1'b1 : node414;
										assign node414 = (inp[0]) ? 1'b0 : 1'b1;
									assign node418 = (inp[0]) ? node420 : 1'b0;
										assign node420 = (inp[4]) ? 1'b0 : node421;
											assign node421 = (inp[2]) ? 1'b0 : 1'b1;
								assign node425 = (inp[4]) ? 1'b0 : node426;
									assign node426 = (inp[1]) ? node428 : 1'b1;
										assign node428 = (inp[0]) ? 1'b1 : 1'b0;
						assign node432 = (inp[7]) ? node468 : node433;
							assign node433 = (inp[6]) ? node451 : node434;
								assign node434 = (inp[4]) ? node444 : node435;
									assign node435 = (inp[1]) ? 1'b0 : node436;
										assign node436 = (inp[2]) ? node440 : node437;
											assign node437 = (inp[11]) ? 1'b0 : 1'b1;
											assign node440 = (inp[11]) ? 1'b1 : 1'b0;
									assign node444 = (inp[1]) ? node448 : node445;
										assign node445 = (inp[0]) ? 1'b0 : 1'b1;
										assign node448 = (inp[11]) ? 1'b0 : 1'b1;
								assign node451 = (inp[1]) ? node463 : node452;
									assign node452 = (inp[4]) ? node458 : node453;
										assign node453 = (inp[11]) ? 1'b0 : node454;
											assign node454 = (inp[0]) ? 1'b0 : 1'b1;
										assign node458 = (inp[2]) ? node460 : 1'b1;
											assign node460 = (inp[11]) ? 1'b0 : 1'b1;
									assign node463 = (inp[0]) ? 1'b1 : node464;
										assign node464 = (inp[2]) ? 1'b1 : 1'b0;
							assign node468 = (inp[1]) ? 1'b0 : node469;
								assign node469 = (inp[11]) ? node481 : node470;
									assign node470 = (inp[0]) ? node476 : node471;
										assign node471 = (inp[6]) ? node473 : 1'b0;
											assign node473 = (inp[2]) ? 1'b0 : 1'b1;
										assign node476 = (inp[4]) ? node478 : 1'b0;
											assign node478 = (inp[6]) ? 1'b0 : 1'b1;
									assign node481 = (inp[4]) ? node485 : node482;
										assign node482 = (inp[6]) ? 1'b1 : 1'b0;
										assign node485 = (inp[6]) ? 1'b0 : node486;
											assign node486 = (inp[0]) ? 1'b0 : 1'b1;
			assign node491 = (inp[2]) ? node763 : node492;
				assign node492 = (inp[6]) ? node638 : node493;
					assign node493 = (inp[0]) ? node567 : node494;
						assign node494 = (inp[4]) ? node530 : node495;
							assign node495 = (inp[1]) ? node511 : node496;
								assign node496 = (inp[8]) ? node506 : node497;
									assign node497 = (inp[7]) ? node501 : node498;
										assign node498 = (inp[5]) ? 1'b0 : 1'b1;
										assign node501 = (inp[10]) ? 1'b0 : node502;
											assign node502 = (inp[11]) ? 1'b1 : 1'b0;
									assign node506 = (inp[7]) ? node508 : 1'b0;
										assign node508 = (inp[11]) ? 1'b0 : 1'b1;
								assign node511 = (inp[10]) ? node517 : node512;
									assign node512 = (inp[8]) ? 1'b1 : node513;
										assign node513 = (inp[5]) ? 1'b0 : 1'b1;
									assign node517 = (inp[11]) ? node523 : node518;
										assign node518 = (inp[7]) ? 1'b0 : node519;
											assign node519 = (inp[5]) ? 1'b1 : 1'b0;
										assign node523 = (inp[7]) ? node527 : node524;
											assign node524 = (inp[8]) ? 1'b0 : 1'b1;
											assign node527 = (inp[5]) ? 1'b1 : 1'b0;
							assign node530 = (inp[5]) ? node554 : node531;
								assign node531 = (inp[8]) ? node545 : node532;
									assign node532 = (inp[1]) ? node538 : node533;
										assign node533 = (inp[11]) ? node535 : 1'b1;
											assign node535 = (inp[7]) ? 1'b1 : 1'b0;
										assign node538 = (inp[11]) ? node542 : node539;
											assign node539 = (inp[7]) ? 1'b1 : 1'b0;
											assign node542 = (inp[10]) ? 1'b1 : 1'b0;
									assign node545 = (inp[11]) ? 1'b0 : node546;
										assign node546 = (inp[10]) ? node550 : node547;
											assign node547 = (inp[7]) ? 1'b0 : 1'b0;
											assign node550 = (inp[1]) ? 1'b1 : 1'b0;
								assign node554 = (inp[7]) ? node556 : 1'b1;
									assign node556 = (inp[10]) ? node562 : node557;
										assign node557 = (inp[8]) ? 1'b0 : node558;
											assign node558 = (inp[1]) ? 1'b0 : 1'b0;
										assign node562 = (inp[8]) ? 1'b1 : node563;
											assign node563 = (inp[1]) ? 1'b1 : 1'b0;
						assign node567 = (inp[8]) ? node601 : node568;
							assign node568 = (inp[10]) ? node586 : node569;
								assign node569 = (inp[1]) ? node579 : node570;
									assign node570 = (inp[11]) ? node572 : 1'b0;
										assign node572 = (inp[4]) ? node576 : node573;
											assign node573 = (inp[5]) ? 1'b0 : 1'b1;
											assign node576 = (inp[5]) ? 1'b1 : 1'b0;
									assign node579 = (inp[11]) ? 1'b0 : node580;
										assign node580 = (inp[4]) ? node582 : 1'b0;
											assign node582 = (inp[5]) ? 1'b0 : 1'b1;
								assign node586 = (inp[11]) ? node594 : node587;
									assign node587 = (inp[4]) ? 1'b1 : node588;
										assign node588 = (inp[7]) ? node590 : 1'b0;
											assign node590 = (inp[1]) ? 1'b1 : 1'b0;
									assign node594 = (inp[7]) ? node596 : 1'b0;
										assign node596 = (inp[4]) ? 1'b0 : node597;
											assign node597 = (inp[1]) ? 1'b0 : 1'b0;
							assign node601 = (inp[10]) ? node621 : node602;
								assign node602 = (inp[5]) ? node612 : node603;
									assign node603 = (inp[11]) ? node605 : 1'b1;
										assign node605 = (inp[4]) ? node609 : node606;
											assign node606 = (inp[1]) ? 1'b0 : 1'b1;
											assign node609 = (inp[7]) ? 1'b0 : 1'b1;
									assign node612 = (inp[7]) ? node614 : 1'b0;
										assign node614 = (inp[11]) ? node618 : node615;
											assign node615 = (inp[1]) ? 1'b1 : 1'b0;
											assign node618 = (inp[1]) ? 1'b0 : 1'b0;
								assign node621 = (inp[1]) ? node631 : node622;
									assign node622 = (inp[11]) ? node624 : 1'b0;
										assign node624 = (inp[7]) ? node628 : node625;
											assign node625 = (inp[5]) ? 1'b1 : 1'b0;
											assign node628 = (inp[5]) ? 1'b0 : 1'b1;
									assign node631 = (inp[11]) ? 1'b1 : node632;
										assign node632 = (inp[4]) ? node634 : 1'b1;
											assign node634 = (inp[7]) ? 1'b0 : 1'b0;
					assign node638 = (inp[8]) ? node700 : node639;
						assign node639 = (inp[7]) ? node669 : node640;
							assign node640 = (inp[1]) ? node658 : node641;
								assign node641 = (inp[11]) ? node647 : node642;
									assign node642 = (inp[10]) ? node644 : 1'b0;
										assign node644 = (inp[4]) ? 1'b1 : 1'b0;
									assign node647 = (inp[4]) ? node653 : node648;
										assign node648 = (inp[0]) ? 1'b1 : node649;
											assign node649 = (inp[5]) ? 1'b0 : 1'b0;
										assign node653 = (inp[5]) ? 1'b1 : node654;
											assign node654 = (inp[10]) ? 1'b1 : 1'b0;
								assign node658 = (inp[5]) ? 1'b0 : node659;
									assign node659 = (inp[4]) ? node663 : node660;
										assign node660 = (inp[10]) ? 1'b0 : 1'b1;
										assign node663 = (inp[10]) ? node665 : 1'b0;
											assign node665 = (inp[11]) ? 1'b1 : 1'b0;
							assign node669 = (inp[11]) ? node685 : node670;
								assign node670 = (inp[4]) ? node678 : node671;
									assign node671 = (inp[10]) ? node673 : 1'b1;
										assign node673 = (inp[5]) ? node675 : 1'b0;
											assign node675 = (inp[0]) ? 1'b1 : 1'b0;
									assign node678 = (inp[5]) ? 1'b1 : node679;
										assign node679 = (inp[1]) ? 1'b1 : node680;
											assign node680 = (inp[0]) ? 1'b0 : 1'b1;
								assign node685 = (inp[4]) ? node693 : node686;
									assign node686 = (inp[1]) ? 1'b1 : node687;
										assign node687 = (inp[0]) ? node689 : 1'b1;
											assign node689 = (inp[5]) ? 1'b0 : 1'b1;
									assign node693 = (inp[0]) ? node695 : 1'b0;
										assign node695 = (inp[1]) ? 1'b0 : node696;
											assign node696 = (inp[5]) ? 1'b0 : 1'b1;
						assign node700 = (inp[1]) ? node738 : node701;
							assign node701 = (inp[10]) ? node715 : node702;
								assign node702 = (inp[11]) ? node710 : node703;
									assign node703 = (inp[0]) ? 1'b0 : node704;
										assign node704 = (inp[5]) ? 1'b0 : node705;
											assign node705 = (inp[4]) ? 1'b1 : 1'b0;
									assign node710 = (inp[0]) ? node712 : 1'b0;
										assign node712 = (inp[5]) ? 1'b1 : 1'b0;
								assign node715 = (inp[0]) ? node725 : node716;
									assign node716 = (inp[5]) ? node722 : node717;
										assign node717 = (inp[4]) ? node719 : 1'b0;
											assign node719 = (inp[11]) ? 1'b1 : 1'b0;
										assign node722 = (inp[11]) ? 1'b0 : 1'b1;
									assign node725 = (inp[5]) ? node733 : node726;
										assign node726 = (inp[4]) ? node730 : node727;
											assign node727 = (inp[7]) ? 1'b0 : 1'b1;
											assign node730 = (inp[7]) ? 1'b0 : 1'b0;
										assign node733 = (inp[11]) ? node735 : 1'b0;
											assign node735 = (inp[7]) ? 1'b0 : 1'b1;
							assign node738 = (inp[7]) ? node750 : node739;
								assign node739 = (inp[11]) ? node741 : 1'b1;
									assign node741 = (inp[10]) ? node745 : node742;
										assign node742 = (inp[4]) ? 1'b0 : 1'b1;
										assign node745 = (inp[4]) ? node747 : 1'b0;
											assign node747 = (inp[0]) ? 1'b1 : 1'b0;
								assign node750 = (inp[4]) ? node756 : node751;
									assign node751 = (inp[0]) ? node753 : 1'b0;
										assign node753 = (inp[5]) ? 1'b1 : 1'b0;
									assign node756 = (inp[0]) ? 1'b0 : node757;
										assign node757 = (inp[10]) ? node759 : 1'b1;
											assign node759 = (inp[11]) ? 1'b1 : 1'b0;
				assign node763 = (inp[0]) ? node877 : node764;
					assign node764 = (inp[7]) ? node814 : node765;
						assign node765 = (inp[5]) ? node797 : node766;
							assign node766 = (inp[8]) ? node780 : node767;
								assign node767 = (inp[10]) ? 1'b1 : node768;
									assign node768 = (inp[1]) ? node774 : node769;
										assign node769 = (inp[11]) ? node771 : 1'b1;
											assign node771 = (inp[6]) ? 1'b1 : 1'b0;
										assign node774 = (inp[6]) ? 1'b0 : node775;
											assign node775 = (inp[4]) ? 1'b0 : 1'b0;
								assign node780 = (inp[11]) ? node790 : node781;
									assign node781 = (inp[4]) ? node783 : 1'b0;
										assign node783 = (inp[10]) ? node787 : node784;
											assign node784 = (inp[6]) ? 1'b1 : 1'b0;
											assign node787 = (inp[6]) ? 1'b0 : 1'b0;
									assign node790 = (inp[4]) ? node792 : 1'b1;
										assign node792 = (inp[1]) ? 1'b0 : node793;
											assign node793 = (inp[10]) ? 1'b0 : 1'b1;
							assign node797 = (inp[11]) ? node807 : node798;
								assign node798 = (inp[6]) ? node804 : node799;
									assign node799 = (inp[4]) ? node801 : 1'b0;
										assign node801 = (inp[1]) ? 1'b0 : 1'b1;
									assign node804 = (inp[10]) ? 1'b0 : 1'b1;
								assign node807 = (inp[8]) ? 1'b0 : node808;
									assign node808 = (inp[10]) ? 1'b0 : node809;
										assign node809 = (inp[1]) ? 1'b0 : 1'b1;
						assign node814 = (inp[4]) ? node852 : node815;
							assign node815 = (inp[8]) ? node835 : node816;
								assign node816 = (inp[5]) ? node826 : node817;
									assign node817 = (inp[1]) ? node821 : node818;
										assign node818 = (inp[10]) ? 1'b1 : 1'b0;
										assign node821 = (inp[10]) ? node823 : 1'b1;
											assign node823 = (inp[6]) ? 1'b1 : 1'b0;
									assign node826 = (inp[1]) ? node830 : node827;
										assign node827 = (inp[11]) ? 1'b0 : 1'b1;
										assign node830 = (inp[11]) ? node832 : 1'b0;
											assign node832 = (inp[10]) ? 1'b0 : 1'b1;
								assign node835 = (inp[1]) ? node845 : node836;
									assign node836 = (inp[5]) ? node842 : node837;
										assign node837 = (inp[10]) ? node839 : 1'b0;
											assign node839 = (inp[6]) ? 1'b0 : 1'b0;
										assign node842 = (inp[10]) ? 1'b0 : 1'b1;
									assign node845 = (inp[5]) ? 1'b1 : node846;
										assign node846 = (inp[6]) ? 1'b0 : node847;
											assign node847 = (inp[11]) ? 1'b1 : 1'b0;
							assign node852 = (inp[6]) ? node860 : node853;
								assign node853 = (inp[11]) ? node855 : 1'b1;
									assign node855 = (inp[1]) ? 1'b1 : node856;
										assign node856 = (inp[5]) ? 1'b1 : 1'b0;
								assign node860 = (inp[1]) ? node870 : node861;
									assign node861 = (inp[10]) ? node863 : 1'b1;
										assign node863 = (inp[8]) ? node867 : node864;
											assign node864 = (inp[11]) ? 1'b1 : 1'b0;
											assign node867 = (inp[11]) ? 1'b0 : 1'b1;
									assign node870 = (inp[5]) ? node874 : node871;
										assign node871 = (inp[8]) ? 1'b0 : 1'b1;
										assign node874 = (inp[8]) ? 1'b1 : 1'b0;
					assign node877 = (inp[7]) ? node941 : node878;
						assign node878 = (inp[4]) ? node910 : node879;
							assign node879 = (inp[8]) ? node893 : node880;
								assign node880 = (inp[1]) ? node888 : node881;
									assign node881 = (inp[5]) ? 1'b1 : node882;
										assign node882 = (inp[11]) ? node884 : 1'b1;
											assign node884 = (inp[6]) ? 1'b1 : 1'b0;
									assign node888 = (inp[5]) ? node890 : 1'b1;
										assign node890 = (inp[6]) ? 1'b0 : 1'b1;
								assign node893 = (inp[10]) ? node903 : node894;
									assign node894 = (inp[1]) ? node896 : 1'b1;
										assign node896 = (inp[11]) ? node900 : node897;
											assign node897 = (inp[5]) ? 1'b1 : 1'b0;
											assign node900 = (inp[5]) ? 1'b0 : 1'b1;
									assign node903 = (inp[6]) ? node905 : 1'b0;
										assign node905 = (inp[1]) ? 1'b1 : node906;
											assign node906 = (inp[11]) ? 1'b1 : 1'b0;
							assign node910 = (inp[6]) ? node926 : node911;
								assign node911 = (inp[5]) ? node921 : node912;
									assign node912 = (inp[10]) ? node916 : node913;
										assign node913 = (inp[11]) ? 1'b0 : 1'b1;
										assign node916 = (inp[11]) ? 1'b1 : node917;
											assign node917 = (inp[1]) ? 1'b1 : 1'b0;
									assign node921 = (inp[10]) ? 1'b0 : node922;
										assign node922 = (inp[1]) ? 1'b0 : 1'b1;
								assign node926 = (inp[11]) ? node934 : node927;
									assign node927 = (inp[1]) ? 1'b1 : node928;
										assign node928 = (inp[10]) ? node930 : 1'b0;
											assign node930 = (inp[5]) ? 1'b0 : 1'b1;
									assign node934 = (inp[10]) ? node936 : 1'b1;
										assign node936 = (inp[8]) ? 1'b1 : node937;
											assign node937 = (inp[5]) ? 1'b1 : 1'b0;
						assign node941 = (inp[8]) ? node985 : node942;
							assign node942 = (inp[10]) ? node962 : node943;
								assign node943 = (inp[4]) ? node955 : node944;
									assign node944 = (inp[1]) ? node950 : node945;
										assign node945 = (inp[11]) ? node947 : 1'b1;
											assign node947 = (inp[6]) ? 1'b1 : 1'b0;
										assign node950 = (inp[5]) ? node952 : 1'b0;
											assign node952 = (inp[11]) ? 1'b1 : 1'b0;
									assign node955 = (inp[5]) ? node957 : 1'b0;
										assign node957 = (inp[1]) ? node959 : 1'b0;
											assign node959 = (inp[6]) ? 1'b0 : 1'b0;
								assign node962 = (inp[11]) ? node976 : node963;
									assign node963 = (inp[5]) ? node969 : node964;
										assign node964 = (inp[1]) ? 1'b1 : node965;
											assign node965 = (inp[6]) ? 1'b1 : 1'b0;
										assign node969 = (inp[4]) ? node973 : node970;
											assign node970 = (inp[6]) ? 1'b1 : 1'b0;
											assign node973 = (inp[1]) ? 1'b0 : 1'b1;
									assign node976 = (inp[5]) ? node982 : node977;
										assign node977 = (inp[6]) ? 1'b0 : node978;
											assign node978 = (inp[1]) ? 1'b1 : 1'b0;
										assign node982 = (inp[6]) ? 1'b1 : 1'b0;
							assign node985 = (inp[1]) ? node995 : node986;
								assign node986 = (inp[10]) ? node988 : 1'b1;
									assign node988 = (inp[11]) ? node990 : 1'b0;
										assign node990 = (inp[5]) ? node992 : 1'b1;
											assign node992 = (inp[6]) ? 1'b1 : 1'b0;
								assign node995 = (inp[11]) ? node1009 : node996;
									assign node996 = (inp[5]) ? node1004 : node997;
										assign node997 = (inp[6]) ? node1001 : node998;
											assign node998 = (inp[10]) ? 1'b1 : 1'b0;
											assign node1001 = (inp[10]) ? 1'b0 : 1'b1;
										assign node1004 = (inp[6]) ? 1'b0 : node1005;
											assign node1005 = (inp[4]) ? 1'b0 : 1'b1;
									assign node1009 = (inp[6]) ? node1011 : 1'b0;
										assign node1011 = (inp[5]) ? node1013 : 1'b1;
											assign node1013 = (inp[4]) ? 1'b1 : 1'b0;
		assign node1016 = (inp[0]) ? node1486 : node1017;
			assign node1017 = (inp[3]) ? node1225 : node1018;
				assign node1018 = (inp[11]) ? node1136 : node1019;
					assign node1019 = (inp[10]) ? node1071 : node1020;
						assign node1020 = (inp[5]) ? node1042 : node1021;
							assign node1021 = (inp[6]) ? node1031 : node1022;
								assign node1022 = (inp[2]) ? 1'b0 : node1023;
									assign node1023 = (inp[7]) ? node1025 : 1'b0;
										assign node1025 = (inp[8]) ? node1027 : 1'b1;
											assign node1027 = (inp[4]) ? 1'b0 : 1'b1;
								assign node1031 = (inp[8]) ? 1'b1 : node1032;
									assign node1032 = (inp[4]) ? 1'b1 : node1033;
										assign node1033 = (inp[7]) ? node1037 : node1034;
											assign node1034 = (inp[2]) ? 1'b1 : 1'b0;
											assign node1037 = (inp[1]) ? 1'b0 : 1'b0;
							assign node1042 = (inp[4]) ? node1054 : node1043;
								assign node1043 = (inp[7]) ? node1049 : node1044;
									assign node1044 = (inp[6]) ? 1'b0 : node1045;
										assign node1045 = (inp[2]) ? 1'b1 : 1'b0;
									assign node1049 = (inp[8]) ? node1051 : 1'b1;
										assign node1051 = (inp[2]) ? 1'b0 : 1'b1;
								assign node1054 = (inp[7]) ? node1064 : node1055;
									assign node1055 = (inp[6]) ? node1061 : node1056;
										assign node1056 = (inp[1]) ? 1'b0 : node1057;
											assign node1057 = (inp[8]) ? 1'b0 : 1'b1;
										assign node1061 = (inp[2]) ? 1'b0 : 1'b1;
									assign node1064 = (inp[1]) ? node1066 : 1'b0;
										assign node1066 = (inp[6]) ? 1'b0 : node1067;
											assign node1067 = (inp[8]) ? 1'b0 : 1'b1;
						assign node1071 = (inp[1]) ? node1103 : node1072;
							assign node1072 = (inp[2]) ? node1088 : node1073;
								assign node1073 = (inp[5]) ? node1075 : 1'b1;
									assign node1075 = (inp[6]) ? node1081 : node1076;
										assign node1076 = (inp[8]) ? 1'b0 : node1077;
											assign node1077 = (inp[7]) ? 1'b0 : 1'b1;
										assign node1081 = (inp[4]) ? node1085 : node1082;
											assign node1082 = (inp[7]) ? 1'b0 : 1'b1;
											assign node1085 = (inp[7]) ? 1'b1 : 1'b0;
								assign node1088 = (inp[7]) ? node1096 : node1089;
									assign node1089 = (inp[8]) ? 1'b1 : node1090;
										assign node1090 = (inp[6]) ? node1092 : 1'b0;
											assign node1092 = (inp[5]) ? 1'b1 : 1'b0;
									assign node1096 = (inp[6]) ? 1'b0 : node1097;
										assign node1097 = (inp[4]) ? 1'b0 : node1098;
											assign node1098 = (inp[5]) ? 1'b1 : 1'b0;
							assign node1103 = (inp[2]) ? node1121 : node1104;
								assign node1104 = (inp[5]) ? node1114 : node1105;
									assign node1105 = (inp[7]) ? node1107 : 1'b1;
										assign node1107 = (inp[4]) ? node1111 : node1108;
											assign node1108 = (inp[6]) ? 1'b0 : 1'b1;
											assign node1111 = (inp[6]) ? 1'b1 : 1'b0;
									assign node1114 = (inp[7]) ? node1118 : node1115;
										assign node1115 = (inp[4]) ? 1'b0 : 1'b1;
										assign node1118 = (inp[4]) ? 1'b1 : 1'b0;
								assign node1121 = (inp[6]) ? node1131 : node1122;
									assign node1122 = (inp[5]) ? node1126 : node1123;
										assign node1123 = (inp[7]) ? 1'b0 : 1'b1;
										assign node1126 = (inp[4]) ? 1'b1 : node1127;
											assign node1127 = (inp[8]) ? 1'b1 : 1'b0;
									assign node1131 = (inp[7]) ? 1'b1 : node1132;
										assign node1132 = (inp[5]) ? 1'b1 : 1'b0;
					assign node1136 = (inp[7]) ? node1164 : node1137;
						assign node1137 = (inp[2]) ? node1157 : node1138;
							assign node1138 = (inp[5]) ? node1146 : node1139;
								assign node1139 = (inp[6]) ? node1141 : 1'b1;
									assign node1141 = (inp[1]) ? 1'b1 : node1142;
										assign node1142 = (inp[4]) ? 1'b1 : 1'b0;
								assign node1146 = (inp[4]) ? node1152 : node1147;
									assign node1147 = (inp[6]) ? 1'b1 : node1148;
										assign node1148 = (inp[10]) ? 1'b0 : 1'b1;
									assign node1152 = (inp[8]) ? node1154 : 1'b0;
										assign node1154 = (inp[1]) ? 1'b1 : 1'b0;
							assign node1157 = (inp[5]) ? node1159 : 1'b1;
								assign node1159 = (inp[6]) ? 1'b1 : node1160;
									assign node1160 = (inp[8]) ? 1'b0 : 1'b1;
						assign node1164 = (inp[10]) ? node1190 : node1165;
							assign node1165 = (inp[2]) ? node1181 : node1166;
								assign node1166 = (inp[5]) ? node1172 : node1167;
									assign node1167 = (inp[6]) ? node1169 : 1'b0;
										assign node1169 = (inp[8]) ? 1'b1 : 1'b0;
									assign node1172 = (inp[4]) ? 1'b1 : node1173;
										assign node1173 = (inp[8]) ? node1177 : node1174;
											assign node1174 = (inp[1]) ? 1'b1 : 1'b0;
											assign node1177 = (inp[1]) ? 1'b0 : 1'b1;
								assign node1181 = (inp[5]) ? node1183 : 1'b1;
									assign node1183 = (inp[4]) ? 1'b1 : node1184;
										assign node1184 = (inp[8]) ? 1'b1 : node1185;
											assign node1185 = (inp[6]) ? 1'b1 : 1'b0;
							assign node1190 = (inp[8]) ? node1206 : node1191;
								assign node1191 = (inp[4]) ? node1201 : node1192;
									assign node1192 = (inp[5]) ? node1198 : node1193;
										assign node1193 = (inp[6]) ? 1'b0 : node1194;
											assign node1194 = (inp[2]) ? 1'b0 : 1'b1;
										assign node1198 = (inp[2]) ? 1'b1 : 1'b0;
									assign node1201 = (inp[1]) ? node1203 : 1'b0;
										assign node1203 = (inp[2]) ? 1'b0 : 1'b1;
								assign node1206 = (inp[1]) ? node1220 : node1207;
									assign node1207 = (inp[5]) ? node1213 : node1208;
										assign node1208 = (inp[4]) ? 1'b0 : node1209;
											assign node1209 = (inp[2]) ? 1'b1 : 1'b0;
										assign node1213 = (inp[2]) ? node1217 : node1214;
											assign node1214 = (inp[4]) ? 1'b1 : 1'b0;
											assign node1217 = (inp[6]) ? 1'b0 : 1'b0;
									assign node1220 = (inp[5]) ? node1222 : 1'b1;
										assign node1222 = (inp[4]) ? 1'b1 : 1'b0;
				assign node1225 = (inp[2]) ? node1343 : node1226;
					assign node1226 = (inp[7]) ? node1276 : node1227;
						assign node1227 = (inp[10]) ? node1261 : node1228;
							assign node1228 = (inp[5]) ? node1248 : node1229;
								assign node1229 = (inp[1]) ? node1241 : node1230;
									assign node1230 = (inp[4]) ? node1236 : node1231;
										assign node1231 = (inp[11]) ? 1'b0 : node1232;
											assign node1232 = (inp[6]) ? 1'b0 : 1'b1;
										assign node1236 = (inp[6]) ? 1'b1 : node1237;
											assign node1237 = (inp[11]) ? 1'b0 : 1'b1;
									assign node1241 = (inp[6]) ? 1'b0 : node1242;
										assign node1242 = (inp[4]) ? 1'b0 : node1243;
											assign node1243 = (inp[11]) ? 1'b0 : 1'b1;
								assign node1248 = (inp[11]) ? node1256 : node1249;
									assign node1249 = (inp[1]) ? 1'b0 : node1250;
										assign node1250 = (inp[4]) ? 1'b1 : node1251;
											assign node1251 = (inp[6]) ? 1'b0 : 1'b1;
									assign node1256 = (inp[8]) ? 1'b1 : node1257;
										assign node1257 = (inp[4]) ? 1'b0 : 1'b1;
							assign node1261 = (inp[4]) ? node1271 : node1262;
								assign node1262 = (inp[6]) ? 1'b1 : node1263;
									assign node1263 = (inp[5]) ? node1265 : 1'b0;
										assign node1265 = (inp[8]) ? node1267 : 1'b0;
											assign node1267 = (inp[1]) ? 1'b0 : 1'b1;
								assign node1271 = (inp[1]) ? node1273 : 1'b0;
									assign node1273 = (inp[5]) ? 1'b0 : 1'b1;
						assign node1276 = (inp[10]) ? node1314 : node1277;
							assign node1277 = (inp[1]) ? node1297 : node1278;
								assign node1278 = (inp[4]) ? node1290 : node1279;
									assign node1279 = (inp[8]) ? node1285 : node1280;
										assign node1280 = (inp[5]) ? 1'b0 : node1281;
											assign node1281 = (inp[6]) ? 1'b1 : 1'b0;
										assign node1285 = (inp[6]) ? 1'b0 : node1286;
											assign node1286 = (inp[11]) ? 1'b0 : 1'b0;
									assign node1290 = (inp[6]) ? node1292 : 1'b0;
										assign node1292 = (inp[8]) ? 1'b0 : node1293;
											assign node1293 = (inp[5]) ? 1'b1 : 1'b0;
								assign node1297 = (inp[11]) ? node1305 : node1298;
									assign node1298 = (inp[4]) ? 1'b0 : node1299;
										assign node1299 = (inp[5]) ? node1301 : 1'b1;
											assign node1301 = (inp[6]) ? 1'b0 : 1'b0;
									assign node1305 = (inp[5]) ? 1'b1 : node1306;
										assign node1306 = (inp[4]) ? node1310 : node1307;
											assign node1307 = (inp[8]) ? 1'b0 : 1'b0;
											assign node1310 = (inp[8]) ? 1'b1 : 1'b0;
							assign node1314 = (inp[5]) ? node1336 : node1315;
								assign node1315 = (inp[11]) ? node1325 : node1316;
									assign node1316 = (inp[6]) ? 1'b1 : node1317;
										assign node1317 = (inp[1]) ? node1321 : node1318;
											assign node1318 = (inp[4]) ? 1'b1 : 1'b0;
											assign node1321 = (inp[4]) ? 1'b0 : 1'b1;
									assign node1325 = (inp[6]) ? node1331 : node1326;
										assign node1326 = (inp[4]) ? node1328 : 1'b1;
											assign node1328 = (inp[8]) ? 1'b0 : 1'b1;
										assign node1331 = (inp[1]) ? 1'b0 : node1332;
											assign node1332 = (inp[4]) ? 1'b0 : 1'b1;
								assign node1336 = (inp[6]) ? node1338 : 1'b1;
									assign node1338 = (inp[8]) ? 1'b1 : node1339;
										assign node1339 = (inp[4]) ? 1'b0 : 1'b1;
					assign node1343 = (inp[4]) ? node1407 : node1344;
						assign node1344 = (inp[11]) ? node1384 : node1345;
							assign node1345 = (inp[10]) ? node1365 : node1346;
								assign node1346 = (inp[7]) ? node1352 : node1347;
									assign node1347 = (inp[6]) ? node1349 : 1'b1;
										assign node1349 = (inp[5]) ? 1'b0 : 1'b1;
									assign node1352 = (inp[8]) ? node1358 : node1353;
										assign node1353 = (inp[5]) ? 1'b0 : node1354;
											assign node1354 = (inp[1]) ? 1'b1 : 1'b0;
										assign node1358 = (inp[5]) ? node1362 : node1359;
											assign node1359 = (inp[1]) ? 1'b0 : 1'b1;
											assign node1362 = (inp[1]) ? 1'b1 : 1'b0;
								assign node1365 = (inp[1]) ? node1377 : node1366;
									assign node1366 = (inp[7]) ? node1372 : node1367;
										assign node1367 = (inp[6]) ? node1369 : 1'b0;
											assign node1369 = (inp[8]) ? 1'b0 : 1'b1;
										assign node1372 = (inp[5]) ? 1'b1 : node1373;
											assign node1373 = (inp[6]) ? 1'b1 : 1'b0;
									assign node1377 = (inp[6]) ? node1379 : 1'b0;
										assign node1379 = (inp[5]) ? node1381 : 1'b0;
											assign node1381 = (inp[7]) ? 1'b0 : 1'b1;
							assign node1384 = (inp[6]) ? node1394 : node1385;
								assign node1385 = (inp[5]) ? 1'b1 : node1386;
									assign node1386 = (inp[7]) ? node1388 : 1'b0;
										assign node1388 = (inp[10]) ? 1'b1 : node1389;
											assign node1389 = (inp[1]) ? 1'b0 : 1'b1;
								assign node1394 = (inp[7]) ? node1396 : 1'b1;
									assign node1396 = (inp[10]) ? node1402 : node1397;
										assign node1397 = (inp[5]) ? node1399 : 1'b1;
											assign node1399 = (inp[1]) ? 1'b0 : 1'b0;
										assign node1402 = (inp[5]) ? 1'b1 : node1403;
											assign node1403 = (inp[8]) ? 1'b1 : 1'b0;
						assign node1407 = (inp[1]) ? node1449 : node1408;
							assign node1408 = (inp[6]) ? node1430 : node1409;
								assign node1409 = (inp[10]) ? node1423 : node1410;
									assign node1410 = (inp[8]) ? node1416 : node1411;
										assign node1411 = (inp[11]) ? 1'b0 : node1412;
											assign node1412 = (inp[7]) ? 1'b0 : 1'b0;
										assign node1416 = (inp[7]) ? node1420 : node1417;
											assign node1417 = (inp[5]) ? 1'b1 : 1'b0;
											assign node1420 = (inp[5]) ? 1'b0 : 1'b1;
									assign node1423 = (inp[7]) ? node1425 : 1'b0;
										assign node1425 = (inp[8]) ? node1427 : 1'b0;
											assign node1427 = (inp[11]) ? 1'b1 : 1'b0;
								assign node1430 = (inp[11]) ? node1442 : node1431;
									assign node1431 = (inp[8]) ? node1437 : node1432;
										assign node1432 = (inp[10]) ? 1'b1 : node1433;
											assign node1433 = (inp[7]) ? 1'b1 : 1'b0;
										assign node1437 = (inp[7]) ? node1439 : 1'b1;
											assign node1439 = (inp[5]) ? 1'b1 : 1'b0;
									assign node1442 = (inp[5]) ? node1444 : 1'b0;
										assign node1444 = (inp[7]) ? node1446 : 1'b1;
											assign node1446 = (inp[10]) ? 1'b0 : 1'b0;
							assign node1449 = (inp[8]) ? node1471 : node1450;
								assign node1450 = (inp[6]) ? node1462 : node1451;
									assign node1451 = (inp[10]) ? node1457 : node1452;
										assign node1452 = (inp[11]) ? 1'b0 : node1453;
											assign node1453 = (inp[5]) ? 1'b1 : 1'b0;
										assign node1457 = (inp[7]) ? 1'b1 : node1458;
											assign node1458 = (inp[11]) ? 1'b1 : 1'b0;
									assign node1462 = (inp[11]) ? node1466 : node1463;
										assign node1463 = (inp[10]) ? 1'b0 : 1'b1;
										assign node1466 = (inp[5]) ? node1468 : 1'b1;
											assign node1468 = (inp[10]) ? 1'b1 : 1'b0;
								assign node1471 = (inp[5]) ? node1479 : node1472;
									assign node1472 = (inp[7]) ? 1'b0 : node1473;
										assign node1473 = (inp[10]) ? 1'b1 : node1474;
											assign node1474 = (inp[11]) ? 1'b1 : 1'b0;
									assign node1479 = (inp[10]) ? node1483 : node1480;
										assign node1480 = (inp[6]) ? 1'b1 : 1'b0;
										assign node1483 = (inp[6]) ? 1'b0 : 1'b1;
			assign node1486 = (inp[6]) ? node1736 : node1487;
				assign node1487 = (inp[5]) ? node1607 : node1488;
					assign node1488 = (inp[10]) ? node1550 : node1489;
						assign node1489 = (inp[4]) ? node1519 : node1490;
							assign node1490 = (inp[3]) ? node1508 : node1491;
								assign node1491 = (inp[11]) ? node1499 : node1492;
									assign node1492 = (inp[7]) ? node1494 : 1'b1;
										assign node1494 = (inp[1]) ? node1496 : 1'b0;
											assign node1496 = (inp[2]) ? 1'b1 : 1'b0;
									assign node1499 = (inp[7]) ? node1501 : 1'b0;
										assign node1501 = (inp[1]) ? node1505 : node1502;
											assign node1502 = (inp[2]) ? 1'b1 : 1'b0;
											assign node1505 = (inp[2]) ? 1'b0 : 1'b1;
								assign node1508 = (inp[11]) ? node1510 : 1'b0;
									assign node1510 = (inp[2]) ? node1516 : node1511;
										assign node1511 = (inp[7]) ? node1513 : 1'b1;
											assign node1513 = (inp[1]) ? 1'b1 : 1'b0;
										assign node1516 = (inp[7]) ? 1'b1 : 1'b0;
							assign node1519 = (inp[11]) ? node1537 : node1520;
								assign node1520 = (inp[3]) ? node1532 : node1521;
									assign node1521 = (inp[2]) ? node1527 : node1522;
										assign node1522 = (inp[8]) ? 1'b1 : node1523;
											assign node1523 = (inp[7]) ? 1'b1 : 1'b0;
										assign node1527 = (inp[7]) ? 1'b0 : node1528;
											assign node1528 = (inp[8]) ? 1'b0 : 1'b1;
									assign node1532 = (inp[7]) ? node1534 : 1'b1;
										assign node1534 = (inp[2]) ? 1'b1 : 1'b0;
								assign node1537 = (inp[7]) ? node1543 : node1538;
									assign node1538 = (inp[3]) ? 1'b0 : node1539;
										assign node1539 = (inp[1]) ? 1'b1 : 1'b0;
									assign node1543 = (inp[8]) ? 1'b1 : node1544;
										assign node1544 = (inp[2]) ? node1546 : 1'b1;
											assign node1546 = (inp[3]) ? 1'b0 : 1'b1;
						assign node1550 = (inp[2]) ? node1584 : node1551;
							assign node1551 = (inp[3]) ? node1573 : node1552;
								assign node1552 = (inp[7]) ? node1558 : node1553;
									assign node1553 = (inp[4]) ? node1555 : 1'b0;
										assign node1555 = (inp[1]) ? 1'b1 : 1'b0;
									assign node1558 = (inp[8]) ? node1566 : node1559;
										assign node1559 = (inp[11]) ? node1563 : node1560;
											assign node1560 = (inp[1]) ? 1'b1 : 1'b0;
											assign node1563 = (inp[1]) ? 1'b0 : 1'b1;
										assign node1566 = (inp[4]) ? node1570 : node1567;
											assign node1567 = (inp[1]) ? 1'b0 : 1'b1;
											assign node1570 = (inp[11]) ? 1'b0 : 1'b0;
								assign node1573 = (inp[4]) ? node1577 : node1574;
									assign node1574 = (inp[7]) ? 1'b0 : 1'b1;
									assign node1577 = (inp[7]) ? node1579 : 1'b0;
										assign node1579 = (inp[8]) ? node1581 : 1'b0;
											assign node1581 = (inp[11]) ? 1'b1 : 1'b0;
							assign node1584 = (inp[8]) ? node1592 : node1585;
								assign node1585 = (inp[11]) ? 1'b0 : node1586;
									assign node1586 = (inp[3]) ? 1'b0 : node1587;
										assign node1587 = (inp[1]) ? 1'b1 : 1'b0;
								assign node1592 = (inp[7]) ? node1598 : node1593;
									assign node1593 = (inp[4]) ? node1595 : 1'b0;
										assign node1595 = (inp[3]) ? 1'b0 : 1'b1;
									assign node1598 = (inp[3]) ? node1600 : 1'b0;
										assign node1600 = (inp[11]) ? node1604 : node1601;
											assign node1601 = (inp[1]) ? 1'b0 : 1'b1;
											assign node1604 = (inp[1]) ? 1'b1 : 1'b0;
					assign node1607 = (inp[4]) ? node1669 : node1608;
						assign node1608 = (inp[10]) ? node1644 : node1609;
							assign node1609 = (inp[7]) ? node1623 : node1610;
								assign node1610 = (inp[3]) ? 1'b1 : node1611;
									assign node1611 = (inp[2]) ? node1617 : node1612;
										assign node1612 = (inp[8]) ? node1614 : 1'b0;
											assign node1614 = (inp[11]) ? 1'b1 : 1'b0;
										assign node1617 = (inp[1]) ? node1619 : 1'b1;
											assign node1619 = (inp[8]) ? 1'b1 : 1'b0;
								assign node1623 = (inp[2]) ? node1635 : node1624;
									assign node1624 = (inp[8]) ? node1630 : node1625;
										assign node1625 = (inp[1]) ? node1627 : 1'b1;
											assign node1627 = (inp[11]) ? 1'b0 : 1'b0;
										assign node1630 = (inp[1]) ? node1632 : 1'b0;
											assign node1632 = (inp[3]) ? 1'b0 : 1'b0;
									assign node1635 = (inp[8]) ? node1639 : node1636;
										assign node1636 = (inp[11]) ? 1'b0 : 1'b1;
										assign node1639 = (inp[1]) ? 1'b0 : node1640;
											assign node1640 = (inp[11]) ? 1'b1 : 1'b0;
							assign node1644 = (inp[7]) ? node1664 : node1645;
								assign node1645 = (inp[11]) ? node1655 : node1646;
									assign node1646 = (inp[1]) ? 1'b1 : node1647;
										assign node1647 = (inp[8]) ? node1651 : node1648;
											assign node1648 = (inp[3]) ? 1'b1 : 1'b0;
											assign node1651 = (inp[3]) ? 1'b0 : 1'b1;
									assign node1655 = (inp[1]) ? node1661 : node1656;
										assign node1656 = (inp[2]) ? 1'b1 : node1657;
											assign node1657 = (inp[3]) ? 1'b1 : 1'b0;
										assign node1661 = (inp[2]) ? 1'b0 : 1'b1;
								assign node1664 = (inp[3]) ? node1666 : 1'b1;
									assign node1666 = (inp[1]) ? 1'b0 : 1'b1;
						assign node1669 = (inp[2]) ? node1701 : node1670;
							assign node1670 = (inp[1]) ? node1686 : node1671;
								assign node1671 = (inp[7]) ? node1677 : node1672;
									assign node1672 = (inp[8]) ? 1'b1 : node1673;
										assign node1673 = (inp[10]) ? 1'b0 : 1'b1;
									assign node1677 = (inp[3]) ? node1681 : node1678;
										assign node1678 = (inp[10]) ? 1'b1 : 1'b0;
										assign node1681 = (inp[11]) ? 1'b0 : node1682;
											assign node1682 = (inp[8]) ? 1'b1 : 1'b0;
								assign node1686 = (inp[3]) ? node1694 : node1687;
									assign node1687 = (inp[7]) ? node1689 : 1'b0;
										assign node1689 = (inp[8]) ? 1'b0 : node1690;
											assign node1690 = (inp[11]) ? 1'b0 : 1'b0;
									assign node1694 = (inp[7]) ? node1696 : 1'b1;
										assign node1696 = (inp[10]) ? 1'b0 : node1697;
											assign node1697 = (inp[11]) ? 1'b0 : 1'b1;
							assign node1701 = (inp[1]) ? node1721 : node1702;
								assign node1702 = (inp[7]) ? node1712 : node1703;
									assign node1703 = (inp[3]) ? 1'b0 : node1704;
										assign node1704 = (inp[8]) ? node1708 : node1705;
											assign node1705 = (inp[10]) ? 1'b0 : 1'b1;
											assign node1708 = (inp[11]) ? 1'b0 : 1'b1;
									assign node1712 = (inp[10]) ? 1'b0 : node1713;
										assign node1713 = (inp[11]) ? node1717 : node1714;
											assign node1714 = (inp[8]) ? 1'b1 : 1'b0;
											assign node1717 = (inp[8]) ? 1'b0 : 1'b1;
								assign node1721 = (inp[10]) ? node1729 : node1722;
									assign node1722 = (inp[3]) ? node1724 : 1'b0;
										assign node1724 = (inp[7]) ? node1726 : 1'b1;
											assign node1726 = (inp[8]) ? 1'b0 : 1'b0;
									assign node1729 = (inp[7]) ? 1'b1 : node1730;
										assign node1730 = (inp[11]) ? 1'b0 : node1731;
											assign node1731 = (inp[3]) ? 1'b0 : 1'b1;
				assign node1736 = (inp[3]) ? node1876 : node1737;
					assign node1737 = (inp[2]) ? node1803 : node1738;
						assign node1738 = (inp[8]) ? node1772 : node1739;
							assign node1739 = (inp[11]) ? node1753 : node1740;
								assign node1740 = (inp[10]) ? node1746 : node1741;
									assign node1741 = (inp[4]) ? node1743 : 1'b1;
										assign node1743 = (inp[5]) ? 1'b1 : 1'b0;
									assign node1746 = (inp[4]) ? node1748 : 1'b0;
										assign node1748 = (inp[1]) ? node1750 : 1'b1;
											assign node1750 = (inp[7]) ? 1'b1 : 1'b0;
								assign node1753 = (inp[10]) ? node1761 : node1754;
									assign node1754 = (inp[7]) ? 1'b0 : node1755;
										assign node1755 = (inp[4]) ? node1757 : 1'b0;
											assign node1757 = (inp[1]) ? 1'b0 : 1'b1;
									assign node1761 = (inp[4]) ? node1767 : node1762;
										assign node1762 = (inp[5]) ? node1764 : 1'b1;
											assign node1764 = (inp[7]) ? 1'b1 : 1'b0;
										assign node1767 = (inp[5]) ? node1769 : 1'b0;
											assign node1769 = (inp[7]) ? 1'b0 : 1'b0;
							assign node1772 = (inp[4]) ? node1788 : node1773;
								assign node1773 = (inp[10]) ? node1783 : node1774;
									assign node1774 = (inp[7]) ? node1780 : node1775;
										assign node1775 = (inp[5]) ? node1777 : 1'b1;
											assign node1777 = (inp[11]) ? 1'b0 : 1'b1;
										assign node1780 = (inp[5]) ? 1'b1 : 1'b0;
									assign node1783 = (inp[7]) ? 1'b0 : node1784;
										assign node1784 = (inp[5]) ? 1'b0 : 1'b1;
								assign node1788 = (inp[10]) ? node1796 : node1789;
									assign node1789 = (inp[11]) ? 1'b1 : node1790;
										assign node1790 = (inp[7]) ? 1'b0 : node1791;
											assign node1791 = (inp[5]) ? 1'b1 : 1'b0;
									assign node1796 = (inp[7]) ? 1'b1 : node1797;
										assign node1797 = (inp[11]) ? node1799 : 1'b1;
											assign node1799 = (inp[1]) ? 1'b0 : 1'b0;
						assign node1803 = (inp[8]) ? node1849 : node1804;
							assign node1804 = (inp[4]) ? node1826 : node1805;
								assign node1805 = (inp[10]) ? node1813 : node1806;
									assign node1806 = (inp[1]) ? 1'b0 : node1807;
										assign node1807 = (inp[7]) ? node1809 : 1'b0;
											assign node1809 = (inp[11]) ? 1'b1 : 1'b0;
									assign node1813 = (inp[1]) ? node1819 : node1814;
										assign node1814 = (inp[5]) ? 1'b0 : node1815;
											assign node1815 = (inp[11]) ? 1'b0 : 1'b0;
										assign node1819 = (inp[5]) ? node1823 : node1820;
											assign node1820 = (inp[11]) ? 1'b0 : 1'b0;
											assign node1823 = (inp[11]) ? 1'b0 : 1'b1;
								assign node1826 = (inp[10]) ? node1838 : node1827;
									assign node1827 = (inp[11]) ? node1833 : node1828;
										assign node1828 = (inp[7]) ? node1830 : 1'b1;
											assign node1830 = (inp[5]) ? 1'b0 : 1'b1;
										assign node1833 = (inp[5]) ? 1'b1 : node1834;
											assign node1834 = (inp[7]) ? 1'b1 : 1'b0;
									assign node1838 = (inp[1]) ? node1844 : node1839;
										assign node1839 = (inp[7]) ? node1841 : 1'b1;
											assign node1841 = (inp[5]) ? 1'b1 : 1'b0;
										assign node1844 = (inp[7]) ? node1846 : 1'b0;
											assign node1846 = (inp[5]) ? 1'b0 : 1'b0;
							assign node1849 = (inp[11]) ? node1861 : node1850;
								assign node1850 = (inp[7]) ? 1'b0 : node1851;
									assign node1851 = (inp[5]) ? 1'b0 : node1852;
										assign node1852 = (inp[4]) ? node1856 : node1853;
											assign node1853 = (inp[1]) ? 1'b0 : 1'b0;
											assign node1856 = (inp[1]) ? 1'b0 : 1'b1;
								assign node1861 = (inp[5]) ? node1869 : node1862;
									assign node1862 = (inp[10]) ? 1'b0 : node1863;
										assign node1863 = (inp[7]) ? node1865 : 1'b1;
											assign node1865 = (inp[4]) ? 1'b0 : 1'b1;
									assign node1869 = (inp[10]) ? 1'b1 : node1870;
										assign node1870 = (inp[4]) ? node1872 : 1'b0;
											assign node1872 = (inp[7]) ? 1'b0 : 1'b0;
					assign node1876 = (inp[5]) ? node1934 : node1877;
						assign node1877 = (inp[1]) ? node1903 : node1878;
							assign node1878 = (inp[7]) ? node1890 : node1879;
								assign node1879 = (inp[11]) ? 1'b1 : node1880;
									assign node1880 = (inp[10]) ? node1886 : node1881;
										assign node1881 = (inp[4]) ? 1'b1 : node1882;
											assign node1882 = (inp[2]) ? 1'b0 : 1'b1;
										assign node1886 = (inp[2]) ? 1'b1 : 1'b0;
								assign node1890 = (inp[8]) ? node1900 : node1891;
									assign node1891 = (inp[11]) ? 1'b1 : node1892;
										assign node1892 = (inp[4]) ? node1896 : node1893;
											assign node1893 = (inp[2]) ? 1'b0 : 1'b0;
											assign node1896 = (inp[10]) ? 1'b0 : 1'b1;
									assign node1900 = (inp[2]) ? 1'b1 : 1'b0;
							assign node1903 = (inp[10]) ? node1919 : node1904;
								assign node1904 = (inp[4]) ? node1912 : node1905;
									assign node1905 = (inp[7]) ? node1907 : 1'b0;
										assign node1907 = (inp[11]) ? node1909 : 1'b0;
											assign node1909 = (inp[2]) ? 1'b1 : 1'b0;
									assign node1912 = (inp[2]) ? 1'b0 : node1913;
										assign node1913 = (inp[7]) ? node1915 : 1'b1;
											assign node1915 = (inp[8]) ? 1'b1 : 1'b0;
								assign node1919 = (inp[2]) ? node1927 : node1920;
									assign node1920 = (inp[11]) ? 1'b1 : node1921;
										assign node1921 = (inp[8]) ? 1'b0 : node1922;
											assign node1922 = (inp[4]) ? 1'b0 : 1'b0;
									assign node1927 = (inp[11]) ? node1929 : 1'b1;
										assign node1929 = (inp[7]) ? node1931 : 1'b0;
											assign node1931 = (inp[8]) ? 1'b1 : 1'b0;
						assign node1934 = (inp[1]) ? node1958 : node1935;
							assign node1935 = (inp[11]) ? node1949 : node1936;
								assign node1936 = (inp[10]) ? node1942 : node1937;
									assign node1937 = (inp[7]) ? node1939 : 1'b1;
										assign node1939 = (inp[2]) ? 1'b1 : 1'b0;
									assign node1942 = (inp[7]) ? node1944 : 1'b0;
										assign node1944 = (inp[4]) ? 1'b1 : node1945;
											assign node1945 = (inp[2]) ? 1'b0 : 1'b1;
								assign node1949 = (inp[7]) ? node1951 : 1'b0;
									assign node1951 = (inp[2]) ? node1953 : 1'b0;
										assign node1953 = (inp[8]) ? node1955 : 1'b0;
											assign node1955 = (inp[4]) ? 1'b0 : 1'b0;
							assign node1958 = (inp[11]) ? node1974 : node1959;
								assign node1959 = (inp[10]) ? node1967 : node1960;
									assign node1960 = (inp[7]) ? 1'b1 : node1961;
										assign node1961 = (inp[4]) ? node1963 : 1'b0;
											assign node1963 = (inp[2]) ? 1'b1 : 1'b0;
									assign node1967 = (inp[2]) ? node1971 : node1968;
										assign node1968 = (inp[4]) ? 1'b1 : 1'b0;
										assign node1971 = (inp[4]) ? 1'b0 : 1'b1;
								assign node1974 = (inp[7]) ? node1980 : node1975;
									assign node1975 = (inp[4]) ? node1977 : 1'b1;
										assign node1977 = (inp[2]) ? 1'b0 : 1'b1;
									assign node1980 = (inp[2]) ? node1988 : node1981;
										assign node1981 = (inp[10]) ? node1985 : node1982;
											assign node1982 = (inp[8]) ? 1'b0 : 1'b0;
											assign node1985 = (inp[4]) ? 1'b0 : 1'b0;
										assign node1988 = (inp[4]) ? node1990 : 1'b1;
											assign node1990 = (inp[10]) ? 1'b0 : 1'b0;

endmodule