module dtc_split125_bm22 (
	input  wire [11-1:0] inp,
	output wire [11-1:0] outp
);

	wire [11-1:0] node1;
	wire [11-1:0] node2;
	wire [11-1:0] node3;
	wire [11-1:0] node4;
	wire [11-1:0] node5;
	wire [11-1:0] node6;
	wire [11-1:0] node7;
	wire [11-1:0] node12;
	wire [11-1:0] node13;
	wire [11-1:0] node15;
	wire [11-1:0] node16;
	wire [11-1:0] node21;
	wire [11-1:0] node22;
	wire [11-1:0] node23;
	wire [11-1:0] node25;
	wire [11-1:0] node28;
	wire [11-1:0] node30;
	wire [11-1:0] node32;
	wire [11-1:0] node35;
	wire [11-1:0] node36;
	wire [11-1:0] node37;
	wire [11-1:0] node40;
	wire [11-1:0] node41;
	wire [11-1:0] node43;
	wire [11-1:0] node47;
	wire [11-1:0] node49;
	wire [11-1:0] node52;
	wire [11-1:0] node53;
	wire [11-1:0] node54;
	wire [11-1:0] node55;
	wire [11-1:0] node58;
	wire [11-1:0] node61;
	wire [11-1:0] node63;
	wire [11-1:0] node65;
	wire [11-1:0] node68;
	wire [11-1:0] node69;
	wire [11-1:0] node70;
	wire [11-1:0] node71;
	wire [11-1:0] node72;
	wire [11-1:0] node76;
	wire [11-1:0] node79;
	wire [11-1:0] node81;
	wire [11-1:0] node82;
	wire [11-1:0] node85;
	wire [11-1:0] node88;
	wire [11-1:0] node89;
	wire [11-1:0] node90;
	wire [11-1:0] node93;
	wire [11-1:0] node94;
	wire [11-1:0] node98;
	wire [11-1:0] node101;
	wire [11-1:0] node102;
	wire [11-1:0] node103;
	wire [11-1:0] node104;
	wire [11-1:0] node105;
	wire [11-1:0] node106;
	wire [11-1:0] node108;
	wire [11-1:0] node111;
	wire [11-1:0] node114;
	wire [11-1:0] node116;
	wire [11-1:0] node119;
	wire [11-1:0] node120;
	wire [11-1:0] node124;
	wire [11-1:0] node125;
	wire [11-1:0] node126;
	wire [11-1:0] node127;
	wire [11-1:0] node129;
	wire [11-1:0] node134;
	wire [11-1:0] node135;
	wire [11-1:0] node138;
	wire [11-1:0] node141;
	wire [11-1:0] node142;
	wire [11-1:0] node144;
	wire [11-1:0] node145;
	wire [11-1:0] node147;
	wire [11-1:0] node148;
	wire [11-1:0] node149;
	wire [11-1:0] node154;
	wire [11-1:0] node155;
	wire [11-1:0] node159;
	wire [11-1:0] node160;
	wire [11-1:0] node161;
	wire [11-1:0] node164;
	wire [11-1:0] node166;
	wire [11-1:0] node169;
	wire [11-1:0] node170;
	wire [11-1:0] node173;
	wire [11-1:0] node175;
	wire [11-1:0] node177;
	wire [11-1:0] node180;
	wire [11-1:0] node181;
	wire [11-1:0] node182;
	wire [11-1:0] node183;
	wire [11-1:0] node184;
	wire [11-1:0] node185;
	wire [11-1:0] node187;
	wire [11-1:0] node189;
	wire [11-1:0] node190;
	wire [11-1:0] node194;
	wire [11-1:0] node197;
	wire [11-1:0] node198;
	wire [11-1:0] node199;
	wire [11-1:0] node203;
	wire [11-1:0] node204;
	wire [11-1:0] node205;
	wire [11-1:0] node208;
	wire [11-1:0] node212;
	wire [11-1:0] node213;
	wire [11-1:0] node214;
	wire [11-1:0] node215;
	wire [11-1:0] node219;
	wire [11-1:0] node221;
	wire [11-1:0] node222;
	wire [11-1:0] node226;
	wire [11-1:0] node227;
	wire [11-1:0] node229;
	wire [11-1:0] node231;
	wire [11-1:0] node234;
	wire [11-1:0] node235;
	wire [11-1:0] node237;
	wire [11-1:0] node241;
	wire [11-1:0] node242;
	wire [11-1:0] node243;
	wire [11-1:0] node244;
	wire [11-1:0] node246;
	wire [11-1:0] node250;
	wire [11-1:0] node251;
	wire [11-1:0] node254;
	wire [11-1:0] node256;
	wire [11-1:0] node259;
	wire [11-1:0] node260;
	wire [11-1:0] node261;
	wire [11-1:0] node262;
	wire [11-1:0] node266;
	wire [11-1:0] node269;
	wire [11-1:0] node270;
	wire [11-1:0] node272;
	wire [11-1:0] node274;
	wire [11-1:0] node276;
	wire [11-1:0] node280;
	wire [11-1:0] node281;
	wire [11-1:0] node282;
	wire [11-1:0] node283;
	wire [11-1:0] node284;
	wire [11-1:0] node288;
	wire [11-1:0] node289;
	wire [11-1:0] node291;
	wire [11-1:0] node293;
	wire [11-1:0] node294;
	wire [11-1:0] node298;
	wire [11-1:0] node299;
	wire [11-1:0] node300;
	wire [11-1:0] node301;
	wire [11-1:0] node306;
	wire [11-1:0] node309;
	wire [11-1:0] node310;
	wire [11-1:0] node311;
	wire [11-1:0] node312;
	wire [11-1:0] node315;
	wire [11-1:0] node316;
	wire [11-1:0] node320;
	wire [11-1:0] node321;
	wire [11-1:0] node325;
	wire [11-1:0] node326;
	wire [11-1:0] node329;
	wire [11-1:0] node331;
	wire [11-1:0] node332;
	wire [11-1:0] node336;
	wire [11-1:0] node337;
	wire [11-1:0] node338;
	wire [11-1:0] node339;
	wire [11-1:0] node340;
	wire [11-1:0] node342;
	wire [11-1:0] node346;
	wire [11-1:0] node348;
	wire [11-1:0] node349;
	wire [11-1:0] node353;
	wire [11-1:0] node354;
	wire [11-1:0] node356;
	wire [11-1:0] node360;
	wire [11-1:0] node361;
	wire [11-1:0] node362;
	wire [11-1:0] node364;
	wire [11-1:0] node365;
	wire [11-1:0] node367;
	wire [11-1:0] node371;
	wire [11-1:0] node374;
	wire [11-1:0] node376;

	assign outp = (inp[4]) ? node180 : node1;
		assign node1 = (inp[0]) ? node101 : node2;
			assign node2 = (inp[6]) ? node52 : node3;
				assign node3 = (inp[5]) ? node21 : node4;
					assign node4 = (inp[3]) ? node12 : node5;
						assign node5 = (inp[7]) ? 11'b00011111111 : node6;
							assign node6 = (inp[1]) ? 11'b00011111111 : node7;
								assign node7 = (inp[9]) ? 11'b00111111111 : 11'b01111111111;
						assign node12 = (inp[10]) ? 11'b00001111111 : node13;
							assign node13 = (inp[9]) ? node15 : 11'b00011111111;
								assign node15 = (inp[2]) ? 11'b00001111111 : node16;
									assign node16 = (inp[8]) ? 11'b00001111111 : 11'b00011111111;
					assign node21 = (inp[2]) ? node35 : node22;
						assign node22 = (inp[1]) ? node28 : node23;
							assign node23 = (inp[10]) ? node25 : 11'b00011111111;
								assign node25 = (inp[8]) ? 11'b00001111111 : 11'b00011111111;
							assign node28 = (inp[10]) ? node30 : 11'b00001111111;
								assign node30 = (inp[7]) ? node32 : 11'b00011111111;
									assign node32 = (inp[3]) ? 11'b00000111111 : 11'b00001111111;
						assign node35 = (inp[1]) ? node47 : node36;
							assign node36 = (inp[9]) ? node40 : node37;
								assign node37 = (inp[3]) ? 11'b00001111111 : 11'b00011111111;
								assign node40 = (inp[7]) ? 11'b00000111111 : node41;
									assign node41 = (inp[3]) ? node43 : 11'b00001111111;
										assign node43 = (inp[8]) ? 11'b00000111111 : 11'b00001111111;
							assign node47 = (inp[9]) ? node49 : 11'b00000011111;
								assign node49 = (inp[8]) ? 11'b00000001111 : 11'b00000011111;
				assign node52 = (inp[9]) ? node68 : node53;
					assign node53 = (inp[10]) ? node61 : node54;
						assign node54 = (inp[8]) ? node58 : node55;
							assign node55 = (inp[7]) ? 11'b00001111111 : 11'b00011111111;
							assign node58 = (inp[5]) ? 11'b00001111111 : 11'b00000111111;
						assign node61 = (inp[1]) ? node63 : 11'b00001111111;
							assign node63 = (inp[7]) ? node65 : 11'b00000111111;
								assign node65 = (inp[3]) ? 11'b00000011111 : 11'b00000111111;
					assign node68 = (inp[2]) ? node88 : node69;
						assign node69 = (inp[7]) ? node79 : node70;
							assign node70 = (inp[10]) ? node76 : node71;
								assign node71 = (inp[8]) ? 11'b00000111111 : node72;
									assign node72 = (inp[1]) ? 11'b00001111111 : 11'b00011111111;
								assign node76 = (inp[3]) ? 11'b00000011111 : 11'b00000111111;
							assign node79 = (inp[5]) ? node81 : 11'b00000111111;
								assign node81 = (inp[1]) ? node85 : node82;
									assign node82 = (inp[10]) ? 11'b00000011111 : 11'b00000111111;
									assign node85 = (inp[10]) ? 11'b00000001111 : 11'b00000011111;
						assign node88 = (inp[5]) ? node98 : node89;
							assign node89 = (inp[3]) ? node93 : node90;
								assign node90 = (inp[10]) ? 11'b00000011111 : 11'b00000111111;
								assign node93 = (inp[1]) ? 11'b00000011111 : node94;
									assign node94 = (inp[10]) ? 11'b00000001111 : 11'b00000011111;
							assign node98 = (inp[3]) ? 11'b00000000111 : 11'b00000001111;
			assign node101 = (inp[5]) ? node141 : node102;
				assign node102 = (inp[3]) ? node124 : node103;
					assign node103 = (inp[8]) ? node119 : node104;
						assign node104 = (inp[2]) ? node114 : node105;
							assign node105 = (inp[7]) ? node111 : node106;
								assign node106 = (inp[10]) ? node108 : 11'b00011111111;
									assign node108 = (inp[9]) ? 11'b00001111111 : 11'b00011111111;
								assign node111 = (inp[6]) ? 11'b00011111111 : 11'b00111111111;
							assign node114 = (inp[6]) ? node116 : 11'b00001111111;
								assign node116 = (inp[9]) ? 11'b00000111111 : 11'b00001111111;
						assign node119 = (inp[10]) ? 11'b00000111111 : node120;
							assign node120 = (inp[7]) ? 11'b00000111111 : 11'b00001111111;
					assign node124 = (inp[6]) ? node134 : node125;
						assign node125 = (inp[9]) ? 11'b00001111111 : node126;
							assign node126 = (inp[1]) ? 11'b00000111111 : node127;
								assign node127 = (inp[8]) ? node129 : 11'b00000111111;
									assign node129 = (inp[10]) ? 11'b00000011111 : 11'b00000111111;
						assign node134 = (inp[1]) ? node138 : node135;
							assign node135 = (inp[9]) ? 11'b00000011111 : 11'b00000111111;
							assign node138 = (inp[9]) ? 11'b00000001111 : 11'b00000011111;
				assign node141 = (inp[9]) ? node159 : node142;
					assign node142 = (inp[2]) ? node144 : 11'b00000111111;
						assign node144 = (inp[3]) ? node154 : node145;
							assign node145 = (inp[8]) ? node147 : 11'b00000111111;
								assign node147 = (inp[1]) ? 11'b00000001111 : node148;
									assign node148 = (inp[6]) ? 11'b00000011111 : node149;
										assign node149 = (inp[7]) ? 11'b00000011111 : 11'b00000111111;
							assign node154 = (inp[10]) ? 11'b00000001111 : node155;
								assign node155 = (inp[6]) ? 11'b00000001111 : 11'b00000011111;
					assign node159 = (inp[1]) ? node169 : node160;
						assign node160 = (inp[3]) ? node164 : node161;
							assign node161 = (inp[10]) ? 11'b00000011111 : 11'b00000111111;
							assign node164 = (inp[10]) ? node166 : 11'b00000001111;
								assign node166 = (inp[8]) ? 11'b00000001111 : 11'b00000000111;
						assign node169 = (inp[6]) ? node173 : node170;
							assign node170 = (inp[7]) ? 11'b00000011111 : 11'b00000000111;
							assign node173 = (inp[10]) ? node175 : 11'b00000000111;
								assign node175 = (inp[3]) ? node177 : 11'b00000000111;
									assign node177 = (inp[8]) ? 11'b00000000001 : 11'b00000000111;
		assign node180 = (inp[3]) ? node280 : node181;
			assign node181 = (inp[8]) ? node241 : node182;
				assign node182 = (inp[10]) ? node212 : node183;
					assign node183 = (inp[9]) ? node197 : node184;
						assign node184 = (inp[6]) ? node194 : node185;
							assign node185 = (inp[7]) ? node187 : 11'b00111111111;
								assign node187 = (inp[0]) ? node189 : 11'b00011111111;
									assign node189 = (inp[2]) ? 11'b00001111111 : node190;
										assign node190 = (inp[1]) ? 11'b00001111111 : 11'b00011111111;
							assign node194 = (inp[7]) ? 11'b00000111111 : 11'b00001111111;
						assign node197 = (inp[0]) ? node203 : node198;
							assign node198 = (inp[1]) ? 11'b00000111111 : node199;
								assign node199 = (inp[7]) ? 11'b00001111111 : 11'b00011111111;
							assign node203 = (inp[7]) ? 11'b00000011111 : node204;
								assign node204 = (inp[1]) ? node208 : node205;
									assign node205 = (inp[2]) ? 11'b00000111111 : 11'b00001111111;
									assign node208 = (inp[2]) ? 11'b00000011111 : 11'b00000111111;
					assign node212 = (inp[0]) ? node226 : node213;
						assign node213 = (inp[1]) ? node219 : node214;
							assign node214 = (inp[5]) ? 11'b00000111111 : node215;
								assign node215 = (inp[6]) ? 11'b00000111111 : 11'b00001111111;
							assign node219 = (inp[7]) ? node221 : 11'b00000111111;
								assign node221 = (inp[6]) ? 11'b00000011111 : node222;
									assign node222 = (inp[2]) ? 11'b00000011111 : 11'b00000111111;
						assign node226 = (inp[5]) ? node234 : node227;
							assign node227 = (inp[1]) ? node229 : 11'b00000011111;
								assign node229 = (inp[9]) ? node231 : 11'b00000011111;
									assign node231 = (inp[2]) ? 11'b00000001111 : 11'b00000011111;
							assign node234 = (inp[9]) ? 11'b00000011111 : node235;
								assign node235 = (inp[7]) ? node237 : 11'b00000111111;
									assign node237 = (inp[2]) ? 11'b00000011111 : 11'b00000111111;
				assign node241 = (inp[1]) ? node259 : node242;
					assign node242 = (inp[9]) ? node250 : node243;
						assign node243 = (inp[2]) ? 11'b00000011111 : node244;
							assign node244 = (inp[0]) ? node246 : 11'b00001111111;
								assign node246 = (inp[10]) ? 11'b00001111111 : 11'b00000111111;
						assign node250 = (inp[6]) ? node254 : node251;
							assign node251 = (inp[10]) ? 11'b00000011111 : 11'b00000111111;
							assign node254 = (inp[7]) ? node256 : 11'b00000011111;
								assign node256 = (inp[2]) ? 11'b00000001111 : 11'b00000011111;
					assign node259 = (inp[6]) ? node269 : node260;
						assign node260 = (inp[5]) ? node266 : node261;
							assign node261 = (inp[10]) ? 11'b00000011111 : node262;
								assign node262 = (inp[2]) ? 11'b00000011111 : 11'b00000111111;
							assign node266 = (inp[7]) ? 11'b00000001111 : 11'b00000011111;
						assign node269 = (inp[5]) ? 11'b00000001111 : node270;
							assign node270 = (inp[0]) ? node272 : 11'b00000011111;
								assign node272 = (inp[2]) ? node274 : 11'b00000111111;
									assign node274 = (inp[7]) ? node276 : 11'b00000001111;
										assign node276 = (inp[9]) ? 11'b00000000011 : 11'b00000000111;
			assign node280 = (inp[1]) ? node336 : node281;
				assign node281 = (inp[0]) ? node309 : node282;
					assign node282 = (inp[5]) ? node288 : node283;
						assign node283 = (inp[10]) ? 11'b00000111111 : node284;
							assign node284 = (inp[6]) ? 11'b00001111111 : 11'b00011111111;
						assign node288 = (inp[6]) ? node298 : node289;
							assign node289 = (inp[10]) ? node291 : 11'b00001111111;
								assign node291 = (inp[7]) ? node293 : 11'b00000111111;
									assign node293 = (inp[9]) ? 11'b00000011111 : node294;
										assign node294 = (inp[2]) ? 11'b00000011111 : 11'b00000111111;
							assign node298 = (inp[9]) ? node306 : node299;
								assign node299 = (inp[7]) ? 11'b00000011111 : node300;
									assign node300 = (inp[10]) ? 11'b00000011111 : node301;
										assign node301 = (inp[2]) ? 11'b00000011111 : 11'b00000111111;
								assign node306 = (inp[10]) ? 11'b00000000111 : 11'b00000011111;
					assign node309 = (inp[5]) ? node325 : node310;
						assign node310 = (inp[6]) ? node320 : node311;
							assign node311 = (inp[8]) ? node315 : node312;
								assign node312 = (inp[9]) ? 11'b00000111111 : 11'b00001111111;
								assign node315 = (inp[10]) ? 11'b00000011111 : node316;
									assign node316 = (inp[9]) ? 11'b00000011111 : 11'b00000111111;
							assign node320 = (inp[7]) ? 11'b00000011111 : node321;
								assign node321 = (inp[10]) ? 11'b00000001111 : 11'b00000011111;
						assign node325 = (inp[8]) ? node329 : node326;
							assign node326 = (inp[9]) ? 11'b00000001111 : 11'b00000111111;
							assign node329 = (inp[10]) ? node331 : 11'b00000001111;
								assign node331 = (inp[7]) ? 11'b00000000111 : node332;
									assign node332 = (inp[2]) ? 11'b00000000111 : 11'b00000001111;
				assign node336 = (inp[6]) ? node360 : node337;
					assign node337 = (inp[2]) ? node353 : node338;
						assign node338 = (inp[7]) ? node346 : node339;
							assign node339 = (inp[8]) ? 11'b00000011111 : node340;
								assign node340 = (inp[5]) ? node342 : 11'b00001111111;
									assign node342 = (inp[10]) ? 11'b00000011111 : 11'b00000111111;
							assign node346 = (inp[0]) ? node348 : 11'b00000011111;
								assign node348 = (inp[8]) ? 11'b00000001111 : node349;
									assign node349 = (inp[9]) ? 11'b00000011111 : 11'b00000001111;
						assign node353 = (inp[5]) ? 11'b00000000011 : node354;
							assign node354 = (inp[8]) ? node356 : 11'b00000011111;
								assign node356 = (inp[7]) ? 11'b00000000111 : 11'b00000001111;
					assign node360 = (inp[0]) ? node374 : node361;
						assign node361 = (inp[9]) ? node371 : node362;
							assign node362 = (inp[2]) ? node364 : 11'b00000011111;
								assign node364 = (inp[5]) ? 11'b00000001111 : node365;
									assign node365 = (inp[10]) ? node367 : 11'b00000011111;
										assign node367 = (inp[7]) ? 11'b00000001111 : 11'b00000011111;
							assign node371 = (inp[5]) ? 11'b00000000111 : 11'b00000001111;
						assign node374 = (inp[8]) ? node376 : 11'b00000000111;
							assign node376 = (inp[2]) ? 11'b00000000011 : 11'b00000000111;

endmodule