module dtc_split875_bm96 (
	input  wire [12-1:0] inp,
	output wire [3-1:0] outp
);

	wire [3-1:0] node2;
	wire [3-1:0] node3;
	wire [3-1:0] node5;
	wire [3-1:0] node7;
	wire [3-1:0] node9;
	wire [3-1:0] node11;
	wire [3-1:0] node12;
	wire [3-1:0] node14;
	wire [3-1:0] node18;
	wire [3-1:0] node19;
	wire [3-1:0] node20;
	wire [3-1:0] node21;
	wire [3-1:0] node23;
	wire [3-1:0] node24;
	wire [3-1:0] node27;
	wire [3-1:0] node31;
	wire [3-1:0] node32;
	wire [3-1:0] node33;
	wire [3-1:0] node34;
	wire [3-1:0] node35;
	wire [3-1:0] node36;
	wire [3-1:0] node39;
	wire [3-1:0] node42;
	wire [3-1:0] node44;
	wire [3-1:0] node46;
	wire [3-1:0] node49;
	wire [3-1:0] node50;
	wire [3-1:0] node51;
	wire [3-1:0] node55;
	wire [3-1:0] node56;
	wire [3-1:0] node57;
	wire [3-1:0] node60;
	wire [3-1:0] node63;
	wire [3-1:0] node64;
	wire [3-1:0] node67;
	wire [3-1:0] node70;
	wire [3-1:0] node71;
	wire [3-1:0] node73;
	wire [3-1:0] node75;
	wire [3-1:0] node77;
	wire [3-1:0] node80;
	wire [3-1:0] node81;
	wire [3-1:0] node83;
	wire [3-1:0] node86;
	wire [3-1:0] node87;
	wire [3-1:0] node88;
	wire [3-1:0] node92;
	wire [3-1:0] node94;
	wire [3-1:0] node97;
	wire [3-1:0] node98;
	wire [3-1:0] node100;
	wire [3-1:0] node102;
	wire [3-1:0] node104;
	wire [3-1:0] node106;
	wire [3-1:0] node109;
	wire [3-1:0] node110;
	wire [3-1:0] node111;
	wire [3-1:0] node112;
	wire [3-1:0] node113;
	wire [3-1:0] node115;
	wire [3-1:0] node118;
	wire [3-1:0] node120;
	wire [3-1:0] node123;
	wire [3-1:0] node124;
	wire [3-1:0] node127;
	wire [3-1:0] node130;
	wire [3-1:0] node132;
	wire [3-1:0] node133;
	wire [3-1:0] node137;
	wire [3-1:0] node139;
	wire [3-1:0] node141;
	wire [3-1:0] node142;
	wire [3-1:0] node146;
	wire [3-1:0] node147;
	wire [3-1:0] node148;
	wire [3-1:0] node149;
	wire [3-1:0] node151;
	wire [3-1:0] node152;
	wire [3-1:0] node153;
	wire [3-1:0] node154;
	wire [3-1:0] node157;
	wire [3-1:0] node160;
	wire [3-1:0] node161;
	wire [3-1:0] node164;
	wire [3-1:0] node167;
	wire [3-1:0] node168;
	wire [3-1:0] node170;
	wire [3-1:0] node172;
	wire [3-1:0] node175;
	wire [3-1:0] node176;
	wire [3-1:0] node177;
	wire [3-1:0] node180;
	wire [3-1:0] node183;
	wire [3-1:0] node184;
	wire [3-1:0] node187;
	wire [3-1:0] node190;
	wire [3-1:0] node191;
	wire [3-1:0] node192;
	wire [3-1:0] node195;
	wire [3-1:0] node198;
	wire [3-1:0] node199;
	wire [3-1:0] node202;
	wire [3-1:0] node205;
	wire [3-1:0] node206;
	wire [3-1:0] node207;
	wire [3-1:0] node208;
	wire [3-1:0] node209;
	wire [3-1:0] node212;
	wire [3-1:0] node214;
	wire [3-1:0] node217;
	wire [3-1:0] node218;
	wire [3-1:0] node222;
	wire [3-1:0] node223;
	wire [3-1:0] node226;
	wire [3-1:0] node228;
	wire [3-1:0] node231;
	wire [3-1:0] node232;
	wire [3-1:0] node234;
	wire [3-1:0] node236;
	wire [3-1:0] node238;
	wire [3-1:0] node241;
	wire [3-1:0] node242;
	wire [3-1:0] node245;
	wire [3-1:0] node247;
	wire [3-1:0] node250;
	wire [3-1:0] node251;
	wire [3-1:0] node252;
	wire [3-1:0] node254;
	wire [3-1:0] node256;
	wire [3-1:0] node258;
	wire [3-1:0] node260;
	wire [3-1:0] node263;
	wire [3-1:0] node264;
	wire [3-1:0] node265;
	wire [3-1:0] node266;
	wire [3-1:0] node270;
	wire [3-1:0] node272;
	wire [3-1:0] node274;
	wire [3-1:0] node278;
	wire [3-1:0] node279;
	wire [3-1:0] node280;
	wire [3-1:0] node282;
	wire [3-1:0] node284;
	wire [3-1:0] node286;
	wire [3-1:0] node289;
	wire [3-1:0] node291;
	wire [3-1:0] node293;
	wire [3-1:0] node295;
	wire [3-1:0] node298;
	wire [3-1:0] node299;
	wire [3-1:0] node300;
	wire [3-1:0] node301;
	wire [3-1:0] node304;
	wire [3-1:0] node307;
	wire [3-1:0] node308;
	wire [3-1:0] node310;
	wire [3-1:0] node314;
	wire [3-1:0] node316;
	wire [3-1:0] node317;
	wire [3-1:0] node319;

	assign outp = (inp[6]) ? node2 : 3'b000;
		assign node2 = (inp[7]) ? node18 : node3;
			assign node3 = (inp[2]) ? node5 : 3'b000;
				assign node5 = (inp[1]) ? node7 : 3'b000;
					assign node7 = (inp[8]) ? node9 : 3'b000;
						assign node9 = (inp[4]) ? node11 : 3'b000;
							assign node11 = (inp[9]) ? 3'b000 : node12;
								assign node12 = (inp[3]) ? node14 : 3'b000;
									assign node14 = (inp[10]) ? 3'b000 : 3'b100;
			assign node18 = (inp[3]) ? node146 : node19;
				assign node19 = (inp[4]) ? node31 : node20;
					assign node20 = (inp[1]) ? 3'b011 : node21;
						assign node21 = (inp[9]) ? node23 : 3'b011;
							assign node23 = (inp[10]) ? node27 : node24;
								assign node24 = (inp[5]) ? 3'b011 : 3'b111;
								assign node27 = (inp[5]) ? 3'b101 : 3'b011;
					assign node31 = (inp[1]) ? node97 : node32;
						assign node32 = (inp[0]) ? node70 : node33;
							assign node33 = (inp[9]) ? node49 : node34;
								assign node34 = (inp[11]) ? node42 : node35;
									assign node35 = (inp[8]) ? node39 : node36;
										assign node36 = (inp[10]) ? 3'b010 : 3'b001;
										assign node39 = (inp[10]) ? 3'b001 : 3'b010;
									assign node42 = (inp[8]) ? node44 : 3'b010;
										assign node44 = (inp[2]) ? node46 : 3'b010;
											assign node46 = (inp[10]) ? 3'b010 : 3'b001;
								assign node49 = (inp[5]) ? node55 : node50;
									assign node50 = (inp[10]) ? 3'b001 : node51;
										assign node51 = (inp[11]) ? 3'b001 : 3'b010;
									assign node55 = (inp[8]) ? node63 : node56;
										assign node56 = (inp[11]) ? node60 : node57;
											assign node57 = (inp[10]) ? 3'b001 : 3'b010;
											assign node60 = (inp[10]) ? 3'b010 : 3'b001;
										assign node63 = (inp[11]) ? node67 : node64;
											assign node64 = (inp[10]) ? 3'b001 : 3'b010;
											assign node67 = (inp[10]) ? 3'b010 : 3'b001;
							assign node70 = (inp[9]) ? node80 : node71;
								assign node71 = (inp[10]) ? node73 : 3'b001;
									assign node73 = (inp[8]) ? node75 : 3'b001;
										assign node75 = (inp[11]) ? node77 : 3'b001;
											assign node77 = (inp[5]) ? 3'b010 : 3'b001;
								assign node80 = (inp[11]) ? node86 : node81;
									assign node81 = (inp[10]) ? node83 : 3'b110;
										assign node83 = (inp[5]) ? 3'b001 : 3'b101;
									assign node86 = (inp[5]) ? node92 : node87;
										assign node87 = (inp[10]) ? 3'b001 : node88;
											assign node88 = (inp[8]) ? 3'b101 : 3'b001;
										assign node92 = (inp[10]) ? node94 : 3'b001;
											assign node94 = (inp[8]) ? 3'b110 : 3'b010;
						assign node97 = (inp[0]) ? node109 : node98;
							assign node98 = (inp[5]) ? node100 : 3'b010;
								assign node100 = (inp[10]) ? node102 : 3'b010;
									assign node102 = (inp[9]) ? node104 : 3'b010;
										assign node104 = (inp[8]) ? node106 : 3'b010;
											assign node106 = (inp[11]) ? 3'b001 : 3'b010;
							assign node109 = (inp[9]) ? node137 : node110;
								assign node110 = (inp[11]) ? node130 : node111;
									assign node111 = (inp[5]) ? node123 : node112;
										assign node112 = (inp[2]) ? node118 : node113;
											assign node113 = (inp[10]) ? node115 : 3'b010;
												assign node115 = (inp[8]) ? 3'b010 : 3'b001;
											assign node118 = (inp[10]) ? node120 : 3'b001;
												assign node120 = (inp[8]) ? 3'b010 : 3'b001;
										assign node123 = (inp[8]) ? node127 : node124;
											assign node124 = (inp[10]) ? 3'b001 : 3'b010;
											assign node127 = (inp[10]) ? 3'b010 : 3'b001;
									assign node130 = (inp[2]) ? node132 : 3'b001;
										assign node132 = (inp[10]) ? 3'b001 : node133;
											assign node133 = (inp[8]) ? 3'b010 : 3'b001;
								assign node137 = (inp[8]) ? node139 : 3'b010;
									assign node139 = (inp[2]) ? node141 : 3'b010;
										assign node141 = (inp[10]) ? 3'b010 : node142;
											assign node142 = (inp[11]) ? 3'b010 : 3'b001;
				assign node146 = (inp[1]) ? node250 : node147;
					assign node147 = (inp[4]) ? node205 : node148;
						assign node148 = (inp[10]) ? node190 : node149;
							assign node149 = (inp[9]) ? node151 : 3'b111;
								assign node151 = (inp[5]) ? node167 : node152;
									assign node152 = (inp[2]) ? node160 : node153;
										assign node153 = (inp[0]) ? node157 : node154;
											assign node154 = (inp[11]) ? 3'b111 : 3'b110;
											assign node157 = (inp[11]) ? 3'b110 : 3'b111;
										assign node160 = (inp[11]) ? node164 : node161;
											assign node161 = (inp[0]) ? 3'b111 : 3'b110;
											assign node164 = (inp[0]) ? 3'b110 : 3'b111;
									assign node167 = (inp[8]) ? node175 : node168;
										assign node168 = (inp[2]) ? node170 : 3'b111;
											assign node170 = (inp[0]) ? node172 : 3'b111;
												assign node172 = (inp[11]) ? 3'b110 : 3'b111;
										assign node175 = (inp[2]) ? node183 : node176;
											assign node176 = (inp[11]) ? node180 : node177;
												assign node177 = (inp[0]) ? 3'b111 : 3'b110;
												assign node180 = (inp[0]) ? 3'b110 : 3'b111;
											assign node183 = (inp[0]) ? node187 : node184;
												assign node184 = (inp[11]) ? 3'b111 : 3'b110;
												assign node187 = (inp[11]) ? 3'b110 : 3'b111;
							assign node190 = (inp[5]) ? node198 : node191;
								assign node191 = (inp[0]) ? node195 : node192;
									assign node192 = (inp[9]) ? 3'b111 : 3'b110;
									assign node195 = (inp[9]) ? 3'b110 : 3'b111;
								assign node198 = (inp[9]) ? node202 : node199;
									assign node199 = (inp[0]) ? 3'b111 : 3'b110;
									assign node202 = (inp[0]) ? 3'b010 : 3'b011;
						assign node205 = (inp[0]) ? node231 : node206;
							assign node206 = (inp[9]) ? node222 : node207;
								assign node207 = (inp[10]) ? node217 : node208;
									assign node208 = (inp[11]) ? node212 : node209;
										assign node209 = (inp[8]) ? 3'b011 : 3'b111;
										assign node212 = (inp[8]) ? node214 : 3'b011;
											assign node214 = (inp[2]) ? 3'b111 : 3'b011;
									assign node217 = (inp[11]) ? 3'b001 : node218;
										assign node218 = (inp[8]) ? 3'b101 : 3'b001;
								assign node222 = (inp[11]) ? node226 : node223;
									assign node223 = (inp[10]) ? 3'b110 : 3'b001;
									assign node226 = (inp[5]) ? node228 : 3'b110;
										assign node228 = (inp[10]) ? 3'b010 : 3'b110;
							assign node231 = (inp[9]) ? node241 : node232;
								assign node232 = (inp[8]) ? node234 : 3'b110;
									assign node234 = (inp[11]) ? node236 : 3'b110;
										assign node236 = (inp[10]) ? node238 : 3'b110;
											assign node238 = (inp[5]) ? 3'b010 : 3'b110;
								assign node241 = (inp[10]) ? node245 : node242;
									assign node242 = (inp[11]) ? 3'b100 : 3'b010;
									assign node245 = (inp[11]) ? node247 : 3'b100;
										assign node247 = (inp[5]) ? 3'b000 : 3'b100;
					assign node250 = (inp[4]) ? node278 : node251;
						assign node251 = (inp[0]) ? node263 : node252;
							assign node252 = (inp[9]) ? node254 : 3'b100;
								assign node254 = (inp[5]) ? node256 : 3'b101;
									assign node256 = (inp[8]) ? node258 : 3'b101;
										assign node258 = (inp[10]) ? node260 : 3'b101;
											assign node260 = (inp[11]) ? 3'b100 : 3'b101;
							assign node263 = (inp[9]) ? 3'b100 : node264;
								assign node264 = (inp[11]) ? node270 : node265;
									assign node265 = (inp[8]) ? 3'b101 : node266;
										assign node266 = (inp[10]) ? 3'b100 : 3'b101;
									assign node270 = (inp[2]) ? node272 : 3'b100;
										assign node272 = (inp[8]) ? node274 : 3'b100;
											assign node274 = (inp[10]) ? 3'b100 : 3'b101;
						assign node278 = (inp[0]) ? node298 : node279;
							assign node279 = (inp[9]) ? node289 : node280;
								assign node280 = (inp[11]) ? node282 : 3'b001;
									assign node282 = (inp[5]) ? node284 : 3'b001;
										assign node284 = (inp[10]) ? node286 : 3'b001;
											assign node286 = (inp[8]) ? 3'b000 : 3'b001;
								assign node289 = (inp[5]) ? node291 : 3'b010;
									assign node291 = (inp[11]) ? node293 : 3'b010;
										assign node293 = (inp[8]) ? node295 : 3'b010;
											assign node295 = (inp[10]) ? 3'b100 : 3'b010;
							assign node298 = (inp[9]) ? node314 : node299;
								assign node299 = (inp[11]) ? node307 : node300;
									assign node300 = (inp[8]) ? node304 : node301;
										assign node301 = (inp[10]) ? 3'b100 : 3'b010;
										assign node304 = (inp[10]) ? 3'b010 : 3'b110;
									assign node307 = (inp[10]) ? 3'b100 : node308;
										assign node308 = (inp[2]) ? node310 : 3'b100;
											assign node310 = (inp[8]) ? 3'b010 : 3'b100;
								assign node314 = (inp[2]) ? node316 : 3'b000;
									assign node316 = (inp[10]) ? 3'b000 : node317;
										assign node317 = (inp[8]) ? node319 : 3'b000;
											assign node319 = (inp[11]) ? 3'b000 : 3'b100;

endmodule