module dtc_split5_bm24 (
	input  wire [13-1:0] inp,
	output wire [13-1:0] outp
);

	wire [13-1:0] node1;
	wire [13-1:0] node2;
	wire [13-1:0] node3;
	wire [13-1:0] node4;
	wire [13-1:0] node5;
	wire [13-1:0] node6;
	wire [13-1:0] node7;
	wire [13-1:0] node8;
	wire [13-1:0] node9;
	wire [13-1:0] node10;
	wire [13-1:0] node13;
	wire [13-1:0] node16;
	wire [13-1:0] node17;
	wire [13-1:0] node20;
	wire [13-1:0] node23;
	wire [13-1:0] node24;
	wire [13-1:0] node26;
	wire [13-1:0] node29;
	wire [13-1:0] node30;
	wire [13-1:0] node33;
	wire [13-1:0] node36;
	wire [13-1:0] node37;
	wire [13-1:0] node38;
	wire [13-1:0] node40;
	wire [13-1:0] node43;
	wire [13-1:0] node44;
	wire [13-1:0] node47;
	wire [13-1:0] node50;
	wire [13-1:0] node51;
	wire [13-1:0] node53;
	wire [13-1:0] node56;
	wire [13-1:0] node57;
	wire [13-1:0] node61;
	wire [13-1:0] node62;
	wire [13-1:0] node63;
	wire [13-1:0] node64;
	wire [13-1:0] node65;
	wire [13-1:0] node68;
	wire [13-1:0] node71;
	wire [13-1:0] node72;
	wire [13-1:0] node75;
	wire [13-1:0] node78;
	wire [13-1:0] node79;
	wire [13-1:0] node80;
	wire [13-1:0] node83;
	wire [13-1:0] node86;
	wire [13-1:0] node87;
	wire [13-1:0] node90;
	wire [13-1:0] node93;
	wire [13-1:0] node94;
	wire [13-1:0] node95;
	wire [13-1:0] node96;
	wire [13-1:0] node99;
	wire [13-1:0] node102;
	wire [13-1:0] node103;
	wire [13-1:0] node106;
	wire [13-1:0] node109;
	wire [13-1:0] node110;
	wire [13-1:0] node111;
	wire [13-1:0] node115;
	wire [13-1:0] node116;
	wire [13-1:0] node119;
	wire [13-1:0] node122;
	wire [13-1:0] node123;
	wire [13-1:0] node124;
	wire [13-1:0] node125;
	wire [13-1:0] node126;
	wire [13-1:0] node127;
	wire [13-1:0] node130;
	wire [13-1:0] node133;
	wire [13-1:0] node134;
	wire [13-1:0] node137;
	wire [13-1:0] node140;
	wire [13-1:0] node141;
	wire [13-1:0] node142;
	wire [13-1:0] node145;
	wire [13-1:0] node148;
	wire [13-1:0] node149;
	wire [13-1:0] node152;
	wire [13-1:0] node155;
	wire [13-1:0] node156;
	wire [13-1:0] node157;
	wire [13-1:0] node158;
	wire [13-1:0] node161;
	wire [13-1:0] node164;
	wire [13-1:0] node165;
	wire [13-1:0] node168;
	wire [13-1:0] node171;
	wire [13-1:0] node172;
	wire [13-1:0] node173;
	wire [13-1:0] node176;
	wire [13-1:0] node179;
	wire [13-1:0] node180;
	wire [13-1:0] node184;
	wire [13-1:0] node185;
	wire [13-1:0] node186;
	wire [13-1:0] node187;
	wire [13-1:0] node188;
	wire [13-1:0] node191;
	wire [13-1:0] node194;
	wire [13-1:0] node195;
	wire [13-1:0] node198;
	wire [13-1:0] node201;
	wire [13-1:0] node202;
	wire [13-1:0] node203;
	wire [13-1:0] node206;
	wire [13-1:0] node209;
	wire [13-1:0] node210;
	wire [13-1:0] node213;
	wire [13-1:0] node216;
	wire [13-1:0] node217;
	wire [13-1:0] node218;
	wire [13-1:0] node219;
	wire [13-1:0] node222;
	wire [13-1:0] node225;
	wire [13-1:0] node227;
	wire [13-1:0] node230;
	wire [13-1:0] node231;
	wire [13-1:0] node232;
	wire [13-1:0] node235;
	wire [13-1:0] node238;
	wire [13-1:0] node239;
	wire [13-1:0] node242;
	wire [13-1:0] node245;
	wire [13-1:0] node246;
	wire [13-1:0] node247;
	wire [13-1:0] node248;
	wire [13-1:0] node249;
	wire [13-1:0] node250;
	wire [13-1:0] node252;
	wire [13-1:0] node255;
	wire [13-1:0] node256;
	wire [13-1:0] node259;
	wire [13-1:0] node262;
	wire [13-1:0] node263;
	wire [13-1:0] node264;
	wire [13-1:0] node267;
	wire [13-1:0] node270;
	wire [13-1:0] node271;
	wire [13-1:0] node275;
	wire [13-1:0] node276;
	wire [13-1:0] node277;
	wire [13-1:0] node278;
	wire [13-1:0] node281;
	wire [13-1:0] node284;
	wire [13-1:0] node285;
	wire [13-1:0] node288;
	wire [13-1:0] node291;
	wire [13-1:0] node292;
	wire [13-1:0] node294;
	wire [13-1:0] node297;
	wire [13-1:0] node298;
	wire [13-1:0] node301;
	wire [13-1:0] node304;
	wire [13-1:0] node305;
	wire [13-1:0] node306;
	wire [13-1:0] node307;
	wire [13-1:0] node308;
	wire [13-1:0] node311;
	wire [13-1:0] node314;
	wire [13-1:0] node315;
	wire [13-1:0] node318;
	wire [13-1:0] node321;
	wire [13-1:0] node322;
	wire [13-1:0] node323;
	wire [13-1:0] node326;
	wire [13-1:0] node329;
	wire [13-1:0] node330;
	wire [13-1:0] node333;
	wire [13-1:0] node336;
	wire [13-1:0] node337;
	wire [13-1:0] node338;
	wire [13-1:0] node340;
	wire [13-1:0] node343;
	wire [13-1:0] node344;
	wire [13-1:0] node347;
	wire [13-1:0] node350;
	wire [13-1:0] node351;
	wire [13-1:0] node352;
	wire [13-1:0] node355;
	wire [13-1:0] node358;
	wire [13-1:0] node359;
	wire [13-1:0] node362;
	wire [13-1:0] node365;
	wire [13-1:0] node366;
	wire [13-1:0] node367;
	wire [13-1:0] node368;
	wire [13-1:0] node369;
	wire [13-1:0] node370;
	wire [13-1:0] node373;
	wire [13-1:0] node376;
	wire [13-1:0] node378;
	wire [13-1:0] node381;
	wire [13-1:0] node382;
	wire [13-1:0] node383;
	wire [13-1:0] node386;
	wire [13-1:0] node389;
	wire [13-1:0] node390;
	wire [13-1:0] node393;
	wire [13-1:0] node396;
	wire [13-1:0] node397;
	wire [13-1:0] node398;
	wire [13-1:0] node399;
	wire [13-1:0] node402;
	wire [13-1:0] node405;
	wire [13-1:0] node406;
	wire [13-1:0] node409;
	wire [13-1:0] node412;
	wire [13-1:0] node413;
	wire [13-1:0] node414;
	wire [13-1:0] node417;
	wire [13-1:0] node420;
	wire [13-1:0] node421;
	wire [13-1:0] node424;
	wire [13-1:0] node427;
	wire [13-1:0] node428;
	wire [13-1:0] node429;
	wire [13-1:0] node430;
	wire [13-1:0] node431;
	wire [13-1:0] node434;
	wire [13-1:0] node437;
	wire [13-1:0] node438;
	wire [13-1:0] node441;
	wire [13-1:0] node444;
	wire [13-1:0] node445;
	wire [13-1:0] node446;
	wire [13-1:0] node449;
	wire [13-1:0] node452;
	wire [13-1:0] node453;
	wire [13-1:0] node456;
	wire [13-1:0] node459;
	wire [13-1:0] node460;
	wire [13-1:0] node461;
	wire [13-1:0] node463;
	wire [13-1:0] node466;
	wire [13-1:0] node467;
	wire [13-1:0] node470;
	wire [13-1:0] node473;
	wire [13-1:0] node474;
	wire [13-1:0] node476;
	wire [13-1:0] node479;
	wire [13-1:0] node480;
	wire [13-1:0] node483;
	wire [13-1:0] node486;
	wire [13-1:0] node487;
	wire [13-1:0] node488;
	wire [13-1:0] node489;
	wire [13-1:0] node490;
	wire [13-1:0] node491;
	wire [13-1:0] node492;
	wire [13-1:0] node493;
	wire [13-1:0] node496;
	wire [13-1:0] node499;
	wire [13-1:0] node500;
	wire [13-1:0] node503;
	wire [13-1:0] node506;
	wire [13-1:0] node507;
	wire [13-1:0] node508;
	wire [13-1:0] node511;
	wire [13-1:0] node514;
	wire [13-1:0] node515;
	wire [13-1:0] node518;
	wire [13-1:0] node521;
	wire [13-1:0] node522;
	wire [13-1:0] node523;
	wire [13-1:0] node524;
	wire [13-1:0] node527;
	wire [13-1:0] node530;
	wire [13-1:0] node531;
	wire [13-1:0] node534;
	wire [13-1:0] node537;
	wire [13-1:0] node538;
	wire [13-1:0] node539;
	wire [13-1:0] node542;
	wire [13-1:0] node545;
	wire [13-1:0] node546;
	wire [13-1:0] node549;
	wire [13-1:0] node552;
	wire [13-1:0] node553;
	wire [13-1:0] node554;
	wire [13-1:0] node555;
	wire [13-1:0] node556;
	wire [13-1:0] node559;
	wire [13-1:0] node562;
	wire [13-1:0] node563;
	wire [13-1:0] node567;
	wire [13-1:0] node568;
	wire [13-1:0] node569;
	wire [13-1:0] node572;
	wire [13-1:0] node575;
	wire [13-1:0] node576;
	wire [13-1:0] node579;
	wire [13-1:0] node582;
	wire [13-1:0] node583;
	wire [13-1:0] node584;
	wire [13-1:0] node585;
	wire [13-1:0] node588;
	wire [13-1:0] node591;
	wire [13-1:0] node592;
	wire [13-1:0] node595;
	wire [13-1:0] node598;
	wire [13-1:0] node599;
	wire [13-1:0] node600;
	wire [13-1:0] node604;
	wire [13-1:0] node605;
	wire [13-1:0] node608;
	wire [13-1:0] node611;
	wire [13-1:0] node612;
	wire [13-1:0] node613;
	wire [13-1:0] node614;
	wire [13-1:0] node615;
	wire [13-1:0] node616;
	wire [13-1:0] node619;
	wire [13-1:0] node622;
	wire [13-1:0] node624;
	wire [13-1:0] node627;
	wire [13-1:0] node628;
	wire [13-1:0] node629;
	wire [13-1:0] node632;
	wire [13-1:0] node635;
	wire [13-1:0] node636;
	wire [13-1:0] node639;
	wire [13-1:0] node642;
	wire [13-1:0] node643;
	wire [13-1:0] node644;
	wire [13-1:0] node645;
	wire [13-1:0] node648;
	wire [13-1:0] node651;
	wire [13-1:0] node652;
	wire [13-1:0] node655;
	wire [13-1:0] node658;
	wire [13-1:0] node659;
	wire [13-1:0] node660;
	wire [13-1:0] node663;
	wire [13-1:0] node666;
	wire [13-1:0] node668;
	wire [13-1:0] node671;
	wire [13-1:0] node672;
	wire [13-1:0] node673;
	wire [13-1:0] node674;
	wire [13-1:0] node675;
	wire [13-1:0] node678;
	wire [13-1:0] node681;
	wire [13-1:0] node682;
	wire [13-1:0] node686;
	wire [13-1:0] node687;
	wire [13-1:0] node688;
	wire [13-1:0] node691;
	wire [13-1:0] node694;
	wire [13-1:0] node695;
	wire [13-1:0] node698;
	wire [13-1:0] node701;
	wire [13-1:0] node702;
	wire [13-1:0] node703;
	wire [13-1:0] node704;
	wire [13-1:0] node707;
	wire [13-1:0] node710;
	wire [13-1:0] node711;
	wire [13-1:0] node714;
	wire [13-1:0] node717;
	wire [13-1:0] node718;
	wire [13-1:0] node720;
	wire [13-1:0] node723;
	wire [13-1:0] node724;
	wire [13-1:0] node727;
	wire [13-1:0] node730;
	wire [13-1:0] node731;
	wire [13-1:0] node732;
	wire [13-1:0] node733;
	wire [13-1:0] node734;
	wire [13-1:0] node735;
	wire [13-1:0] node736;
	wire [13-1:0] node739;
	wire [13-1:0] node742;
	wire [13-1:0] node743;
	wire [13-1:0] node747;
	wire [13-1:0] node748;
	wire [13-1:0] node749;
	wire [13-1:0] node752;
	wire [13-1:0] node755;
	wire [13-1:0] node757;
	wire [13-1:0] node760;
	wire [13-1:0] node761;
	wire [13-1:0] node762;
	wire [13-1:0] node763;
	wire [13-1:0] node766;
	wire [13-1:0] node769;
	wire [13-1:0] node770;
	wire [13-1:0] node773;
	wire [13-1:0] node776;
	wire [13-1:0] node777;
	wire [13-1:0] node778;
	wire [13-1:0] node782;
	wire [13-1:0] node783;
	wire [13-1:0] node786;
	wire [13-1:0] node789;
	wire [13-1:0] node790;
	wire [13-1:0] node791;
	wire [13-1:0] node792;
	wire [13-1:0] node793;
	wire [13-1:0] node796;
	wire [13-1:0] node799;
	wire [13-1:0] node800;
	wire [13-1:0] node803;
	wire [13-1:0] node806;
	wire [13-1:0] node807;
	wire [13-1:0] node808;
	wire [13-1:0] node811;
	wire [13-1:0] node814;
	wire [13-1:0] node815;
	wire [13-1:0] node818;
	wire [13-1:0] node821;
	wire [13-1:0] node822;
	wire [13-1:0] node823;
	wire [13-1:0] node824;
	wire [13-1:0] node827;
	wire [13-1:0] node830;
	wire [13-1:0] node832;
	wire [13-1:0] node835;
	wire [13-1:0] node836;
	wire [13-1:0] node837;
	wire [13-1:0] node840;
	wire [13-1:0] node843;
	wire [13-1:0] node845;
	wire [13-1:0] node848;
	wire [13-1:0] node849;
	wire [13-1:0] node850;
	wire [13-1:0] node851;
	wire [13-1:0] node852;
	wire [13-1:0] node853;
	wire [13-1:0] node856;
	wire [13-1:0] node859;
	wire [13-1:0] node860;
	wire [13-1:0] node863;
	wire [13-1:0] node866;
	wire [13-1:0] node867;
	wire [13-1:0] node868;
	wire [13-1:0] node871;
	wire [13-1:0] node874;
	wire [13-1:0] node875;
	wire [13-1:0] node878;
	wire [13-1:0] node881;
	wire [13-1:0] node882;
	wire [13-1:0] node883;
	wire [13-1:0] node884;
	wire [13-1:0] node887;
	wire [13-1:0] node890;
	wire [13-1:0] node891;
	wire [13-1:0] node894;
	wire [13-1:0] node897;
	wire [13-1:0] node898;
	wire [13-1:0] node899;
	wire [13-1:0] node903;
	wire [13-1:0] node904;
	wire [13-1:0] node907;
	wire [13-1:0] node910;
	wire [13-1:0] node911;
	wire [13-1:0] node912;
	wire [13-1:0] node913;
	wire [13-1:0] node914;
	wire [13-1:0] node917;
	wire [13-1:0] node920;
	wire [13-1:0] node921;
	wire [13-1:0] node924;
	wire [13-1:0] node927;
	wire [13-1:0] node928;
	wire [13-1:0] node929;
	wire [13-1:0] node932;
	wire [13-1:0] node935;
	wire [13-1:0] node936;
	wire [13-1:0] node939;
	wire [13-1:0] node942;
	wire [13-1:0] node943;
	wire [13-1:0] node944;
	wire [13-1:0] node945;
	wire [13-1:0] node948;
	wire [13-1:0] node951;
	wire [13-1:0] node952;
	wire [13-1:0] node955;
	wire [13-1:0] node958;
	wire [13-1:0] node959;
	wire [13-1:0] node960;
	wire [13-1:0] node963;
	wire [13-1:0] node966;
	wire [13-1:0] node967;
	wire [13-1:0] node970;
	wire [13-1:0] node973;
	wire [13-1:0] node974;
	wire [13-1:0] node975;
	wire [13-1:0] node976;
	wire [13-1:0] node977;
	wire [13-1:0] node978;
	wire [13-1:0] node979;
	wire [13-1:0] node980;
	wire [13-1:0] node981;
	wire [13-1:0] node984;
	wire [13-1:0] node987;
	wire [13-1:0] node988;
	wire [13-1:0] node991;
	wire [13-1:0] node994;
	wire [13-1:0] node995;
	wire [13-1:0] node997;
	wire [13-1:0] node1000;
	wire [13-1:0] node1001;
	wire [13-1:0] node1004;
	wire [13-1:0] node1007;
	wire [13-1:0] node1008;
	wire [13-1:0] node1009;
	wire [13-1:0] node1010;
	wire [13-1:0] node1013;
	wire [13-1:0] node1016;
	wire [13-1:0] node1017;
	wire [13-1:0] node1020;
	wire [13-1:0] node1023;
	wire [13-1:0] node1024;
	wire [13-1:0] node1025;
	wire [13-1:0] node1028;
	wire [13-1:0] node1031;
	wire [13-1:0] node1032;
	wire [13-1:0] node1035;
	wire [13-1:0] node1038;
	wire [13-1:0] node1039;
	wire [13-1:0] node1040;
	wire [13-1:0] node1041;
	wire [13-1:0] node1042;
	wire [13-1:0] node1045;
	wire [13-1:0] node1048;
	wire [13-1:0] node1049;
	wire [13-1:0] node1052;
	wire [13-1:0] node1055;
	wire [13-1:0] node1056;
	wire [13-1:0] node1057;
	wire [13-1:0] node1060;
	wire [13-1:0] node1063;
	wire [13-1:0] node1064;
	wire [13-1:0] node1067;
	wire [13-1:0] node1070;
	wire [13-1:0] node1071;
	wire [13-1:0] node1072;
	wire [13-1:0] node1074;
	wire [13-1:0] node1077;
	wire [13-1:0] node1078;
	wire [13-1:0] node1082;
	wire [13-1:0] node1083;
	wire [13-1:0] node1084;
	wire [13-1:0] node1087;
	wire [13-1:0] node1090;
	wire [13-1:0] node1091;
	wire [13-1:0] node1094;
	wire [13-1:0] node1097;
	wire [13-1:0] node1098;
	wire [13-1:0] node1099;
	wire [13-1:0] node1100;
	wire [13-1:0] node1101;
	wire [13-1:0] node1102;
	wire [13-1:0] node1105;
	wire [13-1:0] node1108;
	wire [13-1:0] node1109;
	wire [13-1:0] node1112;
	wire [13-1:0] node1115;
	wire [13-1:0] node1116;
	wire [13-1:0] node1117;
	wire [13-1:0] node1120;
	wire [13-1:0] node1123;
	wire [13-1:0] node1124;
	wire [13-1:0] node1127;
	wire [13-1:0] node1130;
	wire [13-1:0] node1131;
	wire [13-1:0] node1132;
	wire [13-1:0] node1133;
	wire [13-1:0] node1136;
	wire [13-1:0] node1140;
	wire [13-1:0] node1141;
	wire [13-1:0] node1142;
	wire [13-1:0] node1145;
	wire [13-1:0] node1148;
	wire [13-1:0] node1149;
	wire [13-1:0] node1152;
	wire [13-1:0] node1155;
	wire [13-1:0] node1156;
	wire [13-1:0] node1157;
	wire [13-1:0] node1158;
	wire [13-1:0] node1159;
	wire [13-1:0] node1162;
	wire [13-1:0] node1165;
	wire [13-1:0] node1167;
	wire [13-1:0] node1170;
	wire [13-1:0] node1171;
	wire [13-1:0] node1172;
	wire [13-1:0] node1175;
	wire [13-1:0] node1178;
	wire [13-1:0] node1179;
	wire [13-1:0] node1182;
	wire [13-1:0] node1185;
	wire [13-1:0] node1186;
	wire [13-1:0] node1187;
	wire [13-1:0] node1188;
	wire [13-1:0] node1191;
	wire [13-1:0] node1194;
	wire [13-1:0] node1195;
	wire [13-1:0] node1199;
	wire [13-1:0] node1200;
	wire [13-1:0] node1201;
	wire [13-1:0] node1204;
	wire [13-1:0] node1207;
	wire [13-1:0] node1208;
	wire [13-1:0] node1211;
	wire [13-1:0] node1214;
	wire [13-1:0] node1215;
	wire [13-1:0] node1216;
	wire [13-1:0] node1217;
	wire [13-1:0] node1218;
	wire [13-1:0] node1219;
	wire [13-1:0] node1220;
	wire [13-1:0] node1224;
	wire [13-1:0] node1225;
	wire [13-1:0] node1228;
	wire [13-1:0] node1231;
	wire [13-1:0] node1232;
	wire [13-1:0] node1233;
	wire [13-1:0] node1236;
	wire [13-1:0] node1239;
	wire [13-1:0] node1240;
	wire [13-1:0] node1243;
	wire [13-1:0] node1246;
	wire [13-1:0] node1247;
	wire [13-1:0] node1248;
	wire [13-1:0] node1250;
	wire [13-1:0] node1253;
	wire [13-1:0] node1254;
	wire [13-1:0] node1257;
	wire [13-1:0] node1260;
	wire [13-1:0] node1261;
	wire [13-1:0] node1263;
	wire [13-1:0] node1266;
	wire [13-1:0] node1268;
	wire [13-1:0] node1271;
	wire [13-1:0] node1272;
	wire [13-1:0] node1273;
	wire [13-1:0] node1274;
	wire [13-1:0] node1275;
	wire [13-1:0] node1278;
	wire [13-1:0] node1281;
	wire [13-1:0] node1282;
	wire [13-1:0] node1285;
	wire [13-1:0] node1288;
	wire [13-1:0] node1289;
	wire [13-1:0] node1290;
	wire [13-1:0] node1293;
	wire [13-1:0] node1296;
	wire [13-1:0] node1297;
	wire [13-1:0] node1300;
	wire [13-1:0] node1303;
	wire [13-1:0] node1304;
	wire [13-1:0] node1305;
	wire [13-1:0] node1306;
	wire [13-1:0] node1309;
	wire [13-1:0] node1312;
	wire [13-1:0] node1313;
	wire [13-1:0] node1316;
	wire [13-1:0] node1319;
	wire [13-1:0] node1320;
	wire [13-1:0] node1321;
	wire [13-1:0] node1324;
	wire [13-1:0] node1327;
	wire [13-1:0] node1328;
	wire [13-1:0] node1331;
	wire [13-1:0] node1334;
	wire [13-1:0] node1335;
	wire [13-1:0] node1336;
	wire [13-1:0] node1337;
	wire [13-1:0] node1338;
	wire [13-1:0] node1339;
	wire [13-1:0] node1342;
	wire [13-1:0] node1345;
	wire [13-1:0] node1346;
	wire [13-1:0] node1349;
	wire [13-1:0] node1352;
	wire [13-1:0] node1353;
	wire [13-1:0] node1354;
	wire [13-1:0] node1357;
	wire [13-1:0] node1360;
	wire [13-1:0] node1361;
	wire [13-1:0] node1364;
	wire [13-1:0] node1367;
	wire [13-1:0] node1368;
	wire [13-1:0] node1369;
	wire [13-1:0] node1370;
	wire [13-1:0] node1373;
	wire [13-1:0] node1376;
	wire [13-1:0] node1377;
	wire [13-1:0] node1380;
	wire [13-1:0] node1383;
	wire [13-1:0] node1384;
	wire [13-1:0] node1385;
	wire [13-1:0] node1388;
	wire [13-1:0] node1391;
	wire [13-1:0] node1392;
	wire [13-1:0] node1395;
	wire [13-1:0] node1398;
	wire [13-1:0] node1399;
	wire [13-1:0] node1400;
	wire [13-1:0] node1401;
	wire [13-1:0] node1402;
	wire [13-1:0] node1405;
	wire [13-1:0] node1408;
	wire [13-1:0] node1409;
	wire [13-1:0] node1412;
	wire [13-1:0] node1415;
	wire [13-1:0] node1416;
	wire [13-1:0] node1417;
	wire [13-1:0] node1420;
	wire [13-1:0] node1423;
	wire [13-1:0] node1424;
	wire [13-1:0] node1427;
	wire [13-1:0] node1430;
	wire [13-1:0] node1431;
	wire [13-1:0] node1432;
	wire [13-1:0] node1433;
	wire [13-1:0] node1436;
	wire [13-1:0] node1439;
	wire [13-1:0] node1440;
	wire [13-1:0] node1443;
	wire [13-1:0] node1446;
	wire [13-1:0] node1447;
	wire [13-1:0] node1448;
	wire [13-1:0] node1451;
	wire [13-1:0] node1454;
	wire [13-1:0] node1455;
	wire [13-1:0] node1458;
	wire [13-1:0] node1461;
	wire [13-1:0] node1462;
	wire [13-1:0] node1463;
	wire [13-1:0] node1464;
	wire [13-1:0] node1465;
	wire [13-1:0] node1466;
	wire [13-1:0] node1467;
	wire [13-1:0] node1468;
	wire [13-1:0] node1472;
	wire [13-1:0] node1473;
	wire [13-1:0] node1476;
	wire [13-1:0] node1479;
	wire [13-1:0] node1480;
	wire [13-1:0] node1481;
	wire [13-1:0] node1484;
	wire [13-1:0] node1487;
	wire [13-1:0] node1488;
	wire [13-1:0] node1491;
	wire [13-1:0] node1494;
	wire [13-1:0] node1495;
	wire [13-1:0] node1496;
	wire [13-1:0] node1497;
	wire [13-1:0] node1500;
	wire [13-1:0] node1503;
	wire [13-1:0] node1504;
	wire [13-1:0] node1508;
	wire [13-1:0] node1509;
	wire [13-1:0] node1510;
	wire [13-1:0] node1514;
	wire [13-1:0] node1515;
	wire [13-1:0] node1518;
	wire [13-1:0] node1521;
	wire [13-1:0] node1522;
	wire [13-1:0] node1523;
	wire [13-1:0] node1524;
	wire [13-1:0] node1525;
	wire [13-1:0] node1528;
	wire [13-1:0] node1531;
	wire [13-1:0] node1532;
	wire [13-1:0] node1535;
	wire [13-1:0] node1538;
	wire [13-1:0] node1539;
	wire [13-1:0] node1540;
	wire [13-1:0] node1543;
	wire [13-1:0] node1546;
	wire [13-1:0] node1547;
	wire [13-1:0] node1550;
	wire [13-1:0] node1553;
	wire [13-1:0] node1554;
	wire [13-1:0] node1555;
	wire [13-1:0] node1556;
	wire [13-1:0] node1559;
	wire [13-1:0] node1562;
	wire [13-1:0] node1563;
	wire [13-1:0] node1566;
	wire [13-1:0] node1569;
	wire [13-1:0] node1570;
	wire [13-1:0] node1571;
	wire [13-1:0] node1574;
	wire [13-1:0] node1577;
	wire [13-1:0] node1578;
	wire [13-1:0] node1581;
	wire [13-1:0] node1584;
	wire [13-1:0] node1585;
	wire [13-1:0] node1586;
	wire [13-1:0] node1587;
	wire [13-1:0] node1588;
	wire [13-1:0] node1589;
	wire [13-1:0] node1592;
	wire [13-1:0] node1595;
	wire [13-1:0] node1596;
	wire [13-1:0] node1599;
	wire [13-1:0] node1602;
	wire [13-1:0] node1603;
	wire [13-1:0] node1604;
	wire [13-1:0] node1607;
	wire [13-1:0] node1610;
	wire [13-1:0] node1611;
	wire [13-1:0] node1614;
	wire [13-1:0] node1617;
	wire [13-1:0] node1618;
	wire [13-1:0] node1619;
	wire [13-1:0] node1620;
	wire [13-1:0] node1623;
	wire [13-1:0] node1626;
	wire [13-1:0] node1627;
	wire [13-1:0] node1630;
	wire [13-1:0] node1633;
	wire [13-1:0] node1634;
	wire [13-1:0] node1635;
	wire [13-1:0] node1638;
	wire [13-1:0] node1641;
	wire [13-1:0] node1642;
	wire [13-1:0] node1645;
	wire [13-1:0] node1648;
	wire [13-1:0] node1649;
	wire [13-1:0] node1650;
	wire [13-1:0] node1651;
	wire [13-1:0] node1653;
	wire [13-1:0] node1656;
	wire [13-1:0] node1657;
	wire [13-1:0] node1660;
	wire [13-1:0] node1663;
	wire [13-1:0] node1664;
	wire [13-1:0] node1665;
	wire [13-1:0] node1668;
	wire [13-1:0] node1671;
	wire [13-1:0] node1672;
	wire [13-1:0] node1675;
	wire [13-1:0] node1678;
	wire [13-1:0] node1679;
	wire [13-1:0] node1680;
	wire [13-1:0] node1681;
	wire [13-1:0] node1684;
	wire [13-1:0] node1687;
	wire [13-1:0] node1688;
	wire [13-1:0] node1691;
	wire [13-1:0] node1694;
	wire [13-1:0] node1695;
	wire [13-1:0] node1696;
	wire [13-1:0] node1699;
	wire [13-1:0] node1702;
	wire [13-1:0] node1703;
	wire [13-1:0] node1706;
	wire [13-1:0] node1709;
	wire [13-1:0] node1710;
	wire [13-1:0] node1711;
	wire [13-1:0] node1712;
	wire [13-1:0] node1713;
	wire [13-1:0] node1714;
	wire [13-1:0] node1715;
	wire [13-1:0] node1718;
	wire [13-1:0] node1721;
	wire [13-1:0] node1722;
	wire [13-1:0] node1726;
	wire [13-1:0] node1727;
	wire [13-1:0] node1728;
	wire [13-1:0] node1731;
	wire [13-1:0] node1734;
	wire [13-1:0] node1735;
	wire [13-1:0] node1738;
	wire [13-1:0] node1741;
	wire [13-1:0] node1742;
	wire [13-1:0] node1743;
	wire [13-1:0] node1744;
	wire [13-1:0] node1747;
	wire [13-1:0] node1750;
	wire [13-1:0] node1751;
	wire [13-1:0] node1754;
	wire [13-1:0] node1757;
	wire [13-1:0] node1758;
	wire [13-1:0] node1760;
	wire [13-1:0] node1763;
	wire [13-1:0] node1764;
	wire [13-1:0] node1767;
	wire [13-1:0] node1770;
	wire [13-1:0] node1771;
	wire [13-1:0] node1772;
	wire [13-1:0] node1773;
	wire [13-1:0] node1775;
	wire [13-1:0] node1778;
	wire [13-1:0] node1779;
	wire [13-1:0] node1782;
	wire [13-1:0] node1785;
	wire [13-1:0] node1786;
	wire [13-1:0] node1787;
	wire [13-1:0] node1790;
	wire [13-1:0] node1793;
	wire [13-1:0] node1794;
	wire [13-1:0] node1797;
	wire [13-1:0] node1800;
	wire [13-1:0] node1801;
	wire [13-1:0] node1802;
	wire [13-1:0] node1803;
	wire [13-1:0] node1806;
	wire [13-1:0] node1809;
	wire [13-1:0] node1810;
	wire [13-1:0] node1813;
	wire [13-1:0] node1816;
	wire [13-1:0] node1817;
	wire [13-1:0] node1818;
	wire [13-1:0] node1821;
	wire [13-1:0] node1824;
	wire [13-1:0] node1825;
	wire [13-1:0] node1828;
	wire [13-1:0] node1831;
	wire [13-1:0] node1832;
	wire [13-1:0] node1833;
	wire [13-1:0] node1834;
	wire [13-1:0] node1835;
	wire [13-1:0] node1838;
	wire [13-1:0] node1839;
	wire [13-1:0] node1842;
	wire [13-1:0] node1845;
	wire [13-1:0] node1846;
	wire [13-1:0] node1847;
	wire [13-1:0] node1850;
	wire [13-1:0] node1853;
	wire [13-1:0] node1854;
	wire [13-1:0] node1857;
	wire [13-1:0] node1860;
	wire [13-1:0] node1861;
	wire [13-1:0] node1862;
	wire [13-1:0] node1863;
	wire [13-1:0] node1866;
	wire [13-1:0] node1869;
	wire [13-1:0] node1870;
	wire [13-1:0] node1873;
	wire [13-1:0] node1876;
	wire [13-1:0] node1877;
	wire [13-1:0] node1878;
	wire [13-1:0] node1881;
	wire [13-1:0] node1884;
	wire [13-1:0] node1885;
	wire [13-1:0] node1888;
	wire [13-1:0] node1891;
	wire [13-1:0] node1892;
	wire [13-1:0] node1893;
	wire [13-1:0] node1894;
	wire [13-1:0] node1895;
	wire [13-1:0] node1898;
	wire [13-1:0] node1901;
	wire [13-1:0] node1902;
	wire [13-1:0] node1905;
	wire [13-1:0] node1908;
	wire [13-1:0] node1909;
	wire [13-1:0] node1910;
	wire [13-1:0] node1913;
	wire [13-1:0] node1916;
	wire [13-1:0] node1917;
	wire [13-1:0] node1920;
	wire [13-1:0] node1923;
	wire [13-1:0] node1924;
	wire [13-1:0] node1925;
	wire [13-1:0] node1926;
	wire [13-1:0] node1929;
	wire [13-1:0] node1932;
	wire [13-1:0] node1934;
	wire [13-1:0] node1937;
	wire [13-1:0] node1938;
	wire [13-1:0] node1939;
	wire [13-1:0] node1942;
	wire [13-1:0] node1945;
	wire [13-1:0] node1946;
	wire [13-1:0] node1949;
	wire [13-1:0] node1952;
	wire [13-1:0] node1953;
	wire [13-1:0] node1954;
	wire [13-1:0] node1955;
	wire [13-1:0] node1956;
	wire [13-1:0] node1957;
	wire [13-1:0] node1958;
	wire [13-1:0] node1959;
	wire [13-1:0] node1960;
	wire [13-1:0] node1961;
	wire [13-1:0] node1964;
	wire [13-1:0] node1967;
	wire [13-1:0] node1968;
	wire [13-1:0] node1971;
	wire [13-1:0] node1974;
	wire [13-1:0] node1975;
	wire [13-1:0] node1976;
	wire [13-1:0] node1979;
	wire [13-1:0] node1982;
	wire [13-1:0] node1983;
	wire [13-1:0] node1986;
	wire [13-1:0] node1989;
	wire [13-1:0] node1990;
	wire [13-1:0] node1991;
	wire [13-1:0] node1993;
	wire [13-1:0] node1996;
	wire [13-1:0] node1997;
	wire [13-1:0] node2000;
	wire [13-1:0] node2003;
	wire [13-1:0] node2004;
	wire [13-1:0] node2005;
	wire [13-1:0] node2008;
	wire [13-1:0] node2011;
	wire [13-1:0] node2013;
	wire [13-1:0] node2016;
	wire [13-1:0] node2017;
	wire [13-1:0] node2018;
	wire [13-1:0] node2019;
	wire [13-1:0] node2020;
	wire [13-1:0] node2023;
	wire [13-1:0] node2026;
	wire [13-1:0] node2027;
	wire [13-1:0] node2030;
	wire [13-1:0] node2033;
	wire [13-1:0] node2034;
	wire [13-1:0] node2035;
	wire [13-1:0] node2038;
	wire [13-1:0] node2041;
	wire [13-1:0] node2042;
	wire [13-1:0] node2045;
	wire [13-1:0] node2048;
	wire [13-1:0] node2049;
	wire [13-1:0] node2050;
	wire [13-1:0] node2051;
	wire [13-1:0] node2054;
	wire [13-1:0] node2057;
	wire [13-1:0] node2058;
	wire [13-1:0] node2061;
	wire [13-1:0] node2064;
	wire [13-1:0] node2065;
	wire [13-1:0] node2067;
	wire [13-1:0] node2070;
	wire [13-1:0] node2072;
	wire [13-1:0] node2075;
	wire [13-1:0] node2076;
	wire [13-1:0] node2077;
	wire [13-1:0] node2078;
	wire [13-1:0] node2079;
	wire [13-1:0] node2080;
	wire [13-1:0] node2083;
	wire [13-1:0] node2086;
	wire [13-1:0] node2087;
	wire [13-1:0] node2090;
	wire [13-1:0] node2093;
	wire [13-1:0] node2094;
	wire [13-1:0] node2096;
	wire [13-1:0] node2099;
	wire [13-1:0] node2100;
	wire [13-1:0] node2103;
	wire [13-1:0] node2106;
	wire [13-1:0] node2107;
	wire [13-1:0] node2108;
	wire [13-1:0] node2109;
	wire [13-1:0] node2112;
	wire [13-1:0] node2115;
	wire [13-1:0] node2116;
	wire [13-1:0] node2119;
	wire [13-1:0] node2122;
	wire [13-1:0] node2123;
	wire [13-1:0] node2124;
	wire [13-1:0] node2127;
	wire [13-1:0] node2130;
	wire [13-1:0] node2131;
	wire [13-1:0] node2134;
	wire [13-1:0] node2137;
	wire [13-1:0] node2138;
	wire [13-1:0] node2139;
	wire [13-1:0] node2140;
	wire [13-1:0] node2141;
	wire [13-1:0] node2144;
	wire [13-1:0] node2147;
	wire [13-1:0] node2148;
	wire [13-1:0] node2151;
	wire [13-1:0] node2154;
	wire [13-1:0] node2155;
	wire [13-1:0] node2156;
	wire [13-1:0] node2159;
	wire [13-1:0] node2162;
	wire [13-1:0] node2163;
	wire [13-1:0] node2166;
	wire [13-1:0] node2169;
	wire [13-1:0] node2170;
	wire [13-1:0] node2171;
	wire [13-1:0] node2172;
	wire [13-1:0] node2175;
	wire [13-1:0] node2178;
	wire [13-1:0] node2179;
	wire [13-1:0] node2182;
	wire [13-1:0] node2185;
	wire [13-1:0] node2186;
	wire [13-1:0] node2187;
	wire [13-1:0] node2190;
	wire [13-1:0] node2193;
	wire [13-1:0] node2195;
	wire [13-1:0] node2198;
	wire [13-1:0] node2199;
	wire [13-1:0] node2200;
	wire [13-1:0] node2201;
	wire [13-1:0] node2202;
	wire [13-1:0] node2203;
	wire [13-1:0] node2204;
	wire [13-1:0] node2207;
	wire [13-1:0] node2210;
	wire [13-1:0] node2211;
	wire [13-1:0] node2214;
	wire [13-1:0] node2217;
	wire [13-1:0] node2218;
	wire [13-1:0] node2219;
	wire [13-1:0] node2222;
	wire [13-1:0] node2225;
	wire [13-1:0] node2226;
	wire [13-1:0] node2229;
	wire [13-1:0] node2232;
	wire [13-1:0] node2233;
	wire [13-1:0] node2234;
	wire [13-1:0] node2235;
	wire [13-1:0] node2239;
	wire [13-1:0] node2240;
	wire [13-1:0] node2244;
	wire [13-1:0] node2245;
	wire [13-1:0] node2246;
	wire [13-1:0] node2249;
	wire [13-1:0] node2252;
	wire [13-1:0] node2253;
	wire [13-1:0] node2256;
	wire [13-1:0] node2259;
	wire [13-1:0] node2260;
	wire [13-1:0] node2261;
	wire [13-1:0] node2262;
	wire [13-1:0] node2263;
	wire [13-1:0] node2266;
	wire [13-1:0] node2269;
	wire [13-1:0] node2270;
	wire [13-1:0] node2273;
	wire [13-1:0] node2276;
	wire [13-1:0] node2277;
	wire [13-1:0] node2278;
	wire [13-1:0] node2281;
	wire [13-1:0] node2284;
	wire [13-1:0] node2285;
	wire [13-1:0] node2288;
	wire [13-1:0] node2291;
	wire [13-1:0] node2292;
	wire [13-1:0] node2293;
	wire [13-1:0] node2295;
	wire [13-1:0] node2298;
	wire [13-1:0] node2299;
	wire [13-1:0] node2302;
	wire [13-1:0] node2305;
	wire [13-1:0] node2306;
	wire [13-1:0] node2307;
	wire [13-1:0] node2310;
	wire [13-1:0] node2313;
	wire [13-1:0] node2314;
	wire [13-1:0] node2317;
	wire [13-1:0] node2320;
	wire [13-1:0] node2321;
	wire [13-1:0] node2322;
	wire [13-1:0] node2323;
	wire [13-1:0] node2324;
	wire [13-1:0] node2325;
	wire [13-1:0] node2328;
	wire [13-1:0] node2331;
	wire [13-1:0] node2332;
	wire [13-1:0] node2335;
	wire [13-1:0] node2338;
	wire [13-1:0] node2339;
	wire [13-1:0] node2340;
	wire [13-1:0] node2343;
	wire [13-1:0] node2346;
	wire [13-1:0] node2347;
	wire [13-1:0] node2350;
	wire [13-1:0] node2353;
	wire [13-1:0] node2354;
	wire [13-1:0] node2355;
	wire [13-1:0] node2356;
	wire [13-1:0] node2359;
	wire [13-1:0] node2362;
	wire [13-1:0] node2363;
	wire [13-1:0] node2366;
	wire [13-1:0] node2369;
	wire [13-1:0] node2370;
	wire [13-1:0] node2371;
	wire [13-1:0] node2374;
	wire [13-1:0] node2377;
	wire [13-1:0] node2378;
	wire [13-1:0] node2382;
	wire [13-1:0] node2383;
	wire [13-1:0] node2384;
	wire [13-1:0] node2385;
	wire [13-1:0] node2386;
	wire [13-1:0] node2389;
	wire [13-1:0] node2392;
	wire [13-1:0] node2393;
	wire [13-1:0] node2396;
	wire [13-1:0] node2399;
	wire [13-1:0] node2400;
	wire [13-1:0] node2401;
	wire [13-1:0] node2404;
	wire [13-1:0] node2407;
	wire [13-1:0] node2408;
	wire [13-1:0] node2412;
	wire [13-1:0] node2413;
	wire [13-1:0] node2414;
	wire [13-1:0] node2415;
	wire [13-1:0] node2418;
	wire [13-1:0] node2421;
	wire [13-1:0] node2422;
	wire [13-1:0] node2425;
	wire [13-1:0] node2428;
	wire [13-1:0] node2429;
	wire [13-1:0] node2430;
	wire [13-1:0] node2433;
	wire [13-1:0] node2436;
	wire [13-1:0] node2438;
	wire [13-1:0] node2441;
	wire [13-1:0] node2442;
	wire [13-1:0] node2443;
	wire [13-1:0] node2444;
	wire [13-1:0] node2445;
	wire [13-1:0] node2446;
	wire [13-1:0] node2447;
	wire [13-1:0] node2448;
	wire [13-1:0] node2451;
	wire [13-1:0] node2454;
	wire [13-1:0] node2455;
	wire [13-1:0] node2459;
	wire [13-1:0] node2460;
	wire [13-1:0] node2461;
	wire [13-1:0] node2464;
	wire [13-1:0] node2467;
	wire [13-1:0] node2468;
	wire [13-1:0] node2472;
	wire [13-1:0] node2473;
	wire [13-1:0] node2474;
	wire [13-1:0] node2475;
	wire [13-1:0] node2479;
	wire [13-1:0] node2480;
	wire [13-1:0] node2483;
	wire [13-1:0] node2486;
	wire [13-1:0] node2487;
	wire [13-1:0] node2488;
	wire [13-1:0] node2491;
	wire [13-1:0] node2494;
	wire [13-1:0] node2495;
	wire [13-1:0] node2498;
	wire [13-1:0] node2501;
	wire [13-1:0] node2502;
	wire [13-1:0] node2503;
	wire [13-1:0] node2504;
	wire [13-1:0] node2505;
	wire [13-1:0] node2508;
	wire [13-1:0] node2511;
	wire [13-1:0] node2512;
	wire [13-1:0] node2515;
	wire [13-1:0] node2518;
	wire [13-1:0] node2519;
	wire [13-1:0] node2520;
	wire [13-1:0] node2523;
	wire [13-1:0] node2526;
	wire [13-1:0] node2527;
	wire [13-1:0] node2530;
	wire [13-1:0] node2533;
	wire [13-1:0] node2534;
	wire [13-1:0] node2535;
	wire [13-1:0] node2536;
	wire [13-1:0] node2539;
	wire [13-1:0] node2542;
	wire [13-1:0] node2543;
	wire [13-1:0] node2546;
	wire [13-1:0] node2549;
	wire [13-1:0] node2550;
	wire [13-1:0] node2551;
	wire [13-1:0] node2554;
	wire [13-1:0] node2557;
	wire [13-1:0] node2558;
	wire [13-1:0] node2561;
	wire [13-1:0] node2564;
	wire [13-1:0] node2565;
	wire [13-1:0] node2566;
	wire [13-1:0] node2567;
	wire [13-1:0] node2568;
	wire [13-1:0] node2569;
	wire [13-1:0] node2572;
	wire [13-1:0] node2575;
	wire [13-1:0] node2576;
	wire [13-1:0] node2579;
	wire [13-1:0] node2582;
	wire [13-1:0] node2583;
	wire [13-1:0] node2585;
	wire [13-1:0] node2588;
	wire [13-1:0] node2589;
	wire [13-1:0] node2593;
	wire [13-1:0] node2594;
	wire [13-1:0] node2595;
	wire [13-1:0] node2596;
	wire [13-1:0] node2599;
	wire [13-1:0] node2602;
	wire [13-1:0] node2604;
	wire [13-1:0] node2607;
	wire [13-1:0] node2608;
	wire [13-1:0] node2609;
	wire [13-1:0] node2612;
	wire [13-1:0] node2615;
	wire [13-1:0] node2616;
	wire [13-1:0] node2619;
	wire [13-1:0] node2622;
	wire [13-1:0] node2623;
	wire [13-1:0] node2624;
	wire [13-1:0] node2625;
	wire [13-1:0] node2627;
	wire [13-1:0] node2630;
	wire [13-1:0] node2631;
	wire [13-1:0] node2634;
	wire [13-1:0] node2637;
	wire [13-1:0] node2638;
	wire [13-1:0] node2639;
	wire [13-1:0] node2642;
	wire [13-1:0] node2645;
	wire [13-1:0] node2646;
	wire [13-1:0] node2649;
	wire [13-1:0] node2652;
	wire [13-1:0] node2653;
	wire [13-1:0] node2654;
	wire [13-1:0] node2655;
	wire [13-1:0] node2659;
	wire [13-1:0] node2660;
	wire [13-1:0] node2663;
	wire [13-1:0] node2666;
	wire [13-1:0] node2667;
	wire [13-1:0] node2668;
	wire [13-1:0] node2671;
	wire [13-1:0] node2674;
	wire [13-1:0] node2675;
	wire [13-1:0] node2678;
	wire [13-1:0] node2681;
	wire [13-1:0] node2682;
	wire [13-1:0] node2683;
	wire [13-1:0] node2684;
	wire [13-1:0] node2685;
	wire [13-1:0] node2686;
	wire [13-1:0] node2687;
	wire [13-1:0] node2690;
	wire [13-1:0] node2693;
	wire [13-1:0] node2694;
	wire [13-1:0] node2697;
	wire [13-1:0] node2700;
	wire [13-1:0] node2701;
	wire [13-1:0] node2702;
	wire [13-1:0] node2705;
	wire [13-1:0] node2708;
	wire [13-1:0] node2709;
	wire [13-1:0] node2712;
	wire [13-1:0] node2715;
	wire [13-1:0] node2716;
	wire [13-1:0] node2717;
	wire [13-1:0] node2718;
	wire [13-1:0] node2721;
	wire [13-1:0] node2724;
	wire [13-1:0] node2725;
	wire [13-1:0] node2728;
	wire [13-1:0] node2731;
	wire [13-1:0] node2732;
	wire [13-1:0] node2733;
	wire [13-1:0] node2736;
	wire [13-1:0] node2739;
	wire [13-1:0] node2740;
	wire [13-1:0] node2743;
	wire [13-1:0] node2746;
	wire [13-1:0] node2747;
	wire [13-1:0] node2748;
	wire [13-1:0] node2749;
	wire [13-1:0] node2751;
	wire [13-1:0] node2754;
	wire [13-1:0] node2755;
	wire [13-1:0] node2758;
	wire [13-1:0] node2761;
	wire [13-1:0] node2762;
	wire [13-1:0] node2764;
	wire [13-1:0] node2767;
	wire [13-1:0] node2768;
	wire [13-1:0] node2771;
	wire [13-1:0] node2774;
	wire [13-1:0] node2775;
	wire [13-1:0] node2776;
	wire [13-1:0] node2777;
	wire [13-1:0] node2781;
	wire [13-1:0] node2782;
	wire [13-1:0] node2785;
	wire [13-1:0] node2788;
	wire [13-1:0] node2789;
	wire [13-1:0] node2790;
	wire [13-1:0] node2793;
	wire [13-1:0] node2796;
	wire [13-1:0] node2797;
	wire [13-1:0] node2800;
	wire [13-1:0] node2803;
	wire [13-1:0] node2804;
	wire [13-1:0] node2805;
	wire [13-1:0] node2806;
	wire [13-1:0] node2807;
	wire [13-1:0] node2808;
	wire [13-1:0] node2811;
	wire [13-1:0] node2814;
	wire [13-1:0] node2815;
	wire [13-1:0] node2818;
	wire [13-1:0] node2821;
	wire [13-1:0] node2822;
	wire [13-1:0] node2823;
	wire [13-1:0] node2826;
	wire [13-1:0] node2829;
	wire [13-1:0] node2830;
	wire [13-1:0] node2833;
	wire [13-1:0] node2836;
	wire [13-1:0] node2837;
	wire [13-1:0] node2838;
	wire [13-1:0] node2839;
	wire [13-1:0] node2842;
	wire [13-1:0] node2845;
	wire [13-1:0] node2846;
	wire [13-1:0] node2849;
	wire [13-1:0] node2852;
	wire [13-1:0] node2853;
	wire [13-1:0] node2855;
	wire [13-1:0] node2858;
	wire [13-1:0] node2859;
	wire [13-1:0] node2862;
	wire [13-1:0] node2865;
	wire [13-1:0] node2866;
	wire [13-1:0] node2867;
	wire [13-1:0] node2868;
	wire [13-1:0] node2869;
	wire [13-1:0] node2872;
	wire [13-1:0] node2875;
	wire [13-1:0] node2876;
	wire [13-1:0] node2879;
	wire [13-1:0] node2882;
	wire [13-1:0] node2883;
	wire [13-1:0] node2885;
	wire [13-1:0] node2888;
	wire [13-1:0] node2889;
	wire [13-1:0] node2892;
	wire [13-1:0] node2895;
	wire [13-1:0] node2896;
	wire [13-1:0] node2897;
	wire [13-1:0] node2899;
	wire [13-1:0] node2902;
	wire [13-1:0] node2903;
	wire [13-1:0] node2906;
	wire [13-1:0] node2909;
	wire [13-1:0] node2910;
	wire [13-1:0] node2912;
	wire [13-1:0] node2915;
	wire [13-1:0] node2916;
	wire [13-1:0] node2919;
	wire [13-1:0] node2922;
	wire [13-1:0] node2923;
	wire [13-1:0] node2924;
	wire [13-1:0] node2925;
	wire [13-1:0] node2926;
	wire [13-1:0] node2927;
	wire [13-1:0] node2928;
	wire [13-1:0] node2929;
	wire [13-1:0] node2930;
	wire [13-1:0] node2933;
	wire [13-1:0] node2936;
	wire [13-1:0] node2937;
	wire [13-1:0] node2940;
	wire [13-1:0] node2943;
	wire [13-1:0] node2944;
	wire [13-1:0] node2945;
	wire [13-1:0] node2948;
	wire [13-1:0] node2951;
	wire [13-1:0] node2952;
	wire [13-1:0] node2956;
	wire [13-1:0] node2957;
	wire [13-1:0] node2958;
	wire [13-1:0] node2959;
	wire [13-1:0] node2962;
	wire [13-1:0] node2965;
	wire [13-1:0] node2966;
	wire [13-1:0] node2969;
	wire [13-1:0] node2972;
	wire [13-1:0] node2973;
	wire [13-1:0] node2974;
	wire [13-1:0] node2977;
	wire [13-1:0] node2980;
	wire [13-1:0] node2981;
	wire [13-1:0] node2984;
	wire [13-1:0] node2987;
	wire [13-1:0] node2988;
	wire [13-1:0] node2989;
	wire [13-1:0] node2990;
	wire [13-1:0] node2991;
	wire [13-1:0] node2995;
	wire [13-1:0] node2996;
	wire [13-1:0] node2999;
	wire [13-1:0] node3002;
	wire [13-1:0] node3003;
	wire [13-1:0] node3004;
	wire [13-1:0] node3007;
	wire [13-1:0] node3010;
	wire [13-1:0] node3011;
	wire [13-1:0] node3014;
	wire [13-1:0] node3017;
	wire [13-1:0] node3018;
	wire [13-1:0] node3019;
	wire [13-1:0] node3020;
	wire [13-1:0] node3023;
	wire [13-1:0] node3026;
	wire [13-1:0] node3027;
	wire [13-1:0] node3030;
	wire [13-1:0] node3033;
	wire [13-1:0] node3034;
	wire [13-1:0] node3035;
	wire [13-1:0] node3038;
	wire [13-1:0] node3041;
	wire [13-1:0] node3042;
	wire [13-1:0] node3045;
	wire [13-1:0] node3048;
	wire [13-1:0] node3049;
	wire [13-1:0] node3050;
	wire [13-1:0] node3051;
	wire [13-1:0] node3052;
	wire [13-1:0] node3053;
	wire [13-1:0] node3057;
	wire [13-1:0] node3058;
	wire [13-1:0] node3062;
	wire [13-1:0] node3063;
	wire [13-1:0] node3065;
	wire [13-1:0] node3068;
	wire [13-1:0] node3069;
	wire [13-1:0] node3072;
	wire [13-1:0] node3075;
	wire [13-1:0] node3076;
	wire [13-1:0] node3077;
	wire [13-1:0] node3078;
	wire [13-1:0] node3081;
	wire [13-1:0] node3084;
	wire [13-1:0] node3085;
	wire [13-1:0] node3088;
	wire [13-1:0] node3091;
	wire [13-1:0] node3092;
	wire [13-1:0] node3093;
	wire [13-1:0] node3096;
	wire [13-1:0] node3099;
	wire [13-1:0] node3100;
	wire [13-1:0] node3103;
	wire [13-1:0] node3106;
	wire [13-1:0] node3107;
	wire [13-1:0] node3108;
	wire [13-1:0] node3109;
	wire [13-1:0] node3111;
	wire [13-1:0] node3114;
	wire [13-1:0] node3115;
	wire [13-1:0] node3118;
	wire [13-1:0] node3121;
	wire [13-1:0] node3122;
	wire [13-1:0] node3123;
	wire [13-1:0] node3126;
	wire [13-1:0] node3129;
	wire [13-1:0] node3130;
	wire [13-1:0] node3133;
	wire [13-1:0] node3136;
	wire [13-1:0] node3137;
	wire [13-1:0] node3138;
	wire [13-1:0] node3139;
	wire [13-1:0] node3142;
	wire [13-1:0] node3145;
	wire [13-1:0] node3146;
	wire [13-1:0] node3149;
	wire [13-1:0] node3152;
	wire [13-1:0] node3153;
	wire [13-1:0] node3155;
	wire [13-1:0] node3158;
	wire [13-1:0] node3159;
	wire [13-1:0] node3162;
	wire [13-1:0] node3165;
	wire [13-1:0] node3166;
	wire [13-1:0] node3167;
	wire [13-1:0] node3168;
	wire [13-1:0] node3169;
	wire [13-1:0] node3170;
	wire [13-1:0] node3171;
	wire [13-1:0] node3175;
	wire [13-1:0] node3176;
	wire [13-1:0] node3179;
	wire [13-1:0] node3182;
	wire [13-1:0] node3183;
	wire [13-1:0] node3184;
	wire [13-1:0] node3187;
	wire [13-1:0] node3190;
	wire [13-1:0] node3191;
	wire [13-1:0] node3194;
	wire [13-1:0] node3197;
	wire [13-1:0] node3198;
	wire [13-1:0] node3199;
	wire [13-1:0] node3200;
	wire [13-1:0] node3204;
	wire [13-1:0] node3205;
	wire [13-1:0] node3208;
	wire [13-1:0] node3211;
	wire [13-1:0] node3212;
	wire [13-1:0] node3213;
	wire [13-1:0] node3216;
	wire [13-1:0] node3219;
	wire [13-1:0] node3220;
	wire [13-1:0] node3223;
	wire [13-1:0] node3226;
	wire [13-1:0] node3227;
	wire [13-1:0] node3228;
	wire [13-1:0] node3229;
	wire [13-1:0] node3230;
	wire [13-1:0] node3233;
	wire [13-1:0] node3236;
	wire [13-1:0] node3237;
	wire [13-1:0] node3240;
	wire [13-1:0] node3243;
	wire [13-1:0] node3244;
	wire [13-1:0] node3245;
	wire [13-1:0] node3248;
	wire [13-1:0] node3251;
	wire [13-1:0] node3252;
	wire [13-1:0] node3255;
	wire [13-1:0] node3258;
	wire [13-1:0] node3259;
	wire [13-1:0] node3260;
	wire [13-1:0] node3261;
	wire [13-1:0] node3264;
	wire [13-1:0] node3267;
	wire [13-1:0] node3268;
	wire [13-1:0] node3271;
	wire [13-1:0] node3274;
	wire [13-1:0] node3275;
	wire [13-1:0] node3276;
	wire [13-1:0] node3279;
	wire [13-1:0] node3282;
	wire [13-1:0] node3283;
	wire [13-1:0] node3286;
	wire [13-1:0] node3289;
	wire [13-1:0] node3290;
	wire [13-1:0] node3291;
	wire [13-1:0] node3292;
	wire [13-1:0] node3293;
	wire [13-1:0] node3294;
	wire [13-1:0] node3297;
	wire [13-1:0] node3301;
	wire [13-1:0] node3302;
	wire [13-1:0] node3303;
	wire [13-1:0] node3306;
	wire [13-1:0] node3309;
	wire [13-1:0] node3310;
	wire [13-1:0] node3313;
	wire [13-1:0] node3316;
	wire [13-1:0] node3317;
	wire [13-1:0] node3318;
	wire [13-1:0] node3319;
	wire [13-1:0] node3322;
	wire [13-1:0] node3325;
	wire [13-1:0] node3326;
	wire [13-1:0] node3329;
	wire [13-1:0] node3332;
	wire [13-1:0] node3333;
	wire [13-1:0] node3334;
	wire [13-1:0] node3337;
	wire [13-1:0] node3340;
	wire [13-1:0] node3341;
	wire [13-1:0] node3344;
	wire [13-1:0] node3347;
	wire [13-1:0] node3348;
	wire [13-1:0] node3349;
	wire [13-1:0] node3350;
	wire [13-1:0] node3351;
	wire [13-1:0] node3354;
	wire [13-1:0] node3357;
	wire [13-1:0] node3358;
	wire [13-1:0] node3362;
	wire [13-1:0] node3363;
	wire [13-1:0] node3364;
	wire [13-1:0] node3367;
	wire [13-1:0] node3370;
	wire [13-1:0] node3371;
	wire [13-1:0] node3374;
	wire [13-1:0] node3377;
	wire [13-1:0] node3378;
	wire [13-1:0] node3379;
	wire [13-1:0] node3380;
	wire [13-1:0] node3383;
	wire [13-1:0] node3386;
	wire [13-1:0] node3387;
	wire [13-1:0] node3390;
	wire [13-1:0] node3393;
	wire [13-1:0] node3394;
	wire [13-1:0] node3395;
	wire [13-1:0] node3398;
	wire [13-1:0] node3401;
	wire [13-1:0] node3402;
	wire [13-1:0] node3405;
	wire [13-1:0] node3408;
	wire [13-1:0] node3409;
	wire [13-1:0] node3410;
	wire [13-1:0] node3411;
	wire [13-1:0] node3412;
	wire [13-1:0] node3413;
	wire [13-1:0] node3414;
	wire [13-1:0] node3415;
	wire [13-1:0] node3418;
	wire [13-1:0] node3421;
	wire [13-1:0] node3423;
	wire [13-1:0] node3426;
	wire [13-1:0] node3427;
	wire [13-1:0] node3428;
	wire [13-1:0] node3431;
	wire [13-1:0] node3434;
	wire [13-1:0] node3435;
	wire [13-1:0] node3438;
	wire [13-1:0] node3441;
	wire [13-1:0] node3442;
	wire [13-1:0] node3443;
	wire [13-1:0] node3444;
	wire [13-1:0] node3448;
	wire [13-1:0] node3449;
	wire [13-1:0] node3452;
	wire [13-1:0] node3455;
	wire [13-1:0] node3456;
	wire [13-1:0] node3457;
	wire [13-1:0] node3460;
	wire [13-1:0] node3463;
	wire [13-1:0] node3464;
	wire [13-1:0] node3467;
	wire [13-1:0] node3470;
	wire [13-1:0] node3471;
	wire [13-1:0] node3472;
	wire [13-1:0] node3473;
	wire [13-1:0] node3474;
	wire [13-1:0] node3477;
	wire [13-1:0] node3480;
	wire [13-1:0] node3481;
	wire [13-1:0] node3484;
	wire [13-1:0] node3487;
	wire [13-1:0] node3488;
	wire [13-1:0] node3489;
	wire [13-1:0] node3492;
	wire [13-1:0] node3495;
	wire [13-1:0] node3496;
	wire [13-1:0] node3499;
	wire [13-1:0] node3502;
	wire [13-1:0] node3503;
	wire [13-1:0] node3504;
	wire [13-1:0] node3506;
	wire [13-1:0] node3509;
	wire [13-1:0] node3510;
	wire [13-1:0] node3513;
	wire [13-1:0] node3516;
	wire [13-1:0] node3517;
	wire [13-1:0] node3518;
	wire [13-1:0] node3521;
	wire [13-1:0] node3524;
	wire [13-1:0] node3526;
	wire [13-1:0] node3529;
	wire [13-1:0] node3530;
	wire [13-1:0] node3531;
	wire [13-1:0] node3532;
	wire [13-1:0] node3533;
	wire [13-1:0] node3534;
	wire [13-1:0] node3537;
	wire [13-1:0] node3540;
	wire [13-1:0] node3542;
	wire [13-1:0] node3545;
	wire [13-1:0] node3546;
	wire [13-1:0] node3547;
	wire [13-1:0] node3550;
	wire [13-1:0] node3553;
	wire [13-1:0] node3554;
	wire [13-1:0] node3557;
	wire [13-1:0] node3560;
	wire [13-1:0] node3561;
	wire [13-1:0] node3562;
	wire [13-1:0] node3563;
	wire [13-1:0] node3566;
	wire [13-1:0] node3569;
	wire [13-1:0] node3570;
	wire [13-1:0] node3573;
	wire [13-1:0] node3576;
	wire [13-1:0] node3577;
	wire [13-1:0] node3578;
	wire [13-1:0] node3581;
	wire [13-1:0] node3584;
	wire [13-1:0] node3585;
	wire [13-1:0] node3588;
	wire [13-1:0] node3591;
	wire [13-1:0] node3592;
	wire [13-1:0] node3593;
	wire [13-1:0] node3594;
	wire [13-1:0] node3595;
	wire [13-1:0] node3598;
	wire [13-1:0] node3601;
	wire [13-1:0] node3602;
	wire [13-1:0] node3605;
	wire [13-1:0] node3608;
	wire [13-1:0] node3609;
	wire [13-1:0] node3610;
	wire [13-1:0] node3613;
	wire [13-1:0] node3616;
	wire [13-1:0] node3617;
	wire [13-1:0] node3620;
	wire [13-1:0] node3623;
	wire [13-1:0] node3624;
	wire [13-1:0] node3625;
	wire [13-1:0] node3626;
	wire [13-1:0] node3629;
	wire [13-1:0] node3632;
	wire [13-1:0] node3633;
	wire [13-1:0] node3636;
	wire [13-1:0] node3639;
	wire [13-1:0] node3640;
	wire [13-1:0] node3641;
	wire [13-1:0] node3644;
	wire [13-1:0] node3647;
	wire [13-1:0] node3648;
	wire [13-1:0] node3651;
	wire [13-1:0] node3654;
	wire [13-1:0] node3655;
	wire [13-1:0] node3656;
	wire [13-1:0] node3657;
	wire [13-1:0] node3658;
	wire [13-1:0] node3659;
	wire [13-1:0] node3660;
	wire [13-1:0] node3663;
	wire [13-1:0] node3666;
	wire [13-1:0] node3667;
	wire [13-1:0] node3671;
	wire [13-1:0] node3672;
	wire [13-1:0] node3673;
	wire [13-1:0] node3676;
	wire [13-1:0] node3679;
	wire [13-1:0] node3680;
	wire [13-1:0] node3683;
	wire [13-1:0] node3686;
	wire [13-1:0] node3687;
	wire [13-1:0] node3688;
	wire [13-1:0] node3689;
	wire [13-1:0] node3692;
	wire [13-1:0] node3695;
	wire [13-1:0] node3697;
	wire [13-1:0] node3700;
	wire [13-1:0] node3701;
	wire [13-1:0] node3703;
	wire [13-1:0] node3706;
	wire [13-1:0] node3707;
	wire [13-1:0] node3710;
	wire [13-1:0] node3713;
	wire [13-1:0] node3714;
	wire [13-1:0] node3715;
	wire [13-1:0] node3716;
	wire [13-1:0] node3717;
	wire [13-1:0] node3720;
	wire [13-1:0] node3723;
	wire [13-1:0] node3724;
	wire [13-1:0] node3727;
	wire [13-1:0] node3730;
	wire [13-1:0] node3731;
	wire [13-1:0] node3732;
	wire [13-1:0] node3735;
	wire [13-1:0] node3738;
	wire [13-1:0] node3739;
	wire [13-1:0] node3742;
	wire [13-1:0] node3745;
	wire [13-1:0] node3746;
	wire [13-1:0] node3747;
	wire [13-1:0] node3748;
	wire [13-1:0] node3751;
	wire [13-1:0] node3754;
	wire [13-1:0] node3755;
	wire [13-1:0] node3758;
	wire [13-1:0] node3761;
	wire [13-1:0] node3762;
	wire [13-1:0] node3763;
	wire [13-1:0] node3766;
	wire [13-1:0] node3769;
	wire [13-1:0] node3770;
	wire [13-1:0] node3773;
	wire [13-1:0] node3776;
	wire [13-1:0] node3777;
	wire [13-1:0] node3778;
	wire [13-1:0] node3779;
	wire [13-1:0] node3780;
	wire [13-1:0] node3781;
	wire [13-1:0] node3785;
	wire [13-1:0] node3786;
	wire [13-1:0] node3789;
	wire [13-1:0] node3792;
	wire [13-1:0] node3793;
	wire [13-1:0] node3794;
	wire [13-1:0] node3797;
	wire [13-1:0] node3800;
	wire [13-1:0] node3801;
	wire [13-1:0] node3804;
	wire [13-1:0] node3807;
	wire [13-1:0] node3808;
	wire [13-1:0] node3809;
	wire [13-1:0] node3810;
	wire [13-1:0] node3813;
	wire [13-1:0] node3817;
	wire [13-1:0] node3818;
	wire [13-1:0] node3819;
	wire [13-1:0] node3822;
	wire [13-1:0] node3825;
	wire [13-1:0] node3827;
	wire [13-1:0] node3830;
	wire [13-1:0] node3831;
	wire [13-1:0] node3832;
	wire [13-1:0] node3833;
	wire [13-1:0] node3834;
	wire [13-1:0] node3837;
	wire [13-1:0] node3840;
	wire [13-1:0] node3842;
	wire [13-1:0] node3845;
	wire [13-1:0] node3846;
	wire [13-1:0] node3847;
	wire [13-1:0] node3850;
	wire [13-1:0] node3853;
	wire [13-1:0] node3854;
	wire [13-1:0] node3857;
	wire [13-1:0] node3860;
	wire [13-1:0] node3861;
	wire [13-1:0] node3862;
	wire [13-1:0] node3863;
	wire [13-1:0] node3866;
	wire [13-1:0] node3869;
	wire [13-1:0] node3870;
	wire [13-1:0] node3873;
	wire [13-1:0] node3876;
	wire [13-1:0] node3877;
	wire [13-1:0] node3878;
	wire [13-1:0] node3881;
	wire [13-1:0] node3884;
	wire [13-1:0] node3885;
	wire [13-1:0] node3888;

	assign outp = (inp[12]) ? node1952 : node1;
		assign node1 = (inp[4]) ? node973 : node2;
			assign node2 = (inp[6]) ? node486 : node3;
				assign node3 = (inp[1]) ? node245 : node4;
					assign node4 = (inp[11]) ? node122 : node5;
						assign node5 = (inp[3]) ? node61 : node6;
							assign node6 = (inp[8]) ? node36 : node7;
								assign node7 = (inp[0]) ? node23 : node8;
									assign node8 = (inp[5]) ? node16 : node9;
										assign node9 = (inp[7]) ? node13 : node10;
											assign node10 = (inp[10]) ? 13'b0011111111111 : 13'b0111111111111;
											assign node13 = (inp[2]) ? 13'b0001111111111 : 13'b0011111111111;
										assign node16 = (inp[9]) ? node20 : node17;
											assign node17 = (inp[10]) ? 13'b0001111111111 : 13'b0011111111111;
											assign node20 = (inp[7]) ? 13'b0000011111111 : 13'b0001111111111;
									assign node23 = (inp[7]) ? node29 : node24;
										assign node24 = (inp[5]) ? node26 : 13'b0001111111111;
											assign node26 = (inp[9]) ? 13'b0001111111111 : 13'b0001111111111;
										assign node29 = (inp[9]) ? node33 : node30;
											assign node30 = (inp[5]) ? 13'b0000111111111 : 13'b0001111111111;
											assign node33 = (inp[2]) ? 13'b0000011111111 : 13'b0000111111111;
								assign node36 = (inp[10]) ? node50 : node37;
									assign node37 = (inp[0]) ? node43 : node38;
										assign node38 = (inp[5]) ? node40 : 13'b0011111111111;
											assign node40 = (inp[2]) ? 13'b0000111111111 : 13'b0001111111111;
										assign node43 = (inp[2]) ? node47 : node44;
											assign node44 = (inp[7]) ? 13'b0000111111111 : 13'b0001111111111;
											assign node47 = (inp[7]) ? 13'b0000111111111 : 13'b0000111111111;
									assign node50 = (inp[9]) ? node56 : node51;
										assign node51 = (inp[7]) ? node53 : 13'b0001111111111;
											assign node53 = (inp[5]) ? 13'b0000011111111 : 13'b0000111111111;
										assign node56 = (inp[7]) ? 13'b0000001111111 : node57;
											assign node57 = (inp[2]) ? 13'b0000011111111 : 13'b0000111111111;
							assign node61 = (inp[7]) ? node93 : node62;
								assign node62 = (inp[0]) ? node78 : node63;
									assign node63 = (inp[10]) ? node71 : node64;
										assign node64 = (inp[5]) ? node68 : node65;
											assign node65 = (inp[8]) ? 13'b0001111111111 : 13'b0011111111111;
											assign node68 = (inp[8]) ? 13'b0000111111111 : 13'b0001111111111;
										assign node71 = (inp[2]) ? node75 : node72;
											assign node72 = (inp[9]) ? 13'b0000111111111 : 13'b0001111111111;
											assign node75 = (inp[5]) ? 13'b0000011111111 : 13'b0000111111111;
									assign node78 = (inp[2]) ? node86 : node79;
										assign node79 = (inp[9]) ? node83 : node80;
											assign node80 = (inp[5]) ? 13'b0000111111111 : 13'b0001111111111;
											assign node83 = (inp[10]) ? 13'b0000011111111 : 13'b0000111111111;
										assign node86 = (inp[10]) ? node90 : node87;
											assign node87 = (inp[8]) ? 13'b0000011111111 : 13'b0000111111111;
											assign node90 = (inp[5]) ? 13'b0000001111111 : 13'b0000011111111;
								assign node93 = (inp[9]) ? node109 : node94;
									assign node94 = (inp[8]) ? node102 : node95;
										assign node95 = (inp[10]) ? node99 : node96;
											assign node96 = (inp[0]) ? 13'b0000111111111 : 13'b0001111111111;
											assign node99 = (inp[2]) ? 13'b0000011111111 : 13'b0000111111111;
										assign node102 = (inp[2]) ? node106 : node103;
											assign node103 = (inp[0]) ? 13'b0000011111111 : 13'b0000111111111;
											assign node106 = (inp[0]) ? 13'b0000001111111 : 13'b0000011111111;
									assign node109 = (inp[5]) ? node115 : node110;
										assign node110 = (inp[0]) ? 13'b0000001111111 : node111;
											assign node111 = (inp[2]) ? 13'b0000001111111 : 13'b0000111111111;
										assign node115 = (inp[2]) ? node119 : node116;
											assign node116 = (inp[8]) ? 13'b0000001111111 : 13'b0000011111111;
											assign node119 = (inp[10]) ? 13'b0000000111111 : 13'b0000001111111;
						assign node122 = (inp[8]) ? node184 : node123;
							assign node123 = (inp[5]) ? node155 : node124;
								assign node124 = (inp[9]) ? node140 : node125;
									assign node125 = (inp[7]) ? node133 : node126;
										assign node126 = (inp[2]) ? node130 : node127;
											assign node127 = (inp[10]) ? 13'b0001111111111 : 13'b0011111111111;
											assign node130 = (inp[10]) ? 13'b0000111111111 : 13'b0001111111111;
										assign node133 = (inp[2]) ? node137 : node134;
											assign node134 = (inp[10]) ? 13'b0000111111111 : 13'b0001111111111;
											assign node137 = (inp[0]) ? 13'b0000011111111 : 13'b0000111111111;
									assign node140 = (inp[3]) ? node148 : node141;
										assign node141 = (inp[0]) ? node145 : node142;
											assign node142 = (inp[10]) ? 13'b0000111111111 : 13'b0001111111111;
											assign node145 = (inp[10]) ? 13'b0000011111111 : 13'b0000111111111;
										assign node148 = (inp[10]) ? node152 : node149;
											assign node149 = (inp[2]) ? 13'b0000011111111 : 13'b0000011111111;
											assign node152 = (inp[7]) ? 13'b0000001111111 : 13'b0000011111111;
								assign node155 = (inp[0]) ? node171 : node156;
									assign node156 = (inp[3]) ? node164 : node157;
										assign node157 = (inp[9]) ? node161 : node158;
											assign node158 = (inp[2]) ? 13'b0000111111111 : 13'b0001111111111;
											assign node161 = (inp[10]) ? 13'b0000011111111 : 13'b0000111111111;
										assign node164 = (inp[10]) ? node168 : node165;
											assign node165 = (inp[2]) ? 13'b0000011111111 : 13'b0000111111111;
											assign node168 = (inp[9]) ? 13'b0000001111111 : 13'b0000011111111;
									assign node171 = (inp[10]) ? node179 : node172;
										assign node172 = (inp[7]) ? node176 : node173;
											assign node173 = (inp[9]) ? 13'b0000011111111 : 13'b0000111111111;
											assign node176 = (inp[9]) ? 13'b0000001111111 : 13'b0000011111111;
										assign node179 = (inp[7]) ? 13'b0000001111111 : node180;
											assign node180 = (inp[3]) ? 13'b0000001111111 : 13'b0000001111111;
							assign node184 = (inp[2]) ? node216 : node185;
								assign node185 = (inp[7]) ? node201 : node186;
									assign node186 = (inp[9]) ? node194 : node187;
										assign node187 = (inp[0]) ? node191 : node188;
											assign node188 = (inp[5]) ? 13'b0000111111111 : 13'b0001111111111;
											assign node191 = (inp[5]) ? 13'b0000011111111 : 13'b0000111111111;
										assign node194 = (inp[3]) ? node198 : node195;
											assign node195 = (inp[10]) ? 13'b0000011111111 : 13'b0000111111111;
											assign node198 = (inp[0]) ? 13'b0000001111111 : 13'b0000001111111;
									assign node201 = (inp[0]) ? node209 : node202;
										assign node202 = (inp[3]) ? node206 : node203;
											assign node203 = (inp[5]) ? 13'b0000011111111 : 13'b0000011111111;
											assign node206 = (inp[10]) ? 13'b0000001111111 : 13'b0000011111111;
										assign node209 = (inp[3]) ? node213 : node210;
											assign node210 = (inp[5]) ? 13'b0000001111111 : 13'b0000011111111;
											assign node213 = (inp[9]) ? 13'b0000000111111 : 13'b0000001111111;
								assign node216 = (inp[10]) ? node230 : node217;
									assign node217 = (inp[0]) ? node225 : node218;
										assign node218 = (inp[9]) ? node222 : node219;
											assign node219 = (inp[3]) ? 13'b0000011111111 : 13'b0000111111111;
											assign node222 = (inp[7]) ? 13'b0000001111111 : 13'b0000011111111;
										assign node225 = (inp[7]) ? node227 : 13'b0000001111111;
											assign node227 = (inp[3]) ? 13'b0000000111111 : 13'b0000001111111;
									assign node230 = (inp[3]) ? node238 : node231;
										assign node231 = (inp[5]) ? node235 : node232;
											assign node232 = (inp[9]) ? 13'b0000001111111 : 13'b0000011111111;
											assign node235 = (inp[0]) ? 13'b0000000111111 : 13'b0000001111111;
										assign node238 = (inp[9]) ? node242 : node239;
											assign node239 = (inp[7]) ? 13'b0000000111111 : 13'b0000001111111;
											assign node242 = (inp[0]) ? 13'b0000000011111 : 13'b0000000111111;
					assign node245 = (inp[8]) ? node365 : node246;
						assign node246 = (inp[9]) ? node304 : node247;
							assign node247 = (inp[0]) ? node275 : node248;
								assign node248 = (inp[7]) ? node262 : node249;
									assign node249 = (inp[3]) ? node255 : node250;
										assign node250 = (inp[11]) ? node252 : 13'b0001111111111;
											assign node252 = (inp[2]) ? 13'b0000111111111 : 13'b0001111111111;
										assign node255 = (inp[10]) ? node259 : node256;
											assign node256 = (inp[5]) ? 13'b0000111111111 : 13'b0000111111111;
											assign node259 = (inp[5]) ? 13'b0000011111111 : 13'b0000111111111;
									assign node262 = (inp[3]) ? node270 : node263;
										assign node263 = (inp[5]) ? node267 : node264;
											assign node264 = (inp[2]) ? 13'b0000111111111 : 13'b0000111111111;
											assign node267 = (inp[2]) ? 13'b0000011111111 : 13'b0000111111111;
										assign node270 = (inp[10]) ? 13'b0000011111111 : node271;
											assign node271 = (inp[11]) ? 13'b0000011111111 : 13'b0000111111111;
								assign node275 = (inp[3]) ? node291 : node276;
									assign node276 = (inp[7]) ? node284 : node277;
										assign node277 = (inp[2]) ? node281 : node278;
											assign node278 = (inp[10]) ? 13'b0000111111111 : 13'b0001111111111;
											assign node281 = (inp[11]) ? 13'b0000011111111 : 13'b0000111111111;
										assign node284 = (inp[5]) ? node288 : node285;
											assign node285 = (inp[10]) ? 13'b0000001111111 : 13'b0000111111111;
											assign node288 = (inp[11]) ? 13'b0000001111111 : 13'b0000011111111;
									assign node291 = (inp[5]) ? node297 : node292;
										assign node292 = (inp[2]) ? node294 : 13'b0000111111111;
											assign node294 = (inp[10]) ? 13'b0000001111111 : 13'b0000011111111;
										assign node297 = (inp[11]) ? node301 : node298;
											assign node298 = (inp[2]) ? 13'b0000001111111 : 13'b0000001111111;
											assign node301 = (inp[7]) ? 13'b0000000111111 : 13'b0000001111111;
							assign node304 = (inp[7]) ? node336 : node305;
								assign node305 = (inp[3]) ? node321 : node306;
									assign node306 = (inp[11]) ? node314 : node307;
										assign node307 = (inp[2]) ? node311 : node308;
											assign node308 = (inp[0]) ? 13'b0000111111111 : 13'b0001111111111;
											assign node311 = (inp[0]) ? 13'b0000011111111 : 13'b0000111111111;
										assign node314 = (inp[5]) ? node318 : node315;
											assign node315 = (inp[0]) ? 13'b0000011111111 : 13'b0000111111111;
											assign node318 = (inp[10]) ? 13'b0000001111111 : 13'b0000011111111;
									assign node321 = (inp[5]) ? node329 : node322;
										assign node322 = (inp[0]) ? node326 : node323;
											assign node323 = (inp[11]) ? 13'b0000011111111 : 13'b0000111111111;
											assign node326 = (inp[10]) ? 13'b0000001111111 : 13'b0000011111111;
										assign node329 = (inp[10]) ? node333 : node330;
											assign node330 = (inp[2]) ? 13'b0000000111111 : 13'b0000011111111;
											assign node333 = (inp[0]) ? 13'b0000000111111 : 13'b0000001111111;
								assign node336 = (inp[2]) ? node350 : node337;
									assign node337 = (inp[0]) ? node343 : node338;
										assign node338 = (inp[5]) ? node340 : 13'b0000111111111;
											assign node340 = (inp[10]) ? 13'b0000001111111 : 13'b0000011111111;
										assign node343 = (inp[3]) ? node347 : node344;
											assign node344 = (inp[5]) ? 13'b0000001111111 : 13'b0000011111111;
											assign node347 = (inp[11]) ? 13'b0000000111111 : 13'b0000001111111;
									assign node350 = (inp[0]) ? node358 : node351;
										assign node351 = (inp[5]) ? node355 : node352;
											assign node352 = (inp[3]) ? 13'b0000001111111 : 13'b0000001111111;
											assign node355 = (inp[3]) ? 13'b0000000111111 : 13'b0000001111111;
										assign node358 = (inp[3]) ? node362 : node359;
											assign node359 = (inp[5]) ? 13'b0000000111111 : 13'b0000001111111;
											assign node362 = (inp[10]) ? 13'b0000000011111 : 13'b0000000111111;
						assign node365 = (inp[3]) ? node427 : node366;
							assign node366 = (inp[2]) ? node396 : node367;
								assign node367 = (inp[7]) ? node381 : node368;
									assign node368 = (inp[0]) ? node376 : node369;
										assign node369 = (inp[10]) ? node373 : node370;
											assign node370 = (inp[9]) ? 13'b0000111111111 : 13'b0001111111111;
											assign node373 = (inp[9]) ? 13'b0000011111111 : 13'b0000111111111;
										assign node376 = (inp[5]) ? node378 : 13'b0000111111111;
											assign node378 = (inp[11]) ? 13'b0000001111111 : 13'b0000011111111;
									assign node381 = (inp[5]) ? node389 : node382;
										assign node382 = (inp[9]) ? node386 : node383;
											assign node383 = (inp[0]) ? 13'b0000011111111 : 13'b0000111111111;
											assign node386 = (inp[11]) ? 13'b0000001111111 : 13'b0000011111111;
										assign node389 = (inp[9]) ? node393 : node390;
											assign node390 = (inp[11]) ? 13'b0000001111111 : 13'b0000011111111;
											assign node393 = (inp[11]) ? 13'b0000000111111 : 13'b0000001111111;
								assign node396 = (inp[0]) ? node412 : node397;
									assign node397 = (inp[11]) ? node405 : node398;
										assign node398 = (inp[9]) ? node402 : node399;
											assign node399 = (inp[5]) ? 13'b0000011111111 : 13'b0000111111111;
											assign node402 = (inp[7]) ? 13'b0000001111111 : 13'b0000011111111;
										assign node405 = (inp[5]) ? node409 : node406;
											assign node406 = (inp[10]) ? 13'b0000001111111 : 13'b0000001111111;
											assign node409 = (inp[10]) ? 13'b0000000111111 : 13'b0000001111111;
									assign node412 = (inp[9]) ? node420 : node413;
										assign node413 = (inp[10]) ? node417 : node414;
											assign node414 = (inp[7]) ? 13'b0000001111111 : 13'b0000011111111;
											assign node417 = (inp[7]) ? 13'b0000000111111 : 13'b0000001111111;
										assign node420 = (inp[11]) ? node424 : node421;
											assign node421 = (inp[7]) ? 13'b0000000011111 : 13'b0000001111111;
											assign node424 = (inp[10]) ? 13'b0000000011111 : 13'b0000000011111;
							assign node427 = (inp[9]) ? node459 : node428;
								assign node428 = (inp[11]) ? node444 : node429;
									assign node429 = (inp[10]) ? node437 : node430;
										assign node430 = (inp[7]) ? node434 : node431;
											assign node431 = (inp[5]) ? 13'b0000011111111 : 13'b0000111111111;
											assign node434 = (inp[0]) ? 13'b0000000111111 : 13'b0000011111111;
										assign node437 = (inp[0]) ? node441 : node438;
											assign node438 = (inp[7]) ? 13'b0000001111111 : 13'b0000011111111;
											assign node441 = (inp[7]) ? 13'b0000000111111 : 13'b0000001111111;
									assign node444 = (inp[2]) ? node452 : node445;
										assign node445 = (inp[7]) ? node449 : node446;
											assign node446 = (inp[10]) ? 13'b0000001111111 : 13'b0000001111111;
											assign node449 = (inp[5]) ? 13'b0000000111111 : 13'b0000001111111;
										assign node452 = (inp[0]) ? node456 : node453;
											assign node453 = (inp[10]) ? 13'b0000000111111 : 13'b0000001111111;
											assign node456 = (inp[10]) ? 13'b0000000011111 : 13'b0000000111111;
								assign node459 = (inp[0]) ? node473 : node460;
									assign node460 = (inp[5]) ? node466 : node461;
										assign node461 = (inp[2]) ? node463 : 13'b0000011111111;
											assign node463 = (inp[11]) ? 13'b0000000111111 : 13'b0000001111111;
										assign node466 = (inp[11]) ? node470 : node467;
											assign node467 = (inp[10]) ? 13'b0000000111111 : 13'b0000001111111;
											assign node470 = (inp[2]) ? 13'b0000000011111 : 13'b0000000011111;
									assign node473 = (inp[7]) ? node479 : node474;
										assign node474 = (inp[11]) ? node476 : 13'b0000000111111;
											assign node476 = (inp[10]) ? 13'b0000000011111 : 13'b0000000111111;
										assign node479 = (inp[5]) ? node483 : node480;
											assign node480 = (inp[2]) ? 13'b0000000011111 : 13'b0000000111111;
											assign node483 = (inp[2]) ? 13'b0000000001111 : 13'b0000000001111;
				assign node486 = (inp[5]) ? node730 : node487;
					assign node487 = (inp[1]) ? node611 : node488;
						assign node488 = (inp[2]) ? node552 : node489;
							assign node489 = (inp[7]) ? node521 : node490;
								assign node490 = (inp[8]) ? node506 : node491;
									assign node491 = (inp[10]) ? node499 : node492;
										assign node492 = (inp[0]) ? node496 : node493;
											assign node493 = (inp[11]) ? 13'b0001111111111 : 13'b0111111111111;
											assign node496 = (inp[11]) ? 13'b0000011111111 : 13'b0001111111111;
										assign node499 = (inp[11]) ? node503 : node500;
											assign node500 = (inp[0]) ? 13'b0000111111111 : 13'b0001111111111;
											assign node503 = (inp[0]) ? 13'b0000011111111 : 13'b0000111111111;
									assign node506 = (inp[0]) ? node514 : node507;
										assign node507 = (inp[9]) ? node511 : node508;
											assign node508 = (inp[11]) ? 13'b0000111111111 : 13'b0000111111111;
											assign node511 = (inp[11]) ? 13'b0000011111111 : 13'b0000111111111;
										assign node514 = (inp[11]) ? node518 : node515;
											assign node515 = (inp[10]) ? 13'b0000011111111 : 13'b0000111111111;
											assign node518 = (inp[9]) ? 13'b0000001111111 : 13'b0000011111111;
								assign node521 = (inp[10]) ? node537 : node522;
									assign node522 = (inp[0]) ? node530 : node523;
										assign node523 = (inp[9]) ? node527 : node524;
											assign node524 = (inp[3]) ? 13'b0000111111111 : 13'b0001111111111;
											assign node527 = (inp[8]) ? 13'b0000011111111 : 13'b0000111111111;
										assign node530 = (inp[3]) ? node534 : node531;
											assign node531 = (inp[11]) ? 13'b0000011111111 : 13'b0000111111111;
											assign node534 = (inp[11]) ? 13'b0000000111111 : 13'b0000011111111;
									assign node537 = (inp[8]) ? node545 : node538;
										assign node538 = (inp[9]) ? node542 : node539;
											assign node539 = (inp[11]) ? 13'b0000011111111 : 13'b0000111111111;
											assign node542 = (inp[3]) ? 13'b0000001111111 : 13'b0000011111111;
										assign node545 = (inp[0]) ? node549 : node546;
											assign node546 = (inp[11]) ? 13'b0000001111111 : 13'b0000011111111;
											assign node549 = (inp[9]) ? 13'b0000000111111 : 13'b0000000111111;
							assign node552 = (inp[9]) ? node582 : node553;
								assign node553 = (inp[7]) ? node567 : node554;
									assign node554 = (inp[3]) ? node562 : node555;
										assign node555 = (inp[11]) ? node559 : node556;
											assign node556 = (inp[0]) ? 13'b0000111111111 : 13'b0001111111111;
											assign node559 = (inp[0]) ? 13'b0000011111111 : 13'b0000111111111;
										assign node562 = (inp[11]) ? 13'b0000011111111 : node563;
											assign node563 = (inp[10]) ? 13'b0000011111111 : 13'b0000111111111;
									assign node567 = (inp[0]) ? node575 : node568;
										assign node568 = (inp[11]) ? node572 : node569;
											assign node569 = (inp[10]) ? 13'b0000011111111 : 13'b0000111111111;
											assign node572 = (inp[10]) ? 13'b0000001111111 : 13'b0000011111111;
										assign node575 = (inp[11]) ? node579 : node576;
											assign node576 = (inp[3]) ? 13'b0000001111111 : 13'b0000011111111;
											assign node579 = (inp[8]) ? 13'b0000000011111 : 13'b0000001111111;
								assign node582 = (inp[8]) ? node598 : node583;
									assign node583 = (inp[0]) ? node591 : node584;
										assign node584 = (inp[10]) ? node588 : node585;
											assign node585 = (inp[7]) ? 13'b0000001111111 : 13'b0000111111111;
											assign node588 = (inp[3]) ? 13'b0000001111111 : 13'b0000011111111;
										assign node591 = (inp[11]) ? node595 : node592;
											assign node592 = (inp[7]) ? 13'b0000001111111 : 13'b0000011111111;
											assign node595 = (inp[3]) ? 13'b0000000111111 : 13'b0000001111111;
									assign node598 = (inp[3]) ? node604 : node599;
										assign node599 = (inp[0]) ? 13'b0000001111111 : node600;
											assign node600 = (inp[10]) ? 13'b0000001111111 : 13'b0000011111111;
										assign node604 = (inp[10]) ? node608 : node605;
											assign node605 = (inp[0]) ? 13'b0000000111111 : 13'b0000001111111;
											assign node608 = (inp[11]) ? 13'b0000000011111 : 13'b0000000111111;
						assign node611 = (inp[2]) ? node671 : node612;
							assign node612 = (inp[9]) ? node642 : node613;
								assign node613 = (inp[7]) ? node627 : node614;
									assign node614 = (inp[3]) ? node622 : node615;
										assign node615 = (inp[10]) ? node619 : node616;
											assign node616 = (inp[8]) ? 13'b0000111111111 : 13'b0001111111111;
											assign node619 = (inp[8]) ? 13'b0000011111111 : 13'b0000111111111;
										assign node622 = (inp[11]) ? node624 : 13'b0000111111111;
											assign node624 = (inp[0]) ? 13'b0000011111111 : 13'b0000011111111;
									assign node627 = (inp[11]) ? node635 : node628;
										assign node628 = (inp[8]) ? node632 : node629;
											assign node629 = (inp[10]) ? 13'b0000011111111 : 13'b0000111111111;
											assign node632 = (inp[3]) ? 13'b0000001111111 : 13'b0000111111111;
										assign node635 = (inp[0]) ? node639 : node636;
											assign node636 = (inp[3]) ? 13'b0000001111111 : 13'b0000001111111;
											assign node639 = (inp[3]) ? 13'b0000001111111 : 13'b0000011111111;
								assign node642 = (inp[7]) ? node658 : node643;
									assign node643 = (inp[8]) ? node651 : node644;
										assign node644 = (inp[10]) ? node648 : node645;
											assign node645 = (inp[11]) ? 13'b0000011111111 : 13'b0000011111111;
											assign node648 = (inp[0]) ? 13'b0000001111111 : 13'b0000011111111;
										assign node651 = (inp[11]) ? node655 : node652;
											assign node652 = (inp[10]) ? 13'b0000001111111 : 13'b0000011111111;
											assign node655 = (inp[3]) ? 13'b0000000111111 : 13'b0000001111111;
									assign node658 = (inp[10]) ? node666 : node659;
										assign node659 = (inp[0]) ? node663 : node660;
											assign node660 = (inp[11]) ? 13'b0000001111111 : 13'b0000001111111;
											assign node663 = (inp[3]) ? 13'b0000000111111 : 13'b0000001111111;
										assign node666 = (inp[8]) ? node668 : 13'b0000001111111;
											assign node668 = (inp[3]) ? 13'b0000000011111 : 13'b0000000111111;
							assign node671 = (inp[3]) ? node701 : node672;
								assign node672 = (inp[10]) ? node686 : node673;
									assign node673 = (inp[8]) ? node681 : node674;
										assign node674 = (inp[9]) ? node678 : node675;
											assign node675 = (inp[0]) ? 13'b0000001111111 : 13'b0000111111111;
											assign node678 = (inp[0]) ? 13'b0000001111111 : 13'b0000011111111;
										assign node681 = (inp[0]) ? 13'b0000000111111 : node682;
											assign node682 = (inp[7]) ? 13'b0000001111111 : 13'b0000011111111;
									assign node686 = (inp[8]) ? node694 : node687;
										assign node687 = (inp[0]) ? node691 : node688;
											assign node688 = (inp[7]) ? 13'b0000001111111 : 13'b0000011111111;
											assign node691 = (inp[9]) ? 13'b0000000111111 : 13'b0000001111111;
										assign node694 = (inp[9]) ? node698 : node695;
											assign node695 = (inp[0]) ? 13'b0000000111111 : 13'b0000001111111;
											assign node698 = (inp[7]) ? 13'b0000000011111 : 13'b0000000111111;
								assign node701 = (inp[9]) ? node717 : node702;
									assign node702 = (inp[7]) ? node710 : node703;
										assign node703 = (inp[8]) ? node707 : node704;
											assign node704 = (inp[10]) ? 13'b0000001111111 : 13'b0000011111111;
											assign node707 = (inp[0]) ? 13'b0000000111111 : 13'b0000001111111;
										assign node710 = (inp[0]) ? node714 : node711;
											assign node711 = (inp[8]) ? 13'b0000000011111 : 13'b0000001111111;
											assign node714 = (inp[10]) ? 13'b0000000011111 : 13'b0000000111111;
									assign node717 = (inp[7]) ? node723 : node718;
										assign node718 = (inp[0]) ? node720 : 13'b0000000111111;
											assign node720 = (inp[10]) ? 13'b0000000001111 : 13'b0000000111111;
										assign node723 = (inp[8]) ? node727 : node724;
											assign node724 = (inp[10]) ? 13'b0000000001111 : 13'b0000000111111;
											assign node727 = (inp[0]) ? 13'b0000000001111 : 13'b0000000001111;
					assign node730 = (inp[10]) ? node848 : node731;
						assign node731 = (inp[11]) ? node789 : node732;
							assign node732 = (inp[3]) ? node760 : node733;
								assign node733 = (inp[8]) ? node747 : node734;
									assign node734 = (inp[9]) ? node742 : node735;
										assign node735 = (inp[2]) ? node739 : node736;
											assign node736 = (inp[7]) ? 13'b0000111111111 : 13'b0001111111111;
											assign node739 = (inp[7]) ? 13'b0000011111111 : 13'b0000111111111;
										assign node742 = (inp[2]) ? 13'b0000001111111 : node743;
											assign node743 = (inp[0]) ? 13'b0000011111111 : 13'b0000111111111;
									assign node747 = (inp[1]) ? node755 : node748;
										assign node748 = (inp[7]) ? node752 : node749;
											assign node749 = (inp[2]) ? 13'b0000011111111 : 13'b0000111111111;
											assign node752 = (inp[2]) ? 13'b0000001111111 : 13'b0000011111111;
										assign node755 = (inp[2]) ? node757 : 13'b0000001111111;
											assign node757 = (inp[9]) ? 13'b0000000111111 : 13'b0000001111111;
								assign node760 = (inp[8]) ? node776 : node761;
									assign node761 = (inp[9]) ? node769 : node762;
										assign node762 = (inp[7]) ? node766 : node763;
											assign node763 = (inp[2]) ? 13'b0000011111111 : 13'b0000111111111;
											assign node766 = (inp[1]) ? 13'b0000001111111 : 13'b0000011111111;
										assign node769 = (inp[0]) ? node773 : node770;
											assign node770 = (inp[7]) ? 13'b0000001111111 : 13'b0000011111111;
											assign node773 = (inp[2]) ? 13'b0000000111111 : 13'b0000001111111;
									assign node776 = (inp[1]) ? node782 : node777;
										assign node777 = (inp[0]) ? 13'b0000001111111 : node778;
											assign node778 = (inp[7]) ? 13'b0000001111111 : 13'b0000011111111;
										assign node782 = (inp[7]) ? node786 : node783;
											assign node783 = (inp[2]) ? 13'b0000000111111 : 13'b0000001111111;
											assign node786 = (inp[2]) ? 13'b0000000011111 : 13'b0000000111111;
							assign node789 = (inp[9]) ? node821 : node790;
								assign node790 = (inp[0]) ? node806 : node791;
									assign node791 = (inp[1]) ? node799 : node792;
										assign node792 = (inp[2]) ? node796 : node793;
											assign node793 = (inp[3]) ? 13'b0000011111111 : 13'b0000111111111;
											assign node796 = (inp[3]) ? 13'b0000001111111 : 13'b0000011111111;
										assign node799 = (inp[3]) ? node803 : node800;
											assign node800 = (inp[2]) ? 13'b0000001111111 : 13'b0000011111111;
											assign node803 = (inp[7]) ? 13'b0000000111111 : 13'b0000001111111;
									assign node806 = (inp[7]) ? node814 : node807;
										assign node807 = (inp[8]) ? node811 : node808;
											assign node808 = (inp[2]) ? 13'b0000001111111 : 13'b0000011111111;
											assign node811 = (inp[3]) ? 13'b0000000111111 : 13'b0000001111111;
										assign node814 = (inp[2]) ? node818 : node815;
											assign node815 = (inp[8]) ? 13'b0000000111111 : 13'b0000001111111;
											assign node818 = (inp[1]) ? 13'b0000000001111 : 13'b0000000111111;
								assign node821 = (inp[0]) ? node835 : node822;
									assign node822 = (inp[1]) ? node830 : node823;
										assign node823 = (inp[2]) ? node827 : node824;
											assign node824 = (inp[8]) ? 13'b0000001111111 : 13'b0000011111111;
											assign node827 = (inp[3]) ? 13'b0000000111111 : 13'b0000001111111;
										assign node830 = (inp[2]) ? node832 : 13'b0000000111111;
											assign node832 = (inp[7]) ? 13'b0000000011111 : 13'b0000001111111;
									assign node835 = (inp[2]) ? node843 : node836;
										assign node836 = (inp[3]) ? node840 : node837;
											assign node837 = (inp[7]) ? 13'b0000000111111 : 13'b0000011111111;
											assign node840 = (inp[8]) ? 13'b0000000011111 : 13'b0000000111111;
										assign node843 = (inp[1]) ? node845 : 13'b0000000011111;
											assign node845 = (inp[7]) ? 13'b0000000001111 : 13'b0000000011111;
						assign node848 = (inp[7]) ? node910 : node849;
							assign node849 = (inp[3]) ? node881 : node850;
								assign node850 = (inp[2]) ? node866 : node851;
									assign node851 = (inp[11]) ? node859 : node852;
										assign node852 = (inp[0]) ? node856 : node853;
											assign node853 = (inp[9]) ? 13'b0000011111111 : 13'b0000111111111;
											assign node856 = (inp[1]) ? 13'b0000001111111 : 13'b0000011111111;
										assign node859 = (inp[1]) ? node863 : node860;
											assign node860 = (inp[9]) ? 13'b0000001111111 : 13'b0000011111111;
											assign node863 = (inp[8]) ? 13'b0000000111111 : 13'b0000001111111;
									assign node866 = (inp[8]) ? node874 : node867;
										assign node867 = (inp[11]) ? node871 : node868;
											assign node868 = (inp[0]) ? 13'b0000001111111 : 13'b0000011111111;
											assign node871 = (inp[0]) ? 13'b0000000111111 : 13'b0000001111111;
										assign node874 = (inp[11]) ? node878 : node875;
											assign node875 = (inp[0]) ? 13'b0000000111111 : 13'b0000001111111;
											assign node878 = (inp[9]) ? 13'b0000000011111 : 13'b0000000111111;
								assign node881 = (inp[9]) ? node897 : node882;
									assign node882 = (inp[8]) ? node890 : node883;
										assign node883 = (inp[1]) ? node887 : node884;
											assign node884 = (inp[0]) ? 13'b0000001111111 : 13'b0000001111111;
											assign node887 = (inp[0]) ? 13'b0000000011111 : 13'b0000001111111;
										assign node890 = (inp[2]) ? node894 : node891;
											assign node891 = (inp[11]) ? 13'b0000000111111 : 13'b0000001111111;
											assign node894 = (inp[11]) ? 13'b0000000001111 : 13'b0000000111111;
									assign node897 = (inp[0]) ? node903 : node898;
										assign node898 = (inp[1]) ? 13'b0000000011111 : node899;
											assign node899 = (inp[8]) ? 13'b0000000111111 : 13'b0000001111111;
										assign node903 = (inp[11]) ? node907 : node904;
											assign node904 = (inp[2]) ? 13'b0000000011111 : 13'b0000000111111;
											assign node907 = (inp[2]) ? 13'b0000000001111 : 13'b0000000011111;
							assign node910 = (inp[11]) ? node942 : node911;
								assign node911 = (inp[0]) ? node927 : node912;
									assign node912 = (inp[9]) ? node920 : node913;
										assign node913 = (inp[2]) ? node917 : node914;
											assign node914 = (inp[1]) ? 13'b0000001111111 : 13'b0000011111111;
											assign node917 = (inp[3]) ? 13'b0000000111111 : 13'b0000001111111;
										assign node920 = (inp[1]) ? node924 : node921;
											assign node921 = (inp[2]) ? 13'b0000000111111 : 13'b0000001111111;
											assign node924 = (inp[8]) ? 13'b0000000011111 : 13'b0000000111111;
									assign node927 = (inp[1]) ? node935 : node928;
										assign node928 = (inp[9]) ? node932 : node929;
											assign node929 = (inp[3]) ? 13'b0000000111111 : 13'b0000011111111;
											assign node932 = (inp[3]) ? 13'b0000000011111 : 13'b0000000111111;
										assign node935 = (inp[8]) ? node939 : node936;
											assign node936 = (inp[2]) ? 13'b0000000011111 : 13'b0000000111111;
											assign node939 = (inp[3]) ? 13'b0000000001111 : 13'b0000000011111;
								assign node942 = (inp[9]) ? node958 : node943;
									assign node943 = (inp[2]) ? node951 : node944;
										assign node944 = (inp[8]) ? node948 : node945;
											assign node945 = (inp[1]) ? 13'b0000000111111 : 13'b0000000111111;
											assign node948 = (inp[1]) ? 13'b0000000011111 : 13'b0000000111111;
										assign node951 = (inp[3]) ? node955 : node952;
											assign node952 = (inp[8]) ? 13'b0000000011111 : 13'b0000000111111;
											assign node955 = (inp[8]) ? 13'b0000000001111 : 13'b0000000011111;
									assign node958 = (inp[3]) ? node966 : node959;
										assign node959 = (inp[2]) ? node963 : node960;
											assign node960 = (inp[8]) ? 13'b0000000011111 : 13'b0000000111111;
											assign node963 = (inp[1]) ? 13'b0000000001111 : 13'b0000000011111;
										assign node966 = (inp[2]) ? node970 : node967;
											assign node967 = (inp[1]) ? 13'b0000000001111 : 13'b0000000011111;
											assign node970 = (inp[0]) ? 13'b0000000000111 : 13'b0000000001111;
			assign node973 = (inp[9]) ? node1461 : node974;
				assign node974 = (inp[8]) ? node1214 : node975;
					assign node975 = (inp[0]) ? node1097 : node976;
						assign node976 = (inp[1]) ? node1038 : node977;
							assign node977 = (inp[5]) ? node1007 : node978;
								assign node978 = (inp[6]) ? node994 : node979;
									assign node979 = (inp[7]) ? node987 : node980;
										assign node980 = (inp[3]) ? node984 : node981;
											assign node981 = (inp[2]) ? 13'b0001111111111 : 13'b0011111111111;
											assign node984 = (inp[11]) ? 13'b0000111111111 : 13'b0001111111111;
										assign node987 = (inp[11]) ? node991 : node988;
											assign node988 = (inp[3]) ? 13'b0000111111111 : 13'b0001111111111;
											assign node991 = (inp[10]) ? 13'b0000011111111 : 13'b0000111111111;
									assign node994 = (inp[3]) ? node1000 : node995;
										assign node995 = (inp[7]) ? node997 : 13'b0001111111111;
											assign node997 = (inp[2]) ? 13'b0000011111111 : 13'b0000111111111;
										assign node1000 = (inp[2]) ? node1004 : node1001;
											assign node1001 = (inp[7]) ? 13'b0000011111111 : 13'b0000111111111;
											assign node1004 = (inp[10]) ? 13'b0000001111111 : 13'b0000011111111;
								assign node1007 = (inp[7]) ? node1023 : node1008;
									assign node1008 = (inp[6]) ? node1016 : node1009;
										assign node1009 = (inp[11]) ? node1013 : node1010;
											assign node1010 = (inp[10]) ? 13'b0000111111111 : 13'b0001111111111;
											assign node1013 = (inp[10]) ? 13'b0000011111111 : 13'b0000111111111;
										assign node1016 = (inp[3]) ? node1020 : node1017;
											assign node1017 = (inp[10]) ? 13'b0000011111111 : 13'b0000111111111;
											assign node1020 = (inp[2]) ? 13'b0000001111111 : 13'b0000011111111;
									assign node1023 = (inp[11]) ? node1031 : node1024;
										assign node1024 = (inp[2]) ? node1028 : node1025;
											assign node1025 = (inp[6]) ? 13'b0000011111111 : 13'b0000011111111;
											assign node1028 = (inp[3]) ? 13'b0000001111111 : 13'b0000001111111;
										assign node1031 = (inp[2]) ? node1035 : node1032;
											assign node1032 = (inp[3]) ? 13'b0000001111111 : 13'b0000011111111;
											assign node1035 = (inp[10]) ? 13'b0000000111111 : 13'b0000011111111;
							assign node1038 = (inp[3]) ? node1070 : node1039;
								assign node1039 = (inp[10]) ? node1055 : node1040;
									assign node1040 = (inp[2]) ? node1048 : node1041;
										assign node1041 = (inp[7]) ? node1045 : node1042;
											assign node1042 = (inp[6]) ? 13'b0000111111111 : 13'b0001111111111;
											assign node1045 = (inp[6]) ? 13'b0000011111111 : 13'b0000111111111;
										assign node1048 = (inp[5]) ? node1052 : node1049;
											assign node1049 = (inp[11]) ? 13'b0000011111111 : 13'b0000111111111;
											assign node1052 = (inp[6]) ? 13'b0000001111111 : 13'b0000011111111;
									assign node1055 = (inp[6]) ? node1063 : node1056;
										assign node1056 = (inp[5]) ? node1060 : node1057;
											assign node1057 = (inp[11]) ? 13'b0000011111111 : 13'b0000111111111;
											assign node1060 = (inp[11]) ? 13'b0000001111111 : 13'b0000011111111;
										assign node1063 = (inp[2]) ? node1067 : node1064;
											assign node1064 = (inp[11]) ? 13'b0000000111111 : 13'b0000011111111;
											assign node1067 = (inp[7]) ? 13'b0000000111111 : 13'b0000001111111;
								assign node1070 = (inp[7]) ? node1082 : node1071;
									assign node1071 = (inp[10]) ? node1077 : node1072;
										assign node1072 = (inp[2]) ? node1074 : 13'b0000011111111;
											assign node1074 = (inp[11]) ? 13'b0000001111111 : 13'b0000011111111;
										assign node1077 = (inp[11]) ? 13'b0000001111111 : node1078;
											assign node1078 = (inp[2]) ? 13'b0000001111111 : 13'b0000011111111;
									assign node1082 = (inp[2]) ? node1090 : node1083;
										assign node1083 = (inp[6]) ? node1087 : node1084;
											assign node1084 = (inp[10]) ? 13'b0000001111111 : 13'b0000011111111;
											assign node1087 = (inp[5]) ? 13'b0000000111111 : 13'b0000000111111;
										assign node1090 = (inp[11]) ? node1094 : node1091;
											assign node1091 = (inp[5]) ? 13'b0000000111111 : 13'b0000001111111;
											assign node1094 = (inp[5]) ? 13'b0000000011111 : 13'b0000000111111;
						assign node1097 = (inp[6]) ? node1155 : node1098;
							assign node1098 = (inp[7]) ? node1130 : node1099;
								assign node1099 = (inp[11]) ? node1115 : node1100;
									assign node1100 = (inp[1]) ? node1108 : node1101;
										assign node1101 = (inp[2]) ? node1105 : node1102;
											assign node1102 = (inp[5]) ? 13'b0000111111111 : 13'b0001111111111;
											assign node1105 = (inp[3]) ? 13'b0000001111111 : 13'b0000111111111;
										assign node1108 = (inp[5]) ? node1112 : node1109;
											assign node1109 = (inp[3]) ? 13'b0000011111111 : 13'b0000111111111;
											assign node1112 = (inp[3]) ? 13'b0000001111111 : 13'b0000001111111;
									assign node1115 = (inp[3]) ? node1123 : node1116;
										assign node1116 = (inp[1]) ? node1120 : node1117;
											assign node1117 = (inp[10]) ? 13'b0000011111111 : 13'b0000111111111;
											assign node1120 = (inp[5]) ? 13'b0000001111111 : 13'b0000011111111;
										assign node1123 = (inp[5]) ? node1127 : node1124;
											assign node1124 = (inp[10]) ? 13'b0000001111111 : 13'b0000011111111;
											assign node1127 = (inp[2]) ? 13'b0000000111111 : 13'b0000001111111;
								assign node1130 = (inp[5]) ? node1140 : node1131;
									assign node1131 = (inp[3]) ? 13'b0000001111111 : node1132;
										assign node1132 = (inp[1]) ? node1136 : node1133;
											assign node1133 = (inp[11]) ? 13'b0000011111111 : 13'b0000011111111;
											assign node1136 = (inp[11]) ? 13'b0000001111111 : 13'b0000011111111;
									assign node1140 = (inp[2]) ? node1148 : node1141;
										assign node1141 = (inp[10]) ? node1145 : node1142;
											assign node1142 = (inp[11]) ? 13'b0000001111111 : 13'b0000011111111;
											assign node1145 = (inp[11]) ? 13'b0000000111111 : 13'b0000001111111;
										assign node1148 = (inp[3]) ? node1152 : node1149;
											assign node1149 = (inp[10]) ? 13'b0000000111111 : 13'b0000001111111;
											assign node1152 = (inp[1]) ? 13'b0000000011111 : 13'b0000000111111;
							assign node1155 = (inp[10]) ? node1185 : node1156;
								assign node1156 = (inp[2]) ? node1170 : node1157;
									assign node1157 = (inp[5]) ? node1165 : node1158;
										assign node1158 = (inp[1]) ? node1162 : node1159;
											assign node1159 = (inp[7]) ? 13'b0000011111111 : 13'b0000111111111;
											assign node1162 = (inp[3]) ? 13'b0000001111111 : 13'b0000011111111;
										assign node1165 = (inp[11]) ? node1167 : 13'b0000011111111;
											assign node1167 = (inp[7]) ? 13'b0000000111111 : 13'b0000001111111;
									assign node1170 = (inp[7]) ? node1178 : node1171;
										assign node1171 = (inp[11]) ? node1175 : node1172;
											assign node1172 = (inp[1]) ? 13'b0000001111111 : 13'b0000011111111;
											assign node1175 = (inp[1]) ? 13'b0000000111111 : 13'b0000001111111;
										assign node1178 = (inp[11]) ? node1182 : node1179;
											assign node1179 = (inp[3]) ? 13'b0000000111111 : 13'b0000011111111;
											assign node1182 = (inp[5]) ? 13'b0000000011111 : 13'b0000000111111;
								assign node1185 = (inp[5]) ? node1199 : node1186;
									assign node1186 = (inp[1]) ? node1194 : node1187;
										assign node1187 = (inp[7]) ? node1191 : node1188;
											assign node1188 = (inp[11]) ? 13'b0000001111111 : 13'b0000011111111;
											assign node1191 = (inp[2]) ? 13'b0000000111111 : 13'b0000000111111;
										assign node1194 = (inp[11]) ? 13'b0000000011111 : node1195;
											assign node1195 = (inp[2]) ? 13'b0000000111111 : 13'b0000000111111;
									assign node1199 = (inp[2]) ? node1207 : node1200;
										assign node1200 = (inp[11]) ? node1204 : node1201;
											assign node1201 = (inp[7]) ? 13'b0000000111111 : 13'b0000000111111;
											assign node1204 = (inp[1]) ? 13'b0000000001111 : 13'b0000000111111;
										assign node1207 = (inp[1]) ? node1211 : node1208;
											assign node1208 = (inp[7]) ? 13'b0000000011111 : 13'b0000000011111;
											assign node1211 = (inp[11]) ? 13'b0000000000111 : 13'b0000000011111;
					assign node1214 = (inp[0]) ? node1334 : node1215;
						assign node1215 = (inp[2]) ? node1271 : node1216;
							assign node1216 = (inp[11]) ? node1246 : node1217;
								assign node1217 = (inp[7]) ? node1231 : node1218;
									assign node1218 = (inp[6]) ? node1224 : node1219;
										assign node1219 = (inp[5]) ? 13'b0000111111111 : node1220;
											assign node1220 = (inp[10]) ? 13'b0000111111111 : 13'b0001111111111;
										assign node1224 = (inp[10]) ? node1228 : node1225;
											assign node1225 = (inp[3]) ? 13'b0000011111111 : 13'b0000111111111;
											assign node1228 = (inp[5]) ? 13'b0000001111111 : 13'b0000011111111;
									assign node1231 = (inp[10]) ? node1239 : node1232;
										assign node1232 = (inp[3]) ? node1236 : node1233;
											assign node1233 = (inp[1]) ? 13'b0000011111111 : 13'b0000111111111;
											assign node1236 = (inp[5]) ? 13'b0000001111111 : 13'b0000011111111;
										assign node1239 = (inp[6]) ? node1243 : node1240;
											assign node1240 = (inp[5]) ? 13'b0000001111111 : 13'b0000011111111;
											assign node1243 = (inp[3]) ? 13'b0000000111111 : 13'b0000001111111;
								assign node1246 = (inp[10]) ? node1260 : node1247;
									assign node1247 = (inp[1]) ? node1253 : node1248;
										assign node1248 = (inp[5]) ? node1250 : 13'b0000111111111;
											assign node1250 = (inp[7]) ? 13'b0000001111111 : 13'b0000011111111;
										assign node1253 = (inp[3]) ? node1257 : node1254;
											assign node1254 = (inp[7]) ? 13'b0000001111111 : 13'b0000011111111;
											assign node1257 = (inp[5]) ? 13'b0000000111111 : 13'b0000001111111;
									assign node1260 = (inp[1]) ? node1266 : node1261;
										assign node1261 = (inp[7]) ? node1263 : 13'b0000001111111;
											assign node1263 = (inp[6]) ? 13'b0000000111111 : 13'b0000001111111;
										assign node1266 = (inp[3]) ? node1268 : 13'b0000000111111;
											assign node1268 = (inp[5]) ? 13'b0000000011111 : 13'b0000000111111;
							assign node1271 = (inp[5]) ? node1303 : node1272;
								assign node1272 = (inp[6]) ? node1288 : node1273;
									assign node1273 = (inp[3]) ? node1281 : node1274;
										assign node1274 = (inp[11]) ? node1278 : node1275;
											assign node1275 = (inp[7]) ? 13'b0000011111111 : 13'b0000111111111;
											assign node1278 = (inp[1]) ? 13'b0000001111111 : 13'b0000011111111;
										assign node1281 = (inp[10]) ? node1285 : node1282;
											assign node1282 = (inp[11]) ? 13'b0000001111111 : 13'b0000111111111;
											assign node1285 = (inp[11]) ? 13'b0000000111111 : 13'b0000001111111;
									assign node1288 = (inp[10]) ? node1296 : node1289;
										assign node1289 = (inp[7]) ? node1293 : node1290;
											assign node1290 = (inp[11]) ? 13'b0000001111111 : 13'b0000011111111;
											assign node1293 = (inp[1]) ? 13'b0000000011111 : 13'b0000001111111;
										assign node1296 = (inp[11]) ? node1300 : node1297;
											assign node1297 = (inp[1]) ? 13'b0000000111111 : 13'b0000001111111;
											assign node1300 = (inp[7]) ? 13'b0000000011111 : 13'b0000000111111;
								assign node1303 = (inp[7]) ? node1319 : node1304;
									assign node1304 = (inp[6]) ? node1312 : node1305;
										assign node1305 = (inp[3]) ? node1309 : node1306;
											assign node1306 = (inp[1]) ? 13'b0000001111111 : 13'b0000001111111;
											assign node1309 = (inp[11]) ? 13'b0000000111111 : 13'b0000001111111;
										assign node1312 = (inp[10]) ? node1316 : node1313;
											assign node1313 = (inp[1]) ? 13'b0000000111111 : 13'b0000000111111;
											assign node1316 = (inp[3]) ? 13'b0000000011111 : 13'b0000000111111;
									assign node1319 = (inp[6]) ? node1327 : node1320;
										assign node1320 = (inp[1]) ? node1324 : node1321;
											assign node1321 = (inp[10]) ? 13'b0000000111111 : 13'b0000001111111;
											assign node1324 = (inp[10]) ? 13'b0000000011111 : 13'b0000000111111;
										assign node1327 = (inp[10]) ? node1331 : node1328;
											assign node1328 = (inp[11]) ? 13'b0000000011111 : 13'b0000000111111;
											assign node1331 = (inp[3]) ? 13'b0000000001111 : 13'b0000000011111;
						assign node1334 = (inp[7]) ? node1398 : node1335;
							assign node1335 = (inp[11]) ? node1367 : node1336;
								assign node1336 = (inp[2]) ? node1352 : node1337;
									assign node1337 = (inp[5]) ? node1345 : node1338;
										assign node1338 = (inp[3]) ? node1342 : node1339;
											assign node1339 = (inp[10]) ? 13'b0000011111111 : 13'b0000111111111;
											assign node1342 = (inp[1]) ? 13'b0000001111111 : 13'b0000011111111;
										assign node1345 = (inp[10]) ? node1349 : node1346;
											assign node1346 = (inp[6]) ? 13'b0000001111111 : 13'b0000011111111;
											assign node1349 = (inp[3]) ? 13'b0000000111111 : 13'b0000001111111;
									assign node1352 = (inp[5]) ? node1360 : node1353;
										assign node1353 = (inp[3]) ? node1357 : node1354;
											assign node1354 = (inp[1]) ? 13'b0000001111111 : 13'b0000011111111;
											assign node1357 = (inp[1]) ? 13'b0000000111111 : 13'b0000001111111;
										assign node1360 = (inp[1]) ? node1364 : node1361;
											assign node1361 = (inp[3]) ? 13'b0000000111111 : 13'b0000001111111;
											assign node1364 = (inp[10]) ? 13'b0000000001111 : 13'b0000000111111;
								assign node1367 = (inp[6]) ? node1383 : node1368;
									assign node1368 = (inp[2]) ? node1376 : node1369;
										assign node1369 = (inp[5]) ? node1373 : node1370;
											assign node1370 = (inp[1]) ? 13'b0000001111111 : 13'b0000111111111;
											assign node1373 = (inp[1]) ? 13'b0000000111111 : 13'b0000001111111;
										assign node1376 = (inp[3]) ? node1380 : node1377;
											assign node1377 = (inp[10]) ? 13'b0000000011111 : 13'b0000001111111;
											assign node1380 = (inp[5]) ? 13'b0000000011111 : 13'b0000000111111;
									assign node1383 = (inp[5]) ? node1391 : node1384;
										assign node1384 = (inp[3]) ? node1388 : node1385;
											assign node1385 = (inp[10]) ? 13'b0000000111111 : 13'b0000000111111;
											assign node1388 = (inp[1]) ? 13'b0000000011111 : 13'b0000000111111;
										assign node1391 = (inp[3]) ? node1395 : node1392;
											assign node1392 = (inp[10]) ? 13'b0000000011111 : 13'b0000000111111;
											assign node1395 = (inp[1]) ? 13'b0000000001111 : 13'b0000000011111;
							assign node1398 = (inp[10]) ? node1430 : node1399;
								assign node1399 = (inp[1]) ? node1415 : node1400;
									assign node1400 = (inp[6]) ? node1408 : node1401;
										assign node1401 = (inp[11]) ? node1405 : node1402;
											assign node1402 = (inp[2]) ? 13'b0000001111111 : 13'b0000011111111;
											assign node1405 = (inp[2]) ? 13'b0000000111111 : 13'b0000001111111;
										assign node1408 = (inp[5]) ? node1412 : node1409;
											assign node1409 = (inp[3]) ? 13'b0000000111111 : 13'b0000001111111;
											assign node1412 = (inp[2]) ? 13'b0000000011111 : 13'b0000000111111;
									assign node1415 = (inp[3]) ? node1423 : node1416;
										assign node1416 = (inp[5]) ? node1420 : node1417;
											assign node1417 = (inp[2]) ? 13'b0000000111111 : 13'b0000001111111;
											assign node1420 = (inp[6]) ? 13'b0000000011111 : 13'b0000000111111;
										assign node1423 = (inp[5]) ? node1427 : node1424;
											assign node1424 = (inp[11]) ? 13'b0000000011111 : 13'b0000000111111;
											assign node1427 = (inp[2]) ? 13'b0000000001111 : 13'b0000000011111;
								assign node1430 = (inp[2]) ? node1446 : node1431;
									assign node1431 = (inp[11]) ? node1439 : node1432;
										assign node1432 = (inp[5]) ? node1436 : node1433;
											assign node1433 = (inp[6]) ? 13'b0000000111111 : 13'b0000011111111;
											assign node1436 = (inp[6]) ? 13'b0000000011111 : 13'b0000000111111;
										assign node1439 = (inp[1]) ? node1443 : node1440;
											assign node1440 = (inp[6]) ? 13'b0000000011111 : 13'b0000000111111;
											assign node1443 = (inp[5]) ? 13'b0000000000111 : 13'b0000000011111;
									assign node1446 = (inp[11]) ? node1454 : node1447;
										assign node1447 = (inp[6]) ? node1451 : node1448;
											assign node1448 = (inp[5]) ? 13'b0000000011111 : 13'b0000000111111;
											assign node1451 = (inp[1]) ? 13'b0000000001111 : 13'b0000000001111;
										assign node1454 = (inp[1]) ? node1458 : node1455;
											assign node1455 = (inp[5]) ? 13'b0000000001111 : 13'b0000000001111;
											assign node1458 = (inp[3]) ? 13'b0000000000111 : 13'b0000000000111;
				assign node1461 = (inp[11]) ? node1709 : node1462;
					assign node1462 = (inp[5]) ? node1584 : node1463;
						assign node1463 = (inp[6]) ? node1521 : node1464;
							assign node1464 = (inp[7]) ? node1494 : node1465;
								assign node1465 = (inp[10]) ? node1479 : node1466;
									assign node1466 = (inp[8]) ? node1472 : node1467;
										assign node1467 = (inp[0]) ? 13'b0000111111111 : node1468;
											assign node1468 = (inp[3]) ? 13'b0000111111111 : 13'b0001111111111;
										assign node1472 = (inp[2]) ? node1476 : node1473;
											assign node1473 = (inp[1]) ? 13'b0000011111111 : 13'b0000111111111;
											assign node1476 = (inp[3]) ? 13'b0000001111111 : 13'b0000011111111;
									assign node1479 = (inp[2]) ? node1487 : node1480;
										assign node1480 = (inp[8]) ? node1484 : node1481;
											assign node1481 = (inp[1]) ? 13'b0000111111111 : 13'b0001111111111;
											assign node1484 = (inp[1]) ? 13'b0000001111111 : 13'b0000011111111;
										assign node1487 = (inp[1]) ? node1491 : node1488;
											assign node1488 = (inp[8]) ? 13'b0000001111111 : 13'b0000011111111;
											assign node1491 = (inp[0]) ? 13'b0000000111111 : 13'b0000001111111;
								assign node1494 = (inp[0]) ? node1508 : node1495;
									assign node1495 = (inp[8]) ? node1503 : node1496;
										assign node1496 = (inp[1]) ? node1500 : node1497;
											assign node1497 = (inp[10]) ? 13'b0000011111111 : 13'b0000111111111;
											assign node1500 = (inp[2]) ? 13'b0000001111111 : 13'b0000011111111;
										assign node1503 = (inp[10]) ? 13'b0000001111111 : node1504;
											assign node1504 = (inp[3]) ? 13'b0000001111111 : 13'b0000011111111;
									assign node1508 = (inp[2]) ? node1514 : node1509;
										assign node1509 = (inp[10]) ? 13'b0000001111111 : node1510;
											assign node1510 = (inp[8]) ? 13'b0000001111111 : 13'b0000111111111;
										assign node1514 = (inp[8]) ? node1518 : node1515;
											assign node1515 = (inp[10]) ? 13'b0000000111111 : 13'b0000000111111;
											assign node1518 = (inp[10]) ? 13'b0000000001111 : 13'b0000000111111;
							assign node1521 = (inp[1]) ? node1553 : node1522;
								assign node1522 = (inp[8]) ? node1538 : node1523;
									assign node1523 = (inp[3]) ? node1531 : node1524;
										assign node1524 = (inp[10]) ? node1528 : node1525;
											assign node1525 = (inp[7]) ? 13'b0000011111111 : 13'b0000111111111;
											assign node1528 = (inp[0]) ? 13'b0000001111111 : 13'b0000011111111;
										assign node1531 = (inp[0]) ? node1535 : node1532;
											assign node1532 = (inp[10]) ? 13'b0000001111111 : 13'b0000011111111;
											assign node1535 = (inp[7]) ? 13'b0000000111111 : 13'b0000001111111;
									assign node1538 = (inp[10]) ? node1546 : node1539;
										assign node1539 = (inp[3]) ? node1543 : node1540;
											assign node1540 = (inp[2]) ? 13'b0000001111111 : 13'b0000011111111;
											assign node1543 = (inp[7]) ? 13'b0000000111111 : 13'b0000001111111;
										assign node1546 = (inp[7]) ? node1550 : node1547;
											assign node1547 = (inp[0]) ? 13'b0000000111111 : 13'b0000011111111;
											assign node1550 = (inp[3]) ? 13'b0000000011111 : 13'b0000000111111;
								assign node1553 = (inp[2]) ? node1569 : node1554;
									assign node1554 = (inp[7]) ? node1562 : node1555;
										assign node1555 = (inp[0]) ? node1559 : node1556;
											assign node1556 = (inp[8]) ? 13'b0000001111111 : 13'b0000011111111;
											assign node1559 = (inp[10]) ? 13'b0000000011111 : 13'b0000001111111;
										assign node1562 = (inp[10]) ? node1566 : node1563;
											assign node1563 = (inp[3]) ? 13'b0000000111111 : 13'b0000001111111;
											assign node1566 = (inp[0]) ? 13'b0000000011111 : 13'b0000000111111;
									assign node1569 = (inp[7]) ? node1577 : node1570;
										assign node1570 = (inp[8]) ? node1574 : node1571;
											assign node1571 = (inp[0]) ? 13'b0000000111111 : 13'b0000001111111;
											assign node1574 = (inp[0]) ? 13'b0000000011111 : 13'b0000000011111;
										assign node1577 = (inp[3]) ? node1581 : node1578;
											assign node1578 = (inp[0]) ? 13'b0000000011111 : 13'b0000000111111;
											assign node1581 = (inp[8]) ? 13'b0000000000111 : 13'b0000000011111;
						assign node1584 = (inp[1]) ? node1648 : node1585;
							assign node1585 = (inp[8]) ? node1617 : node1586;
								assign node1586 = (inp[2]) ? node1602 : node1587;
									assign node1587 = (inp[6]) ? node1595 : node1588;
										assign node1588 = (inp[3]) ? node1592 : node1589;
											assign node1589 = (inp[10]) ? 13'b0000011111111 : 13'b0000111111111;
											assign node1592 = (inp[10]) ? 13'b0000001111111 : 13'b0000011111111;
										assign node1595 = (inp[7]) ? node1599 : node1596;
											assign node1596 = (inp[3]) ? 13'b0000001111111 : 13'b0000011111111;
											assign node1599 = (inp[10]) ? 13'b0000001111111 : 13'b0000000111111;
									assign node1602 = (inp[7]) ? node1610 : node1603;
										assign node1603 = (inp[3]) ? node1607 : node1604;
											assign node1604 = (inp[6]) ? 13'b0000011111111 : 13'b0000011111111;
											assign node1607 = (inp[0]) ? 13'b0000000111111 : 13'b0000001111111;
										assign node1610 = (inp[0]) ? node1614 : node1611;
											assign node1611 = (inp[6]) ? 13'b0000000011111 : 13'b0000001111111;
											assign node1614 = (inp[10]) ? 13'b0000000011111 : 13'b0000000111111;
								assign node1617 = (inp[7]) ? node1633 : node1618;
									assign node1618 = (inp[2]) ? node1626 : node1619;
										assign node1619 = (inp[3]) ? node1623 : node1620;
											assign node1620 = (inp[6]) ? 13'b0000001111111 : 13'b0000111111111;
											assign node1623 = (inp[0]) ? 13'b0000000111111 : 13'b0000001111111;
										assign node1626 = (inp[0]) ? node1630 : node1627;
											assign node1627 = (inp[6]) ? 13'b0000000111111 : 13'b0000000111111;
											assign node1630 = (inp[6]) ? 13'b0000000011111 : 13'b0000000111111;
									assign node1633 = (inp[3]) ? node1641 : node1634;
										assign node1634 = (inp[0]) ? node1638 : node1635;
											assign node1635 = (inp[6]) ? 13'b0000000111111 : 13'b0000001111111;
											assign node1638 = (inp[2]) ? 13'b0000000001111 : 13'b0000000111111;
										assign node1641 = (inp[10]) ? node1645 : node1642;
											assign node1642 = (inp[0]) ? 13'b0000000011111 : 13'b0000000111111;
											assign node1645 = (inp[0]) ? 13'b0000000000111 : 13'b0000000011111;
							assign node1648 = (inp[0]) ? node1678 : node1649;
								assign node1649 = (inp[10]) ? node1663 : node1650;
									assign node1650 = (inp[6]) ? node1656 : node1651;
										assign node1651 = (inp[8]) ? node1653 : 13'b0000001111111;
											assign node1653 = (inp[2]) ? 13'b0000000111111 : 13'b0000001111111;
										assign node1656 = (inp[7]) ? node1660 : node1657;
											assign node1657 = (inp[3]) ? 13'b0000000111111 : 13'b0000001111111;
											assign node1660 = (inp[2]) ? 13'b0000000011111 : 13'b0000000111111;
									assign node1663 = (inp[6]) ? node1671 : node1664;
										assign node1664 = (inp[3]) ? node1668 : node1665;
											assign node1665 = (inp[2]) ? 13'b0000000111111 : 13'b0000001111111;
											assign node1668 = (inp[8]) ? 13'b0000000011111 : 13'b0000000111111;
										assign node1671 = (inp[7]) ? node1675 : node1672;
											assign node1672 = (inp[3]) ? 13'b0000000011111 : 13'b0000000111111;
											assign node1675 = (inp[2]) ? 13'b0000000001111 : 13'b0000000011111;
								assign node1678 = (inp[7]) ? node1694 : node1679;
									assign node1679 = (inp[2]) ? node1687 : node1680;
										assign node1680 = (inp[3]) ? node1684 : node1681;
											assign node1681 = (inp[6]) ? 13'b0000000111111 : 13'b0000000111111;
											assign node1684 = (inp[6]) ? 13'b0000000011111 : 13'b0000000111111;
										assign node1687 = (inp[6]) ? node1691 : node1688;
											assign node1688 = (inp[8]) ? 13'b0000000011111 : 13'b0000000111111;
											assign node1691 = (inp[8]) ? 13'b0000000001111 : 13'b0000000011111;
									assign node1694 = (inp[2]) ? node1702 : node1695;
										assign node1695 = (inp[6]) ? node1699 : node1696;
											assign node1696 = (inp[8]) ? 13'b0000000011111 : 13'b0000001111111;
											assign node1699 = (inp[8]) ? 13'b0000000001111 : 13'b0000000011111;
										assign node1702 = (inp[10]) ? node1706 : node1703;
											assign node1703 = (inp[3]) ? 13'b0000000001111 : 13'b0000000011111;
											assign node1706 = (inp[8]) ? 13'b0000000000111 : 13'b0000000001111;
					assign node1709 = (inp[5]) ? node1831 : node1710;
						assign node1710 = (inp[3]) ? node1770 : node1711;
							assign node1711 = (inp[0]) ? node1741 : node1712;
								assign node1712 = (inp[7]) ? node1726 : node1713;
									assign node1713 = (inp[8]) ? node1721 : node1714;
										assign node1714 = (inp[10]) ? node1718 : node1715;
											assign node1715 = (inp[1]) ? 13'b0000111111111 : 13'b0000111111111;
											assign node1718 = (inp[6]) ? 13'b0000011111111 : 13'b0000011111111;
										assign node1721 = (inp[6]) ? 13'b0000000111111 : node1722;
											assign node1722 = (inp[2]) ? 13'b0000001111111 : 13'b0000011111111;
									assign node1726 = (inp[1]) ? node1734 : node1727;
										assign node1727 = (inp[10]) ? node1731 : node1728;
											assign node1728 = (inp[2]) ? 13'b0000001111111 : 13'b0000011111111;
											assign node1731 = (inp[2]) ? 13'b0000000111111 : 13'b0000001111111;
										assign node1734 = (inp[6]) ? node1738 : node1735;
											assign node1735 = (inp[10]) ? 13'b0000000111111 : 13'b0000000111111;
											assign node1738 = (inp[2]) ? 13'b0000000011111 : 13'b0000000111111;
								assign node1741 = (inp[2]) ? node1757 : node1742;
									assign node1742 = (inp[10]) ? node1750 : node1743;
										assign node1743 = (inp[7]) ? node1747 : node1744;
											assign node1744 = (inp[1]) ? 13'b0000001111111 : 13'b0000011111111;
											assign node1747 = (inp[8]) ? 13'b0000000111111 : 13'b0000001111111;
										assign node1750 = (inp[1]) ? node1754 : node1751;
											assign node1751 = (inp[8]) ? 13'b0000000111111 : 13'b0000001111111;
											assign node1754 = (inp[7]) ? 13'b0000000011111 : 13'b0000000111111;
									assign node1757 = (inp[8]) ? node1763 : node1758;
										assign node1758 = (inp[10]) ? node1760 : 13'b0000001111111;
											assign node1760 = (inp[1]) ? 13'b0000000011111 : 13'b0000000111111;
										assign node1763 = (inp[6]) ? node1767 : node1764;
											assign node1764 = (inp[10]) ? 13'b0000000011111 : 13'b0000000111111;
											assign node1767 = (inp[1]) ? 13'b0000000000111 : 13'b0000000011111;
							assign node1770 = (inp[7]) ? node1800 : node1771;
								assign node1771 = (inp[2]) ? node1785 : node1772;
									assign node1772 = (inp[1]) ? node1778 : node1773;
										assign node1773 = (inp[0]) ? node1775 : 13'b0000011111111;
											assign node1775 = (inp[6]) ? 13'b0000000111111 : 13'b0000001111111;
										assign node1778 = (inp[8]) ? node1782 : node1779;
											assign node1779 = (inp[10]) ? 13'b0000000111111 : 13'b0000001111111;
											assign node1782 = (inp[0]) ? 13'b0000000011111 : 13'b0000000111111;
									assign node1785 = (inp[1]) ? node1793 : node1786;
										assign node1786 = (inp[6]) ? node1790 : node1787;
											assign node1787 = (inp[10]) ? 13'b0000000111111 : 13'b0000000111111;
											assign node1790 = (inp[0]) ? 13'b0000000011111 : 13'b0000001111111;
										assign node1793 = (inp[0]) ? node1797 : node1794;
											assign node1794 = (inp[6]) ? 13'b0000000001111 : 13'b0000000111111;
											assign node1797 = (inp[8]) ? 13'b0000000000111 : 13'b0000000011111;
								assign node1800 = (inp[10]) ? node1816 : node1801;
									assign node1801 = (inp[6]) ? node1809 : node1802;
										assign node1802 = (inp[0]) ? node1806 : node1803;
											assign node1803 = (inp[1]) ? 13'b0000000111111 : 13'b0000000111111;
											assign node1806 = (inp[8]) ? 13'b0000000011111 : 13'b0000000111111;
										assign node1809 = (inp[8]) ? node1813 : node1810;
											assign node1810 = (inp[0]) ? 13'b0000000011111 : 13'b0000000111111;
											assign node1813 = (inp[2]) ? 13'b0000000001111 : 13'b0000000001111;
									assign node1816 = (inp[0]) ? node1824 : node1817;
										assign node1817 = (inp[8]) ? node1821 : node1818;
											assign node1818 = (inp[6]) ? 13'b0000000011111 : 13'b0000000111111;
											assign node1821 = (inp[6]) ? 13'b0000000000111 : 13'b0000000011111;
										assign node1824 = (inp[2]) ? node1828 : node1825;
											assign node1825 = (inp[6]) ? 13'b0000000001111 : 13'b0000000001111;
											assign node1828 = (inp[8]) ? 13'b0000000000111 : 13'b0000000001111;
						assign node1831 = (inp[1]) ? node1891 : node1832;
							assign node1832 = (inp[10]) ? node1860 : node1833;
								assign node1833 = (inp[6]) ? node1845 : node1834;
									assign node1834 = (inp[8]) ? node1838 : node1835;
										assign node1835 = (inp[7]) ? 13'b0000001111111 : 13'b0000011111111;
										assign node1838 = (inp[3]) ? node1842 : node1839;
											assign node1839 = (inp[0]) ? 13'b0000000111111 : 13'b0000001111111;
											assign node1842 = (inp[0]) ? 13'b0000000011111 : 13'b0000000111111;
									assign node1845 = (inp[8]) ? node1853 : node1846;
										assign node1846 = (inp[0]) ? node1850 : node1847;
											assign node1847 = (inp[7]) ? 13'b0000000111111 : 13'b0000011111111;
											assign node1850 = (inp[3]) ? 13'b0000000011111 : 13'b0000000111111;
										assign node1853 = (inp[0]) ? node1857 : node1854;
											assign node1854 = (inp[7]) ? 13'b0000000011111 : 13'b0000000111111;
											assign node1857 = (inp[3]) ? 13'b0000000000111 : 13'b0000000011111;
								assign node1860 = (inp[6]) ? node1876 : node1861;
									assign node1861 = (inp[0]) ? node1869 : node1862;
										assign node1862 = (inp[7]) ? node1866 : node1863;
											assign node1863 = (inp[2]) ? 13'b0000000111111 : 13'b0000001111111;
											assign node1866 = (inp[3]) ? 13'b0000000011111 : 13'b0000000011111;
										assign node1869 = (inp[3]) ? node1873 : node1870;
											assign node1870 = (inp[8]) ? 13'b0000000011111 : 13'b0000000011111;
											assign node1873 = (inp[2]) ? 13'b0000000011111 : 13'b0000000001111;
									assign node1876 = (inp[2]) ? node1884 : node1877;
										assign node1877 = (inp[7]) ? node1881 : node1878;
											assign node1878 = (inp[0]) ? 13'b0000000011111 : 13'b0000000111111;
											assign node1881 = (inp[8]) ? 13'b0000000001111 : 13'b0000000011111;
										assign node1884 = (inp[8]) ? node1888 : node1885;
											assign node1885 = (inp[0]) ? 13'b0000000001111 : 13'b0000000011111;
											assign node1888 = (inp[0]) ? 13'b0000000000111 : 13'b0000000000111;
							assign node1891 = (inp[0]) ? node1923 : node1892;
								assign node1892 = (inp[7]) ? node1908 : node1893;
									assign node1893 = (inp[2]) ? node1901 : node1894;
										assign node1894 = (inp[8]) ? node1898 : node1895;
											assign node1895 = (inp[3]) ? 13'b0000000111111 : 13'b0000001111111;
											assign node1898 = (inp[3]) ? 13'b0000000001111 : 13'b0000000111111;
										assign node1901 = (inp[3]) ? node1905 : node1902;
											assign node1902 = (inp[6]) ? 13'b0000000011111 : 13'b0000000011111;
											assign node1905 = (inp[10]) ? 13'b0000000001111 : 13'b0000000011111;
									assign node1908 = (inp[6]) ? node1916 : node1909;
										assign node1909 = (inp[8]) ? node1913 : node1910;
											assign node1910 = (inp[3]) ? 13'b0000000011111 : 13'b0000000111111;
											assign node1913 = (inp[2]) ? 13'b0000000001111 : 13'b0000000011111;
										assign node1916 = (inp[3]) ? node1920 : node1917;
											assign node1917 = (inp[8]) ? 13'b0000000001111 : 13'b0000000011111;
											assign node1920 = (inp[2]) ? 13'b0000000000111 : 13'b0000000001111;
								assign node1923 = (inp[10]) ? node1937 : node1924;
									assign node1924 = (inp[8]) ? node1932 : node1925;
										assign node1925 = (inp[2]) ? node1929 : node1926;
											assign node1926 = (inp[6]) ? 13'b0000000011111 : 13'b0000000111111;
											assign node1929 = (inp[7]) ? 13'b0000000001111 : 13'b0000000011111;
										assign node1932 = (inp[7]) ? node1934 : 13'b0000000001111;
											assign node1934 = (inp[3]) ? 13'b0000000000111 : 13'b0000000000111;
									assign node1937 = (inp[2]) ? node1945 : node1938;
										assign node1938 = (inp[7]) ? node1942 : node1939;
											assign node1939 = (inp[6]) ? 13'b0000000001111 : 13'b0000000011111;
											assign node1942 = (inp[6]) ? 13'b0000000000111 : 13'b0000000001111;
										assign node1945 = (inp[7]) ? node1949 : node1946;
											assign node1946 = (inp[6]) ? 13'b0000000000111 : 13'b0000000000111;
											assign node1949 = (inp[3]) ? 13'b0000000000011 : 13'b0000000000111;
		assign node1952 = (inp[8]) ? node2922 : node1953;
			assign node1953 = (inp[2]) ? node2441 : node1954;
				assign node1954 = (inp[3]) ? node2198 : node1955;
					assign node1955 = (inp[0]) ? node2075 : node1956;
						assign node1956 = (inp[9]) ? node2016 : node1957;
							assign node1957 = (inp[5]) ? node1989 : node1958;
								assign node1958 = (inp[4]) ? node1974 : node1959;
									assign node1959 = (inp[11]) ? node1967 : node1960;
										assign node1960 = (inp[10]) ? node1964 : node1961;
											assign node1961 = (inp[6]) ? 13'b0001111111111 : 13'b0011111111111;
											assign node1964 = (inp[1]) ? 13'b0000111111111 : 13'b0001111111111;
										assign node1967 = (inp[10]) ? node1971 : node1968;
											assign node1968 = (inp[7]) ? 13'b0000111111111 : 13'b0001111111111;
											assign node1971 = (inp[1]) ? 13'b0000001111111 : 13'b0000111111111;
									assign node1974 = (inp[10]) ? node1982 : node1975;
										assign node1975 = (inp[7]) ? node1979 : node1976;
											assign node1976 = (inp[6]) ? 13'b0000111111111 : 13'b0001111111111;
											assign node1979 = (inp[1]) ? 13'b0000011111111 : 13'b0000111111111;
										assign node1982 = (inp[11]) ? node1986 : node1983;
											assign node1983 = (inp[1]) ? 13'b0000011111111 : 13'b0000111111111;
											assign node1986 = (inp[7]) ? 13'b0000001111111 : 13'b0000011111111;
								assign node1989 = (inp[4]) ? node2003 : node1990;
									assign node1990 = (inp[11]) ? node1996 : node1991;
										assign node1991 = (inp[7]) ? node1993 : 13'b0000111111111;
											assign node1993 = (inp[10]) ? 13'b0000011111111 : 13'b0000111111111;
										assign node1996 = (inp[6]) ? node2000 : node1997;
											assign node1997 = (inp[7]) ? 13'b0000011111111 : 13'b0000111111111;
											assign node2000 = (inp[1]) ? 13'b0000001111111 : 13'b0000011111111;
									assign node2003 = (inp[1]) ? node2011 : node2004;
										assign node2004 = (inp[6]) ? node2008 : node2005;
											assign node2005 = (inp[10]) ? 13'b0000111111111 : 13'b0001111111111;
											assign node2008 = (inp[10]) ? 13'b0000000111111 : 13'b0000011111111;
										assign node2011 = (inp[7]) ? node2013 : 13'b0000001111111;
											assign node2013 = (inp[11]) ? 13'b0000000111111 : 13'b0000001111111;
							assign node2016 = (inp[1]) ? node2048 : node2017;
								assign node2017 = (inp[4]) ? node2033 : node2018;
									assign node2018 = (inp[5]) ? node2026 : node2019;
										assign node2019 = (inp[10]) ? node2023 : node2020;
											assign node2020 = (inp[6]) ? 13'b0000111111111 : 13'b0001111111111;
											assign node2023 = (inp[7]) ? 13'b0000011111111 : 13'b0000111111111;
										assign node2026 = (inp[7]) ? node2030 : node2027;
											assign node2027 = (inp[10]) ? 13'b0000011111111 : 13'b0000011111111;
											assign node2030 = (inp[11]) ? 13'b0000001111111 : 13'b0000011111111;
									assign node2033 = (inp[5]) ? node2041 : node2034;
										assign node2034 = (inp[10]) ? node2038 : node2035;
											assign node2035 = (inp[6]) ? 13'b0000011111111 : 13'b0000111111111;
											assign node2038 = (inp[6]) ? 13'b0000001111111 : 13'b0000011111111;
										assign node2041 = (inp[11]) ? node2045 : node2042;
											assign node2042 = (inp[6]) ? 13'b0000001111111 : 13'b0000011111111;
											assign node2045 = (inp[7]) ? 13'b0000000111111 : 13'b0000001111111;
								assign node2048 = (inp[5]) ? node2064 : node2049;
									assign node2049 = (inp[10]) ? node2057 : node2050;
										assign node2050 = (inp[6]) ? node2054 : node2051;
											assign node2051 = (inp[4]) ? 13'b0000011111111 : 13'b0000111111111;
											assign node2054 = (inp[11]) ? 13'b0000000111111 : 13'b0000011111111;
										assign node2057 = (inp[7]) ? node2061 : node2058;
											assign node2058 = (inp[4]) ? 13'b0000001111111 : 13'b0000001111111;
											assign node2061 = (inp[11]) ? 13'b0000000111111 : 13'b0000001111111;
									assign node2064 = (inp[10]) ? node2070 : node2065;
										assign node2065 = (inp[7]) ? node2067 : 13'b0000001111111;
											assign node2067 = (inp[11]) ? 13'b0000000011111 : 13'b0000001111111;
										assign node2070 = (inp[4]) ? node2072 : 13'b0000000111111;
											assign node2072 = (inp[7]) ? 13'b0000000001111 : 13'b0000000011111;
						assign node2075 = (inp[7]) ? node2137 : node2076;
							assign node2076 = (inp[5]) ? node2106 : node2077;
								assign node2077 = (inp[10]) ? node2093 : node2078;
									assign node2078 = (inp[4]) ? node2086 : node2079;
										assign node2079 = (inp[1]) ? node2083 : node2080;
											assign node2080 = (inp[11]) ? 13'b0000111111111 : 13'b0001111111111;
											assign node2083 = (inp[6]) ? 13'b0000001111111 : 13'b0000111111111;
										assign node2086 = (inp[11]) ? node2090 : node2087;
											assign node2087 = (inp[6]) ? 13'b0000011111111 : 13'b0000111111111;
											assign node2090 = (inp[6]) ? 13'b0000001111111 : 13'b0000011111111;
									assign node2093 = (inp[11]) ? node2099 : node2094;
										assign node2094 = (inp[1]) ? node2096 : 13'b0000011111111;
											assign node2096 = (inp[6]) ? 13'b0000001111111 : 13'b0000011111111;
										assign node2099 = (inp[4]) ? node2103 : node2100;
											assign node2100 = (inp[1]) ? 13'b0000001111111 : 13'b0000001111111;
											assign node2103 = (inp[1]) ? 13'b0000000111111 : 13'b0000001111111;
								assign node2106 = (inp[6]) ? node2122 : node2107;
									assign node2107 = (inp[9]) ? node2115 : node2108;
										assign node2108 = (inp[4]) ? node2112 : node2109;
											assign node2109 = (inp[1]) ? 13'b0000011111111 : 13'b0000111111111;
											assign node2112 = (inp[10]) ? 13'b0000001111111 : 13'b0000011111111;
										assign node2115 = (inp[1]) ? node2119 : node2116;
											assign node2116 = (inp[4]) ? 13'b0000001111111 : 13'b0000011111111;
											assign node2119 = (inp[10]) ? 13'b0000000111111 : 13'b0000001111111;
									assign node2122 = (inp[4]) ? node2130 : node2123;
										assign node2123 = (inp[11]) ? node2127 : node2124;
											assign node2124 = (inp[10]) ? 13'b0000001111111 : 13'b0000001111111;
											assign node2127 = (inp[1]) ? 13'b0000000111111 : 13'b0000001111111;
										assign node2130 = (inp[1]) ? node2134 : node2131;
											assign node2131 = (inp[10]) ? 13'b0000000111111 : 13'b0000001111111;
											assign node2134 = (inp[11]) ? 13'b0000000011111 : 13'b0000000111111;
							assign node2137 = (inp[1]) ? node2169 : node2138;
								assign node2138 = (inp[6]) ? node2154 : node2139;
									assign node2139 = (inp[11]) ? node2147 : node2140;
										assign node2140 = (inp[10]) ? node2144 : node2141;
											assign node2141 = (inp[9]) ? 13'b0000011111111 : 13'b0000111111111;
											assign node2144 = (inp[5]) ? 13'b0000001111111 : 13'b0000011111111;
										assign node2147 = (inp[4]) ? node2151 : node2148;
											assign node2148 = (inp[10]) ? 13'b0000001111111 : 13'b0000011111111;
											assign node2151 = (inp[10]) ? 13'b0000000111111 : 13'b0000001111111;
									assign node2154 = (inp[10]) ? node2162 : node2155;
										assign node2155 = (inp[4]) ? node2159 : node2156;
											assign node2156 = (inp[11]) ? 13'b0000001111111 : 13'b0000011111111;
											assign node2159 = (inp[11]) ? 13'b0000000111111 : 13'b0000001111111;
										assign node2162 = (inp[5]) ? node2166 : node2163;
											assign node2163 = (inp[4]) ? 13'b0000000111111 : 13'b0000001111111;
											assign node2166 = (inp[11]) ? 13'b0000000011111 : 13'b0000000111111;
								assign node2169 = (inp[4]) ? node2185 : node2170;
									assign node2170 = (inp[5]) ? node2178 : node2171;
										assign node2171 = (inp[6]) ? node2175 : node2172;
											assign node2172 = (inp[9]) ? 13'b0000001111111 : 13'b0000011111111;
											assign node2175 = (inp[9]) ? 13'b0000000111111 : 13'b0000001111111;
										assign node2178 = (inp[11]) ? node2182 : node2179;
											assign node2179 = (inp[10]) ? 13'b0000000111111 : 13'b0000001111111;
											assign node2182 = (inp[9]) ? 13'b0000000011111 : 13'b0000000011111;
									assign node2185 = (inp[6]) ? node2193 : node2186;
										assign node2186 = (inp[10]) ? node2190 : node2187;
											assign node2187 = (inp[9]) ? 13'b0000000011111 : 13'b0000001111111;
											assign node2190 = (inp[11]) ? 13'b0000000011111 : 13'b0000000111111;
										assign node2193 = (inp[11]) ? node2195 : 13'b0000000011111;
											assign node2195 = (inp[5]) ? 13'b0000000001111 : 13'b0000000011111;
					assign node2198 = (inp[6]) ? node2320 : node2199;
						assign node2199 = (inp[4]) ? node2259 : node2200;
							assign node2200 = (inp[9]) ? node2232 : node2201;
								assign node2201 = (inp[5]) ? node2217 : node2202;
									assign node2202 = (inp[11]) ? node2210 : node2203;
										assign node2203 = (inp[10]) ? node2207 : node2204;
											assign node2204 = (inp[7]) ? 13'b0000111111111 : 13'b0001111111111;
											assign node2207 = (inp[0]) ? 13'b0000011111111 : 13'b0000111111111;
										assign node2210 = (inp[1]) ? node2214 : node2211;
											assign node2211 = (inp[0]) ? 13'b0000011111111 : 13'b0000111111111;
											assign node2214 = (inp[10]) ? 13'b0000001111111 : 13'b0000011111111;
									assign node2217 = (inp[0]) ? node2225 : node2218;
										assign node2218 = (inp[1]) ? node2222 : node2219;
											assign node2219 = (inp[7]) ? 13'b0000011111111 : 13'b0000111111111;
											assign node2222 = (inp[7]) ? 13'b0000001111111 : 13'b0000011111111;
										assign node2225 = (inp[10]) ? node2229 : node2226;
											assign node2226 = (inp[7]) ? 13'b0000001111111 : 13'b0000011111111;
											assign node2229 = (inp[11]) ? 13'b0000000111111 : 13'b0000001111111;
								assign node2232 = (inp[7]) ? node2244 : node2233;
									assign node2233 = (inp[0]) ? node2239 : node2234;
										assign node2234 = (inp[11]) ? 13'b0000011111111 : node2235;
											assign node2235 = (inp[1]) ? 13'b0000011111111 : 13'b0000111111111;
										assign node2239 = (inp[11]) ? 13'b0000001111111 : node2240;
											assign node2240 = (inp[5]) ? 13'b0000001111111 : 13'b0000011111111;
									assign node2244 = (inp[11]) ? node2252 : node2245;
										assign node2245 = (inp[10]) ? node2249 : node2246;
											assign node2246 = (inp[5]) ? 13'b0000001111111 : 13'b0000011111111;
											assign node2249 = (inp[0]) ? 13'b0000000111111 : 13'b0000011111111;
										assign node2252 = (inp[1]) ? node2256 : node2253;
											assign node2253 = (inp[10]) ? 13'b0000000111111 : 13'b0000000111111;
											assign node2256 = (inp[5]) ? 13'b0000000011111 : 13'b0000000111111;
							assign node2259 = (inp[1]) ? node2291 : node2260;
								assign node2260 = (inp[7]) ? node2276 : node2261;
									assign node2261 = (inp[11]) ? node2269 : node2262;
										assign node2262 = (inp[0]) ? node2266 : node2263;
											assign node2263 = (inp[10]) ? 13'b0000011111111 : 13'b0000111111111;
											assign node2266 = (inp[9]) ? 13'b0000001111111 : 13'b0000011111111;
										assign node2269 = (inp[0]) ? node2273 : node2270;
											assign node2270 = (inp[10]) ? 13'b0000001111111 : 13'b0000011111111;
											assign node2273 = (inp[10]) ? 13'b0000000011111 : 13'b0000001111111;
									assign node2276 = (inp[0]) ? node2284 : node2277;
										assign node2277 = (inp[9]) ? node2281 : node2278;
											assign node2278 = (inp[10]) ? 13'b0000001111111 : 13'b0000011111111;
											assign node2281 = (inp[11]) ? 13'b0000000111111 : 13'b0000001111111;
										assign node2284 = (inp[10]) ? node2288 : node2285;
											assign node2285 = (inp[11]) ? 13'b0000000111111 : 13'b0000001111111;
											assign node2288 = (inp[9]) ? 13'b0000000001111 : 13'b0000000111111;
								assign node2291 = (inp[5]) ? node2305 : node2292;
									assign node2292 = (inp[0]) ? node2298 : node2293;
										assign node2293 = (inp[9]) ? node2295 : 13'b0000001111111;
											assign node2295 = (inp[10]) ? 13'b0000000111111 : 13'b0000001111111;
										assign node2298 = (inp[9]) ? node2302 : node2299;
											assign node2299 = (inp[11]) ? 13'b0000000111111 : 13'b0000001111111;
											assign node2302 = (inp[7]) ? 13'b0000000001111 : 13'b0000000111111;
									assign node2305 = (inp[10]) ? node2313 : node2306;
										assign node2306 = (inp[7]) ? node2310 : node2307;
											assign node2307 = (inp[9]) ? 13'b0000000111111 : 13'b0000001111111;
											assign node2310 = (inp[11]) ? 13'b0000000011111 : 13'b0000000111111;
										assign node2313 = (inp[11]) ? node2317 : node2314;
											assign node2314 = (inp[9]) ? 13'b0000000011111 : 13'b0000000111111;
											assign node2317 = (inp[0]) ? 13'b0000000001111 : 13'b0000000011111;
						assign node2320 = (inp[0]) ? node2382 : node2321;
							assign node2321 = (inp[5]) ? node2353 : node2322;
								assign node2322 = (inp[4]) ? node2338 : node2323;
									assign node2323 = (inp[7]) ? node2331 : node2324;
										assign node2324 = (inp[10]) ? node2328 : node2325;
											assign node2325 = (inp[9]) ? 13'b0000011111111 : 13'b0000111111111;
											assign node2328 = (inp[11]) ? 13'b0000001111111 : 13'b0000011111111;
										assign node2331 = (inp[9]) ? node2335 : node2332;
											assign node2332 = (inp[1]) ? 13'b0000000111111 : 13'b0000011111111;
											assign node2335 = (inp[11]) ? 13'b0000000111111 : 13'b0000001111111;
									assign node2338 = (inp[10]) ? node2346 : node2339;
										assign node2339 = (inp[11]) ? node2343 : node2340;
											assign node2340 = (inp[9]) ? 13'b0000001111111 : 13'b0000011111111;
											assign node2343 = (inp[1]) ? 13'b0000000111111 : 13'b0000001111111;
										assign node2346 = (inp[11]) ? node2350 : node2347;
											assign node2347 = (inp[7]) ? 13'b0000000111111 : 13'b0000001111111;
											assign node2350 = (inp[7]) ? 13'b0000000001111 : 13'b0000000111111;
								assign node2353 = (inp[10]) ? node2369 : node2354;
									assign node2354 = (inp[11]) ? node2362 : node2355;
										assign node2355 = (inp[4]) ? node2359 : node2356;
											assign node2356 = (inp[9]) ? 13'b0000001111111 : 13'b0000011111111;
											assign node2359 = (inp[1]) ? 13'b0000000111111 : 13'b0000001111111;
										assign node2362 = (inp[7]) ? node2366 : node2363;
											assign node2363 = (inp[4]) ? 13'b0000000111111 : 13'b0000001111111;
											assign node2366 = (inp[4]) ? 13'b0000000011111 : 13'b0000000111111;
									assign node2369 = (inp[4]) ? node2377 : node2370;
										assign node2370 = (inp[11]) ? node2374 : node2371;
											assign node2371 = (inp[1]) ? 13'b0000000111111 : 13'b0000000111111;
											assign node2374 = (inp[1]) ? 13'b0000000011111 : 13'b0000000111111;
										assign node2377 = (inp[9]) ? 13'b0000000011111 : node2378;
											assign node2378 = (inp[11]) ? 13'b0000000011111 : 13'b0000000111111;
							assign node2382 = (inp[1]) ? node2412 : node2383;
								assign node2383 = (inp[11]) ? node2399 : node2384;
									assign node2384 = (inp[10]) ? node2392 : node2385;
										assign node2385 = (inp[7]) ? node2389 : node2386;
											assign node2386 = (inp[9]) ? 13'b0000001111111 : 13'b0000011111111;
											assign node2389 = (inp[4]) ? 13'b0000000111111 : 13'b0000001111111;
										assign node2392 = (inp[9]) ? node2396 : node2393;
											assign node2393 = (inp[5]) ? 13'b0000000111111 : 13'b0000001111111;
											assign node2396 = (inp[4]) ? 13'b0000000011111 : 13'b0000000111111;
									assign node2399 = (inp[7]) ? node2407 : node2400;
										assign node2400 = (inp[4]) ? node2404 : node2401;
											assign node2401 = (inp[9]) ? 13'b0000000111111 : 13'b0000001111111;
											assign node2404 = (inp[10]) ? 13'b0000000011111 : 13'b0000000111111;
										assign node2407 = (inp[10]) ? 13'b0000000011111 : node2408;
											assign node2408 = (inp[4]) ? 13'b0000000011111 : 13'b0000000111111;
								assign node2412 = (inp[11]) ? node2428 : node2413;
									assign node2413 = (inp[7]) ? node2421 : node2414;
										assign node2414 = (inp[9]) ? node2418 : node2415;
											assign node2415 = (inp[5]) ? 13'b0000000111111 : 13'b0000001111111;
											assign node2418 = (inp[4]) ? 13'b0000000011111 : 13'b0000000111111;
										assign node2421 = (inp[10]) ? node2425 : node2422;
											assign node2422 = (inp[4]) ? 13'b0000000011111 : 13'b0000000111111;
											assign node2425 = (inp[5]) ? 13'b0000000001111 : 13'b0000000011111;
									assign node2428 = (inp[10]) ? node2436 : node2429;
										assign node2429 = (inp[4]) ? node2433 : node2430;
											assign node2430 = (inp[9]) ? 13'b0000000011111 : 13'b0000000111111;
											assign node2433 = (inp[9]) ? 13'b0000000001111 : 13'b0000000011111;
										assign node2436 = (inp[7]) ? node2438 : 13'b0000000001111;
											assign node2438 = (inp[5]) ? 13'b0000000000011 : 13'b0000000000111;
				assign node2441 = (inp[0]) ? node2681 : node2442;
					assign node2442 = (inp[7]) ? node2564 : node2443;
						assign node2443 = (inp[5]) ? node2501 : node2444;
							assign node2444 = (inp[3]) ? node2472 : node2445;
								assign node2445 = (inp[9]) ? node2459 : node2446;
									assign node2446 = (inp[1]) ? node2454 : node2447;
										assign node2447 = (inp[6]) ? node2451 : node2448;
											assign node2448 = (inp[11]) ? 13'b0000111111111 : 13'b0001111111111;
											assign node2451 = (inp[10]) ? 13'b0000011111111 : 13'b0000111111111;
										assign node2454 = (inp[6]) ? 13'b0000001111111 : node2455;
											assign node2455 = (inp[4]) ? 13'b0000011111111 : 13'b0000111111111;
									assign node2459 = (inp[4]) ? node2467 : node2460;
										assign node2460 = (inp[10]) ? node2464 : node2461;
											assign node2461 = (inp[6]) ? 13'b0000011111111 : 13'b0000111111111;
											assign node2464 = (inp[11]) ? 13'b0000001111111 : 13'b0000001111111;
										assign node2467 = (inp[6]) ? 13'b0000001111111 : node2468;
											assign node2468 = (inp[1]) ? 13'b0000001111111 : 13'b0000001111111;
								assign node2472 = (inp[10]) ? node2486 : node2473;
									assign node2473 = (inp[1]) ? node2479 : node2474;
										assign node2474 = (inp[11]) ? 13'b0000011111111 : node2475;
											assign node2475 = (inp[4]) ? 13'b0000011111111 : 13'b0000111111111;
										assign node2479 = (inp[9]) ? node2483 : node2480;
											assign node2480 = (inp[11]) ? 13'b0000001111111 : 13'b0000011111111;
											assign node2483 = (inp[4]) ? 13'b0000000111111 : 13'b0000001111111;
									assign node2486 = (inp[4]) ? node2494 : node2487;
										assign node2487 = (inp[9]) ? node2491 : node2488;
											assign node2488 = (inp[11]) ? 13'b0000001111111 : 13'b0000001111111;
											assign node2491 = (inp[11]) ? 13'b0000000111111 : 13'b0000001111111;
										assign node2494 = (inp[11]) ? node2498 : node2495;
											assign node2495 = (inp[6]) ? 13'b0000000111111 : 13'b0000001111111;
											assign node2498 = (inp[1]) ? 13'b0000000001111 : 13'b0000000111111;
							assign node2501 = (inp[9]) ? node2533 : node2502;
								assign node2502 = (inp[6]) ? node2518 : node2503;
									assign node2503 = (inp[1]) ? node2511 : node2504;
										assign node2504 = (inp[3]) ? node2508 : node2505;
											assign node2505 = (inp[10]) ? 13'b0000011111111 : 13'b0000111111111;
											assign node2508 = (inp[4]) ? 13'b0000001111111 : 13'b0000011111111;
										assign node2511 = (inp[10]) ? node2515 : node2512;
											assign node2512 = (inp[3]) ? 13'b0000001111111 : 13'b0000011111111;
											assign node2515 = (inp[3]) ? 13'b0000000011111 : 13'b0000001111111;
									assign node2518 = (inp[3]) ? node2526 : node2519;
										assign node2519 = (inp[10]) ? node2523 : node2520;
											assign node2520 = (inp[4]) ? 13'b0000001111111 : 13'b0000011111111;
											assign node2523 = (inp[1]) ? 13'b0000000111111 : 13'b0000001111111;
										assign node2526 = (inp[4]) ? node2530 : node2527;
											assign node2527 = (inp[1]) ? 13'b0000000111111 : 13'b0000011111111;
											assign node2530 = (inp[1]) ? 13'b0000000011111 : 13'b0000000111111;
								assign node2533 = (inp[10]) ? node2549 : node2534;
									assign node2534 = (inp[4]) ? node2542 : node2535;
										assign node2535 = (inp[3]) ? node2539 : node2536;
											assign node2536 = (inp[6]) ? 13'b0000001111111 : 13'b0000111111111;
											assign node2539 = (inp[11]) ? 13'b0000000111111 : 13'b0000001111111;
										assign node2542 = (inp[6]) ? node2546 : node2543;
											assign node2543 = (inp[11]) ? 13'b0000000011111 : 13'b0000001111111;
											assign node2546 = (inp[3]) ? 13'b0000000011111 : 13'b0000000111111;
									assign node2549 = (inp[1]) ? node2557 : node2550;
										assign node2550 = (inp[3]) ? node2554 : node2551;
											assign node2551 = (inp[4]) ? 13'b0000000111111 : 13'b0000001111111;
											assign node2554 = (inp[6]) ? 13'b0000000011111 : 13'b0000000111111;
										assign node2557 = (inp[3]) ? node2561 : node2558;
											assign node2558 = (inp[4]) ? 13'b0000000011111 : 13'b0000000011111;
											assign node2561 = (inp[4]) ? 13'b0000000000111 : 13'b0000000011111;
						assign node2564 = (inp[3]) ? node2622 : node2565;
							assign node2565 = (inp[9]) ? node2593 : node2566;
								assign node2566 = (inp[6]) ? node2582 : node2567;
									assign node2567 = (inp[11]) ? node2575 : node2568;
										assign node2568 = (inp[1]) ? node2572 : node2569;
											assign node2569 = (inp[5]) ? 13'b0000011111111 : 13'b0000111111111;
											assign node2572 = (inp[4]) ? 13'b0000001111111 : 13'b0000011111111;
										assign node2575 = (inp[1]) ? node2579 : node2576;
											assign node2576 = (inp[5]) ? 13'b0000001111111 : 13'b0000011111111;
											assign node2579 = (inp[5]) ? 13'b0000000011111 : 13'b0000001111111;
									assign node2582 = (inp[10]) ? node2588 : node2583;
										assign node2583 = (inp[5]) ? node2585 : 13'b0000011111111;
											assign node2585 = (inp[4]) ? 13'b0000000111111 : 13'b0000001111111;
										assign node2588 = (inp[11]) ? 13'b0000000111111 : node2589;
											assign node2589 = (inp[1]) ? 13'b0000000111111 : 13'b0000001111111;
								assign node2593 = (inp[5]) ? node2607 : node2594;
									assign node2594 = (inp[6]) ? node2602 : node2595;
										assign node2595 = (inp[10]) ? node2599 : node2596;
											assign node2596 = (inp[4]) ? 13'b0000001111111 : 13'b0000011111111;
											assign node2599 = (inp[4]) ? 13'b0000000111111 : 13'b0000000111111;
										assign node2602 = (inp[11]) ? node2604 : 13'b0000000111111;
											assign node2604 = (inp[10]) ? 13'b0000000011111 : 13'b0000000111111;
									assign node2607 = (inp[4]) ? node2615 : node2608;
										assign node2608 = (inp[1]) ? node2612 : node2609;
											assign node2609 = (inp[11]) ? 13'b0000000111111 : 13'b0000000111111;
											assign node2612 = (inp[6]) ? 13'b0000000011111 : 13'b0000000111111;
										assign node2615 = (inp[1]) ? node2619 : node2616;
											assign node2616 = (inp[6]) ? 13'b0000000011111 : 13'b0000000111111;
											assign node2619 = (inp[10]) ? 13'b0000000000111 : 13'b0000000001111;
							assign node2622 = (inp[1]) ? node2652 : node2623;
								assign node2623 = (inp[5]) ? node2637 : node2624;
									assign node2624 = (inp[11]) ? node2630 : node2625;
										assign node2625 = (inp[4]) ? node2627 : 13'b0000001111111;
											assign node2627 = (inp[10]) ? 13'b0000000111111 : 13'b0000001111111;
										assign node2630 = (inp[6]) ? node2634 : node2631;
											assign node2631 = (inp[9]) ? 13'b0000000111111 : 13'b0000001111111;
											assign node2634 = (inp[10]) ? 13'b0000000001111 : 13'b0000000011111;
									assign node2637 = (inp[4]) ? node2645 : node2638;
										assign node2638 = (inp[11]) ? node2642 : node2639;
											assign node2639 = (inp[6]) ? 13'b0000000111111 : 13'b0000001111111;
											assign node2642 = (inp[10]) ? 13'b0000000011111 : 13'b0000000111111;
										assign node2645 = (inp[9]) ? node2649 : node2646;
											assign node2646 = (inp[11]) ? 13'b0000000011111 : 13'b0000000011111;
											assign node2649 = (inp[10]) ? 13'b0000000001111 : 13'b0000000011111;
								assign node2652 = (inp[10]) ? node2666 : node2653;
									assign node2653 = (inp[9]) ? node2659 : node2654;
										assign node2654 = (inp[4]) ? 13'b0000000011111 : node2655;
											assign node2655 = (inp[11]) ? 13'b0000000111111 : 13'b0000001111111;
										assign node2659 = (inp[6]) ? node2663 : node2660;
											assign node2660 = (inp[5]) ? 13'b0000000011111 : 13'b0000000111111;
											assign node2663 = (inp[11]) ? 13'b0000000001111 : 13'b0000000011111;
									assign node2666 = (inp[9]) ? node2674 : node2667;
										assign node2667 = (inp[4]) ? node2671 : node2668;
											assign node2668 = (inp[6]) ? 13'b0000000011111 : 13'b0000000011111;
											assign node2671 = (inp[6]) ? 13'b0000000001111 : 13'b0000000011111;
										assign node2674 = (inp[11]) ? node2678 : node2675;
											assign node2675 = (inp[4]) ? 13'b0000000001111 : 13'b0000000011111;
											assign node2678 = (inp[5]) ? 13'b0000000000111 : 13'b0000000001111;
					assign node2681 = (inp[4]) ? node2803 : node2682;
						assign node2682 = (inp[9]) ? node2746 : node2683;
							assign node2683 = (inp[5]) ? node2715 : node2684;
								assign node2684 = (inp[1]) ? node2700 : node2685;
									assign node2685 = (inp[7]) ? node2693 : node2686;
										assign node2686 = (inp[10]) ? node2690 : node2687;
											assign node2687 = (inp[6]) ? 13'b0000011111111 : 13'b0000111111111;
											assign node2690 = (inp[3]) ? 13'b0000001111111 : 13'b0000011111111;
										assign node2693 = (inp[6]) ? node2697 : node2694;
											assign node2694 = (inp[11]) ? 13'b0000001111111 : 13'b0000011111111;
											assign node2697 = (inp[3]) ? 13'b0000000111111 : 13'b0000001111111;
									assign node2700 = (inp[11]) ? node2708 : node2701;
										assign node2701 = (inp[3]) ? node2705 : node2702;
											assign node2702 = (inp[7]) ? 13'b0000001111111 : 13'b0000011111111;
											assign node2705 = (inp[6]) ? 13'b0000000111111 : 13'b0000001111111;
										assign node2708 = (inp[7]) ? node2712 : node2709;
											assign node2709 = (inp[3]) ? 13'b0000000011111 : 13'b0000001111111;
											assign node2712 = (inp[6]) ? 13'b0000000011111 : 13'b0000000111111;
								assign node2715 = (inp[10]) ? node2731 : node2716;
									assign node2716 = (inp[7]) ? node2724 : node2717;
										assign node2717 = (inp[1]) ? node2721 : node2718;
											assign node2718 = (inp[6]) ? 13'b0000001111111 : 13'b0000011111111;
											assign node2721 = (inp[6]) ? 13'b0000000111111 : 13'b0000001111111;
										assign node2724 = (inp[6]) ? node2728 : node2725;
											assign node2725 = (inp[11]) ? 13'b0000000111111 : 13'b0000001111111;
											assign node2728 = (inp[11]) ? 13'b0000000011111 : 13'b0000000011111;
									assign node2731 = (inp[1]) ? node2739 : node2732;
										assign node2732 = (inp[6]) ? node2736 : node2733;
											assign node2733 = (inp[3]) ? 13'b0000000111111 : 13'b0000001111111;
											assign node2736 = (inp[3]) ? 13'b0000000011111 : 13'b0000000111111;
										assign node2739 = (inp[6]) ? node2743 : node2740;
											assign node2740 = (inp[11]) ? 13'b0000000011111 : 13'b0000000111111;
											assign node2743 = (inp[11]) ? 13'b0000000000111 : 13'b0000000011111;
							assign node2746 = (inp[6]) ? node2774 : node2747;
								assign node2747 = (inp[10]) ? node2761 : node2748;
									assign node2748 = (inp[11]) ? node2754 : node2749;
										assign node2749 = (inp[7]) ? node2751 : 13'b0000001111111;
											assign node2751 = (inp[1]) ? 13'b0000000111111 : 13'b0000001111111;
										assign node2754 = (inp[7]) ? node2758 : node2755;
											assign node2755 = (inp[1]) ? 13'b0000000111111 : 13'b0000001111111;
											assign node2758 = (inp[3]) ? 13'b0000000011111 : 13'b0000000011111;
									assign node2761 = (inp[5]) ? node2767 : node2762;
										assign node2762 = (inp[1]) ? node2764 : 13'b0000000111111;
											assign node2764 = (inp[7]) ? 13'b0000000011111 : 13'b0000000111111;
										assign node2767 = (inp[3]) ? node2771 : node2768;
											assign node2768 = (inp[7]) ? 13'b0000000011111 : 13'b0000000111111;
											assign node2771 = (inp[11]) ? 13'b0000000001111 : 13'b0000000011111;
								assign node2774 = (inp[5]) ? node2788 : node2775;
									assign node2775 = (inp[3]) ? node2781 : node2776;
										assign node2776 = (inp[1]) ? 13'b0000000111111 : node2777;
											assign node2777 = (inp[11]) ? 13'b0000000111111 : 13'b0000001111111;
										assign node2781 = (inp[7]) ? node2785 : node2782;
											assign node2782 = (inp[1]) ? 13'b0000000001111 : 13'b0000000111111;
											assign node2785 = (inp[1]) ? 13'b0000000001111 : 13'b0000000001111;
									assign node2788 = (inp[10]) ? node2796 : node2789;
										assign node2789 = (inp[11]) ? node2793 : node2790;
											assign node2790 = (inp[3]) ? 13'b0000000011111 : 13'b0000000011111;
											assign node2793 = (inp[1]) ? 13'b0000000001111 : 13'b0000000011111;
										assign node2796 = (inp[11]) ? node2800 : node2797;
											assign node2797 = (inp[7]) ? 13'b0000000001111 : 13'b0000000001111;
											assign node2800 = (inp[1]) ? 13'b0000000000111 : 13'b0000000001111;
						assign node2803 = (inp[11]) ? node2865 : node2804;
							assign node2804 = (inp[7]) ? node2836 : node2805;
								assign node2805 = (inp[9]) ? node2821 : node2806;
									assign node2806 = (inp[6]) ? node2814 : node2807;
										assign node2807 = (inp[3]) ? node2811 : node2808;
											assign node2808 = (inp[5]) ? 13'b0000001111111 : 13'b0000011111111;
											assign node2811 = (inp[1]) ? 13'b0000000111111 : 13'b0000001111111;
										assign node2814 = (inp[10]) ? node2818 : node2815;
											assign node2815 = (inp[1]) ? 13'b0000000111111 : 13'b0000000111111;
											assign node2818 = (inp[3]) ? 13'b0000000011111 : 13'b0000000111111;
									assign node2821 = (inp[5]) ? node2829 : node2822;
										assign node2822 = (inp[6]) ? node2826 : node2823;
											assign node2823 = (inp[3]) ? 13'b0000000111111 : 13'b0000001111111;
											assign node2826 = (inp[10]) ? 13'b0000000011111 : 13'b0000000111111;
										assign node2829 = (inp[3]) ? node2833 : node2830;
											assign node2830 = (inp[1]) ? 13'b0000000011111 : 13'b0000000111111;
											assign node2833 = (inp[1]) ? 13'b0000000001111 : 13'b0000000011111;
								assign node2836 = (inp[3]) ? node2852 : node2837;
									assign node2837 = (inp[6]) ? node2845 : node2838;
										assign node2838 = (inp[5]) ? node2842 : node2839;
											assign node2839 = (inp[10]) ? 13'b0000000111111 : 13'b0000001111111;
											assign node2842 = (inp[10]) ? 13'b0000000011111 : 13'b0000000111111;
										assign node2845 = (inp[10]) ? node2849 : node2846;
											assign node2846 = (inp[9]) ? 13'b0000000011111 : 13'b0000000011111;
											assign node2849 = (inp[5]) ? 13'b0000000001111 : 13'b0000000001111;
									assign node2852 = (inp[5]) ? node2858 : node2853;
										assign node2853 = (inp[10]) ? node2855 : 13'b0000000011111;
											assign node2855 = (inp[1]) ? 13'b0000000001111 : 13'b0000000001111;
										assign node2858 = (inp[1]) ? node2862 : node2859;
											assign node2859 = (inp[6]) ? 13'b0000000001111 : 13'b0000000011111;
											assign node2862 = (inp[9]) ? 13'b0000000000011 : 13'b0000000001111;
							assign node2865 = (inp[10]) ? node2895 : node2866;
								assign node2866 = (inp[9]) ? node2882 : node2867;
									assign node2867 = (inp[1]) ? node2875 : node2868;
										assign node2868 = (inp[7]) ? node2872 : node2869;
											assign node2869 = (inp[5]) ? 13'b0000000111111 : 13'b0000001111111;
											assign node2872 = (inp[6]) ? 13'b0000000011111 : 13'b0000000111111;
										assign node2875 = (inp[3]) ? node2879 : node2876;
											assign node2876 = (inp[6]) ? 13'b0000000011111 : 13'b0000000111111;
											assign node2879 = (inp[7]) ? 13'b0000000000111 : 13'b0000000011111;
									assign node2882 = (inp[1]) ? node2888 : node2883;
										assign node2883 = (inp[6]) ? node2885 : 13'b0000000011111;
											assign node2885 = (inp[3]) ? 13'b0000000001111 : 13'b0000000011111;
										assign node2888 = (inp[6]) ? node2892 : node2889;
											assign node2889 = (inp[7]) ? 13'b0000000001111 : 13'b0000000001111;
											assign node2892 = (inp[3]) ? 13'b0000000000111 : 13'b0000000001111;
								assign node2895 = (inp[3]) ? node2909 : node2896;
									assign node2896 = (inp[7]) ? node2902 : node2897;
										assign node2897 = (inp[1]) ? node2899 : 13'b0000000011111;
											assign node2899 = (inp[6]) ? 13'b0000000001111 : 13'b0000000011111;
										assign node2902 = (inp[9]) ? node2906 : node2903;
											assign node2903 = (inp[1]) ? 13'b0000000001111 : 13'b0000000001111;
											assign node2906 = (inp[6]) ? 13'b0000000000111 : 13'b0000000001111;
									assign node2909 = (inp[5]) ? node2915 : node2910;
										assign node2910 = (inp[1]) ? node2912 : 13'b0000000001111;
											assign node2912 = (inp[6]) ? 13'b0000000000111 : 13'b0000000001111;
										assign node2915 = (inp[9]) ? node2919 : node2916;
											assign node2916 = (inp[7]) ? 13'b0000000000111 : 13'b0000000000111;
											assign node2919 = (inp[6]) ? 13'b0000000000001 : 13'b0000000000111;
			assign node2922 = (inp[7]) ? node3408 : node2923;
				assign node2923 = (inp[6]) ? node3165 : node2924;
					assign node2924 = (inp[5]) ? node3048 : node2925;
						assign node2925 = (inp[10]) ? node2987 : node2926;
							assign node2926 = (inp[9]) ? node2956 : node2927;
								assign node2927 = (inp[3]) ? node2943 : node2928;
									assign node2928 = (inp[0]) ? node2936 : node2929;
										assign node2929 = (inp[1]) ? node2933 : node2930;
											assign node2930 = (inp[2]) ? 13'b0000111111111 : 13'b0001111111111;
											assign node2933 = (inp[2]) ? 13'b0000011111111 : 13'b0000111111111;
										assign node2936 = (inp[11]) ? node2940 : node2937;
											assign node2937 = (inp[4]) ? 13'b0000011111111 : 13'b0000111111111;
											assign node2940 = (inp[1]) ? 13'b0000001111111 : 13'b0000011111111;
									assign node2943 = (inp[0]) ? node2951 : node2944;
										assign node2944 = (inp[1]) ? node2948 : node2945;
											assign node2945 = (inp[4]) ? 13'b0000011111111 : 13'b0000111111111;
											assign node2948 = (inp[11]) ? 13'b0000000111111 : 13'b0000011111111;
										assign node2951 = (inp[11]) ? 13'b0000001111111 : node2952;
											assign node2952 = (inp[4]) ? 13'b0000001111111 : 13'b0000011111111;
								assign node2956 = (inp[2]) ? node2972 : node2957;
									assign node2957 = (inp[0]) ? node2965 : node2958;
										assign node2958 = (inp[3]) ? node2962 : node2959;
											assign node2959 = (inp[11]) ? 13'b0000011111111 : 13'b0000111111111;
											assign node2962 = (inp[4]) ? 13'b0000001111111 : 13'b0000011111111;
										assign node2965 = (inp[4]) ? node2969 : node2966;
											assign node2966 = (inp[11]) ? 13'b0000001111111 : 13'b0000011111111;
											assign node2969 = (inp[11]) ? 13'b0000000111111 : 13'b0000001111111;
									assign node2972 = (inp[11]) ? node2980 : node2973;
										assign node2973 = (inp[1]) ? node2977 : node2974;
											assign node2974 = (inp[0]) ? 13'b0000001111111 : 13'b0000111111111;
											assign node2977 = (inp[4]) ? 13'b0000000111111 : 13'b0000001111111;
										assign node2980 = (inp[4]) ? node2984 : node2981;
											assign node2981 = (inp[0]) ? 13'b0000000111111 : 13'b0000001111111;
											assign node2984 = (inp[1]) ? 13'b0000000011111 : 13'b0000000111111;
							assign node2987 = (inp[3]) ? node3017 : node2988;
								assign node2988 = (inp[11]) ? node3002 : node2989;
									assign node2989 = (inp[4]) ? node2995 : node2990;
										assign node2990 = (inp[0]) ? 13'b0000011111111 : node2991;
											assign node2991 = (inp[2]) ? 13'b0000011111111 : 13'b0000111111111;
										assign node2995 = (inp[1]) ? node2999 : node2996;
											assign node2996 = (inp[9]) ? 13'b0000001111111 : 13'b0000001111111;
											assign node2999 = (inp[0]) ? 13'b0000000111111 : 13'b0000001111111;
									assign node3002 = (inp[0]) ? node3010 : node3003;
										assign node3003 = (inp[4]) ? node3007 : node3004;
											assign node3004 = (inp[1]) ? 13'b0000001111111 : 13'b0000011111111;
											assign node3007 = (inp[1]) ? 13'b0000000111111 : 13'b0000001111111;
										assign node3010 = (inp[2]) ? node3014 : node3011;
											assign node3011 = (inp[1]) ? 13'b0000000011111 : 13'b0000001111111;
											assign node3014 = (inp[9]) ? 13'b0000000011111 : 13'b0000000111111;
								assign node3017 = (inp[1]) ? node3033 : node3018;
									assign node3018 = (inp[4]) ? node3026 : node3019;
										assign node3019 = (inp[0]) ? node3023 : node3020;
											assign node3020 = (inp[9]) ? 13'b0000001111111 : 13'b0000001111111;
											assign node3023 = (inp[11]) ? 13'b0000000111111 : 13'b0000001111111;
										assign node3026 = (inp[2]) ? node3030 : node3027;
											assign node3027 = (inp[0]) ? 13'b0000000111111 : 13'b0000001111111;
											assign node3030 = (inp[11]) ? 13'b0000000011111 : 13'b0000000111111;
									assign node3033 = (inp[4]) ? node3041 : node3034;
										assign node3034 = (inp[0]) ? node3038 : node3035;
											assign node3035 = (inp[11]) ? 13'b0000000111111 : 13'b0000001111111;
											assign node3038 = (inp[9]) ? 13'b0000000011111 : 13'b0000000111111;
										assign node3041 = (inp[2]) ? node3045 : node3042;
											assign node3042 = (inp[9]) ? 13'b0000000011111 : 13'b0000000111111;
											assign node3045 = (inp[9]) ? 13'b0000000000111 : 13'b0000000011111;
						assign node3048 = (inp[9]) ? node3106 : node3049;
							assign node3049 = (inp[10]) ? node3075 : node3050;
								assign node3050 = (inp[2]) ? node3062 : node3051;
									assign node3051 = (inp[3]) ? node3057 : node3052;
										assign node3052 = (inp[1]) ? 13'b0000011111111 : node3053;
											assign node3053 = (inp[0]) ? 13'b0000011111111 : 13'b0000111111111;
										assign node3057 = (inp[11]) ? 13'b0000001111111 : node3058;
											assign node3058 = (inp[1]) ? 13'b0000001111111 : 13'b0000011111111;
									assign node3062 = (inp[1]) ? node3068 : node3063;
										assign node3063 = (inp[4]) ? node3065 : 13'b0000011111111;
											assign node3065 = (inp[0]) ? 13'b0000000111111 : 13'b0000001111111;
										assign node3068 = (inp[4]) ? node3072 : node3069;
											assign node3069 = (inp[3]) ? 13'b0000000111111 : 13'b0000001111111;
											assign node3072 = (inp[0]) ? 13'b0000000011111 : 13'b0000000111111;
								assign node3075 = (inp[2]) ? node3091 : node3076;
									assign node3076 = (inp[3]) ? node3084 : node3077;
										assign node3077 = (inp[0]) ? node3081 : node3078;
											assign node3078 = (inp[4]) ? 13'b0000001111111 : 13'b0000011111111;
											assign node3081 = (inp[1]) ? 13'b0000000011111 : 13'b0000001111111;
										assign node3084 = (inp[11]) ? node3088 : node3085;
											assign node3085 = (inp[1]) ? 13'b0000000111111 : 13'b0000001111111;
											assign node3088 = (inp[4]) ? 13'b0000000011111 : 13'b0000000111111;
									assign node3091 = (inp[4]) ? node3099 : node3092;
										assign node3092 = (inp[3]) ? node3096 : node3093;
											assign node3093 = (inp[11]) ? 13'b0000000111111 : 13'b0000001111111;
											assign node3096 = (inp[0]) ? 13'b0000000011111 : 13'b0000000111111;
										assign node3099 = (inp[1]) ? node3103 : node3100;
											assign node3100 = (inp[11]) ? 13'b0000000011111 : 13'b0000000111111;
											assign node3103 = (inp[3]) ? 13'b0000000001111 : 13'b0000000011111;
							assign node3106 = (inp[2]) ? node3136 : node3107;
								assign node3107 = (inp[4]) ? node3121 : node3108;
									assign node3108 = (inp[10]) ? node3114 : node3109;
										assign node3109 = (inp[11]) ? node3111 : 13'b0000001111111;
											assign node3111 = (inp[1]) ? 13'b0000000111111 : 13'b0000011111111;
										assign node3114 = (inp[0]) ? node3118 : node3115;
											assign node3115 = (inp[1]) ? 13'b0000000111111 : 13'b0000001111111;
											assign node3118 = (inp[11]) ? 13'b0000000011111 : 13'b0000000111111;
									assign node3121 = (inp[0]) ? node3129 : node3122;
										assign node3122 = (inp[1]) ? node3126 : node3123;
											assign node3123 = (inp[10]) ? 13'b0000000111111 : 13'b0000000111111;
											assign node3126 = (inp[11]) ? 13'b0000000011111 : 13'b0000000111111;
										assign node3129 = (inp[10]) ? node3133 : node3130;
											assign node3130 = (inp[11]) ? 13'b0000000011111 : 13'b0000000111111;
											assign node3133 = (inp[11]) ? 13'b0000000001111 : 13'b0000000011111;
								assign node3136 = (inp[11]) ? node3152 : node3137;
									assign node3137 = (inp[4]) ? node3145 : node3138;
										assign node3138 = (inp[1]) ? node3142 : node3139;
											assign node3139 = (inp[10]) ? 13'b0000000111111 : 13'b0000000111111;
											assign node3142 = (inp[0]) ? 13'b0000000011111 : 13'b0000000111111;
										assign node3145 = (inp[3]) ? node3149 : node3146;
											assign node3146 = (inp[10]) ? 13'b0000000011111 : 13'b0000000111111;
											assign node3149 = (inp[10]) ? 13'b0000000001111 : 13'b0000000011111;
									assign node3152 = (inp[0]) ? node3158 : node3153;
										assign node3153 = (inp[1]) ? node3155 : 13'b0000000111111;
											assign node3155 = (inp[3]) ? 13'b0000000001111 : 13'b0000000011111;
										assign node3158 = (inp[4]) ? node3162 : node3159;
											assign node3159 = (inp[10]) ? 13'b0000000001111 : 13'b0000000011111;
											assign node3162 = (inp[1]) ? 13'b0000000000111 : 13'b0000000001111;
					assign node3165 = (inp[10]) ? node3289 : node3166;
						assign node3166 = (inp[3]) ? node3226 : node3167;
							assign node3167 = (inp[5]) ? node3197 : node3168;
								assign node3168 = (inp[4]) ? node3182 : node3169;
									assign node3169 = (inp[0]) ? node3175 : node3170;
										assign node3170 = (inp[1]) ? 13'b0000001111111 : node3171;
											assign node3171 = (inp[11]) ? 13'b0000011111111 : 13'b0000111111111;
										assign node3175 = (inp[1]) ? node3179 : node3176;
											assign node3176 = (inp[11]) ? 13'b0000000111111 : 13'b0000001111111;
											assign node3179 = (inp[2]) ? 13'b0000001111111 : 13'b0000001111111;
									assign node3182 = (inp[9]) ? node3190 : node3183;
										assign node3183 = (inp[1]) ? node3187 : node3184;
											assign node3184 = (inp[11]) ? 13'b0000001111111 : 13'b0000011111111;
											assign node3187 = (inp[0]) ? 13'b0000000111111 : 13'b0000001111111;
										assign node3190 = (inp[1]) ? node3194 : node3191;
											assign node3191 = (inp[2]) ? 13'b0000000111111 : 13'b0000000111111;
											assign node3194 = (inp[11]) ? 13'b0000000011111 : 13'b0000001111111;
								assign node3197 = (inp[4]) ? node3211 : node3198;
									assign node3198 = (inp[9]) ? node3204 : node3199;
										assign node3199 = (inp[0]) ? 13'b0000001111111 : node3200;
											assign node3200 = (inp[1]) ? 13'b0000001111111 : 13'b0000011111111;
										assign node3204 = (inp[2]) ? node3208 : node3205;
											assign node3205 = (inp[1]) ? 13'b0000000111111 : 13'b0000001111111;
											assign node3208 = (inp[11]) ? 13'b0000000011111 : 13'b0000000111111;
									assign node3211 = (inp[0]) ? node3219 : node3212;
										assign node3212 = (inp[9]) ? node3216 : node3213;
											assign node3213 = (inp[11]) ? 13'b0000000111111 : 13'b0000001111111;
											assign node3216 = (inp[2]) ? 13'b0000000011111 : 13'b0000000111111;
										assign node3219 = (inp[1]) ? node3223 : node3220;
											assign node3220 = (inp[2]) ? 13'b0000000011111 : 13'b0000000111111;
											assign node3223 = (inp[9]) ? 13'b0000000000111 : 13'b0000000011111;
							assign node3226 = (inp[2]) ? node3258 : node3227;
								assign node3227 = (inp[11]) ? node3243 : node3228;
									assign node3228 = (inp[4]) ? node3236 : node3229;
										assign node3229 = (inp[0]) ? node3233 : node3230;
											assign node3230 = (inp[5]) ? 13'b0000001111111 : 13'b0000011111111;
											assign node3233 = (inp[1]) ? 13'b0000000111111 : 13'b0000001111111;
										assign node3236 = (inp[9]) ? node3240 : node3237;
											assign node3237 = (inp[1]) ? 13'b0000000111111 : 13'b0000000111111;
											assign node3240 = (inp[5]) ? 13'b0000000001111 : 13'b0000000011111;
									assign node3243 = (inp[1]) ? node3251 : node3244;
										assign node3244 = (inp[5]) ? node3248 : node3245;
											assign node3245 = (inp[4]) ? 13'b0000000111111 : 13'b0000001111111;
											assign node3248 = (inp[0]) ? 13'b0000000011111 : 13'b0000000111111;
										assign node3251 = (inp[9]) ? node3255 : node3252;
											assign node3252 = (inp[0]) ? 13'b0000000011111 : 13'b0000000111111;
											assign node3255 = (inp[0]) ? 13'b0000000001111 : 13'b0000000011111;
								assign node3258 = (inp[9]) ? node3274 : node3259;
									assign node3259 = (inp[11]) ? node3267 : node3260;
										assign node3260 = (inp[0]) ? node3264 : node3261;
											assign node3261 = (inp[1]) ? 13'b0000000111111 : 13'b0000001111111;
											assign node3264 = (inp[1]) ? 13'b0000000011111 : 13'b0000000111111;
										assign node3267 = (inp[4]) ? node3271 : node3268;
											assign node3268 = (inp[0]) ? 13'b0000000011111 : 13'b0000000111111;
											assign node3271 = (inp[1]) ? 13'b0000000001111 : 13'b0000000011111;
									assign node3274 = (inp[0]) ? node3282 : node3275;
										assign node3275 = (inp[4]) ? node3279 : node3276;
											assign node3276 = (inp[11]) ? 13'b0000000011111 : 13'b0000000111111;
											assign node3279 = (inp[1]) ? 13'b0000000001111 : 13'b0000000011111;
										assign node3282 = (inp[4]) ? node3286 : node3283;
											assign node3283 = (inp[5]) ? 13'b0000000001111 : 13'b0000000011111;
											assign node3286 = (inp[11]) ? 13'b0000000000111 : 13'b0000000001111;
						assign node3289 = (inp[5]) ? node3347 : node3290;
							assign node3290 = (inp[1]) ? node3316 : node3291;
								assign node3291 = (inp[0]) ? node3301 : node3292;
									assign node3292 = (inp[9]) ? 13'b0000000111111 : node3293;
										assign node3293 = (inp[3]) ? node3297 : node3294;
											assign node3294 = (inp[4]) ? 13'b0000000111111 : 13'b0000011111111;
											assign node3297 = (inp[11]) ? 13'b0000000111111 : 13'b0000001111111;
									assign node3301 = (inp[4]) ? node3309 : node3302;
										assign node3302 = (inp[11]) ? node3306 : node3303;
											assign node3303 = (inp[9]) ? 13'b0000000111111 : 13'b0000001111111;
											assign node3306 = (inp[2]) ? 13'b0000000011111 : 13'b0000000111111;
										assign node3309 = (inp[3]) ? node3313 : node3310;
											assign node3310 = (inp[11]) ? 13'b0000000011111 : 13'b0000000111111;
											assign node3313 = (inp[11]) ? 13'b0000000001111 : 13'b0000000011111;
								assign node3316 = (inp[3]) ? node3332 : node3317;
									assign node3317 = (inp[2]) ? node3325 : node3318;
										assign node3318 = (inp[9]) ? node3322 : node3319;
											assign node3319 = (inp[4]) ? 13'b0000000111111 : 13'b0000001111111;
											assign node3322 = (inp[0]) ? 13'b0000000011111 : 13'b0000000111111;
										assign node3325 = (inp[0]) ? node3329 : node3326;
											assign node3326 = (inp[9]) ? 13'b0000000011111 : 13'b0000000111111;
											assign node3329 = (inp[9]) ? 13'b0000000001111 : 13'b0000000011111;
									assign node3332 = (inp[9]) ? node3340 : node3333;
										assign node3333 = (inp[11]) ? node3337 : node3334;
											assign node3334 = (inp[0]) ? 13'b0000000011111 : 13'b0000000111111;
											assign node3337 = (inp[4]) ? 13'b0000000001111 : 13'b0000000011111;
										assign node3340 = (inp[4]) ? node3344 : node3341;
											assign node3341 = (inp[0]) ? 13'b0000000001111 : 13'b0000000011111;
											assign node3344 = (inp[11]) ? 13'b0000000000111 : 13'b0000000001111;
							assign node3347 = (inp[2]) ? node3377 : node3348;
								assign node3348 = (inp[9]) ? node3362 : node3349;
									assign node3349 = (inp[3]) ? node3357 : node3350;
										assign node3350 = (inp[1]) ? node3354 : node3351;
											assign node3351 = (inp[0]) ? 13'b0000000111111 : 13'b0000000111111;
											assign node3354 = (inp[4]) ? 13'b0000000011111 : 13'b0000000111111;
										assign node3357 = (inp[0]) ? 13'b0000000011111 : node3358;
											assign node3358 = (inp[11]) ? 13'b0000000011111 : 13'b0000000111111;
									assign node3362 = (inp[0]) ? node3370 : node3363;
										assign node3363 = (inp[4]) ? node3367 : node3364;
											assign node3364 = (inp[11]) ? 13'b0000000011111 : 13'b0000000111111;
											assign node3367 = (inp[3]) ? 13'b0000000001111 : 13'b0000000011111;
										assign node3370 = (inp[4]) ? node3374 : node3371;
											assign node3371 = (inp[1]) ? 13'b0000000001111 : 13'b0000000011111;
											assign node3374 = (inp[11]) ? 13'b0000000000111 : 13'b0000000001111;
								assign node3377 = (inp[4]) ? node3393 : node3378;
									assign node3378 = (inp[11]) ? node3386 : node3379;
										assign node3379 = (inp[9]) ? node3383 : node3380;
											assign node3380 = (inp[0]) ? 13'b0000000011111 : 13'b0000000111111;
											assign node3383 = (inp[3]) ? 13'b0000000001111 : 13'b0000000011111;
										assign node3386 = (inp[0]) ? node3390 : node3387;
											assign node3387 = (inp[9]) ? 13'b0000000001111 : 13'b0000000011111;
											assign node3390 = (inp[3]) ? 13'b0000000000111 : 13'b0000000001111;
									assign node3393 = (inp[0]) ? node3401 : node3394;
										assign node3394 = (inp[3]) ? node3398 : node3395;
											assign node3395 = (inp[9]) ? 13'b0000000001111 : 13'b0000000001111;
											assign node3398 = (inp[9]) ? 13'b0000000000111 : 13'b0000000001111;
										assign node3401 = (inp[9]) ? node3405 : node3402;
											assign node3402 = (inp[1]) ? 13'b0000000000111 : 13'b0000000000111;
											assign node3405 = (inp[3]) ? 13'b0000000000011 : 13'b0000000000111;
				assign node3408 = (inp[1]) ? node3654 : node3409;
					assign node3409 = (inp[5]) ? node3529 : node3410;
						assign node3410 = (inp[2]) ? node3470 : node3411;
							assign node3411 = (inp[3]) ? node3441 : node3412;
								assign node3412 = (inp[11]) ? node3426 : node3413;
									assign node3413 = (inp[6]) ? node3421 : node3414;
										assign node3414 = (inp[4]) ? node3418 : node3415;
											assign node3415 = (inp[10]) ? 13'b0000011111111 : 13'b0000111111111;
											assign node3418 = (inp[0]) ? 13'b0000001111111 : 13'b0000011111111;
										assign node3421 = (inp[4]) ? node3423 : 13'b0000001111111;
											assign node3423 = (inp[9]) ? 13'b0000000111111 : 13'b0000001111111;
									assign node3426 = (inp[0]) ? node3434 : node3427;
										assign node3427 = (inp[6]) ? node3431 : node3428;
											assign node3428 = (inp[4]) ? 13'b0000001111111 : 13'b0000001111111;
											assign node3431 = (inp[10]) ? 13'b0000000011111 : 13'b0000001111111;
										assign node3434 = (inp[10]) ? node3438 : node3435;
											assign node3435 = (inp[9]) ? 13'b0000000111111 : 13'b0000001111111;
											assign node3438 = (inp[9]) ? 13'b0000000011111 : 13'b0000000111111;
								assign node3441 = (inp[4]) ? node3455 : node3442;
									assign node3442 = (inp[6]) ? node3448 : node3443;
										assign node3443 = (inp[0]) ? 13'b0000001111111 : node3444;
											assign node3444 = (inp[10]) ? 13'b0000000111111 : 13'b0000001111111;
										assign node3448 = (inp[10]) ? node3452 : node3449;
											assign node3449 = (inp[9]) ? 13'b0000000111111 : 13'b0000001111111;
											assign node3452 = (inp[0]) ? 13'b0000000011111 : 13'b0000000111111;
									assign node3455 = (inp[0]) ? node3463 : node3456;
										assign node3456 = (inp[6]) ? node3460 : node3457;
											assign node3457 = (inp[10]) ? 13'b0000000111111 : 13'b0000011111111;
											assign node3460 = (inp[9]) ? 13'b0000000011111 : 13'b0000000111111;
										assign node3463 = (inp[11]) ? node3467 : node3464;
											assign node3464 = (inp[9]) ? 13'b0000000011111 : 13'b0000000111111;
											assign node3467 = (inp[6]) ? 13'b0000000001111 : 13'b0000000011111;
							assign node3470 = (inp[3]) ? node3502 : node3471;
								assign node3471 = (inp[6]) ? node3487 : node3472;
									assign node3472 = (inp[9]) ? node3480 : node3473;
										assign node3473 = (inp[10]) ? node3477 : node3474;
											assign node3474 = (inp[0]) ? 13'b0000001111111 : 13'b0000011111111;
											assign node3477 = (inp[11]) ? 13'b0000000111111 : 13'b0000001111111;
										assign node3480 = (inp[11]) ? node3484 : node3481;
											assign node3481 = (inp[10]) ? 13'b0000000111111 : 13'b0000000111111;
											assign node3484 = (inp[10]) ? 13'b0000000011111 : 13'b0000000111111;
									assign node3487 = (inp[4]) ? node3495 : node3488;
										assign node3488 = (inp[9]) ? node3492 : node3489;
											assign node3489 = (inp[0]) ? 13'b0000000111111 : 13'b0000001111111;
											assign node3492 = (inp[0]) ? 13'b0000000011111 : 13'b0000000111111;
										assign node3495 = (inp[11]) ? node3499 : node3496;
											assign node3496 = (inp[9]) ? 13'b0000000011111 : 13'b0000000111111;
											assign node3499 = (inp[0]) ? 13'b0000000001111 : 13'b0000000011111;
								assign node3502 = (inp[4]) ? node3516 : node3503;
									assign node3503 = (inp[0]) ? node3509 : node3504;
										assign node3504 = (inp[11]) ? node3506 : 13'b0000001111111;
											assign node3506 = (inp[6]) ? 13'b0000000011111 : 13'b0000000111111;
										assign node3509 = (inp[9]) ? node3513 : node3510;
											assign node3510 = (inp[6]) ? 13'b0000000011111 : 13'b0000000011111;
											assign node3513 = (inp[6]) ? 13'b0000000001111 : 13'b0000000011111;
									assign node3516 = (inp[6]) ? node3524 : node3517;
										assign node3517 = (inp[9]) ? node3521 : node3518;
											assign node3518 = (inp[11]) ? 13'b0000000011111 : 13'b0000000111111;
											assign node3521 = (inp[10]) ? 13'b0000000001111 : 13'b0000000011111;
										assign node3524 = (inp[10]) ? node3526 : 13'b0000000001111;
											assign node3526 = (inp[11]) ? 13'b0000000000111 : 13'b0000000001111;
						assign node3529 = (inp[3]) ? node3591 : node3530;
							assign node3530 = (inp[6]) ? node3560 : node3531;
								assign node3531 = (inp[11]) ? node3545 : node3532;
									assign node3532 = (inp[0]) ? node3540 : node3533;
										assign node3533 = (inp[9]) ? node3537 : node3534;
											assign node3534 = (inp[4]) ? 13'b0000001111111 : 13'b0000011111111;
											assign node3537 = (inp[10]) ? 13'b0000000011111 : 13'b0000000111111;
										assign node3540 = (inp[2]) ? node3542 : 13'b0000000111111;
											assign node3542 = (inp[4]) ? 13'b0000000011111 : 13'b0000000111111;
									assign node3545 = (inp[4]) ? node3553 : node3546;
										assign node3546 = (inp[10]) ? node3550 : node3547;
											assign node3547 = (inp[2]) ? 13'b0000000111111 : 13'b0000001111111;
											assign node3550 = (inp[0]) ? 13'b0000000011111 : 13'b0000000111111;
										assign node3553 = (inp[2]) ? node3557 : node3554;
											assign node3554 = (inp[10]) ? 13'b0000000011111 : 13'b0000000111111;
											assign node3557 = (inp[9]) ? 13'b0000000001111 : 13'b0000000011111;
								assign node3560 = (inp[0]) ? node3576 : node3561;
									assign node3561 = (inp[4]) ? node3569 : node3562;
										assign node3562 = (inp[9]) ? node3566 : node3563;
											assign node3563 = (inp[10]) ? 13'b0000000111111 : 13'b0000001111111;
											assign node3566 = (inp[10]) ? 13'b0000000011111 : 13'b0000000111111;
										assign node3569 = (inp[10]) ? node3573 : node3570;
											assign node3570 = (inp[11]) ? 13'b0000000011111 : 13'b0000000111111;
											assign node3573 = (inp[2]) ? 13'b0000000001111 : 13'b0000000011111;
									assign node3576 = (inp[9]) ? node3584 : node3577;
										assign node3577 = (inp[4]) ? node3581 : node3578;
											assign node3578 = (inp[11]) ? 13'b0000000011111 : 13'b0000000111111;
											assign node3581 = (inp[2]) ? 13'b0000000001111 : 13'b0000000011111;
										assign node3584 = (inp[4]) ? node3588 : node3585;
											assign node3585 = (inp[10]) ? 13'b0000000001111 : 13'b0000000001111;
											assign node3588 = (inp[2]) ? 13'b0000000000111 : 13'b0000000001111;
							assign node3591 = (inp[4]) ? node3623 : node3592;
								assign node3592 = (inp[11]) ? node3608 : node3593;
									assign node3593 = (inp[9]) ? node3601 : node3594;
										assign node3594 = (inp[6]) ? node3598 : node3595;
											assign node3595 = (inp[0]) ? 13'b0000000111111 : 13'b0000001111111;
											assign node3598 = (inp[2]) ? 13'b0000000011111 : 13'b0000000111111;
										assign node3601 = (inp[10]) ? node3605 : node3602;
											assign node3602 = (inp[2]) ? 13'b0000000011111 : 13'b0000000011111;
											assign node3605 = (inp[6]) ? 13'b0000000001111 : 13'b0000000011111;
									assign node3608 = (inp[9]) ? node3616 : node3609;
										assign node3609 = (inp[0]) ? node3613 : node3610;
											assign node3610 = (inp[10]) ? 13'b0000000001111 : 13'b0000000111111;
											assign node3613 = (inp[2]) ? 13'b0000000001111 : 13'b0000000011111;
										assign node3616 = (inp[6]) ? node3620 : node3617;
											assign node3617 = (inp[0]) ? 13'b0000000001111 : 13'b0000000011111;
											assign node3620 = (inp[2]) ? 13'b0000000000111 : 13'b0000000001111;
								assign node3623 = (inp[6]) ? node3639 : node3624;
									assign node3624 = (inp[2]) ? node3632 : node3625;
										assign node3625 = (inp[9]) ? node3629 : node3626;
											assign node3626 = (inp[0]) ? 13'b0000000011111 : 13'b0000000111111;
											assign node3629 = (inp[10]) ? 13'b0000000001111 : 13'b0000000011111;
										assign node3632 = (inp[10]) ? node3636 : node3633;
											assign node3633 = (inp[0]) ? 13'b0000000001111 : 13'b0000000011111;
											assign node3636 = (inp[11]) ? 13'b0000000000111 : 13'b0000000001111;
									assign node3639 = (inp[0]) ? node3647 : node3640;
										assign node3640 = (inp[11]) ? node3644 : node3641;
											assign node3641 = (inp[10]) ? 13'b0000000001111 : 13'b0000000011111;
											assign node3644 = (inp[9]) ? 13'b0000000000111 : 13'b0000000000111;
										assign node3647 = (inp[11]) ? node3651 : node3648;
											assign node3648 = (inp[9]) ? 13'b0000000000111 : 13'b0000000001111;
											assign node3651 = (inp[9]) ? 13'b0000000000011 : 13'b0000000000111;
					assign node3654 = (inp[4]) ? node3776 : node3655;
						assign node3655 = (inp[10]) ? node3713 : node3656;
							assign node3656 = (inp[2]) ? node3686 : node3657;
								assign node3657 = (inp[9]) ? node3671 : node3658;
									assign node3658 = (inp[6]) ? node3666 : node3659;
										assign node3659 = (inp[3]) ? node3663 : node3660;
											assign node3660 = (inp[5]) ? 13'b0000001111111 : 13'b0000001111111;
											assign node3663 = (inp[0]) ? 13'b0000000111111 : 13'b0000001111111;
										assign node3666 = (inp[5]) ? 13'b0000000111111 : node3667;
											assign node3667 = (inp[0]) ? 13'b0000000111111 : 13'b0000001111111;
									assign node3671 = (inp[11]) ? node3679 : node3672;
										assign node3672 = (inp[5]) ? node3676 : node3673;
											assign node3673 = (inp[3]) ? 13'b0000000111111 : 13'b0000001111111;
											assign node3676 = (inp[0]) ? 13'b0000000011111 : 13'b0000000111111;
										assign node3679 = (inp[5]) ? node3683 : node3680;
											assign node3680 = (inp[6]) ? 13'b0000000011111 : 13'b0000000011111;
											assign node3683 = (inp[3]) ? 13'b0000000000111 : 13'b0000000011111;
								assign node3686 = (inp[3]) ? node3700 : node3687;
									assign node3687 = (inp[6]) ? node3695 : node3688;
										assign node3688 = (inp[5]) ? node3692 : node3689;
											assign node3689 = (inp[0]) ? 13'b0000000111111 : 13'b0000001111111;
											assign node3692 = (inp[11]) ? 13'b0000000001111 : 13'b0000000111111;
										assign node3695 = (inp[9]) ? node3697 : 13'b0000000011111;
											assign node3697 = (inp[0]) ? 13'b0000000001111 : 13'b0000000011111;
									assign node3700 = (inp[5]) ? node3706 : node3701;
										assign node3701 = (inp[11]) ? node3703 : 13'b0000000111111;
											assign node3703 = (inp[9]) ? 13'b0000000001111 : 13'b0000000011111;
										assign node3706 = (inp[11]) ? node3710 : node3707;
											assign node3707 = (inp[9]) ? 13'b0000000001111 : 13'b0000000111111;
											assign node3710 = (inp[0]) ? 13'b0000000000111 : 13'b0000000001111;
							assign node3713 = (inp[0]) ? node3745 : node3714;
								assign node3714 = (inp[11]) ? node3730 : node3715;
									assign node3715 = (inp[5]) ? node3723 : node3716;
										assign node3716 = (inp[9]) ? node3720 : node3717;
											assign node3717 = (inp[3]) ? 13'b0000000111111 : 13'b0000001111111;
											assign node3720 = (inp[2]) ? 13'b0000000011111 : 13'b0000000111111;
										assign node3723 = (inp[6]) ? node3727 : node3724;
											assign node3724 = (inp[3]) ? 13'b0000000011111 : 13'b0000000111111;
											assign node3727 = (inp[9]) ? 13'b0000000001111 : 13'b0000000011111;
									assign node3730 = (inp[6]) ? node3738 : node3731;
										assign node3731 = (inp[9]) ? node3735 : node3732;
											assign node3732 = (inp[5]) ? 13'b0000000011111 : 13'b0000000111111;
											assign node3735 = (inp[5]) ? 13'b0000000001111 : 13'b0000000011111;
										assign node3738 = (inp[3]) ? node3742 : node3739;
											assign node3739 = (inp[9]) ? 13'b0000000001111 : 13'b0000000011111;
											assign node3742 = (inp[9]) ? 13'b0000000000011 : 13'b0000000001111;
								assign node3745 = (inp[3]) ? node3761 : node3746;
									assign node3746 = (inp[2]) ? node3754 : node3747;
										assign node3747 = (inp[11]) ? node3751 : node3748;
											assign node3748 = (inp[6]) ? 13'b0000000011111 : 13'b0000000111111;
											assign node3751 = (inp[6]) ? 13'b0000000000111 : 13'b0000000011111;
										assign node3754 = (inp[9]) ? node3758 : node3755;
											assign node3755 = (inp[11]) ? 13'b0000000001111 : 13'b0000000011111;
											assign node3758 = (inp[5]) ? 13'b0000000000111 : 13'b0000000000111;
									assign node3761 = (inp[2]) ? node3769 : node3762;
										assign node3762 = (inp[5]) ? node3766 : node3763;
											assign node3763 = (inp[6]) ? 13'b0000000001111 : 13'b0000000001111;
											assign node3766 = (inp[6]) ? 13'b0000000000111 : 13'b0000000000111;
										assign node3769 = (inp[11]) ? node3773 : node3770;
											assign node3770 = (inp[5]) ? 13'b0000000000111 : 13'b0000000001111;
											assign node3773 = (inp[9]) ? 13'b0000000000011 : 13'b0000000000111;
						assign node3776 = (inp[11]) ? node3830 : node3777;
							assign node3777 = (inp[10]) ? node3807 : node3778;
								assign node3778 = (inp[0]) ? node3792 : node3779;
									assign node3779 = (inp[2]) ? node3785 : node3780;
										assign node3780 = (inp[5]) ? 13'b0000000011111 : node3781;
											assign node3781 = (inp[3]) ? 13'b0000000111111 : 13'b0000001111111;
										assign node3785 = (inp[5]) ? node3789 : node3786;
											assign node3786 = (inp[3]) ? 13'b0000000011111 : 13'b0000000011111;
											assign node3789 = (inp[6]) ? 13'b0000000000111 : 13'b0000000011111;
									assign node3792 = (inp[6]) ? node3800 : node3793;
										assign node3793 = (inp[2]) ? node3797 : node3794;
											assign node3794 = (inp[5]) ? 13'b0000000011111 : 13'b0000000111111;
											assign node3797 = (inp[5]) ? 13'b0000000001111 : 13'b0000000001111;
										assign node3800 = (inp[9]) ? node3804 : node3801;
											assign node3801 = (inp[3]) ? 13'b0000000001111 : 13'b0000000011111;
											assign node3804 = (inp[2]) ? 13'b0000000000111 : 13'b0000000001111;
								assign node3807 = (inp[6]) ? node3817 : node3808;
									assign node3808 = (inp[5]) ? 13'b0000000001111 : node3809;
										assign node3809 = (inp[0]) ? node3813 : node3810;
											assign node3810 = (inp[2]) ? 13'b0000000111111 : 13'b0000000011111;
											assign node3813 = (inp[9]) ? 13'b0000000001111 : 13'b0000000011111;
									assign node3817 = (inp[9]) ? node3825 : node3818;
										assign node3818 = (inp[0]) ? node3822 : node3819;
											assign node3819 = (inp[3]) ? 13'b0000000001111 : 13'b0000000011111;
											assign node3822 = (inp[5]) ? 13'b0000000000111 : 13'b0000000001111;
										assign node3825 = (inp[2]) ? node3827 : 13'b0000000001111;
											assign node3827 = (inp[3]) ? 13'b0000000000011 : 13'b0000000000011;
							assign node3830 = (inp[3]) ? node3860 : node3831;
								assign node3831 = (inp[0]) ? node3845 : node3832;
									assign node3832 = (inp[5]) ? node3840 : node3833;
										assign node3833 = (inp[6]) ? node3837 : node3834;
											assign node3834 = (inp[10]) ? 13'b0000000011111 : 13'b0000000111111;
											assign node3837 = (inp[10]) ? 13'b0000000000111 : 13'b0000000011111;
										assign node3840 = (inp[6]) ? node3842 : 13'b0000000001111;
											assign node3842 = (inp[10]) ? 13'b0000000000011 : 13'b0000000001111;
									assign node3845 = (inp[9]) ? node3853 : node3846;
										assign node3846 = (inp[10]) ? node3850 : node3847;
											assign node3847 = (inp[5]) ? 13'b0000000001111 : 13'b0000000001111;
											assign node3850 = (inp[5]) ? 13'b0000000000111 : 13'b0000000001111;
										assign node3853 = (inp[2]) ? node3857 : node3854;
											assign node3854 = (inp[5]) ? 13'b0000000000111 : 13'b0000000001111;
											assign node3857 = (inp[6]) ? 13'b0000000000011 : 13'b0000000000111;
								assign node3860 = (inp[9]) ? node3876 : node3861;
									assign node3861 = (inp[6]) ? node3869 : node3862;
										assign node3862 = (inp[2]) ? node3866 : node3863;
											assign node3863 = (inp[5]) ? 13'b0000000001111 : 13'b0000000011111;
											assign node3866 = (inp[0]) ? 13'b0000000000111 : 13'b0000000001111;
										assign node3869 = (inp[0]) ? node3873 : node3870;
											assign node3870 = (inp[5]) ? 13'b0000000000111 : 13'b0000000000111;
											assign node3873 = (inp[10]) ? 13'b0000000000011 : 13'b0000000000111;
									assign node3876 = (inp[5]) ? node3884 : node3877;
										assign node3877 = (inp[10]) ? node3881 : node3878;
											assign node3878 = (inp[6]) ? 13'b0000000000111 : 13'b0000000000111;
											assign node3881 = (inp[6]) ? 13'b0000000000011 : 13'b0000000000111;
										assign node3884 = (inp[2]) ? node3888 : node3885;
											assign node3885 = (inp[0]) ? 13'b0000000000011 : 13'b0000000000111;
											assign node3888 = (inp[10]) ? 13'b0000000000001 : 13'b0000000000011;

endmodule