module dtc_split75_bm78 (
	input  wire [12-1:0] inp,
	output wire [3-1:0] outp
);

	wire [3-1:0] node1;
	wire [3-1:0] node2;
	wire [3-1:0] node3;
	wire [3-1:0] node4;
	wire [3-1:0] node5;
	wire [3-1:0] node6;
	wire [3-1:0] node7;
	wire [3-1:0] node8;
	wire [3-1:0] node9;
	wire [3-1:0] node11;
	wire [3-1:0] node12;
	wire [3-1:0] node15;
	wire [3-1:0] node18;
	wire [3-1:0] node19;
	wire [3-1:0] node20;
	wire [3-1:0] node25;
	wire [3-1:0] node26;
	wire [3-1:0] node27;
	wire [3-1:0] node30;
	wire [3-1:0] node34;
	wire [3-1:0] node35;
	wire [3-1:0] node36;
	wire [3-1:0] node37;
	wire [3-1:0] node39;
	wire [3-1:0] node42;
	wire [3-1:0] node45;
	wire [3-1:0] node47;
	wire [3-1:0] node49;
	wire [3-1:0] node52;
	wire [3-1:0] node53;
	wire [3-1:0] node54;
	wire [3-1:0] node55;
	wire [3-1:0] node60;
	wire [3-1:0] node62;
	wire [3-1:0] node65;
	wire [3-1:0] node66;
	wire [3-1:0] node67;
	wire [3-1:0] node68;
	wire [3-1:0] node70;
	wire [3-1:0] node73;
	wire [3-1:0] node74;
	wire [3-1:0] node77;
	wire [3-1:0] node80;
	wire [3-1:0] node81;
	wire [3-1:0] node83;
	wire [3-1:0] node84;
	wire [3-1:0] node88;
	wire [3-1:0] node89;
	wire [3-1:0] node91;
	wire [3-1:0] node95;
	wire [3-1:0] node96;
	wire [3-1:0] node97;
	wire [3-1:0] node99;
	wire [3-1:0] node101;
	wire [3-1:0] node104;
	wire [3-1:0] node105;
	wire [3-1:0] node107;
	wire [3-1:0] node111;
	wire [3-1:0] node113;
	wire [3-1:0] node114;
	wire [3-1:0] node117;
	wire [3-1:0] node120;
	wire [3-1:0] node121;
	wire [3-1:0] node122;
	wire [3-1:0] node123;
	wire [3-1:0] node124;
	wire [3-1:0] node125;
	wire [3-1:0] node126;
	wire [3-1:0] node129;
	wire [3-1:0] node132;
	wire [3-1:0] node134;
	wire [3-1:0] node137;
	wire [3-1:0] node138;
	wire [3-1:0] node141;
	wire [3-1:0] node143;
	wire [3-1:0] node146;
	wire [3-1:0] node147;
	wire [3-1:0] node148;
	wire [3-1:0] node151;
	wire [3-1:0] node154;
	wire [3-1:0] node155;
	wire [3-1:0] node157;
	wire [3-1:0] node160;
	wire [3-1:0] node163;
	wire [3-1:0] node164;
	wire [3-1:0] node165;
	wire [3-1:0] node166;
	wire [3-1:0] node167;
	wire [3-1:0] node170;
	wire [3-1:0] node173;
	wire [3-1:0] node174;
	wire [3-1:0] node177;
	wire [3-1:0] node180;
	wire [3-1:0] node182;
	wire [3-1:0] node185;
	wire [3-1:0] node186;
	wire [3-1:0] node187;
	wire [3-1:0] node191;
	wire [3-1:0] node192;
	wire [3-1:0] node195;
	wire [3-1:0] node198;
	wire [3-1:0] node199;
	wire [3-1:0] node200;
	wire [3-1:0] node201;
	wire [3-1:0] node204;
	wire [3-1:0] node205;
	wire [3-1:0] node206;
	wire [3-1:0] node211;
	wire [3-1:0] node212;
	wire [3-1:0] node214;
	wire [3-1:0] node215;
	wire [3-1:0] node219;
	wire [3-1:0] node220;
	wire [3-1:0] node221;
	wire [3-1:0] node225;
	wire [3-1:0] node226;
	wire [3-1:0] node230;
	wire [3-1:0] node231;
	wire [3-1:0] node232;
	wire [3-1:0] node233;
	wire [3-1:0] node235;
	wire [3-1:0] node238;
	wire [3-1:0] node241;
	wire [3-1:0] node242;
	wire [3-1:0] node246;
	wire [3-1:0] node247;
	wire [3-1:0] node248;
	wire [3-1:0] node251;
	wire [3-1:0] node252;
	wire [3-1:0] node256;
	wire [3-1:0] node257;
	wire [3-1:0] node258;
	wire [3-1:0] node262;
	wire [3-1:0] node263;
	wire [3-1:0] node267;
	wire [3-1:0] node268;
	wire [3-1:0] node269;
	wire [3-1:0] node270;
	wire [3-1:0] node271;
	wire [3-1:0] node272;
	wire [3-1:0] node273;
	wire [3-1:0] node274;
	wire [3-1:0] node278;
	wire [3-1:0] node279;
	wire [3-1:0] node283;
	wire [3-1:0] node284;
	wire [3-1:0] node288;
	wire [3-1:0] node289;
	wire [3-1:0] node290;
	wire [3-1:0] node291;
	wire [3-1:0] node297;
	wire [3-1:0] node298;
	wire [3-1:0] node299;
	wire [3-1:0] node301;
	wire [3-1:0] node304;
	wire [3-1:0] node305;
	wire [3-1:0] node308;
	wire [3-1:0] node309;
	wire [3-1:0] node313;
	wire [3-1:0] node314;
	wire [3-1:0] node315;
	wire [3-1:0] node318;
	wire [3-1:0] node321;
	wire [3-1:0] node323;
	wire [3-1:0] node326;
	wire [3-1:0] node327;
	wire [3-1:0] node328;
	wire [3-1:0] node330;
	wire [3-1:0] node332;
	wire [3-1:0] node337;
	wire [3-1:0] node338;
	wire [3-1:0] node339;
	wire [3-1:0] node340;
	wire [3-1:0] node342;
	wire [3-1:0] node345;
	wire [3-1:0] node346;
	wire [3-1:0] node347;
	wire [3-1:0] node350;
	wire [3-1:0] node353;
	wire [3-1:0] node354;
	wire [3-1:0] node358;
	wire [3-1:0] node359;
	wire [3-1:0] node360;
	wire [3-1:0] node361;
	wire [3-1:0] node364;
	wire [3-1:0] node365;
	wire [3-1:0] node371;
	wire [3-1:0] node372;
	wire [3-1:0] node373;
	wire [3-1:0] node374;
	wire [3-1:0] node375;
	wire [3-1:0] node378;
	wire [3-1:0] node379;
	wire [3-1:0] node383;
	wire [3-1:0] node384;
	wire [3-1:0] node385;
	wire [3-1:0] node388;
	wire [3-1:0] node391;
	wire [3-1:0] node392;
	wire [3-1:0] node396;
	wire [3-1:0] node397;
	wire [3-1:0] node398;
	wire [3-1:0] node400;
	wire [3-1:0] node403;
	wire [3-1:0] node404;
	wire [3-1:0] node408;
	wire [3-1:0] node410;
	wire [3-1:0] node411;
	wire [3-1:0] node414;
	wire [3-1:0] node417;
	wire [3-1:0] node418;
	wire [3-1:0] node419;
	wire [3-1:0] node420;
	wire [3-1:0] node421;
	wire [3-1:0] node425;
	wire [3-1:0] node426;
	wire [3-1:0] node431;
	wire [3-1:0] node432;
	wire [3-1:0] node436;
	wire [3-1:0] node437;
	wire [3-1:0] node438;
	wire [3-1:0] node439;
	wire [3-1:0] node440;
	wire [3-1:0] node441;
	wire [3-1:0] node442;
	wire [3-1:0] node445;
	wire [3-1:0] node447;
	wire [3-1:0] node450;
	wire [3-1:0] node451;
	wire [3-1:0] node452;
	wire [3-1:0] node455;
	wire [3-1:0] node458;
	wire [3-1:0] node459;
	wire [3-1:0] node462;
	wire [3-1:0] node464;
	wire [3-1:0] node467;
	wire [3-1:0] node468;
	wire [3-1:0] node469;
	wire [3-1:0] node472;
	wire [3-1:0] node473;
	wire [3-1:0] node476;
	wire [3-1:0] node479;
	wire [3-1:0] node480;
	wire [3-1:0] node481;
	wire [3-1:0] node485;
	wire [3-1:0] node486;
	wire [3-1:0] node487;
	wire [3-1:0] node492;
	wire [3-1:0] node493;
	wire [3-1:0] node494;
	wire [3-1:0] node495;
	wire [3-1:0] node497;
	wire [3-1:0] node500;
	wire [3-1:0] node501;
	wire [3-1:0] node505;
	wire [3-1:0] node506;
	wire [3-1:0] node507;
	wire [3-1:0] node508;
	wire [3-1:0] node514;
	wire [3-1:0] node515;
	wire [3-1:0] node516;
	wire [3-1:0] node517;
	wire [3-1:0] node520;
	wire [3-1:0] node522;
	wire [3-1:0] node525;
	wire [3-1:0] node526;
	wire [3-1:0] node530;
	wire [3-1:0] node532;
	wire [3-1:0] node533;
	wire [3-1:0] node537;
	wire [3-1:0] node538;
	wire [3-1:0] node539;
	wire [3-1:0] node540;
	wire [3-1:0] node541;
	wire [3-1:0] node542;
	wire [3-1:0] node543;
	wire [3-1:0] node546;
	wire [3-1:0] node549;
	wire [3-1:0] node550;
	wire [3-1:0] node556;
	wire [3-1:0] node557;
	wire [3-1:0] node558;
	wire [3-1:0] node559;
	wire [3-1:0] node560;
	wire [3-1:0] node564;
	wire [3-1:0] node565;
	wire [3-1:0] node568;
	wire [3-1:0] node571;
	wire [3-1:0] node573;
	wire [3-1:0] node575;
	wire [3-1:0] node578;
	wire [3-1:0] node579;
	wire [3-1:0] node580;
	wire [3-1:0] node581;
	wire [3-1:0] node585;
	wire [3-1:0] node587;
	wire [3-1:0] node590;
	wire [3-1:0] node591;
	wire [3-1:0] node593;
	wire [3-1:0] node596;
	wire [3-1:0] node597;
	wire [3-1:0] node601;
	wire [3-1:0] node602;
	wire [3-1:0] node603;
	wire [3-1:0] node605;
	wire [3-1:0] node611;
	wire [3-1:0] node612;
	wire [3-1:0] node614;
	wire [3-1:0] node615;
	wire [3-1:0] node616;
	wire [3-1:0] node618;
	wire [3-1:0] node619;
	wire [3-1:0] node620;
	wire [3-1:0] node621;
	wire [3-1:0] node624;
	wire [3-1:0] node626;
	wire [3-1:0] node629;
	wire [3-1:0] node630;
	wire [3-1:0] node633;
	wire [3-1:0] node636;
	wire [3-1:0] node638;
	wire [3-1:0] node640;
	wire [3-1:0] node643;
	wire [3-1:0] node644;
	wire [3-1:0] node645;
	wire [3-1:0] node646;
	wire [3-1:0] node649;
	wire [3-1:0] node650;
	wire [3-1:0] node653;
	wire [3-1:0] node657;
	wire [3-1:0] node658;
	wire [3-1:0] node659;
	wire [3-1:0] node661;
	wire [3-1:0] node662;
	wire [3-1:0] node665;
	wire [3-1:0] node668;
	wire [3-1:0] node671;
	wire [3-1:0] node672;
	wire [3-1:0] node673;
	wire [3-1:0] node675;
	wire [3-1:0] node678;
	wire [3-1:0] node681;
	wire [3-1:0] node682;
	wire [3-1:0] node683;
	wire [3-1:0] node686;
	wire [3-1:0] node689;
	wire [3-1:0] node692;
	wire [3-1:0] node694;
	wire [3-1:0] node695;
	wire [3-1:0] node696;
	wire [3-1:0] node698;
	wire [3-1:0] node700;
	wire [3-1:0] node702;
	wire [3-1:0] node706;
	wire [3-1:0] node708;
	wire [3-1:0] node710;
	wire [3-1:0] node711;
	wire [3-1:0] node715;
	wire [3-1:0] node716;
	wire [3-1:0] node717;
	wire [3-1:0] node718;
	wire [3-1:0] node719;
	wire [3-1:0] node720;
	wire [3-1:0] node721;
	wire [3-1:0] node723;
	wire [3-1:0] node724;
	wire [3-1:0] node727;
	wire [3-1:0] node731;
	wire [3-1:0] node733;
	wire [3-1:0] node736;
	wire [3-1:0] node737;
	wire [3-1:0] node738;
	wire [3-1:0] node739;
	wire [3-1:0] node742;
	wire [3-1:0] node745;
	wire [3-1:0] node746;
	wire [3-1:0] node749;
	wire [3-1:0] node752;
	wire [3-1:0] node753;
	wire [3-1:0] node754;
	wire [3-1:0] node755;
	wire [3-1:0] node759;
	wire [3-1:0] node762;
	wire [3-1:0] node763;
	wire [3-1:0] node766;
	wire [3-1:0] node769;
	wire [3-1:0] node770;
	wire [3-1:0] node771;
	wire [3-1:0] node773;
	wire [3-1:0] node775;
	wire [3-1:0] node778;
	wire [3-1:0] node779;
	wire [3-1:0] node781;
	wire [3-1:0] node785;
	wire [3-1:0] node787;
	wire [3-1:0] node789;
	wire [3-1:0] node791;
	wire [3-1:0] node795;
	wire [3-1:0] node796;
	wire [3-1:0] node797;
	wire [3-1:0] node798;
	wire [3-1:0] node799;
	wire [3-1:0] node800;
	wire [3-1:0] node801;
	wire [3-1:0] node803;
	wire [3-1:0] node806;
	wire [3-1:0] node809;
	wire [3-1:0] node810;
	wire [3-1:0] node813;
	wire [3-1:0] node814;
	wire [3-1:0] node818;
	wire [3-1:0] node820;
	wire [3-1:0] node823;
	wire [3-1:0] node824;
	wire [3-1:0] node825;
	wire [3-1:0] node826;
	wire [3-1:0] node827;
	wire [3-1:0] node832;
	wire [3-1:0] node833;
	wire [3-1:0] node835;
	wire [3-1:0] node839;
	wire [3-1:0] node840;
	wire [3-1:0] node842;
	wire [3-1:0] node845;
	wire [3-1:0] node846;
	wire [3-1:0] node849;
	wire [3-1:0] node852;
	wire [3-1:0] node853;
	wire [3-1:0] node854;
	wire [3-1:0] node855;
	wire [3-1:0] node856;
	wire [3-1:0] node857;
	wire [3-1:0] node861;
	wire [3-1:0] node862;
	wire [3-1:0] node866;
	wire [3-1:0] node867;
	wire [3-1:0] node872;
	wire [3-1:0] node873;
	wire [3-1:0] node874;
	wire [3-1:0] node875;
	wire [3-1:0] node876;
	wire [3-1:0] node880;
	wire [3-1:0] node881;
	wire [3-1:0] node885;
	wire [3-1:0] node886;
	wire [3-1:0] node890;
	wire [3-1:0] node891;
	wire [3-1:0] node893;
	wire [3-1:0] node894;
	wire [3-1:0] node898;
	wire [3-1:0] node899;
	wire [3-1:0] node902;
	wire [3-1:0] node904;
	wire [3-1:0] node907;
	wire [3-1:0] node908;
	wire [3-1:0] node912;
	wire [3-1:0] node913;
	wire [3-1:0] node914;
	wire [3-1:0] node916;
	wire [3-1:0] node917;
	wire [3-1:0] node919;
	wire [3-1:0] node921;
	wire [3-1:0] node926;
	wire [3-1:0] node927;
	wire [3-1:0] node928;
	wire [3-1:0] node929;
	wire [3-1:0] node930;
	wire [3-1:0] node932;
	wire [3-1:0] node933;
	wire [3-1:0] node934;
	wire [3-1:0] node936;
	wire [3-1:0] node939;
	wire [3-1:0] node941;
	wire [3-1:0] node948;
	wire [3-1:0] node949;
	wire [3-1:0] node950;
	wire [3-1:0] node951;
	wire [3-1:0] node952;
	wire [3-1:0] node953;
	wire [3-1:0] node954;
	wire [3-1:0] node956;
	wire [3-1:0] node958;
	wire [3-1:0] node961;
	wire [3-1:0] node962;
	wire [3-1:0] node965;
	wire [3-1:0] node968;
	wire [3-1:0] node969;
	wire [3-1:0] node971;
	wire [3-1:0] node973;
	wire [3-1:0] node976;
	wire [3-1:0] node977;
	wire [3-1:0] node978;
	wire [3-1:0] node982;
	wire [3-1:0] node984;
	wire [3-1:0] node987;
	wire [3-1:0] node989;
	wire [3-1:0] node991;
	wire [3-1:0] node994;
	wire [3-1:0] node995;
	wire [3-1:0] node996;
	wire [3-1:0] node997;
	wire [3-1:0] node999;
	wire [3-1:0] node1000;
	wire [3-1:0] node1003;
	wire [3-1:0] node1006;
	wire [3-1:0] node1007;
	wire [3-1:0] node1010;
	wire [3-1:0] node1013;
	wire [3-1:0] node1014;
	wire [3-1:0] node1015;
	wire [3-1:0] node1017;
	wire [3-1:0] node1020;
	wire [3-1:0] node1022;
	wire [3-1:0] node1025;
	wire [3-1:0] node1027;
	wire [3-1:0] node1029;
	wire [3-1:0] node1032;
	wire [3-1:0] node1033;
	wire [3-1:0] node1034;
	wire [3-1:0] node1036;
	wire [3-1:0] node1039;
	wire [3-1:0] node1040;
	wire [3-1:0] node1041;
	wire [3-1:0] node1046;
	wire [3-1:0] node1047;
	wire [3-1:0] node1048;
	wire [3-1:0] node1051;
	wire [3-1:0] node1054;
	wire [3-1:0] node1055;
	wire [3-1:0] node1059;
	wire [3-1:0] node1060;
	wire [3-1:0] node1061;
	wire [3-1:0] node1062;
	wire [3-1:0] node1063;
	wire [3-1:0] node1065;
	wire [3-1:0] node1066;
	wire [3-1:0] node1070;
	wire [3-1:0] node1071;
	wire [3-1:0] node1072;
	wire [3-1:0] node1076;
	wire [3-1:0] node1078;
	wire [3-1:0] node1081;
	wire [3-1:0] node1082;
	wire [3-1:0] node1083;
	wire [3-1:0] node1084;
	wire [3-1:0] node1089;
	wire [3-1:0] node1090;
	wire [3-1:0] node1092;
	wire [3-1:0] node1096;
	wire [3-1:0] node1097;
	wire [3-1:0] node1098;
	wire [3-1:0] node1100;
	wire [3-1:0] node1103;
	wire [3-1:0] node1104;
	wire [3-1:0] node1106;
	wire [3-1:0] node1110;
	wire [3-1:0] node1112;
	wire [3-1:0] node1113;
	wire [3-1:0] node1114;
	wire [3-1:0] node1119;
	wire [3-1:0] node1120;
	wire [3-1:0] node1121;
	wire [3-1:0] node1122;
	wire [3-1:0] node1123;
	wire [3-1:0] node1128;
	wire [3-1:0] node1129;
	wire [3-1:0] node1130;
	wire [3-1:0] node1131;
	wire [3-1:0] node1135;
	wire [3-1:0] node1137;
	wire [3-1:0] node1140;
	wire [3-1:0] node1141;
	wire [3-1:0] node1146;
	wire [3-1:0] node1148;
	wire [3-1:0] node1149;
	wire [3-1:0] node1150;
	wire [3-1:0] node1151;
	wire [3-1:0] node1153;
	wire [3-1:0] node1155;
	wire [3-1:0] node1158;
	wire [3-1:0] node1159;
	wire [3-1:0] node1161;
	wire [3-1:0] node1164;
	wire [3-1:0] node1166;
	wire [3-1:0] node1170;
	wire [3-1:0] node1171;
	wire [3-1:0] node1172;
	wire [3-1:0] node1173;
	wire [3-1:0] node1175;
	wire [3-1:0] node1178;
	wire [3-1:0] node1179;
	wire [3-1:0] node1182;
	wire [3-1:0] node1183;
	wire [3-1:0] node1188;
	wire [3-1:0] node1189;
	wire [3-1:0] node1191;
	wire [3-1:0] node1193;
	wire [3-1:0] node1196;
	wire [3-1:0] node1197;
	wire [3-1:0] node1200;
	wire [3-1:0] node1201;

	assign outp = (inp[3]) ? node912 : node1;
		assign node1 = (inp[4]) ? node611 : node2;
			assign node2 = (inp[0]) ? node436 : node3;
				assign node3 = (inp[6]) ? node267 : node4;
					assign node4 = (inp[9]) ? node120 : node5;
						assign node5 = (inp[1]) ? node65 : node6;
							assign node6 = (inp[2]) ? node34 : node7;
								assign node7 = (inp[7]) ? node25 : node8;
									assign node8 = (inp[8]) ? node18 : node9;
										assign node9 = (inp[11]) ? node11 : 3'b000;
											assign node11 = (inp[10]) ? node15 : node12;
												assign node12 = (inp[5]) ? 3'b000 : 3'b100;
												assign node15 = (inp[5]) ? 3'b100 : 3'b000;
										assign node18 = (inp[10]) ? 3'b100 : node19;
											assign node19 = (inp[11]) ? 3'b000 : node20;
												assign node20 = (inp[5]) ? 3'b000 : 3'b100;
									assign node25 = (inp[5]) ? 3'b000 : node26;
										assign node26 = (inp[8]) ? node30 : node27;
											assign node27 = (inp[10]) ? 3'b100 : 3'b000;
											assign node30 = (inp[10]) ? 3'b010 : 3'b100;
								assign node34 = (inp[5]) ? node52 : node35;
									assign node35 = (inp[10]) ? node45 : node36;
										assign node36 = (inp[7]) ? node42 : node37;
											assign node37 = (inp[11]) ? node39 : 3'b000;
												assign node39 = (inp[8]) ? 3'b100 : 3'b000;
											assign node42 = (inp[8]) ? 3'b000 : 3'b100;
										assign node45 = (inp[7]) ? node47 : 3'b100;
											assign node47 = (inp[11]) ? node49 : 3'b100;
												assign node49 = (inp[8]) ? 3'b110 : 3'b010;
									assign node52 = (inp[11]) ? node60 : node53;
										assign node53 = (inp[7]) ? 3'b000 : node54;
											assign node54 = (inp[8]) ? 3'b100 : node55;
												assign node55 = (inp[10]) ? 3'b100 : 3'b000;
										assign node60 = (inp[10]) ? node62 : 3'b100;
											assign node62 = (inp[7]) ? 3'b100 : 3'b000;
							assign node65 = (inp[2]) ? node95 : node66;
								assign node66 = (inp[10]) ? node80 : node67;
									assign node67 = (inp[7]) ? node73 : node68;
										assign node68 = (inp[8]) ? node70 : 3'b000;
											assign node70 = (inp[11]) ? 3'b000 : 3'b100;
										assign node73 = (inp[5]) ? node77 : node74;
											assign node74 = (inp[11]) ? 3'b000 : 3'b010;
											assign node77 = (inp[11]) ? 3'b100 : 3'b000;
									assign node80 = (inp[7]) ? node88 : node81;
										assign node81 = (inp[5]) ? node83 : 3'b010;
											assign node83 = (inp[8]) ? 3'b100 : node84;
												assign node84 = (inp[11]) ? 3'b100 : 3'b000;
										assign node88 = (inp[5]) ? 3'b010 : node89;
											assign node89 = (inp[8]) ? node91 : 3'b110;
												assign node91 = (inp[11]) ? 3'b001 : 3'b011;
								assign node95 = (inp[5]) ? node111 : node96;
									assign node96 = (inp[10]) ? node104 : node97;
										assign node97 = (inp[7]) ? node99 : 3'b010;
											assign node99 = (inp[8]) ? node101 : 3'b110;
												assign node101 = (inp[11]) ? 3'b111 : 3'b110;
										assign node104 = (inp[7]) ? 3'b101 : node105;
											assign node105 = (inp[11]) ? node107 : 3'b110;
												assign node107 = (inp[8]) ? 3'b001 : 3'b110;
									assign node111 = (inp[11]) ? node113 : 3'b100;
										assign node113 = (inp[7]) ? node117 : node114;
											assign node114 = (inp[10]) ? 3'b010 : 3'b100;
											assign node117 = (inp[10]) ? 3'b110 : 3'b010;
						assign node120 = (inp[1]) ? node198 : node121;
							assign node121 = (inp[5]) ? node163 : node122;
								assign node122 = (inp[10]) ? node146 : node123;
									assign node123 = (inp[2]) ? node137 : node124;
										assign node124 = (inp[7]) ? node132 : node125;
											assign node125 = (inp[8]) ? node129 : node126;
												assign node126 = (inp[11]) ? 3'b110 : 3'b010;
												assign node129 = (inp[11]) ? 3'b010 : 3'b110;
											assign node132 = (inp[11]) ? node134 : 3'b010;
												assign node134 = (inp[8]) ? 3'b100 : 3'b010;
										assign node137 = (inp[7]) ? node141 : node138;
											assign node138 = (inp[11]) ? 3'b110 : 3'b010;
											assign node141 = (inp[11]) ? node143 : 3'b110;
												assign node143 = (inp[8]) ? 3'b111 : 3'b110;
									assign node146 = (inp[7]) ? node154 : node147;
										assign node147 = (inp[8]) ? node151 : node148;
											assign node148 = (inp[2]) ? 3'b110 : 3'b010;
											assign node151 = (inp[2]) ? 3'b001 : 3'b110;
										assign node154 = (inp[2]) ? node160 : node155;
											assign node155 = (inp[8]) ? node157 : 3'b110;
												assign node157 = (inp[11]) ? 3'b001 : 3'b011;
											assign node160 = (inp[11]) ? 3'b101 : 3'b001;
								assign node163 = (inp[10]) ? node185 : node164;
									assign node164 = (inp[11]) ? node180 : node165;
										assign node165 = (inp[8]) ? node173 : node166;
											assign node166 = (inp[2]) ? node170 : node167;
												assign node167 = (inp[7]) ? 3'b000 : 3'b010;
												assign node170 = (inp[7]) ? 3'b100 : 3'b000;
											assign node173 = (inp[2]) ? node177 : node174;
												assign node174 = (inp[7]) ? 3'b100 : 3'b000;
												assign node177 = (inp[7]) ? 3'b000 : 3'b100;
										assign node180 = (inp[2]) ? node182 : 3'b100;
											assign node182 = (inp[7]) ? 3'b010 : 3'b100;
									assign node185 = (inp[7]) ? node191 : node186;
										assign node186 = (inp[2]) ? 3'b010 : node187;
											assign node187 = (inp[11]) ? 3'b100 : 3'b000;
										assign node191 = (inp[11]) ? node195 : node192;
											assign node192 = (inp[2]) ? 3'b100 : 3'b110;
											assign node195 = (inp[2]) ? 3'b110 : 3'b010;
							assign node198 = (inp[5]) ? node230 : node199;
								assign node199 = (inp[2]) ? node211 : node200;
									assign node200 = (inp[7]) ? node204 : node201;
										assign node201 = (inp[10]) ? 3'b101 : 3'b110;
										assign node204 = (inp[10]) ? 3'b011 : node205;
											assign node205 = (inp[8]) ? 3'b101 : node206;
												assign node206 = (inp[11]) ? 3'b101 : 3'b001;
									assign node211 = (inp[10]) ? node219 : node212;
										assign node212 = (inp[7]) ? node214 : 3'b101;
											assign node214 = (inp[8]) ? 3'b011 : node215;
												assign node215 = (inp[11]) ? 3'b011 : 3'b101;
										assign node219 = (inp[7]) ? node225 : node220;
											assign node220 = (inp[11]) ? 3'b011 : node221;
												assign node221 = (inp[8]) ? 3'b011 : 3'b101;
											assign node225 = (inp[8]) ? 3'b111 : node226;
												assign node226 = (inp[11]) ? 3'b111 : 3'b011;
								assign node230 = (inp[10]) ? node246 : node231;
									assign node231 = (inp[8]) ? node241 : node232;
										assign node232 = (inp[2]) ? node238 : node233;
											assign node233 = (inp[7]) ? node235 : 3'b100;
												assign node235 = (inp[11]) ? 3'b110 : 3'b010;
											assign node238 = (inp[7]) ? 3'b001 : 3'b010;
										assign node241 = (inp[11]) ? 3'b110 : node242;
											assign node242 = (inp[7]) ? 3'b100 : 3'b110;
									assign node246 = (inp[7]) ? node256 : node247;
										assign node247 = (inp[2]) ? node251 : node248;
											assign node248 = (inp[8]) ? 3'b110 : 3'b010;
											assign node251 = (inp[11]) ? 3'b001 : node252;
												assign node252 = (inp[8]) ? 3'b001 : 3'b110;
										assign node256 = (inp[11]) ? node262 : node257;
											assign node257 = (inp[2]) ? 3'b101 : node258;
												assign node258 = (inp[8]) ? 3'b001 : 3'b100;
											assign node262 = (inp[2]) ? 3'b011 : node263;
												assign node263 = (inp[8]) ? 3'b101 : 3'b001;
					assign node267 = (inp[9]) ? node337 : node268;
						assign node268 = (inp[1]) ? node326 : node269;
							assign node269 = (inp[5]) ? node297 : node270;
								assign node270 = (inp[7]) ? node288 : node271;
									assign node271 = (inp[2]) ? node283 : node272;
										assign node272 = (inp[10]) ? node278 : node273;
											assign node273 = (inp[11]) ? 3'b010 : node274;
												assign node274 = (inp[8]) ? 3'b010 : 3'b011;
											assign node278 = (inp[11]) ? 3'b011 : node279;
												assign node279 = (inp[8]) ? 3'b011 : 3'b010;
										assign node283 = (inp[11]) ? 3'b011 : node284;
											assign node284 = (inp[8]) ? 3'b011 : 3'b010;
									assign node288 = (inp[8]) ? 3'b011 : node289;
										assign node289 = (inp[11]) ? 3'b011 : node290;
											assign node290 = (inp[10]) ? 3'b011 : node291;
												assign node291 = (inp[2]) ? 3'b011 : 3'b010;
								assign node297 = (inp[7]) ? node313 : node298;
									assign node298 = (inp[2]) ? node304 : node299;
										assign node299 = (inp[11]) ? node301 : 3'b011;
											assign node301 = (inp[8]) ? 3'b011 : 3'b010;
										assign node304 = (inp[11]) ? node308 : node305;
											assign node305 = (inp[10]) ? 3'b010 : 3'b011;
											assign node308 = (inp[10]) ? 3'b011 : node309;
												assign node309 = (inp[8]) ? 3'b010 : 3'b011;
									assign node313 = (inp[8]) ? node321 : node314;
										assign node314 = (inp[10]) ? node318 : node315;
											assign node315 = (inp[2]) ? 3'b010 : 3'b011;
											assign node318 = (inp[2]) ? 3'b011 : 3'b010;
										assign node321 = (inp[11]) ? node323 : 3'b010;
											assign node323 = (inp[2]) ? 3'b011 : 3'b010;
							assign node326 = (inp[11]) ? 3'b011 : node327;
								assign node327 = (inp[7]) ? 3'b011 : node328;
									assign node328 = (inp[5]) ? node330 : 3'b011;
										assign node330 = (inp[8]) ? node332 : 3'b011;
											assign node332 = (inp[2]) ? 3'b011 : 3'b010;
						assign node337 = (inp[5]) ? node371 : node338;
							assign node338 = (inp[1]) ? node358 : node339;
								assign node339 = (inp[2]) ? node345 : node340;
									assign node340 = (inp[11]) ? node342 : 3'b011;
										assign node342 = (inp[8]) ? 3'b011 : 3'b111;
									assign node345 = (inp[10]) ? node353 : node346;
										assign node346 = (inp[7]) ? node350 : node347;
											assign node347 = (inp[11]) ? 3'b111 : 3'b011;
											assign node350 = (inp[11]) ? 3'b011 : 3'b111;
										assign node353 = (inp[7]) ? 3'b111 : node354;
											assign node354 = (inp[11]) ? 3'b011 : 3'b111;
								assign node358 = (inp[2]) ? 3'b111 : node359;
									assign node359 = (inp[10]) ? 3'b111 : node360;
										assign node360 = (inp[7]) ? node364 : node361;
											assign node361 = (inp[11]) ? 3'b011 : 3'b101;
											assign node364 = (inp[8]) ? 3'b111 : node365;
												assign node365 = (inp[11]) ? 3'b111 : 3'b011;
							assign node371 = (inp[7]) ? node417 : node372;
								assign node372 = (inp[11]) ? node396 : node373;
									assign node373 = (inp[10]) ? node383 : node374;
										assign node374 = (inp[8]) ? node378 : node375;
											assign node375 = (inp[2]) ? 3'b101 : 3'b111;
											assign node378 = (inp[2]) ? 3'b101 : node379;
												assign node379 = (inp[1]) ? 3'b001 : 3'b101;
										assign node383 = (inp[8]) ? node391 : node384;
											assign node384 = (inp[2]) ? node388 : node385;
												assign node385 = (inp[1]) ? 3'b101 : 3'b001;
												assign node388 = (inp[1]) ? 3'b011 : 3'b111;
											assign node391 = (inp[2]) ? 3'b001 : node392;
												assign node392 = (inp[1]) ? 3'b111 : 3'b011;
									assign node396 = (inp[1]) ? node408 : node397;
										assign node397 = (inp[8]) ? node403 : node398;
											assign node398 = (inp[2]) ? node400 : 3'b101;
												assign node400 = (inp[10]) ? 3'b011 : 3'b101;
											assign node403 = (inp[10]) ? 3'b111 : node404;
												assign node404 = (inp[2]) ? 3'b111 : 3'b001;
										assign node408 = (inp[10]) ? node410 : 3'b011;
											assign node410 = (inp[8]) ? node414 : node411;
												assign node411 = (inp[2]) ? 3'b011 : 3'b101;
												assign node414 = (inp[2]) ? 3'b111 : 3'b011;
								assign node417 = (inp[10]) ? node431 : node418;
									assign node418 = (inp[8]) ? 3'b011 : node419;
										assign node419 = (inp[2]) ? node425 : node420;
											assign node420 = (inp[1]) ? 3'b111 : node421;
												assign node421 = (inp[11]) ? 3'b111 : 3'b011;
											assign node425 = (inp[1]) ? 3'b011 : node426;
												assign node426 = (inp[11]) ? 3'b011 : 3'b111;
									assign node431 = (inp[2]) ? 3'b111 : node432;
										assign node432 = (inp[8]) ? 3'b111 : 3'b011;
				assign node436 = (inp[6]) ? 3'b111 : node437;
					assign node437 = (inp[1]) ? node537 : node438;
						assign node438 = (inp[9]) ? node492 : node439;
							assign node439 = (inp[7]) ? node467 : node440;
								assign node440 = (inp[10]) ? node450 : node441;
									assign node441 = (inp[5]) ? node445 : node442;
										assign node442 = (inp[11]) ? 3'b110 : 3'b010;
										assign node445 = (inp[11]) ? node447 : 3'b110;
											assign node447 = (inp[2]) ? 3'b110 : 3'b010;
									assign node450 = (inp[5]) ? node458 : node451;
										assign node451 = (inp[2]) ? node455 : node452;
											assign node452 = (inp[11]) ? 3'b101 : 3'b001;
											assign node455 = (inp[11]) ? 3'b011 : 3'b101;
										assign node458 = (inp[2]) ? node462 : node459;
											assign node459 = (inp[11]) ? 3'b110 : 3'b010;
											assign node462 = (inp[11]) ? node464 : 3'b110;
												assign node464 = (inp[8]) ? 3'b101 : 3'b001;
								assign node467 = (inp[2]) ? node479 : node468;
									assign node468 = (inp[5]) ? node472 : node469;
										assign node469 = (inp[11]) ? 3'b101 : 3'b001;
										assign node472 = (inp[10]) ? node476 : node473;
											assign node473 = (inp[11]) ? 3'b111 : 3'b011;
											assign node476 = (inp[11]) ? 3'b001 : 3'b011;
									assign node479 = (inp[11]) ? node485 : node480;
										assign node480 = (inp[5]) ? 3'b101 : node481;
											assign node481 = (inp[10]) ? 3'b111 : 3'b101;
										assign node485 = (inp[10]) ? 3'b111 : node486;
											assign node486 = (inp[8]) ? 3'b011 : node487;
												assign node487 = (inp[5]) ? 3'b001 : 3'b011;
							assign node492 = (inp[5]) ? node514 : node493;
								assign node493 = (inp[10]) ? node505 : node494;
									assign node494 = (inp[7]) ? node500 : node495;
										assign node495 = (inp[2]) ? node497 : 3'b011;
											assign node497 = (inp[8]) ? 3'b111 : 3'b011;
										assign node500 = (inp[11]) ? 3'b111 : node501;
											assign node501 = (inp[8]) ? 3'b111 : 3'b011;
									assign node505 = (inp[11]) ? 3'b111 : node506;
										assign node506 = (inp[7]) ? 3'b111 : node507;
											assign node507 = (inp[8]) ? 3'b111 : node508;
												assign node508 = (inp[2]) ? 3'b111 : 3'b011;
								assign node514 = (inp[2]) ? node530 : node515;
									assign node515 = (inp[11]) ? node525 : node516;
										assign node516 = (inp[10]) ? node520 : node517;
											assign node517 = (inp[8]) ? 3'b001 : 3'b101;
											assign node520 = (inp[7]) ? node522 : 3'b101;
												assign node522 = (inp[8]) ? 3'b111 : 3'b011;
										assign node525 = (inp[7]) ? 3'b011 : node526;
											assign node526 = (inp[8]) ? 3'b011 : 3'b001;
									assign node530 = (inp[10]) ? node532 : 3'b011;
										assign node532 = (inp[7]) ? 3'b111 : node533;
											assign node533 = (inp[8]) ? 3'b111 : 3'b011;
						assign node537 = (inp[9]) ? node601 : node538;
							assign node538 = (inp[5]) ? node556 : node539;
								assign node539 = (inp[11]) ? 3'b111 : node540;
									assign node540 = (inp[8]) ? 3'b111 : node541;
										assign node541 = (inp[10]) ? node549 : node542;
											assign node542 = (inp[2]) ? node546 : node543;
												assign node543 = (inp[7]) ? 3'b011 : 3'b111;
												assign node546 = (inp[7]) ? 3'b111 : 3'b011;
											assign node549 = (inp[7]) ? 3'b111 : node550;
												assign node550 = (inp[2]) ? 3'b111 : 3'b011;
								assign node556 = (inp[7]) ? node578 : node557;
									assign node557 = (inp[2]) ? node571 : node558;
										assign node558 = (inp[8]) ? node564 : node559;
											assign node559 = (inp[10]) ? 3'b101 : node560;
												assign node560 = (inp[11]) ? 3'b001 : 3'b101;
											assign node564 = (inp[11]) ? node568 : node565;
												assign node565 = (inp[10]) ? 3'b101 : 3'b001;
												assign node568 = (inp[10]) ? 3'b011 : 3'b111;
										assign node571 = (inp[10]) ? node573 : 3'b001;
											assign node573 = (inp[8]) ? node575 : 3'b011;
												assign node575 = (inp[11]) ? 3'b111 : 3'b011;
									assign node578 = (inp[2]) ? node590 : node579;
										assign node579 = (inp[11]) ? node585 : node580;
											assign node580 = (inp[10]) ? 3'b111 : node581;
												assign node581 = (inp[8]) ? 3'b011 : 3'b111;
											assign node585 = (inp[10]) ? node587 : 3'b111;
												assign node587 = (inp[8]) ? 3'b111 : 3'b011;
										assign node590 = (inp[10]) ? node596 : node591;
											assign node591 = (inp[11]) ? node593 : 3'b011;
												assign node593 = (inp[8]) ? 3'b111 : 3'b011;
											assign node596 = (inp[11]) ? 3'b111 : node597;
												assign node597 = (inp[8]) ? 3'b011 : 3'b111;
							assign node601 = (inp[10]) ? 3'b111 : node602;
								assign node602 = (inp[7]) ? 3'b111 : node603;
									assign node603 = (inp[5]) ? node605 : 3'b111;
										assign node605 = (inp[2]) ? 3'b111 : 3'b011;
			assign node611 = (inp[0]) ? node715 : node612;
				assign node612 = (inp[9]) ? node614 : 3'b000;
					assign node614 = (inp[6]) ? node692 : node615;
						assign node615 = (inp[7]) ? node643 : node616;
							assign node616 = (inp[1]) ? node618 : 3'b000;
								assign node618 = (inp[5]) ? node636 : node619;
									assign node619 = (inp[10]) ? node629 : node620;
										assign node620 = (inp[2]) ? node624 : node621;
											assign node621 = (inp[8]) ? 3'b100 : 3'b000;
											assign node624 = (inp[8]) ? node626 : 3'b100;
												assign node626 = (inp[11]) ? 3'b010 : 3'b100;
										assign node629 = (inp[8]) ? node633 : node630;
											assign node630 = (inp[2]) ? 3'b010 : 3'b100;
											assign node633 = (inp[2]) ? 3'b110 : 3'b010;
									assign node636 = (inp[2]) ? node638 : 3'b000;
										assign node638 = (inp[11]) ? node640 : 3'b000;
											assign node640 = (inp[10]) ? 3'b100 : 3'b000;
							assign node643 = (inp[2]) ? node657 : node644;
								assign node644 = (inp[5]) ? 3'b100 : node645;
									assign node645 = (inp[10]) ? node649 : node646;
										assign node646 = (inp[8]) ? 3'b000 : 3'b100;
										assign node649 = (inp[1]) ? node653 : node650;
											assign node650 = (inp[8]) ? 3'b100 : 3'b000;
											assign node653 = (inp[8]) ? 3'b110 : 3'b010;
								assign node657 = (inp[10]) ? node671 : node658;
									assign node658 = (inp[5]) ? node668 : node659;
										assign node659 = (inp[1]) ? node661 : 3'b100;
											assign node661 = (inp[11]) ? node665 : node662;
												assign node662 = (inp[8]) ? 3'b110 : 3'b010;
												assign node665 = (inp[8]) ? 3'b101 : 3'b110;
										assign node668 = (inp[11]) ? 3'b000 : 3'b100;
									assign node671 = (inp[1]) ? node681 : node672;
										assign node672 = (inp[8]) ? node678 : node673;
											assign node673 = (inp[11]) ? node675 : 3'b000;
												assign node675 = (inp[5]) ? 3'b000 : 3'b100;
											assign node678 = (inp[5]) ? 3'b000 : 3'b010;
										assign node681 = (inp[5]) ? node689 : node682;
											assign node682 = (inp[8]) ? node686 : node683;
												assign node683 = (inp[11]) ? 3'b110 : 3'b010;
												assign node686 = (inp[11]) ? 3'b001 : 3'b010;
											assign node689 = (inp[11]) ? 3'b010 : 3'b100;
						assign node692 = (inp[1]) ? node694 : 3'b000;
							assign node694 = (inp[7]) ? node706 : node695;
								assign node695 = (inp[5]) ? 3'b000 : node696;
									assign node696 = (inp[11]) ? node698 : 3'b000;
										assign node698 = (inp[8]) ? node700 : 3'b000;
											assign node700 = (inp[2]) ? node702 : 3'b001;
												assign node702 = (inp[10]) ? 3'b000 : 3'b001;
								assign node706 = (inp[5]) ? node708 : 3'b001;
									assign node708 = (inp[2]) ? node710 : 3'b000;
										assign node710 = (inp[8]) ? 3'b001 : node711;
											assign node711 = (inp[11]) ? 3'b001 : 3'b000;
				assign node715 = (inp[9]) ? node795 : node716;
					assign node716 = (inp[6]) ? 3'b000 : node717;
						assign node717 = (inp[7]) ? node769 : node718;
							assign node718 = (inp[1]) ? node736 : node719;
								assign node719 = (inp[5]) ? node731 : node720;
									assign node720 = (inp[2]) ? 3'b010 : node721;
										assign node721 = (inp[8]) ? node723 : 3'b100;
											assign node723 = (inp[10]) ? node727 : node724;
												assign node724 = (inp[11]) ? 3'b000 : 3'b100;
												assign node727 = (inp[11]) ? 3'b010 : 3'b110;
									assign node731 = (inp[2]) ? node733 : 3'b000;
										assign node733 = (inp[11]) ? 3'b100 : 3'b000;
								assign node736 = (inp[5]) ? node752 : node737;
									assign node737 = (inp[10]) ? node745 : node738;
										assign node738 = (inp[2]) ? node742 : node739;
											assign node739 = (inp[8]) ? 3'b110 : 3'b010;
											assign node742 = (inp[11]) ? 3'b111 : 3'b110;
										assign node745 = (inp[2]) ? node749 : node746;
											assign node746 = (inp[8]) ? 3'b001 : 3'b110;
											assign node749 = (inp[8]) ? 3'b101 : 3'b001;
									assign node752 = (inp[11]) ? node762 : node753;
										assign node753 = (inp[8]) ? node759 : node754;
											assign node754 = (inp[10]) ? 3'b100 : node755;
												assign node755 = (inp[2]) ? 3'b100 : 3'b000;
											assign node759 = (inp[10]) ? 3'b110 : 3'b010;
										assign node762 = (inp[2]) ? node766 : node763;
											assign node763 = (inp[10]) ? 3'b010 : 3'b100;
											assign node766 = (inp[10]) ? 3'b110 : 3'b010;
							assign node769 = (inp[5]) ? node785 : node770;
								assign node770 = (inp[10]) ? node778 : node771;
									assign node771 = (inp[2]) ? node773 : 3'b110;
										assign node773 = (inp[1]) ? node775 : 3'b110;
											assign node775 = (inp[8]) ? 3'b110 : 3'b111;
									assign node778 = (inp[1]) ? 3'b111 : node779;
										assign node779 = (inp[8]) ? node781 : 3'b110;
											assign node781 = (inp[2]) ? 3'b111 : 3'b110;
								assign node785 = (inp[11]) ? node787 : 3'b110;
									assign node787 = (inp[10]) ? node789 : 3'b110;
										assign node789 = (inp[2]) ? node791 : 3'b110;
											assign node791 = (inp[1]) ? 3'b111 : 3'b110;
					assign node795 = (inp[6]) ? node907 : node796;
						assign node796 = (inp[1]) ? node852 : node797;
							assign node797 = (inp[5]) ? node823 : node798;
								assign node798 = (inp[7]) ? node818 : node799;
									assign node799 = (inp[2]) ? node809 : node800;
										assign node800 = (inp[10]) ? node806 : node801;
											assign node801 = (inp[8]) ? node803 : 3'b010;
												assign node803 = (inp[11]) ? 3'b110 : 3'b010;
											assign node806 = (inp[8]) ? 3'b001 : 3'b110;
										assign node809 = (inp[10]) ? node813 : node810;
											assign node810 = (inp[11]) ? 3'b111 : 3'b110;
											assign node813 = (inp[11]) ? 3'b101 : node814;
												assign node814 = (inp[8]) ? 3'b101 : 3'b001;
									assign node818 = (inp[11]) ? node820 : 3'b101;
										assign node820 = (inp[2]) ? 3'b011 : 3'b101;
								assign node823 = (inp[2]) ? node839 : node824;
									assign node824 = (inp[10]) ? node832 : node825;
										assign node825 = (inp[8]) ? 3'b100 : node826;
											assign node826 = (inp[11]) ? 3'b100 : node827;
												assign node827 = (inp[7]) ? 3'b100 : 3'b000;
										assign node832 = (inp[11]) ? 3'b010 : node833;
											assign node833 = (inp[8]) ? node835 : 3'b100;
												assign node835 = (inp[7]) ? 3'b110 : 3'b000;
									assign node839 = (inp[7]) ? node845 : node840;
										assign node840 = (inp[10]) ? node842 : 3'b010;
											assign node842 = (inp[8]) ? 3'b110 : 3'b010;
										assign node845 = (inp[11]) ? node849 : node846;
											assign node846 = (inp[8]) ? 3'b111 : 3'b110;
											assign node849 = (inp[10]) ? 3'b001 : 3'b011;
							assign node852 = (inp[5]) ? node872 : node853;
								assign node853 = (inp[7]) ? 3'b111 : node854;
									assign node854 = (inp[11]) ? node866 : node855;
										assign node855 = (inp[10]) ? node861 : node856;
											assign node856 = (inp[8]) ? 3'b101 : node857;
												assign node857 = (inp[2]) ? 3'b101 : 3'b001;
											assign node861 = (inp[2]) ? 3'b011 : node862;
												assign node862 = (inp[8]) ? 3'b011 : 3'b101;
										assign node866 = (inp[2]) ? 3'b011 : node867;
											assign node867 = (inp[8]) ? 3'b011 : 3'b101;
								assign node872 = (inp[7]) ? node890 : node873;
									assign node873 = (inp[2]) ? node885 : node874;
										assign node874 = (inp[10]) ? node880 : node875;
											assign node875 = (inp[8]) ? 3'b110 : node876;
												assign node876 = (inp[11]) ? 3'b110 : 3'b010;
											assign node880 = (inp[11]) ? 3'b001 : node881;
												assign node881 = (inp[8]) ? 3'b001 : 3'b110;
										assign node885 = (inp[10]) ? 3'b101 : node886;
											assign node886 = (inp[8]) ? 3'b011 : 3'b001;
									assign node890 = (inp[10]) ? node898 : node891;
										assign node891 = (inp[8]) ? node893 : 3'b001;
											assign node893 = (inp[2]) ? 3'b101 : node894;
												assign node894 = (inp[11]) ? 3'b011 : 3'b001;
										assign node898 = (inp[2]) ? node902 : node899;
											assign node899 = (inp[8]) ? 3'b011 : 3'b101;
											assign node902 = (inp[8]) ? node904 : 3'b011;
												assign node904 = (inp[11]) ? 3'b111 : 3'b011;
						assign node907 = (inp[10]) ? 3'b111 : node908;
							assign node908 = (inp[7]) ? 3'b111 : 3'b011;
		assign node912 = (inp[0]) ? node926 : node913;
			assign node913 = (inp[4]) ? 3'b000 : node914;
				assign node914 = (inp[8]) ? node916 : 3'b000;
					assign node916 = (inp[6]) ? 3'b000 : node917;
						assign node917 = (inp[9]) ? node919 : 3'b000;
							assign node919 = (inp[7]) ? node921 : 3'b000;
								assign node921 = (inp[11]) ? 3'b100 : 3'b000;
			assign node926 = (inp[9]) ? node948 : node927;
				assign node927 = (inp[6]) ? 3'b000 : node928;
					assign node928 = (inp[4]) ? 3'b000 : node929;
						assign node929 = (inp[7]) ? 3'b100 : node930;
							assign node930 = (inp[1]) ? node932 : 3'b000;
								assign node932 = (inp[5]) ? 3'b000 : node933;
									assign node933 = (inp[2]) ? node939 : node934;
										assign node934 = (inp[10]) ? node936 : 3'b000;
											assign node936 = (inp[8]) ? 3'b100 : 3'b000;
										assign node939 = (inp[11]) ? node941 : 3'b100;
											assign node941 = (inp[8]) ? 3'b000 : 3'b100;
				assign node948 = (inp[4]) ? node1146 : node949;
					assign node949 = (inp[6]) ? node1059 : node950;
						assign node950 = (inp[1]) ? node994 : node951;
							assign node951 = (inp[5]) ? node987 : node952;
								assign node952 = (inp[2]) ? node968 : node953;
									assign node953 = (inp[7]) ? node961 : node954;
										assign node954 = (inp[8]) ? node956 : 3'b000;
											assign node956 = (inp[11]) ? node958 : 3'b000;
												assign node958 = (inp[10]) ? 3'b100 : 3'b000;
										assign node961 = (inp[8]) ? node965 : node962;
											assign node962 = (inp[10]) ? 3'b100 : 3'b000;
											assign node965 = (inp[10]) ? 3'b010 : 3'b100;
									assign node968 = (inp[11]) ? node976 : node969;
										assign node969 = (inp[8]) ? node971 : 3'b100;
											assign node971 = (inp[7]) ? node973 : 3'b010;
												assign node973 = (inp[10]) ? 3'b100 : 3'b000;
										assign node976 = (inp[7]) ? node982 : node977;
											assign node977 = (inp[10]) ? 3'b010 : node978;
												assign node978 = (inp[8]) ? 3'b100 : 3'b000;
											assign node982 = (inp[10]) ? node984 : 3'b010;
												assign node984 = (inp[8]) ? 3'b110 : 3'b010;
								assign node987 = (inp[2]) ? node989 : 3'b000;
									assign node989 = (inp[7]) ? node991 : 3'b000;
										assign node991 = (inp[11]) ? 3'b100 : 3'b000;
							assign node994 = (inp[5]) ? node1032 : node995;
								assign node995 = (inp[8]) ? node1013 : node996;
									assign node996 = (inp[10]) ? node1006 : node997;
										assign node997 = (inp[11]) ? node999 : 3'b010;
											assign node999 = (inp[7]) ? node1003 : node1000;
												assign node1000 = (inp[2]) ? 3'b010 : 3'b100;
												assign node1003 = (inp[2]) ? 3'b110 : 3'b010;
										assign node1006 = (inp[2]) ? node1010 : node1007;
											assign node1007 = (inp[7]) ? 3'b110 : 3'b010;
											assign node1010 = (inp[7]) ? 3'b101 : 3'b110;
									assign node1013 = (inp[11]) ? node1025 : node1014;
										assign node1014 = (inp[2]) ? node1020 : node1015;
											assign node1015 = (inp[7]) ? node1017 : 3'b010;
												assign node1017 = (inp[10]) ? 3'b011 : 3'b010;
											assign node1020 = (inp[7]) ? node1022 : 3'b010;
												assign node1022 = (inp[10]) ? 3'b101 : 3'b110;
										assign node1025 = (inp[2]) ? node1027 : 3'b100;
											assign node1027 = (inp[7]) ? node1029 : 3'b001;
												assign node1029 = (inp[10]) ? 3'b101 : 3'b111;
								assign node1032 = (inp[11]) ? node1046 : node1033;
									assign node1033 = (inp[2]) ? node1039 : node1034;
										assign node1034 = (inp[10]) ? node1036 : 3'b000;
											assign node1036 = (inp[8]) ? 3'b010 : 3'b000;
										assign node1039 = (inp[7]) ? 3'b100 : node1040;
											assign node1040 = (inp[10]) ? 3'b100 : node1041;
												assign node1041 = (inp[8]) ? 3'b100 : 3'b000;
									assign node1046 = (inp[10]) ? node1054 : node1047;
										assign node1047 = (inp[2]) ? node1051 : node1048;
											assign node1048 = (inp[7]) ? 3'b100 : 3'b000;
											assign node1051 = (inp[7]) ? 3'b010 : 3'b100;
										assign node1054 = (inp[2]) ? 3'b010 : node1055;
											assign node1055 = (inp[7]) ? 3'b010 : 3'b100;
						assign node1059 = (inp[7]) ? node1119 : node1060;
							assign node1060 = (inp[1]) ? node1096 : node1061;
								assign node1061 = (inp[2]) ? node1081 : node1062;
									assign node1062 = (inp[10]) ? node1070 : node1063;
										assign node1063 = (inp[5]) ? node1065 : 3'b010;
											assign node1065 = (inp[11]) ? 3'b010 : node1066;
												assign node1066 = (inp[8]) ? 3'b010 : 3'b011;
										assign node1070 = (inp[11]) ? node1076 : node1071;
											assign node1071 = (inp[8]) ? 3'b011 : node1072;
												assign node1072 = (inp[5]) ? 3'b011 : 3'b010;
											assign node1076 = (inp[8]) ? node1078 : 3'b011;
												assign node1078 = (inp[5]) ? 3'b010 : 3'b011;
									assign node1081 = (inp[5]) ? node1089 : node1082;
										assign node1082 = (inp[8]) ? 3'b011 : node1083;
											assign node1083 = (inp[11]) ? 3'b011 : node1084;
												assign node1084 = (inp[10]) ? 3'b011 : 3'b010;
										assign node1089 = (inp[10]) ? 3'b010 : node1090;
											assign node1090 = (inp[11]) ? node1092 : 3'b011;
												assign node1092 = (inp[8]) ? 3'b010 : 3'b011;
								assign node1096 = (inp[2]) ? node1110 : node1097;
									assign node1097 = (inp[5]) ? node1103 : node1098;
										assign node1098 = (inp[11]) ? node1100 : 3'b001;
											assign node1100 = (inp[8]) ? 3'b011 : 3'b001;
										assign node1103 = (inp[10]) ? 3'b011 : node1104;
											assign node1104 = (inp[8]) ? node1106 : 3'b010;
												assign node1106 = (inp[11]) ? 3'b011 : 3'b010;
									assign node1110 = (inp[11]) ? node1112 : 3'b011;
										assign node1112 = (inp[5]) ? 3'b001 : node1113;
											assign node1113 = (inp[8]) ? 3'b011 : node1114;
												assign node1114 = (inp[10]) ? 3'b011 : 3'b001;
							assign node1119 = (inp[1]) ? 3'b101 : node1120;
								assign node1120 = (inp[5]) ? node1128 : node1121;
									assign node1121 = (inp[10]) ? 3'b101 : node1122;
										assign node1122 = (inp[8]) ? 3'b101 : node1123;
											assign node1123 = (inp[11]) ? 3'b101 : 3'b100;
									assign node1128 = (inp[11]) ? node1140 : node1129;
										assign node1129 = (inp[8]) ? node1135 : node1130;
											assign node1130 = (inp[2]) ? 3'b101 : node1131;
												assign node1131 = (inp[10]) ? 3'b100 : 3'b101;
											assign node1135 = (inp[10]) ? node1137 : 3'b100;
												assign node1137 = (inp[2]) ? 3'b100 : 3'b101;
										assign node1140 = (inp[8]) ? 3'b101 : node1141;
											assign node1141 = (inp[2]) ? 3'b100 : 3'b101;
					assign node1146 = (inp[1]) ? node1148 : 3'b000;
						assign node1148 = (inp[6]) ? node1170 : node1149;
							assign node1149 = (inp[5]) ? 3'b000 : node1150;
								assign node1150 = (inp[7]) ? node1158 : node1151;
									assign node1151 = (inp[11]) ? node1153 : 3'b000;
										assign node1153 = (inp[8]) ? node1155 : 3'b000;
											assign node1155 = (inp[10]) ? 3'b100 : 3'b000;
									assign node1158 = (inp[2]) ? node1164 : node1159;
										assign node1159 = (inp[8]) ? node1161 : 3'b000;
											assign node1161 = (inp[10]) ? 3'b100 : 3'b000;
										assign node1164 = (inp[11]) ? node1166 : 3'b100;
											assign node1166 = (inp[8]) ? 3'b010 : 3'b100;
							assign node1170 = (inp[5]) ? node1188 : node1171;
								assign node1171 = (inp[7]) ? 3'b110 : node1172;
									assign node1172 = (inp[2]) ? node1178 : node1173;
										assign node1173 = (inp[8]) ? node1175 : 3'b100;
											assign node1175 = (inp[11]) ? 3'b010 : 3'b100;
										assign node1178 = (inp[8]) ? node1182 : node1179;
											assign node1179 = (inp[10]) ? 3'b010 : 3'b100;
											assign node1182 = (inp[10]) ? 3'b000 : node1183;
												assign node1183 = (inp[11]) ? 3'b010 : 3'b000;
								assign node1188 = (inp[2]) ? node1196 : node1189;
									assign node1189 = (inp[8]) ? node1191 : 3'b000;
										assign node1191 = (inp[11]) ? node1193 : 3'b000;
											assign node1193 = (inp[7]) ? 3'b100 : 3'b000;
									assign node1196 = (inp[7]) ? node1200 : node1197;
										assign node1197 = (inp[11]) ? 3'b100 : 3'b000;
										assign node1200 = (inp[8]) ? 3'b010 : node1201;
											assign node1201 = (inp[11]) ? 3'b010 : 3'b100;

endmodule