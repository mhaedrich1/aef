module dtc_split125_bm61 (
	input  wire [12-1:0] inp,
	output wire [11-1:0] outp
);

	wire [11-1:0] node1;
	wire [11-1:0] node2;
	wire [11-1:0] node3;
	wire [11-1:0] node4;
	wire [11-1:0] node5;
	wire [11-1:0] node6;
	wire [11-1:0] node7;
	wire [11-1:0] node8;
	wire [11-1:0] node9;
	wire [11-1:0] node14;
	wire [11-1:0] node15;
	wire [11-1:0] node18;
	wire [11-1:0] node19;
	wire [11-1:0] node20;
	wire [11-1:0] node25;
	wire [11-1:0] node26;
	wire [11-1:0] node28;
	wire [11-1:0] node30;
	wire [11-1:0] node33;
	wire [11-1:0] node34;
	wire [11-1:0] node37;
	wire [11-1:0] node39;
	wire [11-1:0] node42;
	wire [11-1:0] node43;
	wire [11-1:0] node44;
	wire [11-1:0] node47;
	wire [11-1:0] node49;
	wire [11-1:0] node51;
	wire [11-1:0] node52;
	wire [11-1:0] node56;
	wire [11-1:0] node57;
	wire [11-1:0] node59;
	wire [11-1:0] node62;
	wire [11-1:0] node65;
	wire [11-1:0] node66;
	wire [11-1:0] node67;
	wire [11-1:0] node68;
	wire [11-1:0] node69;
	wire [11-1:0] node72;
	wire [11-1:0] node75;
	wire [11-1:0] node76;
	wire [11-1:0] node77;
	wire [11-1:0] node80;
	wire [11-1:0] node83;
	wire [11-1:0] node84;
	wire [11-1:0] node85;
	wire [11-1:0] node88;
	wire [11-1:0] node91;
	wire [11-1:0] node94;
	wire [11-1:0] node95;
	wire [11-1:0] node96;
	wire [11-1:0] node97;
	wire [11-1:0] node101;
	wire [11-1:0] node104;
	wire [11-1:0] node105;
	wire [11-1:0] node108;
	wire [11-1:0] node111;
	wire [11-1:0] node112;
	wire [11-1:0] node113;
	wire [11-1:0] node114;
	wire [11-1:0] node116;
	wire [11-1:0] node119;
	wire [11-1:0] node122;
	wire [11-1:0] node125;
	wire [11-1:0] node126;
	wire [11-1:0] node127;
	wire [11-1:0] node130;
	wire [11-1:0] node131;
	wire [11-1:0] node134;
	wire [11-1:0] node137;
	wire [11-1:0] node138;
	wire [11-1:0] node142;
	wire [11-1:0] node143;
	wire [11-1:0] node144;
	wire [11-1:0] node145;
	wire [11-1:0] node146;
	wire [11-1:0] node147;
	wire [11-1:0] node150;
	wire [11-1:0] node153;
	wire [11-1:0] node154;
	wire [11-1:0] node157;
	wire [11-1:0] node158;
	wire [11-1:0] node162;
	wire [11-1:0] node163;
	wire [11-1:0] node164;
	wire [11-1:0] node168;
	wire [11-1:0] node170;
	wire [11-1:0] node171;
	wire [11-1:0] node175;
	wire [11-1:0] node176;
	wire [11-1:0] node177;
	wire [11-1:0] node180;
	wire [11-1:0] node183;
	wire [11-1:0] node184;
	wire [11-1:0] node185;
	wire [11-1:0] node189;
	wire [11-1:0] node190;
	wire [11-1:0] node191;
	wire [11-1:0] node193;
	wire [11-1:0] node197;
	wire [11-1:0] node199;
	wire [11-1:0] node202;
	wire [11-1:0] node203;
	wire [11-1:0] node204;
	wire [11-1:0] node205;
	wire [11-1:0] node206;
	wire [11-1:0] node210;
	wire [11-1:0] node211;
	wire [11-1:0] node214;
	wire [11-1:0] node217;
	wire [11-1:0] node218;
	wire [11-1:0] node221;
	wire [11-1:0] node223;
	wire [11-1:0] node226;
	wire [11-1:0] node227;
	wire [11-1:0] node228;
	wire [11-1:0] node230;
	wire [11-1:0] node233;
	wire [11-1:0] node234;
	wire [11-1:0] node235;
	wire [11-1:0] node236;
	wire [11-1:0] node239;
	wire [11-1:0] node242;
	wire [11-1:0] node243;
	wire [11-1:0] node247;
	wire [11-1:0] node248;
	wire [11-1:0] node252;
	wire [11-1:0] node253;
	wire [11-1:0] node254;
	wire [11-1:0] node255;
	wire [11-1:0] node259;
	wire [11-1:0] node261;
	wire [11-1:0] node264;
	wire [11-1:0] node265;
	wire [11-1:0] node266;
	wire [11-1:0] node270;
	wire [11-1:0] node273;
	wire [11-1:0] node274;
	wire [11-1:0] node275;
	wire [11-1:0] node276;
	wire [11-1:0] node277;
	wire [11-1:0] node278;
	wire [11-1:0] node279;
	wire [11-1:0] node280;
	wire [11-1:0] node283;
	wire [11-1:0] node286;
	wire [11-1:0] node289;
	wire [11-1:0] node292;
	wire [11-1:0] node294;
	wire [11-1:0] node295;
	wire [11-1:0] node298;
	wire [11-1:0] node300;
	wire [11-1:0] node303;
	wire [11-1:0] node304;
	wire [11-1:0] node305;
	wire [11-1:0] node307;
	wire [11-1:0] node310;
	wire [11-1:0] node313;
	wire [11-1:0] node314;
	wire [11-1:0] node316;
	wire [11-1:0] node318;
	wire [11-1:0] node319;
	wire [11-1:0] node323;
	wire [11-1:0] node324;
	wire [11-1:0] node328;
	wire [11-1:0] node329;
	wire [11-1:0] node330;
	wire [11-1:0] node331;
	wire [11-1:0] node332;
	wire [11-1:0] node335;
	wire [11-1:0] node338;
	wire [11-1:0] node341;
	wire [11-1:0] node343;
	wire [11-1:0] node346;
	wire [11-1:0] node347;
	wire [11-1:0] node348;
	wire [11-1:0] node349;
	wire [11-1:0] node353;
	wire [11-1:0] node354;
	wire [11-1:0] node357;
	wire [11-1:0] node360;
	wire [11-1:0] node361;
	wire [11-1:0] node362;
	wire [11-1:0] node365;
	wire [11-1:0] node368;
	wire [11-1:0] node370;
	wire [11-1:0] node373;
	wire [11-1:0] node374;
	wire [11-1:0] node375;
	wire [11-1:0] node376;
	wire [11-1:0] node377;
	wire [11-1:0] node378;
	wire [11-1:0] node381;
	wire [11-1:0] node384;
	wire [11-1:0] node387;
	wire [11-1:0] node388;
	wire [11-1:0] node389;
	wire [11-1:0] node392;
	wire [11-1:0] node395;
	wire [11-1:0] node396;
	wire [11-1:0] node400;
	wire [11-1:0] node401;
	wire [11-1:0] node402;
	wire [11-1:0] node403;
	wire [11-1:0] node406;
	wire [11-1:0] node408;
	wire [11-1:0] node411;
	wire [11-1:0] node412;
	wire [11-1:0] node416;
	wire [11-1:0] node418;
	wire [11-1:0] node419;
	wire [11-1:0] node420;
	wire [11-1:0] node422;
	wire [11-1:0] node426;
	wire [11-1:0] node429;
	wire [11-1:0] node430;
	wire [11-1:0] node431;
	wire [11-1:0] node432;
	wire [11-1:0] node433;
	wire [11-1:0] node436;
	wire [11-1:0] node437;
	wire [11-1:0] node441;
	wire [11-1:0] node442;
	wire [11-1:0] node445;
	wire [11-1:0] node446;
	wire [11-1:0] node450;
	wire [11-1:0] node451;
	wire [11-1:0] node452;
	wire [11-1:0] node454;
	wire [11-1:0] node458;
	wire [11-1:0] node459;
	wire [11-1:0] node460;
	wire [11-1:0] node464;
	wire [11-1:0] node465;
	wire [11-1:0] node469;
	wire [11-1:0] node470;
	wire [11-1:0] node471;
	wire [11-1:0] node474;
	wire [11-1:0] node476;
	wire [11-1:0] node477;
	wire [11-1:0] node481;
	wire [11-1:0] node482;
	wire [11-1:0] node483;
	wire [11-1:0] node484;
	wire [11-1:0] node487;
	wire [11-1:0] node488;
	wire [11-1:0] node492;
	wire [11-1:0] node494;
	wire [11-1:0] node497;
	wire [11-1:0] node499;
	wire [11-1:0] node500;
	wire [11-1:0] node503;
	wire [11-1:0] node506;
	wire [11-1:0] node507;
	wire [11-1:0] node508;
	wire [11-1:0] node509;
	wire [11-1:0] node510;
	wire [11-1:0] node511;
	wire [11-1:0] node512;
	wire [11-1:0] node514;
	wire [11-1:0] node516;
	wire [11-1:0] node519;
	wire [11-1:0] node521;
	wire [11-1:0] node522;
	wire [11-1:0] node523;
	wire [11-1:0] node526;
	wire [11-1:0] node527;
	wire [11-1:0] node532;
	wire [11-1:0] node534;
	wire [11-1:0] node535;
	wire [11-1:0] node539;
	wire [11-1:0] node540;
	wire [11-1:0] node541;
	wire [11-1:0] node542;
	wire [11-1:0] node546;
	wire [11-1:0] node549;
	wire [11-1:0] node550;
	wire [11-1:0] node551;
	wire [11-1:0] node552;
	wire [11-1:0] node555;
	wire [11-1:0] node559;
	wire [11-1:0] node561;
	wire [11-1:0] node562;
	wire [11-1:0] node566;
	wire [11-1:0] node567;
	wire [11-1:0] node568;
	wire [11-1:0] node569;
	wire [11-1:0] node571;
	wire [11-1:0] node572;
	wire [11-1:0] node575;
	wire [11-1:0] node578;
	wire [11-1:0] node579;
	wire [11-1:0] node581;
	wire [11-1:0] node584;
	wire [11-1:0] node587;
	wire [11-1:0] node588;
	wire [11-1:0] node590;
	wire [11-1:0] node593;
	wire [11-1:0] node594;
	wire [11-1:0] node598;
	wire [11-1:0] node599;
	wire [11-1:0] node600;
	wire [11-1:0] node601;
	wire [11-1:0] node602;
	wire [11-1:0] node605;
	wire [11-1:0] node606;
	wire [11-1:0] node611;
	wire [11-1:0] node612;
	wire [11-1:0] node615;
	wire [11-1:0] node616;
	wire [11-1:0] node617;
	wire [11-1:0] node621;
	wire [11-1:0] node624;
	wire [11-1:0] node625;
	wire [11-1:0] node628;
	wire [11-1:0] node629;
	wire [11-1:0] node632;
	wire [11-1:0] node634;
	wire [11-1:0] node637;
	wire [11-1:0] node638;
	wire [11-1:0] node639;
	wire [11-1:0] node640;
	wire [11-1:0] node641;
	wire [11-1:0] node643;
	wire [11-1:0] node644;
	wire [11-1:0] node648;
	wire [11-1:0] node649;
	wire [11-1:0] node653;
	wire [11-1:0] node654;
	wire [11-1:0] node655;
	wire [11-1:0] node657;
	wire [11-1:0] node660;
	wire [11-1:0] node664;
	wire [11-1:0] node665;
	wire [11-1:0] node667;
	wire [11-1:0] node669;
	wire [11-1:0] node672;
	wire [11-1:0] node673;
	wire [11-1:0] node674;
	wire [11-1:0] node677;
	wire [11-1:0] node680;
	wire [11-1:0] node682;
	wire [11-1:0] node685;
	wire [11-1:0] node686;
	wire [11-1:0] node687;
	wire [11-1:0] node688;
	wire [11-1:0] node689;
	wire [11-1:0] node693;
	wire [11-1:0] node694;
	wire [11-1:0] node698;
	wire [11-1:0] node699;
	wire [11-1:0] node700;
	wire [11-1:0] node701;
	wire [11-1:0] node705;
	wire [11-1:0] node708;
	wire [11-1:0] node709;
	wire [11-1:0] node712;
	wire [11-1:0] node715;
	wire [11-1:0] node716;
	wire [11-1:0] node717;
	wire [11-1:0] node718;
	wire [11-1:0] node722;
	wire [11-1:0] node724;
	wire [11-1:0] node726;
	wire [11-1:0] node729;
	wire [11-1:0] node730;
	wire [11-1:0] node731;
	wire [11-1:0] node733;
	wire [11-1:0] node737;
	wire [11-1:0] node739;
	wire [11-1:0] node741;
	wire [11-1:0] node743;
	wire [11-1:0] node746;
	wire [11-1:0] node747;
	wire [11-1:0] node748;
	wire [11-1:0] node749;
	wire [11-1:0] node750;
	wire [11-1:0] node751;
	wire [11-1:0] node752;
	wire [11-1:0] node756;
	wire [11-1:0] node759;
	wire [11-1:0] node760;
	wire [11-1:0] node762;
	wire [11-1:0] node764;
	wire [11-1:0] node768;
	wire [11-1:0] node769;
	wire [11-1:0] node770;
	wire [11-1:0] node771;
	wire [11-1:0] node772;
	wire [11-1:0] node773;
	wire [11-1:0] node774;
	wire [11-1:0] node781;
	wire [11-1:0] node782;
	wire [11-1:0] node783;
	wire [11-1:0] node784;
	wire [11-1:0] node787;
	wire [11-1:0] node791;
	wire [11-1:0] node793;
	wire [11-1:0] node796;
	wire [11-1:0] node797;
	wire [11-1:0] node799;
	wire [11-1:0] node800;
	wire [11-1:0] node804;
	wire [11-1:0] node805;
	wire [11-1:0] node806;
	wire [11-1:0] node809;
	wire [11-1:0] node812;
	wire [11-1:0] node815;
	wire [11-1:0] node816;
	wire [11-1:0] node817;
	wire [11-1:0] node818;
	wire [11-1:0] node819;
	wire [11-1:0] node822;
	wire [11-1:0] node825;
	wire [11-1:0] node828;
	wire [11-1:0] node829;
	wire [11-1:0] node831;
	wire [11-1:0] node832;
	wire [11-1:0] node835;
	wire [11-1:0] node838;
	wire [11-1:0] node841;
	wire [11-1:0] node842;
	wire [11-1:0] node843;
	wire [11-1:0] node846;
	wire [11-1:0] node847;
	wire [11-1:0] node848;
	wire [11-1:0] node852;
	wire [11-1:0] node855;
	wire [11-1:0] node856;
	wire [11-1:0] node857;
	wire [11-1:0] node858;
	wire [11-1:0] node862;
	wire [11-1:0] node864;
	wire [11-1:0] node867;
	wire [11-1:0] node869;
	wire [11-1:0] node870;
	wire [11-1:0] node874;
	wire [11-1:0] node875;
	wire [11-1:0] node876;
	wire [11-1:0] node877;
	wire [11-1:0] node878;
	wire [11-1:0] node879;
	wire [11-1:0] node881;
	wire [11-1:0] node882;
	wire [11-1:0] node885;
	wire [11-1:0] node888;
	wire [11-1:0] node891;
	wire [11-1:0] node893;
	wire [11-1:0] node896;
	wire [11-1:0] node897;
	wire [11-1:0] node898;
	wire [11-1:0] node899;
	wire [11-1:0] node900;
	wire [11-1:0] node904;
	wire [11-1:0] node907;
	wire [11-1:0] node908;
	wire [11-1:0] node911;
	wire [11-1:0] node914;
	wire [11-1:0] node916;
	wire [11-1:0] node919;
	wire [11-1:0] node920;
	wire [11-1:0] node921;
	wire [11-1:0] node922;
	wire [11-1:0] node923;
	wire [11-1:0] node924;
	wire [11-1:0] node928;
	wire [11-1:0] node931;
	wire [11-1:0] node932;
	wire [11-1:0] node936;
	wire [11-1:0] node937;
	wire [11-1:0] node940;
	wire [11-1:0] node943;
	wire [11-1:0] node944;
	wire [11-1:0] node945;
	wire [11-1:0] node946;
	wire [11-1:0] node947;
	wire [11-1:0] node951;
	wire [11-1:0] node954;
	wire [11-1:0] node955;
	wire [11-1:0] node959;
	wire [11-1:0] node960;
	wire [11-1:0] node963;
	wire [11-1:0] node966;
	wire [11-1:0] node967;
	wire [11-1:0] node968;
	wire [11-1:0] node969;
	wire [11-1:0] node971;
	wire [11-1:0] node974;
	wire [11-1:0] node976;
	wire [11-1:0] node978;
	wire [11-1:0] node981;
	wire [11-1:0] node982;
	wire [11-1:0] node983;
	wire [11-1:0] node987;
	wire [11-1:0] node989;
	wire [11-1:0] node990;
	wire [11-1:0] node994;
	wire [11-1:0] node995;
	wire [11-1:0] node996;
	wire [11-1:0] node997;
	wire [11-1:0] node1000;
	wire [11-1:0] node1003;
	wire [11-1:0] node1006;
	wire [11-1:0] node1007;
	wire [11-1:0] node1009;
	wire [11-1:0] node1011;
	wire [11-1:0] node1014;
	wire [11-1:0] node1016;
	wire [11-1:0] node1018;

	assign outp = (inp[1]) ? node506 : node1;
		assign node1 = (inp[7]) ? node273 : node2;
			assign node2 = (inp[2]) ? node142 : node3;
				assign node3 = (inp[0]) ? node65 : node4;
					assign node4 = (inp[6]) ? node42 : node5;
						assign node5 = (inp[5]) ? node25 : node6;
							assign node6 = (inp[4]) ? node14 : node7;
								assign node7 = (inp[8]) ? 11'b11111101111 : node8;
									assign node8 = (inp[10]) ? 11'b11000101011 : node9;
										assign node9 = (inp[3]) ? 11'b11001101111 : 11'b01001101011;
								assign node14 = (inp[11]) ? node18 : node15;
									assign node15 = (inp[8]) ? 11'b01010001011 : 11'b11100001011;
									assign node18 = (inp[9]) ? 11'b01000011111 : node19;
										assign node19 = (inp[10]) ? 11'b11111011101 : node20;
											assign node20 = (inp[8]) ? 11'b01110101101 : 11'b11111001111;
							assign node25 = (inp[9]) ? node33 : node26;
								assign node26 = (inp[10]) ? node28 : 11'b01000011011;
									assign node28 = (inp[3]) ? node30 : 11'b11010011010;
										assign node30 = (inp[8]) ? 11'b01001011000 : 11'b01010011010;
								assign node33 = (inp[10]) ? node37 : node34;
									assign node34 = (inp[3]) ? 11'b11100111110 : 11'b01111011110;
									assign node37 = (inp[11]) ? node39 : 11'b01101101100;
										assign node39 = (inp[8]) ? 11'b11110001000 : 11'b01110001000;
						assign node42 = (inp[5]) ? node56 : node43;
							assign node43 = (inp[11]) ? node47 : node44;
								assign node44 = (inp[8]) ? 11'b11100001100 : 11'b11011100100;
								assign node47 = (inp[9]) ? node49 : 11'b01001111101;
									assign node49 = (inp[10]) ? node51 : 11'b01111111001;
										assign node51 = (inp[4]) ? 11'b11111111001 : node52;
											assign node52 = (inp[8]) ? 11'b11011011100 : 11'b11110111101;
							assign node56 = (inp[3]) ? node62 : node57;
								assign node57 = (inp[10]) ? node59 : 11'b01010101001;
									assign node59 = (inp[11]) ? 11'b11110101101 : 11'b11010101111;
								assign node62 = (inp[4]) ? 11'b11100111101 : 11'b01110011101;
					assign node65 = (inp[5]) ? node111 : node66;
						assign node66 = (inp[3]) ? node94 : node67;
							assign node67 = (inp[9]) ? node75 : node68;
								assign node68 = (inp[10]) ? node72 : node69;
									assign node69 = (inp[4]) ? 11'b01110111011 : 11'b01100011011;
									assign node72 = (inp[6]) ? 11'b01100101111 : 11'b01001001101;
								assign node75 = (inp[10]) ? node83 : node76;
									assign node76 = (inp[11]) ? node80 : node77;
										assign node77 = (inp[4]) ? 11'b01101011101 : 11'b01110101101;
										assign node80 = (inp[4]) ? 11'b01011001101 : 11'b01011011100;
									assign node83 = (inp[8]) ? node91 : node84;
										assign node84 = (inp[4]) ? node88 : node85;
											assign node85 = (inp[11]) ? 11'b01000101001 : 11'b01000111001;
											assign node88 = (inp[6]) ? 11'b01100001001 : 11'b01110001001;
										assign node91 = (inp[6]) ? 11'b01101011000 : 11'b01111111001;
							assign node94 = (inp[4]) ? node104 : node95;
								assign node95 = (inp[11]) ? node101 : node96;
									assign node96 = (inp[8]) ? 11'b01001001000 : node97;
										assign node97 = (inp[10]) ? 11'b01000100010 : 11'b01001100000;
									assign node101 = (inp[9]) ? 11'b01010101011 : 11'b01001101001;
								assign node104 = (inp[10]) ? node108 : node105;
									assign node105 = (inp[6]) ? 11'b01111011000 : 11'b01001011001;
									assign node108 = (inp[8]) ? 11'b01110001001 : 11'b01000001001;
						assign node111 = (inp[6]) ? node125 : node112;
							assign node112 = (inp[10]) ? node122 : node113;
								assign node113 = (inp[8]) ? node119 : node114;
									assign node114 = (inp[3]) ? node116 : 11'b01111111110;
										assign node116 = (inp[9]) ? 11'b01001001010 : 11'b01001011010;
									assign node119 = (inp[3]) ? 11'b01110111010 : 11'b01010101010;
								assign node122 = (inp[11]) ? 11'b01100001110 : 11'b01101011110;
							assign node125 = (inp[3]) ? node137 : node126;
								assign node126 = (inp[4]) ? node130 : node127;
									assign node127 = (inp[11]) ? 11'b01101011101 : 11'b01011001001;
									assign node130 = (inp[11]) ? node134 : node131;
										assign node131 = (inp[10]) ? 11'b01001111111 : 11'b01100101011;
										assign node134 = (inp[10]) ? 11'b01110101100 : 11'b01101101110;
								assign node137 = (inp[8]) ? 11'b01100001001 : node138;
									assign node138 = (inp[10]) ? 11'b01110101011 : 11'b01100001011;
				assign node142 = (inp[0]) ? node202 : node143;
					assign node143 = (inp[5]) ? node175 : node144;
						assign node144 = (inp[10]) ? node162 : node145;
							assign node145 = (inp[3]) ? node153 : node146;
								assign node146 = (inp[4]) ? node150 : node147;
									assign node147 = (inp[8]) ? 11'b01001010011 : 11'b01111001010;
									assign node150 = (inp[8]) ? 11'b01111110110 : 11'b01110100101;
								assign node153 = (inp[11]) ? node157 : node154;
									assign node154 = (inp[4]) ? 11'b11110000100 : 11'b11011000010;
									assign node157 = (inp[4]) ? 11'b11101000101 : node158;
										assign node158 = (inp[6]) ? 11'b11000000101 : 11'b11010110001;
							assign node162 = (inp[6]) ? node168 : node163;
								assign node163 = (inp[11]) ? 11'b11000100001 : node164;
									assign node164 = (inp[8]) ? 11'b01101100011 : 11'b01000100001;
								assign node168 = (inp[8]) ? node170 : 11'b01000111010;
									assign node170 = (inp[11]) ? 11'b11101110110 : node171;
										assign node171 = (inp[9]) ? 11'b11110000011 : 11'b11000110111;
						assign node175 = (inp[9]) ? node183 : node176;
							assign node176 = (inp[3]) ? node180 : node177;
								assign node177 = (inp[10]) ? 11'b11110001110 : 11'b01001010110;
								assign node180 = (inp[10]) ? 11'b01111110010 : 11'b11110100010;
							assign node183 = (inp[11]) ? node189 : node184;
								assign node184 = (inp[3]) ? 11'b11101010101 : node185;
									assign node185 = (inp[10]) ? 11'b11010110000 : 11'b01110110001;
								assign node189 = (inp[6]) ? node197 : node190;
									assign node190 = (inp[4]) ? 11'b11001100000 : node191;
										assign node191 = (inp[10]) ? node193 : 11'b01011000000;
											assign node193 = (inp[3]) ? 11'b01011000100 : 11'b11010000110;
									assign node197 = (inp[4]) ? node199 : 11'b11110110101;
										assign node199 = (inp[10]) ? 11'b01010000000 : 11'b11010000010;
					assign node202 = (inp[6]) ? node226 : node203;
						assign node203 = (inp[10]) ? node217 : node204;
							assign node204 = (inp[5]) ? node210 : node205;
								assign node205 = (inp[3]) ? 11'b01100010011 : node206;
									assign node206 = (inp[9]) ? 11'b01101010111 : 11'b01001100011;
								assign node210 = (inp[9]) ? node214 : node211;
									assign node211 = (inp[4]) ? 11'b01110100010 : 11'b01110000010;
									assign node214 = (inp[3]) ? 11'b01111010011 : 11'b01010000111;
							assign node217 = (inp[3]) ? node221 : node218;
								assign node218 = (inp[9]) ? 11'b01111000001 : 11'b01010110100;
								assign node221 = (inp[8]) ? node223 : 11'b01010100011;
									assign node223 = (inp[11]) ? 11'b01001100011 : 11'b01010100011;
						assign node226 = (inp[8]) ? node252 : node227;
							assign node227 = (inp[5]) ? node233 : node228;
								assign node228 = (inp[9]) ? node230 : 11'b01111101100;
									assign node230 = (inp[3]) ? 11'b01101101010 : 11'b01101101000;
								assign node233 = (inp[11]) ? node247 : node234;
									assign node234 = (inp[9]) ? node242 : node235;
										assign node235 = (inp[3]) ? node239 : node236;
											assign node236 = (inp[4]) ? 11'b01101001000 : 11'b01101001110;
											assign node239 = (inp[10]) ? 11'b01001001000 : 11'b01101011000;
										assign node242 = (inp[4]) ? 11'b01111110111 : node243;
											assign node243 = (inp[3]) ? 11'b01110011000 : 11'b01110011010;
									assign node247 = (inp[10]) ? 11'b01110000111 : node248;
										assign node248 = (inp[3]) ? 11'b01010010011 : 11'b01111010001;
							assign node252 = (inp[4]) ? node264 : node253;
								assign node253 = (inp[11]) ? node259 : node254;
									assign node254 = (inp[9]) ? 11'b01110000100 : node255;
										assign node255 = (inp[5]) ? 11'b01111000000 : 11'b01110000001;
									assign node259 = (inp[5]) ? node261 : 11'b01111100000;
										assign node261 = (inp[9]) ? 11'b01001000010 : 11'b01101100010;
								assign node264 = (inp[5]) ? node270 : node265;
									assign node265 = (inp[11]) ? 11'b01100110010 : node266;
										assign node266 = (inp[9]) ? 11'b01000010001 : 11'b01010110001;
									assign node270 = (inp[11]) ? 11'b01001000110 : 11'b01001110100;
			assign node273 = (inp[6]) ? node373 : node274;
				assign node274 = (inp[2]) ? node328 : node275;
					assign node275 = (inp[5]) ? node303 : node276;
						assign node276 = (inp[10]) ? node292 : node277;
							assign node277 = (inp[0]) ? node289 : node278;
								assign node278 = (inp[9]) ? node286 : node279;
									assign node279 = (inp[8]) ? node283 : node280;
										assign node280 = (inp[3]) ? 11'b11100100101 : 11'b01010100111;
										assign node283 = (inp[4]) ? 11'b01111100110 : 11'b11111100010;
									assign node286 = (inp[4]) ? 11'b01100100100 : 11'b11100100100;
								assign node289 = (inp[9]) ? 11'b01010110010 : 11'b01100010010;
							assign node292 = (inp[3]) ? node294 : 11'b01001010000;
								assign node294 = (inp[11]) ? node298 : node295;
									assign node295 = (inp[0]) ? 11'b01000100001 : 11'b01000100010;
									assign node298 = (inp[8]) ? node300 : 11'b01011100001;
										assign node300 = (inp[9]) ? 11'b00001101001 : 11'b00000101001;
						assign node303 = (inp[8]) ? node313 : node304;
							assign node304 = (inp[11]) ? node310 : node305;
								assign node305 = (inp[4]) ? node307 : 11'b01011010011;
									assign node307 = (inp[0]) ? 11'b01010010101 : 11'b01001010101;
								assign node310 = (inp[10]) ? 11'b11010000110 : 11'b01010110000;
							assign node313 = (inp[4]) ? node323 : node314;
								assign node314 = (inp[0]) ? node316 : 11'b10000111001;
									assign node316 = (inp[10]) ? node318 : 11'b00100101011;
										assign node318 = (inp[3]) ? 11'b00000101011 : node319;
											assign node319 = (inp[11]) ? 11'b00011101001 : 11'b00010101101;
								assign node323 = (inp[10]) ? 11'b00101001001 : node324;
									assign node324 = (inp[9]) ? 11'b00110011101 : 11'b10110111101;
					assign node328 = (inp[4]) ? node346 : node329;
						assign node329 = (inp[0]) ? node341 : node330;
							assign node330 = (inp[9]) ? node338 : node331;
								assign node331 = (inp[3]) ? node335 : node332;
									assign node332 = (inp[8]) ? 11'b00111101001 : 11'b10101001000;
									assign node335 = (inp[11]) ? 11'b00111011110 : 11'b00001011101;
								assign node338 = (inp[8]) ? 11'b10110011111 : 11'b10110001101;
							assign node341 = (inp[9]) ? node343 : 11'b00110111011;
								assign node343 = (inp[8]) ? 11'b00010001010 : 11'b00100111010;
						assign node346 = (inp[10]) ? node360 : node347;
							assign node347 = (inp[0]) ? node353 : node348;
								assign node348 = (inp[3]) ? 11'b10000011100 : node349;
									assign node349 = (inp[9]) ? 11'b00000111100 : 11'b00001111110;
								assign node353 = (inp[9]) ? node357 : node354;
									assign node354 = (inp[11]) ? 11'b00100111001 : 11'b00000101010;
									assign node357 = (inp[3]) ? 11'b00111101000 : 11'b00101111100;
							assign node360 = (inp[5]) ? node368 : node361;
								assign node361 = (inp[8]) ? node365 : node362;
									assign node362 = (inp[3]) ? 11'b00001111010 : 11'b10001111000;
									assign node365 = (inp[3]) ? 11'b00001101011 : 11'b00011111001;
								assign node368 = (inp[0]) ? node370 : 11'b10110101011;
									assign node370 = (inp[3]) ? 11'b00001001010 : 11'b00010001010;
				assign node373 = (inp[8]) ? node429 : node374;
					assign node374 = (inp[0]) ? node400 : node375;
						assign node375 = (inp[5]) ? node387 : node376;
							assign node376 = (inp[2]) ? node384 : node377;
								assign node377 = (inp[3]) ? node381 : node378;
									assign node378 = (inp[4]) ? 11'b10010111100 : 11'b10011101000;
									assign node381 = (inp[9]) ? 11'b00001111100 : 11'b00000101110;
								assign node384 = (inp[4]) ? 11'b10010110001 : 11'b10011010101;
							assign node387 = (inp[4]) ? node395 : node388;
								assign node388 = (inp[3]) ? node392 : node389;
									assign node389 = (inp[9]) ? 11'b00101110011 : 11'b00100110001;
									assign node392 = (inp[10]) ? 11'b00101110101 : 11'b10001110001;
								assign node395 = (inp[9]) ? 11'b10000000001 : node396;
									assign node396 = (inp[2]) ? 11'b00110010111 : 11'b10010000111;
						assign node400 = (inp[2]) ? node416 : node401;
							assign node401 = (inp[5]) ? node411 : node402;
								assign node402 = (inp[10]) ? node406 : node403;
									assign node403 = (inp[9]) ? 11'b00001100101 : 11'b00000011010;
									assign node406 = (inp[11]) ? node408 : 11'b00001001000;
										assign node408 = (inp[9]) ? 11'b00000001010 : 11'b00101001010;
								assign node411 = (inp[11]) ? 11'b00000100001 : node412;
									assign node412 = (inp[3]) ? 11'b00110000011 : 11'b00111100101;
							assign node416 = (inp[3]) ? node418 : 11'b00010000100;
								assign node418 = (inp[5]) ? node426 : node419;
									assign node419 = (inp[11]) ? 11'b00101000001 : node420;
										assign node420 = (inp[10]) ? node422 : 11'b00110100001;
											assign node422 = (inp[9]) ? 11'b00001100001 : 11'b00100100001;
									assign node426 = (inp[9]) ? 11'b00000000001 : 11'b00010010001;
					assign node429 = (inp[5]) ? node469 : node430;
						assign node430 = (inp[10]) ? node450 : node431;
							assign node431 = (inp[2]) ? node441 : node432;
								assign node432 = (inp[11]) ? node436 : node433;
									assign node433 = (inp[9]) ? 11'b00010010001 : 11'b00110100001;
									assign node436 = (inp[9]) ? 11'b00110110010 : node437;
										assign node437 = (inp[4]) ? 11'b00110110010 : 11'b00111110010;
								assign node441 = (inp[3]) ? node445 : node442;
									assign node442 = (inp[0]) ? 11'b00011110100 : 11'b00011010000;
									assign node445 = (inp[9]) ? 11'b00100100010 : node446;
										assign node446 = (inp[0]) ? 11'b00011110010 : 11'b10111100110;
							assign node450 = (inp[11]) ? node458 : node451;
								assign node451 = (inp[9]) ? 11'b00001100010 : node452;
									assign node452 = (inp[3]) ? node454 : 11'b00111000101;
										assign node454 = (inp[4]) ? 11'b00011000001 : 11'b00011000011;
								assign node458 = (inp[0]) ? node464 : node459;
									assign node459 = (inp[4]) ? 11'b00101010010 : node460;
										assign node460 = (inp[3]) ? 11'b00111110100 : 11'b10101100000;
									assign node464 = (inp[4]) ? 11'b00010100100 : node465;
										assign node465 = (inp[3]) ? 11'b00011100010 : 11'b00110000010;
						assign node469 = (inp[11]) ? node481 : node470;
							assign node470 = (inp[3]) ? node474 : node471;
								assign node471 = (inp[0]) ? 11'b00011100110 : 11'b10011110010;
								assign node474 = (inp[2]) ? node476 : 11'b00110010100;
									assign node476 = (inp[0]) ? 11'b00101110000 : node477;
										assign node477 = (inp[4]) ? 11'b10101110100 : 11'b10111110000;
							assign node481 = (inp[3]) ? node497 : node482;
								assign node482 = (inp[10]) ? node492 : node483;
									assign node483 = (inp[2]) ? node487 : node484;
										assign node484 = (inp[0]) ? 11'b00011110100 : 11'b00001100010;
										assign node487 = (inp[9]) ? 11'b00000010110 : node488;
											assign node488 = (inp[4]) ? 11'b00001010010 : 11'b00101010010;
									assign node492 = (inp[9]) ? node494 : 11'b00001000110;
										assign node494 = (inp[2]) ? 11'b00000000010 : 11'b10100000010;
								assign node497 = (inp[9]) ? node499 : 11'b00101000000;
									assign node499 = (inp[2]) ? node503 : node500;
										assign node500 = (inp[10]) ? 11'b00000000000 : 11'b10110000000;
										assign node503 = (inp[10]) ? 11'b00000000100 : 11'b00000010000;
		assign node506 = (inp[7]) ? node746 : node507;
			assign node507 = (inp[6]) ? node637 : node508;
				assign node508 = (inp[8]) ? node566 : node509;
					assign node509 = (inp[3]) ? node539 : node510;
						assign node510 = (inp[9]) ? node532 : node511;
							assign node511 = (inp[10]) ? node519 : node512;
								assign node512 = (inp[11]) ? node514 : 11'b00001001010;
									assign node514 = (inp[2]) ? node516 : 11'b00100011001;
										assign node516 = (inp[0]) ? 11'b00010111011 : 11'b00100101011;
								assign node519 = (inp[0]) ? node521 : 11'b10001111011;
									assign node521 = (inp[11]) ? 11'b00111001111 : node522;
										assign node522 = (inp[4]) ? node526 : node523;
											assign node523 = (inp[5]) ? 11'b00110001111 : 11'b00001101111;
											assign node526 = (inp[2]) ? 11'b00011111101 : node527;
												assign node527 = (inp[5]) ? 11'b00011111111 : 11'b00001111111;
							assign node532 = (inp[11]) ? node534 : 11'b10110011100;
								assign node534 = (inp[5]) ? 11'b00111001001 : node535;
									assign node535 = (inp[2]) ? 11'b00111001011 : 11'b00110001011;
						assign node539 = (inp[0]) ? node549 : node540;
							assign node540 = (inp[11]) ? node546 : node541;
								assign node541 = (inp[2]) ? 11'b00110011110 : node542;
									assign node542 = (inp[5]) ? 11'b10000111111 : 11'b00000111101;
								assign node546 = (inp[2]) ? 11'b00010101001 : 11'b00000001101;
							assign node549 = (inp[5]) ? node559 : node550;
								assign node550 = (inp[2]) ? 11'b00100111011 : node551;
									assign node551 = (inp[9]) ? node555 : node552;
										assign node552 = (inp[4]) ? 11'b00101101001 : 11'b00001101001;
										assign node555 = (inp[10]) ? 11'b00000101001 : 11'b00100101001;
								assign node559 = (inp[4]) ? node561 : 11'b00110001001;
									assign node561 = (inp[10]) ? 11'b00111101001 : node562;
										assign node562 = (inp[2]) ? 11'b00011111001 : 11'b00111111001;
					assign node566 = (inp[5]) ? node598 : node567;
						assign node567 = (inp[2]) ? node587 : node568;
							assign node568 = (inp[9]) ? node578 : node569;
								assign node569 = (inp[10]) ? node571 : 11'b00000001011;
									assign node571 = (inp[4]) ? node575 : node572;
										assign node572 = (inp[3]) ? 11'b00011011110 : 11'b00110111100;
										assign node575 = (inp[11]) ? 11'b00000001110 : 11'b00101111110;
								assign node578 = (inp[11]) ? node584 : node579;
									assign node579 = (inp[4]) ? node581 : 11'b10111101100;
										assign node581 = (inp[3]) ? 11'b10011111010 : 11'b00011111110;
									assign node584 = (inp[3]) ? 11'b00101011100 : 11'b10001011110;
							assign node587 = (inp[10]) ? node593 : node588;
								assign node588 = (inp[4]) ? node590 : 11'b10001001111;
									assign node590 = (inp[0]) ? 11'b00001011111 : 11'b10101011011;
								assign node593 = (inp[4]) ? 11'b00000101000 : node594;
									assign node594 = (inp[9]) ? 11'b00111011001 : 11'b00110011101;
						assign node598 = (inp[0]) ? node624 : node599;
							assign node599 = (inp[9]) ? node611 : node600;
								assign node600 = (inp[3]) ? 11'b10011101000 : node601;
									assign node601 = (inp[4]) ? node605 : node602;
										assign node602 = (inp[10]) ? 11'b10100011000 : 11'b00100111000;
										assign node605 = (inp[2]) ? 11'b00010111110 : node606;
											assign node606 = (inp[11]) ? 11'b00101011100 : 11'b00111111100;
								assign node611 = (inp[2]) ? node615 : node612;
									assign node612 = (inp[11]) ? 11'b00110001000 : 11'b00101101000;
									assign node615 = (inp[10]) ? node621 : node616;
										assign node616 = (inp[3]) ? 11'b10001001000 : node617;
											assign node617 = (inp[4]) ? 11'b00000001100 : 11'b00100001000;
										assign node621 = (inp[3]) ? 11'b00000101100 : 11'b10001001110;
							assign node624 = (inp[11]) ? node628 : node625;
								assign node625 = (inp[4]) ? 11'b00111011110 : 11'b00010001110;
								assign node628 = (inp[2]) ? node632 : node629;
									assign node629 = (inp[9]) ? 11'b00001001010 : 11'b00001011000;
									assign node632 = (inp[9]) ? node634 : 11'b00010001110;
										assign node634 = (inp[10]) ? 11'b00010001000 : 11'b00010001100;
				assign node637 = (inp[2]) ? node685 : node638;
					assign node638 = (inp[8]) ? node664 : node639;
						assign node639 = (inp[5]) ? node653 : node640;
							assign node640 = (inp[9]) ? node648 : node641;
								assign node641 = (inp[0]) ? node643 : 11'b10010101100;
									assign node643 = (inp[3]) ? 11'b00001101010 : node644;
										assign node644 = (inp[10]) ? 11'b00011111110 : 11'b00010101010;
								assign node648 = (inp[3]) ? 11'b00111111000 : node649;
									assign node649 = (inp[4]) ? 11'b10101101010 : 11'b00001101000;
							assign node653 = (inp[3]) ? 11'b00110100001 : node654;
								assign node654 = (inp[9]) ? node660 : node655;
									assign node655 = (inp[10]) ? node657 : 11'b00010011100;
										assign node657 = (inp[4]) ? 11'b00111100111 : 11'b00000110111;
									assign node660 = (inp[0]) ? 11'b00101100101 : 11'b00101110111;
						assign node664 = (inp[0]) ? node672 : node665;
							assign node665 = (inp[11]) ? node667 : 11'b00101100111;
								assign node667 = (inp[10]) ? node669 : 11'b10101010001;
									assign node669 = (inp[5]) ? 11'b00110000001 : 11'b00100010101;
							assign node672 = (inp[11]) ? node680 : node673;
								assign node673 = (inp[10]) ? node677 : node674;
									assign node674 = (inp[9]) ? 11'b00011010011 : 11'b00000010011;
									assign node677 = (inp[9]) ? 11'b00101010011 : 11'b00111000111;
								assign node680 = (inp[9]) ? node682 : 11'b00011100111;
									assign node682 = (inp[3]) ? 11'b00001000011 : 11'b00001100011;
					assign node685 = (inp[5]) ? node715 : node686;
						assign node686 = (inp[0]) ? node698 : node687;
							assign node687 = (inp[8]) ? node693 : node688;
								assign node688 = (inp[9]) ? 11'b10001110010 : node689;
									assign node689 = (inp[3]) ? 11'b10010100100 : 11'b10101100000;
								assign node693 = (inp[11]) ? 11'b00110110100 : node694;
									assign node694 = (inp[10]) ? 11'b00000000100 : 11'b00000100110;
							assign node698 = (inp[10]) ? node708 : node699;
								assign node699 = (inp[9]) ? node705 : node700;
									assign node700 = (inp[3]) ? 11'b00011110000 : node701;
										assign node701 = (inp[4]) ? 11'b00101110000 : 11'b00001110010;
									assign node705 = (inp[8]) ? 11'b00011110100 : 11'b00110110000;
								assign node708 = (inp[9]) ? node712 : node709;
									assign node709 = (inp[4]) ? 11'b00000010111 : 11'b00001000011;
									assign node712 = (inp[8]) ? 11'b00101110000 : 11'b00001100000;
						assign node715 = (inp[10]) ? node729 : node716;
							assign node716 = (inp[4]) ? node722 : node717;
								assign node717 = (inp[8]) ? 11'b00100110000 : node718;
									assign node718 = (inp[9]) ? 11'b10111010110 : 11'b00110000010;
								assign node722 = (inp[0]) ? node724 : 11'b00010000110;
									assign node724 = (inp[8]) ? node726 : 11'b00011010010;
										assign node726 = (inp[11]) ? 11'b00000010010 : 11'b00010000010;
							assign node729 = (inp[0]) ? node737 : node730;
								assign node730 = (inp[11]) ? 11'b10101000110 : node731;
									assign node731 = (inp[4]) ? node733 : 11'b00001010100;
										assign node733 = (inp[3]) ? 11'b00110010000 : 11'b10010010000;
								assign node737 = (inp[11]) ? node739 : 11'b00011000100;
									assign node739 = (inp[8]) ? node741 : 11'b00011000000;
										assign node741 = (inp[4]) ? node743 : 11'b00001000000;
											assign node743 = (inp[3]) ? 11'b00000000000 : 11'b00000000100;
			assign node746 = (inp[6]) ? node874 : node747;
				assign node747 = (inp[2]) ? node815 : node748;
					assign node748 = (inp[5]) ? node768 : node749;
						assign node749 = (inp[8]) ? node759 : node750;
							assign node750 = (inp[4]) ? node756 : node751;
								assign node751 = (inp[9]) ? 11'b00011100001 : node752;
									assign node752 = (inp[11]) ? 11'b00011100011 : 11'b00001100011;
								assign node756 = (inp[0]) ? 11'b00000110011 : 11'b10110110011;
							assign node759 = (inp[9]) ? 11'b10010100011 : node760;
								assign node760 = (inp[11]) ? node762 : 11'b10111110111;
									assign node762 = (inp[0]) ? node764 : 11'b00000110111;
										assign node764 = (inp[3]) ? 11'b00110100011 : 11'b00110110111;
						assign node768 = (inp[4]) ? node796 : node769;
							assign node769 = (inp[10]) ? node781 : node770;
								assign node770 = (inp[3]) ? 11'b10010110101 : node771;
									assign node771 = (inp[0]) ? 11'b00001010101 : node772;
										assign node772 = (inp[8]) ? 11'b00000110001 : node773;
											assign node773 = (inp[9]) ? 11'b00011010001 : node774;
												assign node774 = (inp[11]) ? 11'b00010010001 : 11'b00010110001;
								assign node781 = (inp[3]) ? node791 : node782;
									assign node782 = (inp[9]) ? 11'b00101010011 : node783;
										assign node783 = (inp[11]) ? node787 : node784;
											assign node784 = (inp[8]) ? 11'b00010100111 : 11'b00101000111;
											assign node787 = (inp[8]) ? 11'b00111010101 : 11'b00011010111;
									assign node791 = (inp[0]) ? node793 : 11'b00001000111;
										assign node793 = (inp[9]) ? 11'b00011000001 : 11'b00001000001;
							assign node796 = (inp[11]) ? node804 : node797;
								assign node797 = (inp[0]) ? node799 : 11'b10000000111;
									assign node799 = (inp[3]) ? 11'b00110010011 : node800;
										assign node800 = (inp[10]) ? 11'b00001010001 : 11'b00011010111;
								assign node804 = (inp[3]) ? node812 : node805;
									assign node805 = (inp[0]) ? node809 : node806;
										assign node806 = (inp[8]) ? 11'b00110000111 : 11'b00000000111;
										assign node809 = (inp[8]) ? 11'b00010000111 : 11'b00110000001;
									assign node812 = (inp[10]) ? 11'b00000000001 : 11'b10110000001;
					assign node815 = (inp[8]) ? node841 : node816;
						assign node816 = (inp[11]) ? node828 : node817;
							assign node817 = (inp[5]) ? node825 : node818;
								assign node818 = (inp[4]) ? node822 : node819;
									assign node819 = (inp[9]) ? 11'b00111000001 : 11'b00011000101;
									assign node822 = (inp[10]) ? 11'b00000000001 : 11'b00010000111;
								assign node825 = (inp[9]) ? 11'b10010100100 : 11'b00110100010;
							assign node828 = (inp[0]) ? node838 : node829;
								assign node829 = (inp[3]) ? node831 : 11'b10011110000;
									assign node831 = (inp[5]) ? node835 : node832;
										assign node832 = (inp[4]) ? 11'b10111110010 : 11'b10000000101;
										assign node835 = (inp[9]) ? 11'b10111110110 : 11'b00111100110;
								assign node838 = (inp[3]) ? 11'b00101110000 : 11'b00001100010;
						assign node841 = (inp[9]) ? node855 : node842;
							assign node842 = (inp[0]) ? node846 : node843;
								assign node843 = (inp[11]) ? 11'b00101010100 : 11'b10101000110;
								assign node846 = (inp[10]) ? node852 : node847;
									assign node847 = (inp[11]) ? 11'b00001000000 : node848;
										assign node848 = (inp[5]) ? 11'b00001000000 : 11'b00011010000;
									assign node852 = (inp[11]) ? 11'b00110000010 : 11'b00101010100;
							assign node855 = (inp[5]) ? node867 : node856;
								assign node856 = (inp[11]) ? node862 : node857;
									assign node857 = (inp[3]) ? 11'b00000110000 : node858;
										assign node858 = (inp[0]) ? 11'b00110100100 : 11'b00100100000;
									assign node862 = (inp[10]) ? node864 : 11'b10100010010;
										assign node864 = (inp[4]) ? 11'b00010000000 : 11'b00100000010;
								assign node867 = (inp[0]) ? node869 : 11'b00000000100;
									assign node869 = (inp[10]) ? 11'b00010000000 : node870;
										assign node870 = (inp[4]) ? 11'b00010000100 : 11'b00010010100;
				assign node874 = (inp[2]) ? node966 : node875;
					assign node875 = (inp[8]) ? node919 : node876;
						assign node876 = (inp[11]) ? node896 : node877;
							assign node877 = (inp[5]) ? node891 : node878;
								assign node878 = (inp[3]) ? node888 : node879;
									assign node879 = (inp[9]) ? node881 : 11'b00011100010;
										assign node881 = (inp[0]) ? node885 : node882;
											assign node882 = (inp[10]) ? 11'b10111100000 : 11'b00111100100;
											assign node885 = (inp[10]) ? 11'b00111110000 : 11'b00111110100;
									assign node888 = (inp[4]) ? 11'b00101100000 : 11'b00001110000;
								assign node891 = (inp[9]) ? node893 : 11'b00001110100;
									assign node893 = (inp[3]) ? 11'b10011110110 : 11'b10101100110;
							assign node896 = (inp[0]) ? node914 : node897;
								assign node897 = (inp[4]) ? node907 : node898;
									assign node898 = (inp[3]) ? node904 : node899;
										assign node899 = (inp[10]) ? 11'b10000100010 : node900;
											assign node900 = (inp[5]) ? 11'b00001110010 : 11'b00001100000;
										assign node904 = (inp[9]) ? 11'b00000100110 : 11'b00010110110;
									assign node907 = (inp[9]) ? node911 : node908;
										assign node908 = (inp[10]) ? 11'b10000100110 : 11'b10110100110;
										assign node911 = (inp[3]) ? 11'b00100110000 : 11'b00010110110;
								assign node914 = (inp[5]) ? node916 : 11'b00000110000;
									assign node916 = (inp[10]) ? 11'b00000100000 : 11'b00100100100;
						assign node919 = (inp[0]) ? node943 : node920;
							assign node920 = (inp[11]) ? node936 : node921;
								assign node921 = (inp[5]) ? node931 : node922;
									assign node922 = (inp[4]) ? node928 : node923;
										assign node923 = (inp[10]) ? 11'b00100110100 : node924;
											assign node924 = (inp[3]) ? 11'b10100100010 : 11'b00010100010;
										assign node928 = (inp[10]) ? 11'b10011000010 : 11'b10001010010;
									assign node931 = (inp[4]) ? 11'b10110000000 : node932;
										assign node932 = (inp[3]) ? 11'b10011010000 : 11'b10101010000;
								assign node936 = (inp[10]) ? node940 : node937;
									assign node937 = (inp[3]) ? 11'b10101000100 : 11'b00111010000;
									assign node940 = (inp[4]) ? 11'b10100000100 : 11'b10100000110;
							assign node943 = (inp[5]) ? node959 : node944;
								assign node944 = (inp[9]) ? node954 : node945;
									assign node945 = (inp[4]) ? node951 : node946;
										assign node946 = (inp[3]) ? 11'b00000100010 : node947;
											assign node947 = (inp[10]) ? 11'b00110100110 : 11'b00110100010;
										assign node951 = (inp[11]) ? 11'b00111010010 : 11'b00111000010;
									assign node954 = (inp[10]) ? 11'b00011000010 : node955;
										assign node955 = (inp[4]) ? 11'b00001010110 : 11'b00101010000;
								assign node959 = (inp[4]) ? node963 : node960;
									assign node960 = (inp[10]) ? 11'b00000000010 : 11'b00010010010;
									assign node963 = (inp[9]) ? 11'b00000010100 : 11'b00000000100;
					assign node966 = (inp[8]) ? node994 : node967;
						assign node967 = (inp[5]) ? node981 : node968;
							assign node968 = (inp[4]) ? node974 : node969;
								assign node969 = (inp[9]) ? node971 : 11'b00001000110;
									assign node971 = (inp[10]) ? 11'b00011000010 : 11'b00111000010;
								assign node974 = (inp[10]) ? node976 : 11'b10111000100;
									assign node976 = (inp[9]) ? node978 : 11'b00011010000;
										assign node978 = (inp[11]) ? 11'b10001010000 : 11'b00101010000;
							assign node981 = (inp[11]) ? node987 : node982;
								assign node982 = (inp[4]) ? 11'b00100010110 : node983;
									assign node983 = (inp[3]) ? 11'b00001010100 : 11'b00101010000;
								assign node987 = (inp[10]) ? node989 : 11'b00110010100;
									assign node989 = (inp[4]) ? 11'b10100000000 : node990;
										assign node990 = (inp[0]) ? 11'b00110000000 : 11'b10010010000;
						assign node994 = (inp[11]) ? node1006 : node995;
							assign node995 = (inp[10]) ? node1003 : node996;
								assign node996 = (inp[0]) ? node1000 : node997;
									assign node997 = (inp[4]) ? 11'b00000000110 : 11'b00110000010;
									assign node1000 = (inp[3]) ? 11'b00110010000 : 11'b00010000000;
								assign node1003 = (inp[5]) ? 11'b00010010100 : 11'b10010010110;
							assign node1006 = (inp[9]) ? node1014 : node1007;
								assign node1007 = (inp[0]) ? node1009 : 11'b10100010000;
									assign node1009 = (inp[10]) ? node1011 : 11'b00100010000;
										assign node1011 = (inp[3]) ? 11'b00100000000 : 11'b00000000100;
								assign node1014 = (inp[5]) ? node1016 : 11'b00100000100;
									assign node1016 = (inp[4]) ? node1018 : 11'b00000000100;
										assign node1018 = (inp[3]) ? 11'b00000000000 : 11'b00000000100;

endmodule