module dtc_split5_bm65 (
	input  wire [16-1:0] inp,
	output wire [4-1:0] outp
);

	wire [4-1:0] node1;
	wire [4-1:0] node2;
	wire [4-1:0] node3;
	wire [4-1:0] node4;
	wire [4-1:0] node5;
	wire [4-1:0] node6;
	wire [4-1:0] node7;
	wire [4-1:0] node8;
	wire [4-1:0] node9;
	wire [4-1:0] node10;
	wire [4-1:0] node11;
	wire [4-1:0] node12;
	wire [4-1:0] node13;
	wire [4-1:0] node14;
	wire [4-1:0] node19;
	wire [4-1:0] node20;
	wire [4-1:0] node24;
	wire [4-1:0] node25;
	wire [4-1:0] node26;
	wire [4-1:0] node30;
	wire [4-1:0] node32;
	wire [4-1:0] node36;
	wire [4-1:0] node37;
	wire [4-1:0] node38;
	wire [4-1:0] node39;
	wire [4-1:0] node41;
	wire [4-1:0] node42;
	wire [4-1:0] node44;
	wire [4-1:0] node48;
	wire [4-1:0] node49;
	wire [4-1:0] node50;
	wire [4-1:0] node55;
	wire [4-1:0] node56;
	wire [4-1:0] node57;
	wire [4-1:0] node58;
	wire [4-1:0] node62;
	wire [4-1:0] node64;
	wire [4-1:0] node67;
	wire [4-1:0] node68;
	wire [4-1:0] node72;
	wire [4-1:0] node73;
	wire [4-1:0] node74;
	wire [4-1:0] node75;
	wire [4-1:0] node78;
	wire [4-1:0] node81;
	wire [4-1:0] node82;
	wire [4-1:0] node83;
	wire [4-1:0] node88;
	wire [4-1:0] node89;
	wire [4-1:0] node90;
	wire [4-1:0] node94;
	wire [4-1:0] node96;
	wire [4-1:0] node99;
	wire [4-1:0] node100;
	wire [4-1:0] node101;
	wire [4-1:0] node102;
	wire [4-1:0] node103;
	wire [4-1:0] node104;
	wire [4-1:0] node107;
	wire [4-1:0] node110;
	wire [4-1:0] node111;
	wire [4-1:0] node112;
	wire [4-1:0] node116;
	wire [4-1:0] node117;
	wire [4-1:0] node121;
	wire [4-1:0] node122;
	wire [4-1:0] node124;
	wire [4-1:0] node125;
	wire [4-1:0] node129;
	wire [4-1:0] node130;
	wire [4-1:0] node134;
	wire [4-1:0] node135;
	wire [4-1:0] node136;
	wire [4-1:0] node137;
	wire [4-1:0] node139;
	wire [4-1:0] node142;
	wire [4-1:0] node145;
	wire [4-1:0] node146;
	wire [4-1:0] node148;
	wire [4-1:0] node151;
	wire [4-1:0] node152;
	wire [4-1:0] node156;
	wire [4-1:0] node157;
	wire [4-1:0] node160;
	wire [4-1:0] node161;
	wire [4-1:0] node162;
	wire [4-1:0] node166;
	wire [4-1:0] node169;
	wire [4-1:0] node170;
	wire [4-1:0] node171;
	wire [4-1:0] node172;
	wire [4-1:0] node173;
	wire [4-1:0] node174;
	wire [4-1:0] node179;
	wire [4-1:0] node181;
	wire [4-1:0] node182;
	wire [4-1:0] node186;
	wire [4-1:0] node187;
	wire [4-1:0] node188;
	wire [4-1:0] node190;
	wire [4-1:0] node193;
	wire [4-1:0] node194;
	wire [4-1:0] node198;
	wire [4-1:0] node199;
	wire [4-1:0] node203;
	wire [4-1:0] node204;
	wire [4-1:0] node205;
	wire [4-1:0] node206;
	wire [4-1:0] node209;
	wire [4-1:0] node212;
	wire [4-1:0] node213;
	wire [4-1:0] node216;
	wire [4-1:0] node219;
	wire [4-1:0] node220;
	wire [4-1:0] node223;
	wire [4-1:0] node225;
	wire [4-1:0] node229;
	wire [4-1:0] node230;
	wire [4-1:0] node231;
	wire [4-1:0] node232;
	wire [4-1:0] node233;
	wire [4-1:0] node234;
	wire [4-1:0] node235;
	wire [4-1:0] node237;
	wire [4-1:0] node241;
	wire [4-1:0] node243;
	wire [4-1:0] node246;
	wire [4-1:0] node247;
	wire [4-1:0] node248;
	wire [4-1:0] node249;
	wire [4-1:0] node251;
	wire [4-1:0] node254;
	wire [4-1:0] node256;
	wire [4-1:0] node259;
	wire [4-1:0] node260;
	wire [4-1:0] node264;
	wire [4-1:0] node265;
	wire [4-1:0] node266;
	wire [4-1:0] node268;
	wire [4-1:0] node272;
	wire [4-1:0] node275;
	wire [4-1:0] node276;
	wire [4-1:0] node277;
	wire [4-1:0] node279;
	wire [4-1:0] node282;
	wire [4-1:0] node283;
	wire [4-1:0] node286;
	wire [4-1:0] node287;
	wire [4-1:0] node291;
	wire [4-1:0] node292;
	wire [4-1:0] node294;
	wire [4-1:0] node295;
	wire [4-1:0] node299;
	wire [4-1:0] node300;
	wire [4-1:0] node304;
	wire [4-1:0] node305;
	wire [4-1:0] node306;
	wire [4-1:0] node307;
	wire [4-1:0] node308;
	wire [4-1:0] node309;
	wire [4-1:0] node311;
	wire [4-1:0] node314;
	wire [4-1:0] node317;
	wire [4-1:0] node318;
	wire [4-1:0] node321;
	wire [4-1:0] node323;
	wire [4-1:0] node326;
	wire [4-1:0] node327;
	wire [4-1:0] node328;
	wire [4-1:0] node332;
	wire [4-1:0] node333;
	wire [4-1:0] node337;
	wire [4-1:0] node338;
	wire [4-1:0] node339;
	wire [4-1:0] node340;
	wire [4-1:0] node343;
	wire [4-1:0] node346;
	wire [4-1:0] node347;
	wire [4-1:0] node351;
	wire [4-1:0] node352;
	wire [4-1:0] node353;
	wire [4-1:0] node355;
	wire [4-1:0] node359;
	wire [4-1:0] node361;
	wire [4-1:0] node364;
	wire [4-1:0] node365;
	wire [4-1:0] node366;
	wire [4-1:0] node367;
	wire [4-1:0] node368;
	wire [4-1:0] node371;
	wire [4-1:0] node372;
	wire [4-1:0] node373;
	wire [4-1:0] node377;
	wire [4-1:0] node380;
	wire [4-1:0] node383;
	wire [4-1:0] node384;
	wire [4-1:0] node385;
	wire [4-1:0] node389;
	wire [4-1:0] node392;
	wire [4-1:0] node393;
	wire [4-1:0] node394;
	wire [4-1:0] node395;
	wire [4-1:0] node399;
	wire [4-1:0] node401;
	wire [4-1:0] node402;
	wire [4-1:0] node406;
	wire [4-1:0] node407;
	wire [4-1:0] node408;
	wire [4-1:0] node412;
	wire [4-1:0] node415;
	wire [4-1:0] node416;
	wire [4-1:0] node417;
	wire [4-1:0] node418;
	wire [4-1:0] node419;
	wire [4-1:0] node420;
	wire [4-1:0] node422;
	wire [4-1:0] node424;
	wire [4-1:0] node427;
	wire [4-1:0] node428;
	wire [4-1:0] node430;
	wire [4-1:0] node434;
	wire [4-1:0] node435;
	wire [4-1:0] node438;
	wire [4-1:0] node441;
	wire [4-1:0] node442;
	wire [4-1:0] node443;
	wire [4-1:0] node444;
	wire [4-1:0] node446;
	wire [4-1:0] node449;
	wire [4-1:0] node450;
	wire [4-1:0] node454;
	wire [4-1:0] node456;
	wire [4-1:0] node459;
	wire [4-1:0] node460;
	wire [4-1:0] node463;
	wire [4-1:0] node465;
	wire [4-1:0] node468;
	wire [4-1:0] node469;
	wire [4-1:0] node470;
	wire [4-1:0] node472;
	wire [4-1:0] node473;
	wire [4-1:0] node477;
	wire [4-1:0] node479;
	wire [4-1:0] node480;
	wire [4-1:0] node484;
	wire [4-1:0] node485;
	wire [4-1:0] node486;
	wire [4-1:0] node490;
	wire [4-1:0] node491;
	wire [4-1:0] node493;
	wire [4-1:0] node496;
	wire [4-1:0] node499;
	wire [4-1:0] node500;
	wire [4-1:0] node501;
	wire [4-1:0] node502;
	wire [4-1:0] node503;
	wire [4-1:0] node505;
	wire [4-1:0] node509;
	wire [4-1:0] node510;
	wire [4-1:0] node514;
	wire [4-1:0] node515;
	wire [4-1:0] node516;
	wire [4-1:0] node517;
	wire [4-1:0] node521;
	wire [4-1:0] node523;
	wire [4-1:0] node526;
	wire [4-1:0] node527;
	wire [4-1:0] node529;
	wire [4-1:0] node532;
	wire [4-1:0] node534;
	wire [4-1:0] node537;
	wire [4-1:0] node538;
	wire [4-1:0] node539;
	wire [4-1:0] node540;
	wire [4-1:0] node541;
	wire [4-1:0] node545;
	wire [4-1:0] node546;
	wire [4-1:0] node547;
	wire [4-1:0] node552;
	wire [4-1:0] node554;
	wire [4-1:0] node555;
	wire [4-1:0] node558;
	wire [4-1:0] node559;
	wire [4-1:0] node563;
	wire [4-1:0] node564;
	wire [4-1:0] node565;
	wire [4-1:0] node567;
	wire [4-1:0] node570;
	wire [4-1:0] node571;
	wire [4-1:0] node575;
	wire [4-1:0] node576;
	wire [4-1:0] node577;
	wire [4-1:0] node580;
	wire [4-1:0] node581;
	wire [4-1:0] node585;
	wire [4-1:0] node586;
	wire [4-1:0] node588;
	wire [4-1:0] node589;
	wire [4-1:0] node595;
	wire [4-1:0] node596;
	wire [4-1:0] node597;
	wire [4-1:0] node599;
	wire [4-1:0] node600;
	wire [4-1:0] node601;
	wire [4-1:0] node602;
	wire [4-1:0] node603;
	wire [4-1:0] node604;
	wire [4-1:0] node606;
	wire [4-1:0] node608;
	wire [4-1:0] node611;
	wire [4-1:0] node613;
	wire [4-1:0] node614;
	wire [4-1:0] node617;
	wire [4-1:0] node620;
	wire [4-1:0] node621;
	wire [4-1:0] node622;
	wire [4-1:0] node625;
	wire [4-1:0] node628;
	wire [4-1:0] node630;
	wire [4-1:0] node632;
	wire [4-1:0] node636;
	wire [4-1:0] node637;
	wire [4-1:0] node638;
	wire [4-1:0] node639;
	wire [4-1:0] node640;
	wire [4-1:0] node644;
	wire [4-1:0] node645;
	wire [4-1:0] node649;
	wire [4-1:0] node650;
	wire [4-1:0] node651;
	wire [4-1:0] node653;
	wire [4-1:0] node655;
	wire [4-1:0] node658;
	wire [4-1:0] node659;
	wire [4-1:0] node663;
	wire [4-1:0] node664;
	wire [4-1:0] node666;
	wire [4-1:0] node669;
	wire [4-1:0] node670;
	wire [4-1:0] node674;
	wire [4-1:0] node675;
	wire [4-1:0] node677;
	wire [4-1:0] node678;
	wire [4-1:0] node681;
	wire [4-1:0] node683;
	wire [4-1:0] node684;
	wire [4-1:0] node688;
	wire [4-1:0] node689;
	wire [4-1:0] node690;
	wire [4-1:0] node693;
	wire [4-1:0] node694;
	wire [4-1:0] node698;
	wire [4-1:0] node700;
	wire [4-1:0] node704;
	wire [4-1:0] node705;
	wire [4-1:0] node706;
	wire [4-1:0] node707;
	wire [4-1:0] node708;
	wire [4-1:0] node709;
	wire [4-1:0] node710;
	wire [4-1:0] node712;
	wire [4-1:0] node716;
	wire [4-1:0] node717;
	wire [4-1:0] node721;
	wire [4-1:0] node722;
	wire [4-1:0] node723;
	wire [4-1:0] node725;
	wire [4-1:0] node728;
	wire [4-1:0] node729;
	wire [4-1:0] node730;
	wire [4-1:0] node735;
	wire [4-1:0] node736;
	wire [4-1:0] node738;
	wire [4-1:0] node741;
	wire [4-1:0] node742;
	wire [4-1:0] node746;
	wire [4-1:0] node747;
	wire [4-1:0] node748;
	wire [4-1:0] node749;
	wire [4-1:0] node751;
	wire [4-1:0] node753;
	wire [4-1:0] node754;
	wire [4-1:0] node757;
	wire [4-1:0] node760;
	wire [4-1:0] node762;
	wire [4-1:0] node764;
	wire [4-1:0] node767;
	wire [4-1:0] node768;
	wire [4-1:0] node769;
	wire [4-1:0] node771;
	wire [4-1:0] node774;
	wire [4-1:0] node776;
	wire [4-1:0] node779;
	wire [4-1:0] node780;
	wire [4-1:0] node783;
	wire [4-1:0] node785;
	wire [4-1:0] node788;
	wire [4-1:0] node789;
	wire [4-1:0] node790;
	wire [4-1:0] node791;
	wire [4-1:0] node793;
	wire [4-1:0] node796;
	wire [4-1:0] node799;
	wire [4-1:0] node800;
	wire [4-1:0] node803;
	wire [4-1:0] node806;
	wire [4-1:0] node807;
	wire [4-1:0] node808;
	wire [4-1:0] node811;
	wire [4-1:0] node812;
	wire [4-1:0] node816;
	wire [4-1:0] node818;
	wire [4-1:0] node819;
	wire [4-1:0] node821;
	wire [4-1:0] node824;
	wire [4-1:0] node825;
	wire [4-1:0] node829;
	wire [4-1:0] node830;
	wire [4-1:0] node831;
	wire [4-1:0] node832;
	wire [4-1:0] node834;
	wire [4-1:0] node835;
	wire [4-1:0] node837;
	wire [4-1:0] node840;
	wire [4-1:0] node843;
	wire [4-1:0] node844;
	wire [4-1:0] node848;
	wire [4-1:0] node849;
	wire [4-1:0] node850;
	wire [4-1:0] node851;
	wire [4-1:0] node853;
	wire [4-1:0] node857;
	wire [4-1:0] node859;
	wire [4-1:0] node862;
	wire [4-1:0] node863;
	wire [4-1:0] node864;
	wire [4-1:0] node865;
	wire [4-1:0] node869;
	wire [4-1:0] node870;
	wire [4-1:0] node874;
	wire [4-1:0] node875;
	wire [4-1:0] node876;
	wire [4-1:0] node880;
	wire [4-1:0] node883;
	wire [4-1:0] node884;
	wire [4-1:0] node885;
	wire [4-1:0] node886;
	wire [4-1:0] node887;
	wire [4-1:0] node889;
	wire [4-1:0] node892;
	wire [4-1:0] node893;
	wire [4-1:0] node895;
	wire [4-1:0] node899;
	wire [4-1:0] node901;
	wire [4-1:0] node903;
	wire [4-1:0] node906;
	wire [4-1:0] node907;
	wire [4-1:0] node908;
	wire [4-1:0] node911;
	wire [4-1:0] node913;
	wire [4-1:0] node916;
	wire [4-1:0] node917;
	wire [4-1:0] node918;
	wire [4-1:0] node922;
	wire [4-1:0] node925;
	wire [4-1:0] node926;
	wire [4-1:0] node927;
	wire [4-1:0] node928;
	wire [4-1:0] node930;
	wire [4-1:0] node933;
	wire [4-1:0] node934;
	wire [4-1:0] node938;
	wire [4-1:0] node939;
	wire [4-1:0] node942;
	wire [4-1:0] node944;
	wire [4-1:0] node947;
	wire [4-1:0] node948;
	wire [4-1:0] node949;
	wire [4-1:0] node952;
	wire [4-1:0] node954;
	wire [4-1:0] node957;
	wire [4-1:0] node958;
	wire [4-1:0] node959;
	wire [4-1:0] node963;
	wire [4-1:0] node965;
	wire [4-1:0] node968;
	wire [4-1:0] node970;
	wire [4-1:0] node971;
	wire [4-1:0] node972;
	wire [4-1:0] node973;
	wire [4-1:0] node974;
	wire [4-1:0] node975;
	wire [4-1:0] node979;
	wire [4-1:0] node980;
	wire [4-1:0] node982;
	wire [4-1:0] node985;
	wire [4-1:0] node987;
	wire [4-1:0] node990;
	wire [4-1:0] node991;
	wire [4-1:0] node992;
	wire [4-1:0] node995;
	wire [4-1:0] node996;
	wire [4-1:0] node999;
	wire [4-1:0] node1002;
	wire [4-1:0] node1003;
	wire [4-1:0] node1004;
	wire [4-1:0] node1008;
	wire [4-1:0] node1009;
	wire [4-1:0] node1014;
	wire [4-1:0] node1015;
	wire [4-1:0] node1016;
	wire [4-1:0] node1017;
	wire [4-1:0] node1018;
	wire [4-1:0] node1022;
	wire [4-1:0] node1023;
	wire [4-1:0] node1024;
	wire [4-1:0] node1029;
	wire [4-1:0] node1030;
	wire [4-1:0] node1031;
	wire [4-1:0] node1035;
	wire [4-1:0] node1037;
	wire [4-1:0] node1040;
	wire [4-1:0] node1041;
	wire [4-1:0] node1042;
	wire [4-1:0] node1043;
	wire [4-1:0] node1045;
	wire [4-1:0] node1049;
	wire [4-1:0] node1051;
	wire [4-1:0] node1054;
	wire [4-1:0] node1055;
	wire [4-1:0] node1056;
	wire [4-1:0] node1057;
	wire [4-1:0] node1061;
	wire [4-1:0] node1064;
	wire [4-1:0] node1065;
	wire [4-1:0] node1066;
	wire [4-1:0] node1068;
	wire [4-1:0] node1071;
	wire [4-1:0] node1076;
	wire [4-1:0] node1077;
	wire [4-1:0] node1078;
	wire [4-1:0] node1079;
	wire [4-1:0] node1080;
	wire [4-1:0] node1081;
	wire [4-1:0] node1082;
	wire [4-1:0] node1083;
	wire [4-1:0] node1084;
	wire [4-1:0] node1086;
	wire [4-1:0] node1089;
	wire [4-1:0] node1090;
	wire [4-1:0] node1091;
	wire [4-1:0] node1095;
	wire [4-1:0] node1096;
	wire [4-1:0] node1097;
	wire [4-1:0] node1100;
	wire [4-1:0] node1103;
	wire [4-1:0] node1106;
	wire [4-1:0] node1107;
	wire [4-1:0] node1108;
	wire [4-1:0] node1109;
	wire [4-1:0] node1111;
	wire [4-1:0] node1114;
	wire [4-1:0] node1115;
	wire [4-1:0] node1119;
	wire [4-1:0] node1120;
	wire [4-1:0] node1124;
	wire [4-1:0] node1125;
	wire [4-1:0] node1127;
	wire [4-1:0] node1130;
	wire [4-1:0] node1131;
	wire [4-1:0] node1132;
	wire [4-1:0] node1133;
	wire [4-1:0] node1139;
	wire [4-1:0] node1140;
	wire [4-1:0] node1141;
	wire [4-1:0] node1142;
	wire [4-1:0] node1144;
	wire [4-1:0] node1147;
	wire [4-1:0] node1148;
	wire [4-1:0] node1151;
	wire [4-1:0] node1152;
	wire [4-1:0] node1155;
	wire [4-1:0] node1158;
	wire [4-1:0] node1159;
	wire [4-1:0] node1160;
	wire [4-1:0] node1162;
	wire [4-1:0] node1163;
	wire [4-1:0] node1166;
	wire [4-1:0] node1170;
	wire [4-1:0] node1171;
	wire [4-1:0] node1173;
	wire [4-1:0] node1176;
	wire [4-1:0] node1178;
	wire [4-1:0] node1179;
	wire [4-1:0] node1182;
	wire [4-1:0] node1185;
	wire [4-1:0] node1186;
	wire [4-1:0] node1188;
	wire [4-1:0] node1190;
	wire [4-1:0] node1193;
	wire [4-1:0] node1194;
	wire [4-1:0] node1195;
	wire [4-1:0] node1196;
	wire [4-1:0] node1199;
	wire [4-1:0] node1200;
	wire [4-1:0] node1204;
	wire [4-1:0] node1205;
	wire [4-1:0] node1208;
	wire [4-1:0] node1209;
	wire [4-1:0] node1212;
	wire [4-1:0] node1215;
	wire [4-1:0] node1216;
	wire [4-1:0] node1220;
	wire [4-1:0] node1221;
	wire [4-1:0] node1222;
	wire [4-1:0] node1223;
	wire [4-1:0] node1224;
	wire [4-1:0] node1225;
	wire [4-1:0] node1229;
	wire [4-1:0] node1230;
	wire [4-1:0] node1234;
	wire [4-1:0] node1235;
	wire [4-1:0] node1236;
	wire [4-1:0] node1239;
	wire [4-1:0] node1241;
	wire [4-1:0] node1242;
	wire [4-1:0] node1245;
	wire [4-1:0] node1248;
	wire [4-1:0] node1250;
	wire [4-1:0] node1251;
	wire [4-1:0] node1255;
	wire [4-1:0] node1256;
	wire [4-1:0] node1257;
	wire [4-1:0] node1258;
	wire [4-1:0] node1259;
	wire [4-1:0] node1261;
	wire [4-1:0] node1266;
	wire [4-1:0] node1267;
	wire [4-1:0] node1268;
	wire [4-1:0] node1273;
	wire [4-1:0] node1274;
	wire [4-1:0] node1275;
	wire [4-1:0] node1276;
	wire [4-1:0] node1279;
	wire [4-1:0] node1282;
	wire [4-1:0] node1283;
	wire [4-1:0] node1286;
	wire [4-1:0] node1288;
	wire [4-1:0] node1291;
	wire [4-1:0] node1292;
	wire [4-1:0] node1295;
	wire [4-1:0] node1297;
	wire [4-1:0] node1300;
	wire [4-1:0] node1301;
	wire [4-1:0] node1302;
	wire [4-1:0] node1303;
	wire [4-1:0] node1304;
	wire [4-1:0] node1307;
	wire [4-1:0] node1308;
	wire [4-1:0] node1311;
	wire [4-1:0] node1312;
	wire [4-1:0] node1315;
	wire [4-1:0] node1318;
	wire [4-1:0] node1319;
	wire [4-1:0] node1320;
	wire [4-1:0] node1324;
	wire [4-1:0] node1326;
	wire [4-1:0] node1329;
	wire [4-1:0] node1330;
	wire [4-1:0] node1331;
	wire [4-1:0] node1332;
	wire [4-1:0] node1333;
	wire [4-1:0] node1337;
	wire [4-1:0] node1338;
	wire [4-1:0] node1341;
	wire [4-1:0] node1344;
	wire [4-1:0] node1347;
	wire [4-1:0] node1348;
	wire [4-1:0] node1349;
	wire [4-1:0] node1352;
	wire [4-1:0] node1355;
	wire [4-1:0] node1357;
	wire [4-1:0] node1360;
	wire [4-1:0] node1361;
	wire [4-1:0] node1362;
	wire [4-1:0] node1363;
	wire [4-1:0] node1366;
	wire [4-1:0] node1367;
	wire [4-1:0] node1370;
	wire [4-1:0] node1373;
	wire [4-1:0] node1374;
	wire [4-1:0] node1376;
	wire [4-1:0] node1379;
	wire [4-1:0] node1382;
	wire [4-1:0] node1383;
	wire [4-1:0] node1384;
	wire [4-1:0] node1388;
	wire [4-1:0] node1389;
	wire [4-1:0] node1392;
	wire [4-1:0] node1394;
	wire [4-1:0] node1397;
	wire [4-1:0] node1398;
	wire [4-1:0] node1399;
	wire [4-1:0] node1400;
	wire [4-1:0] node1401;
	wire [4-1:0] node1402;
	wire [4-1:0] node1403;
	wire [4-1:0] node1404;
	wire [4-1:0] node1407;
	wire [4-1:0] node1411;
	wire [4-1:0] node1412;
	wire [4-1:0] node1413;
	wire [4-1:0] node1418;
	wire [4-1:0] node1419;
	wire [4-1:0] node1421;
	wire [4-1:0] node1422;
	wire [4-1:0] node1426;
	wire [4-1:0] node1427;
	wire [4-1:0] node1430;
	wire [4-1:0] node1431;
	wire [4-1:0] node1435;
	wire [4-1:0] node1436;
	wire [4-1:0] node1437;
	wire [4-1:0] node1438;
	wire [4-1:0] node1441;
	wire [4-1:0] node1444;
	wire [4-1:0] node1445;
	wire [4-1:0] node1447;
	wire [4-1:0] node1450;
	wire [4-1:0] node1452;
	wire [4-1:0] node1455;
	wire [4-1:0] node1456;
	wire [4-1:0] node1457;
	wire [4-1:0] node1459;
	wire [4-1:0] node1462;
	wire [4-1:0] node1463;
	wire [4-1:0] node1467;
	wire [4-1:0] node1468;
	wire [4-1:0] node1469;
	wire [4-1:0] node1472;
	wire [4-1:0] node1475;
	wire [4-1:0] node1478;
	wire [4-1:0] node1479;
	wire [4-1:0] node1480;
	wire [4-1:0] node1481;
	wire [4-1:0] node1482;
	wire [4-1:0] node1484;
	wire [4-1:0] node1487;
	wire [4-1:0] node1490;
	wire [4-1:0] node1491;
	wire [4-1:0] node1494;
	wire [4-1:0] node1497;
	wire [4-1:0] node1498;
	wire [4-1:0] node1500;
	wire [4-1:0] node1503;
	wire [4-1:0] node1504;
	wire [4-1:0] node1505;
	wire [4-1:0] node1508;
	wire [4-1:0] node1512;
	wire [4-1:0] node1513;
	wire [4-1:0] node1514;
	wire [4-1:0] node1515;
	wire [4-1:0] node1516;
	wire [4-1:0] node1520;
	wire [4-1:0] node1521;
	wire [4-1:0] node1525;
	wire [4-1:0] node1526;
	wire [4-1:0] node1527;
	wire [4-1:0] node1530;
	wire [4-1:0] node1533;
	wire [4-1:0] node1535;
	wire [4-1:0] node1536;
	wire [4-1:0] node1540;
	wire [4-1:0] node1541;
	wire [4-1:0] node1542;
	wire [4-1:0] node1545;
	wire [4-1:0] node1548;
	wire [4-1:0] node1549;
	wire [4-1:0] node1550;
	wire [4-1:0] node1555;
	wire [4-1:0] node1556;
	wire [4-1:0] node1557;
	wire [4-1:0] node1558;
	wire [4-1:0] node1559;
	wire [4-1:0] node1560;
	wire [4-1:0] node1562;
	wire [4-1:0] node1563;
	wire [4-1:0] node1567;
	wire [4-1:0] node1570;
	wire [4-1:0] node1571;
	wire [4-1:0] node1574;
	wire [4-1:0] node1576;
	wire [4-1:0] node1579;
	wire [4-1:0] node1580;
	wire [4-1:0] node1582;
	wire [4-1:0] node1583;
	wire [4-1:0] node1586;
	wire [4-1:0] node1589;
	wire [4-1:0] node1590;
	wire [4-1:0] node1592;
	wire [4-1:0] node1594;
	wire [4-1:0] node1597;
	wire [4-1:0] node1599;
	wire [4-1:0] node1601;
	wire [4-1:0] node1604;
	wire [4-1:0] node1605;
	wire [4-1:0] node1606;
	wire [4-1:0] node1607;
	wire [4-1:0] node1608;
	wire [4-1:0] node1613;
	wire [4-1:0] node1614;
	wire [4-1:0] node1616;
	wire [4-1:0] node1620;
	wire [4-1:0] node1621;
	wire [4-1:0] node1623;
	wire [4-1:0] node1624;
	wire [4-1:0] node1628;
	wire [4-1:0] node1629;
	wire [4-1:0] node1632;
	wire [4-1:0] node1633;
	wire [4-1:0] node1637;
	wire [4-1:0] node1638;
	wire [4-1:0] node1639;
	wire [4-1:0] node1640;
	wire [4-1:0] node1641;
	wire [4-1:0] node1644;
	wire [4-1:0] node1645;
	wire [4-1:0] node1649;
	wire [4-1:0] node1650;
	wire [4-1:0] node1653;
	wire [4-1:0] node1654;
	wire [4-1:0] node1658;
	wire [4-1:0] node1659;
	wire [4-1:0] node1662;
	wire [4-1:0] node1663;
	wire [4-1:0] node1667;
	wire [4-1:0] node1668;
	wire [4-1:0] node1669;
	wire [4-1:0] node1670;
	wire [4-1:0] node1671;
	wire [4-1:0] node1675;
	wire [4-1:0] node1676;
	wire [4-1:0] node1680;
	wire [4-1:0] node1681;
	wire [4-1:0] node1683;
	wire [4-1:0] node1686;
	wire [4-1:0] node1688;
	wire [4-1:0] node1691;
	wire [4-1:0] node1692;
	wire [4-1:0] node1693;
	wire [4-1:0] node1694;
	wire [4-1:0] node1695;
	wire [4-1:0] node1699;
	wire [4-1:0] node1702;
	wire [4-1:0] node1705;
	wire [4-1:0] node1706;
	wire [4-1:0] node1708;
	wire [4-1:0] node1711;
	wire [4-1:0] node1714;
	wire [4-1:0] node1715;
	wire [4-1:0] node1716;
	wire [4-1:0] node1717;
	wire [4-1:0] node1718;
	wire [4-1:0] node1719;
	wire [4-1:0] node1720;
	wire [4-1:0] node1721;
	wire [4-1:0] node1722;
	wire [4-1:0] node1725;
	wire [4-1:0] node1728;
	wire [4-1:0] node1730;
	wire [4-1:0] node1733;
	wire [4-1:0] node1734;
	wire [4-1:0] node1737;
	wire [4-1:0] node1739;
	wire [4-1:0] node1742;
	wire [4-1:0] node1743;
	wire [4-1:0] node1745;
	wire [4-1:0] node1746;
	wire [4-1:0] node1747;
	wire [4-1:0] node1750;
	wire [4-1:0] node1753;
	wire [4-1:0] node1755;
	wire [4-1:0] node1758;
	wire [4-1:0] node1760;
	wire [4-1:0] node1761;
	wire [4-1:0] node1765;
	wire [4-1:0] node1766;
	wire [4-1:0] node1767;
	wire [4-1:0] node1768;
	wire [4-1:0] node1772;
	wire [4-1:0] node1773;
	wire [4-1:0] node1775;
	wire [4-1:0] node1778;
	wire [4-1:0] node1781;
	wire [4-1:0] node1782;
	wire [4-1:0] node1784;
	wire [4-1:0] node1785;
	wire [4-1:0] node1789;
	wire [4-1:0] node1790;
	wire [4-1:0] node1794;
	wire [4-1:0] node1795;
	wire [4-1:0] node1796;
	wire [4-1:0] node1797;
	wire [4-1:0] node1798;
	wire [4-1:0] node1801;
	wire [4-1:0] node1803;
	wire [4-1:0] node1806;
	wire [4-1:0] node1807;
	wire [4-1:0] node1809;
	wire [4-1:0] node1811;
	wire [4-1:0] node1814;
	wire [4-1:0] node1817;
	wire [4-1:0] node1818;
	wire [4-1:0] node1819;
	wire [4-1:0] node1823;
	wire [4-1:0] node1824;
	wire [4-1:0] node1828;
	wire [4-1:0] node1829;
	wire [4-1:0] node1830;
	wire [4-1:0] node1832;
	wire [4-1:0] node1835;
	wire [4-1:0] node1837;
	wire [4-1:0] node1840;
	wire [4-1:0] node1841;
	wire [4-1:0] node1842;
	wire [4-1:0] node1843;
	wire [4-1:0] node1847;
	wire [4-1:0] node1848;
	wire [4-1:0] node1852;
	wire [4-1:0] node1853;
	wire [4-1:0] node1855;
	wire [4-1:0] node1858;
	wire [4-1:0] node1861;
	wire [4-1:0] node1862;
	wire [4-1:0] node1863;
	wire [4-1:0] node1864;
	wire [4-1:0] node1865;
	wire [4-1:0] node1867;
	wire [4-1:0] node1870;
	wire [4-1:0] node1871;
	wire [4-1:0] node1875;
	wire [4-1:0] node1876;
	wire [4-1:0] node1877;
	wire [4-1:0] node1878;
	wire [4-1:0] node1881;
	wire [4-1:0] node1884;
	wire [4-1:0] node1885;
	wire [4-1:0] node1889;
	wire [4-1:0] node1890;
	wire [4-1:0] node1892;
	wire [4-1:0] node1896;
	wire [4-1:0] node1897;
	wire [4-1:0] node1898;
	wire [4-1:0] node1899;
	wire [4-1:0] node1900;
	wire [4-1:0] node1904;
	wire [4-1:0] node1907;
	wire [4-1:0] node1908;
	wire [4-1:0] node1912;
	wire [4-1:0] node1913;
	wire [4-1:0] node1914;
	wire [4-1:0] node1917;
	wire [4-1:0] node1920;
	wire [4-1:0] node1922;
	wire [4-1:0] node1925;
	wire [4-1:0] node1926;
	wire [4-1:0] node1927;
	wire [4-1:0] node1929;
	wire [4-1:0] node1930;
	wire [4-1:0] node1933;
	wire [4-1:0] node1936;
	wire [4-1:0] node1937;
	wire [4-1:0] node1938;
	wire [4-1:0] node1939;
	wire [4-1:0] node1940;
	wire [4-1:0] node1945;
	wire [4-1:0] node1948;
	wire [4-1:0] node1950;
	wire [4-1:0] node1953;
	wire [4-1:0] node1954;
	wire [4-1:0] node1955;
	wire [4-1:0] node1956;
	wire [4-1:0] node1957;
	wire [4-1:0] node1959;
	wire [4-1:0] node1962;
	wire [4-1:0] node1965;
	wire [4-1:0] node1966;
	wire [4-1:0] node1970;
	wire [4-1:0] node1972;
	wire [4-1:0] node1975;
	wire [4-1:0] node1976;
	wire [4-1:0] node1977;
	wire [4-1:0] node1978;
	wire [4-1:0] node1982;
	wire [4-1:0] node1983;
	wire [4-1:0] node1987;
	wire [4-1:0] node1988;
	wire [4-1:0] node1990;
	wire [4-1:0] node1993;
	wire [4-1:0] node1994;
	wire [4-1:0] node1998;
	wire [4-1:0] node1999;
	wire [4-1:0] node2000;
	wire [4-1:0] node2001;
	wire [4-1:0] node2002;
	wire [4-1:0] node2003;
	wire [4-1:0] node2004;
	wire [4-1:0] node2008;
	wire [4-1:0] node2009;
	wire [4-1:0] node2010;
	wire [4-1:0] node2014;
	wire [4-1:0] node2015;
	wire [4-1:0] node2019;
	wire [4-1:0] node2020;
	wire [4-1:0] node2021;
	wire [4-1:0] node2025;
	wire [4-1:0] node2028;
	wire [4-1:0] node2029;
	wire [4-1:0] node2030;
	wire [4-1:0] node2031;
	wire [4-1:0] node2032;
	wire [4-1:0] node2036;
	wire [4-1:0] node2038;
	wire [4-1:0] node2041;
	wire [4-1:0] node2042;
	wire [4-1:0] node2044;
	wire [4-1:0] node2045;
	wire [4-1:0] node2049;
	wire [4-1:0] node2051;
	wire [4-1:0] node2054;
	wire [4-1:0] node2055;
	wire [4-1:0] node2056;
	wire [4-1:0] node2059;
	wire [4-1:0] node2060;
	wire [4-1:0] node2064;
	wire [4-1:0] node2065;
	wire [4-1:0] node2068;
	wire [4-1:0] node2069;
	wire [4-1:0] node2073;
	wire [4-1:0] node2074;
	wire [4-1:0] node2075;
	wire [4-1:0] node2077;
	wire [4-1:0] node2078;
	wire [4-1:0] node2079;
	wire [4-1:0] node2083;
	wire [4-1:0] node2084;
	wire [4-1:0] node2088;
	wire [4-1:0] node2089;
	wire [4-1:0] node2090;
	wire [4-1:0] node2093;
	wire [4-1:0] node2095;
	wire [4-1:0] node2098;
	wire [4-1:0] node2100;
	wire [4-1:0] node2103;
	wire [4-1:0] node2104;
	wire [4-1:0] node2105;
	wire [4-1:0] node2106;
	wire [4-1:0] node2110;
	wire [4-1:0] node2111;
	wire [4-1:0] node2112;
	wire [4-1:0] node2116;
	wire [4-1:0] node2119;
	wire [4-1:0] node2120;
	wire [4-1:0] node2122;
	wire [4-1:0] node2123;
	wire [4-1:0] node2126;
	wire [4-1:0] node2129;
	wire [4-1:0] node2130;
	wire [4-1:0] node2134;
	wire [4-1:0] node2135;
	wire [4-1:0] node2136;
	wire [4-1:0] node2137;
	wire [4-1:0] node2138;
	wire [4-1:0] node2141;
	wire [4-1:0] node2143;
	wire [4-1:0] node2146;
	wire [4-1:0] node2147;
	wire [4-1:0] node2148;
	wire [4-1:0] node2151;
	wire [4-1:0] node2154;
	wire [4-1:0] node2155;
	wire [4-1:0] node2158;
	wire [4-1:0] node2161;
	wire [4-1:0] node2162;
	wire [4-1:0] node2163;
	wire [4-1:0] node2164;
	wire [4-1:0] node2165;
	wire [4-1:0] node2170;
	wire [4-1:0] node2173;
	wire [4-1:0] node2174;
	wire [4-1:0] node2176;
	wire [4-1:0] node2177;
	wire [4-1:0] node2181;
	wire [4-1:0] node2182;
	wire [4-1:0] node2185;
	wire [4-1:0] node2188;
	wire [4-1:0] node2189;
	wire [4-1:0] node2190;
	wire [4-1:0] node2191;
	wire [4-1:0] node2192;
	wire [4-1:0] node2197;
	wire [4-1:0] node2198;
	wire [4-1:0] node2199;
	wire [4-1:0] node2203;
	wire [4-1:0] node2204;
	wire [4-1:0] node2207;
	wire [4-1:0] node2210;
	wire [4-1:0] node2211;
	wire [4-1:0] node2213;
	wire [4-1:0] node2216;
	wire [4-1:0] node2218;
	wire [4-1:0] node2221;
	wire [4-1:0] node2222;
	wire [4-1:0] node2223;
	wire [4-1:0] node2224;
	wire [4-1:0] node2225;
	wire [4-1:0] node2226;
	wire [4-1:0] node2227;
	wire [4-1:0] node2228;
	wire [4-1:0] node2229;
	wire [4-1:0] node2230;
	wire [4-1:0] node2233;
	wire [4-1:0] node2237;
	wire [4-1:0] node2238;
	wire [4-1:0] node2239;
	wire [4-1:0] node2240;
	wire [4-1:0] node2246;
	wire [4-1:0] node2247;
	wire [4-1:0] node2248;
	wire [4-1:0] node2249;
	wire [4-1:0] node2250;
	wire [4-1:0] node2255;
	wire [4-1:0] node2256;
	wire [4-1:0] node2260;
	wire [4-1:0] node2262;
	wire [4-1:0] node2265;
	wire [4-1:0] node2266;
	wire [4-1:0] node2267;
	wire [4-1:0] node2269;
	wire [4-1:0] node2270;
	wire [4-1:0] node2275;
	wire [4-1:0] node2276;
	wire [4-1:0] node2277;
	wire [4-1:0] node2279;
	wire [4-1:0] node2282;
	wire [4-1:0] node2283;
	wire [4-1:0] node2287;
	wire [4-1:0] node2288;
	wire [4-1:0] node2291;
	wire [4-1:0] node2292;
	wire [4-1:0] node2296;
	wire [4-1:0] node2297;
	wire [4-1:0] node2298;
	wire [4-1:0] node2299;
	wire [4-1:0] node2300;
	wire [4-1:0] node2302;
	wire [4-1:0] node2306;
	wire [4-1:0] node2308;
	wire [4-1:0] node2311;
	wire [4-1:0] node2313;
	wire [4-1:0] node2314;
	wire [4-1:0] node2315;
	wire [4-1:0] node2318;
	wire [4-1:0] node2322;
	wire [4-1:0] node2323;
	wire [4-1:0] node2324;
	wire [4-1:0] node2325;
	wire [4-1:0] node2328;
	wire [4-1:0] node2331;
	wire [4-1:0] node2333;
	wire [4-1:0] node2334;
	wire [4-1:0] node2337;
	wire [4-1:0] node2340;
	wire [4-1:0] node2341;
	wire [4-1:0] node2342;
	wire [4-1:0] node2344;
	wire [4-1:0] node2346;
	wire [4-1:0] node2350;
	wire [4-1:0] node2352;
	wire [4-1:0] node2355;
	wire [4-1:0] node2356;
	wire [4-1:0] node2357;
	wire [4-1:0] node2358;
	wire [4-1:0] node2359;
	wire [4-1:0] node2360;
	wire [4-1:0] node2363;
	wire [4-1:0] node2366;
	wire [4-1:0] node2368;
	wire [4-1:0] node2371;
	wire [4-1:0] node2372;
	wire [4-1:0] node2373;
	wire [4-1:0] node2377;
	wire [4-1:0] node2378;
	wire [4-1:0] node2381;
	wire [4-1:0] node2384;
	wire [4-1:0] node2386;
	wire [4-1:0] node2387;
	wire [4-1:0] node2388;
	wire [4-1:0] node2389;
	wire [4-1:0] node2394;
	wire [4-1:0] node2396;
	wire [4-1:0] node2397;
	wire [4-1:0] node2400;
	wire [4-1:0] node2403;
	wire [4-1:0] node2404;
	wire [4-1:0] node2405;
	wire [4-1:0] node2406;
	wire [4-1:0] node2408;
	wire [4-1:0] node2411;
	wire [4-1:0] node2412;
	wire [4-1:0] node2413;
	wire [4-1:0] node2417;
	wire [4-1:0] node2419;
	wire [4-1:0] node2422;
	wire [4-1:0] node2423;
	wire [4-1:0] node2424;
	wire [4-1:0] node2426;
	wire [4-1:0] node2427;
	wire [4-1:0] node2432;
	wire [4-1:0] node2433;
	wire [4-1:0] node2436;
	wire [4-1:0] node2439;
	wire [4-1:0] node2440;
	wire [4-1:0] node2441;
	wire [4-1:0] node2442;
	wire [4-1:0] node2446;
	wire [4-1:0] node2447;
	wire [4-1:0] node2450;
	wire [4-1:0] node2453;
	wire [4-1:0] node2454;
	wire [4-1:0] node2455;
	wire [4-1:0] node2457;
	wire [4-1:0] node2460;
	wire [4-1:0] node2463;
	wire [4-1:0] node2464;
	wire [4-1:0] node2465;
	wire [4-1:0] node2471;
	wire [4-1:0] node2472;
	wire [4-1:0] node2474;
	wire [4-1:0] node2475;
	wire [4-1:0] node2476;
	wire [4-1:0] node2477;
	wire [4-1:0] node2478;
	wire [4-1:0] node2479;
	wire [4-1:0] node2481;
	wire [4-1:0] node2482;
	wire [4-1:0] node2487;
	wire [4-1:0] node2488;
	wire [4-1:0] node2490;
	wire [4-1:0] node2491;
	wire [4-1:0] node2496;
	wire [4-1:0] node2497;
	wire [4-1:0] node2498;
	wire [4-1:0] node2502;
	wire [4-1:0] node2503;
	wire [4-1:0] node2506;
	wire [4-1:0] node2510;
	wire [4-1:0] node2511;
	wire [4-1:0] node2512;
	wire [4-1:0] node2513;
	wire [4-1:0] node2515;
	wire [4-1:0] node2518;
	wire [4-1:0] node2520;
	wire [4-1:0] node2523;
	wire [4-1:0] node2524;
	wire [4-1:0] node2525;
	wire [4-1:0] node2526;
	wire [4-1:0] node2530;
	wire [4-1:0] node2531;
	wire [4-1:0] node2535;
	wire [4-1:0] node2536;
	wire [4-1:0] node2540;
	wire [4-1:0] node2541;
	wire [4-1:0] node2542;
	wire [4-1:0] node2543;
	wire [4-1:0] node2545;
	wire [4-1:0] node2548;
	wire [4-1:0] node2552;
	wire [4-1:0] node2553;
	wire [4-1:0] node2554;
	wire [4-1:0] node2557;
	wire [4-1:0] node2558;
	wire [4-1:0] node2562;
	wire [4-1:0] node2563;
	wire [4-1:0] node2568;
	wire [4-1:0] node2569;
	wire [4-1:0] node2570;
	wire [4-1:0] node2571;
	wire [4-1:0] node2572;
	wire [4-1:0] node2573;
	wire [4-1:0] node2574;
	wire [4-1:0] node2575;
	wire [4-1:0] node2576;
	wire [4-1:0] node2577;
	wire [4-1:0] node2579;
	wire [4-1:0] node2582;
	wire [4-1:0] node2583;
	wire [4-1:0] node2584;
	wire [4-1:0] node2589;
	wire [4-1:0] node2590;
	wire [4-1:0] node2591;
	wire [4-1:0] node2592;
	wire [4-1:0] node2595;
	wire [4-1:0] node2600;
	wire [4-1:0] node2601;
	wire [4-1:0] node2602;
	wire [4-1:0] node2603;
	wire [4-1:0] node2605;
	wire [4-1:0] node2608;
	wire [4-1:0] node2611;
	wire [4-1:0] node2612;
	wire [4-1:0] node2615;
	wire [4-1:0] node2618;
	wire [4-1:0] node2619;
	wire [4-1:0] node2621;
	wire [4-1:0] node2624;
	wire [4-1:0] node2627;
	wire [4-1:0] node2628;
	wire [4-1:0] node2629;
	wire [4-1:0] node2630;
	wire [4-1:0] node2632;
	wire [4-1:0] node2636;
	wire [4-1:0] node2637;
	wire [4-1:0] node2639;
	wire [4-1:0] node2643;
	wire [4-1:0] node2644;
	wire [4-1:0] node2645;
	wire [4-1:0] node2646;
	wire [4-1:0] node2650;
	wire [4-1:0] node2652;
	wire [4-1:0] node2655;
	wire [4-1:0] node2656;
	wire [4-1:0] node2658;
	wire [4-1:0] node2661;
	wire [4-1:0] node2664;
	wire [4-1:0] node2665;
	wire [4-1:0] node2666;
	wire [4-1:0] node2667;
	wire [4-1:0] node2669;
	wire [4-1:0] node2671;
	wire [4-1:0] node2672;
	wire [4-1:0] node2676;
	wire [4-1:0] node2677;
	wire [4-1:0] node2678;
	wire [4-1:0] node2682;
	wire [4-1:0] node2685;
	wire [4-1:0] node2686;
	wire [4-1:0] node2688;
	wire [4-1:0] node2691;
	wire [4-1:0] node2693;
	wire [4-1:0] node2694;
	wire [4-1:0] node2698;
	wire [4-1:0] node2699;
	wire [4-1:0] node2700;
	wire [4-1:0] node2701;
	wire [4-1:0] node2705;
	wire [4-1:0] node2706;
	wire [4-1:0] node2707;
	wire [4-1:0] node2711;
	wire [4-1:0] node2714;
	wire [4-1:0] node2715;
	wire [4-1:0] node2716;
	wire [4-1:0] node2719;
	wire [4-1:0] node2722;
	wire [4-1:0] node2723;
	wire [4-1:0] node2724;
	wire [4-1:0] node2727;
	wire [4-1:0] node2730;
	wire [4-1:0] node2731;
	wire [4-1:0] node2733;
	wire [4-1:0] node2736;
	wire [4-1:0] node2739;
	wire [4-1:0] node2740;
	wire [4-1:0] node2741;
	wire [4-1:0] node2742;
	wire [4-1:0] node2743;
	wire [4-1:0] node2745;
	wire [4-1:0] node2748;
	wire [4-1:0] node2750;
	wire [4-1:0] node2753;
	wire [4-1:0] node2754;
	wire [4-1:0] node2755;
	wire [4-1:0] node2758;
	wire [4-1:0] node2761;
	wire [4-1:0] node2762;
	wire [4-1:0] node2766;
	wire [4-1:0] node2767;
	wire [4-1:0] node2768;
	wire [4-1:0] node2769;
	wire [4-1:0] node2771;
	wire [4-1:0] node2774;
	wire [4-1:0] node2777;
	wire [4-1:0] node2779;
	wire [4-1:0] node2781;
	wire [4-1:0] node2784;
	wire [4-1:0] node2785;
	wire [4-1:0] node2786;
	wire [4-1:0] node2787;
	wire [4-1:0] node2790;
	wire [4-1:0] node2793;
	wire [4-1:0] node2795;
	wire [4-1:0] node2796;
	wire [4-1:0] node2799;
	wire [4-1:0] node2802;
	wire [4-1:0] node2803;
	wire [4-1:0] node2806;
	wire [4-1:0] node2809;
	wire [4-1:0] node2810;
	wire [4-1:0] node2811;
	wire [4-1:0] node2812;
	wire [4-1:0] node2813;
	wire [4-1:0] node2815;
	wire [4-1:0] node2819;
	wire [4-1:0] node2820;
	wire [4-1:0] node2821;
	wire [4-1:0] node2824;
	wire [4-1:0] node2828;
	wire [4-1:0] node2829;
	wire [4-1:0] node2830;
	wire [4-1:0] node2833;
	wire [4-1:0] node2836;
	wire [4-1:0] node2837;
	wire [4-1:0] node2841;
	wire [4-1:0] node2842;
	wire [4-1:0] node2843;
	wire [4-1:0] node2844;
	wire [4-1:0] node2845;
	wire [4-1:0] node2846;
	wire [4-1:0] node2852;
	wire [4-1:0] node2853;
	wire [4-1:0] node2855;
	wire [4-1:0] node2856;
	wire [4-1:0] node2859;
	wire [4-1:0] node2863;
	wire [4-1:0] node2864;
	wire [4-1:0] node2866;
	wire [4-1:0] node2869;
	wire [4-1:0] node2870;
	wire [4-1:0] node2873;
	wire [4-1:0] node2876;
	wire [4-1:0] node2877;
	wire [4-1:0] node2878;
	wire [4-1:0] node2879;
	wire [4-1:0] node2880;
	wire [4-1:0] node2881;
	wire [4-1:0] node2884;
	wire [4-1:0] node2885;
	wire [4-1:0] node2887;
	wire [4-1:0] node2891;
	wire [4-1:0] node2892;
	wire [4-1:0] node2894;
	wire [4-1:0] node2895;
	wire [4-1:0] node2897;
	wire [4-1:0] node2900;
	wire [4-1:0] node2903;
	wire [4-1:0] node2906;
	wire [4-1:0] node2907;
	wire [4-1:0] node2908;
	wire [4-1:0] node2909;
	wire [4-1:0] node2910;
	wire [4-1:0] node2913;
	wire [4-1:0] node2915;
	wire [4-1:0] node2918;
	wire [4-1:0] node2919;
	wire [4-1:0] node2923;
	wire [4-1:0] node2924;
	wire [4-1:0] node2925;
	wire [4-1:0] node2928;
	wire [4-1:0] node2932;
	wire [4-1:0] node2933;
	wire [4-1:0] node2934;
	wire [4-1:0] node2936;
	wire [4-1:0] node2939;
	wire [4-1:0] node2941;
	wire [4-1:0] node2944;
	wire [4-1:0] node2945;
	wire [4-1:0] node2947;
	wire [4-1:0] node2950;
	wire [4-1:0] node2951;
	wire [4-1:0] node2954;
	wire [4-1:0] node2955;
	wire [4-1:0] node2959;
	wire [4-1:0] node2960;
	wire [4-1:0] node2961;
	wire [4-1:0] node2962;
	wire [4-1:0] node2964;
	wire [4-1:0] node2967;
	wire [4-1:0] node2968;
	wire [4-1:0] node2970;
	wire [4-1:0] node2973;
	wire [4-1:0] node2976;
	wire [4-1:0] node2977;
	wire [4-1:0] node2978;
	wire [4-1:0] node2979;
	wire [4-1:0] node2983;
	wire [4-1:0] node2984;
	wire [4-1:0] node2988;
	wire [4-1:0] node2991;
	wire [4-1:0] node2992;
	wire [4-1:0] node2993;
	wire [4-1:0] node2994;
	wire [4-1:0] node2997;
	wire [4-1:0] node3000;
	wire [4-1:0] node3001;
	wire [4-1:0] node3003;
	wire [4-1:0] node3005;
	wire [4-1:0] node3008;
	wire [4-1:0] node3010;
	wire [4-1:0] node3011;
	wire [4-1:0] node3015;
	wire [4-1:0] node3016;
	wire [4-1:0] node3017;
	wire [4-1:0] node3018;
	wire [4-1:0] node3022;
	wire [4-1:0] node3023;
	wire [4-1:0] node3027;
	wire [4-1:0] node3029;
	wire [4-1:0] node3032;
	wire [4-1:0] node3033;
	wire [4-1:0] node3034;
	wire [4-1:0] node3035;
	wire [4-1:0] node3036;
	wire [4-1:0] node3037;
	wire [4-1:0] node3039;
	wire [4-1:0] node3042;
	wire [4-1:0] node3046;
	wire [4-1:0] node3047;
	wire [4-1:0] node3048;
	wire [4-1:0] node3050;
	wire [4-1:0] node3054;
	wire [4-1:0] node3055;
	wire [4-1:0] node3056;
	wire [4-1:0] node3063;
	wire [4-1:0] node3064;
	wire [4-1:0] node3065;
	wire [4-1:0] node3066;
	wire [4-1:0] node3067;
	wire [4-1:0] node3068;
	wire [4-1:0] node3069;
	wire [4-1:0] node3070;
	wire [4-1:0] node3072;
	wire [4-1:0] node3075;
	wire [4-1:0] node3078;
	wire [4-1:0] node3079;
	wire [4-1:0] node3080;
	wire [4-1:0] node3084;
	wire [4-1:0] node3085;
	wire [4-1:0] node3088;
	wire [4-1:0] node3089;
	wire [4-1:0] node3093;
	wire [4-1:0] node3094;
	wire [4-1:0] node3095;
	wire [4-1:0] node3096;
	wire [4-1:0] node3098;
	wire [4-1:0] node3102;
	wire [4-1:0] node3103;
	wire [4-1:0] node3106;
	wire [4-1:0] node3108;
	wire [4-1:0] node3111;
	wire [4-1:0] node3112;
	wire [4-1:0] node3113;
	wire [4-1:0] node3117;
	wire [4-1:0] node3118;
	wire [4-1:0] node3121;
	wire [4-1:0] node3124;
	wire [4-1:0] node3125;
	wire [4-1:0] node3126;
	wire [4-1:0] node3127;
	wire [4-1:0] node3128;
	wire [4-1:0] node3131;
	wire [4-1:0] node3134;
	wire [4-1:0] node3136;
	wire [4-1:0] node3139;
	wire [4-1:0] node3142;
	wire [4-1:0] node3143;
	wire [4-1:0] node3145;
	wire [4-1:0] node3148;
	wire [4-1:0] node3149;
	wire [4-1:0] node3153;
	wire [4-1:0] node3154;
	wire [4-1:0] node3155;
	wire [4-1:0] node3156;
	wire [4-1:0] node3157;
	wire [4-1:0] node3158;
	wire [4-1:0] node3159;
	wire [4-1:0] node3164;
	wire [4-1:0] node3165;
	wire [4-1:0] node3169;
	wire [4-1:0] node3170;
	wire [4-1:0] node3171;
	wire [4-1:0] node3175;
	wire [4-1:0] node3176;
	wire [4-1:0] node3177;
	wire [4-1:0] node3182;
	wire [4-1:0] node3183;
	wire [4-1:0] node3184;
	wire [4-1:0] node3186;
	wire [4-1:0] node3189;
	wire [4-1:0] node3191;
	wire [4-1:0] node3194;
	wire [4-1:0] node3195;
	wire [4-1:0] node3199;
	wire [4-1:0] node3200;
	wire [4-1:0] node3201;
	wire [4-1:0] node3202;
	wire [4-1:0] node3203;
	wire [4-1:0] node3207;
	wire [4-1:0] node3210;
	wire [4-1:0] node3211;
	wire [4-1:0] node3212;
	wire [4-1:0] node3215;
	wire [4-1:0] node3216;
	wire [4-1:0] node3220;
	wire [4-1:0] node3221;
	wire [4-1:0] node3225;
	wire [4-1:0] node3226;
	wire [4-1:0] node3227;
	wire [4-1:0] node3228;
	wire [4-1:0] node3229;
	wire [4-1:0] node3234;
	wire [4-1:0] node3235;
	wire [4-1:0] node3239;
	wire [4-1:0] node3240;
	wire [4-1:0] node3242;
	wire [4-1:0] node3246;
	wire [4-1:0] node3247;
	wire [4-1:0] node3248;
	wire [4-1:0] node3249;
	wire [4-1:0] node3250;
	wire [4-1:0] node3251;
	wire [4-1:0] node3254;
	wire [4-1:0] node3257;
	wire [4-1:0] node3259;
	wire [4-1:0] node3262;
	wire [4-1:0] node3263;
	wire [4-1:0] node3264;
	wire [4-1:0] node3265;
	wire [4-1:0] node3269;
	wire [4-1:0] node3272;
	wire [4-1:0] node3273;
	wire [4-1:0] node3274;
	wire [4-1:0] node3277;
	wire [4-1:0] node3280;
	wire [4-1:0] node3281;
	wire [4-1:0] node3284;
	wire [4-1:0] node3287;
	wire [4-1:0] node3288;
	wire [4-1:0] node3289;
	wire [4-1:0] node3290;
	wire [4-1:0] node3291;
	wire [4-1:0] node3294;
	wire [4-1:0] node3298;
	wire [4-1:0] node3299;
	wire [4-1:0] node3303;
	wire [4-1:0] node3304;
	wire [4-1:0] node3306;
	wire [4-1:0] node3307;
	wire [4-1:0] node3311;
	wire [4-1:0] node3312;
	wire [4-1:0] node3315;
	wire [4-1:0] node3318;
	wire [4-1:0] node3319;
	wire [4-1:0] node3320;
	wire [4-1:0] node3321;
	wire [4-1:0] node3322;
	wire [4-1:0] node3325;
	wire [4-1:0] node3328;
	wire [4-1:0] node3329;
	wire [4-1:0] node3331;
	wire [4-1:0] node3334;
	wire [4-1:0] node3335;
	wire [4-1:0] node3339;
	wire [4-1:0] node3341;
	wire [4-1:0] node3342;
	wire [4-1:0] node3343;
	wire [4-1:0] node3348;
	wire [4-1:0] node3349;
	wire [4-1:0] node3350;
	wire [4-1:0] node3351;
	wire [4-1:0] node3355;
	wire [4-1:0] node3356;
	wire [4-1:0] node3359;
	wire [4-1:0] node3363;
	wire [4-1:0] node3364;
	wire [4-1:0] node3365;
	wire [4-1:0] node3366;
	wire [4-1:0] node3367;
	wire [4-1:0] node3368;
	wire [4-1:0] node3370;
	wire [4-1:0] node3371;
	wire [4-1:0] node3375;
	wire [4-1:0] node3376;
	wire [4-1:0] node3377;
	wire [4-1:0] node3379;
	wire [4-1:0] node3382;
	wire [4-1:0] node3385;
	wire [4-1:0] node3386;
	wire [4-1:0] node3390;
	wire [4-1:0] node3391;
	wire [4-1:0] node3392;
	wire [4-1:0] node3395;
	wire [4-1:0] node3396;
	wire [4-1:0] node3400;
	wire [4-1:0] node3401;
	wire [4-1:0] node3404;
	wire [4-1:0] node3405;
	wire [4-1:0] node3408;
	wire [4-1:0] node3411;
	wire [4-1:0] node3412;
	wire [4-1:0] node3413;
	wire [4-1:0] node3415;
	wire [4-1:0] node3416;
	wire [4-1:0] node3420;
	wire [4-1:0] node3421;
	wire [4-1:0] node3425;
	wire [4-1:0] node3426;
	wire [4-1:0] node3428;
	wire [4-1:0] node3430;
	wire [4-1:0] node3433;
	wire [4-1:0] node3434;
	wire [4-1:0] node3437;
	wire [4-1:0] node3440;
	wire [4-1:0] node3441;
	wire [4-1:0] node3442;
	wire [4-1:0] node3443;
	wire [4-1:0] node3444;
	wire [4-1:0] node3447;
	wire [4-1:0] node3448;
	wire [4-1:0] node3452;
	wire [4-1:0] node3453;
	wire [4-1:0] node3455;
	wire [4-1:0] node3459;
	wire [4-1:0] node3460;
	wire [4-1:0] node3461;
	wire [4-1:0] node3462;
	wire [4-1:0] node3463;
	wire [4-1:0] node3468;
	wire [4-1:0] node3471;
	wire [4-1:0] node3472;
	wire [4-1:0] node3474;
	wire [4-1:0] node3478;
	wire [4-1:0] node3479;
	wire [4-1:0] node3480;
	wire [4-1:0] node3481;
	wire [4-1:0] node3482;
	wire [4-1:0] node3483;
	wire [4-1:0] node3488;
	wire [4-1:0] node3489;
	wire [4-1:0] node3490;
	wire [4-1:0] node3494;
	wire [4-1:0] node3497;
	wire [4-1:0] node3498;
	wire [4-1:0] node3499;
	wire [4-1:0] node3501;
	wire [4-1:0] node3505;
	wire [4-1:0] node3508;
	wire [4-1:0] node3509;
	wire [4-1:0] node3510;
	wire [4-1:0] node3513;
	wire [4-1:0] node3517;
	wire [4-1:0] node3518;
	wire [4-1:0] node3519;
	wire [4-1:0] node3520;
	wire [4-1:0] node3521;
	wire [4-1:0] node3522;
	wire [4-1:0] node3526;
	wire [4-1:0] node3528;
	wire [4-1:0] node3531;
	wire [4-1:0] node3532;
	wire [4-1:0] node3533;
	wire [4-1:0] node3537;
	wire [4-1:0] node3538;
	wire [4-1:0] node3542;
	wire [4-1:0] node3543;
	wire [4-1:0] node3544;
	wire [4-1:0] node3546;
	wire [4-1:0] node3547;
	wire [4-1:0] node3551;
	wire [4-1:0] node3552;
	wire [4-1:0] node3556;
	wire [4-1:0] node3557;
	wire [4-1:0] node3558;
	wire [4-1:0] node3562;
	wire [4-1:0] node3563;
	wire [4-1:0] node3565;
	wire [4-1:0] node3570;
	wire [4-1:0] node3571;
	wire [4-1:0] node3572;
	wire [4-1:0] node3573;
	wire [4-1:0] node3574;
	wire [4-1:0] node3575;
	wire [4-1:0] node3576;
	wire [4-1:0] node3577;
	wire [4-1:0] node3578;
	wire [4-1:0] node3579;
	wire [4-1:0] node3583;
	wire [4-1:0] node3586;
	wire [4-1:0] node3587;
	wire [4-1:0] node3588;
	wire [4-1:0] node3589;
	wire [4-1:0] node3593;
	wire [4-1:0] node3596;
	wire [4-1:0] node3597;
	wire [4-1:0] node3600;
	wire [4-1:0] node3601;
	wire [4-1:0] node3604;
	wire [4-1:0] node3607;
	wire [4-1:0] node3608;
	wire [4-1:0] node3609;
	wire [4-1:0] node3610;
	wire [4-1:0] node3611;
	wire [4-1:0] node3614;
	wire [4-1:0] node3619;
	wire [4-1:0] node3620;
	wire [4-1:0] node3623;
	wire [4-1:0] node3624;
	wire [4-1:0] node3627;
	wire [4-1:0] node3629;
	wire [4-1:0] node3632;
	wire [4-1:0] node3633;
	wire [4-1:0] node3634;
	wire [4-1:0] node3635;
	wire [4-1:0] node3636;
	wire [4-1:0] node3638;
	wire [4-1:0] node3641;
	wire [4-1:0] node3643;
	wire [4-1:0] node3647;
	wire [4-1:0] node3648;
	wire [4-1:0] node3649;
	wire [4-1:0] node3652;
	wire [4-1:0] node3656;
	wire [4-1:0] node3657;
	wire [4-1:0] node3658;
	wire [4-1:0] node3659;
	wire [4-1:0] node3664;
	wire [4-1:0] node3665;
	wire [4-1:0] node3668;
	wire [4-1:0] node3669;
	wire [4-1:0] node3672;
	wire [4-1:0] node3674;
	wire [4-1:0] node3677;
	wire [4-1:0] node3678;
	wire [4-1:0] node3679;
	wire [4-1:0] node3680;
	wire [4-1:0] node3681;
	wire [4-1:0] node3682;
	wire [4-1:0] node3683;
	wire [4-1:0] node3688;
	wire [4-1:0] node3691;
	wire [4-1:0] node3692;
	wire [4-1:0] node3693;
	wire [4-1:0] node3695;
	wire [4-1:0] node3699;
	wire [4-1:0] node3700;
	wire [4-1:0] node3704;
	wire [4-1:0] node3705;
	wire [4-1:0] node3706;
	wire [4-1:0] node3708;
	wire [4-1:0] node3711;
	wire [4-1:0] node3712;
	wire [4-1:0] node3716;
	wire [4-1:0] node3718;
	wire [4-1:0] node3721;
	wire [4-1:0] node3722;
	wire [4-1:0] node3723;
	wire [4-1:0] node3724;
	wire [4-1:0] node3726;
	wire [4-1:0] node3729;
	wire [4-1:0] node3730;
	wire [4-1:0] node3734;
	wire [4-1:0] node3736;
	wire [4-1:0] node3737;
	wire [4-1:0] node3741;
	wire [4-1:0] node3742;
	wire [4-1:0] node3743;
	wire [4-1:0] node3744;
	wire [4-1:0] node3745;
	wire [4-1:0] node3750;
	wire [4-1:0] node3751;
	wire [4-1:0] node3754;
	wire [4-1:0] node3757;
	wire [4-1:0] node3758;
	wire [4-1:0] node3759;
	wire [4-1:0] node3763;
	wire [4-1:0] node3765;
	wire [4-1:0] node3766;
	wire [4-1:0] node3770;
	wire [4-1:0] node3771;
	wire [4-1:0] node3772;
	wire [4-1:0] node3773;
	wire [4-1:0] node3774;
	wire [4-1:0] node3775;
	wire [4-1:0] node3777;
	wire [4-1:0] node3780;
	wire [4-1:0] node3781;
	wire [4-1:0] node3785;
	wire [4-1:0] node3786;
	wire [4-1:0] node3788;
	wire [4-1:0] node3789;
	wire [4-1:0] node3793;
	wire [4-1:0] node3794;
	wire [4-1:0] node3798;
	wire [4-1:0] node3799;
	wire [4-1:0] node3800;
	wire [4-1:0] node3802;
	wire [4-1:0] node3805;
	wire [4-1:0] node3807;
	wire [4-1:0] node3809;
	wire [4-1:0] node3812;
	wire [4-1:0] node3813;
	wire [4-1:0] node3814;
	wire [4-1:0] node3819;
	wire [4-1:0] node3820;
	wire [4-1:0] node3821;
	wire [4-1:0] node3822;
	wire [4-1:0] node3823;
	wire [4-1:0] node3825;
	wire [4-1:0] node3828;
	wire [4-1:0] node3829;
	wire [4-1:0] node3832;
	wire [4-1:0] node3835;
	wire [4-1:0] node3838;
	wire [4-1:0] node3839;
	wire [4-1:0] node3841;
	wire [4-1:0] node3842;
	wire [4-1:0] node3846;
	wire [4-1:0] node3847;
	wire [4-1:0] node3850;
	wire [4-1:0] node3853;
	wire [4-1:0] node3855;
	wire [4-1:0] node3858;
	wire [4-1:0] node3859;
	wire [4-1:0] node3860;
	wire [4-1:0] node3861;
	wire [4-1:0] node3862;
	wire [4-1:0] node3863;
	wire [4-1:0] node3864;
	wire [4-1:0] node3867;
	wire [4-1:0] node3871;
	wire [4-1:0] node3873;
	wire [4-1:0] node3876;
	wire [4-1:0] node3877;
	wire [4-1:0] node3878;
	wire [4-1:0] node3882;
	wire [4-1:0] node3884;
	wire [4-1:0] node3887;
	wire [4-1:0] node3888;
	wire [4-1:0] node3889;
	wire [4-1:0] node3890;
	wire [4-1:0] node3892;
	wire [4-1:0] node3895;
	wire [4-1:0] node3898;
	wire [4-1:0] node3899;
	wire [4-1:0] node3900;
	wire [4-1:0] node3904;
	wire [4-1:0] node3907;
	wire [4-1:0] node3908;
	wire [4-1:0] node3909;
	wire [4-1:0] node3913;
	wire [4-1:0] node3914;
	wire [4-1:0] node3917;
	wire [4-1:0] node3920;
	wire [4-1:0] node3921;
	wire [4-1:0] node3922;
	wire [4-1:0] node3923;
	wire [4-1:0] node3926;
	wire [4-1:0] node3928;
	wire [4-1:0] node3931;
	wire [4-1:0] node3932;
	wire [4-1:0] node3935;
	wire [4-1:0] node3939;
	wire [4-1:0] node3940;
	wire [4-1:0] node3941;
	wire [4-1:0] node3942;
	wire [4-1:0] node3943;
	wire [4-1:0] node3944;
	wire [4-1:0] node3946;
	wire [4-1:0] node3949;
	wire [4-1:0] node3950;
	wire [4-1:0] node3952;
	wire [4-1:0] node3955;
	wire [4-1:0] node3956;
	wire [4-1:0] node3960;
	wire [4-1:0] node3961;
	wire [4-1:0] node3962;
	wire [4-1:0] node3963;
	wire [4-1:0] node3967;
	wire [4-1:0] node3970;
	wire [4-1:0] node3971;
	wire [4-1:0] node3973;
	wire [4-1:0] node3976;
	wire [4-1:0] node3977;
	wire [4-1:0] node3980;
	wire [4-1:0] node3983;
	wire [4-1:0] node3984;
	wire [4-1:0] node3985;
	wire [4-1:0] node3986;
	wire [4-1:0] node3987;
	wire [4-1:0] node3991;
	wire [4-1:0] node3994;
	wire [4-1:0] node3995;
	wire [4-1:0] node3999;
	wire [4-1:0] node4000;
	wire [4-1:0] node4001;
	wire [4-1:0] node4002;
	wire [4-1:0] node4006;
	wire [4-1:0] node4008;
	wire [4-1:0] node4011;
	wire [4-1:0] node4012;
	wire [4-1:0] node4015;
	wire [4-1:0] node4018;
	wire [4-1:0] node4019;
	wire [4-1:0] node4020;
	wire [4-1:0] node4022;
	wire [4-1:0] node4024;
	wire [4-1:0] node4025;
	wire [4-1:0] node4028;
	wire [4-1:0] node4031;
	wire [4-1:0] node4032;
	wire [4-1:0] node4035;
	wire [4-1:0] node4036;
	wire [4-1:0] node4037;
	wire [4-1:0] node4041;
	wire [4-1:0] node4042;
	wire [4-1:0] node4045;
	wire [4-1:0] node4048;
	wire [4-1:0] node4049;
	wire [4-1:0] node4050;
	wire [4-1:0] node4051;
	wire [4-1:0] node4055;
	wire [4-1:0] node4056;
	wire [4-1:0] node4058;
	wire [4-1:0] node4062;
	wire [4-1:0] node4063;
	wire [4-1:0] node4064;
	wire [4-1:0] node4068;
	wire [4-1:0] node4069;
	wire [4-1:0] node4070;
	wire [4-1:0] node4075;
	wire [4-1:0] node4076;
	wire [4-1:0] node4077;
	wire [4-1:0] node4078;
	wire [4-1:0] node4079;
	wire [4-1:0] node4080;
	wire [4-1:0] node4081;
	wire [4-1:0] node4085;
	wire [4-1:0] node4088;
	wire [4-1:0] node4089;
	wire [4-1:0] node4092;
	wire [4-1:0] node4093;
	wire [4-1:0] node4097;
	wire [4-1:0] node4099;
	wire [4-1:0] node4100;
	wire [4-1:0] node4101;
	wire [4-1:0] node4105;
	wire [4-1:0] node4107;
	wire [4-1:0] node4110;
	wire [4-1:0] node4111;
	wire [4-1:0] node4112;
	wire [4-1:0] node4114;
	wire [4-1:0] node4117;
	wire [4-1:0] node4118;
	wire [4-1:0] node4119;
	wire [4-1:0] node4122;
	wire [4-1:0] node4126;
	wire [4-1:0] node4127;
	wire [4-1:0] node4128;
	wire [4-1:0] node4129;
	wire [4-1:0] node4134;
	wire [4-1:0] node4135;
	wire [4-1:0] node4139;
	wire [4-1:0] node4140;
	wire [4-1:0] node4141;
	wire [4-1:0] node4142;
	wire [4-1:0] node4144;
	wire [4-1:0] node4147;
	wire [4-1:0] node4149;
	wire [4-1:0] node4150;
	wire [4-1:0] node4154;
	wire [4-1:0] node4155;
	wire [4-1:0] node4157;
	wire [4-1:0] node4160;
	wire [4-1:0] node4162;
	wire [4-1:0] node4163;
	wire [4-1:0] node4166;
	wire [4-1:0] node4167;
	wire [4-1:0] node4172;
	wire [4-1:0] node4173;
	wire [4-1:0] node4174;
	wire [4-1:0] node4175;
	wire [4-1:0] node4176;
	wire [4-1:0] node4177;
	wire [4-1:0] node4178;
	wire [4-1:0] node4179;
	wire [4-1:0] node4180;
	wire [4-1:0] node4182;
	wire [4-1:0] node4187;
	wire [4-1:0] node4188;
	wire [4-1:0] node4189;
	wire [4-1:0] node4190;
	wire [4-1:0] node4194;
	wire [4-1:0] node4197;
	wire [4-1:0] node4198;
	wire [4-1:0] node4201;
	wire [4-1:0] node4202;
	wire [4-1:0] node4206;
	wire [4-1:0] node4207;
	wire [4-1:0] node4208;
	wire [4-1:0] node4210;
	wire [4-1:0] node4211;
	wire [4-1:0] node4215;
	wire [4-1:0] node4217;
	wire [4-1:0] node4220;
	wire [4-1:0] node4221;
	wire [4-1:0] node4224;
	wire [4-1:0] node4226;
	wire [4-1:0] node4229;
	wire [4-1:0] node4230;
	wire [4-1:0] node4231;
	wire [4-1:0] node4232;
	wire [4-1:0] node4235;
	wire [4-1:0] node4237;
	wire [4-1:0] node4240;
	wire [4-1:0] node4241;
	wire [4-1:0] node4245;
	wire [4-1:0] node4246;
	wire [4-1:0] node4247;
	wire [4-1:0] node4248;
	wire [4-1:0] node4252;
	wire [4-1:0] node4255;
	wire [4-1:0] node4256;
	wire [4-1:0] node4260;
	wire [4-1:0] node4261;
	wire [4-1:0] node4262;
	wire [4-1:0] node4263;
	wire [4-1:0] node4264;
	wire [4-1:0] node4266;
	wire [4-1:0] node4270;
	wire [4-1:0] node4272;
	wire [4-1:0] node4273;
	wire [4-1:0] node4274;
	wire [4-1:0] node4279;
	wire [4-1:0] node4280;
	wire [4-1:0] node4281;
	wire [4-1:0] node4282;
	wire [4-1:0] node4283;
	wire [4-1:0] node4287;
	wire [4-1:0] node4288;
	wire [4-1:0] node4292;
	wire [4-1:0] node4294;
	wire [4-1:0] node4296;
	wire [4-1:0] node4299;
	wire [4-1:0] node4301;
	wire [4-1:0] node4302;
	wire [4-1:0] node4306;
	wire [4-1:0] node4307;
	wire [4-1:0] node4308;
	wire [4-1:0] node4309;
	wire [4-1:0] node4311;
	wire [4-1:0] node4312;
	wire [4-1:0] node4316;
	wire [4-1:0] node4319;
	wire [4-1:0] node4320;
	wire [4-1:0] node4323;
	wire [4-1:0] node4325;
	wire [4-1:0] node4328;
	wire [4-1:0] node4329;
	wire [4-1:0] node4330;
	wire [4-1:0] node4332;
	wire [4-1:0] node4335;
	wire [4-1:0] node4336;
	wire [4-1:0] node4339;
	wire [4-1:0] node4340;
	wire [4-1:0] node4344;
	wire [4-1:0] node4345;
	wire [4-1:0] node4347;
	wire [4-1:0] node4349;
	wire [4-1:0] node4352;
	wire [4-1:0] node4354;
	wire [4-1:0] node4356;
	wire [4-1:0] node4359;
	wire [4-1:0] node4360;
	wire [4-1:0] node4361;
	wire [4-1:0] node4362;
	wire [4-1:0] node4363;
	wire [4-1:0] node4364;
	wire [4-1:0] node4365;
	wire [4-1:0] node4367;
	wire [4-1:0] node4371;
	wire [4-1:0] node4372;
	wire [4-1:0] node4376;
	wire [4-1:0] node4377;
	wire [4-1:0] node4378;
	wire [4-1:0] node4380;
	wire [4-1:0] node4383;
	wire [4-1:0] node4387;
	wire [4-1:0] node4388;
	wire [4-1:0] node4389;
	wire [4-1:0] node4391;
	wire [4-1:0] node4394;
	wire [4-1:0] node4395;
	wire [4-1:0] node4399;
	wire [4-1:0] node4400;
	wire [4-1:0] node4403;
	wire [4-1:0] node4406;
	wire [4-1:0] node4407;
	wire [4-1:0] node4408;
	wire [4-1:0] node4409;
	wire [4-1:0] node4413;
	wire [4-1:0] node4414;
	wire [4-1:0] node4415;
	wire [4-1:0] node4416;
	wire [4-1:0] node4419;
	wire [4-1:0] node4422;
	wire [4-1:0] node4423;
	wire [4-1:0] node4426;
	wire [4-1:0] node4429;
	wire [4-1:0] node4431;
	wire [4-1:0] node4434;
	wire [4-1:0] node4435;
	wire [4-1:0] node4436;
	wire [4-1:0] node4438;
	wire [4-1:0] node4441;
	wire [4-1:0] node4442;
	wire [4-1:0] node4446;
	wire [4-1:0] node4447;
	wire [4-1:0] node4448;
	wire [4-1:0] node4451;
	wire [4-1:0] node4454;
	wire [4-1:0] node4455;
	wire [4-1:0] node4458;
	wire [4-1:0] node4461;
	wire [4-1:0] node4462;
	wire [4-1:0] node4463;
	wire [4-1:0] node4464;
	wire [4-1:0] node4465;
	wire [4-1:0] node4467;
	wire [4-1:0] node4471;
	wire [4-1:0] node4472;
	wire [4-1:0] node4474;
	wire [4-1:0] node4477;
	wire [4-1:0] node4478;
	wire [4-1:0] node4482;
	wire [4-1:0] node4483;
	wire [4-1:0] node4484;
	wire [4-1:0] node4485;
	wire [4-1:0] node4488;
	wire [4-1:0] node4491;
	wire [4-1:0] node4493;
	wire [4-1:0] node4496;
	wire [4-1:0] node4497;
	wire [4-1:0] node4499;
	wire [4-1:0] node4504;
	wire [4-1:0] node4505;
	wire [4-1:0] node4506;
	wire [4-1:0] node4507;
	wire [4-1:0] node4508;
	wire [4-1:0] node4509;
	wire [4-1:0] node4510;
	wire [4-1:0] node4514;
	wire [4-1:0] node4515;
	wire [4-1:0] node4516;
	wire [4-1:0] node4520;
	wire [4-1:0] node4521;
	wire [4-1:0] node4525;
	wire [4-1:0] node4526;
	wire [4-1:0] node4527;
	wire [4-1:0] node4528;
	wire [4-1:0] node4532;
	wire [4-1:0] node4533;
	wire [4-1:0] node4537;
	wire [4-1:0] node4538;
	wire [4-1:0] node4539;
	wire [4-1:0] node4543;
	wire [4-1:0] node4545;
	wire [4-1:0] node4546;
	wire [4-1:0] node4550;
	wire [4-1:0] node4551;
	wire [4-1:0] node4552;
	wire [4-1:0] node4553;
	wire [4-1:0] node4555;
	wire [4-1:0] node4556;
	wire [4-1:0] node4559;
	wire [4-1:0] node4563;
	wire [4-1:0] node4565;
	wire [4-1:0] node4568;
	wire [4-1:0] node4569;
	wire [4-1:0] node4570;
	wire [4-1:0] node4572;
	wire [4-1:0] node4575;
	wire [4-1:0] node4577;
	wire [4-1:0] node4580;
	wire [4-1:0] node4581;
	wire [4-1:0] node4584;
	wire [4-1:0] node4586;
	wire [4-1:0] node4589;
	wire [4-1:0] node4590;
	wire [4-1:0] node4591;
	wire [4-1:0] node4592;
	wire [4-1:0] node4594;
	wire [4-1:0] node4596;
	wire [4-1:0] node4599;
	wire [4-1:0] node4600;
	wire [4-1:0] node4604;
	wire [4-1:0] node4605;
	wire [4-1:0] node4606;
	wire [4-1:0] node4607;
	wire [4-1:0] node4610;
	wire [4-1:0] node4614;
	wire [4-1:0] node4616;
	wire [4-1:0] node4618;
	wire [4-1:0] node4622;
	wire [4-1:0] node4623;
	wire [4-1:0] node4624;
	wire [4-1:0] node4625;
	wire [4-1:0] node4626;
	wire [4-1:0] node4628;
	wire [4-1:0] node4629;
	wire [4-1:0] node4632;
	wire [4-1:0] node4635;
	wire [4-1:0] node4636;
	wire [4-1:0] node4637;
	wire [4-1:0] node4642;
	wire [4-1:0] node4643;
	wire [4-1:0] node4644;
	wire [4-1:0] node4645;
	wire [4-1:0] node4646;
	wire [4-1:0] node4649;
	wire [4-1:0] node4654;
	wire [4-1:0] node4655;
	wire [4-1:0] node4658;
	wire [4-1:0] node4659;
	wire [4-1:0] node4660;
	wire [4-1:0] node4667;
	wire [4-1:0] node4668;
	wire [4-1:0] node4669;
	wire [4-1:0] node4670;
	wire [4-1:0] node4671;
	wire [4-1:0] node4672;
	wire [4-1:0] node4673;
	wire [4-1:0] node4674;
	wire [4-1:0] node4675;
	wire [4-1:0] node4677;
	wire [4-1:0] node4678;
	wire [4-1:0] node4679;
	wire [4-1:0] node4683;
	wire [4-1:0] node4685;
	wire [4-1:0] node4687;
	wire [4-1:0] node4688;
	wire [4-1:0] node4691;
	wire [4-1:0] node4694;
	wire [4-1:0] node4695;
	wire [4-1:0] node4696;
	wire [4-1:0] node4698;
	wire [4-1:0] node4699;
	wire [4-1:0] node4700;
	wire [4-1:0] node4704;
	wire [4-1:0] node4707;
	wire [4-1:0] node4708;
	wire [4-1:0] node4709;
	wire [4-1:0] node4710;
	wire [4-1:0] node4716;
	wire [4-1:0] node4717;
	wire [4-1:0] node4719;
	wire [4-1:0] node4722;
	wire [4-1:0] node4723;
	wire [4-1:0] node4724;
	wire [4-1:0] node4729;
	wire [4-1:0] node4731;
	wire [4-1:0] node4733;
	wire [4-1:0] node4734;
	wire [4-1:0] node4736;
	wire [4-1:0] node4737;
	wire [4-1:0] node4738;
	wire [4-1:0] node4742;
	wire [4-1:0] node4743;
	wire [4-1:0] node4746;
	wire [4-1:0] node4749;
	wire [4-1:0] node4751;
	wire [4-1:0] node4754;
	wire [4-1:0] node4755;
	wire [4-1:0] node4756;
	wire [4-1:0] node4757;
	wire [4-1:0] node4758;
	wire [4-1:0] node4759;
	wire [4-1:0] node4763;
	wire [4-1:0] node4766;
	wire [4-1:0] node4767;
	wire [4-1:0] node4770;
	wire [4-1:0] node4771;
	wire [4-1:0] node4773;
	wire [4-1:0] node4776;
	wire [4-1:0] node4777;
	wire [4-1:0] node4780;
	wire [4-1:0] node4783;
	wire [4-1:0] node4784;
	wire [4-1:0] node4785;
	wire [4-1:0] node4786;
	wire [4-1:0] node4790;
	wire [4-1:0] node4791;
	wire [4-1:0] node4793;
	wire [4-1:0] node4797;
	wire [4-1:0] node4798;
	wire [4-1:0] node4799;
	wire [4-1:0] node4801;
	wire [4-1:0] node4804;
	wire [4-1:0] node4807;
	wire [4-1:0] node4809;
	wire [4-1:0] node4812;
	wire [4-1:0] node4813;
	wire [4-1:0] node4814;
	wire [4-1:0] node4815;
	wire [4-1:0] node4816;
	wire [4-1:0] node4817;
	wire [4-1:0] node4821;
	wire [4-1:0] node4823;
	wire [4-1:0] node4826;
	wire [4-1:0] node4828;
	wire [4-1:0] node4831;
	wire [4-1:0] node4832;
	wire [4-1:0] node4833;
	wire [4-1:0] node4836;
	wire [4-1:0] node4839;
	wire [4-1:0] node4840;
	wire [4-1:0] node4844;
	wire [4-1:0] node4845;
	wire [4-1:0] node4846;
	wire [4-1:0] node4847;
	wire [4-1:0] node4851;
	wire [4-1:0] node4852;
	wire [4-1:0] node4856;
	wire [4-1:0] node4857;
	wire [4-1:0] node4859;
	wire [4-1:0] node4860;
	wire [4-1:0] node4862;
	wire [4-1:0] node4866;
	wire [4-1:0] node4867;
	wire [4-1:0] node4868;
	wire [4-1:0] node4869;
	wire [4-1:0] node4872;
	wire [4-1:0] node4878;
	wire [4-1:0] node4879;
	wire [4-1:0] node4880;
	wire [4-1:0] node4881;
	wire [4-1:0] node4882;
	wire [4-1:0] node4883;
	wire [4-1:0] node4884;
	wire [4-1:0] node4886;
	wire [4-1:0] node4889;
	wire [4-1:0] node4891;
	wire [4-1:0] node4892;
	wire [4-1:0] node4896;
	wire [4-1:0] node4897;
	wire [4-1:0] node4898;
	wire [4-1:0] node4902;
	wire [4-1:0] node4903;
	wire [4-1:0] node4907;
	wire [4-1:0] node4908;
	wire [4-1:0] node4909;
	wire [4-1:0] node4912;
	wire [4-1:0] node4915;
	wire [4-1:0] node4916;
	wire [4-1:0] node4918;
	wire [4-1:0] node4921;
	wire [4-1:0] node4924;
	wire [4-1:0] node4925;
	wire [4-1:0] node4926;
	wire [4-1:0] node4927;
	wire [4-1:0] node4928;
	wire [4-1:0] node4931;
	wire [4-1:0] node4932;
	wire [4-1:0] node4936;
	wire [4-1:0] node4937;
	wire [4-1:0] node4941;
	wire [4-1:0] node4942;
	wire [4-1:0] node4943;
	wire [4-1:0] node4944;
	wire [4-1:0] node4949;
	wire [4-1:0] node4950;
	wire [4-1:0] node4951;
	wire [4-1:0] node4955;
	wire [4-1:0] node4956;
	wire [4-1:0] node4960;
	wire [4-1:0] node4961;
	wire [4-1:0] node4962;
	wire [4-1:0] node4963;
	wire [4-1:0] node4964;
	wire [4-1:0] node4967;
	wire [4-1:0] node4969;
	wire [4-1:0] node4972;
	wire [4-1:0] node4975;
	wire [4-1:0] node4976;
	wire [4-1:0] node4979;
	wire [4-1:0] node4980;
	wire [4-1:0] node4982;
	wire [4-1:0] node4986;
	wire [4-1:0] node4987;
	wire [4-1:0] node4988;
	wire [4-1:0] node4989;
	wire [4-1:0] node4991;
	wire [4-1:0] node4994;
	wire [4-1:0] node4996;
	wire [4-1:0] node5000;
	wire [4-1:0] node5001;
	wire [4-1:0] node5005;
	wire [4-1:0] node5006;
	wire [4-1:0] node5007;
	wire [4-1:0] node5008;
	wire [4-1:0] node5010;
	wire [4-1:0] node5011;
	wire [4-1:0] node5012;
	wire [4-1:0] node5017;
	wire [4-1:0] node5018;
	wire [4-1:0] node5019;
	wire [4-1:0] node5022;
	wire [4-1:0] node5023;
	wire [4-1:0] node5027;
	wire [4-1:0] node5028;
	wire [4-1:0] node5031;
	wire [4-1:0] node5034;
	wire [4-1:0] node5036;
	wire [4-1:0] node5038;
	wire [4-1:0] node5040;
	wire [4-1:0] node5042;
	wire [4-1:0] node5045;
	wire [4-1:0] node5046;
	wire [4-1:0] node5047;
	wire [4-1:0] node5048;
	wire [4-1:0] node5049;
	wire [4-1:0] node5052;
	wire [4-1:0] node5055;
	wire [4-1:0] node5056;
	wire [4-1:0] node5060;
	wire [4-1:0] node5061;
	wire [4-1:0] node5063;
	wire [4-1:0] node5066;
	wire [4-1:0] node5067;
	wire [4-1:0] node5069;
	wire [4-1:0] node5073;
	wire [4-1:0] node5074;
	wire [4-1:0] node5075;
	wire [4-1:0] node5076;
	wire [4-1:0] node5077;
	wire [4-1:0] node5080;
	wire [4-1:0] node5084;
	wire [4-1:0] node5085;
	wire [4-1:0] node5087;
	wire [4-1:0] node5090;
	wire [4-1:0] node5091;
	wire [4-1:0] node5095;
	wire [4-1:0] node5096;
	wire [4-1:0] node5097;
	wire [4-1:0] node5098;
	wire [4-1:0] node5102;
	wire [4-1:0] node5103;
	wire [4-1:0] node5107;
	wire [4-1:0] node5110;
	wire [4-1:0] node5111;
	wire [4-1:0] node5112;
	wire [4-1:0] node5113;
	wire [4-1:0] node5114;
	wire [4-1:0] node5115;
	wire [4-1:0] node5117;
	wire [4-1:0] node5120;
	wire [4-1:0] node5121;
	wire [4-1:0] node5123;
	wire [4-1:0] node5127;
	wire [4-1:0] node5129;
	wire [4-1:0] node5130;
	wire [4-1:0] node5134;
	wire [4-1:0] node5135;
	wire [4-1:0] node5136;
	wire [4-1:0] node5138;
	wire [4-1:0] node5141;
	wire [4-1:0] node5143;
	wire [4-1:0] node5146;
	wire [4-1:0] node5148;
	wire [4-1:0] node5151;
	wire [4-1:0] node5152;
	wire [4-1:0] node5153;
	wire [4-1:0] node5154;
	wire [4-1:0] node5156;
	wire [4-1:0] node5160;
	wire [4-1:0] node5162;
	wire [4-1:0] node5165;
	wire [4-1:0] node5166;
	wire [4-1:0] node5167;
	wire [4-1:0] node5169;
	wire [4-1:0] node5170;
	wire [4-1:0] node5173;
	wire [4-1:0] node5176;
	wire [4-1:0] node5177;
	wire [4-1:0] node5179;
	wire [4-1:0] node5182;
	wire [4-1:0] node5185;
	wire [4-1:0] node5186;
	wire [4-1:0] node5188;
	wire [4-1:0] node5191;
	wire [4-1:0] node5192;
	wire [4-1:0] node5196;
	wire [4-1:0] node5197;
	wire [4-1:0] node5198;
	wire [4-1:0] node5199;
	wire [4-1:0] node5200;
	wire [4-1:0] node5202;
	wire [4-1:0] node5205;
	wire [4-1:0] node5206;
	wire [4-1:0] node5207;
	wire [4-1:0] node5209;
	wire [4-1:0] node5213;
	wire [4-1:0] node5216;
	wire [4-1:0] node5217;
	wire [4-1:0] node5218;
	wire [4-1:0] node5222;
	wire [4-1:0] node5223;
	wire [4-1:0] node5226;
	wire [4-1:0] node5228;
	wire [4-1:0] node5229;
	wire [4-1:0] node5232;
	wire [4-1:0] node5235;
	wire [4-1:0] node5236;
	wire [4-1:0] node5237;
	wire [4-1:0] node5238;
	wire [4-1:0] node5239;
	wire [4-1:0] node5244;
	wire [4-1:0] node5245;
	wire [4-1:0] node5247;
	wire [4-1:0] node5248;
	wire [4-1:0] node5251;
	wire [4-1:0] node5254;
	wire [4-1:0] node5256;
	wire [4-1:0] node5257;
	wire [4-1:0] node5261;
	wire [4-1:0] node5262;
	wire [4-1:0] node5263;
	wire [4-1:0] node5265;
	wire [4-1:0] node5266;
	wire [4-1:0] node5270;
	wire [4-1:0] node5273;
	wire [4-1:0] node5275;
	wire [4-1:0] node5276;
	wire [4-1:0] node5279;
	wire [4-1:0] node5282;
	wire [4-1:0] node5283;
	wire [4-1:0] node5284;
	wire [4-1:0] node5285;
	wire [4-1:0] node5286;
	wire [4-1:0] node5289;
	wire [4-1:0] node5290;
	wire [4-1:0] node5291;
	wire [4-1:0] node5295;
	wire [4-1:0] node5296;
	wire [4-1:0] node5299;
	wire [4-1:0] node5302;
	wire [4-1:0] node5304;
	wire [4-1:0] node5305;
	wire [4-1:0] node5309;
	wire [4-1:0] node5310;
	wire [4-1:0] node5311;
	wire [4-1:0] node5312;
	wire [4-1:0] node5313;
	wire [4-1:0] node5318;
	wire [4-1:0] node5320;
	wire [4-1:0] node5321;
	wire [4-1:0] node5325;
	wire [4-1:0] node5326;
	wire [4-1:0] node5327;
	wire [4-1:0] node5330;
	wire [4-1:0] node5333;
	wire [4-1:0] node5336;
	wire [4-1:0] node5337;
	wire [4-1:0] node5338;
	wire [4-1:0] node5339;
	wire [4-1:0] node5342;
	wire [4-1:0] node5343;
	wire [4-1:0] node5347;
	wire [4-1:0] node5349;
	wire [4-1:0] node5352;
	wire [4-1:0] node5353;
	wire [4-1:0] node5354;
	wire [4-1:0] node5355;
	wire [4-1:0] node5359;
	wire [4-1:0] node5361;
	wire [4-1:0] node5362;
	wire [4-1:0] node5366;
	wire [4-1:0] node5370;
	wire [4-1:0] node5371;
	wire [4-1:0] node5372;
	wire [4-1:0] node5373;
	wire [4-1:0] node5374;
	wire [4-1:0] node5375;
	wire [4-1:0] node5376;
	wire [4-1:0] node5377;
	wire [4-1:0] node5378;
	wire [4-1:0] node5380;
	wire [4-1:0] node5383;
	wire [4-1:0] node5385;
	wire [4-1:0] node5388;
	wire [4-1:0] node5389;
	wire [4-1:0] node5391;
	wire [4-1:0] node5392;
	wire [4-1:0] node5395;
	wire [4-1:0] node5396;
	wire [4-1:0] node5400;
	wire [4-1:0] node5401;
	wire [4-1:0] node5403;
	wire [4-1:0] node5404;
	wire [4-1:0] node5408;
	wire [4-1:0] node5409;
	wire [4-1:0] node5412;
	wire [4-1:0] node5415;
	wire [4-1:0] node5416;
	wire [4-1:0] node5417;
	wire [4-1:0] node5418;
	wire [4-1:0] node5421;
	wire [4-1:0] node5423;
	wire [4-1:0] node5426;
	wire [4-1:0] node5428;
	wire [4-1:0] node5431;
	wire [4-1:0] node5432;
	wire [4-1:0] node5433;
	wire [4-1:0] node5434;
	wire [4-1:0] node5438;
	wire [4-1:0] node5439;
	wire [4-1:0] node5443;
	wire [4-1:0] node5444;
	wire [4-1:0] node5446;
	wire [4-1:0] node5449;
	wire [4-1:0] node5450;
	wire [4-1:0] node5453;
	wire [4-1:0] node5456;
	wire [4-1:0] node5457;
	wire [4-1:0] node5458;
	wire [4-1:0] node5459;
	wire [4-1:0] node5460;
	wire [4-1:0] node5461;
	wire [4-1:0] node5466;
	wire [4-1:0] node5467;
	wire [4-1:0] node5468;
	wire [4-1:0] node5472;
	wire [4-1:0] node5475;
	wire [4-1:0] node5476;
	wire [4-1:0] node5477;
	wire [4-1:0] node5478;
	wire [4-1:0] node5481;
	wire [4-1:0] node5483;
	wire [4-1:0] node5486;
	wire [4-1:0] node5488;
	wire [4-1:0] node5491;
	wire [4-1:0] node5492;
	wire [4-1:0] node5493;
	wire [4-1:0] node5494;
	wire [4-1:0] node5498;
	wire [4-1:0] node5501;
	wire [4-1:0] node5504;
	wire [4-1:0] node5505;
	wire [4-1:0] node5506;
	wire [4-1:0] node5507;
	wire [4-1:0] node5510;
	wire [4-1:0] node5512;
	wire [4-1:0] node5515;
	wire [4-1:0] node5516;
	wire [4-1:0] node5519;
	wire [4-1:0] node5520;
	wire [4-1:0] node5524;
	wire [4-1:0] node5525;
	wire [4-1:0] node5527;
	wire [4-1:0] node5528;
	wire [4-1:0] node5532;
	wire [4-1:0] node5533;
	wire [4-1:0] node5535;
	wire [4-1:0] node5538;
	wire [4-1:0] node5539;
	wire [4-1:0] node5542;
	wire [4-1:0] node5545;
	wire [4-1:0] node5546;
	wire [4-1:0] node5547;
	wire [4-1:0] node5548;
	wire [4-1:0] node5549;
	wire [4-1:0] node5551;
	wire [4-1:0] node5554;
	wire [4-1:0] node5555;
	wire [4-1:0] node5558;
	wire [4-1:0] node5561;
	wire [4-1:0] node5562;
	wire [4-1:0] node5564;
	wire [4-1:0] node5565;
	wire [4-1:0] node5567;
	wire [4-1:0] node5570;
	wire [4-1:0] node5571;
	wire [4-1:0] node5575;
	wire [4-1:0] node5577;
	wire [4-1:0] node5580;
	wire [4-1:0] node5581;
	wire [4-1:0] node5582;
	wire [4-1:0] node5584;
	wire [4-1:0] node5586;
	wire [4-1:0] node5589;
	wire [4-1:0] node5590;
	wire [4-1:0] node5591;
	wire [4-1:0] node5595;
	wire [4-1:0] node5598;
	wire [4-1:0] node5599;
	wire [4-1:0] node5601;
	wire [4-1:0] node5603;
	wire [4-1:0] node5606;
	wire [4-1:0] node5607;
	wire [4-1:0] node5609;
	wire [4-1:0] node5613;
	wire [4-1:0] node5614;
	wire [4-1:0] node5615;
	wire [4-1:0] node5616;
	wire [4-1:0] node5618;
	wire [4-1:0] node5619;
	wire [4-1:0] node5620;
	wire [4-1:0] node5625;
	wire [4-1:0] node5626;
	wire [4-1:0] node5630;
	wire [4-1:0] node5631;
	wire [4-1:0] node5632;
	wire [4-1:0] node5635;
	wire [4-1:0] node5637;
	wire [4-1:0] node5640;
	wire [4-1:0] node5641;
	wire [4-1:0] node5642;
	wire [4-1:0] node5645;
	wire [4-1:0] node5647;
	wire [4-1:0] node5650;
	wire [4-1:0] node5653;
	wire [4-1:0] node5654;
	wire [4-1:0] node5655;
	wire [4-1:0] node5656;
	wire [4-1:0] node5657;
	wire [4-1:0] node5660;
	wire [4-1:0] node5661;
	wire [4-1:0] node5665;
	wire [4-1:0] node5666;
	wire [4-1:0] node5670;
	wire [4-1:0] node5671;
	wire [4-1:0] node5673;
	wire [4-1:0] node5676;
	wire [4-1:0] node5677;
	wire [4-1:0] node5681;
	wire [4-1:0] node5682;
	wire [4-1:0] node5684;
	wire [4-1:0] node5685;
	wire [4-1:0] node5688;
	wire [4-1:0] node5691;
	wire [4-1:0] node5692;
	wire [4-1:0] node5695;
	wire [4-1:0] node5696;
	wire [4-1:0] node5700;
	wire [4-1:0] node5701;
	wire [4-1:0] node5702;
	wire [4-1:0] node5703;
	wire [4-1:0] node5704;
	wire [4-1:0] node5705;
	wire [4-1:0] node5707;
	wire [4-1:0] node5708;
	wire [4-1:0] node5712;
	wire [4-1:0] node5714;
	wire [4-1:0] node5717;
	wire [4-1:0] node5718;
	wire [4-1:0] node5719;
	wire [4-1:0] node5722;
	wire [4-1:0] node5725;
	wire [4-1:0] node5728;
	wire [4-1:0] node5729;
	wire [4-1:0] node5730;
	wire [4-1:0] node5731;
	wire [4-1:0] node5734;
	wire [4-1:0] node5735;
	wire [4-1:0] node5739;
	wire [4-1:0] node5740;
	wire [4-1:0] node5741;
	wire [4-1:0] node5745;
	wire [4-1:0] node5746;
	wire [4-1:0] node5747;
	wire [4-1:0] node5750;
	wire [4-1:0] node5753;
	wire [4-1:0] node5755;
	wire [4-1:0] node5758;
	wire [4-1:0] node5759;
	wire [4-1:0] node5760;
	wire [4-1:0] node5763;
	wire [4-1:0] node5764;
	wire [4-1:0] node5767;
	wire [4-1:0] node5770;
	wire [4-1:0] node5771;
	wire [4-1:0] node5773;
	wire [4-1:0] node5776;
	wire [4-1:0] node5778;
	wire [4-1:0] node5781;
	wire [4-1:0] node5782;
	wire [4-1:0] node5783;
	wire [4-1:0] node5784;
	wire [4-1:0] node5785;
	wire [4-1:0] node5789;
	wire [4-1:0] node5791;
	wire [4-1:0] node5792;
	wire [4-1:0] node5796;
	wire [4-1:0] node5798;
	wire [4-1:0] node5799;
	wire [4-1:0] node5800;
	wire [4-1:0] node5804;
	wire [4-1:0] node5807;
	wire [4-1:0] node5808;
	wire [4-1:0] node5809;
	wire [4-1:0] node5810;
	wire [4-1:0] node5813;
	wire [4-1:0] node5814;
	wire [4-1:0] node5817;
	wire [4-1:0] node5820;
	wire [4-1:0] node5822;
	wire [4-1:0] node5825;
	wire [4-1:0] node5826;
	wire [4-1:0] node5827;
	wire [4-1:0] node5829;
	wire [4-1:0] node5832;
	wire [4-1:0] node5835;
	wire [4-1:0] node5836;
	wire [4-1:0] node5837;
	wire [4-1:0] node5838;
	wire [4-1:0] node5841;
	wire [4-1:0] node5845;
	wire [4-1:0] node5848;
	wire [4-1:0] node5849;
	wire [4-1:0] node5850;
	wire [4-1:0] node5851;
	wire [4-1:0] node5852;
	wire [4-1:0] node5855;
	wire [4-1:0] node5856;
	wire [4-1:0] node5857;
	wire [4-1:0] node5862;
	wire [4-1:0] node5863;
	wire [4-1:0] node5865;
	wire [4-1:0] node5867;
	wire [4-1:0] node5870;
	wire [4-1:0] node5871;
	wire [4-1:0] node5873;
	wire [4-1:0] node5876;
	wire [4-1:0] node5879;
	wire [4-1:0] node5880;
	wire [4-1:0] node5881;
	wire [4-1:0] node5882;
	wire [4-1:0] node5886;
	wire [4-1:0] node5887;
	wire [4-1:0] node5889;
	wire [4-1:0] node5892;
	wire [4-1:0] node5895;
	wire [4-1:0] node5896;
	wire [4-1:0] node5898;
	wire [4-1:0] node5899;
	wire [4-1:0] node5903;
	wire [4-1:0] node5904;
	wire [4-1:0] node5907;
	wire [4-1:0] node5910;
	wire [4-1:0] node5911;
	wire [4-1:0] node5912;
	wire [4-1:0] node5914;
	wire [4-1:0] node5915;
	wire [4-1:0] node5918;
	wire [4-1:0] node5919;
	wire [4-1:0] node5920;
	wire [4-1:0] node5923;
	wire [4-1:0] node5927;
	wire [4-1:0] node5928;
	wire [4-1:0] node5930;
	wire [4-1:0] node5933;
	wire [4-1:0] node5934;
	wire [4-1:0] node5937;
	wire [4-1:0] node5940;
	wire [4-1:0] node5941;
	wire [4-1:0] node5943;
	wire [4-1:0] node5944;
	wire [4-1:0] node5948;
	wire [4-1:0] node5950;
	wire [4-1:0] node5953;
	wire [4-1:0] node5954;
	wire [4-1:0] node5955;
	wire [4-1:0] node5956;
	wire [4-1:0] node5957;
	wire [4-1:0] node5959;
	wire [4-1:0] node5960;
	wire [4-1:0] node5961;
	wire [4-1:0] node5962;
	wire [4-1:0] node5965;
	wire [4-1:0] node5969;
	wire [4-1:0] node5970;
	wire [4-1:0] node5972;
	wire [4-1:0] node5975;
	wire [4-1:0] node5978;
	wire [4-1:0] node5979;
	wire [4-1:0] node5980;
	wire [4-1:0] node5981;
	wire [4-1:0] node5982;
	wire [4-1:0] node5986;
	wire [4-1:0] node5989;
	wire [4-1:0] node5990;
	wire [4-1:0] node5992;
	wire [4-1:0] node5994;
	wire [4-1:0] node5997;
	wire [4-1:0] node5999;
	wire [4-1:0] node6001;
	wire [4-1:0] node6004;
	wire [4-1:0] node6005;
	wire [4-1:0] node6007;
	wire [4-1:0] node6010;
	wire [4-1:0] node6011;
	wire [4-1:0] node6012;
	wire [4-1:0] node6015;
	wire [4-1:0] node6019;
	wire [4-1:0] node6021;
	wire [4-1:0] node6023;
	wire [4-1:0] node6024;
	wire [4-1:0] node6025;
	wire [4-1:0] node6026;
	wire [4-1:0] node6031;
	wire [4-1:0] node6032;
	wire [4-1:0] node6034;
	wire [4-1:0] node6035;
	wire [4-1:0] node6039;
	wire [4-1:0] node6041;
	wire [4-1:0] node6044;
	wire [4-1:0] node6045;
	wire [4-1:0] node6046;
	wire [4-1:0] node6047;
	wire [4-1:0] node6048;
	wire [4-1:0] node6049;
	wire [4-1:0] node6050;
	wire [4-1:0] node6054;
	wire [4-1:0] node6055;
	wire [4-1:0] node6056;
	wire [4-1:0] node6059;
	wire [4-1:0] node6063;
	wire [4-1:0] node6064;
	wire [4-1:0] node6067;
	wire [4-1:0] node6069;
	wire [4-1:0] node6072;
	wire [4-1:0] node6073;
	wire [4-1:0] node6074;
	wire [4-1:0] node6077;
	wire [4-1:0] node6078;
	wire [4-1:0] node6082;
	wire [4-1:0] node6085;
	wire [4-1:0] node6086;
	wire [4-1:0] node6087;
	wire [4-1:0] node6089;
	wire [4-1:0] node6092;
	wire [4-1:0] node6093;
	wire [4-1:0] node6095;
	wire [4-1:0] node6098;
	wire [4-1:0] node6101;
	wire [4-1:0] node6102;
	wire [4-1:0] node6103;
	wire [4-1:0] node6106;
	wire [4-1:0] node6108;
	wire [4-1:0] node6111;
	wire [4-1:0] node6112;
	wire [4-1:0] node6116;
	wire [4-1:0] node6117;
	wire [4-1:0] node6118;
	wire [4-1:0] node6119;
	wire [4-1:0] node6121;
	wire [4-1:0] node6122;
	wire [4-1:0] node6126;
	wire [4-1:0] node6128;
	wire [4-1:0] node6131;
	wire [4-1:0] node6132;
	wire [4-1:0] node6133;
	wire [4-1:0] node6134;
	wire [4-1:0] node6137;
	wire [4-1:0] node6141;
	wire [4-1:0] node6142;
	wire [4-1:0] node6143;
	wire [4-1:0] node6147;
	wire [4-1:0] node6150;
	wire [4-1:0] node6151;
	wire [4-1:0] node6152;
	wire [4-1:0] node6153;
	wire [4-1:0] node6155;
	wire [4-1:0] node6159;
	wire [4-1:0] node6160;
	wire [4-1:0] node6161;
	wire [4-1:0] node6166;
	wire [4-1:0] node6167;
	wire [4-1:0] node6169;
	wire [4-1:0] node6170;
	wire [4-1:0] node6173;
	wire [4-1:0] node6176;
	wire [4-1:0] node6177;
	wire [4-1:0] node6178;
	wire [4-1:0] node6181;
	wire [4-1:0] node6186;
	wire [4-1:0] node6187;
	wire [4-1:0] node6188;
	wire [4-1:0] node6189;
	wire [4-1:0] node6190;
	wire [4-1:0] node6191;
	wire [4-1:0] node6192;
	wire [4-1:0] node6193;
	wire [4-1:0] node6194;
	wire [4-1:0] node6197;
	wire [4-1:0] node6199;
	wire [4-1:0] node6202;
	wire [4-1:0] node6203;
	wire [4-1:0] node6207;
	wire [4-1:0] node6208;
	wire [4-1:0] node6209;
	wire [4-1:0] node6210;
	wire [4-1:0] node6212;
	wire [4-1:0] node6215;
	wire [4-1:0] node6219;
	wire [4-1:0] node6220;
	wire [4-1:0] node6223;
	wire [4-1:0] node6226;
	wire [4-1:0] node6227;
	wire [4-1:0] node6228;
	wire [4-1:0] node6229;
	wire [4-1:0] node6232;
	wire [4-1:0] node6234;
	wire [4-1:0] node6235;
	wire [4-1:0] node6239;
	wire [4-1:0] node6240;
	wire [4-1:0] node6243;
	wire [4-1:0] node6246;
	wire [4-1:0] node6247;
	wire [4-1:0] node6249;
	wire [4-1:0] node6250;
	wire [4-1:0] node6255;
	wire [4-1:0] node6256;
	wire [4-1:0] node6257;
	wire [4-1:0] node6258;
	wire [4-1:0] node6259;
	wire [4-1:0] node6260;
	wire [4-1:0] node6262;
	wire [4-1:0] node6265;
	wire [4-1:0] node6268;
	wire [4-1:0] node6270;
	wire [4-1:0] node6271;
	wire [4-1:0] node6275;
	wire [4-1:0] node6276;
	wire [4-1:0] node6279;
	wire [4-1:0] node6282;
	wire [4-1:0] node6283;
	wire [4-1:0] node6284;
	wire [4-1:0] node6285;
	wire [4-1:0] node6286;
	wire [4-1:0] node6290;
	wire [4-1:0] node6293;
	wire [4-1:0] node6295;
	wire [4-1:0] node6298;
	wire [4-1:0] node6299;
	wire [4-1:0] node6300;
	wire [4-1:0] node6305;
	wire [4-1:0] node6306;
	wire [4-1:0] node6307;
	wire [4-1:0] node6308;
	wire [4-1:0] node6310;
	wire [4-1:0] node6312;
	wire [4-1:0] node6315;
	wire [4-1:0] node6318;
	wire [4-1:0] node6319;
	wire [4-1:0] node6320;
	wire [4-1:0] node6326;
	wire [4-1:0] node6327;
	wire [4-1:0] node6328;
	wire [4-1:0] node6329;
	wire [4-1:0] node6330;
	wire [4-1:0] node6331;
	wire [4-1:0] node6335;
	wire [4-1:0] node6338;
	wire [4-1:0] node6339;
	wire [4-1:0] node6340;
	wire [4-1:0] node6341;
	wire [4-1:0] node6346;
	wire [4-1:0] node6348;
	wire [4-1:0] node6351;
	wire [4-1:0] node6352;
	wire [4-1:0] node6353;
	wire [4-1:0] node6355;
	wire [4-1:0] node6358;
	wire [4-1:0] node6359;
	wire [4-1:0] node6360;
	wire [4-1:0] node6364;
	wire [4-1:0] node6366;
	wire [4-1:0] node6369;
	wire [4-1:0] node6370;
	wire [4-1:0] node6371;
	wire [4-1:0] node6374;
	wire [4-1:0] node6377;
	wire [4-1:0] node6378;
	wire [4-1:0] node6381;
	wire [4-1:0] node6384;
	wire [4-1:0] node6385;
	wire [4-1:0] node6386;
	wire [4-1:0] node6387;
	wire [4-1:0] node6388;
	wire [4-1:0] node6389;
	wire [4-1:0] node6391;
	wire [4-1:0] node6395;
	wire [4-1:0] node6397;
	wire [4-1:0] node6398;
	wire [4-1:0] node6402;
	wire [4-1:0] node6403;
	wire [4-1:0] node6405;
	wire [4-1:0] node6408;
	wire [4-1:0] node6411;
	wire [4-1:0] node6412;
	wire [4-1:0] node6413;
	wire [4-1:0] node6415;
	wire [4-1:0] node6416;
	wire [4-1:0] node6421;
	wire [4-1:0] node6423;
	wire [4-1:0] node6424;
	wire [4-1:0] node6428;
	wire [4-1:0] node6429;
	wire [4-1:0] node6430;
	wire [4-1:0] node6431;
	wire [4-1:0] node6433;
	wire [4-1:0] node6434;
	wire [4-1:0] node6438;
	wire [4-1:0] node6441;
	wire [4-1:0] node6442;
	wire [4-1:0] node6444;
	wire [4-1:0] node6445;
	wire [4-1:0] node6449;
	wire [4-1:0] node6453;
	wire [4-1:0] node6454;
	wire [4-1:0] node6455;
	wire [4-1:0] node6456;
	wire [4-1:0] node6457;
	wire [4-1:0] node6458;
	wire [4-1:0] node6459;
	wire [4-1:0] node6461;
	wire [4-1:0] node6464;
	wire [4-1:0] node6467;
	wire [4-1:0] node6469;
	wire [4-1:0] node6472;
	wire [4-1:0] node6473;
	wire [4-1:0] node6474;
	wire [4-1:0] node6477;
	wire [4-1:0] node6479;
	wire [4-1:0] node6482;
	wire [4-1:0] node6484;
	wire [4-1:0] node6487;
	wire [4-1:0] node6488;
	wire [4-1:0] node6489;
	wire [4-1:0] node6490;
	wire [4-1:0] node6491;
	wire [4-1:0] node6492;
	wire [4-1:0] node6495;
	wire [4-1:0] node6498;
	wire [4-1:0] node6501;
	wire [4-1:0] node6502;
	wire [4-1:0] node6503;
	wire [4-1:0] node6508;
	wire [4-1:0] node6509;
	wire [4-1:0] node6512;
	wire [4-1:0] node6513;
	wire [4-1:0] node6517;
	wire [4-1:0] node6518;
	wire [4-1:0] node6519;
	wire [4-1:0] node6521;
	wire [4-1:0] node6524;
	wire [4-1:0] node6525;
	wire [4-1:0] node6528;
	wire [4-1:0] node6531;
	wire [4-1:0] node6532;
	wire [4-1:0] node6534;
	wire [4-1:0] node6537;
	wire [4-1:0] node6539;
	wire [4-1:0] node6542;
	wire [4-1:0] node6543;
	wire [4-1:0] node6544;
	wire [4-1:0] node6545;
	wire [4-1:0] node6546;
	wire [4-1:0] node6548;
	wire [4-1:0] node6552;
	wire [4-1:0] node6553;
	wire [4-1:0] node6557;
	wire [4-1:0] node6558;
	wire [4-1:0] node6559;
	wire [4-1:0] node6560;
	wire [4-1:0] node6563;
	wire [4-1:0] node6565;
	wire [4-1:0] node6568;
	wire [4-1:0] node6570;
	wire [4-1:0] node6574;
	wire [4-1:0] node6575;
	wire [4-1:0] node6576;
	wire [4-1:0] node6577;
	wire [4-1:0] node6579;
	wire [4-1:0] node6582;
	wire [4-1:0] node6585;
	wire [4-1:0] node6586;
	wire [4-1:0] node6589;
	wire [4-1:0] node6592;
	wire [4-1:0] node6593;
	wire [4-1:0] node6594;
	wire [4-1:0] node6596;
	wire [4-1:0] node6600;
	wire [4-1:0] node6601;
	wire [4-1:0] node6605;
	wire [4-1:0] node6606;
	wire [4-1:0] node6607;
	wire [4-1:0] node6608;
	wire [4-1:0] node6609;
	wire [4-1:0] node6611;
	wire [4-1:0] node6613;
	wire [4-1:0] node6616;
	wire [4-1:0] node6617;
	wire [4-1:0] node6620;
	wire [4-1:0] node6622;
	wire [4-1:0] node6625;
	wire [4-1:0] node6626;
	wire [4-1:0] node6627;
	wire [4-1:0] node6630;
	wire [4-1:0] node6631;
	wire [4-1:0] node6634;
	wire [4-1:0] node6637;
	wire [4-1:0] node6638;
	wire [4-1:0] node6642;
	wire [4-1:0] node6643;
	wire [4-1:0] node6644;
	wire [4-1:0] node6645;
	wire [4-1:0] node6648;
	wire [4-1:0] node6651;
	wire [4-1:0] node6653;
	wire [4-1:0] node6656;
	wire [4-1:0] node6657;
	wire [4-1:0] node6659;
	wire [4-1:0] node6660;
	wire [4-1:0] node6661;
	wire [4-1:0] node6664;
	wire [4-1:0] node6668;
	wire [4-1:0] node6670;
	wire [4-1:0] node6671;
	wire [4-1:0] node6675;
	wire [4-1:0] node6676;
	wire [4-1:0] node6677;
	wire [4-1:0] node6679;
	wire [4-1:0] node6680;
	wire [4-1:0] node6683;
	wire [4-1:0] node6686;
	wire [4-1:0] node6687;
	wire [4-1:0] node6690;
	wire [4-1:0] node6691;
	wire [4-1:0] node6693;
	wire [4-1:0] node6697;
	wire [4-1:0] node6698;
	wire [4-1:0] node6699;
	wire [4-1:0] node6700;
	wire [4-1:0] node6704;
	wire [4-1:0] node6708;
	wire [4-1:0] node6709;
	wire [4-1:0] node6710;
	wire [4-1:0] node6711;
	wire [4-1:0] node6712;
	wire [4-1:0] node6713;
	wire [4-1:0] node6714;
	wire [4-1:0] node6715;
	wire [4-1:0] node6719;
	wire [4-1:0] node6720;
	wire [4-1:0] node6723;
	wire [4-1:0] node6724;
	wire [4-1:0] node6728;
	wire [4-1:0] node6729;
	wire [4-1:0] node6730;
	wire [4-1:0] node6733;
	wire [4-1:0] node6734;
	wire [4-1:0] node6737;
	wire [4-1:0] node6740;
	wire [4-1:0] node6741;
	wire [4-1:0] node6744;
	wire [4-1:0] node6747;
	wire [4-1:0] node6748;
	wire [4-1:0] node6749;
	wire [4-1:0] node6752;
	wire [4-1:0] node6753;
	wire [4-1:0] node6755;
	wire [4-1:0] node6758;
	wire [4-1:0] node6761;
	wire [4-1:0] node6762;
	wire [4-1:0] node6764;
	wire [4-1:0] node6766;
	wire [4-1:0] node6769;
	wire [4-1:0] node6770;
	wire [4-1:0] node6773;
	wire [4-1:0] node6774;
	wire [4-1:0] node6778;
	wire [4-1:0] node6779;
	wire [4-1:0] node6780;
	wire [4-1:0] node6781;
	wire [4-1:0] node6782;
	wire [4-1:0] node6783;
	wire [4-1:0] node6784;
	wire [4-1:0] node6789;
	wire [4-1:0] node6790;
	wire [4-1:0] node6794;
	wire [4-1:0] node6795;
	wire [4-1:0] node6799;
	wire [4-1:0] node6801;
	wire [4-1:0] node6802;
	wire [4-1:0] node6804;
	wire [4-1:0] node6807;
	wire [4-1:0] node6808;
	wire [4-1:0] node6811;
	wire [4-1:0] node6814;
	wire [4-1:0] node6815;
	wire [4-1:0] node6816;
	wire [4-1:0] node6817;
	wire [4-1:0] node6819;
	wire [4-1:0] node6822;
	wire [4-1:0] node6823;
	wire [4-1:0] node6827;
	wire [4-1:0] node6828;
	wire [4-1:0] node6829;
	wire [4-1:0] node6831;
	wire [4-1:0] node6834;
	wire [4-1:0] node6838;
	wire [4-1:0] node6839;
	wire [4-1:0] node6840;
	wire [4-1:0] node6842;
	wire [4-1:0] node6845;
	wire [4-1:0] node6846;
	wire [4-1:0] node6847;
	wire [4-1:0] node6852;
	wire [4-1:0] node6853;
	wire [4-1:0] node6854;
	wire [4-1:0] node6859;
	wire [4-1:0] node6860;
	wire [4-1:0] node6861;
	wire [4-1:0] node6862;
	wire [4-1:0] node6863;
	wire [4-1:0] node6864;
	wire [4-1:0] node6865;
	wire [4-1:0] node6870;
	wire [4-1:0] node6871;
	wire [4-1:0] node6872;
	wire [4-1:0] node6877;
	wire [4-1:0] node6878;
	wire [4-1:0] node6879;
	wire [4-1:0] node6882;
	wire [4-1:0] node6884;
	wire [4-1:0] node6887;
	wire [4-1:0] node6888;
	wire [4-1:0] node6890;
	wire [4-1:0] node6892;
	wire [4-1:0] node6895;
	wire [4-1:0] node6896;
	wire [4-1:0] node6900;
	wire [4-1:0] node6901;
	wire [4-1:0] node6902;
	wire [4-1:0] node6904;
	wire [4-1:0] node6905;
	wire [4-1:0] node6909;
	wire [4-1:0] node6910;
	wire [4-1:0] node6912;
	wire [4-1:0] node6913;
	wire [4-1:0] node6916;
	wire [4-1:0] node6920;
	wire [4-1:0] node6921;
	wire [4-1:0] node6922;
	wire [4-1:0] node6925;
	wire [4-1:0] node6926;
	wire [4-1:0] node6930;
	wire [4-1:0] node6931;
	wire [4-1:0] node6932;
	wire [4-1:0] node6934;
	wire [4-1:0] node6938;
	wire [4-1:0] node6939;
	wire [4-1:0] node6943;
	wire [4-1:0] node6944;
	wire [4-1:0] node6945;
	wire [4-1:0] node6947;
	wire [4-1:0] node6948;
	wire [4-1:0] node6951;
	wire [4-1:0] node6953;
	wire [4-1:0] node6954;
	wire [4-1:0] node6958;
	wire [4-1:0] node6959;
	wire [4-1:0] node6961;
	wire [4-1:0] node6964;
	wire [4-1:0] node6965;
	wire [4-1:0] node6968;
	wire [4-1:0] node6970;
	wire [4-1:0] node6973;
	wire [4-1:0] node6974;
	wire [4-1:0] node6975;
	wire [4-1:0] node6977;
	wire [4-1:0] node6980;
	wire [4-1:0] node6981;
	wire [4-1:0] node6982;
	wire [4-1:0] node6988;
	wire [4-1:0] node6989;
	wire [4-1:0] node6990;
	wire [4-1:0] node6991;
	wire [4-1:0] node6992;
	wire [4-1:0] node6993;
	wire [4-1:0] node6994;
	wire [4-1:0] node6996;
	wire [4-1:0] node6997;
	wire [4-1:0] node7002;
	wire [4-1:0] node7003;
	wire [4-1:0] node7005;
	wire [4-1:0] node7008;
	wire [4-1:0] node7011;
	wire [4-1:0] node7012;
	wire [4-1:0] node7013;
	wire [4-1:0] node7014;
	wire [4-1:0] node7018;
	wire [4-1:0] node7020;
	wire [4-1:0] node7023;
	wire [4-1:0] node7025;
	wire [4-1:0] node7028;
	wire [4-1:0] node7029;
	wire [4-1:0] node7030;
	wire [4-1:0] node7031;
	wire [4-1:0] node7033;
	wire [4-1:0] node7036;
	wire [4-1:0] node7039;
	wire [4-1:0] node7040;
	wire [4-1:0] node7042;
	wire [4-1:0] node7045;
	wire [4-1:0] node7046;
	wire [4-1:0] node7050;
	wire [4-1:0] node7051;
	wire [4-1:0] node7052;
	wire [4-1:0] node7053;
	wire [4-1:0] node7056;
	wire [4-1:0] node7057;
	wire [4-1:0] node7061;
	wire [4-1:0] node7062;
	wire [4-1:0] node7063;
	wire [4-1:0] node7067;
	wire [4-1:0] node7070;
	wire [4-1:0] node7071;
	wire [4-1:0] node7072;
	wire [4-1:0] node7073;
	wire [4-1:0] node7076;
	wire [4-1:0] node7080;
	wire [4-1:0] node7081;
	wire [4-1:0] node7085;
	wire [4-1:0] node7086;
	wire [4-1:0] node7087;
	wire [4-1:0] node7088;
	wire [4-1:0] node7089;
	wire [4-1:0] node7093;
	wire [4-1:0] node7094;
	wire [4-1:0] node7095;
	wire [4-1:0] node7097;
	wire [4-1:0] node7100;
	wire [4-1:0] node7103;
	wire [4-1:0] node7105;
	wire [4-1:0] node7106;
	wire [4-1:0] node7109;
	wire [4-1:0] node7112;
	wire [4-1:0] node7113;
	wire [4-1:0] node7114;
	wire [4-1:0] node7117;
	wire [4-1:0] node7118;
	wire [4-1:0] node7122;
	wire [4-1:0] node7124;
	wire [4-1:0] node7127;
	wire [4-1:0] node7128;
	wire [4-1:0] node7129;
	wire [4-1:0] node7130;
	wire [4-1:0] node7131;
	wire [4-1:0] node7134;
	wire [4-1:0] node7136;
	wire [4-1:0] node7140;
	wire [4-1:0] node7141;
	wire [4-1:0] node7142;
	wire [4-1:0] node7146;
	wire [4-1:0] node7147;
	wire [4-1:0] node7149;
	wire [4-1:0] node7154;
	wire [4-1:0] node7155;
	wire [4-1:0] node7156;
	wire [4-1:0] node7157;
	wire [4-1:0] node7158;
	wire [4-1:0] node7159;
	wire [4-1:0] node7160;
	wire [4-1:0] node7163;
	wire [4-1:0] node7164;
	wire [4-1:0] node7168;
	wire [4-1:0] node7170;
	wire [4-1:0] node7171;
	wire [4-1:0] node7174;
	wire [4-1:0] node7177;
	wire [4-1:0] node7179;
	wire [4-1:0] node7180;
	wire [4-1:0] node7182;
	wire [4-1:0] node7185;
	wire [4-1:0] node7186;
	wire [4-1:0] node7189;
	wire [4-1:0] node7192;
	wire [4-1:0] node7193;
	wire [4-1:0] node7194;
	wire [4-1:0] node7195;
	wire [4-1:0] node7198;
	wire [4-1:0] node7203;
	wire [4-1:0] node7204;
	wire [4-1:0] node7205;
	wire [4-1:0] node7206;
	wire [4-1:0] node7210;
	wire [4-1:0] node7211;
	wire [4-1:0] node7213;
	wire [4-1:0] node7216;
	wire [4-1:0] node7217;
	wire [4-1:0] node7219;
	wire [4-1:0] node7224;
	wire [4-1:0] node7225;
	wire [4-1:0] node7226;
	wire [4-1:0] node7227;
	wire [4-1:0] node7229;
	wire [4-1:0] node7230;
	wire [4-1:0] node7233;
	wire [4-1:0] node7235;
	wire [4-1:0] node7238;
	wire [4-1:0] node7239;
	wire [4-1:0] node7241;
	wire [4-1:0] node7242;
	wire [4-1:0] node7245;
	wire [4-1:0] node7248;
	wire [4-1:0] node7250;
	wire [4-1:0] node7255;
	wire [4-1:0] node7256;
	wire [4-1:0] node7257;
	wire [4-1:0] node7258;
	wire [4-1:0] node7260;
	wire [4-1:0] node7261;
	wire [4-1:0] node7262;
	wire [4-1:0] node7263;
	wire [4-1:0] node7265;
	wire [4-1:0] node7266;
	wire [4-1:0] node7268;
	wire [4-1:0] node7271;
	wire [4-1:0] node7273;
	wire [4-1:0] node7274;
	wire [4-1:0] node7277;
	wire [4-1:0] node7279;
	wire [4-1:0] node7282;
	wire [4-1:0] node7283;
	wire [4-1:0] node7284;
	wire [4-1:0] node7285;
	wire [4-1:0] node7287;
	wire [4-1:0] node7290;
	wire [4-1:0] node7291;
	wire [4-1:0] node7295;
	wire [4-1:0] node7296;
	wire [4-1:0] node7298;
	wire [4-1:0] node7300;
	wire [4-1:0] node7303;
	wire [4-1:0] node7304;
	wire [4-1:0] node7308;
	wire [4-1:0] node7309;
	wire [4-1:0] node7310;
	wire [4-1:0] node7311;
	wire [4-1:0] node7315;
	wire [4-1:0] node7316;
	wire [4-1:0] node7319;
	wire [4-1:0] node7322;
	wire [4-1:0] node7323;
	wire [4-1:0] node7324;
	wire [4-1:0] node7328;
	wire [4-1:0] node7329;
	wire [4-1:0] node7333;
	wire [4-1:0] node7335;
	wire [4-1:0] node7337;
	wire [4-1:0] node7338;
	wire [4-1:0] node7339;
	wire [4-1:0] node7340;
	wire [4-1:0] node7344;
	wire [4-1:0] node7345;
	wire [4-1:0] node7349;
	wire [4-1:0] node7351;
	wire [4-1:0] node7355;
	wire [4-1:0] node7356;
	wire [4-1:0] node7357;
	wire [4-1:0] node7358;
	wire [4-1:0] node7359;
	wire [4-1:0] node7360;
	wire [4-1:0] node7361;
	wire [4-1:0] node7363;
	wire [4-1:0] node7364;
	wire [4-1:0] node7368;
	wire [4-1:0] node7370;
	wire [4-1:0] node7373;
	wire [4-1:0] node7374;
	wire [4-1:0] node7375;
	wire [4-1:0] node7377;
	wire [4-1:0] node7381;
	wire [4-1:0] node7383;
	wire [4-1:0] node7386;
	wire [4-1:0] node7387;
	wire [4-1:0] node7388;
	wire [4-1:0] node7389;
	wire [4-1:0] node7393;
	wire [4-1:0] node7395;
	wire [4-1:0] node7398;
	wire [4-1:0] node7399;
	wire [4-1:0] node7402;
	wire [4-1:0] node7403;
	wire [4-1:0] node7404;
	wire [4-1:0] node7408;
	wire [4-1:0] node7410;
	wire [4-1:0] node7413;
	wire [4-1:0] node7414;
	wire [4-1:0] node7415;
	wire [4-1:0] node7416;
	wire [4-1:0] node7417;
	wire [4-1:0] node7419;
	wire [4-1:0] node7420;
	wire [4-1:0] node7424;
	wire [4-1:0] node7426;
	wire [4-1:0] node7429;
	wire [4-1:0] node7430;
	wire [4-1:0] node7431;
	wire [4-1:0] node7434;
	wire [4-1:0] node7438;
	wire [4-1:0] node7439;
	wire [4-1:0] node7441;
	wire [4-1:0] node7442;
	wire [4-1:0] node7446;
	wire [4-1:0] node7448;
	wire [4-1:0] node7451;
	wire [4-1:0] node7452;
	wire [4-1:0] node7453;
	wire [4-1:0] node7454;
	wire [4-1:0] node7455;
	wire [4-1:0] node7460;
	wire [4-1:0] node7462;
	wire [4-1:0] node7465;
	wire [4-1:0] node7466;
	wire [4-1:0] node7467;
	wire [4-1:0] node7468;
	wire [4-1:0] node7474;
	wire [4-1:0] node7475;
	wire [4-1:0] node7476;
	wire [4-1:0] node7477;
	wire [4-1:0] node7478;
	wire [4-1:0] node7479;
	wire [4-1:0] node7482;
	wire [4-1:0] node7486;
	wire [4-1:0] node7487;
	wire [4-1:0] node7488;
	wire [4-1:0] node7490;
	wire [4-1:0] node7493;
	wire [4-1:0] node7496;
	wire [4-1:0] node7497;
	wire [4-1:0] node7500;
	wire [4-1:0] node7501;
	wire [4-1:0] node7503;
	wire [4-1:0] node7507;
	wire [4-1:0] node7508;
	wire [4-1:0] node7510;
	wire [4-1:0] node7511;
	wire [4-1:0] node7512;
	wire [4-1:0] node7516;
	wire [4-1:0] node7519;
	wire [4-1:0] node7520;
	wire [4-1:0] node7521;
	wire [4-1:0] node7523;
	wire [4-1:0] node7524;
	wire [4-1:0] node7529;
	wire [4-1:0] node7530;
	wire [4-1:0] node7531;
	wire [4-1:0] node7533;
	wire [4-1:0] node7536;
	wire [4-1:0] node7538;
	wire [4-1:0] node7541;
	wire [4-1:0] node7544;
	wire [4-1:0] node7545;
	wire [4-1:0] node7546;
	wire [4-1:0] node7547;
	wire [4-1:0] node7548;
	wire [4-1:0] node7552;
	wire [4-1:0] node7553;
	wire [4-1:0] node7557;
	wire [4-1:0] node7558;
	wire [4-1:0] node7559;
	wire [4-1:0] node7561;
	wire [4-1:0] node7564;
	wire [4-1:0] node7565;
	wire [4-1:0] node7569;
	wire [4-1:0] node7570;
	wire [4-1:0] node7571;
	wire [4-1:0] node7574;
	wire [4-1:0] node7576;
	wire [4-1:0] node7580;
	wire [4-1:0] node7581;
	wire [4-1:0] node7583;
	wire [4-1:0] node7584;
	wire [4-1:0] node7588;
	wire [4-1:0] node7589;
	wire [4-1:0] node7590;
	wire [4-1:0] node7591;
	wire [4-1:0] node7593;
	wire [4-1:0] node7597;
	wire [4-1:0] node7598;
	wire [4-1:0] node7602;
	wire [4-1:0] node7603;
	wire [4-1:0] node7606;
	wire [4-1:0] node7607;
	wire [4-1:0] node7611;
	wire [4-1:0] node7613;
	wire [4-1:0] node7614;
	wire [4-1:0] node7615;
	wire [4-1:0] node7617;
	wire [4-1:0] node7618;
	wire [4-1:0] node7619;
	wire [4-1:0] node7621;
	wire [4-1:0] node7624;
	wire [4-1:0] node7625;
	wire [4-1:0] node7629;
	wire [4-1:0] node7631;
	wire [4-1:0] node7632;
	wire [4-1:0] node7634;
	wire [4-1:0] node7637;
	wire [4-1:0] node7638;
	wire [4-1:0] node7642;
	wire [4-1:0] node7643;
	wire [4-1:0] node7644;
	wire [4-1:0] node7645;
	wire [4-1:0] node7646;
	wire [4-1:0] node7650;
	wire [4-1:0] node7651;
	wire [4-1:0] node7655;
	wire [4-1:0] node7657;
	wire [4-1:0] node7658;
	wire [4-1:0] node7662;
	wire [4-1:0] node7663;
	wire [4-1:0] node7664;
	wire [4-1:0] node7666;
	wire [4-1:0] node7669;
	wire [4-1:0] node7671;
	wire [4-1:0] node7672;
	wire [4-1:0] node7676;
	wire [4-1:0] node7677;
	wire [4-1:0] node7679;
	wire [4-1:0] node7682;
	wire [4-1:0] node7683;
	wire [4-1:0] node7687;
	wire [4-1:0] node7689;
	wire [4-1:0] node7691;
	wire [4-1:0] node7693;
	wire [4-1:0] node7695;
	wire [4-1:0] node7696;
	wire [4-1:0] node7699;
	wire [4-1:0] node7702;
	wire [4-1:0] node7703;
	wire [4-1:0] node7704;
	wire [4-1:0] node7705;
	wire [4-1:0] node7706;
	wire [4-1:0] node7707;
	wire [4-1:0] node7708;
	wire [4-1:0] node7709;
	wire [4-1:0] node7711;
	wire [4-1:0] node7715;
	wire [4-1:0] node7716;
	wire [4-1:0] node7717;
	wire [4-1:0] node7718;
	wire [4-1:0] node7722;
	wire [4-1:0] node7723;
	wire [4-1:0] node7727;
	wire [4-1:0] node7729;
	wire [4-1:0] node7732;
	wire [4-1:0] node7733;
	wire [4-1:0] node7734;
	wire [4-1:0] node7735;
	wire [4-1:0] node7736;
	wire [4-1:0] node7737;
	wire [4-1:0] node7740;
	wire [4-1:0] node7744;
	wire [4-1:0] node7746;
	wire [4-1:0] node7749;
	wire [4-1:0] node7750;
	wire [4-1:0] node7751;
	wire [4-1:0] node7754;
	wire [4-1:0] node7758;
	wire [4-1:0] node7759;
	wire [4-1:0] node7762;
	wire [4-1:0] node7764;
	wire [4-1:0] node7767;
	wire [4-1:0] node7768;
	wire [4-1:0] node7769;
	wire [4-1:0] node7770;
	wire [4-1:0] node7771;
	wire [4-1:0] node7774;
	wire [4-1:0] node7775;
	wire [4-1:0] node7777;
	wire [4-1:0] node7781;
	wire [4-1:0] node7782;
	wire [4-1:0] node7785;
	wire [4-1:0] node7788;
	wire [4-1:0] node7789;
	wire [4-1:0] node7790;
	wire [4-1:0] node7791;
	wire [4-1:0] node7796;
	wire [4-1:0] node7797;
	wire [4-1:0] node7800;
	wire [4-1:0] node7801;
	wire [4-1:0] node7805;
	wire [4-1:0] node7806;
	wire [4-1:0] node7807;
	wire [4-1:0] node7809;
	wire [4-1:0] node7812;
	wire [4-1:0] node7813;
	wire [4-1:0] node7814;
	wire [4-1:0] node7817;
	wire [4-1:0] node7820;
	wire [4-1:0] node7821;
	wire [4-1:0] node7824;
	wire [4-1:0] node7827;
	wire [4-1:0] node7828;
	wire [4-1:0] node7829;
	wire [4-1:0] node7831;
	wire [4-1:0] node7835;
	wire [4-1:0] node7836;
	wire [4-1:0] node7839;
	wire [4-1:0] node7840;
	wire [4-1:0] node7843;
	wire [4-1:0] node7846;
	wire [4-1:0] node7847;
	wire [4-1:0] node7848;
	wire [4-1:0] node7849;
	wire [4-1:0] node7850;
	wire [4-1:0] node7851;
	wire [4-1:0] node7855;
	wire [4-1:0] node7856;
	wire [4-1:0] node7860;
	wire [4-1:0] node7861;
	wire [4-1:0] node7863;
	wire [4-1:0] node7865;
	wire [4-1:0] node7868;
	wire [4-1:0] node7869;
	wire [4-1:0] node7870;
	wire [4-1:0] node7873;
	wire [4-1:0] node7877;
	wire [4-1:0] node7878;
	wire [4-1:0] node7879;
	wire [4-1:0] node7880;
	wire [4-1:0] node7881;
	wire [4-1:0] node7885;
	wire [4-1:0] node7886;
	wire [4-1:0] node7890;
	wire [4-1:0] node7891;
	wire [4-1:0] node7894;
	wire [4-1:0] node7895;
	wire [4-1:0] node7898;
	wire [4-1:0] node7901;
	wire [4-1:0] node7902;
	wire [4-1:0] node7903;
	wire [4-1:0] node7905;
	wire [4-1:0] node7907;
	wire [4-1:0] node7910;
	wire [4-1:0] node7912;
	wire [4-1:0] node7914;
	wire [4-1:0] node7917;
	wire [4-1:0] node7918;
	wire [4-1:0] node7919;
	wire [4-1:0] node7923;
	wire [4-1:0] node7925;
	wire [4-1:0] node7928;
	wire [4-1:0] node7929;
	wire [4-1:0] node7930;
	wire [4-1:0] node7931;
	wire [4-1:0] node7932;
	wire [4-1:0] node7935;
	wire [4-1:0] node7938;
	wire [4-1:0] node7939;
	wire [4-1:0] node7943;
	wire [4-1:0] node7944;
	wire [4-1:0] node7945;
	wire [4-1:0] node7946;
	wire [4-1:0] node7949;
	wire [4-1:0] node7952;
	wire [4-1:0] node7954;
	wire [4-1:0] node7957;
	wire [4-1:0] node7958;
	wire [4-1:0] node7962;
	wire [4-1:0] node7963;
	wire [4-1:0] node7964;
	wire [4-1:0] node7965;
	wire [4-1:0] node7966;
	wire [4-1:0] node7969;
	wire [4-1:0] node7971;
	wire [4-1:0] node7974;
	wire [4-1:0] node7977;
	wire [4-1:0] node7978;
	wire [4-1:0] node7979;
	wire [4-1:0] node7982;
	wire [4-1:0] node7985;
	wire [4-1:0] node7988;
	wire [4-1:0] node7989;
	wire [4-1:0] node7991;
	wire [4-1:0] node7993;
	wire [4-1:0] node7996;
	wire [4-1:0] node7997;
	wire [4-1:0] node7998;
	wire [4-1:0] node8002;
	wire [4-1:0] node8004;
	wire [4-1:0] node8007;
	wire [4-1:0] node8008;
	wire [4-1:0] node8009;
	wire [4-1:0] node8010;
	wire [4-1:0] node8011;
	wire [4-1:0] node8012;
	wire [4-1:0] node8014;
	wire [4-1:0] node8015;
	wire [4-1:0] node8018;
	wire [4-1:0] node8021;
	wire [4-1:0] node8022;
	wire [4-1:0] node8023;
	wire [4-1:0] node8024;
	wire [4-1:0] node8028;
	wire [4-1:0] node8031;
	wire [4-1:0] node8032;
	wire [4-1:0] node8035;
	wire [4-1:0] node8036;
	wire [4-1:0] node8040;
	wire [4-1:0] node8041;
	wire [4-1:0] node8042;
	wire [4-1:0] node8046;
	wire [4-1:0] node8047;
	wire [4-1:0] node8049;
	wire [4-1:0] node8052;
	wire [4-1:0] node8055;
	wire [4-1:0] node8056;
	wire [4-1:0] node8057;
	wire [4-1:0] node8058;
	wire [4-1:0] node8059;
	wire [4-1:0] node8063;
	wire [4-1:0] node8066;
	wire [4-1:0] node8067;
	wire [4-1:0] node8068;
	wire [4-1:0] node8071;
	wire [4-1:0] node8074;
	wire [4-1:0] node8077;
	wire [4-1:0] node8078;
	wire [4-1:0] node8079;
	wire [4-1:0] node8081;
	wire [4-1:0] node8084;
	wire [4-1:0] node8085;
	wire [4-1:0] node8089;
	wire [4-1:0] node8091;
	wire [4-1:0] node8094;
	wire [4-1:0] node8095;
	wire [4-1:0] node8096;
	wire [4-1:0] node8097;
	wire [4-1:0] node8098;
	wire [4-1:0] node8099;
	wire [4-1:0] node8103;
	wire [4-1:0] node8107;
	wire [4-1:0] node8108;
	wire [4-1:0] node8109;
	wire [4-1:0] node8112;
	wire [4-1:0] node8113;
	wire [4-1:0] node8114;
	wire [4-1:0] node8119;
	wire [4-1:0] node8120;
	wire [4-1:0] node8123;
	wire [4-1:0] node8124;
	wire [4-1:0] node8128;
	wire [4-1:0] node8129;
	wire [4-1:0] node8130;
	wire [4-1:0] node8131;
	wire [4-1:0] node8133;
	wire [4-1:0] node8135;
	wire [4-1:0] node8138;
	wire [4-1:0] node8142;
	wire [4-1:0] node8143;
	wire [4-1:0] node8145;
	wire [4-1:0] node8148;
	wire [4-1:0] node8149;
	wire [4-1:0] node8152;
	wire [4-1:0] node8153;
	wire [4-1:0] node8154;
	wire [4-1:0] node8159;
	wire [4-1:0] node8160;
	wire [4-1:0] node8161;
	wire [4-1:0] node8162;
	wire [4-1:0] node8163;
	wire [4-1:0] node8166;
	wire [4-1:0] node8169;
	wire [4-1:0] node8170;
	wire [4-1:0] node8172;
	wire [4-1:0] node8176;
	wire [4-1:0] node8177;
	wire [4-1:0] node8178;
	wire [4-1:0] node8181;
	wire [4-1:0] node8182;
	wire [4-1:0] node8183;
	wire [4-1:0] node8188;
	wire [4-1:0] node8189;
	wire [4-1:0] node8190;
	wire [4-1:0] node8193;
	wire [4-1:0] node8196;
	wire [4-1:0] node8198;
	wire [4-1:0] node8201;
	wire [4-1:0] node8202;
	wire [4-1:0] node8203;
	wire [4-1:0] node8204;
	wire [4-1:0] node8205;
	wire [4-1:0] node8207;
	wire [4-1:0] node8210;
	wire [4-1:0] node8213;
	wire [4-1:0] node8214;
	wire [4-1:0] node8216;
	wire [4-1:0] node8217;
	wire [4-1:0] node8221;
	wire [4-1:0] node8224;
	wire [4-1:0] node8226;
	wire [4-1:0] node8227;
	wire [4-1:0] node8230;
	wire [4-1:0] node8231;
	wire [4-1:0] node8235;
	wire [4-1:0] node8236;
	wire [4-1:0] node8237;
	wire [4-1:0] node8239;
	wire [4-1:0] node8240;
	wire [4-1:0] node8242;
	wire [4-1:0] node8245;
	wire [4-1:0] node8246;
	wire [4-1:0] node8249;
	wire [4-1:0] node8253;
	wire [4-1:0] node8254;
	wire [4-1:0] node8258;
	wire [4-1:0] node8259;
	wire [4-1:0] node8260;
	wire [4-1:0] node8261;
	wire [4-1:0] node8262;
	wire [4-1:0] node8263;
	wire [4-1:0] node8264;
	wire [4-1:0] node8265;
	wire [4-1:0] node8269;
	wire [4-1:0] node8270;
	wire [4-1:0] node8271;
	wire [4-1:0] node8275;
	wire [4-1:0] node8278;
	wire [4-1:0] node8279;
	wire [4-1:0] node8280;
	wire [4-1:0] node8282;
	wire [4-1:0] node8285;
	wire [4-1:0] node8288;
	wire [4-1:0] node8289;
	wire [4-1:0] node8291;
	wire [4-1:0] node8294;
	wire [4-1:0] node8296;
	wire [4-1:0] node8299;
	wire [4-1:0] node8300;
	wire [4-1:0] node8301;
	wire [4-1:0] node8303;
	wire [4-1:0] node8306;
	wire [4-1:0] node8307;
	wire [4-1:0] node8310;
	wire [4-1:0] node8313;
	wire [4-1:0] node8314;
	wire [4-1:0] node8315;
	wire [4-1:0] node8317;
	wire [4-1:0] node8318;
	wire [4-1:0] node8321;
	wire [4-1:0] node8324;
	wire [4-1:0] node8326;
	wire [4-1:0] node8329;
	wire [4-1:0] node8331;
	wire [4-1:0] node8332;
	wire [4-1:0] node8335;
	wire [4-1:0] node8337;
	wire [4-1:0] node8340;
	wire [4-1:0] node8341;
	wire [4-1:0] node8342;
	wire [4-1:0] node8343;
	wire [4-1:0] node8345;
	wire [4-1:0] node8347;
	wire [4-1:0] node8350;
	wire [4-1:0] node8352;
	wire [4-1:0] node8355;
	wire [4-1:0] node8356;
	wire [4-1:0] node8358;
	wire [4-1:0] node8361;
	wire [4-1:0] node8362;
	wire [4-1:0] node8364;
	wire [4-1:0] node8366;
	wire [4-1:0] node8370;
	wire [4-1:0] node8371;
	wire [4-1:0] node8372;
	wire [4-1:0] node8373;
	wire [4-1:0] node8374;
	wire [4-1:0] node8378;
	wire [4-1:0] node8379;
	wire [4-1:0] node8383;
	wire [4-1:0] node8385;
	wire [4-1:0] node8386;
	wire [4-1:0] node8387;
	wire [4-1:0] node8392;
	wire [4-1:0] node8393;
	wire [4-1:0] node8394;
	wire [4-1:0] node8396;
	wire [4-1:0] node8399;
	wire [4-1:0] node8402;
	wire [4-1:0] node8403;
	wire [4-1:0] node8404;
	wire [4-1:0] node8405;
	wire [4-1:0] node8409;
	wire [4-1:0] node8413;
	wire [4-1:0] node8414;
	wire [4-1:0] node8415;
	wire [4-1:0] node8416;
	wire [4-1:0] node8417;
	wire [4-1:0] node8418;
	wire [4-1:0] node8419;
	wire [4-1:0] node8422;
	wire [4-1:0] node8425;
	wire [4-1:0] node8426;
	wire [4-1:0] node8429;
	wire [4-1:0] node8432;
	wire [4-1:0] node8433;
	wire [4-1:0] node8434;
	wire [4-1:0] node8438;
	wire [4-1:0] node8441;
	wire [4-1:0] node8442;
	wire [4-1:0] node8443;
	wire [4-1:0] node8444;
	wire [4-1:0] node8447;
	wire [4-1:0] node8450;
	wire [4-1:0] node8452;
	wire [4-1:0] node8455;
	wire [4-1:0] node8456;
	wire [4-1:0] node8459;
	wire [4-1:0] node8460;
	wire [4-1:0] node8463;
	wire [4-1:0] node8464;
	wire [4-1:0] node8468;
	wire [4-1:0] node8469;
	wire [4-1:0] node8470;
	wire [4-1:0] node8473;
	wire [4-1:0] node8474;
	wire [4-1:0] node8475;
	wire [4-1:0] node8478;
	wire [4-1:0] node8481;
	wire [4-1:0] node8484;
	wire [4-1:0] node8485;
	wire [4-1:0] node8486;
	wire [4-1:0] node8488;
	wire [4-1:0] node8491;
	wire [4-1:0] node8492;
	wire [4-1:0] node8496;
	wire [4-1:0] node8497;
	wire [4-1:0] node8500;
	wire [4-1:0] node8503;
	wire [4-1:0] node8504;
	wire [4-1:0] node8505;
	wire [4-1:0] node8506;
	wire [4-1:0] node8507;
	wire [4-1:0] node8508;
	wire [4-1:0] node8512;
	wire [4-1:0] node8515;
	wire [4-1:0] node8516;
	wire [4-1:0] node8517;
	wire [4-1:0] node8522;
	wire [4-1:0] node8523;
	wire [4-1:0] node8524;
	wire [4-1:0] node8528;
	wire [4-1:0] node8529;
	wire [4-1:0] node8531;
	wire [4-1:0] node8534;
	wire [4-1:0] node8537;
	wire [4-1:0] node8538;
	wire [4-1:0] node8539;
	wire [4-1:0] node8541;
	wire [4-1:0] node8544;
	wire [4-1:0] node8545;
	wire [4-1:0] node8546;
	wire [4-1:0] node8550;
	wire [4-1:0] node8552;
	wire [4-1:0] node8554;
	wire [4-1:0] node8557;
	wire [4-1:0] node8559;
	wire [4-1:0] node8561;
	wire [4-1:0] node8563;
	wire [4-1:0] node8566;
	wire [4-1:0] node8567;
	wire [4-1:0] node8568;
	wire [4-1:0] node8569;
	wire [4-1:0] node8570;
	wire [4-1:0] node8571;
	wire [4-1:0] node8572;
	wire [4-1:0] node8574;
	wire [4-1:0] node8577;
	wire [4-1:0] node8578;
	wire [4-1:0] node8579;
	wire [4-1:0] node8583;
	wire [4-1:0] node8586;
	wire [4-1:0] node8587;
	wire [4-1:0] node8588;
	wire [4-1:0] node8592;
	wire [4-1:0] node8594;
	wire [4-1:0] node8597;
	wire [4-1:0] node8598;
	wire [4-1:0] node8599;
	wire [4-1:0] node8601;
	wire [4-1:0] node8602;
	wire [4-1:0] node8607;
	wire [4-1:0] node8608;
	wire [4-1:0] node8609;
	wire [4-1:0] node8611;
	wire [4-1:0] node8615;
	wire [4-1:0] node8616;
	wire [4-1:0] node8619;
	wire [4-1:0] node8620;
	wire [4-1:0] node8624;
	wire [4-1:0] node8625;
	wire [4-1:0] node8626;
	wire [4-1:0] node8627;
	wire [4-1:0] node8631;
	wire [4-1:0] node8632;
	wire [4-1:0] node8634;
	wire [4-1:0] node8635;
	wire [4-1:0] node8640;
	wire [4-1:0] node8641;
	wire [4-1:0] node8642;
	wire [4-1:0] node8645;
	wire [4-1:0] node8646;
	wire [4-1:0] node8650;
	wire [4-1:0] node8653;
	wire [4-1:0] node8654;
	wire [4-1:0] node8655;
	wire [4-1:0] node8656;
	wire [4-1:0] node8658;
	wire [4-1:0] node8661;
	wire [4-1:0] node8662;
	wire [4-1:0] node8663;
	wire [4-1:0] node8668;
	wire [4-1:0] node8669;
	wire [4-1:0] node8670;
	wire [4-1:0] node8671;
	wire [4-1:0] node8674;
	wire [4-1:0] node8678;
	wire [4-1:0] node8679;
	wire [4-1:0] node8681;
	wire [4-1:0] node8684;
	wire [4-1:0] node8685;
	wire [4-1:0] node8689;
	wire [4-1:0] node8690;
	wire [4-1:0] node8691;
	wire [4-1:0] node8692;
	wire [4-1:0] node8695;
	wire [4-1:0] node8697;
	wire [4-1:0] node8700;
	wire [4-1:0] node8701;
	wire [4-1:0] node8703;
	wire [4-1:0] node8706;
	wire [4-1:0] node8709;
	wire [4-1:0] node8711;
	wire [4-1:0] node8713;
	wire [4-1:0] node8716;
	wire [4-1:0] node8717;
	wire [4-1:0] node8718;
	wire [4-1:0] node8719;
	wire [4-1:0] node8720;
	wire [4-1:0] node8722;
	wire [4-1:0] node8723;
	wire [4-1:0] node8727;
	wire [4-1:0] node8728;
	wire [4-1:0] node8730;
	wire [4-1:0] node8733;
	wire [4-1:0] node8734;
	wire [4-1:0] node8737;
	wire [4-1:0] node8738;
	wire [4-1:0] node8742;
	wire [4-1:0] node8743;
	wire [4-1:0] node8744;
	wire [4-1:0] node8746;
	wire [4-1:0] node8747;
	wire [4-1:0] node8751;
	wire [4-1:0] node8752;
	wire [4-1:0] node8755;
	wire [4-1:0] node8758;
	wire [4-1:0] node8759;
	wire [4-1:0] node8760;
	wire [4-1:0] node8764;
	wire [4-1:0] node8765;
	wire [4-1:0] node8769;
	wire [4-1:0] node8770;
	wire [4-1:0] node8771;
	wire [4-1:0] node8772;
	wire [4-1:0] node8776;
	wire [4-1:0] node8777;
	wire [4-1:0] node8780;
	wire [4-1:0] node8781;
	wire [4-1:0] node8785;
	wire [4-1:0] node8786;
	wire [4-1:0] node8787;
	wire [4-1:0] node8789;
	wire [4-1:0] node8791;
	wire [4-1:0] node8794;
	wire [4-1:0] node8796;
	wire [4-1:0] node8798;
	wire [4-1:0] node8802;
	wire [4-1:0] node8803;
	wire [4-1:0] node8804;
	wire [4-1:0] node8805;
	wire [4-1:0] node8807;
	wire [4-1:0] node8809;
	wire [4-1:0] node8812;
	wire [4-1:0] node8813;
	wire [4-1:0] node8815;
	wire [4-1:0] node8819;
	wire [4-1:0] node8820;
	wire [4-1:0] node8821;
	wire [4-1:0] node8823;
	wire [4-1:0] node8826;
	wire [4-1:0] node8828;
	wire [4-1:0] node8832;
	wire [4-1:0] node8833;
	wire [4-1:0] node8834;
	wire [4-1:0] node8835;
	wire [4-1:0] node8836;
	wire [4-1:0] node8839;
	wire [4-1:0] node8842;
	wire [4-1:0] node8843;
	wire [4-1:0] node8846;
	wire [4-1:0] node8851;
	wire [4-1:0] node8853;
	wire [4-1:0] node8854;
	wire [4-1:0] node8856;
	wire [4-1:0] node8857;
	wire [4-1:0] node8858;
	wire [4-1:0] node8859;
	wire [4-1:0] node8861;
	wire [4-1:0] node8862;
	wire [4-1:0] node8863;
	wire [4-1:0] node8867;
	wire [4-1:0] node8868;
	wire [4-1:0] node8870;
	wire [4-1:0] node8871;
	wire [4-1:0] node8876;
	wire [4-1:0] node8877;
	wire [4-1:0] node8878;
	wire [4-1:0] node8879;
	wire [4-1:0] node8882;
	wire [4-1:0] node8883;
	wire [4-1:0] node8887;
	wire [4-1:0] node8888;
	wire [4-1:0] node8889;
	wire [4-1:0] node8892;
	wire [4-1:0] node8896;
	wire [4-1:0] node8897;
	wire [4-1:0] node8898;
	wire [4-1:0] node8902;
	wire [4-1:0] node8903;
	wire [4-1:0] node8906;
	wire [4-1:0] node8909;
	wire [4-1:0] node8911;
	wire [4-1:0] node8912;
	wire [4-1:0] node8914;
	wire [4-1:0] node8915;
	wire [4-1:0] node8917;
	wire [4-1:0] node8918;
	wire [4-1:0] node8921;
	wire [4-1:0] node8927;
	wire [4-1:0] node8928;
	wire [4-1:0] node8929;
	wire [4-1:0] node8930;
	wire [4-1:0] node8931;
	wire [4-1:0] node8932;
	wire [4-1:0] node8933;
	wire [4-1:0] node8934;
	wire [4-1:0] node8935;
	wire [4-1:0] node8938;
	wire [4-1:0] node8941;
	wire [4-1:0] node8943;
	wire [4-1:0] node8946;
	wire [4-1:0] node8947;
	wire [4-1:0] node8948;
	wire [4-1:0] node8952;
	wire [4-1:0] node8953;
	wire [4-1:0] node8954;
	wire [4-1:0] node8959;
	wire [4-1:0] node8960;
	wire [4-1:0] node8962;
	wire [4-1:0] node8963;
	wire [4-1:0] node8967;
	wire [4-1:0] node8968;
	wire [4-1:0] node8970;
	wire [4-1:0] node8972;
	wire [4-1:0] node8975;
	wire [4-1:0] node8978;
	wire [4-1:0] node8979;
	wire [4-1:0] node8980;
	wire [4-1:0] node8981;
	wire [4-1:0] node8983;
	wire [4-1:0] node8986;
	wire [4-1:0] node8987;
	wire [4-1:0] node8988;
	wire [4-1:0] node8992;
	wire [4-1:0] node8995;
	wire [4-1:0] node8996;
	wire [4-1:0] node8997;
	wire [4-1:0] node9000;
	wire [4-1:0] node9003;
	wire [4-1:0] node9005;
	wire [4-1:0] node9008;
	wire [4-1:0] node9009;
	wire [4-1:0] node9010;
	wire [4-1:0] node9012;
	wire [4-1:0] node9015;
	wire [4-1:0] node9017;
	wire [4-1:0] node9020;
	wire [4-1:0] node9021;
	wire [4-1:0] node9022;
	wire [4-1:0] node9027;
	wire [4-1:0] node9028;
	wire [4-1:0] node9029;
	wire [4-1:0] node9030;
	wire [4-1:0] node9031;
	wire [4-1:0] node9033;
	wire [4-1:0] node9037;
	wire [4-1:0] node9038;
	wire [4-1:0] node9040;
	wire [4-1:0] node9043;
	wire [4-1:0] node9044;
	wire [4-1:0] node9048;
	wire [4-1:0] node9049;
	wire [4-1:0] node9050;
	wire [4-1:0] node9052;
	wire [4-1:0] node9055;
	wire [4-1:0] node9057;
	wire [4-1:0] node9060;
	wire [4-1:0] node9062;
	wire [4-1:0] node9064;
	wire [4-1:0] node9067;
	wire [4-1:0] node9068;
	wire [4-1:0] node9069;
	wire [4-1:0] node9070;
	wire [4-1:0] node9075;
	wire [4-1:0] node9076;
	wire [4-1:0] node9077;
	wire [4-1:0] node9080;
	wire [4-1:0] node9081;
	wire [4-1:0] node9085;
	wire [4-1:0] node9087;
	wire [4-1:0] node9090;
	wire [4-1:0] node9091;
	wire [4-1:0] node9092;
	wire [4-1:0] node9093;
	wire [4-1:0] node9094;
	wire [4-1:0] node9096;
	wire [4-1:0] node9097;
	wire [4-1:0] node9098;
	wire [4-1:0] node9102;
	wire [4-1:0] node9103;
	wire [4-1:0] node9107;
	wire [4-1:0] node9108;
	wire [4-1:0] node9111;
	wire [4-1:0] node9113;
	wire [4-1:0] node9116;
	wire [4-1:0] node9117;
	wire [4-1:0] node9118;
	wire [4-1:0] node9121;
	wire [4-1:0] node9124;
	wire [4-1:0] node9125;
	wire [4-1:0] node9129;
	wire [4-1:0] node9130;
	wire [4-1:0] node9131;
	wire [4-1:0] node9132;
	wire [4-1:0] node9133;
	wire [4-1:0] node9136;
	wire [4-1:0] node9138;
	wire [4-1:0] node9142;
	wire [4-1:0] node9143;
	wire [4-1:0] node9145;
	wire [4-1:0] node9146;
	wire [4-1:0] node9150;
	wire [4-1:0] node9153;
	wire [4-1:0] node9154;
	wire [4-1:0] node9155;
	wire [4-1:0] node9158;
	wire [4-1:0] node9160;
	wire [4-1:0] node9163;
	wire [4-1:0] node9164;
	wire [4-1:0] node9168;
	wire [4-1:0] node9169;
	wire [4-1:0] node9170;
	wire [4-1:0] node9171;
	wire [4-1:0] node9172;
	wire [4-1:0] node9173;
	wire [4-1:0] node9175;
	wire [4-1:0] node9180;
	wire [4-1:0] node9181;
	wire [4-1:0] node9182;
	wire [4-1:0] node9187;
	wire [4-1:0] node9188;
	wire [4-1:0] node9189;
	wire [4-1:0] node9191;
	wire [4-1:0] node9194;
	wire [4-1:0] node9195;
	wire [4-1:0] node9198;
	wire [4-1:0] node9201;
	wire [4-1:0] node9202;
	wire [4-1:0] node9203;
	wire [4-1:0] node9208;
	wire [4-1:0] node9209;
	wire [4-1:0] node9210;
	wire [4-1:0] node9211;
	wire [4-1:0] node9213;
	wire [4-1:0] node9214;
	wire [4-1:0] node9219;
	wire [4-1:0] node9220;
	wire [4-1:0] node9224;
	wire [4-1:0] node9225;
	wire [4-1:0] node9226;
	wire [4-1:0] node9227;
	wire [4-1:0] node9228;
	wire [4-1:0] node9231;
	wire [4-1:0] node9237;
	wire [4-1:0] node9239;
	wire [4-1:0] node9240;
	wire [4-1:0] node9241;
	wire [4-1:0] node9243;
	wire [4-1:0] node9244;
	wire [4-1:0] node9245;
	wire [4-1:0] node9248;
	wire [4-1:0] node9251;
	wire [4-1:0] node9253;
	wire [4-1:0] node9257;
	wire [4-1:0] node9258;
	wire [4-1:0] node9259;
	wire [4-1:0] node9260;
	wire [4-1:0] node9261;
	wire [4-1:0] node9264;
	wire [4-1:0] node9265;
	wire [4-1:0] node9269;
	wire [4-1:0] node9270;
	wire [4-1:0] node9273;
	wire [4-1:0] node9274;
	wire [4-1:0] node9279;
	wire [4-1:0] node9280;
	wire [4-1:0] node9281;
	wire [4-1:0] node9282;
	wire [4-1:0] node9285;
	wire [4-1:0] node9286;
	wire [4-1:0] node9287;
	wire [4-1:0] node9292;
	wire [4-1:0] node9293;
	wire [4-1:0] node9295;
	wire [4-1:0] node9299;
	wire [4-1:0] node9300;
	wire [4-1:0] node9301;
	wire [4-1:0] node9306;
	wire [4-1:0] node9307;
	wire [4-1:0] node9308;
	wire [4-1:0] node9309;
	wire [4-1:0] node9310;
	wire [4-1:0] node9311;
	wire [4-1:0] node9312;
	wire [4-1:0] node9313;
	wire [4-1:0] node9314;
	wire [4-1:0] node9315;
	wire [4-1:0] node9316;
	wire [4-1:0] node9317;
	wire [4-1:0] node9319;
	wire [4-1:0] node9320;
	wire [4-1:0] node9324;
	wire [4-1:0] node9327;
	wire [4-1:0] node9328;
	wire [4-1:0] node9329;
	wire [4-1:0] node9331;
	wire [4-1:0] node9334;
	wire [4-1:0] node9335;
	wire [4-1:0] node9339;
	wire [4-1:0] node9341;
	wire [4-1:0] node9344;
	wire [4-1:0] node9345;
	wire [4-1:0] node9346;
	wire [4-1:0] node9348;
	wire [4-1:0] node9349;
	wire [4-1:0] node9352;
	wire [4-1:0] node9353;
	wire [4-1:0] node9358;
	wire [4-1:0] node9359;
	wire [4-1:0] node9360;
	wire [4-1:0] node9361;
	wire [4-1:0] node9364;
	wire [4-1:0] node9368;
	wire [4-1:0] node9369;
	wire [4-1:0] node9370;
	wire [4-1:0] node9372;
	wire [4-1:0] node9376;
	wire [4-1:0] node9377;
	wire [4-1:0] node9380;
	wire [4-1:0] node9383;
	wire [4-1:0] node9385;
	wire [4-1:0] node9386;
	wire [4-1:0] node9388;
	wire [4-1:0] node9389;
	wire [4-1:0] node9392;
	wire [4-1:0] node9394;
	wire [4-1:0] node9395;
	wire [4-1:0] node9399;
	wire [4-1:0] node9400;
	wire [4-1:0] node9401;
	wire [4-1:0] node9404;
	wire [4-1:0] node9405;
	wire [4-1:0] node9409;
	wire [4-1:0] node9411;
	wire [4-1:0] node9412;
	wire [4-1:0] node9415;
	wire [4-1:0] node9418;
	wire [4-1:0] node9419;
	wire [4-1:0] node9420;
	wire [4-1:0] node9421;
	wire [4-1:0] node9422;
	wire [4-1:0] node9423;
	wire [4-1:0] node9425;
	wire [4-1:0] node9429;
	wire [4-1:0] node9431;
	wire [4-1:0] node9434;
	wire [4-1:0] node9435;
	wire [4-1:0] node9437;
	wire [4-1:0] node9440;
	wire [4-1:0] node9441;
	wire [4-1:0] node9442;
	wire [4-1:0] node9446;
	wire [4-1:0] node9447;
	wire [4-1:0] node9451;
	wire [4-1:0] node9452;
	wire [4-1:0] node9453;
	wire [4-1:0] node9454;
	wire [4-1:0] node9457;
	wire [4-1:0] node9458;
	wire [4-1:0] node9462;
	wire [4-1:0] node9463;
	wire [4-1:0] node9466;
	wire [4-1:0] node9467;
	wire [4-1:0] node9471;
	wire [4-1:0] node9472;
	wire [4-1:0] node9473;
	wire [4-1:0] node9475;
	wire [4-1:0] node9479;
	wire [4-1:0] node9480;
	wire [4-1:0] node9481;
	wire [4-1:0] node9485;
	wire [4-1:0] node9488;
	wire [4-1:0] node9489;
	wire [4-1:0] node9490;
	wire [4-1:0] node9491;
	wire [4-1:0] node9492;
	wire [4-1:0] node9494;
	wire [4-1:0] node9495;
	wire [4-1:0] node9499;
	wire [4-1:0] node9501;
	wire [4-1:0] node9505;
	wire [4-1:0] node9506;
	wire [4-1:0] node9508;
	wire [4-1:0] node9511;
	wire [4-1:0] node9514;
	wire [4-1:0] node9515;
	wire [4-1:0] node9516;
	wire [4-1:0] node9517;
	wire [4-1:0] node9519;
	wire [4-1:0] node9523;
	wire [4-1:0] node9524;
	wire [4-1:0] node9528;
	wire [4-1:0] node9529;
	wire [4-1:0] node9530;
	wire [4-1:0] node9531;
	wire [4-1:0] node9535;
	wire [4-1:0] node9540;
	wire [4-1:0] node9541;
	wire [4-1:0] node9542;
	wire [4-1:0] node9543;
	wire [4-1:0] node9544;
	wire [4-1:0] node9545;
	wire [4-1:0] node9546;
	wire [4-1:0] node9549;
	wire [4-1:0] node9551;
	wire [4-1:0] node9554;
	wire [4-1:0] node9556;
	wire [4-1:0] node9559;
	wire [4-1:0] node9560;
	wire [4-1:0] node9561;
	wire [4-1:0] node9563;
	wire [4-1:0] node9564;
	wire [4-1:0] node9568;
	wire [4-1:0] node9570;
	wire [4-1:0] node9573;
	wire [4-1:0] node9574;
	wire [4-1:0] node9575;
	wire [4-1:0] node9578;
	wire [4-1:0] node9581;
	wire [4-1:0] node9583;
	wire [4-1:0] node9586;
	wire [4-1:0] node9587;
	wire [4-1:0] node9588;
	wire [4-1:0] node9589;
	wire [4-1:0] node9590;
	wire [4-1:0] node9591;
	wire [4-1:0] node9596;
	wire [4-1:0] node9598;
	wire [4-1:0] node9599;
	wire [4-1:0] node9602;
	wire [4-1:0] node9604;
	wire [4-1:0] node9607;
	wire [4-1:0] node9608;
	wire [4-1:0] node9609;
	wire [4-1:0] node9610;
	wire [4-1:0] node9613;
	wire [4-1:0] node9614;
	wire [4-1:0] node9619;
	wire [4-1:0] node9621;
	wire [4-1:0] node9622;
	wire [4-1:0] node9625;
	wire [4-1:0] node9628;
	wire [4-1:0] node9629;
	wire [4-1:0] node9630;
	wire [4-1:0] node9631;
	wire [4-1:0] node9633;
	wire [4-1:0] node9637;
	wire [4-1:0] node9639;
	wire [4-1:0] node9641;
	wire [4-1:0] node9644;
	wire [4-1:0] node9645;
	wire [4-1:0] node9646;
	wire [4-1:0] node9650;
	wire [4-1:0] node9651;
	wire [4-1:0] node9653;
	wire [4-1:0] node9656;
	wire [4-1:0] node9658;
	wire [4-1:0] node9661;
	wire [4-1:0] node9662;
	wire [4-1:0] node9663;
	wire [4-1:0] node9664;
	wire [4-1:0] node9665;
	wire [4-1:0] node9669;
	wire [4-1:0] node9670;
	wire [4-1:0] node9671;
	wire [4-1:0] node9673;
	wire [4-1:0] node9678;
	wire [4-1:0] node9679;
	wire [4-1:0] node9680;
	wire [4-1:0] node9683;
	wire [4-1:0] node9684;
	wire [4-1:0] node9688;
	wire [4-1:0] node9689;
	wire [4-1:0] node9693;
	wire [4-1:0] node9694;
	wire [4-1:0] node9695;
	wire [4-1:0] node9696;
	wire [4-1:0] node9698;
	wire [4-1:0] node9700;
	wire [4-1:0] node9701;
	wire [4-1:0] node9706;
	wire [4-1:0] node9707;
	wire [4-1:0] node9708;
	wire [4-1:0] node9710;
	wire [4-1:0] node9711;
	wire [4-1:0] node9715;
	wire [4-1:0] node9718;
	wire [4-1:0] node9719;
	wire [4-1:0] node9720;
	wire [4-1:0] node9724;
	wire [4-1:0] node9727;
	wire [4-1:0] node9728;
	wire [4-1:0] node9729;
	wire [4-1:0] node9731;
	wire [4-1:0] node9733;
	wire [4-1:0] node9736;
	wire [4-1:0] node9737;
	wire [4-1:0] node9740;
	wire [4-1:0] node9743;
	wire [4-1:0] node9744;
	wire [4-1:0] node9746;
	wire [4-1:0] node9747;
	wire [4-1:0] node9751;
	wire [4-1:0] node9753;
	wire [4-1:0] node9756;
	wire [4-1:0] node9757;
	wire [4-1:0] node9758;
	wire [4-1:0] node9759;
	wire [4-1:0] node9760;
	wire [4-1:0] node9762;
	wire [4-1:0] node9763;
	wire [4-1:0] node9764;
	wire [4-1:0] node9769;
	wire [4-1:0] node9771;
	wire [4-1:0] node9774;
	wire [4-1:0] node9775;
	wire [4-1:0] node9776;
	wire [4-1:0] node9777;
	wire [4-1:0] node9780;
	wire [4-1:0] node9781;
	wire [4-1:0] node9785;
	wire [4-1:0] node9786;
	wire [4-1:0] node9790;
	wire [4-1:0] node9792;
	wire [4-1:0] node9793;
	wire [4-1:0] node9797;
	wire [4-1:0] node9798;
	wire [4-1:0] node9799;
	wire [4-1:0] node9800;
	wire [4-1:0] node9801;
	wire [4-1:0] node9803;
	wire [4-1:0] node9807;
	wire [4-1:0] node9808;
	wire [4-1:0] node9809;
	wire [4-1:0] node9813;
	wire [4-1:0] node9817;
	wire [4-1:0] node9818;
	wire [4-1:0] node9819;
	wire [4-1:0] node9821;
	wire [4-1:0] node9822;
	wire [4-1:0] node9826;
	wire [4-1:0] node9828;
	wire [4-1:0] node9831;
	wire [4-1:0] node9832;
	wire [4-1:0] node9834;
	wire [4-1:0] node9837;
	wire [4-1:0] node9838;
	wire [4-1:0] node9839;
	wire [4-1:0] node9843;
	wire [4-1:0] node9845;
	wire [4-1:0] node9848;
	wire [4-1:0] node9849;
	wire [4-1:0] node9850;
	wire [4-1:0] node9851;
	wire [4-1:0] node9853;
	wire [4-1:0] node9854;
	wire [4-1:0] node9858;
	wire [4-1:0] node9860;
	wire [4-1:0] node9863;
	wire [4-1:0] node9864;
	wire [4-1:0] node9865;
	wire [4-1:0] node9866;
	wire [4-1:0] node9867;
	wire [4-1:0] node9871;
	wire [4-1:0] node9873;
	wire [4-1:0] node9877;
	wire [4-1:0] node9878;
	wire [4-1:0] node9881;
	wire [4-1:0] node9883;
	wire [4-1:0] node9886;
	wire [4-1:0] node9887;
	wire [4-1:0] node9888;
	wire [4-1:0] node9889;
	wire [4-1:0] node9890;
	wire [4-1:0] node9891;
	wire [4-1:0] node9895;
	wire [4-1:0] node9898;
	wire [4-1:0] node9900;
	wire [4-1:0] node9903;
	wire [4-1:0] node9904;
	wire [4-1:0] node9907;
	wire [4-1:0] node9909;
	wire [4-1:0] node9912;
	wire [4-1:0] node9913;
	wire [4-1:0] node9914;
	wire [4-1:0] node9916;
	wire [4-1:0] node9917;
	wire [4-1:0] node9920;
	wire [4-1:0] node9923;
	wire [4-1:0] node9924;
	wire [4-1:0] node9928;
	wire [4-1:0] node9929;
	wire [4-1:0] node9930;
	wire [4-1:0] node9932;
	wire [4-1:0] node9936;
	wire [4-1:0] node9938;
	wire [4-1:0] node9942;
	wire [4-1:0] node9943;
	wire [4-1:0] node9944;
	wire [4-1:0] node9945;
	wire [4-1:0] node9946;
	wire [4-1:0] node9947;
	wire [4-1:0] node9948;
	wire [4-1:0] node9949;
	wire [4-1:0] node9950;
	wire [4-1:0] node9951;
	wire [4-1:0] node9955;
	wire [4-1:0] node9956;
	wire [4-1:0] node9958;
	wire [4-1:0] node9962;
	wire [4-1:0] node9963;
	wire [4-1:0] node9964;
	wire [4-1:0] node9965;
	wire [4-1:0] node9969;
	wire [4-1:0] node9970;
	wire [4-1:0] node9974;
	wire [4-1:0] node9975;
	wire [4-1:0] node9977;
	wire [4-1:0] node9980;
	wire [4-1:0] node9981;
	wire [4-1:0] node9985;
	wire [4-1:0] node9986;
	wire [4-1:0] node9987;
	wire [4-1:0] node9989;
	wire [4-1:0] node9992;
	wire [4-1:0] node9993;
	wire [4-1:0] node9997;
	wire [4-1:0] node9998;
	wire [4-1:0] node9999;
	wire [4-1:0] node10002;
	wire [4-1:0] node10005;
	wire [4-1:0] node10006;
	wire [4-1:0] node10007;
	wire [4-1:0] node10010;
	wire [4-1:0] node10014;
	wire [4-1:0] node10015;
	wire [4-1:0] node10016;
	wire [4-1:0] node10017;
	wire [4-1:0] node10018;
	wire [4-1:0] node10022;
	wire [4-1:0] node10023;
	wire [4-1:0] node10026;
	wire [4-1:0] node10028;
	wire [4-1:0] node10031;
	wire [4-1:0] node10032;
	wire [4-1:0] node10033;
	wire [4-1:0] node10034;
	wire [4-1:0] node10038;
	wire [4-1:0] node10040;
	wire [4-1:0] node10042;
	wire [4-1:0] node10045;
	wire [4-1:0] node10046;
	wire [4-1:0] node10048;
	wire [4-1:0] node10052;
	wire [4-1:0] node10053;
	wire [4-1:0] node10054;
	wire [4-1:0] node10055;
	wire [4-1:0] node10056;
	wire [4-1:0] node10060;
	wire [4-1:0] node10061;
	wire [4-1:0] node10065;
	wire [4-1:0] node10066;
	wire [4-1:0] node10068;
	wire [4-1:0] node10069;
	wire [4-1:0] node10072;
	wire [4-1:0] node10075;
	wire [4-1:0] node10076;
	wire [4-1:0] node10079;
	wire [4-1:0] node10082;
	wire [4-1:0] node10083;
	wire [4-1:0] node10085;
	wire [4-1:0] node10088;
	wire [4-1:0] node10090;
	wire [4-1:0] node10091;
	wire [4-1:0] node10095;
	wire [4-1:0] node10096;
	wire [4-1:0] node10097;
	wire [4-1:0] node10098;
	wire [4-1:0] node10099;
	wire [4-1:0] node10100;
	wire [4-1:0] node10102;
	wire [4-1:0] node10107;
	wire [4-1:0] node10108;
	wire [4-1:0] node10109;
	wire [4-1:0] node10110;
	wire [4-1:0] node10113;
	wire [4-1:0] node10116;
	wire [4-1:0] node10117;
	wire [4-1:0] node10119;
	wire [4-1:0] node10123;
	wire [4-1:0] node10124;
	wire [4-1:0] node10127;
	wire [4-1:0] node10128;
	wire [4-1:0] node10131;
	wire [4-1:0] node10133;
	wire [4-1:0] node10136;
	wire [4-1:0] node10137;
	wire [4-1:0] node10139;
	wire [4-1:0] node10141;
	wire [4-1:0] node10142;
	wire [4-1:0] node10146;
	wire [4-1:0] node10147;
	wire [4-1:0] node10148;
	wire [4-1:0] node10150;
	wire [4-1:0] node10154;
	wire [4-1:0] node10156;
	wire [4-1:0] node10157;
	wire [4-1:0] node10161;
	wire [4-1:0] node10162;
	wire [4-1:0] node10163;
	wire [4-1:0] node10164;
	wire [4-1:0] node10165;
	wire [4-1:0] node10166;
	wire [4-1:0] node10170;
	wire [4-1:0] node10171;
	wire [4-1:0] node10175;
	wire [4-1:0] node10176;
	wire [4-1:0] node10177;
	wire [4-1:0] node10178;
	wire [4-1:0] node10182;
	wire [4-1:0] node10185;
	wire [4-1:0] node10186;
	wire [4-1:0] node10190;
	wire [4-1:0] node10191;
	wire [4-1:0] node10192;
	wire [4-1:0] node10195;
	wire [4-1:0] node10196;
	wire [4-1:0] node10200;
	wire [4-1:0] node10201;
	wire [4-1:0] node10202;
	wire [4-1:0] node10205;
	wire [4-1:0] node10209;
	wire [4-1:0] node10210;
	wire [4-1:0] node10211;
	wire [4-1:0] node10212;
	wire [4-1:0] node10216;
	wire [4-1:0] node10217;
	wire [4-1:0] node10220;
	wire [4-1:0] node10222;
	wire [4-1:0] node10225;
	wire [4-1:0] node10226;
	wire [4-1:0] node10228;
	wire [4-1:0] node10229;
	wire [4-1:0] node10232;
	wire [4-1:0] node10233;
	wire [4-1:0] node10237;
	wire [4-1:0] node10238;
	wire [4-1:0] node10239;
	wire [4-1:0] node10244;
	wire [4-1:0] node10245;
	wire [4-1:0] node10246;
	wire [4-1:0] node10247;
	wire [4-1:0] node10248;
	wire [4-1:0] node10249;
	wire [4-1:0] node10251;
	wire [4-1:0] node10254;
	wire [4-1:0] node10255;
	wire [4-1:0] node10256;
	wire [4-1:0] node10259;
	wire [4-1:0] node10263;
	wire [4-1:0] node10264;
	wire [4-1:0] node10266;
	wire [4-1:0] node10269;
	wire [4-1:0] node10271;
	wire [4-1:0] node10273;
	wire [4-1:0] node10276;
	wire [4-1:0] node10277;
	wire [4-1:0] node10278;
	wire [4-1:0] node10279;
	wire [4-1:0] node10280;
	wire [4-1:0] node10283;
	wire [4-1:0] node10286;
	wire [4-1:0] node10289;
	wire [4-1:0] node10290;
	wire [4-1:0] node10291;
	wire [4-1:0] node10294;
	wire [4-1:0] node10297;
	wire [4-1:0] node10300;
	wire [4-1:0] node10301;
	wire [4-1:0] node10302;
	wire [4-1:0] node10304;
	wire [4-1:0] node10308;
	wire [4-1:0] node10309;
	wire [4-1:0] node10311;
	wire [4-1:0] node10314;
	wire [4-1:0] node10317;
	wire [4-1:0] node10318;
	wire [4-1:0] node10319;
	wire [4-1:0] node10320;
	wire [4-1:0] node10321;
	wire [4-1:0] node10322;
	wire [4-1:0] node10323;
	wire [4-1:0] node10326;
	wire [4-1:0] node10330;
	wire [4-1:0] node10333;
	wire [4-1:0] node10334;
	wire [4-1:0] node10337;
	wire [4-1:0] node10338;
	wire [4-1:0] node10339;
	wire [4-1:0] node10344;
	wire [4-1:0] node10345;
	wire [4-1:0] node10346;
	wire [4-1:0] node10349;
	wire [4-1:0] node10350;
	wire [4-1:0] node10354;
	wire [4-1:0] node10355;
	wire [4-1:0] node10356;
	wire [4-1:0] node10360;
	wire [4-1:0] node10363;
	wire [4-1:0] node10364;
	wire [4-1:0] node10365;
	wire [4-1:0] node10366;
	wire [4-1:0] node10367;
	wire [4-1:0] node10371;
	wire [4-1:0] node10373;
	wire [4-1:0] node10376;
	wire [4-1:0] node10377;
	wire [4-1:0] node10380;
	wire [4-1:0] node10383;
	wire [4-1:0] node10384;
	wire [4-1:0] node10385;
	wire [4-1:0] node10387;
	wire [4-1:0] node10391;
	wire [4-1:0] node10392;
	wire [4-1:0] node10393;
	wire [4-1:0] node10397;
	wire [4-1:0] node10399;
	wire [4-1:0] node10402;
	wire [4-1:0] node10403;
	wire [4-1:0] node10404;
	wire [4-1:0] node10405;
	wire [4-1:0] node10407;
	wire [4-1:0] node10410;
	wire [4-1:0] node10411;
	wire [4-1:0] node10412;
	wire [4-1:0] node10413;
	wire [4-1:0] node10415;
	wire [4-1:0] node10419;
	wire [4-1:0] node10422;
	wire [4-1:0] node10423;
	wire [4-1:0] node10427;
	wire [4-1:0] node10428;
	wire [4-1:0] node10429;
	wire [4-1:0] node10431;
	wire [4-1:0] node10432;
	wire [4-1:0] node10435;
	wire [4-1:0] node10438;
	wire [4-1:0] node10439;
	wire [4-1:0] node10441;
	wire [4-1:0] node10442;
	wire [4-1:0] node10445;
	wire [4-1:0] node10448;
	wire [4-1:0] node10449;
	wire [4-1:0] node10451;
	wire [4-1:0] node10455;
	wire [4-1:0] node10456;
	wire [4-1:0] node10457;
	wire [4-1:0] node10458;
	wire [4-1:0] node10463;
	wire [4-1:0] node10464;
	wire [4-1:0] node10466;
	wire [4-1:0] node10469;
	wire [4-1:0] node10470;
	wire [4-1:0] node10474;
	wire [4-1:0] node10475;
	wire [4-1:0] node10476;
	wire [4-1:0] node10477;
	wire [4-1:0] node10479;
	wire [4-1:0] node10481;
	wire [4-1:0] node10484;
	wire [4-1:0] node10485;
	wire [4-1:0] node10487;
	wire [4-1:0] node10490;
	wire [4-1:0] node10491;
	wire [4-1:0] node10494;
	wire [4-1:0] node10497;
	wire [4-1:0] node10498;
	wire [4-1:0] node10501;
	wire [4-1:0] node10502;
	wire [4-1:0] node10506;
	wire [4-1:0] node10507;
	wire [4-1:0] node10509;
	wire [4-1:0] node10511;
	wire [4-1:0] node10514;
	wire [4-1:0] node10516;
	wire [4-1:0] node10519;
	wire [4-1:0] node10520;
	wire [4-1:0] node10521;
	wire [4-1:0] node10522;
	wire [4-1:0] node10523;
	wire [4-1:0] node10524;
	wire [4-1:0] node10525;
	wire [4-1:0] node10527;
	wire [4-1:0] node10530;
	wire [4-1:0] node10532;
	wire [4-1:0] node10535;
	wire [4-1:0] node10536;
	wire [4-1:0] node10537;
	wire [4-1:0] node10541;
	wire [4-1:0] node10542;
	wire [4-1:0] node10544;
	wire [4-1:0] node10547;
	wire [4-1:0] node10551;
	wire [4-1:0] node10552;
	wire [4-1:0] node10553;
	wire [4-1:0] node10554;
	wire [4-1:0] node10555;
	wire [4-1:0] node10557;
	wire [4-1:0] node10558;
	wire [4-1:0] node10561;
	wire [4-1:0] node10564;
	wire [4-1:0] node10565;
	wire [4-1:0] node10568;
	wire [4-1:0] node10570;
	wire [4-1:0] node10573;
	wire [4-1:0] node10574;
	wire [4-1:0] node10575;
	wire [4-1:0] node10578;
	wire [4-1:0] node10579;
	wire [4-1:0] node10583;
	wire [4-1:0] node10584;
	wire [4-1:0] node10588;
	wire [4-1:0] node10589;
	wire [4-1:0] node10591;
	wire [4-1:0] node10593;
	wire [4-1:0] node10596;
	wire [4-1:0] node10598;
	wire [4-1:0] node10600;
	wire [4-1:0] node10603;
	wire [4-1:0] node10604;
	wire [4-1:0] node10605;
	wire [4-1:0] node10606;
	wire [4-1:0] node10610;
	wire [4-1:0] node10611;
	wire [4-1:0] node10614;
	wire [4-1:0] node10616;
	wire [4-1:0] node10619;
	wire [4-1:0] node10620;
	wire [4-1:0] node10621;
	wire [4-1:0] node10622;
	wire [4-1:0] node10626;
	wire [4-1:0] node10629;
	wire [4-1:0] node10631;
	wire [4-1:0] node10634;
	wire [4-1:0] node10635;
	wire [4-1:0] node10636;
	wire [4-1:0] node10637;
	wire [4-1:0] node10638;
	wire [4-1:0] node10639;
	wire [4-1:0] node10640;
	wire [4-1:0] node10643;
	wire [4-1:0] node10646;
	wire [4-1:0] node10647;
	wire [4-1:0] node10651;
	wire [4-1:0] node10653;
	wire [4-1:0] node10654;
	wire [4-1:0] node10656;
	wire [4-1:0] node10660;
	wire [4-1:0] node10661;
	wire [4-1:0] node10662;
	wire [4-1:0] node10663;
	wire [4-1:0] node10664;
	wire [4-1:0] node10667;
	wire [4-1:0] node10671;
	wire [4-1:0] node10674;
	wire [4-1:0] node10676;
	wire [4-1:0] node10679;
	wire [4-1:0] node10680;
	wire [4-1:0] node10681;
	wire [4-1:0] node10683;
	wire [4-1:0] node10684;
	wire [4-1:0] node10687;
	wire [4-1:0] node10690;
	wire [4-1:0] node10692;
	wire [4-1:0] node10694;
	wire [4-1:0] node10697;
	wire [4-1:0] node10698;
	wire [4-1:0] node10699;
	wire [4-1:0] node10700;
	wire [4-1:0] node10704;
	wire [4-1:0] node10705;
	wire [4-1:0] node10709;
	wire [4-1:0] node10710;
	wire [4-1:0] node10714;
	wire [4-1:0] node10715;
	wire [4-1:0] node10716;
	wire [4-1:0] node10717;
	wire [4-1:0] node10718;
	wire [4-1:0] node10719;
	wire [4-1:0] node10724;
	wire [4-1:0] node10726;
	wire [4-1:0] node10729;
	wire [4-1:0] node10730;
	wire [4-1:0] node10731;
	wire [4-1:0] node10734;
	wire [4-1:0] node10737;
	wire [4-1:0] node10738;
	wire [4-1:0] node10742;
	wire [4-1:0] node10743;
	wire [4-1:0] node10744;
	wire [4-1:0] node10745;
	wire [4-1:0] node10747;
	wire [4-1:0] node10751;
	wire [4-1:0] node10752;
	wire [4-1:0] node10754;
	wire [4-1:0] node10757;
	wire [4-1:0] node10758;
	wire [4-1:0] node10762;
	wire [4-1:0] node10763;
	wire [4-1:0] node10765;
	wire [4-1:0] node10766;
	wire [4-1:0] node10770;
	wire [4-1:0] node10771;
	wire [4-1:0] node10776;
	wire [4-1:0] node10777;
	wire [4-1:0] node10778;
	wire [4-1:0] node10779;
	wire [4-1:0] node10780;
	wire [4-1:0] node10781;
	wire [4-1:0] node10782;
	wire [4-1:0] node10783;
	wire [4-1:0] node10784;
	wire [4-1:0] node10785;
	wire [4-1:0] node10789;
	wire [4-1:0] node10790;
	wire [4-1:0] node10794;
	wire [4-1:0] node10795;
	wire [4-1:0] node10796;
	wire [4-1:0] node10799;
	wire [4-1:0] node10802;
	wire [4-1:0] node10805;
	wire [4-1:0] node10806;
	wire [4-1:0] node10807;
	wire [4-1:0] node10810;
	wire [4-1:0] node10813;
	wire [4-1:0] node10814;
	wire [4-1:0] node10815;
	wire [4-1:0] node10818;
	wire [4-1:0] node10820;
	wire [4-1:0] node10823;
	wire [4-1:0] node10824;
	wire [4-1:0] node10828;
	wire [4-1:0] node10829;
	wire [4-1:0] node10830;
	wire [4-1:0] node10831;
	wire [4-1:0] node10832;
	wire [4-1:0] node10833;
	wire [4-1:0] node10838;
	wire [4-1:0] node10841;
	wire [4-1:0] node10843;
	wire [4-1:0] node10845;
	wire [4-1:0] node10848;
	wire [4-1:0] node10849;
	wire [4-1:0] node10850;
	wire [4-1:0] node10855;
	wire [4-1:0] node10856;
	wire [4-1:0] node10857;
	wire [4-1:0] node10858;
	wire [4-1:0] node10859;
	wire [4-1:0] node10860;
	wire [4-1:0] node10864;
	wire [4-1:0] node10866;
	wire [4-1:0] node10869;
	wire [4-1:0] node10871;
	wire [4-1:0] node10872;
	wire [4-1:0] node10875;
	wire [4-1:0] node10878;
	wire [4-1:0] node10879;
	wire [4-1:0] node10880;
	wire [4-1:0] node10883;
	wire [4-1:0] node10886;
	wire [4-1:0] node10887;
	wire [4-1:0] node10888;
	wire [4-1:0] node10892;
	wire [4-1:0] node10893;
	wire [4-1:0] node10897;
	wire [4-1:0] node10898;
	wire [4-1:0] node10899;
	wire [4-1:0] node10900;
	wire [4-1:0] node10902;
	wire [4-1:0] node10903;
	wire [4-1:0] node10907;
	wire [4-1:0] node10910;
	wire [4-1:0] node10912;
	wire [4-1:0] node10915;
	wire [4-1:0] node10916;
	wire [4-1:0] node10917;
	wire [4-1:0] node10918;
	wire [4-1:0] node10922;
	wire [4-1:0] node10925;
	wire [4-1:0] node10926;
	wire [4-1:0] node10927;
	wire [4-1:0] node10932;
	wire [4-1:0] node10933;
	wire [4-1:0] node10934;
	wire [4-1:0] node10935;
	wire [4-1:0] node10936;
	wire [4-1:0] node10938;
	wire [4-1:0] node10939;
	wire [4-1:0] node10942;
	wire [4-1:0] node10945;
	wire [4-1:0] node10946;
	wire [4-1:0] node10948;
	wire [4-1:0] node10950;
	wire [4-1:0] node10953;
	wire [4-1:0] node10954;
	wire [4-1:0] node10958;
	wire [4-1:0] node10959;
	wire [4-1:0] node10960;
	wire [4-1:0] node10961;
	wire [4-1:0] node10962;
	wire [4-1:0] node10965;
	wire [4-1:0] node10968;
	wire [4-1:0] node10971;
	wire [4-1:0] node10972;
	wire [4-1:0] node10975;
	wire [4-1:0] node10977;
	wire [4-1:0] node10980;
	wire [4-1:0] node10982;
	wire [4-1:0] node10985;
	wire [4-1:0] node10986;
	wire [4-1:0] node10987;
	wire [4-1:0] node10988;
	wire [4-1:0] node10989;
	wire [4-1:0] node10993;
	wire [4-1:0] node10996;
	wire [4-1:0] node10997;
	wire [4-1:0] node11000;
	wire [4-1:0] node11002;
	wire [4-1:0] node11005;
	wire [4-1:0] node11006;
	wire [4-1:0] node11007;
	wire [4-1:0] node11010;
	wire [4-1:0] node11013;
	wire [4-1:0] node11014;
	wire [4-1:0] node11015;
	wire [4-1:0] node11019;
	wire [4-1:0] node11020;
	wire [4-1:0] node11024;
	wire [4-1:0] node11025;
	wire [4-1:0] node11026;
	wire [4-1:0] node11027;
	wire [4-1:0] node11028;
	wire [4-1:0] node11029;
	wire [4-1:0] node11033;
	wire [4-1:0] node11035;
	wire [4-1:0] node11038;
	wire [4-1:0] node11039;
	wire [4-1:0] node11040;
	wire [4-1:0] node11042;
	wire [4-1:0] node11046;
	wire [4-1:0] node11049;
	wire [4-1:0] node11050;
	wire [4-1:0] node11052;
	wire [4-1:0] node11055;
	wire [4-1:0] node11056;
	wire [4-1:0] node11059;
	wire [4-1:0] node11060;
	wire [4-1:0] node11064;
	wire [4-1:0] node11065;
	wire [4-1:0] node11066;
	wire [4-1:0] node11067;
	wire [4-1:0] node11068;
	wire [4-1:0] node11072;
	wire [4-1:0] node11073;
	wire [4-1:0] node11076;
	wire [4-1:0] node11079;
	wire [4-1:0] node11080;
	wire [4-1:0] node11083;
	wire [4-1:0] node11086;
	wire [4-1:0] node11087;
	wire [4-1:0] node11088;
	wire [4-1:0] node11089;
	wire [4-1:0] node11092;
	wire [4-1:0] node11094;
	wire [4-1:0] node11097;
	wire [4-1:0] node11098;
	wire [4-1:0] node11101;
	wire [4-1:0] node11105;
	wire [4-1:0] node11106;
	wire [4-1:0] node11107;
	wire [4-1:0] node11108;
	wire [4-1:0] node11109;
	wire [4-1:0] node11110;
	wire [4-1:0] node11111;
	wire [4-1:0] node11114;
	wire [4-1:0] node11115;
	wire [4-1:0] node11117;
	wire [4-1:0] node11120;
	wire [4-1:0] node11123;
	wire [4-1:0] node11124;
	wire [4-1:0] node11125;
	wire [4-1:0] node11126;
	wire [4-1:0] node11130;
	wire [4-1:0] node11133;
	wire [4-1:0] node11134;
	wire [4-1:0] node11135;
	wire [4-1:0] node11139;
	wire [4-1:0] node11140;
	wire [4-1:0] node11143;
	wire [4-1:0] node11146;
	wire [4-1:0] node11147;
	wire [4-1:0] node11148;
	wire [4-1:0] node11151;
	wire [4-1:0] node11154;
	wire [4-1:0] node11155;
	wire [4-1:0] node11156;
	wire [4-1:0] node11160;
	wire [4-1:0] node11161;
	wire [4-1:0] node11165;
	wire [4-1:0] node11166;
	wire [4-1:0] node11167;
	wire [4-1:0] node11168;
	wire [4-1:0] node11170;
	wire [4-1:0] node11173;
	wire [4-1:0] node11174;
	wire [4-1:0] node11178;
	wire [4-1:0] node11179;
	wire [4-1:0] node11181;
	wire [4-1:0] node11184;
	wire [4-1:0] node11185;
	wire [4-1:0] node11189;
	wire [4-1:0] node11190;
	wire [4-1:0] node11194;
	wire [4-1:0] node11195;
	wire [4-1:0] node11196;
	wire [4-1:0] node11197;
	wire [4-1:0] node11198;
	wire [4-1:0] node11199;
	wire [4-1:0] node11203;
	wire [4-1:0] node11204;
	wire [4-1:0] node11206;
	wire [4-1:0] node11210;
	wire [4-1:0] node11211;
	wire [4-1:0] node11212;
	wire [4-1:0] node11213;
	wire [4-1:0] node11217;
	wire [4-1:0] node11219;
	wire [4-1:0] node11223;
	wire [4-1:0] node11224;
	wire [4-1:0] node11225;
	wire [4-1:0] node11229;
	wire [4-1:0] node11230;
	wire [4-1:0] node11231;
	wire [4-1:0] node11232;
	wire [4-1:0] node11236;
	wire [4-1:0] node11238;
	wire [4-1:0] node11241;
	wire [4-1:0] node11244;
	wire [4-1:0] node11245;
	wire [4-1:0] node11246;
	wire [4-1:0] node11247;
	wire [4-1:0] node11248;
	wire [4-1:0] node11251;
	wire [4-1:0] node11255;
	wire [4-1:0] node11257;
	wire [4-1:0] node11260;
	wire [4-1:0] node11261;
	wire [4-1:0] node11263;
	wire [4-1:0] node11264;
	wire [4-1:0] node11268;
	wire [4-1:0] node11269;
	wire [4-1:0] node11270;
	wire [4-1:0] node11274;
	wire [4-1:0] node11276;
	wire [4-1:0] node11279;
	wire [4-1:0] node11280;
	wire [4-1:0] node11281;
	wire [4-1:0] node11282;
	wire [4-1:0] node11283;
	wire [4-1:0] node11284;
	wire [4-1:0] node11287;
	wire [4-1:0] node11290;
	wire [4-1:0] node11291;
	wire [4-1:0] node11295;
	wire [4-1:0] node11296;
	wire [4-1:0] node11297;
	wire [4-1:0] node11298;
	wire [4-1:0] node11302;
	wire [4-1:0] node11303;
	wire [4-1:0] node11308;
	wire [4-1:0] node11309;
	wire [4-1:0] node11310;
	wire [4-1:0] node11311;
	wire [4-1:0] node11312;
	wire [4-1:0] node11316;
	wire [4-1:0] node11318;
	wire [4-1:0] node11319;
	wire [4-1:0] node11323;
	wire [4-1:0] node11324;
	wire [4-1:0] node11326;
	wire [4-1:0] node11329;
	wire [4-1:0] node11331;
	wire [4-1:0] node11334;
	wire [4-1:0] node11335;
	wire [4-1:0] node11336;
	wire [4-1:0] node11339;
	wire [4-1:0] node11340;
	wire [4-1:0] node11344;
	wire [4-1:0] node11346;
	wire [4-1:0] node11349;
	wire [4-1:0] node11350;
	wire [4-1:0] node11351;
	wire [4-1:0] node11352;
	wire [4-1:0] node11353;
	wire [4-1:0] node11355;
	wire [4-1:0] node11358;
	wire [4-1:0] node11359;
	wire [4-1:0] node11360;
	wire [4-1:0] node11364;
	wire [4-1:0] node11365;
	wire [4-1:0] node11369;
	wire [4-1:0] node11371;
	wire [4-1:0] node11374;
	wire [4-1:0] node11375;
	wire [4-1:0] node11376;
	wire [4-1:0] node11379;
	wire [4-1:0] node11383;
	wire [4-1:0] node11384;
	wire [4-1:0] node11385;
	wire [4-1:0] node11386;
	wire [4-1:0] node11390;
	wire [4-1:0] node11392;
	wire [4-1:0] node11396;
	wire [4-1:0] node11397;
	wire [4-1:0] node11398;
	wire [4-1:0] node11399;
	wire [4-1:0] node11400;
	wire [4-1:0] node11401;
	wire [4-1:0] node11403;
	wire [4-1:0] node11404;
	wire [4-1:0] node11406;
	wire [4-1:0] node11409;
	wire [4-1:0] node11410;
	wire [4-1:0] node11413;
	wire [4-1:0] node11416;
	wire [4-1:0] node11417;
	wire [4-1:0] node11418;
	wire [4-1:0] node11419;
	wire [4-1:0] node11420;
	wire [4-1:0] node11424;
	wire [4-1:0] node11426;
	wire [4-1:0] node11430;
	wire [4-1:0] node11431;
	wire [4-1:0] node11432;
	wire [4-1:0] node11434;
	wire [4-1:0] node11437;
	wire [4-1:0] node11440;
	wire [4-1:0] node11441;
	wire [4-1:0] node11444;
	wire [4-1:0] node11445;
	wire [4-1:0] node11449;
	wire [4-1:0] node11450;
	wire [4-1:0] node11451;
	wire [4-1:0] node11453;
	wire [4-1:0] node11454;
	wire [4-1:0] node11457;
	wire [4-1:0] node11460;
	wire [4-1:0] node11462;
	wire [4-1:0] node11463;
	wire [4-1:0] node11467;
	wire [4-1:0] node11468;
	wire [4-1:0] node11469;
	wire [4-1:0] node11470;
	wire [4-1:0] node11474;
	wire [4-1:0] node11475;
	wire [4-1:0] node11479;
	wire [4-1:0] node11480;
	wire [4-1:0] node11482;
	wire [4-1:0] node11484;
	wire [4-1:0] node11487;
	wire [4-1:0] node11488;
	wire [4-1:0] node11492;
	wire [4-1:0] node11493;
	wire [4-1:0] node11494;
	wire [4-1:0] node11495;
	wire [4-1:0] node11496;
	wire [4-1:0] node11499;
	wire [4-1:0] node11500;
	wire [4-1:0] node11502;
	wire [4-1:0] node11506;
	wire [4-1:0] node11508;
	wire [4-1:0] node11509;
	wire [4-1:0] node11510;
	wire [4-1:0] node11515;
	wire [4-1:0] node11516;
	wire [4-1:0] node11517;
	wire [4-1:0] node11518;
	wire [4-1:0] node11522;
	wire [4-1:0] node11523;
	wire [4-1:0] node11524;
	wire [4-1:0] node11529;
	wire [4-1:0] node11530;
	wire [4-1:0] node11532;
	wire [4-1:0] node11535;
	wire [4-1:0] node11536;
	wire [4-1:0] node11539;
	wire [4-1:0] node11542;
	wire [4-1:0] node11543;
	wire [4-1:0] node11544;
	wire [4-1:0] node11546;
	wire [4-1:0] node11548;
	wire [4-1:0] node11549;
	wire [4-1:0] node11552;
	wire [4-1:0] node11555;
	wire [4-1:0] node11556;
	wire [4-1:0] node11557;
	wire [4-1:0] node11559;
	wire [4-1:0] node11563;
	wire [4-1:0] node11565;
	wire [4-1:0] node11568;
	wire [4-1:0] node11569;
	wire [4-1:0] node11570;
	wire [4-1:0] node11572;
	wire [4-1:0] node11575;
	wire [4-1:0] node11576;
	wire [4-1:0] node11580;
	wire [4-1:0] node11581;
	wire [4-1:0] node11584;
	wire [4-1:0] node11585;
	wire [4-1:0] node11587;
	wire [4-1:0] node11591;
	wire [4-1:0] node11592;
	wire [4-1:0] node11593;
	wire [4-1:0] node11594;
	wire [4-1:0] node11595;
	wire [4-1:0] node11596;
	wire [4-1:0] node11598;
	wire [4-1:0] node11602;
	wire [4-1:0] node11604;
	wire [4-1:0] node11606;
	wire [4-1:0] node11608;
	wire [4-1:0] node11611;
	wire [4-1:0] node11614;
	wire [4-1:0] node11615;
	wire [4-1:0] node11616;
	wire [4-1:0] node11618;
	wire [4-1:0] node11619;
	wire [4-1:0] node11623;
	wire [4-1:0] node11624;
	wire [4-1:0] node11626;
	wire [4-1:0] node11629;
	wire [4-1:0] node11630;
	wire [4-1:0] node11633;
	wire [4-1:0] node11636;
	wire [4-1:0] node11637;
	wire [4-1:0] node11638;
	wire [4-1:0] node11640;
	wire [4-1:0] node11641;
	wire [4-1:0] node11644;
	wire [4-1:0] node11647;
	wire [4-1:0] node11648;
	wire [4-1:0] node11651;
	wire [4-1:0] node11654;
	wire [4-1:0] node11655;
	wire [4-1:0] node11658;
	wire [4-1:0] node11659;
	wire [4-1:0] node11662;
	wire [4-1:0] node11665;
	wire [4-1:0] node11666;
	wire [4-1:0] node11667;
	wire [4-1:0] node11668;
	wire [4-1:0] node11669;
	wire [4-1:0] node11670;
	wire [4-1:0] node11676;
	wire [4-1:0] node11677;
	wire [4-1:0] node11678;
	wire [4-1:0] node11681;
	wire [4-1:0] node11682;
	wire [4-1:0] node11686;
	wire [4-1:0] node11687;
	wire [4-1:0] node11691;
	wire [4-1:0] node11692;
	wire [4-1:0] node11693;
	wire [4-1:0] node11694;
	wire [4-1:0] node11696;
	wire [4-1:0] node11700;
	wire [4-1:0] node11702;
	wire [4-1:0] node11703;
	wire [4-1:0] node11708;
	wire [4-1:0] node11709;
	wire [4-1:0] node11710;
	wire [4-1:0] node11711;
	wire [4-1:0] node11712;
	wire [4-1:0] node11713;
	wire [4-1:0] node11714;
	wire [4-1:0] node11716;
	wire [4-1:0] node11719;
	wire [4-1:0] node11721;
	wire [4-1:0] node11722;
	wire [4-1:0] node11726;
	wire [4-1:0] node11727;
	wire [4-1:0] node11730;
	wire [4-1:0] node11732;
	wire [4-1:0] node11735;
	wire [4-1:0] node11736;
	wire [4-1:0] node11737;
	wire [4-1:0] node11738;
	wire [4-1:0] node11739;
	wire [4-1:0] node11745;
	wire [4-1:0] node11747;
	wire [4-1:0] node11748;
	wire [4-1:0] node11750;
	wire [4-1:0] node11753;
	wire [4-1:0] node11756;
	wire [4-1:0] node11757;
	wire [4-1:0] node11758;
	wire [4-1:0] node11759;
	wire [4-1:0] node11761;
	wire [4-1:0] node11763;
	wire [4-1:0] node11766;
	wire [4-1:0] node11767;
	wire [4-1:0] node11771;
	wire [4-1:0] node11772;
	wire [4-1:0] node11774;
	wire [4-1:0] node11777;
	wire [4-1:0] node11778;
	wire [4-1:0] node11781;
	wire [4-1:0] node11784;
	wire [4-1:0] node11785;
	wire [4-1:0] node11786;
	wire [4-1:0] node11789;
	wire [4-1:0] node11790;
	wire [4-1:0] node11794;
	wire [4-1:0] node11796;
	wire [4-1:0] node11798;
	wire [4-1:0] node11800;
	wire [4-1:0] node11803;
	wire [4-1:0] node11804;
	wire [4-1:0] node11805;
	wire [4-1:0] node11807;
	wire [4-1:0] node11808;
	wire [4-1:0] node11809;
	wire [4-1:0] node11810;
	wire [4-1:0] node11815;
	wire [4-1:0] node11816;
	wire [4-1:0] node11820;
	wire [4-1:0] node11821;
	wire [4-1:0] node11822;
	wire [4-1:0] node11823;
	wire [4-1:0] node11826;
	wire [4-1:0] node11829;
	wire [4-1:0] node11830;
	wire [4-1:0] node11834;
	wire [4-1:0] node11835;
	wire [4-1:0] node11836;
	wire [4-1:0] node11840;
	wire [4-1:0] node11842;
	wire [4-1:0] node11843;
	wire [4-1:0] node11847;
	wire [4-1:0] node11848;
	wire [4-1:0] node11849;
	wire [4-1:0] node11851;
	wire [4-1:0] node11852;
	wire [4-1:0] node11856;
	wire [4-1:0] node11858;
	wire [4-1:0] node11860;
	wire [4-1:0] node11864;
	wire [4-1:0] node11865;
	wire [4-1:0] node11866;
	wire [4-1:0] node11867;
	wire [4-1:0] node11868;
	wire [4-1:0] node11869;
	wire [4-1:0] node11870;
	wire [4-1:0] node11872;
	wire [4-1:0] node11876;
	wire [4-1:0] node11877;
	wire [4-1:0] node11881;
	wire [4-1:0] node11882;
	wire [4-1:0] node11886;
	wire [4-1:0] node11887;
	wire [4-1:0] node11888;
	wire [4-1:0] node11889;
	wire [4-1:0] node11891;
	wire [4-1:0] node11894;
	wire [4-1:0] node11895;
	wire [4-1:0] node11898;
	wire [4-1:0] node11902;
	wire [4-1:0] node11903;
	wire [4-1:0] node11905;
	wire [4-1:0] node11909;
	wire [4-1:0] node11910;
	wire [4-1:0] node11911;
	wire [4-1:0] node11913;
	wire [4-1:0] node11914;
	wire [4-1:0] node11918;
	wire [4-1:0] node11919;
	wire [4-1:0] node11921;
	wire [4-1:0] node11924;
	wire [4-1:0] node11925;
	wire [4-1:0] node11928;
	wire [4-1:0] node11932;
	wire [4-1:0] node11933;
	wire [4-1:0] node11934;
	wire [4-1:0] node11935;
	wire [4-1:0] node11937;
	wire [4-1:0] node11938;
	wire [4-1:0] node11940;
	wire [4-1:0] node11944;
	wire [4-1:0] node11945;
	wire [4-1:0] node11946;
	wire [4-1:0] node11947;
	wire [4-1:0] node11950;
	wire [4-1:0] node11954;
	wire [4-1:0] node11956;
	wire [4-1:0] node11957;
	wire [4-1:0] node11960;
	wire [4-1:0] node11965;
	wire [4-1:0] node11966;
	wire [4-1:0] node11967;
	wire [4-1:0] node11968;
	wire [4-1:0] node11970;
	wire [4-1:0] node11971;
	wire [4-1:0] node11972;
	wire [4-1:0] node11973;
	wire [4-1:0] node11974;
	wire [4-1:0] node11975;
	wire [4-1:0] node11977;
	wire [4-1:0] node11979;
	wire [4-1:0] node11982;
	wire [4-1:0] node11985;
	wire [4-1:0] node11987;
	wire [4-1:0] node11988;
	wire [4-1:0] node11990;
	wire [4-1:0] node11994;
	wire [4-1:0] node11995;
	wire [4-1:0] node11996;
	wire [4-1:0] node11997;
	wire [4-1:0] node11999;
	wire [4-1:0] node12002;
	wire [4-1:0] node12004;
	wire [4-1:0] node12007;
	wire [4-1:0] node12008;
	wire [4-1:0] node12009;
	wire [4-1:0] node12010;
	wire [4-1:0] node12014;
	wire [4-1:0] node12018;
	wire [4-1:0] node12019;
	wire [4-1:0] node12021;
	wire [4-1:0] node12023;
	wire [4-1:0] node12026;
	wire [4-1:0] node12029;
	wire [4-1:0] node12031;
	wire [4-1:0] node12032;
	wire [4-1:0] node12034;
	wire [4-1:0] node12035;
	wire [4-1:0] node12036;
	wire [4-1:0] node12041;
	wire [4-1:0] node12042;
	wire [4-1:0] node12044;
	wire [4-1:0] node12047;
	wire [4-1:0] node12048;
	wire [4-1:0] node12050;
	wire [4-1:0] node12051;
	wire [4-1:0] node12054;
	wire [4-1:0] node12057;
	wire [4-1:0] node12059;
	wire [4-1:0] node12060;
	wire [4-1:0] node12065;
	wire [4-1:0] node12066;
	wire [4-1:0] node12067;
	wire [4-1:0] node12068;
	wire [4-1:0] node12069;
	wire [4-1:0] node12070;
	wire [4-1:0] node12071;
	wire [4-1:0] node12073;
	wire [4-1:0] node12074;
	wire [4-1:0] node12078;
	wire [4-1:0] node12079;
	wire [4-1:0] node12080;
	wire [4-1:0] node12085;
	wire [4-1:0] node12086;
	wire [4-1:0] node12088;
	wire [4-1:0] node12089;
	wire [4-1:0] node12092;
	wire [4-1:0] node12095;
	wire [4-1:0] node12096;
	wire [4-1:0] node12098;
	wire [4-1:0] node12099;
	wire [4-1:0] node12104;
	wire [4-1:0] node12105;
	wire [4-1:0] node12106;
	wire [4-1:0] node12107;
	wire [4-1:0] node12108;
	wire [4-1:0] node12113;
	wire [4-1:0] node12114;
	wire [4-1:0] node12117;
	wire [4-1:0] node12120;
	wire [4-1:0] node12121;
	wire [4-1:0] node12122;
	wire [4-1:0] node12125;
	wire [4-1:0] node12126;
	wire [4-1:0] node12130;
	wire [4-1:0] node12131;
	wire [4-1:0] node12133;
	wire [4-1:0] node12136;
	wire [4-1:0] node12137;
	wire [4-1:0] node12141;
	wire [4-1:0] node12142;
	wire [4-1:0] node12143;
	wire [4-1:0] node12144;
	wire [4-1:0] node12146;
	wire [4-1:0] node12149;
	wire [4-1:0] node12150;
	wire [4-1:0] node12154;
	wire [4-1:0] node12155;
	wire [4-1:0] node12156;
	wire [4-1:0] node12158;
	wire [4-1:0] node12161;
	wire [4-1:0] node12163;
	wire [4-1:0] node12166;
	wire [4-1:0] node12168;
	wire [4-1:0] node12171;
	wire [4-1:0] node12172;
	wire [4-1:0] node12174;
	wire [4-1:0] node12175;
	wire [4-1:0] node12179;
	wire [4-1:0] node12180;
	wire [4-1:0] node12181;
	wire [4-1:0] node12185;
	wire [4-1:0] node12187;
	wire [4-1:0] node12189;
	wire [4-1:0] node12190;
	wire [4-1:0] node12193;
	wire [4-1:0] node12196;
	wire [4-1:0] node12197;
	wire [4-1:0] node12198;
	wire [4-1:0] node12199;
	wire [4-1:0] node12200;
	wire [4-1:0] node12202;
	wire [4-1:0] node12203;
	wire [4-1:0] node12206;
	wire [4-1:0] node12208;
	wire [4-1:0] node12211;
	wire [4-1:0] node12212;
	wire [4-1:0] node12215;
	wire [4-1:0] node12218;
	wire [4-1:0] node12219;
	wire [4-1:0] node12220;
	wire [4-1:0] node12223;
	wire [4-1:0] node12225;
	wire [4-1:0] node12228;
	wire [4-1:0] node12229;
	wire [4-1:0] node12232;
	wire [4-1:0] node12235;
	wire [4-1:0] node12236;
	wire [4-1:0] node12237;
	wire [4-1:0] node12238;
	wire [4-1:0] node12240;
	wire [4-1:0] node12243;
	wire [4-1:0] node12244;
	wire [4-1:0] node12248;
	wire [4-1:0] node12249;
	wire [4-1:0] node12251;
	wire [4-1:0] node12252;
	wire [4-1:0] node12257;
	wire [4-1:0] node12258;
	wire [4-1:0] node12259;
	wire [4-1:0] node12263;
	wire [4-1:0] node12264;
	wire [4-1:0] node12266;
	wire [4-1:0] node12267;
	wire [4-1:0] node12270;
	wire [4-1:0] node12273;
	wire [4-1:0] node12276;
	wire [4-1:0] node12277;
	wire [4-1:0] node12278;
	wire [4-1:0] node12279;
	wire [4-1:0] node12280;
	wire [4-1:0] node12281;
	wire [4-1:0] node12285;
	wire [4-1:0] node12288;
	wire [4-1:0] node12289;
	wire [4-1:0] node12293;
	wire [4-1:0] node12294;
	wire [4-1:0] node12295;
	wire [4-1:0] node12298;
	wire [4-1:0] node12301;
	wire [4-1:0] node12303;
	wire [4-1:0] node12304;
	wire [4-1:0] node12308;
	wire [4-1:0] node12309;
	wire [4-1:0] node12310;
	wire [4-1:0] node12312;
	wire [4-1:0] node12315;
	wire [4-1:0] node12316;
	wire [4-1:0] node12320;
	wire [4-1:0] node12321;
	wire [4-1:0] node12322;
	wire [4-1:0] node12326;
	wire [4-1:0] node12327;
	wire [4-1:0] node12330;
	wire [4-1:0] node12333;
	wire [4-1:0] node12335;
	wire [4-1:0] node12336;
	wire [4-1:0] node12337;
	wire [4-1:0] node12338;
	wire [4-1:0] node12339;
	wire [4-1:0] node12340;
	wire [4-1:0] node12341;
	wire [4-1:0] node12347;
	wire [4-1:0] node12348;
	wire [4-1:0] node12349;
	wire [4-1:0] node12352;
	wire [4-1:0] node12355;
	wire [4-1:0] node12356;
	wire [4-1:0] node12359;
	wire [4-1:0] node12360;
	wire [4-1:0] node12363;
	wire [4-1:0] node12367;
	wire [4-1:0] node12368;
	wire [4-1:0] node12369;
	wire [4-1:0] node12370;
	wire [4-1:0] node12371;
	wire [4-1:0] node12373;
	wire [4-1:0] node12374;
	wire [4-1:0] node12378;
	wire [4-1:0] node12380;
	wire [4-1:0] node12383;
	wire [4-1:0] node12384;
	wire [4-1:0] node12385;
	wire [4-1:0] node12388;
	wire [4-1:0] node12392;
	wire [4-1:0] node12394;
	wire [4-1:0] node12395;
	wire [4-1:0] node12398;
	wire [4-1:0] node12401;
	wire [4-1:0] node12402;
	wire [4-1:0] node12403;
	wire [4-1:0] node12405;
	wire [4-1:0] node12408;
	wire [4-1:0] node12411;
	wire [4-1:0] node12412;
	wire [4-1:0] node12414;
	wire [4-1:0] node12417;
	wire [4-1:0] node12418;
	wire [4-1:0] node12419;
	wire [4-1:0] node12423;
	wire [4-1:0] node12425;
	wire [4-1:0] node12428;
	wire [4-1:0] node12429;
	wire [4-1:0] node12430;
	wire [4-1:0] node12431;
	wire [4-1:0] node12432;
	wire [4-1:0] node12433;
	wire [4-1:0] node12434;
	wire [4-1:0] node12435;
	wire [4-1:0] node12436;
	wire [4-1:0] node12437;
	wire [4-1:0] node12441;
	wire [4-1:0] node12443;
	wire [4-1:0] node12445;
	wire [4-1:0] node12448;
	wire [4-1:0] node12449;
	wire [4-1:0] node12451;
	wire [4-1:0] node12452;
	wire [4-1:0] node12455;
	wire [4-1:0] node12458;
	wire [4-1:0] node12461;
	wire [4-1:0] node12462;
	wire [4-1:0] node12463;
	wire [4-1:0] node12464;
	wire [4-1:0] node12467;
	wire [4-1:0] node12471;
	wire [4-1:0] node12473;
	wire [4-1:0] node12476;
	wire [4-1:0] node12477;
	wire [4-1:0] node12478;
	wire [4-1:0] node12479;
	wire [4-1:0] node12482;
	wire [4-1:0] node12484;
	wire [4-1:0] node12487;
	wire [4-1:0] node12488;
	wire [4-1:0] node12489;
	wire [4-1:0] node12492;
	wire [4-1:0] node12495;
	wire [4-1:0] node12497;
	wire [4-1:0] node12500;
	wire [4-1:0] node12501;
	wire [4-1:0] node12502;
	wire [4-1:0] node12503;
	wire [4-1:0] node12505;
	wire [4-1:0] node12509;
	wire [4-1:0] node12510;
	wire [4-1:0] node12514;
	wire [4-1:0] node12515;
	wire [4-1:0] node12518;
	wire [4-1:0] node12519;
	wire [4-1:0] node12523;
	wire [4-1:0] node12524;
	wire [4-1:0] node12525;
	wire [4-1:0] node12526;
	wire [4-1:0] node12528;
	wire [4-1:0] node12529;
	wire [4-1:0] node12530;
	wire [4-1:0] node12535;
	wire [4-1:0] node12537;
	wire [4-1:0] node12539;
	wire [4-1:0] node12542;
	wire [4-1:0] node12543;
	wire [4-1:0] node12545;
	wire [4-1:0] node12548;
	wire [4-1:0] node12550;
	wire [4-1:0] node12551;
	wire [4-1:0] node12555;
	wire [4-1:0] node12556;
	wire [4-1:0] node12557;
	wire [4-1:0] node12558;
	wire [4-1:0] node12561;
	wire [4-1:0] node12564;
	wire [4-1:0] node12565;
	wire [4-1:0] node12567;
	wire [4-1:0] node12570;
	wire [4-1:0] node12571;
	wire [4-1:0] node12575;
	wire [4-1:0] node12576;
	wire [4-1:0] node12577;
	wire [4-1:0] node12578;
	wire [4-1:0] node12579;
	wire [4-1:0] node12582;
	wire [4-1:0] node12586;
	wire [4-1:0] node12589;
	wire [4-1:0] node12590;
	wire [4-1:0] node12591;
	wire [4-1:0] node12594;
	wire [4-1:0] node12595;
	wire [4-1:0] node12598;
	wire [4-1:0] node12601;
	wire [4-1:0] node12604;
	wire [4-1:0] node12605;
	wire [4-1:0] node12606;
	wire [4-1:0] node12607;
	wire [4-1:0] node12608;
	wire [4-1:0] node12609;
	wire [4-1:0] node12610;
	wire [4-1:0] node12614;
	wire [4-1:0] node12615;
	wire [4-1:0] node12619;
	wire [4-1:0] node12621;
	wire [4-1:0] node12624;
	wire [4-1:0] node12625;
	wire [4-1:0] node12627;
	wire [4-1:0] node12629;
	wire [4-1:0] node12632;
	wire [4-1:0] node12633;
	wire [4-1:0] node12636;
	wire [4-1:0] node12639;
	wire [4-1:0] node12640;
	wire [4-1:0] node12641;
	wire [4-1:0] node12642;
	wire [4-1:0] node12643;
	wire [4-1:0] node12646;
	wire [4-1:0] node12649;
	wire [4-1:0] node12651;
	wire [4-1:0] node12652;
	wire [4-1:0] node12656;
	wire [4-1:0] node12657;
	wire [4-1:0] node12660;
	wire [4-1:0] node12663;
	wire [4-1:0] node12664;
	wire [4-1:0] node12665;
	wire [4-1:0] node12667;
	wire [4-1:0] node12668;
	wire [4-1:0] node12672;
	wire [4-1:0] node12674;
	wire [4-1:0] node12675;
	wire [4-1:0] node12679;
	wire [4-1:0] node12681;
	wire [4-1:0] node12684;
	wire [4-1:0] node12685;
	wire [4-1:0] node12686;
	wire [4-1:0] node12687;
	wire [4-1:0] node12688;
	wire [4-1:0] node12690;
	wire [4-1:0] node12694;
	wire [4-1:0] node12696;
	wire [4-1:0] node12699;
	wire [4-1:0] node12700;
	wire [4-1:0] node12701;
	wire [4-1:0] node12704;
	wire [4-1:0] node12705;
	wire [4-1:0] node12708;
	wire [4-1:0] node12711;
	wire [4-1:0] node12712;
	wire [4-1:0] node12713;
	wire [4-1:0] node12716;
	wire [4-1:0] node12717;
	wire [4-1:0] node12721;
	wire [4-1:0] node12722;
	wire [4-1:0] node12726;
	wire [4-1:0] node12727;
	wire [4-1:0] node12728;
	wire [4-1:0] node12729;
	wire [4-1:0] node12730;
	wire [4-1:0] node12733;
	wire [4-1:0] node12735;
	wire [4-1:0] node12738;
	wire [4-1:0] node12740;
	wire [4-1:0] node12741;
	wire [4-1:0] node12744;
	wire [4-1:0] node12747;
	wire [4-1:0] node12748;
	wire [4-1:0] node12749;
	wire [4-1:0] node12752;
	wire [4-1:0] node12755;
	wire [4-1:0] node12758;
	wire [4-1:0] node12759;
	wire [4-1:0] node12760;
	wire [4-1:0] node12761;
	wire [4-1:0] node12766;
	wire [4-1:0] node12767;
	wire [4-1:0] node12768;
	wire [4-1:0] node12773;
	wire [4-1:0] node12774;
	wire [4-1:0] node12775;
	wire [4-1:0] node12776;
	wire [4-1:0] node12777;
	wire [4-1:0] node12778;
	wire [4-1:0] node12779;
	wire [4-1:0] node12782;
	wire [4-1:0] node12785;
	wire [4-1:0] node12786;
	wire [4-1:0] node12789;
	wire [4-1:0] node12792;
	wire [4-1:0] node12793;
	wire [4-1:0] node12794;
	wire [4-1:0] node12795;
	wire [4-1:0] node12800;
	wire [4-1:0] node12801;
	wire [4-1:0] node12803;
	wire [4-1:0] node12806;
	wire [4-1:0] node12809;
	wire [4-1:0] node12810;
	wire [4-1:0] node12811;
	wire [4-1:0] node12813;
	wire [4-1:0] node12817;
	wire [4-1:0] node12818;
	wire [4-1:0] node12820;
	wire [4-1:0] node12823;
	wire [4-1:0] node12824;
	wire [4-1:0] node12826;
	wire [4-1:0] node12830;
	wire [4-1:0] node12831;
	wire [4-1:0] node12832;
	wire [4-1:0] node12833;
	wire [4-1:0] node12834;
	wire [4-1:0] node12838;
	wire [4-1:0] node12839;
	wire [4-1:0] node12840;
	wire [4-1:0] node12842;
	wire [4-1:0] node12846;
	wire [4-1:0] node12848;
	wire [4-1:0] node12851;
	wire [4-1:0] node12852;
	wire [4-1:0] node12853;
	wire [4-1:0] node12856;
	wire [4-1:0] node12860;
	wire [4-1:0] node12861;
	wire [4-1:0] node12862;
	wire [4-1:0] node12864;
	wire [4-1:0] node12865;
	wire [4-1:0] node12869;
	wire [4-1:0] node12870;
	wire [4-1:0] node12872;
	wire [4-1:0] node12875;
	wire [4-1:0] node12878;
	wire [4-1:0] node12879;
	wire [4-1:0] node12880;
	wire [4-1:0] node12884;
	wire [4-1:0] node12885;
	wire [4-1:0] node12888;
	wire [4-1:0] node12889;
	wire [4-1:0] node12893;
	wire [4-1:0] node12894;
	wire [4-1:0] node12895;
	wire [4-1:0] node12896;
	wire [4-1:0] node12897;
	wire [4-1:0] node12899;
	wire [4-1:0] node12902;
	wire [4-1:0] node12903;
	wire [4-1:0] node12904;
	wire [4-1:0] node12909;
	wire [4-1:0] node12910;
	wire [4-1:0] node12912;
	wire [4-1:0] node12915;
	wire [4-1:0] node12917;
	wire [4-1:0] node12920;
	wire [4-1:0] node12921;
	wire [4-1:0] node12922;
	wire [4-1:0] node12923;
	wire [4-1:0] node12925;
	wire [4-1:0] node12928;
	wire [4-1:0] node12931;
	wire [4-1:0] node12932;
	wire [4-1:0] node12933;
	wire [4-1:0] node12936;
	wire [4-1:0] node12940;
	wire [4-1:0] node12941;
	wire [4-1:0] node12942;
	wire [4-1:0] node12946;
	wire [4-1:0] node12947;
	wire [4-1:0] node12948;
	wire [4-1:0] node12952;
	wire [4-1:0] node12955;
	wire [4-1:0] node12956;
	wire [4-1:0] node12957;
	wire [4-1:0] node12958;
	wire [4-1:0] node12959;
	wire [4-1:0] node12960;
	wire [4-1:0] node12963;
	wire [4-1:0] node12966;
	wire [4-1:0] node12967;
	wire [4-1:0] node12970;
	wire [4-1:0] node12973;
	wire [4-1:0] node12975;
	wire [4-1:0] node12978;
	wire [4-1:0] node12979;
	wire [4-1:0] node12980;
	wire [4-1:0] node12981;
	wire [4-1:0] node12985;
	wire [4-1:0] node12986;
	wire [4-1:0] node12988;
	wire [4-1:0] node12992;
	wire [4-1:0] node12993;
	wire [4-1:0] node12997;
	wire [4-1:0] node12998;
	wire [4-1:0] node12999;
	wire [4-1:0] node13003;
	wire [4-1:0] node13004;
	wire [4-1:0] node13005;
	wire [4-1:0] node13009;
	wire [4-1:0] node13010;
	wire [4-1:0] node13014;
	wire [4-1:0] node13015;
	wire [4-1:0] node13016;
	wire [4-1:0] node13017;
	wire [4-1:0] node13018;
	wire [4-1:0] node13019;
	wire [4-1:0] node13020;
	wire [4-1:0] node13022;
	wire [4-1:0] node13023;
	wire [4-1:0] node13024;
	wire [4-1:0] node13028;
	wire [4-1:0] node13031;
	wire [4-1:0] node13032;
	wire [4-1:0] node13034;
	wire [4-1:0] node13037;
	wire [4-1:0] node13038;
	wire [4-1:0] node13040;
	wire [4-1:0] node13043;
	wire [4-1:0] node13046;
	wire [4-1:0] node13047;
	wire [4-1:0] node13048;
	wire [4-1:0] node13050;
	wire [4-1:0] node13053;
	wire [4-1:0] node13054;
	wire [4-1:0] node13056;
	wire [4-1:0] node13060;
	wire [4-1:0] node13061;
	wire [4-1:0] node13062;
	wire [4-1:0] node13067;
	wire [4-1:0] node13068;
	wire [4-1:0] node13069;
	wire [4-1:0] node13070;
	wire [4-1:0] node13071;
	wire [4-1:0] node13076;
	wire [4-1:0] node13078;
	wire [4-1:0] node13081;
	wire [4-1:0] node13082;
	wire [4-1:0] node13083;
	wire [4-1:0] node13084;
	wire [4-1:0] node13086;
	wire [4-1:0] node13090;
	wire [4-1:0] node13091;
	wire [4-1:0] node13096;
	wire [4-1:0] node13097;
	wire [4-1:0] node13098;
	wire [4-1:0] node13099;
	wire [4-1:0] node13100;
	wire [4-1:0] node13101;
	wire [4-1:0] node13106;
	wire [4-1:0] node13107;
	wire [4-1:0] node13111;
	wire [4-1:0] node13112;
	wire [4-1:0] node13113;
	wire [4-1:0] node13114;
	wire [4-1:0] node13115;
	wire [4-1:0] node13119;
	wire [4-1:0] node13120;
	wire [4-1:0] node13124;
	wire [4-1:0] node13126;
	wire [4-1:0] node13129;
	wire [4-1:0] node13131;
	wire [4-1:0] node13133;
	wire [4-1:0] node13136;
	wire [4-1:0] node13137;
	wire [4-1:0] node13138;
	wire [4-1:0] node13139;
	wire [4-1:0] node13140;
	wire [4-1:0] node13143;
	wire [4-1:0] node13146;
	wire [4-1:0] node13147;
	wire [4-1:0] node13151;
	wire [4-1:0] node13154;
	wire [4-1:0] node13155;
	wire [4-1:0] node13157;
	wire [4-1:0] node13160;
	wire [4-1:0] node13162;
	wire [4-1:0] node13165;
	wire [4-1:0] node13166;
	wire [4-1:0] node13167;
	wire [4-1:0] node13168;
	wire [4-1:0] node13169;
	wire [4-1:0] node13170;
	wire [4-1:0] node13172;
	wire [4-1:0] node13175;
	wire [4-1:0] node13178;
	wire [4-1:0] node13179;
	wire [4-1:0] node13181;
	wire [4-1:0] node13184;
	wire [4-1:0] node13186;
	wire [4-1:0] node13189;
	wire [4-1:0] node13190;
	wire [4-1:0] node13191;
	wire [4-1:0] node13194;
	wire [4-1:0] node13196;
	wire [4-1:0] node13199;
	wire [4-1:0] node13200;
	wire [4-1:0] node13202;
	wire [4-1:0] node13205;
	wire [4-1:0] node13208;
	wire [4-1:0] node13209;
	wire [4-1:0] node13210;
	wire [4-1:0] node13211;
	wire [4-1:0] node13212;
	wire [4-1:0] node13215;
	wire [4-1:0] node13218;
	wire [4-1:0] node13220;
	wire [4-1:0] node13223;
	wire [4-1:0] node13224;
	wire [4-1:0] node13228;
	wire [4-1:0] node13229;
	wire [4-1:0] node13232;
	wire [4-1:0] node13233;
	wire [4-1:0] node13234;
	wire [4-1:0] node13235;
	wire [4-1:0] node13241;
	wire [4-1:0] node13242;
	wire [4-1:0] node13243;
	wire [4-1:0] node13244;
	wire [4-1:0] node13245;
	wire [4-1:0] node13246;
	wire [4-1:0] node13249;
	wire [4-1:0] node13252;
	wire [4-1:0] node13254;
	wire [4-1:0] node13257;
	wire [4-1:0] node13258;
	wire [4-1:0] node13259;
	wire [4-1:0] node13264;
	wire [4-1:0] node13265;
	wire [4-1:0] node13267;
	wire [4-1:0] node13268;
	wire [4-1:0] node13270;
	wire [4-1:0] node13274;
	wire [4-1:0] node13276;
	wire [4-1:0] node13277;
	wire [4-1:0] node13281;
	wire [4-1:0] node13282;
	wire [4-1:0] node13283;
	wire [4-1:0] node13284;
	wire [4-1:0] node13285;
	wire [4-1:0] node13290;
	wire [4-1:0] node13291;
	wire [4-1:0] node13293;
	wire [4-1:0] node13297;
	wire [4-1:0] node13298;
	wire [4-1:0] node13299;
	wire [4-1:0] node13300;
	wire [4-1:0] node13304;
	wire [4-1:0] node13305;
	wire [4-1:0] node13310;
	wire [4-1:0] node13311;
	wire [4-1:0] node13312;
	wire [4-1:0] node13313;
	wire [4-1:0] node13314;
	wire [4-1:0] node13315;
	wire [4-1:0] node13316;
	wire [4-1:0] node13318;
	wire [4-1:0] node13319;
	wire [4-1:0] node13323;
	wire [4-1:0] node13324;
	wire [4-1:0] node13327;
	wire [4-1:0] node13330;
	wire [4-1:0] node13331;
	wire [4-1:0] node13334;
	wire [4-1:0] node13336;
	wire [4-1:0] node13339;
	wire [4-1:0] node13340;
	wire [4-1:0] node13341;
	wire [4-1:0] node13342;
	wire [4-1:0] node13345;
	wire [4-1:0] node13348;
	wire [4-1:0] node13349;
	wire [4-1:0] node13353;
	wire [4-1:0] node13354;
	wire [4-1:0] node13357;
	wire [4-1:0] node13360;
	wire [4-1:0] node13361;
	wire [4-1:0] node13362;
	wire [4-1:0] node13363;
	wire [4-1:0] node13366;
	wire [4-1:0] node13367;
	wire [4-1:0] node13371;
	wire [4-1:0] node13372;
	wire [4-1:0] node13373;
	wire [4-1:0] node13376;
	wire [4-1:0] node13380;
	wire [4-1:0] node13381;
	wire [4-1:0] node13382;
	wire [4-1:0] node13383;
	wire [4-1:0] node13388;
	wire [4-1:0] node13389;
	wire [4-1:0] node13392;
	wire [4-1:0] node13395;
	wire [4-1:0] node13396;
	wire [4-1:0] node13397;
	wire [4-1:0] node13398;
	wire [4-1:0] node13399;
	wire [4-1:0] node13402;
	wire [4-1:0] node13403;
	wire [4-1:0] node13406;
	wire [4-1:0] node13409;
	wire [4-1:0] node13410;
	wire [4-1:0] node13412;
	wire [4-1:0] node13413;
	wire [4-1:0] node13417;
	wire [4-1:0] node13418;
	wire [4-1:0] node13422;
	wire [4-1:0] node13423;
	wire [4-1:0] node13425;
	wire [4-1:0] node13428;
	wire [4-1:0] node13431;
	wire [4-1:0] node13432;
	wire [4-1:0] node13433;
	wire [4-1:0] node13434;
	wire [4-1:0] node13435;
	wire [4-1:0] node13438;
	wire [4-1:0] node13442;
	wire [4-1:0] node13443;
	wire [4-1:0] node13447;
	wire [4-1:0] node13448;
	wire [4-1:0] node13450;
	wire [4-1:0] node13453;
	wire [4-1:0] node13454;
	wire [4-1:0] node13457;
	wire [4-1:0] node13460;
	wire [4-1:0] node13461;
	wire [4-1:0] node13462;
	wire [4-1:0] node13463;
	wire [4-1:0] node13464;
	wire [4-1:0] node13467;
	wire [4-1:0] node13469;
	wire [4-1:0] node13470;
	wire [4-1:0] node13472;
	wire [4-1:0] node13475;
	wire [4-1:0] node13476;
	wire [4-1:0] node13480;
	wire [4-1:0] node13481;
	wire [4-1:0] node13482;
	wire [4-1:0] node13483;
	wire [4-1:0] node13487;
	wire [4-1:0] node13490;
	wire [4-1:0] node13491;
	wire [4-1:0] node13492;
	wire [4-1:0] node13495;
	wire [4-1:0] node13498;
	wire [4-1:0] node13499;
	wire [4-1:0] node13502;
	wire [4-1:0] node13504;
	wire [4-1:0] node13507;
	wire [4-1:0] node13508;
	wire [4-1:0] node13509;
	wire [4-1:0] node13511;
	wire [4-1:0] node13514;
	wire [4-1:0] node13516;
	wire [4-1:0] node13517;
	wire [4-1:0] node13518;
	wire [4-1:0] node13521;
	wire [4-1:0] node13525;
	wire [4-1:0] node13526;
	wire [4-1:0] node13528;
	wire [4-1:0] node13530;
	wire [4-1:0] node13534;
	wire [4-1:0] node13535;
	wire [4-1:0] node13536;
	wire [4-1:0] node13537;
	wire [4-1:0] node13539;
	wire [4-1:0] node13540;
	wire [4-1:0] node13543;
	wire [4-1:0] node13547;
	wire [4-1:0] node13548;
	wire [4-1:0] node13550;
	wire [4-1:0] node13553;
	wire [4-1:0] node13556;
	wire [4-1:0] node13557;
	wire [4-1:0] node13558;
	wire [4-1:0] node13559;
	wire [4-1:0] node13561;
	wire [4-1:0] node13567;
	wire [4-1:0] node13569;
	wire [4-1:0] node13570;
	wire [4-1:0] node13572;
	wire [4-1:0] node13573;
	wire [4-1:0] node13574;
	wire [4-1:0] node13575;
	wire [4-1:0] node13576;
	wire [4-1:0] node13577;
	wire [4-1:0] node13579;
	wire [4-1:0] node13582;
	wire [4-1:0] node13583;
	wire [4-1:0] node13588;
	wire [4-1:0] node13589;
	wire [4-1:0] node13590;
	wire [4-1:0] node13592;
	wire [4-1:0] node13593;
	wire [4-1:0] node13597;
	wire [4-1:0] node13598;
	wire [4-1:0] node13599;
	wire [4-1:0] node13604;
	wire [4-1:0] node13605;
	wire [4-1:0] node13607;
	wire [4-1:0] node13610;
	wire [4-1:0] node13612;
	wire [4-1:0] node13615;
	wire [4-1:0] node13616;
	wire [4-1:0] node13617;
	wire [4-1:0] node13618;
	wire [4-1:0] node13619;
	wire [4-1:0] node13623;
	wire [4-1:0] node13624;
	wire [4-1:0] node13628;
	wire [4-1:0] node13629;
	wire [4-1:0] node13631;
	wire [4-1:0] node13632;
	wire [4-1:0] node13637;
	wire [4-1:0] node13638;
	wire [4-1:0] node13639;
	wire [4-1:0] node13640;
	wire [4-1:0] node13641;
	wire [4-1:0] node13642;
	wire [4-1:0] node13648;
	wire [4-1:0] node13649;
	wire [4-1:0] node13650;
	wire [4-1:0] node13653;
	wire [4-1:0] node13657;
	wire [4-1:0] node13658;
	wire [4-1:0] node13659;
	wire [4-1:0] node13663;
	wire [4-1:0] node13665;
	wire [4-1:0] node13666;
	wire [4-1:0] node13669;
	wire [4-1:0] node13673;
	wire [4-1:0] node13674;
	wire [4-1:0] node13675;
	wire [4-1:0] node13676;
	wire [4-1:0] node13677;
	wire [4-1:0] node13678;
	wire [4-1:0] node13679;
	wire [4-1:0] node13680;
	wire [4-1:0] node13681;
	wire [4-1:0] node13685;
	wire [4-1:0] node13687;
	wire [4-1:0] node13690;
	wire [4-1:0] node13691;
	wire [4-1:0] node13692;
	wire [4-1:0] node13696;
	wire [4-1:0] node13697;
	wire [4-1:0] node13701;
	wire [4-1:0] node13702;
	wire [4-1:0] node13703;
	wire [4-1:0] node13705;
	wire [4-1:0] node13707;
	wire [4-1:0] node13710;
	wire [4-1:0] node13711;
	wire [4-1:0] node13714;
	wire [4-1:0] node13715;
	wire [4-1:0] node13719;
	wire [4-1:0] node13720;
	wire [4-1:0] node13721;
	wire [4-1:0] node13725;
	wire [4-1:0] node13728;
	wire [4-1:0] node13729;
	wire [4-1:0] node13730;
	wire [4-1:0] node13733;
	wire [4-1:0] node13734;
	wire [4-1:0] node13737;
	wire [4-1:0] node13740;
	wire [4-1:0] node13741;
	wire [4-1:0] node13742;
	wire [4-1:0] node13745;
	wire [4-1:0] node13747;
	wire [4-1:0] node13750;
	wire [4-1:0] node13751;
	wire [4-1:0] node13754;
	wire [4-1:0] node13755;
	wire [4-1:0] node13759;
	wire [4-1:0] node13760;
	wire [4-1:0] node13761;
	wire [4-1:0] node13762;
	wire [4-1:0] node13763;
	wire [4-1:0] node13764;
	wire [4-1:0] node13768;
	wire [4-1:0] node13771;
	wire [4-1:0] node13772;
	wire [4-1:0] node13774;
	wire [4-1:0] node13775;
	wire [4-1:0] node13779;
	wire [4-1:0] node13782;
	wire [4-1:0] node13783;
	wire [4-1:0] node13784;
	wire [4-1:0] node13786;
	wire [4-1:0] node13790;
	wire [4-1:0] node13791;
	wire [4-1:0] node13792;
	wire [4-1:0] node13793;
	wire [4-1:0] node13798;
	wire [4-1:0] node13800;
	wire [4-1:0] node13802;
	wire [4-1:0] node13805;
	wire [4-1:0] node13806;
	wire [4-1:0] node13807;
	wire [4-1:0] node13808;
	wire [4-1:0] node13809;
	wire [4-1:0] node13813;
	wire [4-1:0] node13814;
	wire [4-1:0] node13818;
	wire [4-1:0] node13820;
	wire [4-1:0] node13822;
	wire [4-1:0] node13825;
	wire [4-1:0] node13826;
	wire [4-1:0] node13827;
	wire [4-1:0] node13828;
	wire [4-1:0] node13833;
	wire [4-1:0] node13835;
	wire [4-1:0] node13838;
	wire [4-1:0] node13839;
	wire [4-1:0] node13840;
	wire [4-1:0] node13841;
	wire [4-1:0] node13842;
	wire [4-1:0] node13844;
	wire [4-1:0] node13846;
	wire [4-1:0] node13849;
	wire [4-1:0] node13851;
	wire [4-1:0] node13852;
	wire [4-1:0] node13855;
	wire [4-1:0] node13858;
	wire [4-1:0] node13859;
	wire [4-1:0] node13860;
	wire [4-1:0] node13863;
	wire [4-1:0] node13865;
	wire [4-1:0] node13868;
	wire [4-1:0] node13869;
	wire [4-1:0] node13871;
	wire [4-1:0] node13873;
	wire [4-1:0] node13876;
	wire [4-1:0] node13877;
	wire [4-1:0] node13881;
	wire [4-1:0] node13882;
	wire [4-1:0] node13883;
	wire [4-1:0] node13884;
	wire [4-1:0] node13886;
	wire [4-1:0] node13890;
	wire [4-1:0] node13891;
	wire [4-1:0] node13893;
	wire [4-1:0] node13894;
	wire [4-1:0] node13899;
	wire [4-1:0] node13900;
	wire [4-1:0] node13901;
	wire [4-1:0] node13904;
	wire [4-1:0] node13905;
	wire [4-1:0] node13906;
	wire [4-1:0] node13911;
	wire [4-1:0] node13912;
	wire [4-1:0] node13916;
	wire [4-1:0] node13917;
	wire [4-1:0] node13918;
	wire [4-1:0] node13919;
	wire [4-1:0] node13921;
	wire [4-1:0] node13924;
	wire [4-1:0] node13925;
	wire [4-1:0] node13926;
	wire [4-1:0] node13931;
	wire [4-1:0] node13932;
	wire [4-1:0] node13933;
	wire [4-1:0] node13937;
	wire [4-1:0] node13939;
	wire [4-1:0] node13940;
	wire [4-1:0] node13944;
	wire [4-1:0] node13945;
	wire [4-1:0] node13946;
	wire [4-1:0] node13948;
	wire [4-1:0] node13949;
	wire [4-1:0] node13953;
	wire [4-1:0] node13957;
	wire [4-1:0] node13959;
	wire [4-1:0] node13960;
	wire [4-1:0] node13961;
	wire [4-1:0] node13962;
	wire [4-1:0] node13963;
	wire [4-1:0] node13964;
	wire [4-1:0] node13967;
	wire [4-1:0] node13968;
	wire [4-1:0] node13972;
	wire [4-1:0] node13974;
	wire [4-1:0] node13977;
	wire [4-1:0] node13978;
	wire [4-1:0] node13979;
	wire [4-1:0] node13982;
	wire [4-1:0] node13983;
	wire [4-1:0] node13986;
	wire [4-1:0] node13987;
	wire [4-1:0] node13991;
	wire [4-1:0] node13993;
	wire [4-1:0] node13994;
	wire [4-1:0] node13997;
	wire [4-1:0] node14001;
	wire [4-1:0] node14002;
	wire [4-1:0] node14003;
	wire [4-1:0] node14004;
	wire [4-1:0] node14005;
	wire [4-1:0] node14006;
	wire [4-1:0] node14007;
	wire [4-1:0] node14013;
	wire [4-1:0] node14014;
	wire [4-1:0] node14015;
	wire [4-1:0] node14018;
	wire [4-1:0] node14022;
	wire [4-1:0] node14023;
	wire [4-1:0] node14024;
	wire [4-1:0] node14027;
	wire [4-1:0] node14028;
	wire [4-1:0] node14030;
	wire [4-1:0] node14035;
	wire [4-1:0] node14036;
	wire [4-1:0] node14037;
	wire [4-1:0] node14038;
	wire [4-1:0] node14042;
	wire [4-1:0] node14044;
	wire [4-1:0] node14048;
	wire [4-1:0] node14049;
	wire [4-1:0] node14050;
	wire [4-1:0] node14051;
	wire [4-1:0] node14052;
	wire [4-1:0] node14053;
	wire [4-1:0] node14054;
	wire [4-1:0] node14055;
	wire [4-1:0] node14056;
	wire [4-1:0] node14058;
	wire [4-1:0] node14059;
	wire [4-1:0] node14060;
	wire [4-1:0] node14064;
	wire [4-1:0] node14066;
	wire [4-1:0] node14070;
	wire [4-1:0] node14071;
	wire [4-1:0] node14072;
	wire [4-1:0] node14073;
	wire [4-1:0] node14074;
	wire [4-1:0] node14076;
	wire [4-1:0] node14078;
	wire [4-1:0] node14081;
	wire [4-1:0] node14082;
	wire [4-1:0] node14086;
	wire [4-1:0] node14089;
	wire [4-1:0] node14090;
	wire [4-1:0] node14091;
	wire [4-1:0] node14093;
	wire [4-1:0] node14094;
	wire [4-1:0] node14098;
	wire [4-1:0] node14099;
	wire [4-1:0] node14103;
	wire [4-1:0] node14104;
	wire [4-1:0] node14105;
	wire [4-1:0] node14107;
	wire [4-1:0] node14111;
	wire [4-1:0] node14114;
	wire [4-1:0] node14115;
	wire [4-1:0] node14117;
	wire [4-1:0] node14118;
	wire [4-1:0] node14121;
	wire [4-1:0] node14122;
	wire [4-1:0] node14125;
	wire [4-1:0] node14129;
	wire [4-1:0] node14130;
	wire [4-1:0] node14131;
	wire [4-1:0] node14132;
	wire [4-1:0] node14133;
	wire [4-1:0] node14134;
	wire [4-1:0] node14138;
	wire [4-1:0] node14139;
	wire [4-1:0] node14141;
	wire [4-1:0] node14145;
	wire [4-1:0] node14146;
	wire [4-1:0] node14147;
	wire [4-1:0] node14148;
	wire [4-1:0] node14152;
	wire [4-1:0] node14154;
	wire [4-1:0] node14157;
	wire [4-1:0] node14158;
	wire [4-1:0] node14161;
	wire [4-1:0] node14162;
	wire [4-1:0] node14166;
	wire [4-1:0] node14167;
	wire [4-1:0] node14169;
	wire [4-1:0] node14171;
	wire [4-1:0] node14173;
	wire [4-1:0] node14176;
	wire [4-1:0] node14177;
	wire [4-1:0] node14178;
	wire [4-1:0] node14179;
	wire [4-1:0] node14184;
	wire [4-1:0] node14185;
	wire [4-1:0] node14186;
	wire [4-1:0] node14190;
	wire [4-1:0] node14192;
	wire [4-1:0] node14194;
	wire [4-1:0] node14197;
	wire [4-1:0] node14198;
	wire [4-1:0] node14199;
	wire [4-1:0] node14200;
	wire [4-1:0] node14201;
	wire [4-1:0] node14203;
	wire [4-1:0] node14204;
	wire [4-1:0] node14209;
	wire [4-1:0] node14210;
	wire [4-1:0] node14214;
	wire [4-1:0] node14215;
	wire [4-1:0] node14217;
	wire [4-1:0] node14220;
	wire [4-1:0] node14221;
	wire [4-1:0] node14225;
	wire [4-1:0] node14226;
	wire [4-1:0] node14227;
	wire [4-1:0] node14231;
	wire [4-1:0] node14232;
	wire [4-1:0] node14233;
	wire [4-1:0] node14235;
	wire [4-1:0] node14238;
	wire [4-1:0] node14239;
	wire [4-1:0] node14241;
	wire [4-1:0] node14245;
	wire [4-1:0] node14246;
	wire [4-1:0] node14248;
	wire [4-1:0] node14251;
	wire [4-1:0] node14254;
	wire [4-1:0] node14255;
	wire [4-1:0] node14256;
	wire [4-1:0] node14257;
	wire [4-1:0] node14258;
	wire [4-1:0] node14259;
	wire [4-1:0] node14261;
	wire [4-1:0] node14264;
	wire [4-1:0] node14266;
	wire [4-1:0] node14268;
	wire [4-1:0] node14271;
	wire [4-1:0] node14272;
	wire [4-1:0] node14273;
	wire [4-1:0] node14277;
	wire [4-1:0] node14279;
	wire [4-1:0] node14280;
	wire [4-1:0] node14284;
	wire [4-1:0] node14285;
	wire [4-1:0] node14287;
	wire [4-1:0] node14290;
	wire [4-1:0] node14292;
	wire [4-1:0] node14295;
	wire [4-1:0] node14296;
	wire [4-1:0] node14297;
	wire [4-1:0] node14298;
	wire [4-1:0] node14300;
	wire [4-1:0] node14303;
	wire [4-1:0] node14304;
	wire [4-1:0] node14307;
	wire [4-1:0] node14310;
	wire [4-1:0] node14311;
	wire [4-1:0] node14314;
	wire [4-1:0] node14316;
	wire [4-1:0] node14317;
	wire [4-1:0] node14321;
	wire [4-1:0] node14322;
	wire [4-1:0] node14324;
	wire [4-1:0] node14327;
	wire [4-1:0] node14328;
	wire [4-1:0] node14330;
	wire [4-1:0] node14333;
	wire [4-1:0] node14334;
	wire [4-1:0] node14338;
	wire [4-1:0] node14339;
	wire [4-1:0] node14340;
	wire [4-1:0] node14341;
	wire [4-1:0] node14342;
	wire [4-1:0] node14344;
	wire [4-1:0] node14347;
	wire [4-1:0] node14350;
	wire [4-1:0] node14351;
	wire [4-1:0] node14352;
	wire [4-1:0] node14355;
	wire [4-1:0] node14358;
	wire [4-1:0] node14359;
	wire [4-1:0] node14360;
	wire [4-1:0] node14365;
	wire [4-1:0] node14366;
	wire [4-1:0] node14367;
	wire [4-1:0] node14368;
	wire [4-1:0] node14372;
	wire [4-1:0] node14374;
	wire [4-1:0] node14377;
	wire [4-1:0] node14378;
	wire [4-1:0] node14379;
	wire [4-1:0] node14381;
	wire [4-1:0] node14385;
	wire [4-1:0] node14388;
	wire [4-1:0] node14389;
	wire [4-1:0] node14390;
	wire [4-1:0] node14391;
	wire [4-1:0] node14392;
	wire [4-1:0] node14396;
	wire [4-1:0] node14397;
	wire [4-1:0] node14401;
	wire [4-1:0] node14402;
	wire [4-1:0] node14403;
	wire [4-1:0] node14407;
	wire [4-1:0] node14408;
	wire [4-1:0] node14412;
	wire [4-1:0] node14413;
	wire [4-1:0] node14414;
	wire [4-1:0] node14415;
	wire [4-1:0] node14419;
	wire [4-1:0] node14421;
	wire [4-1:0] node14424;
	wire [4-1:0] node14425;
	wire [4-1:0] node14426;
	wire [4-1:0] node14428;
	wire [4-1:0] node14431;
	wire [4-1:0] node14433;
	wire [4-1:0] node14436;
	wire [4-1:0] node14437;
	wire [4-1:0] node14440;
	wire [4-1:0] node14441;
	wire [4-1:0] node14445;
	wire [4-1:0] node14447;
	wire [4-1:0] node14448;
	wire [4-1:0] node14449;
	wire [4-1:0] node14451;
	wire [4-1:0] node14452;
	wire [4-1:0] node14454;
	wire [4-1:0] node14456;
	wire [4-1:0] node14457;
	wire [4-1:0] node14462;
	wire [4-1:0] node14463;
	wire [4-1:0] node14464;
	wire [4-1:0] node14465;
	wire [4-1:0] node14467;
	wire [4-1:0] node14468;
	wire [4-1:0] node14471;
	wire [4-1:0] node14474;
	wire [4-1:0] node14475;
	wire [4-1:0] node14477;
	wire [4-1:0] node14480;
	wire [4-1:0] node14481;
	wire [4-1:0] node14485;
	wire [4-1:0] node14486;
	wire [4-1:0] node14489;
	wire [4-1:0] node14490;
	wire [4-1:0] node14491;
	wire [4-1:0] node14492;
	wire [4-1:0] node14496;
	wire [4-1:0] node14498;
	wire [4-1:0] node14502;
	wire [4-1:0] node14504;
	wire [4-1:0] node14505;
	wire [4-1:0] node14506;
	wire [4-1:0] node14510;
	wire [4-1:0] node14511;
	wire [4-1:0] node14512;
	wire [4-1:0] node14514;
	wire [4-1:0] node14518;
	wire [4-1:0] node14520;
	wire [4-1:0] node14523;
	wire [4-1:0] node14524;
	wire [4-1:0] node14525;
	wire [4-1:0] node14526;
	wire [4-1:0] node14527;
	wire [4-1:0] node14529;
	wire [4-1:0] node14531;
	wire [4-1:0] node14532;
	wire [4-1:0] node14536;
	wire [4-1:0] node14537;
	wire [4-1:0] node14539;
	wire [4-1:0] node14543;
	wire [4-1:0] node14544;
	wire [4-1:0] node14545;
	wire [4-1:0] node14549;
	wire [4-1:0] node14550;
	wire [4-1:0] node14554;
	wire [4-1:0] node14555;
	wire [4-1:0] node14556;
	wire [4-1:0] node14557;
	wire [4-1:0] node14559;
	wire [4-1:0] node14560;
	wire [4-1:0] node14564;
	wire [4-1:0] node14565;
	wire [4-1:0] node14569;
	wire [4-1:0] node14570;
	wire [4-1:0] node14571;
	wire [4-1:0] node14575;
	wire [4-1:0] node14578;
	wire [4-1:0] node14579;
	wire [4-1:0] node14580;
	wire [4-1:0] node14584;
	wire [4-1:0] node14586;
	wire [4-1:0] node14589;
	wire [4-1:0] node14590;
	wire [4-1:0] node14591;
	wire [4-1:0] node14592;
	wire [4-1:0] node14593;
	wire [4-1:0] node14596;
	wire [4-1:0] node14597;
	wire [4-1:0] node14600;
	wire [4-1:0] node14603;
	wire [4-1:0] node14604;
	wire [4-1:0] node14605;
	wire [4-1:0] node14608;
	wire [4-1:0] node14611;
	wire [4-1:0] node14614;
	wire [4-1:0] node14615;
	wire [4-1:0] node14616;
	wire [4-1:0] node14617;
	wire [4-1:0] node14622;
	wire [4-1:0] node14623;
	wire [4-1:0] node14624;
	wire [4-1:0] node14629;
	wire [4-1:0] node14630;
	wire [4-1:0] node14631;
	wire [4-1:0] node14633;
	wire [4-1:0] node14634;
	wire [4-1:0] node14637;
	wire [4-1:0] node14640;
	wire [4-1:0] node14642;
	wire [4-1:0] node14645;
	wire [4-1:0] node14646;
	wire [4-1:0] node14648;
	wire [4-1:0] node14649;
	wire [4-1:0] node14652;
	wire [4-1:0] node14655;
	wire [4-1:0] node14656;
	wire [4-1:0] node14659;
	wire [4-1:0] node14661;
	wire [4-1:0] node14665;
	wire [4-1:0] node14666;
	wire [4-1:0] node14667;
	wire [4-1:0] node14668;
	wire [4-1:0] node14669;
	wire [4-1:0] node14670;
	wire [4-1:0] node14671;
	wire [4-1:0] node14672;
	wire [4-1:0] node14673;
	wire [4-1:0] node14676;
	wire [4-1:0] node14677;
	wire [4-1:0] node14681;
	wire [4-1:0] node14682;
	wire [4-1:0] node14683;
	wire [4-1:0] node14684;
	wire [4-1:0] node14688;
	wire [4-1:0] node14690;
	wire [4-1:0] node14693;
	wire [4-1:0] node14696;
	wire [4-1:0] node14697;
	wire [4-1:0] node14698;
	wire [4-1:0] node14699;
	wire [4-1:0] node14701;
	wire [4-1:0] node14705;
	wire [4-1:0] node14706;
	wire [4-1:0] node14709;
	wire [4-1:0] node14712;
	wire [4-1:0] node14713;
	wire [4-1:0] node14714;
	wire [4-1:0] node14715;
	wire [4-1:0] node14719;
	wire [4-1:0] node14721;
	wire [4-1:0] node14724;
	wire [4-1:0] node14725;
	wire [4-1:0] node14727;
	wire [4-1:0] node14730;
	wire [4-1:0] node14733;
	wire [4-1:0] node14734;
	wire [4-1:0] node14735;
	wire [4-1:0] node14736;
	wire [4-1:0] node14738;
	wire [4-1:0] node14740;
	wire [4-1:0] node14743;
	wire [4-1:0] node14744;
	wire [4-1:0] node14746;
	wire [4-1:0] node14749;
	wire [4-1:0] node14750;
	wire [4-1:0] node14754;
	wire [4-1:0] node14755;
	wire [4-1:0] node14756;
	wire [4-1:0] node14760;
	wire [4-1:0] node14762;
	wire [4-1:0] node14765;
	wire [4-1:0] node14766;
	wire [4-1:0] node14767;
	wire [4-1:0] node14768;
	wire [4-1:0] node14771;
	wire [4-1:0] node14773;
	wire [4-1:0] node14774;
	wire [4-1:0] node14777;
	wire [4-1:0] node14780;
	wire [4-1:0] node14783;
	wire [4-1:0] node14784;
	wire [4-1:0] node14785;
	wire [4-1:0] node14786;
	wire [4-1:0] node14787;
	wire [4-1:0] node14791;
	wire [4-1:0] node14793;
	wire [4-1:0] node14796;
	wire [4-1:0] node14799;
	wire [4-1:0] node14800;
	wire [4-1:0] node14803;
	wire [4-1:0] node14805;
	wire [4-1:0] node14808;
	wire [4-1:0] node14809;
	wire [4-1:0] node14810;
	wire [4-1:0] node14811;
	wire [4-1:0] node14812;
	wire [4-1:0] node14814;
	wire [4-1:0] node14817;
	wire [4-1:0] node14818;
	wire [4-1:0] node14820;
	wire [4-1:0] node14824;
	wire [4-1:0] node14825;
	wire [4-1:0] node14827;
	wire [4-1:0] node14829;
	wire [4-1:0] node14832;
	wire [4-1:0] node14833;
	wire [4-1:0] node14834;
	wire [4-1:0] node14838;
	wire [4-1:0] node14841;
	wire [4-1:0] node14842;
	wire [4-1:0] node14843;
	wire [4-1:0] node14844;
	wire [4-1:0] node14847;
	wire [4-1:0] node14848;
	wire [4-1:0] node14850;
	wire [4-1:0] node14854;
	wire [4-1:0] node14855;
	wire [4-1:0] node14858;
	wire [4-1:0] node14860;
	wire [4-1:0] node14863;
	wire [4-1:0] node14864;
	wire [4-1:0] node14865;
	wire [4-1:0] node14867;
	wire [4-1:0] node14871;
	wire [4-1:0] node14872;
	wire [4-1:0] node14874;
	wire [4-1:0] node14875;
	wire [4-1:0] node14878;
	wire [4-1:0] node14881;
	wire [4-1:0] node14882;
	wire [4-1:0] node14885;
	wire [4-1:0] node14888;
	wire [4-1:0] node14889;
	wire [4-1:0] node14890;
	wire [4-1:0] node14891;
	wire [4-1:0] node14892;
	wire [4-1:0] node14893;
	wire [4-1:0] node14897;
	wire [4-1:0] node14898;
	wire [4-1:0] node14901;
	wire [4-1:0] node14904;
	wire [4-1:0] node14906;
	wire [4-1:0] node14907;
	wire [4-1:0] node14908;
	wire [4-1:0] node14913;
	wire [4-1:0] node14914;
	wire [4-1:0] node14915;
	wire [4-1:0] node14916;
	wire [4-1:0] node14921;
	wire [4-1:0] node14922;
	wire [4-1:0] node14923;
	wire [4-1:0] node14926;
	wire [4-1:0] node14928;
	wire [4-1:0] node14931;
	wire [4-1:0] node14932;
	wire [4-1:0] node14936;
	wire [4-1:0] node14937;
	wire [4-1:0] node14938;
	wire [4-1:0] node14940;
	wire [4-1:0] node14943;
	wire [4-1:0] node14946;
	wire [4-1:0] node14947;
	wire [4-1:0] node14949;
	wire [4-1:0] node14953;
	wire [4-1:0] node14954;
	wire [4-1:0] node14955;
	wire [4-1:0] node14956;
	wire [4-1:0] node14957;
	wire [4-1:0] node14959;
	wire [4-1:0] node14960;
	wire [4-1:0] node14963;
	wire [4-1:0] node14964;
	wire [4-1:0] node14968;
	wire [4-1:0] node14969;
	wire [4-1:0] node14971;
	wire [4-1:0] node14973;
	wire [4-1:0] node14976;
	wire [4-1:0] node14977;
	wire [4-1:0] node14978;
	wire [4-1:0] node14981;
	wire [4-1:0] node14984;
	wire [4-1:0] node14985;
	wire [4-1:0] node14989;
	wire [4-1:0] node14990;
	wire [4-1:0] node14991;
	wire [4-1:0] node14994;
	wire [4-1:0] node14995;
	wire [4-1:0] node14997;
	wire [4-1:0] node15001;
	wire [4-1:0] node15002;
	wire [4-1:0] node15004;
	wire [4-1:0] node15007;
	wire [4-1:0] node15008;
	wire [4-1:0] node15011;
	wire [4-1:0] node15013;
	wire [4-1:0] node15016;
	wire [4-1:0] node15017;
	wire [4-1:0] node15018;
	wire [4-1:0] node15019;
	wire [4-1:0] node15021;
	wire [4-1:0] node15022;
	wire [4-1:0] node15026;
	wire [4-1:0] node15027;
	wire [4-1:0] node15029;
	wire [4-1:0] node15032;
	wire [4-1:0] node15035;
	wire [4-1:0] node15036;
	wire [4-1:0] node15037;
	wire [4-1:0] node15039;
	wire [4-1:0] node15043;
	wire [4-1:0] node15044;
	wire [4-1:0] node15045;
	wire [4-1:0] node15048;
	wire [4-1:0] node15052;
	wire [4-1:0] node15053;
	wire [4-1:0] node15054;
	wire [4-1:0] node15055;
	wire [4-1:0] node15058;
	wire [4-1:0] node15059;
	wire [4-1:0] node15062;
	wire [4-1:0] node15065;
	wire [4-1:0] node15067;
	wire [4-1:0] node15068;
	wire [4-1:0] node15072;
	wire [4-1:0] node15073;
	wire [4-1:0] node15075;
	wire [4-1:0] node15077;
	wire [4-1:0] node15080;
	wire [4-1:0] node15081;
	wire [4-1:0] node15084;
	wire [4-1:0] node15087;
	wire [4-1:0] node15088;
	wire [4-1:0] node15089;
	wire [4-1:0] node15090;
	wire [4-1:0] node15091;
	wire [4-1:0] node15094;
	wire [4-1:0] node15095;
	wire [4-1:0] node15098;
	wire [4-1:0] node15101;
	wire [4-1:0] node15102;
	wire [4-1:0] node15103;
	wire [4-1:0] node15107;
	wire [4-1:0] node15108;
	wire [4-1:0] node15109;
	wire [4-1:0] node15112;
	wire [4-1:0] node15115;
	wire [4-1:0] node15116;
	wire [4-1:0] node15120;
	wire [4-1:0] node15121;
	wire [4-1:0] node15122;
	wire [4-1:0] node15123;
	wire [4-1:0] node15126;
	wire [4-1:0] node15127;
	wire [4-1:0] node15131;
	wire [4-1:0] node15133;
	wire [4-1:0] node15135;
	wire [4-1:0] node15138;
	wire [4-1:0] node15139;
	wire [4-1:0] node15141;
	wire [4-1:0] node15143;
	wire [4-1:0] node15146;
	wire [4-1:0] node15147;
	wire [4-1:0] node15149;
	wire [4-1:0] node15150;
	wire [4-1:0] node15153;
	wire [4-1:0] node15157;
	wire [4-1:0] node15158;
	wire [4-1:0] node15159;
	wire [4-1:0] node15160;
	wire [4-1:0] node15161;
	wire [4-1:0] node15165;
	wire [4-1:0] node15167;
	wire [4-1:0] node15170;
	wire [4-1:0] node15171;
	wire [4-1:0] node15172;
	wire [4-1:0] node15173;
	wire [4-1:0] node15175;
	wire [4-1:0] node15178;
	wire [4-1:0] node15179;
	wire [4-1:0] node15183;
	wire [4-1:0] node15184;
	wire [4-1:0] node15188;
	wire [4-1:0] node15190;
	wire [4-1:0] node15193;
	wire [4-1:0] node15194;
	wire [4-1:0] node15196;
	wire [4-1:0] node15198;
	wire [4-1:0] node15201;
	wire [4-1:0] node15202;
	wire [4-1:0] node15206;
	wire [4-1:0] node15207;
	wire [4-1:0] node15208;
	wire [4-1:0] node15209;
	wire [4-1:0] node15210;
	wire [4-1:0] node15212;
	wire [4-1:0] node15214;
	wire [4-1:0] node15215;
	wire [4-1:0] node15217;
	wire [4-1:0] node15222;
	wire [4-1:0] node15223;
	wire [4-1:0] node15224;
	wire [4-1:0] node15225;
	wire [4-1:0] node15226;
	wire [4-1:0] node15229;
	wire [4-1:0] node15231;
	wire [4-1:0] node15234;
	wire [4-1:0] node15235;
	wire [4-1:0] node15238;
	wire [4-1:0] node15241;
	wire [4-1:0] node15242;
	wire [4-1:0] node15244;
	wire [4-1:0] node15247;
	wire [4-1:0] node15248;
	wire [4-1:0] node15249;
	wire [4-1:0] node15251;
	wire [4-1:0] node15254;
	wire [4-1:0] node15258;
	wire [4-1:0] node15260;
	wire [4-1:0] node15261;
	wire [4-1:0] node15263;
	wire [4-1:0] node15266;
	wire [4-1:0] node15267;
	wire [4-1:0] node15270;
	wire [4-1:0] node15272;
	wire [4-1:0] node15275;
	wire [4-1:0] node15276;
	wire [4-1:0] node15277;
	wire [4-1:0] node15278;
	wire [4-1:0] node15279;
	wire [4-1:0] node15281;
	wire [4-1:0] node15282;
	wire [4-1:0] node15285;
	wire [4-1:0] node15288;
	wire [4-1:0] node15289;
	wire [4-1:0] node15293;
	wire [4-1:0] node15294;
	wire [4-1:0] node15295;
	wire [4-1:0] node15297;
	wire [4-1:0] node15298;
	wire [4-1:0] node15302;
	wire [4-1:0] node15304;
	wire [4-1:0] node15307;
	wire [4-1:0] node15308;
	wire [4-1:0] node15309;
	wire [4-1:0] node15311;
	wire [4-1:0] node15314;
	wire [4-1:0] node15318;
	wire [4-1:0] node15319;
	wire [4-1:0] node15320;
	wire [4-1:0] node15321;
	wire [4-1:0] node15324;
	wire [4-1:0] node15325;
	wire [4-1:0] node15328;
	wire [4-1:0] node15329;
	wire [4-1:0] node15333;
	wire [4-1:0] node15334;
	wire [4-1:0] node15336;
	wire [4-1:0] node15339;
	wire [4-1:0] node15342;
	wire [4-1:0] node15343;
	wire [4-1:0] node15344;
	wire [4-1:0] node15345;
	wire [4-1:0] node15349;
	wire [4-1:0] node15352;
	wire [4-1:0] node15353;
	wire [4-1:0] node15356;
	wire [4-1:0] node15357;
	wire [4-1:0] node15361;
	wire [4-1:0] node15362;
	wire [4-1:0] node15363;
	wire [4-1:0] node15364;
	wire [4-1:0] node15366;
	wire [4-1:0] node15367;
	wire [4-1:0] node15369;
	wire [4-1:0] node15373;
	wire [4-1:0] node15374;
	wire [4-1:0] node15376;
	wire [4-1:0] node15379;
	wire [4-1:0] node15382;
	wire [4-1:0] node15383;
	wire [4-1:0] node15385;
	wire [4-1:0] node15388;
	wire [4-1:0] node15390;
	wire [4-1:0] node15391;
	wire [4-1:0] node15395;
	wire [4-1:0] node15396;
	wire [4-1:0] node15397;
	wire [4-1:0] node15398;
	wire [4-1:0] node15399;
	wire [4-1:0] node15402;
	wire [4-1:0] node15406;
	wire [4-1:0] node15407;
	wire [4-1:0] node15408;
	wire [4-1:0] node15412;
	wire [4-1:0] node15413;
	wire [4-1:0] node15417;
	wire [4-1:0] node15418;
	wire [4-1:0] node15420;
	wire [4-1:0] node15423;
	wire [4-1:0] node15424;
	wire [4-1:0] node15426;
	wire [4-1:0] node15429;
	wire [4-1:0] node15431;
	wire [4-1:0] node15435;
	wire [4-1:0] node15436;
	wire [4-1:0] node15437;
	wire [4-1:0] node15438;
	wire [4-1:0] node15439;
	wire [4-1:0] node15440;
	wire [4-1:0] node15441;
	wire [4-1:0] node15442;
	wire [4-1:0] node15443;
	wire [4-1:0] node15444;
	wire [4-1:0] node15445;
	wire [4-1:0] node15449;
	wire [4-1:0] node15453;
	wire [4-1:0] node15454;
	wire [4-1:0] node15457;
	wire [4-1:0] node15459;
	wire [4-1:0] node15462;
	wire [4-1:0] node15463;
	wire [4-1:0] node15464;
	wire [4-1:0] node15468;
	wire [4-1:0] node15469;
	wire [4-1:0] node15470;
	wire [4-1:0] node15474;
	wire [4-1:0] node15475;
	wire [4-1:0] node15478;
	wire [4-1:0] node15479;
	wire [4-1:0] node15483;
	wire [4-1:0] node15484;
	wire [4-1:0] node15485;
	wire [4-1:0] node15486;
	wire [4-1:0] node15487;
	wire [4-1:0] node15489;
	wire [4-1:0] node15493;
	wire [4-1:0] node15496;
	wire [4-1:0] node15497;
	wire [4-1:0] node15500;
	wire [4-1:0] node15501;
	wire [4-1:0] node15505;
	wire [4-1:0] node15506;
	wire [4-1:0] node15507;
	wire [4-1:0] node15508;
	wire [4-1:0] node15512;
	wire [4-1:0] node15515;
	wire [4-1:0] node15518;
	wire [4-1:0] node15519;
	wire [4-1:0] node15520;
	wire [4-1:0] node15521;
	wire [4-1:0] node15522;
	wire [4-1:0] node15526;
	wire [4-1:0] node15528;
	wire [4-1:0] node15529;
	wire [4-1:0] node15532;
	wire [4-1:0] node15535;
	wire [4-1:0] node15536;
	wire [4-1:0] node15537;
	wire [4-1:0] node15541;
	wire [4-1:0] node15542;
	wire [4-1:0] node15544;
	wire [4-1:0] node15547;
	wire [4-1:0] node15548;
	wire [4-1:0] node15553;
	wire [4-1:0] node15554;
	wire [4-1:0] node15555;
	wire [4-1:0] node15556;
	wire [4-1:0] node15558;
	wire [4-1:0] node15559;
	wire [4-1:0] node15561;
	wire [4-1:0] node15564;
	wire [4-1:0] node15567;
	wire [4-1:0] node15568;
	wire [4-1:0] node15569;
	wire [4-1:0] node15572;
	wire [4-1:0] node15575;
	wire [4-1:0] node15576;
	wire [4-1:0] node15580;
	wire [4-1:0] node15581;
	wire [4-1:0] node15582;
	wire [4-1:0] node15584;
	wire [4-1:0] node15585;
	wire [4-1:0] node15589;
	wire [4-1:0] node15592;
	wire [4-1:0] node15593;
	wire [4-1:0] node15595;
	wire [4-1:0] node15596;
	wire [4-1:0] node15599;
	wire [4-1:0] node15602;
	wire [4-1:0] node15603;
	wire [4-1:0] node15606;
	wire [4-1:0] node15608;
	wire [4-1:0] node15609;
	wire [4-1:0] node15613;
	wire [4-1:0] node15614;
	wire [4-1:0] node15615;
	wire [4-1:0] node15616;
	wire [4-1:0] node15617;
	wire [4-1:0] node15618;
	wire [4-1:0] node15621;
	wire [4-1:0] node15624;
	wire [4-1:0] node15625;
	wire [4-1:0] node15629;
	wire [4-1:0] node15630;
	wire [4-1:0] node15632;
	wire [4-1:0] node15636;
	wire [4-1:0] node15637;
	wire [4-1:0] node15638;
	wire [4-1:0] node15639;
	wire [4-1:0] node15642;
	wire [4-1:0] node15645;
	wire [4-1:0] node15648;
	wire [4-1:0] node15649;
	wire [4-1:0] node15653;
	wire [4-1:0] node15654;
	wire [4-1:0] node15655;
	wire [4-1:0] node15656;
	wire [4-1:0] node15657;
	wire [4-1:0] node15662;
	wire [4-1:0] node15663;
	wire [4-1:0] node15665;
	wire [4-1:0] node15667;
	wire [4-1:0] node15672;
	wire [4-1:0] node15673;
	wire [4-1:0] node15674;
	wire [4-1:0] node15675;
	wire [4-1:0] node15676;
	wire [4-1:0] node15677;
	wire [4-1:0] node15678;
	wire [4-1:0] node15681;
	wire [4-1:0] node15683;
	wire [4-1:0] node15684;
	wire [4-1:0] node15688;
	wire [4-1:0] node15689;
	wire [4-1:0] node15693;
	wire [4-1:0] node15694;
	wire [4-1:0] node15696;
	wire [4-1:0] node15697;
	wire [4-1:0] node15698;
	wire [4-1:0] node15703;
	wire [4-1:0] node15704;
	wire [4-1:0] node15705;
	wire [4-1:0] node15709;
	wire [4-1:0] node15711;
	wire [4-1:0] node15714;
	wire [4-1:0] node15715;
	wire [4-1:0] node15716;
	wire [4-1:0] node15717;
	wire [4-1:0] node15718;
	wire [4-1:0] node15719;
	wire [4-1:0] node15724;
	wire [4-1:0] node15727;
	wire [4-1:0] node15728;
	wire [4-1:0] node15729;
	wire [4-1:0] node15734;
	wire [4-1:0] node15735;
	wire [4-1:0] node15736;
	wire [4-1:0] node15738;
	wire [4-1:0] node15741;
	wire [4-1:0] node15742;
	wire [4-1:0] node15744;
	wire [4-1:0] node15748;
	wire [4-1:0] node15749;
	wire [4-1:0] node15753;
	wire [4-1:0] node15754;
	wire [4-1:0] node15755;
	wire [4-1:0] node15756;
	wire [4-1:0] node15757;
	wire [4-1:0] node15760;
	wire [4-1:0] node15763;
	wire [4-1:0] node15764;
	wire [4-1:0] node15765;
	wire [4-1:0] node15768;
	wire [4-1:0] node15773;
	wire [4-1:0] node15774;
	wire [4-1:0] node15775;
	wire [4-1:0] node15776;
	wire [4-1:0] node15777;
	wire [4-1:0] node15780;
	wire [4-1:0] node15783;
	wire [4-1:0] node15784;
	wire [4-1:0] node15787;
	wire [4-1:0] node15790;
	wire [4-1:0] node15791;
	wire [4-1:0] node15793;
	wire [4-1:0] node15796;
	wire [4-1:0] node15797;
	wire [4-1:0] node15801;
	wire [4-1:0] node15802;
	wire [4-1:0] node15803;
	wire [4-1:0] node15806;
	wire [4-1:0] node15810;
	wire [4-1:0] node15811;
	wire [4-1:0] node15812;
	wire [4-1:0] node15813;
	wire [4-1:0] node15814;
	wire [4-1:0] node15815;
	wire [4-1:0] node15816;
	wire [4-1:0] node15817;
	wire [4-1:0] node15820;
	wire [4-1:0] node15824;
	wire [4-1:0] node15825;
	wire [4-1:0] node15828;
	wire [4-1:0] node15831;
	wire [4-1:0] node15832;
	wire [4-1:0] node15835;
	wire [4-1:0] node15836;
	wire [4-1:0] node15837;
	wire [4-1:0] node15841;
	wire [4-1:0] node15844;
	wire [4-1:0] node15845;
	wire [4-1:0] node15846;
	wire [4-1:0] node15847;
	wire [4-1:0] node15852;
	wire [4-1:0] node15853;
	wire [4-1:0] node15856;
	wire [4-1:0] node15858;
	wire [4-1:0] node15859;
	wire [4-1:0] node15862;
	wire [4-1:0] node15865;
	wire [4-1:0] node15866;
	wire [4-1:0] node15867;
	wire [4-1:0] node15868;
	wire [4-1:0] node15869;
	wire [4-1:0] node15872;
	wire [4-1:0] node15875;
	wire [4-1:0] node15876;
	wire [4-1:0] node15879;
	wire [4-1:0] node15881;
	wire [4-1:0] node15884;
	wire [4-1:0] node15885;
	wire [4-1:0] node15887;
	wire [4-1:0] node15890;
	wire [4-1:0] node15891;
	wire [4-1:0] node15894;
	wire [4-1:0] node15895;
	wire [4-1:0] node15899;
	wire [4-1:0] node15900;
	wire [4-1:0] node15901;
	wire [4-1:0] node15905;
	wire [4-1:0] node15906;
	wire [4-1:0] node15907;
	wire [4-1:0] node15911;
	wire [4-1:0] node15912;
	wire [4-1:0] node15916;
	wire [4-1:0] node15917;
	wire [4-1:0] node15918;
	wire [4-1:0] node15919;
	wire [4-1:0] node15920;
	wire [4-1:0] node15921;
	wire [4-1:0] node15925;
	wire [4-1:0] node15928;
	wire [4-1:0] node15929;
	wire [4-1:0] node15931;
	wire [4-1:0] node15934;
	wire [4-1:0] node15935;
	wire [4-1:0] node15939;
	wire [4-1:0] node15940;
	wire [4-1:0] node15942;
	wire [4-1:0] node15945;
	wire [4-1:0] node15946;
	wire [4-1:0] node15948;
	wire [4-1:0] node15952;
	wire [4-1:0] node15954;
	wire [4-1:0] node15955;
	wire [4-1:0] node15956;
	wire [4-1:0] node15959;
	wire [4-1:0] node15962;
	wire [4-1:0] node15964;
	wire [4-1:0] node15966;
	wire [4-1:0] node15969;
	wire [4-1:0] node15970;
	wire [4-1:0] node15971;
	wire [4-1:0] node15972;
	wire [4-1:0] node15973;
	wire [4-1:0] node15974;
	wire [4-1:0] node15975;
	wire [4-1:0] node15976;
	wire [4-1:0] node15979;
	wire [4-1:0] node15980;
	wire [4-1:0] node15984;
	wire [4-1:0] node15985;
	wire [4-1:0] node15987;
	wire [4-1:0] node15990;
	wire [4-1:0] node15993;
	wire [4-1:0] node15994;
	wire [4-1:0] node15995;
	wire [4-1:0] node15998;
	wire [4-1:0] node16001;
	wire [4-1:0] node16003;
	wire [4-1:0] node16004;
	wire [4-1:0] node16006;
	wire [4-1:0] node16010;
	wire [4-1:0] node16011;
	wire [4-1:0] node16012;
	wire [4-1:0] node16013;
	wire [4-1:0] node16014;
	wire [4-1:0] node16018;
	wire [4-1:0] node16020;
	wire [4-1:0] node16023;
	wire [4-1:0] node16025;
	wire [4-1:0] node16027;
	wire [4-1:0] node16030;
	wire [4-1:0] node16031;
	wire [4-1:0] node16032;
	wire [4-1:0] node16033;
	wire [4-1:0] node16036;
	wire [4-1:0] node16039;
	wire [4-1:0] node16041;
	wire [4-1:0] node16044;
	wire [4-1:0] node16045;
	wire [4-1:0] node16048;
	wire [4-1:0] node16049;
	wire [4-1:0] node16052;
	wire [4-1:0] node16055;
	wire [4-1:0] node16056;
	wire [4-1:0] node16057;
	wire [4-1:0] node16058;
	wire [4-1:0] node16059;
	wire [4-1:0] node16060;
	wire [4-1:0] node16063;
	wire [4-1:0] node16064;
	wire [4-1:0] node16068;
	wire [4-1:0] node16071;
	wire [4-1:0] node16072;
	wire [4-1:0] node16075;
	wire [4-1:0] node16076;
	wire [4-1:0] node16079;
	wire [4-1:0] node16081;
	wire [4-1:0] node16084;
	wire [4-1:0] node16085;
	wire [4-1:0] node16087;
	wire [4-1:0] node16088;
	wire [4-1:0] node16089;
	wire [4-1:0] node16094;
	wire [4-1:0] node16095;
	wire [4-1:0] node16097;
	wire [4-1:0] node16101;
	wire [4-1:0] node16102;
	wire [4-1:0] node16103;
	wire [4-1:0] node16104;
	wire [4-1:0] node16105;
	wire [4-1:0] node16109;
	wire [4-1:0] node16112;
	wire [4-1:0] node16113;
	wire [4-1:0] node16116;
	wire [4-1:0] node16118;
	wire [4-1:0] node16121;
	wire [4-1:0] node16122;
	wire [4-1:0] node16123;
	wire [4-1:0] node16124;
	wire [4-1:0] node16125;
	wire [4-1:0] node16130;
	wire [4-1:0] node16131;
	wire [4-1:0] node16135;
	wire [4-1:0] node16136;
	wire [4-1:0] node16138;
	wire [4-1:0] node16141;
	wire [4-1:0] node16143;
	wire [4-1:0] node16146;
	wire [4-1:0] node16147;
	wire [4-1:0] node16148;
	wire [4-1:0] node16149;
	wire [4-1:0] node16150;
	wire [4-1:0] node16151;
	wire [4-1:0] node16152;
	wire [4-1:0] node16156;
	wire [4-1:0] node16159;
	wire [4-1:0] node16161;
	wire [4-1:0] node16164;
	wire [4-1:0] node16165;
	wire [4-1:0] node16166;
	wire [4-1:0] node16167;
	wire [4-1:0] node16172;
	wire [4-1:0] node16173;
	wire [4-1:0] node16174;
	wire [4-1:0] node16177;
	wire [4-1:0] node16180;
	wire [4-1:0] node16181;
	wire [4-1:0] node16184;
	wire [4-1:0] node16187;
	wire [4-1:0] node16188;
	wire [4-1:0] node16189;
	wire [4-1:0] node16190;
	wire [4-1:0] node16193;
	wire [4-1:0] node16196;
	wire [4-1:0] node16199;
	wire [4-1:0] node16200;
	wire [4-1:0] node16202;
	wire [4-1:0] node16204;
	wire [4-1:0] node16207;
	wire [4-1:0] node16208;
	wire [4-1:0] node16209;
	wire [4-1:0] node16212;
	wire [4-1:0] node16216;
	wire [4-1:0] node16217;
	wire [4-1:0] node16218;
	wire [4-1:0] node16219;
	wire [4-1:0] node16221;
	wire [4-1:0] node16224;
	wire [4-1:0] node16226;
	wire [4-1:0] node16227;
	wire [4-1:0] node16230;
	wire [4-1:0] node16233;
	wire [4-1:0] node16234;
	wire [4-1:0] node16235;
	wire [4-1:0] node16238;
	wire [4-1:0] node16240;
	wire [4-1:0] node16244;
	wire [4-1:0] node16245;
	wire [4-1:0] node16246;
	wire [4-1:0] node16247;
	wire [4-1:0] node16249;
	wire [4-1:0] node16253;
	wire [4-1:0] node16257;
	wire [4-1:0] node16258;
	wire [4-1:0] node16259;
	wire [4-1:0] node16260;
	wire [4-1:0] node16261;
	wire [4-1:0] node16262;
	wire [4-1:0] node16263;
	wire [4-1:0] node16265;
	wire [4-1:0] node16268;
	wire [4-1:0] node16269;
	wire [4-1:0] node16272;
	wire [4-1:0] node16275;
	wire [4-1:0] node16276;
	wire [4-1:0] node16278;
	wire [4-1:0] node16281;
	wire [4-1:0] node16284;
	wire [4-1:0] node16285;
	wire [4-1:0] node16286;
	wire [4-1:0] node16287;
	wire [4-1:0] node16291;
	wire [4-1:0] node16294;
	wire [4-1:0] node16295;
	wire [4-1:0] node16297;
	wire [4-1:0] node16300;
	wire [4-1:0] node16301;
	wire [4-1:0] node16305;
	wire [4-1:0] node16306;
	wire [4-1:0] node16307;
	wire [4-1:0] node16308;
	wire [4-1:0] node16311;
	wire [4-1:0] node16312;
	wire [4-1:0] node16315;
	wire [4-1:0] node16316;
	wire [4-1:0] node16320;
	wire [4-1:0] node16321;
	wire [4-1:0] node16325;
	wire [4-1:0] node16326;
	wire [4-1:0] node16327;
	wire [4-1:0] node16328;
	wire [4-1:0] node16331;
	wire [4-1:0] node16333;
	wire [4-1:0] node16337;
	wire [4-1:0] node16338;
	wire [4-1:0] node16339;
	wire [4-1:0] node16340;
	wire [4-1:0] node16343;
	wire [4-1:0] node16347;
	wire [4-1:0] node16348;
	wire [4-1:0] node16352;
	wire [4-1:0] node16353;
	wire [4-1:0] node16354;
	wire [4-1:0] node16355;
	wire [4-1:0] node16356;
	wire [4-1:0] node16359;
	wire [4-1:0] node16361;
	wire [4-1:0] node16364;
	wire [4-1:0] node16366;
	wire [4-1:0] node16367;
	wire [4-1:0] node16371;
	wire [4-1:0] node16372;
	wire [4-1:0] node16373;
	wire [4-1:0] node16375;
	wire [4-1:0] node16376;
	wire [4-1:0] node16379;
	wire [4-1:0] node16382;
	wire [4-1:0] node16384;
	wire [4-1:0] node16387;
	wire [4-1:0] node16388;
	wire [4-1:0] node16390;
	wire [4-1:0] node16393;
	wire [4-1:0] node16395;
	wire [4-1:0] node16398;
	wire [4-1:0] node16399;
	wire [4-1:0] node16400;
	wire [4-1:0] node16401;
	wire [4-1:0] node16403;
	wire [4-1:0] node16406;
	wire [4-1:0] node16407;
	wire [4-1:0] node16408;
	wire [4-1:0] node16413;
	wire [4-1:0] node16415;
	wire [4-1:0] node16416;
	wire [4-1:0] node16417;
	wire [4-1:0] node16420;
	wire [4-1:0] node16425;
	wire [4-1:0] node16426;
	wire [4-1:0] node16427;
	wire [4-1:0] node16428;
	wire [4-1:0] node16430;
	wire [4-1:0] node16432;
	wire [4-1:0] node16434;
	wire [4-1:0] node16437;
	wire [4-1:0] node16438;
	wire [4-1:0] node16439;
	wire [4-1:0] node16442;
	wire [4-1:0] node16443;
	wire [4-1:0] node16447;
	wire [4-1:0] node16448;
	wire [4-1:0] node16450;
	wire [4-1:0] node16454;
	wire [4-1:0] node16455;
	wire [4-1:0] node16456;
	wire [4-1:0] node16458;
	wire [4-1:0] node16461;
	wire [4-1:0] node16462;
	wire [4-1:0] node16464;
	wire [4-1:0] node16467;
	wire [4-1:0] node16468;
	wire [4-1:0] node16469;
	wire [4-1:0] node16473;
	wire [4-1:0] node16477;
	wire [4-1:0] node16478;
	wire [4-1:0] node16479;
	wire [4-1:0] node16480;
	wire [4-1:0] node16481;
	wire [4-1:0] node16484;
	wire [4-1:0] node16487;
	wire [4-1:0] node16489;
	wire [4-1:0] node16490;
	wire [4-1:0] node16493;
	wire [4-1:0] node16498;
	wire [4-1:0] node16499;
	wire [4-1:0] node16500;
	wire [4-1:0] node16501;
	wire [4-1:0] node16502;
	wire [4-1:0] node16504;
	wire [4-1:0] node16505;
	wire [4-1:0] node16506;
	wire [4-1:0] node16508;
	wire [4-1:0] node16509;
	wire [4-1:0] node16510;
	wire [4-1:0] node16512;
	wire [4-1:0] node16514;
	wire [4-1:0] node16518;
	wire [4-1:0] node16519;
	wire [4-1:0] node16523;
	wire [4-1:0] node16524;
	wire [4-1:0] node16525;
	wire [4-1:0] node16526;
	wire [4-1:0] node16529;
	wire [4-1:0] node16532;
	wire [4-1:0] node16533;
	wire [4-1:0] node16534;
	wire [4-1:0] node16535;
	wire [4-1:0] node16539;
	wire [4-1:0] node16542;
	wire [4-1:0] node16545;
	wire [4-1:0] node16546;
	wire [4-1:0] node16547;
	wire [4-1:0] node16549;
	wire [4-1:0] node16552;
	wire [4-1:0] node16554;
	wire [4-1:0] node16557;
	wire [4-1:0] node16558;
	wire [4-1:0] node16559;
	wire [4-1:0] node16560;
	wire [4-1:0] node16563;
	wire [4-1:0] node16568;
	wire [4-1:0] node16570;
	wire [4-1:0] node16572;
	wire [4-1:0] node16574;
	wire [4-1:0] node16575;
	wire [4-1:0] node16576;
	wire [4-1:0] node16580;
	wire [4-1:0] node16582;
	wire [4-1:0] node16586;
	wire [4-1:0] node16587;
	wire [4-1:0] node16588;
	wire [4-1:0] node16589;
	wire [4-1:0] node16590;
	wire [4-1:0] node16591;
	wire [4-1:0] node16592;
	wire [4-1:0] node16593;
	wire [4-1:0] node16597;
	wire [4-1:0] node16598;
	wire [4-1:0] node16602;
	wire [4-1:0] node16603;
	wire [4-1:0] node16605;
	wire [4-1:0] node16607;
	wire [4-1:0] node16610;
	wire [4-1:0] node16611;
	wire [4-1:0] node16613;
	wire [4-1:0] node16617;
	wire [4-1:0] node16618;
	wire [4-1:0] node16619;
	wire [4-1:0] node16620;
	wire [4-1:0] node16622;
	wire [4-1:0] node16625;
	wire [4-1:0] node16628;
	wire [4-1:0] node16629;
	wire [4-1:0] node16630;
	wire [4-1:0] node16635;
	wire [4-1:0] node16636;
	wire [4-1:0] node16639;
	wire [4-1:0] node16641;
	wire [4-1:0] node16644;
	wire [4-1:0] node16645;
	wire [4-1:0] node16646;
	wire [4-1:0] node16647;
	wire [4-1:0] node16648;
	wire [4-1:0] node16649;
	wire [4-1:0] node16653;
	wire [4-1:0] node16655;
	wire [4-1:0] node16658;
	wire [4-1:0] node16659;
	wire [4-1:0] node16660;
	wire [4-1:0] node16665;
	wire [4-1:0] node16666;
	wire [4-1:0] node16667;
	wire [4-1:0] node16669;
	wire [4-1:0] node16672;
	wire [4-1:0] node16675;
	wire [4-1:0] node16676;
	wire [4-1:0] node16677;
	wire [4-1:0] node16680;
	wire [4-1:0] node16681;
	wire [4-1:0] node16686;
	wire [4-1:0] node16687;
	wire [4-1:0] node16688;
	wire [4-1:0] node16689;
	wire [4-1:0] node16693;
	wire [4-1:0] node16696;
	wire [4-1:0] node16697;
	wire [4-1:0] node16698;
	wire [4-1:0] node16701;
	wire [4-1:0] node16702;
	wire [4-1:0] node16706;
	wire [4-1:0] node16708;
	wire [4-1:0] node16711;
	wire [4-1:0] node16712;
	wire [4-1:0] node16713;
	wire [4-1:0] node16714;
	wire [4-1:0] node16715;
	wire [4-1:0] node16716;
	wire [4-1:0] node16720;
	wire [4-1:0] node16722;
	wire [4-1:0] node16725;
	wire [4-1:0] node16726;
	wire [4-1:0] node16727;
	wire [4-1:0] node16729;
	wire [4-1:0] node16732;
	wire [4-1:0] node16734;
	wire [4-1:0] node16737;
	wire [4-1:0] node16738;
	wire [4-1:0] node16739;
	wire [4-1:0] node16744;
	wire [4-1:0] node16745;
	wire [4-1:0] node16746;
	wire [4-1:0] node16747;
	wire [4-1:0] node16751;
	wire [4-1:0] node16752;
	wire [4-1:0] node16756;
	wire [4-1:0] node16757;
	wire [4-1:0] node16759;
	wire [4-1:0] node16762;
	wire [4-1:0] node16763;
	wire [4-1:0] node16764;
	wire [4-1:0] node16769;
	wire [4-1:0] node16770;
	wire [4-1:0] node16771;
	wire [4-1:0] node16772;
	wire [4-1:0] node16773;
	wire [4-1:0] node16775;
	wire [4-1:0] node16778;
	wire [4-1:0] node16779;
	wire [4-1:0] node16783;
	wire [4-1:0] node16784;
	wire [4-1:0] node16787;
	wire [4-1:0] node16788;
	wire [4-1:0] node16792;
	wire [4-1:0] node16794;
	wire [4-1:0] node16795;
	wire [4-1:0] node16797;
	wire [4-1:0] node16800;
	wire [4-1:0] node16801;
	wire [4-1:0] node16805;
	wire [4-1:0] node16806;
	wire [4-1:0] node16807;
	wire [4-1:0] node16810;
	wire [4-1:0] node16811;
	wire [4-1:0] node16814;
	wire [4-1:0] node16816;
	wire [4-1:0] node16819;
	wire [4-1:0] node16820;
	wire [4-1:0] node16821;
	wire [4-1:0] node16823;
	wire [4-1:0] node16827;
	wire [4-1:0] node16828;
	wire [4-1:0] node16830;
	wire [4-1:0] node16834;
	wire [4-1:0] node16836;
	wire [4-1:0] node16837;
	wire [4-1:0] node16838;
	wire [4-1:0] node16840;
	wire [4-1:0] node16841;
	wire [4-1:0] node16842;
	wire [4-1:0] node16845;
	wire [4-1:0] node16846;
	wire [4-1:0] node16850;
	wire [4-1:0] node16852;
	wire [4-1:0] node16856;
	wire [4-1:0] node16857;
	wire [4-1:0] node16858;
	wire [4-1:0] node16859;
	wire [4-1:0] node16860;
	wire [4-1:0] node16863;
	wire [4-1:0] node16864;
	wire [4-1:0] node16866;
	wire [4-1:0] node16869;
	wire [4-1:0] node16872;
	wire [4-1:0] node16873;
	wire [4-1:0] node16874;
	wire [4-1:0] node16878;
	wire [4-1:0] node16881;
	wire [4-1:0] node16882;
	wire [4-1:0] node16884;
	wire [4-1:0] node16885;
	wire [4-1:0] node16889;
	wire [4-1:0] node16891;
	wire [4-1:0] node16892;
	wire [4-1:0] node16894;
	wire [4-1:0] node16898;
	wire [4-1:0] node16900;
	wire [4-1:0] node16901;
	wire [4-1:0] node16902;
	wire [4-1:0] node16903;
	wire [4-1:0] node16906;
	wire [4-1:0] node16910;
	wire [4-1:0] node16911;
	wire [4-1:0] node16913;
	wire [4-1:0] node16917;
	wire [4-1:0] node16918;
	wire [4-1:0] node16919;
	wire [4-1:0] node16920;
	wire [4-1:0] node16921;
	wire [4-1:0] node16922;
	wire [4-1:0] node16923;
	wire [4-1:0] node16924;
	wire [4-1:0] node16925;
	wire [4-1:0] node16929;
	wire [4-1:0] node16930;
	wire [4-1:0] node16934;
	wire [4-1:0] node16935;
	wire [4-1:0] node16937;
	wire [4-1:0] node16938;
	wire [4-1:0] node16941;
	wire [4-1:0] node16943;
	wire [4-1:0] node16947;
	wire [4-1:0] node16948;
	wire [4-1:0] node16949;
	wire [4-1:0] node16951;
	wire [4-1:0] node16954;
	wire [4-1:0] node16956;
	wire [4-1:0] node16959;
	wire [4-1:0] node16960;
	wire [4-1:0] node16961;
	wire [4-1:0] node16963;
	wire [4-1:0] node16966;
	wire [4-1:0] node16968;
	wire [4-1:0] node16971;
	wire [4-1:0] node16972;
	wire [4-1:0] node16975;
	wire [4-1:0] node16978;
	wire [4-1:0] node16979;
	wire [4-1:0] node16980;
	wire [4-1:0] node16981;
	wire [4-1:0] node16983;
	wire [4-1:0] node16986;
	wire [4-1:0] node16989;
	wire [4-1:0] node16990;
	wire [4-1:0] node16991;
	wire [4-1:0] node16995;
	wire [4-1:0] node16996;
	wire [4-1:0] node16997;
	wire [4-1:0] node17000;
	wire [4-1:0] node17003;
	wire [4-1:0] node17006;
	wire [4-1:0] node17007;
	wire [4-1:0] node17009;
	wire [4-1:0] node17012;
	wire [4-1:0] node17014;
	wire [4-1:0] node17017;
	wire [4-1:0] node17018;
	wire [4-1:0] node17019;
	wire [4-1:0] node17020;
	wire [4-1:0] node17021;
	wire [4-1:0] node17022;
	wire [4-1:0] node17025;
	wire [4-1:0] node17028;
	wire [4-1:0] node17029;
	wire [4-1:0] node17033;
	wire [4-1:0] node17034;
	wire [4-1:0] node17035;
	wire [4-1:0] node17036;
	wire [4-1:0] node17040;
	wire [4-1:0] node17041;
	wire [4-1:0] node17044;
	wire [4-1:0] node17046;
	wire [4-1:0] node17049;
	wire [4-1:0] node17050;
	wire [4-1:0] node17051;
	wire [4-1:0] node17056;
	wire [4-1:0] node17057;
	wire [4-1:0] node17058;
	wire [4-1:0] node17061;
	wire [4-1:0] node17062;
	wire [4-1:0] node17066;
	wire [4-1:0] node17067;
	wire [4-1:0] node17068;
	wire [4-1:0] node17069;
	wire [4-1:0] node17073;
	wire [4-1:0] node17076;
	wire [4-1:0] node17077;
	wire [4-1:0] node17079;
	wire [4-1:0] node17082;
	wire [4-1:0] node17085;
	wire [4-1:0] node17086;
	wire [4-1:0] node17087;
	wire [4-1:0] node17088;
	wire [4-1:0] node17091;
	wire [4-1:0] node17093;
	wire [4-1:0] node17096;
	wire [4-1:0] node17097;
	wire [4-1:0] node17098;
	wire [4-1:0] node17099;
	wire [4-1:0] node17100;
	wire [4-1:0] node17104;
	wire [4-1:0] node17107;
	wire [4-1:0] node17108;
	wire [4-1:0] node17111;
	wire [4-1:0] node17114;
	wire [4-1:0] node17115;
	wire [4-1:0] node17116;
	wire [4-1:0] node17119;
	wire [4-1:0] node17122;
	wire [4-1:0] node17123;
	wire [4-1:0] node17124;
	wire [4-1:0] node17127;
	wire [4-1:0] node17130;
	wire [4-1:0] node17131;
	wire [4-1:0] node17135;
	wire [4-1:0] node17136;
	wire [4-1:0] node17137;
	wire [4-1:0] node17138;
	wire [4-1:0] node17141;
	wire [4-1:0] node17144;
	wire [4-1:0] node17145;
	wire [4-1:0] node17146;
	wire [4-1:0] node17149;
	wire [4-1:0] node17153;
	wire [4-1:0] node17154;
	wire [4-1:0] node17155;
	wire [4-1:0] node17157;
	wire [4-1:0] node17161;
	wire [4-1:0] node17162;
	wire [4-1:0] node17164;
	wire [4-1:0] node17167;
	wire [4-1:0] node17169;
	wire [4-1:0] node17172;
	wire [4-1:0] node17173;
	wire [4-1:0] node17174;
	wire [4-1:0] node17175;
	wire [4-1:0] node17176;
	wire [4-1:0] node17177;
	wire [4-1:0] node17179;
	wire [4-1:0] node17180;
	wire [4-1:0] node17183;
	wire [4-1:0] node17186;
	wire [4-1:0] node17187;
	wire [4-1:0] node17189;
	wire [4-1:0] node17192;
	wire [4-1:0] node17193;
	wire [4-1:0] node17197;
	wire [4-1:0] node17198;
	wire [4-1:0] node17200;
	wire [4-1:0] node17203;
	wire [4-1:0] node17204;
	wire [4-1:0] node17207;
	wire [4-1:0] node17210;
	wire [4-1:0] node17211;
	wire [4-1:0] node17212;
	wire [4-1:0] node17214;
	wire [4-1:0] node17216;
	wire [4-1:0] node17219;
	wire [4-1:0] node17220;
	wire [4-1:0] node17222;
	wire [4-1:0] node17223;
	wire [4-1:0] node17226;
	wire [4-1:0] node17230;
	wire [4-1:0] node17231;
	wire [4-1:0] node17232;
	wire [4-1:0] node17233;
	wire [4-1:0] node17238;
	wire [4-1:0] node17239;
	wire [4-1:0] node17242;
	wire [4-1:0] node17244;
	wire [4-1:0] node17247;
	wire [4-1:0] node17248;
	wire [4-1:0] node17249;
	wire [4-1:0] node17250;
	wire [4-1:0] node17251;
	wire [4-1:0] node17255;
	wire [4-1:0] node17256;
	wire [4-1:0] node17257;
	wire [4-1:0] node17260;
	wire [4-1:0] node17264;
	wire [4-1:0] node17265;
	wire [4-1:0] node17266;
	wire [4-1:0] node17270;
	wire [4-1:0] node17271;
	wire [4-1:0] node17274;
	wire [4-1:0] node17276;
	wire [4-1:0] node17279;
	wire [4-1:0] node17280;
	wire [4-1:0] node17281;
	wire [4-1:0] node17282;
	wire [4-1:0] node17286;
	wire [4-1:0] node17287;
	wire [4-1:0] node17290;
	wire [4-1:0] node17291;
	wire [4-1:0] node17293;
	wire [4-1:0] node17297;
	wire [4-1:0] node17298;
	wire [4-1:0] node17299;
	wire [4-1:0] node17301;
	wire [4-1:0] node17304;
	wire [4-1:0] node17307;
	wire [4-1:0] node17308;
	wire [4-1:0] node17309;
	wire [4-1:0] node17313;
	wire [4-1:0] node17316;
	wire [4-1:0] node17317;
	wire [4-1:0] node17318;
	wire [4-1:0] node17319;
	wire [4-1:0] node17320;
	wire [4-1:0] node17321;
	wire [4-1:0] node17324;
	wire [4-1:0] node17327;
	wire [4-1:0] node17329;
	wire [4-1:0] node17331;
	wire [4-1:0] node17334;
	wire [4-1:0] node17335;
	wire [4-1:0] node17336;
	wire [4-1:0] node17339;
	wire [4-1:0] node17340;
	wire [4-1:0] node17344;
	wire [4-1:0] node17345;
	wire [4-1:0] node17348;
	wire [4-1:0] node17349;
	wire [4-1:0] node17353;
	wire [4-1:0] node17354;
	wire [4-1:0] node17355;
	wire [4-1:0] node17356;
	wire [4-1:0] node17358;
	wire [4-1:0] node17359;
	wire [4-1:0] node17364;
	wire [4-1:0] node17365;
	wire [4-1:0] node17367;
	wire [4-1:0] node17370;
	wire [4-1:0] node17373;
	wire [4-1:0] node17374;
	wire [4-1:0] node17376;
	wire [4-1:0] node17379;
	wire [4-1:0] node17381;
	wire [4-1:0] node17383;
	wire [4-1:0] node17386;
	wire [4-1:0] node17387;
	wire [4-1:0] node17388;
	wire [4-1:0] node17389;
	wire [4-1:0] node17390;
	wire [4-1:0] node17394;
	wire [4-1:0] node17396;
	wire [4-1:0] node17399;
	wire [4-1:0] node17400;
	wire [4-1:0] node17402;
	wire [4-1:0] node17403;
	wire [4-1:0] node17406;
	wire [4-1:0] node17409;
	wire [4-1:0] node17411;
	wire [4-1:0] node17414;
	wire [4-1:0] node17415;
	wire [4-1:0] node17416;
	wire [4-1:0] node17418;
	wire [4-1:0] node17421;
	wire [4-1:0] node17424;
	wire [4-1:0] node17425;
	wire [4-1:0] node17429;
	wire [4-1:0] node17430;
	wire [4-1:0] node17431;
	wire [4-1:0] node17432;
	wire [4-1:0] node17433;
	wire [4-1:0] node17434;
	wire [4-1:0] node17435;
	wire [4-1:0] node17436;
	wire [4-1:0] node17439;
	wire [4-1:0] node17442;
	wire [4-1:0] node17443;
	wire [4-1:0] node17444;
	wire [4-1:0] node17447;
	wire [4-1:0] node17450;
	wire [4-1:0] node17451;
	wire [4-1:0] node17455;
	wire [4-1:0] node17456;
	wire [4-1:0] node17457;
	wire [4-1:0] node17461;
	wire [4-1:0] node17462;
	wire [4-1:0] node17463;
	wire [4-1:0] node17466;
	wire [4-1:0] node17469;
	wire [4-1:0] node17472;
	wire [4-1:0] node17473;
	wire [4-1:0] node17474;
	wire [4-1:0] node17475;
	wire [4-1:0] node17477;
	wire [4-1:0] node17480;
	wire [4-1:0] node17481;
	wire [4-1:0] node17485;
	wire [4-1:0] node17486;
	wire [4-1:0] node17487;
	wire [4-1:0] node17491;
	wire [4-1:0] node17492;
	wire [4-1:0] node17495;
	wire [4-1:0] node17496;
	wire [4-1:0] node17500;
	wire [4-1:0] node17501;
	wire [4-1:0] node17502;
	wire [4-1:0] node17506;
	wire [4-1:0] node17508;
	wire [4-1:0] node17509;
	wire [4-1:0] node17512;
	wire [4-1:0] node17515;
	wire [4-1:0] node17516;
	wire [4-1:0] node17517;
	wire [4-1:0] node17518;
	wire [4-1:0] node17519;
	wire [4-1:0] node17521;
	wire [4-1:0] node17524;
	wire [4-1:0] node17525;
	wire [4-1:0] node17529;
	wire [4-1:0] node17530;
	wire [4-1:0] node17532;
	wire [4-1:0] node17535;
	wire [4-1:0] node17538;
	wire [4-1:0] node17539;
	wire [4-1:0] node17540;
	wire [4-1:0] node17541;
	wire [4-1:0] node17544;
	wire [4-1:0] node17547;
	wire [4-1:0] node17550;
	wire [4-1:0] node17551;
	wire [4-1:0] node17552;
	wire [4-1:0] node17554;
	wire [4-1:0] node17558;
	wire [4-1:0] node17559;
	wire [4-1:0] node17561;
	wire [4-1:0] node17564;
	wire [4-1:0] node17565;
	wire [4-1:0] node17569;
	wire [4-1:0] node17570;
	wire [4-1:0] node17571;
	wire [4-1:0] node17573;
	wire [4-1:0] node17576;
	wire [4-1:0] node17577;
	wire [4-1:0] node17581;
	wire [4-1:0] node17582;
	wire [4-1:0] node17584;
	wire [4-1:0] node17585;
	wire [4-1:0] node17586;
	wire [4-1:0] node17591;
	wire [4-1:0] node17592;
	wire [4-1:0] node17593;
	wire [4-1:0] node17596;
	wire [4-1:0] node17599;
	wire [4-1:0] node17600;
	wire [4-1:0] node17604;
	wire [4-1:0] node17605;
	wire [4-1:0] node17606;
	wire [4-1:0] node17607;
	wire [4-1:0] node17608;
	wire [4-1:0] node17609;
	wire [4-1:0] node17612;
	wire [4-1:0] node17614;
	wire [4-1:0] node17616;
	wire [4-1:0] node17619;
	wire [4-1:0] node17620;
	wire [4-1:0] node17621;
	wire [4-1:0] node17622;
	wire [4-1:0] node17627;
	wire [4-1:0] node17630;
	wire [4-1:0] node17631;
	wire [4-1:0] node17632;
	wire [4-1:0] node17633;
	wire [4-1:0] node17636;
	wire [4-1:0] node17639;
	wire [4-1:0] node17642;
	wire [4-1:0] node17643;
	wire [4-1:0] node17644;
	wire [4-1:0] node17648;
	wire [4-1:0] node17649;
	wire [4-1:0] node17653;
	wire [4-1:0] node17654;
	wire [4-1:0] node17655;
	wire [4-1:0] node17656;
	wire [4-1:0] node17659;
	wire [4-1:0] node17661;
	wire [4-1:0] node17664;
	wire [4-1:0] node17665;
	wire [4-1:0] node17666;
	wire [4-1:0] node17669;
	wire [4-1:0] node17672;
	wire [4-1:0] node17673;
	wire [4-1:0] node17674;
	wire [4-1:0] node17679;
	wire [4-1:0] node17680;
	wire [4-1:0] node17681;
	wire [4-1:0] node17684;
	wire [4-1:0] node17687;
	wire [4-1:0] node17688;
	wire [4-1:0] node17690;
	wire [4-1:0] node17691;
	wire [4-1:0] node17695;
	wire [4-1:0] node17697;
	wire [4-1:0] node17698;
	wire [4-1:0] node17701;
	wire [4-1:0] node17704;
	wire [4-1:0] node17705;
	wire [4-1:0] node17706;
	wire [4-1:0] node17707;
	wire [4-1:0] node17708;
	wire [4-1:0] node17710;
	wire [4-1:0] node17714;
	wire [4-1:0] node17715;
	wire [4-1:0] node17718;
	wire [4-1:0] node17721;
	wire [4-1:0] node17722;
	wire [4-1:0] node17723;
	wire [4-1:0] node17727;
	wire [4-1:0] node17729;
	wire [4-1:0] node17732;
	wire [4-1:0] node17733;
	wire [4-1:0] node17734;
	wire [4-1:0] node17735;
	wire [4-1:0] node17738;
	wire [4-1:0] node17741;
	wire [4-1:0] node17742;
	wire [4-1:0] node17743;
	wire [4-1:0] node17747;
	wire [4-1:0] node17750;
	wire [4-1:0] node17752;
	wire [4-1:0] node17754;
	wire [4-1:0] node17757;
	wire [4-1:0] node17758;
	wire [4-1:0] node17759;
	wire [4-1:0] node17760;
	wire [4-1:0] node17761;
	wire [4-1:0] node17762;
	wire [4-1:0] node17763;
	wire [4-1:0] node17764;
	wire [4-1:0] node17769;
	wire [4-1:0] node17772;
	wire [4-1:0] node17773;
	wire [4-1:0] node17774;
	wire [4-1:0] node17775;
	wire [4-1:0] node17778;
	wire [4-1:0] node17782;
	wire [4-1:0] node17784;
	wire [4-1:0] node17787;
	wire [4-1:0] node17788;
	wire [4-1:0] node17789;
	wire [4-1:0] node17791;
	wire [4-1:0] node17794;
	wire [4-1:0] node17795;
	wire [4-1:0] node17797;
	wire [4-1:0] node17800;
	wire [4-1:0] node17801;
	wire [4-1:0] node17804;
	wire [4-1:0] node17807;
	wire [4-1:0] node17808;
	wire [4-1:0] node17809;
	wire [4-1:0] node17811;
	wire [4-1:0] node17812;
	wire [4-1:0] node17816;
	wire [4-1:0] node17817;
	wire [4-1:0] node17818;
	wire [4-1:0] node17821;
	wire [4-1:0] node17825;
	wire [4-1:0] node17826;
	wire [4-1:0] node17827;
	wire [4-1:0] node17831;
	wire [4-1:0] node17834;
	wire [4-1:0] node17835;
	wire [4-1:0] node17836;
	wire [4-1:0] node17837;
	wire [4-1:0] node17838;
	wire [4-1:0] node17839;
	wire [4-1:0] node17842;
	wire [4-1:0] node17846;
	wire [4-1:0] node17847;
	wire [4-1:0] node17848;
	wire [4-1:0] node17852;
	wire [4-1:0] node17853;
	wire [4-1:0] node17854;
	wire [4-1:0] node17858;
	wire [4-1:0] node17860;
	wire [4-1:0] node17863;
	wire [4-1:0] node17864;
	wire [4-1:0] node17867;
	wire [4-1:0] node17868;
	wire [4-1:0] node17869;
	wire [4-1:0] node17873;
	wire [4-1:0] node17876;
	wire [4-1:0] node17877;
	wire [4-1:0] node17878;
	wire [4-1:0] node17879;
	wire [4-1:0] node17882;
	wire [4-1:0] node17885;
	wire [4-1:0] node17886;
	wire [4-1:0] node17889;
	wire [4-1:0] node17890;
	wire [4-1:0] node17894;
	wire [4-1:0] node17895;
	wire [4-1:0] node17897;
	wire [4-1:0] node17901;
	wire [4-1:0] node17902;
	wire [4-1:0] node17903;
	wire [4-1:0] node17904;
	wire [4-1:0] node17905;
	wire [4-1:0] node17906;
	wire [4-1:0] node17907;
	wire [4-1:0] node17911;
	wire [4-1:0] node17913;
	wire [4-1:0] node17916;
	wire [4-1:0] node17917;
	wire [4-1:0] node17918;
	wire [4-1:0] node17921;
	wire [4-1:0] node17924;
	wire [4-1:0] node17925;
	wire [4-1:0] node17928;
	wire [4-1:0] node17931;
	wire [4-1:0] node17932;
	wire [4-1:0] node17933;
	wire [4-1:0] node17934;
	wire [4-1:0] node17938;
	wire [4-1:0] node17939;
	wire [4-1:0] node17942;
	wire [4-1:0] node17945;
	wire [4-1:0] node17948;
	wire [4-1:0] node17949;
	wire [4-1:0] node17950;
	wire [4-1:0] node17951;
	wire [4-1:0] node17953;
	wire [4-1:0] node17957;
	wire [4-1:0] node17958;
	wire [4-1:0] node17959;
	wire [4-1:0] node17963;
	wire [4-1:0] node17966;
	wire [4-1:0] node17967;
	wire [4-1:0] node17968;
	wire [4-1:0] node17969;
	wire [4-1:0] node17972;
	wire [4-1:0] node17977;
	wire [4-1:0] node17978;
	wire [4-1:0] node17979;
	wire [4-1:0] node17980;
	wire [4-1:0] node17981;
	wire [4-1:0] node17983;
	wire [4-1:0] node17987;
	wire [4-1:0] node17988;
	wire [4-1:0] node17992;
	wire [4-1:0] node17993;
	wire [4-1:0] node17994;
	wire [4-1:0] node17996;
	wire [4-1:0] node18001;
	wire [4-1:0] node18002;
	wire [4-1:0] node18003;
	wire [4-1:0] node18005;
	wire [4-1:0] node18010;
	wire [4-1:0] node18012;
	wire [4-1:0] node18013;
	wire [4-1:0] node18014;
	wire [4-1:0] node18016;
	wire [4-1:0] node18017;
	wire [4-1:0] node18018;
	wire [4-1:0] node18020;
	wire [4-1:0] node18021;
	wire [4-1:0] node18022;
	wire [4-1:0] node18027;
	wire [4-1:0] node18028;
	wire [4-1:0] node18029;
	wire [4-1:0] node18031;
	wire [4-1:0] node18032;
	wire [4-1:0] node18033;
	wire [4-1:0] node18037;
	wire [4-1:0] node18040;
	wire [4-1:0] node18042;
	wire [4-1:0] node18044;
	wire [4-1:0] node18047;
	wire [4-1:0] node18048;
	wire [4-1:0] node18049;
	wire [4-1:0] node18052;
	wire [4-1:0] node18053;
	wire [4-1:0] node18057;
	wire [4-1:0] node18059;
	wire [4-1:0] node18063;
	wire [4-1:0] node18064;
	wire [4-1:0] node18065;
	wire [4-1:0] node18066;
	wire [4-1:0] node18067;
	wire [4-1:0] node18069;
	wire [4-1:0] node18070;
	wire [4-1:0] node18073;
	wire [4-1:0] node18074;
	wire [4-1:0] node18075;
	wire [4-1:0] node18080;
	wire [4-1:0] node18081;
	wire [4-1:0] node18082;
	wire [4-1:0] node18085;
	wire [4-1:0] node18086;
	wire [4-1:0] node18090;
	wire [4-1:0] node18091;
	wire [4-1:0] node18094;
	wire [4-1:0] node18097;
	wire [4-1:0] node18098;
	wire [4-1:0] node18099;
	wire [4-1:0] node18100;
	wire [4-1:0] node18101;
	wire [4-1:0] node18106;
	wire [4-1:0] node18107;
	wire [4-1:0] node18108;
	wire [4-1:0] node18111;
	wire [4-1:0] node18114;
	wire [4-1:0] node18117;
	wire [4-1:0] node18118;
	wire [4-1:0] node18119;
	wire [4-1:0] node18123;
	wire [4-1:0] node18124;
	wire [4-1:0] node18127;
	wire [4-1:0] node18129;
	wire [4-1:0] node18130;
	wire [4-1:0] node18134;
	wire [4-1:0] node18135;
	wire [4-1:0] node18136;
	wire [4-1:0] node18137;
	wire [4-1:0] node18138;
	wire [4-1:0] node18142;
	wire [4-1:0] node18143;
	wire [4-1:0] node18144;
	wire [4-1:0] node18146;
	wire [4-1:0] node18151;
	wire [4-1:0] node18152;
	wire [4-1:0] node18153;
	wire [4-1:0] node18154;
	wire [4-1:0] node18157;
	wire [4-1:0] node18160;
	wire [4-1:0] node18161;
	wire [4-1:0] node18164;
	wire [4-1:0] node18166;
	wire [4-1:0] node18169;
	wire [4-1:0] node18170;
	wire [4-1:0] node18172;
	wire [4-1:0] node18173;
	wire [4-1:0] node18178;
	wire [4-1:0] node18179;
	wire [4-1:0] node18180;
	wire [4-1:0] node18181;
	wire [4-1:0] node18182;
	wire [4-1:0] node18185;
	wire [4-1:0] node18188;
	wire [4-1:0] node18191;
	wire [4-1:0] node18192;
	wire [4-1:0] node18193;
	wire [4-1:0] node18194;
	wire [4-1:0] node18199;
	wire [4-1:0] node18202;
	wire [4-1:0] node18203;
	wire [4-1:0] node18204;
	wire [4-1:0] node18205;
	wire [4-1:0] node18210;
	wire [4-1:0] node18212;
	wire [4-1:0] node18213;
	wire [4-1:0] node18217;
	wire [4-1:0] node18218;
	wire [4-1:0] node18219;
	wire [4-1:0] node18220;
	wire [4-1:0] node18221;
	wire [4-1:0] node18223;
	wire [4-1:0] node18224;
	wire [4-1:0] node18226;
	wire [4-1:0] node18230;
	wire [4-1:0] node18231;
	wire [4-1:0] node18234;
	wire [4-1:0] node18236;
	wire [4-1:0] node18237;
	wire [4-1:0] node18241;
	wire [4-1:0] node18242;
	wire [4-1:0] node18243;
	wire [4-1:0] node18247;
	wire [4-1:0] node18248;
	wire [4-1:0] node18250;
	wire [4-1:0] node18252;
	wire [4-1:0] node18256;
	wire [4-1:0] node18257;
	wire [4-1:0] node18258;
	wire [4-1:0] node18259;
	wire [4-1:0] node18262;
	wire [4-1:0] node18265;
	wire [4-1:0] node18267;
	wire [4-1:0] node18268;
	wire [4-1:0] node18272;
	wire [4-1:0] node18273;
	wire [4-1:0] node18274;
	wire [4-1:0] node18277;
	wire [4-1:0] node18280;
	wire [4-1:0] node18281;
	wire [4-1:0] node18283;
	wire [4-1:0] node18284;
	wire [4-1:0] node18288;
	wire [4-1:0] node18291;
	wire [4-1:0] node18292;
	wire [4-1:0] node18293;
	wire [4-1:0] node18294;
	wire [4-1:0] node18295;
	wire [4-1:0] node18297;
	wire [4-1:0] node18300;
	wire [4-1:0] node18303;
	wire [4-1:0] node18305;
	wire [4-1:0] node18308;
	wire [4-1:0] node18309;
	wire [4-1:0] node18310;
	wire [4-1:0] node18314;
	wire [4-1:0] node18315;
	wire [4-1:0] node18316;
	wire [4-1:0] node18319;
	wire [4-1:0] node18323;
	wire [4-1:0] node18324;
	wire [4-1:0] node18325;
	wire [4-1:0] node18328;
	wire [4-1:0] node18330;
	wire [4-1:0] node18331;
	wire [4-1:0] node18335;
	wire [4-1:0] node18336;
	wire [4-1:0] node18337;
	wire [4-1:0] node18342;
	wire [4-1:0] node18344;
	wire [4-1:0] node18346;
	wire [4-1:0] node18347;
	wire [4-1:0] node18348;
	wire [4-1:0] node18350;
	wire [4-1:0] node18352;
	wire [4-1:0] node18354;
	wire [4-1:0] node18356;
	wire [4-1:0] node18359;
	wire [4-1:0] node18360;
	wire [4-1:0] node18361;
	wire [4-1:0] node18362;
	wire [4-1:0] node18363;
	wire [4-1:0] node18367;
	wire [4-1:0] node18368;
	wire [4-1:0] node18372;
	wire [4-1:0] node18373;
	wire [4-1:0] node18376;
	wire [4-1:0] node18379;
	wire [4-1:0] node18380;
	wire [4-1:0] node18381;
	wire [4-1:0] node18382;
	wire [4-1:0] node18385;
	wire [4-1:0] node18390;
	wire [4-1:0] node18391;
	wire [4-1:0] node18393;
	wire [4-1:0] node18395;
	wire [4-1:0] node18396;
	wire [4-1:0] node18398;

	assign outp = (inp[8]) ? node9306 : node1;
		assign node1 = (inp[9]) ? node4667 : node2;
			assign node2 = (inp[6]) ? node1076 : node3;
				assign node3 = (inp[15]) ? node595 : node4;
					assign node4 = (inp[0]) ? 4'b1101 : node5;
						assign node5 = (inp[5]) ? node229 : node6;
							assign node6 = (inp[2]) ? 4'b1111 : node7;
								assign node7 = (inp[3]) ? node99 : node8;
									assign node8 = (inp[4]) ? node36 : node9;
										assign node9 = (inp[7]) ? 4'b1111 : node10;
											assign node10 = (inp[13]) ? node24 : node11;
												assign node11 = (inp[10]) ? node19 : node12;
													assign node12 = (inp[12]) ? 4'b1111 : node13;
														assign node13 = (inp[14]) ? 4'b1111 : node14;
															assign node14 = (inp[1]) ? 4'b0001 : 4'b0000;
													assign node19 = (inp[1]) ? 4'b0001 : node20;
														assign node20 = (inp[14]) ? 4'b0001 : 4'b0000;
												assign node24 = (inp[1]) ? node30 : node25;
													assign node25 = (inp[11]) ? 4'b1000 : node26;
														assign node26 = (inp[14]) ? 4'b1001 : 4'b1000;
													assign node30 = (inp[12]) ? node32 : 4'b1001;
														assign node32 = (inp[11]) ? 4'b0001 : 4'b1000;
										assign node36 = (inp[1]) ? node72 : node37;
											assign node37 = (inp[11]) ? node55 : node38;
												assign node38 = (inp[14]) ? node48 : node39;
													assign node39 = (inp[12]) ? node41 : 4'b0000;
														assign node41 = (inp[7]) ? 4'b0000 : node42;
															assign node42 = (inp[10]) ? node44 : 4'b1000;
																assign node44 = (inp[13]) ? 4'b1000 : 4'b0000;
													assign node48 = (inp[13]) ? 4'b0001 : node49;
														assign node49 = (inp[7]) ? 4'b1111 : node50;
															assign node50 = (inp[10]) ? 4'b0001 : 4'b1001;
												assign node55 = (inp[13]) ? node67 : node56;
													assign node56 = (inp[7]) ? node62 : node57;
														assign node57 = (inp[10]) ? 4'b0000 : node58;
															assign node58 = (inp[14]) ? 4'b1000 : 4'b0000;
														assign node62 = (inp[12]) ? node64 : 4'b0000;
															assign node64 = (inp[10]) ? 4'b0000 : 4'b1111;
													assign node67 = (inp[10]) ? 4'b1000 : node68;
														assign node68 = (inp[12]) ? 4'b0000 : 4'b1000;
											assign node72 = (inp[11]) ? node88 : node73;
												assign node73 = (inp[14]) ? node81 : node74;
													assign node74 = (inp[12]) ? node78 : node75;
														assign node75 = (inp[7]) ? 4'b1001 : 4'b0001;
														assign node78 = (inp[7]) ? 4'b0001 : 4'b1001;
													assign node81 = (inp[13]) ? 4'b1000 : node82;
														assign node82 = (inp[10]) ? 4'b0000 : node83;
															assign node83 = (inp[12]) ? 4'b1000 : 4'b0000;
												assign node88 = (inp[13]) ? node94 : node89;
													assign node89 = (inp[10]) ? 4'b0001 : node90;
														assign node90 = (inp[12]) ? 4'b1111 : 4'b0001;
													assign node94 = (inp[12]) ? node96 : 4'b1001;
														assign node96 = (inp[10]) ? 4'b1001 : 4'b0001;
									assign node99 = (inp[1]) ? node169 : node100;
										assign node100 = (inp[7]) ? node134 : node101;
											assign node101 = (inp[11]) ? node121 : node102;
												assign node102 = (inp[14]) ? node110 : node103;
													assign node103 = (inp[12]) ? node107 : node104;
														assign node104 = (inp[13]) ? 4'b1100 : 4'b0100;
														assign node107 = (inp[4]) ? 4'b1100 : 4'b1000;
													assign node110 = (inp[4]) ? node116 : node111;
														assign node111 = (inp[13]) ? 4'b0101 : node112;
															assign node112 = (inp[10]) ? 4'b0101 : 4'b1001;
														assign node116 = (inp[12]) ? 4'b1101 : node117;
															assign node117 = (inp[13]) ? 4'b1101 : 4'b0101;
												assign node121 = (inp[13]) ? node129 : node122;
													assign node122 = (inp[12]) ? node124 : 4'b0100;
														assign node124 = (inp[10]) ? 4'b0100 : node125;
															assign node125 = (inp[4]) ? 4'b1100 : 4'b1000;
													assign node129 = (inp[10]) ? 4'b1100 : node130;
														assign node130 = (inp[12]) ? 4'b0100 : 4'b1100;
											assign node134 = (inp[4]) ? node156 : node135;
												assign node135 = (inp[11]) ? node145 : node136;
													assign node136 = (inp[14]) ? node142 : node137;
														assign node137 = (inp[10]) ? node139 : 4'b0000;
															assign node139 = (inp[13]) ? 4'b1000 : 4'b0000;
														assign node142 = (inp[12]) ? 4'b0001 : 4'b1001;
													assign node145 = (inp[13]) ? node151 : node146;
														assign node146 = (inp[12]) ? node148 : 4'b0000;
															assign node148 = (inp[10]) ? 4'b0000 : 4'b1000;
														assign node151 = (inp[10]) ? 4'b1000 : node152;
															assign node152 = (inp[12]) ? 4'b0000 : 4'b1000;
												assign node156 = (inp[14]) ? node160 : node157;
													assign node157 = (inp[13]) ? 4'b1100 : 4'b0100;
													assign node160 = (inp[11]) ? node166 : node161;
														assign node161 = (inp[13]) ? 4'b0101 : node162;
															assign node162 = (inp[10]) ? 4'b0101 : 4'b1001;
														assign node166 = (inp[10]) ? 4'b0100 : 4'b1000;
										assign node169 = (inp[13]) ? node203 : node170;
											assign node170 = (inp[10]) ? node186 : node171;
												assign node171 = (inp[12]) ? node179 : node172;
													assign node172 = (inp[4]) ? 4'b0101 : node173;
														assign node173 = (inp[7]) ? 4'b0001 : node174;
															assign node174 = (inp[14]) ? 4'b0100 : 4'b0101;
													assign node179 = (inp[4]) ? node181 : 4'b1001;
														assign node181 = (inp[7]) ? 4'b1001 : node182;
															assign node182 = (inp[11]) ? 4'b1101 : 4'b1100;
												assign node186 = (inp[11]) ? node198 : node187;
													assign node187 = (inp[14]) ? node193 : node188;
														assign node188 = (inp[7]) ? node190 : 4'b0101;
															assign node190 = (inp[4]) ? 4'b0101 : 4'b0001;
														assign node193 = (inp[4]) ? 4'b0100 : node194;
															assign node194 = (inp[12]) ? 4'b0100 : 4'b0000;
													assign node198 = (inp[4]) ? 4'b0101 : node199;
														assign node199 = (inp[7]) ? 4'b0001 : 4'b0101;
											assign node203 = (inp[10]) ? node219 : node204;
												assign node204 = (inp[12]) ? node212 : node205;
													assign node205 = (inp[14]) ? node209 : node206;
														assign node206 = (inp[7]) ? 4'b1001 : 4'b1101;
														assign node209 = (inp[11]) ? 4'b1101 : 4'b1100;
													assign node212 = (inp[11]) ? node216 : node213;
														assign node213 = (inp[14]) ? 4'b0100 : 4'b0001;
														assign node216 = (inp[4]) ? 4'b0101 : 4'b0001;
												assign node219 = (inp[4]) ? node223 : node220;
													assign node220 = (inp[11]) ? 4'b1001 : 4'b1101;
													assign node223 = (inp[14]) ? node225 : 4'b1101;
														assign node225 = (inp[11]) ? 4'b1101 : 4'b1100;
							assign node229 = (inp[1]) ? node415 : node230;
								assign node230 = (inp[14]) ? node304 : node231;
									assign node231 = (inp[13]) ? node275 : node232;
										assign node232 = (inp[12]) ? node246 : node233;
											assign node233 = (inp[3]) ? node241 : node234;
												assign node234 = (inp[4]) ? 4'b0000 : node235;
													assign node235 = (inp[7]) ? node237 : 4'b0000;
														assign node237 = (inp[2]) ? 4'b1111 : 4'b0100;
												assign node241 = (inp[7]) ? node243 : 4'b0100;
													assign node243 = (inp[4]) ? 4'b0100 : 4'b0000;
											assign node246 = (inp[10]) ? node264 : node247;
												assign node247 = (inp[3]) ? node259 : node248;
													assign node248 = (inp[2]) ? node254 : node249;
														assign node249 = (inp[11]) ? node251 : 4'b1100;
															assign node251 = (inp[4]) ? 4'b1000 : 4'b1100;
														assign node254 = (inp[4]) ? node256 : 4'b1111;
															assign node256 = (inp[7]) ? 4'b1111 : 4'b1000;
													assign node259 = (inp[7]) ? 4'b1000 : node260;
														assign node260 = (inp[4]) ? 4'b1100 : 4'b1000;
												assign node264 = (inp[3]) ? node272 : node265;
													assign node265 = (inp[4]) ? 4'b0000 : node266;
														assign node266 = (inp[7]) ? node268 : 4'b0000;
															assign node268 = (inp[2]) ? 4'b1111 : 4'b0100;
													assign node272 = (inp[2]) ? 4'b0100 : 4'b0000;
										assign node275 = (inp[3]) ? node291 : node276;
											assign node276 = (inp[7]) ? node282 : node277;
												assign node277 = (inp[12]) ? node279 : 4'b1000;
													assign node279 = (inp[10]) ? 4'b1000 : 4'b0000;
												assign node282 = (inp[4]) ? node286 : node283;
													assign node283 = (inp[2]) ? 4'b1111 : 4'b1100;
													assign node286 = (inp[10]) ? 4'b1000 : node287;
														assign node287 = (inp[12]) ? 4'b0000 : 4'b1000;
											assign node291 = (inp[4]) ? node299 : node292;
												assign node292 = (inp[7]) ? node294 : 4'b1100;
													assign node294 = (inp[10]) ? 4'b1000 : node295;
														assign node295 = (inp[12]) ? 4'b0000 : 4'b1000;
												assign node299 = (inp[10]) ? 4'b1100 : node300;
													assign node300 = (inp[12]) ? 4'b0100 : 4'b1100;
									assign node304 = (inp[11]) ? node364 : node305;
										assign node305 = (inp[13]) ? node337 : node306;
											assign node306 = (inp[12]) ? node326 : node307;
												assign node307 = (inp[10]) ? node317 : node308;
													assign node308 = (inp[3]) ? node314 : node309;
														assign node309 = (inp[2]) ? node311 : 4'b1101;
															assign node311 = (inp[4]) ? 4'b1001 : 4'b1111;
														assign node314 = (inp[7]) ? 4'b1001 : 4'b1101;
													assign node317 = (inp[3]) ? node321 : node318;
														assign node318 = (inp[7]) ? 4'b0101 : 4'b0001;
														assign node321 = (inp[7]) ? node323 : 4'b0101;
															assign node323 = (inp[4]) ? 4'b0101 : 4'b0001;
												assign node326 = (inp[3]) ? node332 : node327;
													assign node327 = (inp[4]) ? 4'b1001 : node328;
														assign node328 = (inp[2]) ? 4'b1111 : 4'b1101;
													assign node332 = (inp[7]) ? 4'b1001 : node333;
														assign node333 = (inp[4]) ? 4'b1101 : 4'b1001;
											assign node337 = (inp[12]) ? node351 : node338;
												assign node338 = (inp[10]) ? node346 : node339;
													assign node339 = (inp[3]) ? node343 : node340;
														assign node340 = (inp[4]) ? 4'b0001 : 4'b1111;
														assign node343 = (inp[4]) ? 4'b0101 : 4'b0001;
													assign node346 = (inp[3]) ? 4'b1101 : node347;
														assign node347 = (inp[4]) ? 4'b1001 : 4'b1111;
												assign node351 = (inp[3]) ? node359 : node352;
													assign node352 = (inp[4]) ? 4'b0001 : node353;
														assign node353 = (inp[7]) ? node355 : 4'b0001;
															assign node355 = (inp[2]) ? 4'b1111 : 4'b0101;
													assign node359 = (inp[7]) ? node361 : 4'b0101;
														assign node361 = (inp[4]) ? 4'b0101 : 4'b0001;
										assign node364 = (inp[3]) ? node392 : node365;
											assign node365 = (inp[4]) ? node383 : node366;
												assign node366 = (inp[7]) ? node380 : node367;
													assign node367 = (inp[12]) ? node371 : node368;
														assign node368 = (inp[13]) ? 4'b1000 : 4'b0000;
														assign node371 = (inp[13]) ? node377 : node372;
															assign node372 = (inp[10]) ? 4'b0000 : node373;
																assign node373 = (inp[2]) ? 4'b1111 : 4'b1100;
															assign node377 = (inp[10]) ? 4'b1000 : 4'b0000;
													assign node380 = (inp[2]) ? 4'b1111 : 4'b0100;
												assign node383 = (inp[13]) ? node389 : node384;
													assign node384 = (inp[10]) ? 4'b0000 : node385;
														assign node385 = (inp[12]) ? 4'b1000 : 4'b0000;
													assign node389 = (inp[10]) ? 4'b1000 : 4'b0000;
											assign node392 = (inp[13]) ? node406 : node393;
												assign node393 = (inp[7]) ? node399 : node394;
													assign node394 = (inp[10]) ? 4'b0100 : node395;
														assign node395 = (inp[12]) ? 4'b1100 : 4'b0100;
													assign node399 = (inp[4]) ? node401 : 4'b0000;
														assign node401 = (inp[10]) ? 4'b0100 : node402;
															assign node402 = (inp[12]) ? 4'b1000 : 4'b0100;
												assign node406 = (inp[12]) ? node412 : node407;
													assign node407 = (inp[4]) ? 4'b1100 : node408;
														assign node408 = (inp[7]) ? 4'b1000 : 4'b1100;
													assign node412 = (inp[7]) ? 4'b1100 : 4'b0100;
								assign node415 = (inp[13]) ? node499 : node416;
									assign node416 = (inp[10]) ? node468 : node417;
										assign node417 = (inp[12]) ? node441 : node418;
											assign node418 = (inp[3]) ? node434 : node419;
												assign node419 = (inp[11]) ? node427 : node420;
													assign node420 = (inp[14]) ? node422 : 4'b0001;
														assign node422 = (inp[7]) ? node424 : 4'b0000;
															assign node424 = (inp[4]) ? 4'b0000 : 4'b0100;
													assign node427 = (inp[4]) ? 4'b0001 : node428;
														assign node428 = (inp[7]) ? node430 : 4'b0001;
															assign node430 = (inp[2]) ? 4'b1111 : 4'b0101;
												assign node434 = (inp[11]) ? node438 : node435;
													assign node435 = (inp[14]) ? 4'b0100 : 4'b0101;
													assign node438 = (inp[4]) ? 4'b0101 : 4'b0001;
											assign node441 = (inp[3]) ? node459 : node442;
												assign node442 = (inp[2]) ? node454 : node443;
													assign node443 = (inp[14]) ? node449 : node444;
														assign node444 = (inp[11]) ? node446 : 4'b1101;
															assign node446 = (inp[4]) ? 4'b1001 : 4'b1101;
														assign node449 = (inp[11]) ? 4'b1101 : node450;
															assign node450 = (inp[7]) ? 4'b1100 : 4'b1000;
													assign node454 = (inp[4]) ? node456 : 4'b1111;
														assign node456 = (inp[7]) ? 4'b1111 : 4'b1001;
												assign node459 = (inp[7]) ? node463 : node460;
													assign node460 = (inp[4]) ? 4'b1101 : 4'b1001;
													assign node463 = (inp[14]) ? node465 : 4'b1001;
														assign node465 = (inp[11]) ? 4'b1001 : 4'b1000;
										assign node468 = (inp[3]) ? node484 : node469;
											assign node469 = (inp[14]) ? node477 : node470;
												assign node470 = (inp[7]) ? node472 : 4'b0001;
													assign node472 = (inp[4]) ? 4'b0001 : node473;
														assign node473 = (inp[2]) ? 4'b1111 : 4'b0101;
												assign node477 = (inp[11]) ? node479 : 4'b0000;
													assign node479 = (inp[4]) ? 4'b0001 : node480;
														assign node480 = (inp[7]) ? 4'b0101 : 4'b0001;
											assign node484 = (inp[7]) ? node490 : node485;
												assign node485 = (inp[11]) ? 4'b0101 : node486;
													assign node486 = (inp[14]) ? 4'b0100 : 4'b0101;
												assign node490 = (inp[4]) ? node496 : node491;
													assign node491 = (inp[14]) ? node493 : 4'b0001;
														assign node493 = (inp[11]) ? 4'b0001 : 4'b0000;
													assign node496 = (inp[14]) ? 4'b0100 : 4'b0101;
									assign node499 = (inp[14]) ? node537 : node500;
										assign node500 = (inp[12]) ? node514 : node501;
											assign node501 = (inp[3]) ? node509 : node502;
												assign node502 = (inp[4]) ? 4'b1001 : node503;
													assign node503 = (inp[7]) ? node505 : 4'b1001;
														assign node505 = (inp[2]) ? 4'b1111 : 4'b1101;
												assign node509 = (inp[4]) ? 4'b1101 : node510;
													assign node510 = (inp[7]) ? 4'b1001 : 4'b1101;
											assign node514 = (inp[10]) ? node526 : node515;
												assign node515 = (inp[3]) ? node521 : node516;
													assign node516 = (inp[4]) ? 4'b0001 : node517;
														assign node517 = (inp[7]) ? 4'b1111 : 4'b0001;
													assign node521 = (inp[7]) ? node523 : 4'b0101;
														assign node523 = (inp[4]) ? 4'b0101 : 4'b0001;
												assign node526 = (inp[3]) ? node532 : node527;
													assign node527 = (inp[7]) ? node529 : 4'b1001;
														assign node529 = (inp[4]) ? 4'b1001 : 4'b1101;
													assign node532 = (inp[7]) ? node534 : 4'b1101;
														assign node534 = (inp[2]) ? 4'b1101 : 4'b1001;
										assign node537 = (inp[11]) ? node563 : node538;
											assign node538 = (inp[3]) ? node552 : node539;
												assign node539 = (inp[7]) ? node545 : node540;
													assign node540 = (inp[10]) ? 4'b1000 : node541;
														assign node541 = (inp[12]) ? 4'b0000 : 4'b1000;
													assign node545 = (inp[4]) ? 4'b1000 : node546;
														assign node546 = (inp[2]) ? 4'b1111 : node547;
															assign node547 = (inp[10]) ? 4'b1100 : 4'b0100;
												assign node552 = (inp[7]) ? node554 : 4'b1100;
													assign node554 = (inp[4]) ? node558 : node555;
														assign node555 = (inp[10]) ? 4'b1000 : 4'b0000;
														assign node558 = (inp[10]) ? 4'b1100 : node559;
															assign node559 = (inp[12]) ? 4'b0100 : 4'b1100;
											assign node563 = (inp[12]) ? node575 : node564;
												assign node564 = (inp[3]) ? node570 : node565;
													assign node565 = (inp[7]) ? node567 : 4'b1001;
														assign node567 = (inp[4]) ? 4'b1001 : 4'b1111;
													assign node570 = (inp[4]) ? 4'b1101 : node571;
														assign node571 = (inp[7]) ? 4'b1001 : 4'b1101;
												assign node575 = (inp[10]) ? node585 : node576;
													assign node576 = (inp[7]) ? node580 : node577;
														assign node577 = (inp[3]) ? 4'b0101 : 4'b0001;
														assign node580 = (inp[3]) ? 4'b0001 : node581;
															assign node581 = (inp[4]) ? 4'b0001 : 4'b0101;
													assign node585 = (inp[3]) ? 4'b1101 : node586;
														assign node586 = (inp[7]) ? node588 : 4'b1001;
															assign node588 = (inp[4]) ? 4'b1001 : node589;
																assign node589 = (inp[2]) ? 4'b1111 : 4'b1101;
					assign node595 = (inp[0]) ? 4'b1001 : node596;
						assign node596 = (inp[5]) ? node704 : node597;
							assign node597 = (inp[3]) ? node599 : 4'b1011;
								assign node599 = (inp[2]) ? 4'b1011 : node600;
									assign node600 = (inp[4]) ? node636 : node601;
										assign node601 = (inp[7]) ? 4'b1011 : node602;
											assign node602 = (inp[13]) ? node620 : node603;
												assign node603 = (inp[12]) ? node611 : node604;
													assign node604 = (inp[1]) ? node606 : 4'b0000;
														assign node606 = (inp[14]) ? node608 : 4'b0001;
															assign node608 = (inp[11]) ? 4'b0001 : 4'b0000;
													assign node611 = (inp[10]) ? node613 : 4'b1011;
														assign node613 = (inp[1]) ? node617 : node614;
															assign node614 = (inp[14]) ? 4'b1011 : 4'b0000;
															assign node617 = (inp[11]) ? 4'b0001 : 4'b0000;
												assign node620 = (inp[1]) ? node628 : node621;
													assign node621 = (inp[14]) ? node625 : node622;
														assign node622 = (inp[10]) ? 4'b1000 : 4'b0000;
														assign node625 = (inp[11]) ? 4'b1000 : 4'b1001;
													assign node628 = (inp[12]) ? node630 : 4'b1001;
														assign node630 = (inp[11]) ? node632 : 4'b1000;
															assign node632 = (inp[14]) ? 4'b1001 : 4'b0001;
										assign node636 = (inp[1]) ? node674 : node637;
											assign node637 = (inp[14]) ? node649 : node638;
												assign node638 = (inp[13]) ? node644 : node639;
													assign node639 = (inp[10]) ? 4'b0000 : node640;
														assign node640 = (inp[12]) ? 4'b1000 : 4'b0000;
													assign node644 = (inp[10]) ? 4'b1000 : node645;
														assign node645 = (inp[12]) ? 4'b0000 : 4'b1000;
												assign node649 = (inp[11]) ? node663 : node650;
													assign node650 = (inp[13]) ? node658 : node651;
														assign node651 = (inp[7]) ? node653 : 4'b1001;
															assign node653 = (inp[10]) ? node655 : 4'b1011;
																assign node655 = (inp[12]) ? 4'b1011 : 4'b0001;
														assign node658 = (inp[12]) ? 4'b0001 : node659;
															assign node659 = (inp[10]) ? 4'b1001 : 4'b0001;
													assign node663 = (inp[13]) ? node669 : node664;
														assign node664 = (inp[12]) ? node666 : 4'b0000;
															assign node666 = (inp[10]) ? 4'b0000 : 4'b1011;
														assign node669 = (inp[10]) ? 4'b1000 : node670;
															assign node670 = (inp[7]) ? 4'b0000 : 4'b1000;
											assign node674 = (inp[13]) ? node688 : node675;
												assign node675 = (inp[14]) ? node677 : 4'b0001;
													assign node677 = (inp[11]) ? node681 : node678;
														assign node678 = (inp[10]) ? 4'b0000 : 4'b1000;
														assign node681 = (inp[12]) ? node683 : 4'b0001;
															assign node683 = (inp[7]) ? 4'b1011 : node684;
																assign node684 = (inp[10]) ? 4'b0001 : 4'b1001;
												assign node688 = (inp[10]) ? node698 : node689;
													assign node689 = (inp[12]) ? node693 : node690;
														assign node690 = (inp[11]) ? 4'b1001 : 4'b1000;
														assign node693 = (inp[7]) ? 4'b0001 : node694;
															assign node694 = (inp[11]) ? 4'b0001 : 4'b0000;
													assign node698 = (inp[7]) ? node700 : 4'b1001;
														assign node700 = (inp[14]) ? 4'b1000 : 4'b1001;
							assign node704 = (inp[2]) ? node968 : node705;
								assign node705 = (inp[1]) ? node829 : node706;
									assign node706 = (inp[14]) ? node746 : node707;
										assign node707 = (inp[13]) ? node721 : node708;
											assign node708 = (inp[12]) ? node716 : node709;
												assign node709 = (inp[3]) ? 4'b0000 : node710;
													assign node710 = (inp[7]) ? node712 : 4'b0100;
														assign node712 = (inp[4]) ? 4'b0100 : 4'b0000;
												assign node716 = (inp[10]) ? 4'b0100 : node717;
													assign node717 = (inp[3]) ? 4'b1100 : 4'b1000;
											assign node721 = (inp[10]) ? node735 : node722;
												assign node722 = (inp[12]) ? node728 : node723;
													assign node723 = (inp[4]) ? node725 : 4'b1000;
														assign node725 = (inp[3]) ? 4'b1000 : 4'b1100;
													assign node728 = (inp[3]) ? 4'b0000 : node729;
														assign node729 = (inp[4]) ? 4'b0100 : node730;
															assign node730 = (inp[7]) ? 4'b0000 : 4'b0100;
												assign node735 = (inp[3]) ? node741 : node736;
													assign node736 = (inp[7]) ? node738 : 4'b1100;
														assign node738 = (inp[4]) ? 4'b1100 : 4'b1000;
													assign node741 = (inp[4]) ? 4'b1000 : node742;
														assign node742 = (inp[7]) ? 4'b1100 : 4'b1000;
										assign node746 = (inp[11]) ? node788 : node747;
											assign node747 = (inp[13]) ? node767 : node748;
												assign node748 = (inp[12]) ? node760 : node749;
													assign node749 = (inp[10]) ? node751 : 4'b1101;
														assign node751 = (inp[7]) ? node753 : 4'b0101;
															assign node753 = (inp[4]) ? node757 : node754;
																assign node754 = (inp[3]) ? 4'b0101 : 4'b0001;
																assign node757 = (inp[3]) ? 4'b0001 : 4'b0101;
													assign node760 = (inp[3]) ? node762 : 4'b1001;
														assign node762 = (inp[4]) ? node764 : 4'b1101;
															assign node764 = (inp[7]) ? 4'b1101 : 4'b1001;
												assign node767 = (inp[3]) ? node779 : node768;
													assign node768 = (inp[4]) ? node774 : node769;
														assign node769 = (inp[7]) ? node771 : 4'b0101;
															assign node771 = (inp[12]) ? 4'b0001 : 4'b1001;
														assign node774 = (inp[10]) ? node776 : 4'b0101;
															assign node776 = (inp[12]) ? 4'b0101 : 4'b1101;
													assign node779 = (inp[12]) ? node783 : node780;
														assign node780 = (inp[10]) ? 4'b1001 : 4'b0001;
														assign node783 = (inp[7]) ? node785 : 4'b0001;
															assign node785 = (inp[4]) ? 4'b0001 : 4'b0101;
											assign node788 = (inp[13]) ? node806 : node789;
												assign node789 = (inp[12]) ? node799 : node790;
													assign node790 = (inp[4]) ? node796 : node791;
														assign node791 = (inp[7]) ? node793 : 4'b0100;
															assign node793 = (inp[3]) ? 4'b0100 : 4'b0000;
														assign node796 = (inp[3]) ? 4'b0000 : 4'b0100;
													assign node799 = (inp[10]) ? node803 : node800;
														assign node800 = (inp[4]) ? 4'b1100 : 4'b1000;
														assign node803 = (inp[3]) ? 4'b0000 : 4'b0100;
												assign node806 = (inp[3]) ? node816 : node807;
													assign node807 = (inp[4]) ? node811 : node808;
														assign node808 = (inp[10]) ? 4'b1000 : 4'b1100;
														assign node811 = (inp[10]) ? 4'b1100 : node812;
															assign node812 = (inp[12]) ? 4'b0100 : 4'b1100;
													assign node816 = (inp[12]) ? node818 : 4'b1000;
														assign node818 = (inp[10]) ? node824 : node819;
															assign node819 = (inp[7]) ? node821 : 4'b0000;
																assign node821 = (inp[4]) ? 4'b0000 : 4'b0100;
															assign node824 = (inp[4]) ? 4'b1000 : node825;
																assign node825 = (inp[7]) ? 4'b1100 : 4'b1000;
									assign node829 = (inp[14]) ? node883 : node830;
										assign node830 = (inp[3]) ? node848 : node831;
											assign node831 = (inp[13]) ? node843 : node832;
												assign node832 = (inp[12]) ? node834 : 4'b0101;
													assign node834 = (inp[10]) ? node840 : node835;
														assign node835 = (inp[4]) ? node837 : 4'b1001;
															assign node837 = (inp[7]) ? 4'b1001 : 4'b1101;
														assign node840 = (inp[7]) ? 4'b0001 : 4'b0101;
												assign node843 = (inp[10]) ? 4'b1101 : node844;
													assign node844 = (inp[12]) ? 4'b0101 : 4'b1101;
											assign node848 = (inp[7]) ? node862 : node849;
												assign node849 = (inp[13]) ? node857 : node850;
													assign node850 = (inp[10]) ? 4'b0001 : node851;
														assign node851 = (inp[12]) ? node853 : 4'b0001;
															assign node853 = (inp[11]) ? 4'b1001 : 4'b1101;
													assign node857 = (inp[12]) ? node859 : 4'b1001;
														assign node859 = (inp[10]) ? 4'b1001 : 4'b0001;
												assign node862 = (inp[4]) ? node874 : node863;
													assign node863 = (inp[13]) ? node869 : node864;
														assign node864 = (inp[10]) ? 4'b0101 : node865;
															assign node865 = (inp[12]) ? 4'b1101 : 4'b0101;
														assign node869 = (inp[10]) ? 4'b1101 : node870;
															assign node870 = (inp[12]) ? 4'b0101 : 4'b1101;
													assign node874 = (inp[10]) ? node880 : node875;
														assign node875 = (inp[13]) ? 4'b0001 : node876;
															assign node876 = (inp[12]) ? 4'b1101 : 4'b0001;
														assign node880 = (inp[13]) ? 4'b1001 : 4'b0001;
										assign node883 = (inp[11]) ? node925 : node884;
											assign node884 = (inp[13]) ? node906 : node885;
												assign node885 = (inp[10]) ? node899 : node886;
													assign node886 = (inp[12]) ? node892 : node887;
														assign node887 = (inp[4]) ? node889 : 4'b0100;
															assign node889 = (inp[3]) ? 4'b0000 : 4'b0100;
														assign node892 = (inp[3]) ? 4'b1100 : node893;
															assign node893 = (inp[4]) ? node895 : 4'b1000;
																assign node895 = (inp[7]) ? 4'b1000 : 4'b1100;
													assign node899 = (inp[3]) ? node901 : 4'b0100;
														assign node901 = (inp[7]) ? node903 : 4'b0000;
															assign node903 = (inp[12]) ? 4'b0000 : 4'b0100;
												assign node906 = (inp[12]) ? node916 : node907;
													assign node907 = (inp[3]) ? node911 : node908;
														assign node908 = (inp[7]) ? 4'b1000 : 4'b1100;
														assign node911 = (inp[7]) ? node913 : 4'b1000;
															assign node913 = (inp[4]) ? 4'b1000 : 4'b1100;
													assign node916 = (inp[10]) ? node922 : node917;
														assign node917 = (inp[3]) ? 4'b0000 : node918;
															assign node918 = (inp[7]) ? 4'b0000 : 4'b0100;
														assign node922 = (inp[3]) ? 4'b1000 : 4'b1100;
											assign node925 = (inp[3]) ? node947 : node926;
												assign node926 = (inp[4]) ? node938 : node927;
													assign node927 = (inp[7]) ? node933 : node928;
														assign node928 = (inp[13]) ? node930 : 4'b1001;
															assign node930 = (inp[12]) ? 4'b0101 : 4'b1101;
														assign node933 = (inp[10]) ? 4'b0001 : node934;
															assign node934 = (inp[13]) ? 4'b0001 : 4'b1001;
													assign node938 = (inp[13]) ? node942 : node939;
														assign node939 = (inp[10]) ? 4'b0101 : 4'b1101;
														assign node942 = (inp[12]) ? node944 : 4'b1101;
															assign node944 = (inp[10]) ? 4'b1101 : 4'b0101;
												assign node947 = (inp[4]) ? node957 : node948;
													assign node948 = (inp[12]) ? node952 : node949;
														assign node949 = (inp[13]) ? 4'b1001 : 4'b0001;
														assign node952 = (inp[13]) ? node954 : 4'b1101;
															assign node954 = (inp[7]) ? 4'b0101 : 4'b0001;
													assign node957 = (inp[13]) ? node963 : node958;
														assign node958 = (inp[7]) ? 4'b0001 : node959;
															assign node959 = (inp[12]) ? 4'b1001 : 4'b0001;
														assign node963 = (inp[12]) ? node965 : 4'b1001;
															assign node965 = (inp[10]) ? 4'b1001 : 4'b0001;
								assign node968 = (inp[3]) ? node970 : 4'b1011;
									assign node970 = (inp[4]) ? node1014 : node971;
										assign node971 = (inp[7]) ? 4'b1011 : node972;
											assign node972 = (inp[13]) ? node990 : node973;
												assign node973 = (inp[10]) ? node979 : node974;
													assign node974 = (inp[12]) ? 4'b1011 : node975;
														assign node975 = (inp[1]) ? 4'b0001 : 4'b1011;
													assign node979 = (inp[1]) ? node985 : node980;
														assign node980 = (inp[14]) ? node982 : 4'b0000;
															assign node982 = (inp[11]) ? 4'b0000 : 4'b0001;
														assign node985 = (inp[12]) ? node987 : 4'b0001;
															assign node987 = (inp[11]) ? 4'b0001 : 4'b0000;
												assign node990 = (inp[10]) ? node1002 : node991;
													assign node991 = (inp[14]) ? node995 : node992;
														assign node992 = (inp[1]) ? 4'b1001 : 4'b1000;
														assign node995 = (inp[1]) ? node999 : node996;
															assign node996 = (inp[11]) ? 4'b0000 : 4'b0001;
															assign node999 = (inp[12]) ? 4'b0000 : 4'b1000;
													assign node1002 = (inp[1]) ? node1008 : node1003;
														assign node1003 = (inp[11]) ? 4'b1000 : node1004;
															assign node1004 = (inp[12]) ? 4'b0001 : 4'b1001;
														assign node1008 = (inp[11]) ? 4'b1001 : node1009;
															assign node1009 = (inp[14]) ? 4'b1000 : 4'b1001;
										assign node1014 = (inp[1]) ? node1040 : node1015;
											assign node1015 = (inp[11]) ? node1029 : node1016;
												assign node1016 = (inp[14]) ? node1022 : node1017;
													assign node1017 = (inp[12]) ? 4'b0000 : node1018;
														assign node1018 = (inp[13]) ? 4'b1000 : 4'b0000;
													assign node1022 = (inp[13]) ? 4'b0001 : node1023;
														assign node1023 = (inp[7]) ? 4'b1011 : node1024;
															assign node1024 = (inp[12]) ? 4'b1001 : 4'b0001;
												assign node1029 = (inp[13]) ? node1035 : node1030;
													assign node1030 = (inp[10]) ? 4'b0000 : node1031;
														assign node1031 = (inp[12]) ? 4'b1011 : 4'b0000;
													assign node1035 = (inp[12]) ? node1037 : 4'b1000;
														assign node1037 = (inp[10]) ? 4'b1000 : 4'b0000;
											assign node1040 = (inp[14]) ? node1054 : node1041;
												assign node1041 = (inp[13]) ? node1049 : node1042;
													assign node1042 = (inp[10]) ? 4'b0001 : node1043;
														assign node1043 = (inp[12]) ? node1045 : 4'b0001;
															assign node1045 = (inp[7]) ? 4'b1011 : 4'b1001;
													assign node1049 = (inp[12]) ? node1051 : 4'b1001;
														assign node1051 = (inp[10]) ? 4'b1001 : 4'b0001;
												assign node1054 = (inp[11]) ? node1064 : node1055;
													assign node1055 = (inp[13]) ? node1061 : node1056;
														assign node1056 = (inp[10]) ? 4'b0000 : node1057;
															assign node1057 = (inp[7]) ? 4'b0000 : 4'b1000;
														assign node1061 = (inp[7]) ? 4'b1000 : 4'b0000;
													assign node1064 = (inp[7]) ? 4'b0001 : node1065;
														assign node1065 = (inp[10]) ? node1071 : node1066;
															assign node1066 = (inp[12]) ? node1068 : 4'b0001;
																assign node1068 = (inp[13]) ? 4'b0001 : 4'b1001;
															assign node1071 = (inp[13]) ? 4'b1001 : 4'b0001;
				assign node1076 = (inp[5]) ? node2568 : node1077;
					assign node1077 = (inp[0]) ? node2221 : node1078;
						assign node1078 = (inp[11]) ? node1714 : node1079;
							assign node1079 = (inp[10]) ? node1397 : node1080;
								assign node1080 = (inp[12]) ? node1220 : node1081;
									assign node1081 = (inp[2]) ? node1139 : node1082;
										assign node1082 = (inp[15]) ? node1106 : node1083;
											assign node1083 = (inp[4]) ? node1089 : node1084;
												assign node1084 = (inp[7]) ? node1086 : 4'b0000;
													assign node1086 = (inp[13]) ? 4'b0000 : 4'b0100;
												assign node1089 = (inp[3]) ? node1095 : node1090;
													assign node1090 = (inp[13]) ? 4'b0100 : node1091;
														assign node1091 = (inp[7]) ? 4'b0000 : 4'b0100;
													assign node1095 = (inp[13]) ? node1103 : node1096;
														assign node1096 = (inp[14]) ? node1100 : node1097;
															assign node1097 = (inp[1]) ? 4'b1000 : 4'b0001;
															assign node1100 = (inp[1]) ? 4'b0001 : 4'b0000;
														assign node1103 = (inp[7]) ? 4'b1000 : 4'b0100;
											assign node1106 = (inp[4]) ? node1124 : node1107;
												assign node1107 = (inp[3]) ? node1119 : node1108;
													assign node1108 = (inp[7]) ? node1114 : node1109;
														assign node1109 = (inp[13]) ? node1111 : 4'b1001;
															assign node1111 = (inp[1]) ? 4'b1100 : 4'b0101;
														assign node1114 = (inp[13]) ? 4'b1000 : node1115;
															assign node1115 = (inp[14]) ? 4'b0000 : 4'b0001;
													assign node1119 = (inp[13]) ? 4'b0100 : node1120;
														assign node1120 = (inp[7]) ? 4'b0000 : 4'b0100;
												assign node1124 = (inp[7]) ? node1130 : node1125;
													assign node1125 = (inp[3]) ? node1127 : 4'b0000;
														assign node1127 = (inp[13]) ? 4'b1001 : 4'b0000;
													assign node1130 = (inp[13]) ? 4'b0000 : node1131;
														assign node1131 = (inp[3]) ? 4'b0100 : node1132;
															assign node1132 = (inp[14]) ? 4'b1001 : node1133;
																assign node1133 = (inp[1]) ? 4'b0101 : 4'b0100;
										assign node1139 = (inp[3]) ? node1185 : node1140;
											assign node1140 = (inp[13]) ? node1158 : node1141;
												assign node1141 = (inp[1]) ? node1147 : node1142;
													assign node1142 = (inp[14]) ? node1144 : 4'b0100;
														assign node1144 = (inp[15]) ? 4'b1001 : 4'b1101;
													assign node1147 = (inp[14]) ? node1151 : node1148;
														assign node1148 = (inp[15]) ? 4'b0101 : 4'b0001;
														assign node1151 = (inp[4]) ? node1155 : node1152;
															assign node1152 = (inp[15]) ? 4'b0000 : 4'b0100;
															assign node1155 = (inp[15]) ? 4'b0100 : 4'b0000;
												assign node1158 = (inp[1]) ? node1170 : node1159;
													assign node1159 = (inp[14]) ? 4'b0001 : node1160;
														assign node1160 = (inp[7]) ? node1162 : 4'b1000;
															assign node1162 = (inp[4]) ? node1166 : node1163;
																assign node1163 = (inp[15]) ? 4'b1000 : 4'b1100;
																assign node1166 = (inp[15]) ? 4'b1100 : 4'b1000;
													assign node1170 = (inp[14]) ? node1176 : node1171;
														assign node1171 = (inp[15]) ? node1173 : 4'b1101;
															assign node1173 = (inp[7]) ? 4'b1001 : 4'b1101;
														assign node1176 = (inp[7]) ? node1178 : 4'b1100;
															assign node1178 = (inp[4]) ? node1182 : node1179;
																assign node1179 = (inp[15]) ? 4'b1000 : 4'b1100;
																assign node1182 = (inp[15]) ? 4'b1100 : 4'b1000;
											assign node1185 = (inp[15]) ? node1193 : node1186;
												assign node1186 = (inp[4]) ? node1188 : 4'b0000;
													assign node1188 = (inp[7]) ? node1190 : 4'b0100;
														assign node1190 = (inp[13]) ? 4'b0100 : 4'b0000;
												assign node1193 = (inp[4]) ? node1215 : node1194;
													assign node1194 = (inp[7]) ? node1204 : node1195;
														assign node1195 = (inp[13]) ? node1199 : node1196;
															assign node1196 = (inp[1]) ? 4'b0001 : 4'b0000;
															assign node1199 = (inp[14]) ? 4'b1000 : node1200;
																assign node1200 = (inp[1]) ? 4'b1001 : 4'b1000;
														assign node1204 = (inp[14]) ? node1208 : node1205;
															assign node1205 = (inp[1]) ? 4'b1101 : 4'b1100;
															assign node1208 = (inp[1]) ? node1212 : node1209;
																assign node1209 = (inp[13]) ? 4'b0101 : 4'b1101;
																assign node1212 = (inp[13]) ? 4'b1100 : 4'b0100;
													assign node1215 = (inp[14]) ? 4'b0000 : node1216;
														assign node1216 = (inp[7]) ? 4'b0001 : 4'b0000;
									assign node1220 = (inp[13]) ? node1300 : node1221;
										assign node1221 = (inp[1]) ? node1255 : node1222;
											assign node1222 = (inp[14]) ? node1234 : node1223;
												assign node1223 = (inp[4]) ? node1229 : node1224;
													assign node1224 = (inp[3]) ? 4'b1100 : node1225;
														assign node1225 = (inp[15]) ? 4'b1000 : 4'b1100;
													assign node1229 = (inp[2]) ? 4'b1000 : node1230;
														assign node1230 = (inp[15]) ? 4'b1100 : 4'b1000;
												assign node1234 = (inp[2]) ? node1248 : node1235;
													assign node1235 = (inp[3]) ? node1239 : node1236;
														assign node1236 = (inp[15]) ? 4'b1001 : 4'b1101;
														assign node1239 = (inp[7]) ? node1241 : 4'b1100;
															assign node1241 = (inp[15]) ? node1245 : node1242;
																assign node1242 = (inp[4]) ? 4'b1000 : 4'b1100;
																assign node1245 = (inp[4]) ? 4'b1100 : 4'b1000;
													assign node1248 = (inp[7]) ? node1250 : 4'b1001;
														assign node1250 = (inp[15]) ? 4'b1101 : node1251;
															assign node1251 = (inp[3]) ? 4'b1001 : 4'b1101;
											assign node1255 = (inp[3]) ? node1273 : node1256;
												assign node1256 = (inp[14]) ? node1266 : node1257;
													assign node1257 = (inp[7]) ? 4'b1101 : node1258;
														assign node1258 = (inp[15]) ? 4'b1001 : node1259;
															assign node1259 = (inp[2]) ? node1261 : 4'b0100;
																assign node1261 = (inp[4]) ? 4'b1001 : 4'b1101;
													assign node1266 = (inp[15]) ? 4'b1000 : node1267;
														assign node1267 = (inp[2]) ? 4'b1100 : node1268;
															assign node1268 = (inp[4]) ? 4'b0100 : 4'b0000;
												assign node1273 = (inp[7]) ? node1291 : node1274;
													assign node1274 = (inp[14]) ? node1282 : node1275;
														assign node1275 = (inp[4]) ? node1279 : node1276;
															assign node1276 = (inp[15]) ? 4'b0100 : 4'b0000;
															assign node1279 = (inp[15]) ? 4'b0000 : 4'b0100;
														assign node1282 = (inp[2]) ? node1286 : node1283;
															assign node1283 = (inp[4]) ? 4'b0001 : 4'b0000;
															assign node1286 = (inp[4]) ? node1288 : 4'b0000;
																assign node1288 = (inp[15]) ? 4'b0000 : 4'b0100;
													assign node1291 = (inp[2]) ? node1295 : node1292;
														assign node1292 = (inp[14]) ? 4'b0100 : 4'b0000;
														assign node1295 = (inp[15]) ? node1297 : 4'b0000;
															assign node1297 = (inp[14]) ? 4'b1100 : 4'b1101;
										assign node1300 = (inp[2]) ? node1360 : node1301;
											assign node1301 = (inp[7]) ? node1329 : node1302;
												assign node1302 = (inp[15]) ? node1318 : node1303;
													assign node1303 = (inp[4]) ? node1307 : node1304;
														assign node1304 = (inp[1]) ? 4'b0000 : 4'b1000;
														assign node1307 = (inp[3]) ? node1311 : node1308;
															assign node1308 = (inp[1]) ? 4'b0100 : 4'b1100;
															assign node1311 = (inp[1]) ? node1315 : node1312;
																assign node1312 = (inp[14]) ? 4'b0100 : 4'b0101;
																assign node1315 = (inp[14]) ? 4'b1101 : 4'b1100;
													assign node1318 = (inp[4]) ? node1324 : node1319;
														assign node1319 = (inp[3]) ? 4'b1100 : node1320;
															assign node1320 = (inp[14]) ? 4'b0101 : 4'b0100;
														assign node1324 = (inp[3]) ? node1326 : 4'b0000;
															assign node1326 = (inp[1]) ? 4'b1001 : 4'b0001;
												assign node1329 = (inp[14]) ? node1347 : node1330;
													assign node1330 = (inp[3]) ? node1344 : node1331;
														assign node1331 = (inp[1]) ? node1337 : node1332;
															assign node1332 = (inp[4]) ? 4'b0100 : node1333;
																assign node1333 = (inp[15]) ? 4'b0000 : 4'b0100;
															assign node1337 = (inp[4]) ? node1341 : node1338;
																assign node1338 = (inp[15]) ? 4'b0001 : 4'b0000;
																assign node1341 = (inp[15]) ? 4'b0000 : 4'b0100;
														assign node1344 = (inp[4]) ? 4'b1100 : 4'b0100;
													assign node1347 = (inp[1]) ? node1355 : node1348;
														assign node1348 = (inp[4]) ? node1352 : node1349;
															assign node1349 = (inp[3]) ? 4'b1000 : 4'b0001;
															assign node1352 = (inp[3]) ? 4'b0000 : 4'b1000;
														assign node1355 = (inp[3]) ? node1357 : 4'b0000;
															assign node1357 = (inp[15]) ? 4'b0100 : 4'b0000;
											assign node1360 = (inp[3]) ? node1382 : node1361;
												assign node1361 = (inp[15]) ? node1373 : node1362;
													assign node1362 = (inp[4]) ? node1366 : node1363;
														assign node1363 = (inp[1]) ? 4'b0101 : 4'b0100;
														assign node1366 = (inp[14]) ? node1370 : node1367;
															assign node1367 = (inp[1]) ? 4'b0001 : 4'b0000;
															assign node1370 = (inp[1]) ? 4'b0000 : 4'b0001;
													assign node1373 = (inp[4]) ? node1379 : node1374;
														assign node1374 = (inp[14]) ? node1376 : 4'b0000;
															assign node1376 = (inp[7]) ? 4'b0001 : 4'b0101;
														assign node1379 = (inp[7]) ? 4'b0101 : 4'b0100;
												assign node1382 = (inp[14]) ? node1388 : node1383;
													assign node1383 = (inp[15]) ? 4'b0000 : node1384;
														assign node1384 = (inp[4]) ? 4'b1000 : 4'b0000;
													assign node1388 = (inp[1]) ? node1392 : node1389;
														assign node1389 = (inp[4]) ? 4'b1100 : 4'b0001;
														assign node1392 = (inp[15]) ? node1394 : 4'b0100;
															assign node1394 = (inp[4]) ? 4'b0000 : 4'b0100;
								assign node1397 = (inp[13]) ? node1555 : node1398;
									assign node1398 = (inp[7]) ? node1478 : node1399;
										assign node1399 = (inp[2]) ? node1435 : node1400;
											assign node1400 = (inp[1]) ? node1418 : node1401;
												assign node1401 = (inp[12]) ? node1411 : node1402;
													assign node1402 = (inp[15]) ? 4'b1000 : node1403;
														assign node1403 = (inp[3]) ? node1407 : node1404;
															assign node1404 = (inp[4]) ? 4'b1100 : 4'b1000;
															assign node1407 = (inp[4]) ? 4'b1001 : 4'b1000;
													assign node1411 = (inp[4]) ? 4'b0100 : node1412;
														assign node1412 = (inp[3]) ? 4'b0100 : node1413;
															assign node1413 = (inp[15]) ? 4'b1001 : 4'b0000;
												assign node1418 = (inp[4]) ? node1426 : node1419;
													assign node1419 = (inp[15]) ? node1421 : 4'b1000;
														assign node1421 = (inp[3]) ? 4'b1100 : node1422;
															assign node1422 = (inp[12]) ? 4'b0101 : 4'b0100;
													assign node1426 = (inp[3]) ? node1430 : node1427;
														assign node1427 = (inp[15]) ? 4'b1000 : 4'b1100;
														assign node1430 = (inp[14]) ? 4'b0101 : node1431;
															assign node1431 = (inp[15]) ? 4'b0000 : 4'b0100;
											assign node1435 = (inp[3]) ? node1455 : node1436;
												assign node1436 = (inp[15]) ? node1444 : node1437;
													assign node1437 = (inp[14]) ? node1441 : node1438;
														assign node1438 = (inp[1]) ? 4'b0001 : 4'b0000;
														assign node1441 = (inp[1]) ? 4'b0000 : 4'b0001;
													assign node1444 = (inp[12]) ? node1450 : node1445;
														assign node1445 = (inp[14]) ? node1447 : 4'b0101;
															assign node1447 = (inp[1]) ? 4'b0100 : 4'b0101;
														assign node1450 = (inp[14]) ? node1452 : 4'b0100;
															assign node1452 = (inp[1]) ? 4'b0100 : 4'b1001;
												assign node1455 = (inp[15]) ? node1467 : node1456;
													assign node1456 = (inp[4]) ? node1462 : node1457;
														assign node1457 = (inp[12]) ? node1459 : 4'b1000;
															assign node1459 = (inp[1]) ? 4'b1000 : 4'b0000;
														assign node1462 = (inp[1]) ? 4'b1100 : node1463;
															assign node1463 = (inp[12]) ? 4'b0100 : 4'b1100;
													assign node1467 = (inp[4]) ? node1475 : node1468;
														assign node1468 = (inp[1]) ? node1472 : node1469;
															assign node1469 = (inp[14]) ? 4'b1101 : 4'b0000;
															assign node1472 = (inp[14]) ? 4'b0000 : 4'b0001;
														assign node1475 = (inp[1]) ? 4'b1000 : 4'b0000;
										assign node1478 = (inp[3]) ? node1512 : node1479;
											assign node1479 = (inp[15]) ? node1497 : node1480;
												assign node1480 = (inp[4]) ? node1490 : node1481;
													assign node1481 = (inp[1]) ? node1487 : node1482;
														assign node1482 = (inp[14]) ? node1484 : 4'b0100;
															assign node1484 = (inp[12]) ? 4'b1101 : 4'b0101;
														assign node1487 = (inp[14]) ? 4'b0100 : 4'b0101;
													assign node1490 = (inp[14]) ? node1494 : node1491;
														assign node1491 = (inp[1]) ? 4'b1000 : 4'b0000;
														assign node1494 = (inp[12]) ? 4'b1101 : 4'b0001;
												assign node1497 = (inp[4]) ? node1503 : node1498;
													assign node1498 = (inp[1]) ? node1500 : 4'b0000;
														assign node1500 = (inp[14]) ? 4'b0000 : 4'b0001;
													assign node1503 = (inp[12]) ? 4'b0100 : node1504;
														assign node1504 = (inp[1]) ? node1508 : node1505;
															assign node1505 = (inp[14]) ? 4'b0101 : 4'b0100;
															assign node1508 = (inp[14]) ? 4'b0100 : 4'b0101;
											assign node1512 = (inp[15]) ? node1540 : node1513;
												assign node1513 = (inp[1]) ? node1525 : node1514;
													assign node1514 = (inp[4]) ? node1520 : node1515;
														assign node1515 = (inp[2]) ? 4'b1001 : node1516;
															assign node1516 = (inp[14]) ? 4'b0100 : 4'b1100;
														assign node1520 = (inp[2]) ? 4'b0000 : node1521;
															assign node1521 = (inp[14]) ? 4'b1000 : 4'b1001;
													assign node1525 = (inp[12]) ? node1533 : node1526;
														assign node1526 = (inp[4]) ? node1530 : node1527;
															assign node1527 = (inp[14]) ? 4'b0000 : 4'b0001;
															assign node1530 = (inp[14]) ? 4'b0001 : 4'b0000;
														assign node1533 = (inp[4]) ? node1535 : 4'b0001;
															assign node1535 = (inp[14]) ? 4'b1001 : node1536;
																assign node1536 = (inp[2]) ? 4'b1000 : 4'b0000;
												assign node1540 = (inp[2]) ? node1548 : node1541;
													assign node1541 = (inp[4]) ? node1545 : node1542;
														assign node1542 = (inp[1]) ? 4'b1000 : 4'b0000;
														assign node1545 = (inp[1]) ? 4'b1100 : 4'b0100;
													assign node1548 = (inp[4]) ? 4'b0001 : node1549;
														assign node1549 = (inp[1]) ? 4'b0100 : node1550;
															assign node1550 = (inp[12]) ? 4'b1101 : 4'b0101;
									assign node1555 = (inp[1]) ? node1637 : node1556;
										assign node1556 = (inp[12]) ? node1604 : node1557;
											assign node1557 = (inp[2]) ? node1579 : node1558;
												assign node1558 = (inp[4]) ? node1570 : node1559;
													assign node1559 = (inp[15]) ? node1567 : node1560;
														assign node1560 = (inp[3]) ? node1562 : 4'b1000;
															assign node1562 = (inp[7]) ? 4'b1000 : node1563;
																assign node1563 = (inp[14]) ? 4'b0000 : 4'b0001;
														assign node1567 = (inp[3]) ? 4'b1100 : 4'b1101;
													assign node1570 = (inp[3]) ? node1574 : node1571;
														assign node1571 = (inp[15]) ? 4'b1000 : 4'b1100;
														assign node1574 = (inp[15]) ? node1576 : 4'b0101;
															assign node1576 = (inp[14]) ? 4'b0000 : 4'b0001;
												assign node1579 = (inp[14]) ? node1589 : node1580;
													assign node1580 = (inp[4]) ? node1582 : 4'b1000;
														assign node1582 = (inp[3]) ? node1586 : node1583;
															assign node1583 = (inp[7]) ? 4'b1100 : 4'b1000;
															assign node1586 = (inp[15]) ? 4'b1000 : 4'b1100;
													assign node1589 = (inp[3]) ? node1597 : node1590;
														assign node1590 = (inp[7]) ? node1592 : 4'b1001;
															assign node1592 = (inp[4]) ? node1594 : 4'b1101;
																assign node1594 = (inp[15]) ? 4'b1101 : 4'b1001;
														assign node1597 = (inp[7]) ? node1599 : 4'b1000;
															assign node1599 = (inp[4]) ? node1601 : 4'b1101;
																assign node1601 = (inp[15]) ? 4'b1000 : 4'b1100;
											assign node1604 = (inp[15]) ? node1620 : node1605;
												assign node1605 = (inp[4]) ? node1613 : node1606;
													assign node1606 = (inp[3]) ? 4'b0000 : node1607;
														assign node1607 = (inp[14]) ? 4'b0101 : node1608;
															assign node1608 = (inp[7]) ? 4'b1100 : 4'b1000;
													assign node1613 = (inp[7]) ? 4'b0100 : node1614;
														assign node1614 = (inp[2]) ? node1616 : 4'b0100;
															assign node1616 = (inp[3]) ? 4'b0100 : 4'b1000;
												assign node1620 = (inp[14]) ? node1628 : node1621;
													assign node1621 = (inp[4]) ? node1623 : 4'b1000;
														assign node1623 = (inp[2]) ? 4'b0000 : node1624;
															assign node1624 = (inp[3]) ? 4'b0001 : 4'b0000;
													assign node1628 = (inp[3]) ? node1632 : node1629;
														assign node1629 = (inp[7]) ? 4'b0001 : 4'b0101;
														assign node1632 = (inp[4]) ? 4'b0000 : node1633;
															assign node1633 = (inp[2]) ? 4'b0101 : 4'b0100;
										assign node1637 = (inp[14]) ? node1667 : node1638;
											assign node1638 = (inp[3]) ? node1658 : node1639;
												assign node1639 = (inp[2]) ? node1649 : node1640;
													assign node1640 = (inp[15]) ? node1644 : node1641;
														assign node1641 = (inp[4]) ? 4'b1100 : 4'b1000;
														assign node1644 = (inp[4]) ? 4'b1000 : node1645;
															assign node1645 = (inp[12]) ? 4'b1001 : 4'b1101;
													assign node1649 = (inp[7]) ? node1653 : node1650;
														assign node1650 = (inp[15]) ? 4'b1101 : 4'b1001;
														assign node1653 = (inp[15]) ? 4'b1001 : node1654;
															assign node1654 = (inp[12]) ? 4'b1101 : 4'b1001;
												assign node1658 = (inp[15]) ? node1662 : node1659;
													assign node1659 = (inp[4]) ? 4'b1100 : 4'b1000;
													assign node1662 = (inp[4]) ? 4'b1000 : node1663;
														assign node1663 = (inp[2]) ? 4'b1101 : 4'b1100;
											assign node1667 = (inp[3]) ? node1691 : node1668;
												assign node1668 = (inp[15]) ? node1680 : node1669;
													assign node1669 = (inp[12]) ? node1675 : node1670;
														assign node1670 = (inp[4]) ? 4'b1100 : node1671;
															assign node1671 = (inp[2]) ? 4'b1100 : 4'b1000;
														assign node1675 = (inp[2]) ? 4'b1000 : node1676;
															assign node1676 = (inp[4]) ? 4'b1100 : 4'b1000;
													assign node1680 = (inp[7]) ? node1686 : node1681;
														assign node1681 = (inp[4]) ? node1683 : 4'b1100;
															assign node1683 = (inp[2]) ? 4'b1100 : 4'b1000;
														assign node1686 = (inp[4]) ? node1688 : 4'b1000;
															assign node1688 = (inp[2]) ? 4'b1100 : 4'b1000;
												assign node1691 = (inp[2]) ? node1705 : node1692;
													assign node1692 = (inp[12]) ? node1702 : node1693;
														assign node1693 = (inp[4]) ? node1699 : node1694;
															assign node1694 = (inp[15]) ? 4'b1100 : node1695;
																assign node1695 = (inp[7]) ? 4'b1000 : 4'b1001;
															assign node1699 = (inp[15]) ? 4'b1001 : 4'b1101;
														assign node1702 = (inp[15]) ? 4'b0001 : 4'b0101;
													assign node1705 = (inp[4]) ? node1711 : node1706;
														assign node1706 = (inp[7]) ? node1708 : 4'b1000;
															assign node1708 = (inp[12]) ? 4'b1100 : 4'b1000;
														assign node1711 = (inp[15]) ? 4'b1000 : 4'b1100;
							assign node1714 = (inp[1]) ? node1998 : node1715;
								assign node1715 = (inp[3]) ? node1861 : node1716;
									assign node1716 = (inp[2]) ? node1794 : node1717;
										assign node1717 = (inp[15]) ? node1765 : node1718;
											assign node1718 = (inp[4]) ? node1742 : node1719;
												assign node1719 = (inp[13]) ? node1733 : node1720;
													assign node1720 = (inp[7]) ? node1728 : node1721;
														assign node1721 = (inp[12]) ? node1725 : node1722;
															assign node1722 = (inp[14]) ? 4'b0001 : 4'b1001;
															assign node1725 = (inp[10]) ? 4'b0001 : 4'b1100;
														assign node1728 = (inp[12]) ? node1730 : 4'b0100;
															assign node1730 = (inp[14]) ? 4'b1100 : 4'b0100;
													assign node1733 = (inp[12]) ? node1737 : node1734;
														assign node1734 = (inp[10]) ? 4'b1001 : 4'b0001;
														assign node1737 = (inp[7]) ? node1739 : 4'b1001;
															assign node1739 = (inp[14]) ? 4'b0001 : 4'b0100;
												assign node1742 = (inp[13]) ? node1758 : node1743;
													assign node1743 = (inp[7]) ? node1745 : 4'b1001;
														assign node1745 = (inp[14]) ? node1753 : node1746;
															assign node1746 = (inp[12]) ? node1750 : node1747;
																assign node1747 = (inp[10]) ? 4'b1001 : 4'b0001;
																assign node1750 = (inp[10]) ? 4'b0001 : 4'b1001;
															assign node1753 = (inp[10]) ? node1755 : 4'b0001;
																assign node1755 = (inp[12]) ? 4'b0001 : 4'b1001;
													assign node1758 = (inp[14]) ? node1760 : 4'b0101;
														assign node1760 = (inp[10]) ? 4'b1101 : node1761;
															assign node1761 = (inp[12]) ? 4'b1101 : 4'b0101;
											assign node1765 = (inp[4]) ? node1781 : node1766;
												assign node1766 = (inp[7]) ? node1772 : node1767;
													assign node1767 = (inp[10]) ? 4'b0100 : node1768;
														assign node1768 = (inp[13]) ? 4'b1100 : 4'b1000;
													assign node1772 = (inp[10]) ? node1778 : node1773;
														assign node1773 = (inp[12]) ? node1775 : 4'b1000;
															assign node1775 = (inp[13]) ? 4'b0000 : 4'b1000;
														assign node1778 = (inp[12]) ? 4'b1000 : 4'b0000;
												assign node1781 = (inp[12]) ? node1789 : node1782;
													assign node1782 = (inp[10]) ? node1784 : 4'b0001;
														assign node1784 = (inp[13]) ? 4'b1001 : node1785;
															assign node1785 = (inp[7]) ? 4'b0100 : 4'b1001;
													assign node1789 = (inp[7]) ? 4'b0100 : node1790;
														assign node1790 = (inp[10]) ? 4'b0001 : 4'b1100;
										assign node1794 = (inp[13]) ? node1828 : node1795;
											assign node1795 = (inp[10]) ? node1817 : node1796;
												assign node1796 = (inp[12]) ? node1806 : node1797;
													assign node1797 = (inp[7]) ? node1801 : node1798;
														assign node1798 = (inp[15]) ? 4'b0100 : 4'b0000;
														assign node1801 = (inp[14]) ? node1803 : 4'b0100;
															assign node1803 = (inp[15]) ? 4'b0000 : 4'b0100;
													assign node1806 = (inp[15]) ? node1814 : node1807;
														assign node1807 = (inp[14]) ? node1809 : 4'b1100;
															assign node1809 = (inp[4]) ? node1811 : 4'b1100;
																assign node1811 = (inp[7]) ? 4'b1100 : 4'b1000;
														assign node1814 = (inp[7]) ? 4'b1000 : 4'b1100;
												assign node1817 = (inp[15]) ? node1823 : node1818;
													assign node1818 = (inp[4]) ? 4'b0000 : node1819;
														assign node1819 = (inp[7]) ? 4'b0100 : 4'b0000;
													assign node1823 = (inp[4]) ? 4'b0100 : node1824;
														assign node1824 = (inp[7]) ? 4'b0000 : 4'b0100;
											assign node1828 = (inp[12]) ? node1840 : node1829;
												assign node1829 = (inp[15]) ? node1835 : node1830;
													assign node1830 = (inp[7]) ? node1832 : 4'b1000;
														assign node1832 = (inp[4]) ? 4'b1000 : 4'b1100;
													assign node1835 = (inp[7]) ? node1837 : 4'b1100;
														assign node1837 = (inp[4]) ? 4'b1100 : 4'b1000;
												assign node1840 = (inp[10]) ? node1852 : node1841;
													assign node1841 = (inp[15]) ? node1847 : node1842;
														assign node1842 = (inp[4]) ? 4'b0000 : node1843;
															assign node1843 = (inp[7]) ? 4'b0100 : 4'b0000;
														assign node1847 = (inp[4]) ? 4'b0100 : node1848;
															assign node1848 = (inp[7]) ? 4'b0000 : 4'b0100;
													assign node1852 = (inp[15]) ? node1858 : node1853;
														assign node1853 = (inp[7]) ? node1855 : 4'b1000;
															assign node1855 = (inp[4]) ? 4'b1000 : 4'b1100;
														assign node1858 = (inp[7]) ? 4'b1000 : 4'b1100;
									assign node1861 = (inp[10]) ? node1925 : node1862;
										assign node1862 = (inp[12]) ? node1896 : node1863;
											assign node1863 = (inp[7]) ? node1875 : node1864;
												assign node1864 = (inp[14]) ? node1870 : node1865;
													assign node1865 = (inp[4]) ? node1867 : 4'b0001;
														assign node1867 = (inp[15]) ? 4'b0001 : 4'b0101;
													assign node1870 = (inp[15]) ? 4'b0101 : node1871;
														assign node1871 = (inp[4]) ? 4'b0101 : 4'b0001;
												assign node1875 = (inp[2]) ? node1889 : node1876;
													assign node1876 = (inp[4]) ? node1884 : node1877;
														assign node1877 = (inp[15]) ? node1881 : node1878;
															assign node1878 = (inp[13]) ? 4'b0001 : 4'b0101;
															assign node1881 = (inp[13]) ? 4'b0101 : 4'b0001;
														assign node1884 = (inp[15]) ? 4'b0001 : node1885;
															assign node1885 = (inp[13]) ? 4'b1000 : 4'b0000;
													assign node1889 = (inp[13]) ? 4'b1100 : node1890;
														assign node1890 = (inp[15]) ? node1892 : 4'b0000;
															assign node1892 = (inp[14]) ? 4'b0100 : 4'b0000;
											assign node1896 = (inp[2]) ? node1912 : node1897;
												assign node1897 = (inp[15]) ? node1907 : node1898;
													assign node1898 = (inp[4]) ? node1904 : node1899;
														assign node1899 = (inp[7]) ? 4'b1101 : node1900;
															assign node1900 = (inp[13]) ? 4'b1001 : 4'b1101;
														assign node1904 = (inp[7]) ? 4'b1000 : 4'b0000;
													assign node1907 = (inp[13]) ? 4'b1101 : node1908;
														assign node1908 = (inp[4]) ? 4'b1101 : 4'b1001;
												assign node1912 = (inp[15]) ? node1920 : node1913;
													assign node1913 = (inp[4]) ? node1917 : node1914;
														assign node1914 = (inp[7]) ? 4'b0000 : 4'b1000;
														assign node1917 = (inp[13]) ? 4'b1101 : 4'b1001;
													assign node1920 = (inp[13]) ? node1922 : 4'b1100;
														assign node1922 = (inp[14]) ? 4'b0000 : 4'b0100;
										assign node1925 = (inp[12]) ? node1953 : node1926;
											assign node1926 = (inp[4]) ? node1936 : node1927;
												assign node1927 = (inp[15]) ? node1929 : 4'b1001;
													assign node1929 = (inp[2]) ? node1933 : node1930;
														assign node1930 = (inp[7]) ? 4'b1001 : 4'b1101;
														assign node1933 = (inp[7]) ? 4'b1100 : 4'b1000;
												assign node1936 = (inp[2]) ? node1948 : node1937;
													assign node1937 = (inp[13]) ? node1945 : node1938;
														assign node1938 = (inp[14]) ? 4'b0000 : node1939;
															assign node1939 = (inp[15]) ? 4'b1101 : node1940;
																assign node1940 = (inp[7]) ? 4'b0000 : 4'b0100;
														assign node1945 = (inp[15]) ? 4'b1000 : 4'b1100;
													assign node1948 = (inp[15]) ? node1950 : 4'b1101;
														assign node1950 = (inp[7]) ? 4'b0000 : 4'b1001;
											assign node1953 = (inp[2]) ? node1975 : node1954;
												assign node1954 = (inp[4]) ? node1970 : node1955;
													assign node1955 = (inp[15]) ? node1965 : node1956;
														assign node1956 = (inp[14]) ? node1962 : node1957;
															assign node1957 = (inp[13]) ? node1959 : 4'b0001;
																assign node1959 = (inp[7]) ? 4'b0001 : 4'b0000;
															assign node1962 = (inp[13]) ? 4'b0001 : 4'b0101;
														assign node1965 = (inp[13]) ? 4'b0101 : node1966;
															assign node1966 = (inp[7]) ? 4'b0001 : 4'b0101;
													assign node1970 = (inp[13]) ? node1972 : 4'b0101;
														assign node1972 = (inp[15]) ? 4'b0000 : 4'b0100;
												assign node1975 = (inp[4]) ? node1987 : node1976;
													assign node1976 = (inp[15]) ? node1982 : node1977;
														assign node1977 = (inp[14]) ? 4'b0001 : node1978;
															assign node1978 = (inp[7]) ? 4'b0000 : 4'b0001;
														assign node1982 = (inp[13]) ? 4'b1000 : node1983;
															assign node1983 = (inp[7]) ? 4'b0100 : 4'b0000;
													assign node1987 = (inp[15]) ? node1993 : node1988;
														assign node1988 = (inp[7]) ? node1990 : 4'b0101;
															assign node1990 = (inp[13]) ? 4'b0101 : 4'b0001;
														assign node1993 = (inp[13]) ? 4'b0001 : node1994;
															assign node1994 = (inp[7]) ? 4'b0000 : 4'b0001;
								assign node1998 = (inp[10]) ? node2134 : node1999;
									assign node1999 = (inp[3]) ? node2073 : node2000;
										assign node2000 = (inp[2]) ? node2028 : node2001;
											assign node2001 = (inp[4]) ? node2019 : node2002;
												assign node2002 = (inp[15]) ? node2008 : node2003;
													assign node2003 = (inp[13]) ? 4'b0001 : node2004;
														assign node2004 = (inp[7]) ? 4'b1101 : 4'b0001;
													assign node2008 = (inp[7]) ? node2014 : node2009;
														assign node2009 = (inp[12]) ? 4'b1001 : node2010;
															assign node2010 = (inp[13]) ? 4'b1101 : 4'b0101;
														assign node2014 = (inp[13]) ? 4'b1001 : node2015;
															assign node2015 = (inp[14]) ? 4'b1001 : 4'b0001;
												assign node2019 = (inp[15]) ? node2025 : node2020;
													assign node2020 = (inp[13]) ? 4'b0101 : node2021;
														assign node2021 = (inp[7]) ? 4'b0001 : 4'b0101;
													assign node2025 = (inp[13]) ? 4'b0001 : 4'b0101;
											assign node2028 = (inp[15]) ? node2054 : node2029;
												assign node2029 = (inp[7]) ? node2041 : node2030;
													assign node2030 = (inp[4]) ? node2036 : node2031;
														assign node2031 = (inp[12]) ? 4'b1101 : node2032;
															assign node2032 = (inp[13]) ? 4'b1001 : 4'b0001;
														assign node2036 = (inp[12]) ? node2038 : 4'b1001;
															assign node2038 = (inp[13]) ? 4'b0001 : 4'b1001;
													assign node2041 = (inp[4]) ? node2049 : node2042;
														assign node2042 = (inp[14]) ? node2044 : 4'b1101;
															assign node2044 = (inp[12]) ? 4'b0101 : node2045;
																assign node2045 = (inp[13]) ? 4'b1101 : 4'b0101;
														assign node2049 = (inp[12]) ? node2051 : 4'b0001;
															assign node2051 = (inp[13]) ? 4'b0001 : 4'b1101;
												assign node2054 = (inp[7]) ? node2064 : node2055;
													assign node2055 = (inp[12]) ? node2059 : node2056;
														assign node2056 = (inp[13]) ? 4'b1101 : 4'b0101;
														assign node2059 = (inp[13]) ? 4'b0101 : node2060;
															assign node2060 = (inp[4]) ? 4'b1101 : 4'b1001;
													assign node2064 = (inp[4]) ? node2068 : node2065;
														assign node2065 = (inp[12]) ? 4'b0001 : 4'b1001;
														assign node2068 = (inp[14]) ? 4'b1001 : node2069;
															assign node2069 = (inp[13]) ? 4'b1101 : 4'b0101;
										assign node2073 = (inp[15]) ? node2103 : node2074;
											assign node2074 = (inp[4]) ? node2088 : node2075;
												assign node2075 = (inp[14]) ? node2077 : 4'b0001;
													assign node2077 = (inp[12]) ? node2083 : node2078;
														assign node2078 = (inp[13]) ? 4'b0001 : node2079;
															assign node2079 = (inp[2]) ? 4'b0001 : 4'b0101;
														assign node2083 = (inp[13]) ? 4'b0001 : node2084;
															assign node2084 = (inp[2]) ? 4'b1001 : 4'b0001;
												assign node2088 = (inp[2]) ? node2098 : node2089;
													assign node2089 = (inp[13]) ? node2093 : node2090;
														assign node2090 = (inp[7]) ? 4'b0001 : 4'b1001;
														assign node2093 = (inp[12]) ? node2095 : 4'b0101;
															assign node2095 = (inp[7]) ? 4'b1001 : 4'b1101;
													assign node2098 = (inp[7]) ? node2100 : 4'b0101;
														assign node2100 = (inp[13]) ? 4'b0101 : 4'b0001;
											assign node2103 = (inp[4]) ? node2119 : node2104;
												assign node2104 = (inp[2]) ? node2110 : node2105;
													assign node2105 = (inp[13]) ? 4'b0101 : node2106;
														assign node2106 = (inp[7]) ? 4'b0001 : 4'b0101;
													assign node2110 = (inp[12]) ? node2116 : node2111;
														assign node2111 = (inp[13]) ? 4'b1001 : node2112;
															assign node2112 = (inp[7]) ? 4'b0101 : 4'b0001;
														assign node2116 = (inp[13]) ? 4'b0101 : 4'b1101;
												assign node2119 = (inp[13]) ? node2129 : node2120;
													assign node2120 = (inp[7]) ? node2122 : 4'b0001;
														assign node2122 = (inp[12]) ? node2126 : node2123;
															assign node2123 = (inp[2]) ? 4'b0001 : 4'b0101;
															assign node2126 = (inp[2]) ? 4'b1101 : 4'b0101;
													assign node2129 = (inp[7]) ? 4'b0001 : node2130;
														assign node2130 = (inp[2]) ? 4'b0001 : 4'b1001;
									assign node2134 = (inp[13]) ? node2188 : node2135;
										assign node2135 = (inp[2]) ? node2161 : node2136;
											assign node2136 = (inp[15]) ? node2146 : node2137;
												assign node2137 = (inp[7]) ? node2141 : node2138;
													assign node2138 = (inp[4]) ? 4'b1101 : 4'b1001;
													assign node2141 = (inp[4]) ? node2143 : 4'b0101;
														assign node2143 = (inp[3]) ? 4'b0001 : 4'b1001;
												assign node2146 = (inp[3]) ? node2154 : node2147;
													assign node2147 = (inp[4]) ? node2151 : node2148;
														assign node2148 = (inp[7]) ? 4'b0001 : 4'b0101;
														assign node2151 = (inp[7]) ? 4'b0101 : 4'b1001;
													assign node2154 = (inp[7]) ? node2158 : node2155;
														assign node2155 = (inp[4]) ? 4'b0001 : 4'b1101;
														assign node2158 = (inp[4]) ? 4'b1101 : 4'b1001;
											assign node2161 = (inp[3]) ? node2173 : node2162;
												assign node2162 = (inp[15]) ? node2170 : node2163;
													assign node2163 = (inp[12]) ? 4'b0001 : node2164;
														assign node2164 = (inp[4]) ? 4'b0001 : node2165;
															assign node2165 = (inp[7]) ? 4'b0101 : 4'b0001;
													assign node2170 = (inp[7]) ? 4'b0001 : 4'b0101;
												assign node2173 = (inp[7]) ? node2181 : node2174;
													assign node2174 = (inp[12]) ? node2176 : 4'b1001;
														assign node2176 = (inp[14]) ? 4'b0001 : node2177;
															assign node2177 = (inp[4]) ? 4'b1101 : 4'b1001;
													assign node2181 = (inp[4]) ? node2185 : node2182;
														assign node2182 = (inp[15]) ? 4'b0101 : 4'b0001;
														assign node2185 = (inp[15]) ? 4'b0001 : 4'b1001;
										assign node2188 = (inp[4]) ? node2210 : node2189;
											assign node2189 = (inp[15]) ? node2197 : node2190;
												assign node2190 = (inp[3]) ? 4'b1001 : node2191;
													assign node2191 = (inp[14]) ? 4'b1001 : node2192;
														assign node2192 = (inp[7]) ? 4'b1101 : 4'b1001;
												assign node2197 = (inp[2]) ? node2203 : node2198;
													assign node2198 = (inp[3]) ? 4'b1101 : node2199;
														assign node2199 = (inp[7]) ? 4'b1001 : 4'b1101;
													assign node2203 = (inp[7]) ? node2207 : node2204;
														assign node2204 = (inp[3]) ? 4'b1001 : 4'b1101;
														assign node2207 = (inp[3]) ? 4'b1101 : 4'b1001;
											assign node2210 = (inp[15]) ? node2216 : node2211;
												assign node2211 = (inp[2]) ? node2213 : 4'b1101;
													assign node2213 = (inp[3]) ? 4'b1101 : 4'b1001;
												assign node2216 = (inp[2]) ? node2218 : 4'b1001;
													assign node2218 = (inp[3]) ? 4'b1001 : 4'b1101;
						assign node2221 = (inp[15]) ? node2471 : node2222;
							assign node2222 = (inp[2]) ? 4'b1101 : node2223;
								assign node2223 = (inp[13]) ? node2355 : node2224;
									assign node2224 = (inp[10]) ? node2296 : node2225;
										assign node2225 = (inp[12]) ? node2265 : node2226;
											assign node2226 = (inp[1]) ? node2246 : node2227;
												assign node2227 = (inp[14]) ? node2237 : node2228;
													assign node2228 = (inp[4]) ? 4'b0000 : node2229;
														assign node2229 = (inp[7]) ? node2233 : node2230;
															assign node2230 = (inp[11]) ? 4'b0000 : 4'b0100;
															assign node2233 = (inp[3]) ? 4'b0000 : 4'b1101;
													assign node2237 = (inp[11]) ? 4'b0100 : node2238;
														assign node2238 = (inp[3]) ? 4'b1001 : node2239;
															assign node2239 = (inp[7]) ? 4'b1101 : node2240;
																assign node2240 = (inp[4]) ? 4'b1001 : 4'b1101;
												assign node2246 = (inp[11]) ? node2260 : node2247;
													assign node2247 = (inp[4]) ? node2255 : node2248;
														assign node2248 = (inp[14]) ? 4'b1101 : node2249;
															assign node2249 = (inp[3]) ? 4'b0001 : node2250;
																assign node2250 = (inp[7]) ? 4'b1101 : 4'b0001;
														assign node2255 = (inp[3]) ? 4'b0101 : node2256;
															assign node2256 = (inp[14]) ? 4'b0000 : 4'b0001;
													assign node2260 = (inp[3]) ? node2262 : 4'b0001;
														assign node2262 = (inp[4]) ? 4'b0101 : 4'b0001;
											assign node2265 = (inp[3]) ? node2275 : node2266;
												assign node2266 = (inp[7]) ? 4'b1101 : node2267;
													assign node2267 = (inp[4]) ? node2269 : 4'b1101;
														assign node2269 = (inp[14]) ? 4'b1001 : node2270;
															assign node2270 = (inp[1]) ? 4'b1001 : 4'b1000;
												assign node2275 = (inp[1]) ? node2287 : node2276;
													assign node2276 = (inp[11]) ? node2282 : node2277;
														assign node2277 = (inp[14]) ? node2279 : 4'b1000;
															assign node2279 = (inp[7]) ? 4'b1001 : 4'b1101;
														assign node2282 = (inp[7]) ? 4'b1000 : node2283;
															assign node2283 = (inp[4]) ? 4'b1100 : 4'b1000;
													assign node2287 = (inp[11]) ? node2291 : node2288;
														assign node2288 = (inp[14]) ? 4'b1000 : 4'b1001;
														assign node2291 = (inp[7]) ? 4'b1001 : node2292;
															assign node2292 = (inp[4]) ? 4'b1101 : 4'b1001;
										assign node2296 = (inp[3]) ? node2322 : node2297;
											assign node2297 = (inp[7]) ? node2311 : node2298;
												assign node2298 = (inp[1]) ? node2306 : node2299;
													assign node2299 = (inp[11]) ? 4'b0000 : node2300;
														assign node2300 = (inp[14]) ? node2302 : 4'b0000;
															assign node2302 = (inp[12]) ? 4'b1001 : 4'b0001;
													assign node2306 = (inp[14]) ? node2308 : 4'b0001;
														assign node2308 = (inp[11]) ? 4'b0001 : 4'b0000;
												assign node2311 = (inp[4]) ? node2313 : 4'b1101;
													assign node2313 = (inp[11]) ? 4'b0000 : node2314;
														assign node2314 = (inp[14]) ? node2318 : node2315;
															assign node2315 = (inp[1]) ? 4'b0001 : 4'b0000;
															assign node2318 = (inp[1]) ? 4'b0000 : 4'b0001;
											assign node2322 = (inp[4]) ? node2340 : node2323;
												assign node2323 = (inp[7]) ? node2331 : node2324;
													assign node2324 = (inp[12]) ? node2328 : node2325;
														assign node2325 = (inp[1]) ? 4'b0101 : 4'b0100;
														assign node2328 = (inp[14]) ? 4'b1001 : 4'b0101;
													assign node2331 = (inp[14]) ? node2333 : 4'b0001;
														assign node2333 = (inp[1]) ? node2337 : node2334;
															assign node2334 = (inp[11]) ? 4'b0000 : 4'b1001;
															assign node2337 = (inp[11]) ? 4'b0001 : 4'b0000;
												assign node2340 = (inp[1]) ? node2350 : node2341;
													assign node2341 = (inp[11]) ? 4'b0100 : node2342;
														assign node2342 = (inp[14]) ? node2344 : 4'b0100;
															assign node2344 = (inp[12]) ? node2346 : 4'b0101;
																assign node2346 = (inp[7]) ? 4'b1001 : 4'b1101;
													assign node2350 = (inp[14]) ? node2352 : 4'b0101;
														assign node2352 = (inp[11]) ? 4'b0101 : 4'b0100;
									assign node2355 = (inp[3]) ? node2403 : node2356;
										assign node2356 = (inp[7]) ? node2384 : node2357;
											assign node2357 = (inp[1]) ? node2371 : node2358;
												assign node2358 = (inp[11]) ? node2366 : node2359;
													assign node2359 = (inp[14]) ? node2363 : node2360;
														assign node2360 = (inp[12]) ? 4'b0000 : 4'b1000;
														assign node2363 = (inp[10]) ? 4'b1001 : 4'b0001;
													assign node2366 = (inp[12]) ? node2368 : 4'b1000;
														assign node2368 = (inp[10]) ? 4'b1000 : 4'b0000;
												assign node2371 = (inp[14]) ? node2377 : node2372;
													assign node2372 = (inp[10]) ? 4'b1001 : node2373;
														assign node2373 = (inp[12]) ? 4'b0001 : 4'b1001;
													assign node2377 = (inp[11]) ? node2381 : node2378;
														assign node2378 = (inp[12]) ? 4'b0000 : 4'b1000;
														assign node2381 = (inp[12]) ? 4'b0001 : 4'b1001;
											assign node2384 = (inp[4]) ? node2386 : 4'b1101;
												assign node2386 = (inp[10]) ? node2394 : node2387;
													assign node2387 = (inp[12]) ? 4'b0001 : node2388;
														assign node2388 = (inp[1]) ? 4'b1000 : node2389;
															assign node2389 = (inp[14]) ? 4'b0001 : 4'b1000;
													assign node2394 = (inp[14]) ? node2396 : 4'b1000;
														assign node2396 = (inp[11]) ? node2400 : node2397;
															assign node2397 = (inp[1]) ? 4'b1000 : 4'b1001;
															assign node2400 = (inp[1]) ? 4'b1001 : 4'b1000;
										assign node2403 = (inp[1]) ? node2439 : node2404;
											assign node2404 = (inp[14]) ? node2422 : node2405;
												assign node2405 = (inp[7]) ? node2411 : node2406;
													assign node2406 = (inp[12]) ? node2408 : 4'b1100;
														assign node2408 = (inp[10]) ? 4'b1100 : 4'b0100;
													assign node2411 = (inp[4]) ? node2417 : node2412;
														assign node2412 = (inp[10]) ? 4'b1000 : node2413;
															assign node2413 = (inp[12]) ? 4'b0000 : 4'b1000;
														assign node2417 = (inp[12]) ? node2419 : 4'b1100;
															assign node2419 = (inp[10]) ? 4'b1100 : 4'b0100;
												assign node2422 = (inp[11]) ? node2432 : node2423;
													assign node2423 = (inp[12]) ? 4'b0101 : node2424;
														assign node2424 = (inp[10]) ? node2426 : 4'b0101;
															assign node2426 = (inp[4]) ? 4'b1101 : node2427;
																assign node2427 = (inp[7]) ? 4'b1001 : 4'b1101;
													assign node2432 = (inp[10]) ? node2436 : node2433;
														assign node2433 = (inp[12]) ? 4'b0100 : 4'b1100;
														assign node2436 = (inp[7]) ? 4'b1000 : 4'b1100;
											assign node2439 = (inp[14]) ? node2453 : node2440;
												assign node2440 = (inp[12]) ? node2446 : node2441;
													assign node2441 = (inp[4]) ? 4'b1101 : node2442;
														assign node2442 = (inp[10]) ? 4'b1001 : 4'b1101;
													assign node2446 = (inp[10]) ? node2450 : node2447;
														assign node2447 = (inp[4]) ? 4'b0101 : 4'b0001;
														assign node2450 = (inp[7]) ? 4'b1001 : 4'b1101;
												assign node2453 = (inp[11]) ? node2463 : node2454;
													assign node2454 = (inp[7]) ? node2460 : node2455;
														assign node2455 = (inp[12]) ? node2457 : 4'b1100;
															assign node2457 = (inp[4]) ? 4'b1100 : 4'b0100;
														assign node2460 = (inp[4]) ? 4'b1100 : 4'b1000;
													assign node2463 = (inp[10]) ? 4'b1101 : node2464;
														assign node2464 = (inp[12]) ? 4'b0101 : node2465;
															assign node2465 = (inp[4]) ? 4'b1101 : 4'b1001;
							assign node2471 = (inp[2]) ? 4'b1001 : node2472;
								assign node2472 = (inp[3]) ? node2474 : 4'b1001;
									assign node2474 = (inp[4]) ? node2510 : node2475;
										assign node2475 = (inp[7]) ? 4'b1001 : node2476;
											assign node2476 = (inp[13]) ? node2496 : node2477;
												assign node2477 = (inp[10]) ? node2487 : node2478;
													assign node2478 = (inp[12]) ? 4'b1001 : node2479;
														assign node2479 = (inp[1]) ? node2481 : 4'b1001;
															assign node2481 = (inp[11]) ? 4'b0001 : node2482;
																assign node2482 = (inp[14]) ? 4'b0000 : 4'b0001;
													assign node2487 = (inp[1]) ? 4'b0001 : node2488;
														assign node2488 = (inp[14]) ? node2490 : 4'b0000;
															assign node2490 = (inp[11]) ? 4'b0000 : node2491;
																assign node2491 = (inp[12]) ? 4'b1001 : 4'b0001;
												assign node2496 = (inp[1]) ? node2502 : node2497;
													assign node2497 = (inp[10]) ? 4'b1000 : node2498;
														assign node2498 = (inp[12]) ? 4'b0000 : 4'b1000;
													assign node2502 = (inp[14]) ? node2506 : node2503;
														assign node2503 = (inp[12]) ? 4'b0001 : 4'b1001;
														assign node2506 = (inp[11]) ? 4'b1001 : 4'b1000;
										assign node2510 = (inp[1]) ? node2540 : node2511;
											assign node2511 = (inp[14]) ? node2523 : node2512;
												assign node2512 = (inp[13]) ? node2518 : node2513;
													assign node2513 = (inp[12]) ? node2515 : 4'b0000;
														assign node2515 = (inp[10]) ? 4'b0000 : 4'b1000;
													assign node2518 = (inp[12]) ? node2520 : 4'b1000;
														assign node2520 = (inp[10]) ? 4'b1000 : 4'b0000;
												assign node2523 = (inp[11]) ? node2535 : node2524;
													assign node2524 = (inp[13]) ? node2530 : node2525;
														assign node2525 = (inp[7]) ? 4'b1001 : node2526;
															assign node2526 = (inp[10]) ? 4'b0001 : 4'b1001;
														assign node2530 = (inp[12]) ? 4'b0001 : node2531;
															assign node2531 = (inp[10]) ? 4'b1001 : 4'b0001;
													assign node2535 = (inp[13]) ? 4'b1000 : node2536;
														assign node2536 = (inp[12]) ? 4'b1000 : 4'b0000;
											assign node2540 = (inp[13]) ? node2552 : node2541;
												assign node2541 = (inp[11]) ? 4'b0001 : node2542;
													assign node2542 = (inp[14]) ? node2548 : node2543;
														assign node2543 = (inp[12]) ? node2545 : 4'b0001;
															assign node2545 = (inp[10]) ? 4'b0001 : 4'b1001;
														assign node2548 = (inp[7]) ? 4'b1001 : 4'b0000;
												assign node2552 = (inp[10]) ? node2562 : node2553;
													assign node2553 = (inp[12]) ? node2557 : node2554;
														assign node2554 = (inp[14]) ? 4'b1000 : 4'b1001;
														assign node2557 = (inp[11]) ? 4'b0001 : node2558;
															assign node2558 = (inp[14]) ? 4'b0000 : 4'b0001;
													assign node2562 = (inp[11]) ? 4'b1001 : node2563;
														assign node2563 = (inp[14]) ? 4'b1000 : 4'b1001;
					assign node2568 = (inp[3]) ? node3570 : node2569;
						assign node2569 = (inp[4]) ? node3063 : node2570;
							assign node2570 = (inp[0]) ? node2876 : node2571;
								assign node2571 = (inp[11]) ? node2739 : node2572;
									assign node2572 = (inp[2]) ? node2664 : node2573;
										assign node2573 = (inp[10]) ? node2627 : node2574;
											assign node2574 = (inp[14]) ? node2600 : node2575;
												assign node2575 = (inp[1]) ? node2589 : node2576;
													assign node2576 = (inp[12]) ? node2582 : node2577;
														assign node2577 = (inp[7]) ? node2579 : 4'b0101;
															assign node2579 = (inp[13]) ? 4'b1101 : 4'b0001;
														assign node2582 = (inp[7]) ? 4'b1001 : node2583;
															assign node2583 = (inp[15]) ? 4'b0101 : node2584;
																assign node2584 = (inp[13]) ? 4'b1001 : 4'b1101;
													assign node2589 = (inp[12]) ? 4'b0001 : node2590;
														assign node2590 = (inp[13]) ? 4'b1101 : node2591;
															assign node2591 = (inp[7]) ? node2595 : node2592;
																assign node2592 = (inp[15]) ? 4'b1100 : 4'b1001;
																assign node2595 = (inp[15]) ? 4'b1000 : 4'b1100;
												assign node2600 = (inp[1]) ? node2618 : node2601;
													assign node2601 = (inp[15]) ? node2611 : node2602;
														assign node2602 = (inp[12]) ? node2608 : node2603;
															assign node2603 = (inp[7]) ? node2605 : 4'b0001;
																assign node2605 = (inp[13]) ? 4'b0001 : 4'b0100;
															assign node2608 = (inp[7]) ? 4'b1100 : 4'b1001;
														assign node2611 = (inp[7]) ? node2615 : node2612;
															assign node2612 = (inp[12]) ? 4'b1000 : 4'b0100;
															assign node2615 = (inp[12]) ? 4'b0100 : 4'b1100;
													assign node2618 = (inp[13]) ? node2624 : node2619;
														assign node2619 = (inp[15]) ? node2621 : 4'b0101;
															assign node2621 = (inp[7]) ? 4'b0001 : 4'b0101;
														assign node2624 = (inp[12]) ? 4'b0001 : 4'b1001;
											assign node2627 = (inp[15]) ? node2643 : node2628;
												assign node2628 = (inp[13]) ? node2636 : node2629;
													assign node2629 = (inp[7]) ? 4'b0001 : node2630;
														assign node2630 = (inp[1]) ? node2632 : 4'b0001;
															assign node2632 = (inp[12]) ? 4'b0001 : 4'b1001;
													assign node2636 = (inp[7]) ? 4'b0101 : node2637;
														assign node2637 = (inp[12]) ? node2639 : 4'b0101;
															assign node2639 = (inp[14]) ? 4'b0000 : 4'b0001;
												assign node2643 = (inp[13]) ? node2655 : node2644;
													assign node2644 = (inp[1]) ? node2650 : node2645;
														assign node2645 = (inp[7]) ? 4'b1001 : node2646;
															assign node2646 = (inp[14]) ? 4'b1100 : 4'b1101;
														assign node2650 = (inp[14]) ? node2652 : 4'b0100;
															assign node2652 = (inp[12]) ? 4'b1101 : 4'b0101;
													assign node2655 = (inp[1]) ? node2661 : node2656;
														assign node2656 = (inp[12]) ? node2658 : 4'b0001;
															assign node2658 = (inp[7]) ? 4'b0100 : 4'b1001;
														assign node2661 = (inp[12]) ? 4'b0001 : 4'b1001;
										assign node2664 = (inp[15]) ? node2698 : node2665;
											assign node2665 = (inp[13]) ? node2685 : node2666;
												assign node2666 = (inp[7]) ? node2676 : node2667;
													assign node2667 = (inp[12]) ? node2669 : 4'b0001;
														assign node2669 = (inp[10]) ? node2671 : 4'b1100;
															assign node2671 = (inp[14]) ? 4'b1001 : node2672;
																assign node2672 = (inp[1]) ? 4'b0000 : 4'b1001;
													assign node2676 = (inp[1]) ? node2682 : node2677;
														assign node2677 = (inp[12]) ? 4'b0100 : node2678;
															assign node2678 = (inp[10]) ? 4'b1100 : 4'b0100;
														assign node2682 = (inp[10]) ? 4'b0000 : 4'b0100;
												assign node2685 = (inp[14]) ? node2691 : node2686;
													assign node2686 = (inp[1]) ? node2688 : 4'b0001;
														assign node2688 = (inp[7]) ? 4'b1000 : 4'b0100;
													assign node2691 = (inp[1]) ? node2693 : 4'b1000;
														assign node2693 = (inp[7]) ? 4'b1001 : node2694;
															assign node2694 = (inp[10]) ? 4'b1101 : 4'b1001;
											assign node2698 = (inp[10]) ? node2714 : node2699;
												assign node2699 = (inp[1]) ? node2705 : node2700;
													assign node2700 = (inp[7]) ? 4'b1000 : node2701;
														assign node2701 = (inp[13]) ? 4'b1100 : 4'b0100;
													assign node2705 = (inp[7]) ? node2711 : node2706;
														assign node2706 = (inp[12]) ? 4'b0100 : node2707;
															assign node2707 = (inp[14]) ? 4'b0100 : 4'b0000;
														assign node2711 = (inp[13]) ? 4'b0100 : 4'b0000;
												assign node2714 = (inp[12]) ? node2722 : node2715;
													assign node2715 = (inp[7]) ? node2719 : node2716;
														assign node2716 = (inp[13]) ? 4'b1001 : 4'b1100;
														assign node2719 = (inp[13]) ? 4'b1100 : 4'b1000;
													assign node2722 = (inp[1]) ? node2730 : node2723;
														assign node2723 = (inp[7]) ? node2727 : node2724;
															assign node2724 = (inp[13]) ? 4'b0001 : 4'b0100;
															assign node2727 = (inp[13]) ? 4'b0100 : 4'b0000;
														assign node2730 = (inp[14]) ? node2736 : node2731;
															assign node2731 = (inp[7]) ? node2733 : 4'b1100;
																assign node2733 = (inp[13]) ? 4'b1100 : 4'b1000;
															assign node2736 = (inp[13]) ? 4'b0001 : 4'b1100;
									assign node2739 = (inp[1]) ? node2809 : node2740;
										assign node2740 = (inp[2]) ? node2766 : node2741;
											assign node2741 = (inp[13]) ? node2753 : node2742;
												assign node2742 = (inp[15]) ? node2748 : node2743;
													assign node2743 = (inp[7]) ? node2745 : 4'b0001;
														assign node2745 = (inp[10]) ? 4'b0001 : 4'b0100;
													assign node2748 = (inp[7]) ? node2750 : 4'b0100;
														assign node2750 = (inp[10]) ? 4'b1000 : 4'b0000;
												assign node2753 = (inp[15]) ? node2761 : node2754;
													assign node2754 = (inp[7]) ? node2758 : node2755;
														assign node2755 = (inp[10]) ? 4'b0000 : 4'b0101;
														assign node2758 = (inp[10]) ? 4'b0101 : 4'b0001;
													assign node2761 = (inp[10]) ? 4'b0001 : node2762;
														assign node2762 = (inp[7]) ? 4'b1100 : 4'b0001;
											assign node2766 = (inp[15]) ? node2784 : node2767;
												assign node2767 = (inp[13]) ? node2777 : node2768;
													assign node2768 = (inp[12]) ? node2774 : node2769;
														assign node2769 = (inp[7]) ? node2771 : 4'b0000;
															assign node2771 = (inp[14]) ? 4'b0101 : 4'b0000;
														assign node2774 = (inp[10]) ? 4'b0101 : 4'b1101;
													assign node2777 = (inp[10]) ? node2779 : 4'b1000;
														assign node2779 = (inp[12]) ? node2781 : 4'b1000;
															assign node2781 = (inp[7]) ? 4'b0000 : 4'b0100;
												assign node2784 = (inp[13]) ? node2802 : node2785;
													assign node2785 = (inp[7]) ? node2793 : node2786;
														assign node2786 = (inp[10]) ? node2790 : node2787;
															assign node2787 = (inp[12]) ? 4'b1001 : 4'b0101;
															assign node2790 = (inp[12]) ? 4'b0101 : 4'b1101;
														assign node2793 = (inp[14]) ? node2795 : 4'b0001;
															assign node2795 = (inp[10]) ? node2799 : node2796;
																assign node2796 = (inp[12]) ? 4'b1001 : 4'b0001;
																assign node2799 = (inp[12]) ? 4'b0001 : 4'b1001;
													assign node2802 = (inp[10]) ? node2806 : node2803;
														assign node2803 = (inp[12]) ? 4'b1101 : 4'b0101;
														assign node2806 = (inp[7]) ? 4'b0101 : 4'b0000;
										assign node2809 = (inp[2]) ? node2841 : node2810;
											assign node2810 = (inp[13]) ? node2828 : node2811;
												assign node2811 = (inp[15]) ? node2819 : node2812;
													assign node2812 = (inp[10]) ? 4'b1001 : node2813;
														assign node2813 = (inp[7]) ? node2815 : 4'b1001;
															assign node2815 = (inp[12]) ? 4'b0101 : 4'b1101;
													assign node2819 = (inp[10]) ? 4'b0101 : node2820;
														assign node2820 = (inp[14]) ? node2824 : node2821;
															assign node2821 = (inp[12]) ? 4'b0001 : 4'b1001;
															assign node2824 = (inp[12]) ? 4'b0101 : 4'b1101;
												assign node2828 = (inp[15]) ? node2836 : node2829;
													assign node2829 = (inp[7]) ? node2833 : node2830;
														assign node2830 = (inp[10]) ? 4'b1001 : 4'b1101;
														assign node2833 = (inp[10]) ? 4'b1101 : 4'b1001;
													assign node2836 = (inp[10]) ? 4'b1001 : node2837;
														assign node2837 = (inp[7]) ? 4'b0101 : 4'b1001;
											assign node2841 = (inp[10]) ? node2863 : node2842;
												assign node2842 = (inp[15]) ? node2852 : node2843;
													assign node2843 = (inp[7]) ? 4'b0101 : node2844;
														assign node2844 = (inp[14]) ? 4'b1001 : node2845;
															assign node2845 = (inp[13]) ? 4'b0101 : node2846;
																assign node2846 = (inp[12]) ? 4'b0001 : 4'b1001;
													assign node2852 = (inp[12]) ? 4'b0101 : node2853;
														assign node2853 = (inp[14]) ? node2855 : 4'b0101;
															assign node2855 = (inp[13]) ? node2859 : node2856;
																assign node2856 = (inp[7]) ? 4'b0001 : 4'b0101;
																assign node2859 = (inp[7]) ? 4'b0101 : 4'b0001;
												assign node2863 = (inp[15]) ? node2869 : node2864;
													assign node2864 = (inp[13]) ? node2866 : 4'b0001;
														assign node2866 = (inp[7]) ? 4'b1001 : 4'b1101;
													assign node2869 = (inp[7]) ? node2873 : node2870;
														assign node2870 = (inp[13]) ? 4'b1001 : 4'b1101;
														assign node2873 = (inp[14]) ? 4'b1101 : 4'b1001;
								assign node2876 = (inp[2]) ? node3032 : node2877;
									assign node2877 = (inp[7]) ? node2959 : node2878;
										assign node2878 = (inp[15]) ? node2906 : node2879;
											assign node2879 = (inp[11]) ? node2891 : node2880;
												assign node2880 = (inp[10]) ? node2884 : node2881;
													assign node2881 = (inp[14]) ? 4'b1101 : 4'b0000;
													assign node2884 = (inp[13]) ? 4'b1000 : node2885;
														assign node2885 = (inp[12]) ? node2887 : 4'b1000;
															assign node2887 = (inp[1]) ? 4'b1000 : 4'b0000;
												assign node2891 = (inp[1]) ? node2903 : node2892;
													assign node2892 = (inp[14]) ? node2894 : 4'b1001;
														assign node2894 = (inp[10]) ? node2900 : node2895;
															assign node2895 = (inp[12]) ? node2897 : 4'b0001;
																assign node2897 = (inp[13]) ? 4'b1001 : 4'b1100;
															assign node2900 = (inp[12]) ? 4'b0001 : 4'b1001;
													assign node2903 = (inp[10]) ? 4'b1001 : 4'b0001;
											assign node2906 = (inp[13]) ? node2932 : node2907;
												assign node2907 = (inp[10]) ? node2923 : node2908;
													assign node2908 = (inp[12]) ? node2918 : node2909;
														assign node2909 = (inp[14]) ? node2913 : node2910;
															assign node2910 = (inp[1]) ? 4'b0101 : 4'b0100;
															assign node2913 = (inp[1]) ? node2915 : 4'b1001;
																assign node2915 = (inp[11]) ? 4'b0101 : 4'b0100;
														assign node2918 = (inp[11]) ? 4'b1000 : node2919;
															assign node2919 = (inp[1]) ? 4'b1000 : 4'b1001;
													assign node2923 = (inp[11]) ? 4'b0101 : node2924;
														assign node2924 = (inp[14]) ? node2928 : node2925;
															assign node2925 = (inp[1]) ? 4'b0101 : 4'b0100;
															assign node2928 = (inp[1]) ? 4'b0100 : 4'b0101;
												assign node2932 = (inp[12]) ? node2944 : node2933;
													assign node2933 = (inp[1]) ? node2939 : node2934;
														assign node2934 = (inp[14]) ? node2936 : 4'b1100;
															assign node2936 = (inp[11]) ? 4'b1100 : 4'b0101;
														assign node2939 = (inp[14]) ? node2941 : 4'b1101;
															assign node2941 = (inp[11]) ? 4'b1101 : 4'b1100;
													assign node2944 = (inp[10]) ? node2950 : node2945;
														assign node2945 = (inp[1]) ? node2947 : 4'b0100;
															assign node2947 = (inp[14]) ? 4'b0100 : 4'b0101;
														assign node2950 = (inp[1]) ? node2954 : node2951;
															assign node2951 = (inp[14]) ? 4'b0101 : 4'b1100;
															assign node2954 = (inp[11]) ? 4'b1101 : node2955;
																assign node2955 = (inp[14]) ? 4'b1100 : 4'b1101;
										assign node2959 = (inp[15]) ? node2991 : node2960;
											assign node2960 = (inp[13]) ? node2976 : node2961;
												assign node2961 = (inp[1]) ? node2967 : node2962;
													assign node2962 = (inp[12]) ? node2964 : 4'b0100;
														assign node2964 = (inp[10]) ? 4'b0100 : 4'b1100;
													assign node2967 = (inp[10]) ? node2973 : node2968;
														assign node2968 = (inp[12]) ? node2970 : 4'b0101;
															assign node2970 = (inp[11]) ? 4'b1101 : 4'b1100;
														assign node2973 = (inp[14]) ? 4'b0100 : 4'b0101;
												assign node2976 = (inp[11]) ? node2988 : node2977;
													assign node2977 = (inp[10]) ? node2983 : node2978;
														assign node2978 = (inp[1]) ? 4'b0000 : node2979;
															assign node2979 = (inp[14]) ? 4'b0000 : 4'b0100;
														assign node2983 = (inp[1]) ? 4'b1000 : node2984;
															assign node2984 = (inp[12]) ? 4'b0000 : 4'b1000;
													assign node2988 = (inp[10]) ? 4'b1001 : 4'b0001;
											assign node2991 = (inp[1]) ? node3015 : node2992;
												assign node2992 = (inp[14]) ? node3000 : node2993;
													assign node2993 = (inp[13]) ? node2997 : node2994;
														assign node2994 = (inp[10]) ? 4'b0000 : 4'b1000;
														assign node2997 = (inp[10]) ? 4'b1000 : 4'b0000;
													assign node3000 = (inp[11]) ? node3008 : node3001;
														assign node3001 = (inp[10]) ? node3003 : 4'b0001;
															assign node3003 = (inp[12]) ? node3005 : 4'b1001;
																assign node3005 = (inp[13]) ? 4'b0001 : 4'b1001;
														assign node3008 = (inp[12]) ? node3010 : 4'b0000;
															assign node3010 = (inp[10]) ? 4'b0000 : node3011;
																assign node3011 = (inp[13]) ? 4'b0000 : 4'b1000;
												assign node3015 = (inp[11]) ? node3027 : node3016;
													assign node3016 = (inp[14]) ? node3022 : node3017;
														assign node3017 = (inp[13]) ? 4'b1001 : node3018;
															assign node3018 = (inp[10]) ? 4'b0001 : 4'b1001;
														assign node3022 = (inp[13]) ? 4'b1000 : node3023;
															assign node3023 = (inp[10]) ? 4'b0000 : 4'b1000;
													assign node3027 = (inp[13]) ? node3029 : 4'b0001;
														assign node3029 = (inp[12]) ? 4'b0001 : 4'b1001;
									assign node3032 = (inp[15]) ? 4'b1001 : node3033;
										assign node3033 = (inp[7]) ? 4'b1101 : node3034;
											assign node3034 = (inp[13]) ? node3046 : node3035;
												assign node3035 = (inp[12]) ? 4'b1101 : node3036;
													assign node3036 = (inp[1]) ? node3042 : node3037;
														assign node3037 = (inp[14]) ? node3039 : 4'b0000;
															assign node3039 = (inp[10]) ? 4'b0001 : 4'b1101;
														assign node3042 = (inp[14]) ? 4'b0000 : 4'b0001;
												assign node3046 = (inp[1]) ? node3054 : node3047;
													assign node3047 = (inp[14]) ? 4'b0000 : node3048;
														assign node3048 = (inp[12]) ? node3050 : 4'b1000;
															assign node3050 = (inp[10]) ? 4'b1000 : 4'b0000;
													assign node3054 = (inp[10]) ? 4'b1001 : node3055;
														assign node3055 = (inp[12]) ? 4'b0001 : node3056;
															assign node3056 = (inp[11]) ? 4'b1001 : 4'b1000;
							assign node3063 = (inp[2]) ? node3363 : node3064;
								assign node3064 = (inp[11]) ? node3246 : node3065;
									assign node3065 = (inp[0]) ? node3153 : node3066;
										assign node3066 = (inp[13]) ? node3124 : node3067;
											assign node3067 = (inp[15]) ? node3093 : node3068;
												assign node3068 = (inp[10]) ? node3078 : node3069;
													assign node3069 = (inp[1]) ? node3075 : node3070;
														assign node3070 = (inp[14]) ? node3072 : 4'b0000;
															assign node3072 = (inp[12]) ? 4'b1001 : 4'b0001;
														assign node3075 = (inp[14]) ? 4'b1000 : 4'b1001;
													assign node3078 = (inp[7]) ? node3084 : node3079;
														assign node3079 = (inp[14]) ? 4'b0101 : node3080;
															assign node3080 = (inp[12]) ? 4'b0100 : 4'b1100;
														assign node3084 = (inp[1]) ? node3088 : node3085;
															assign node3085 = (inp[14]) ? 4'b0001 : 4'b1000;
															assign node3088 = (inp[12]) ? 4'b1000 : node3089;
																assign node3089 = (inp[14]) ? 4'b0100 : 4'b0101;
												assign node3093 = (inp[7]) ? node3111 : node3094;
													assign node3094 = (inp[10]) ? node3102 : node3095;
														assign node3095 = (inp[14]) ? 4'b1001 : node3096;
															assign node3096 = (inp[12]) ? node3098 : 4'b0101;
																assign node3098 = (inp[1]) ? 4'b0101 : 4'b1001;
														assign node3102 = (inp[1]) ? node3106 : node3103;
															assign node3103 = (inp[12]) ? 4'b0001 : 4'b1000;
															assign node3106 = (inp[12]) ? node3108 : 4'b0001;
																assign node3108 = (inp[14]) ? 4'b1000 : 4'b1001;
													assign node3111 = (inp[10]) ? node3117 : node3112;
														assign node3112 = (inp[14]) ? 4'b0001 : node3113;
															assign node3113 = (inp[12]) ? 4'b0001 : 4'b1001;
														assign node3117 = (inp[12]) ? node3121 : node3118;
															assign node3118 = (inp[1]) ? 4'b0001 : 4'b0101;
															assign node3121 = (inp[1]) ? 4'b0101 : 4'b1001;
											assign node3124 = (inp[1]) ? node3142 : node3125;
												assign node3125 = (inp[14]) ? node3139 : node3126;
													assign node3126 = (inp[15]) ? node3134 : node3127;
														assign node3127 = (inp[7]) ? node3131 : node3128;
															assign node3128 = (inp[12]) ? 4'b0001 : 4'b1001;
															assign node3131 = (inp[10]) ? 4'b1000 : 4'b0000;
														assign node3134 = (inp[10]) ? node3136 : 4'b1000;
															assign node3136 = (inp[12]) ? 4'b1000 : 4'b0100;
													assign node3139 = (inp[15]) ? 4'b1001 : 4'b1000;
												assign node3142 = (inp[7]) ? node3148 : node3143;
													assign node3143 = (inp[10]) ? node3145 : 4'b0101;
														assign node3145 = (inp[12]) ? 4'b0000 : 4'b0001;
													assign node3148 = (inp[14]) ? 4'b0000 : node3149;
														assign node3149 = (inp[15]) ? 4'b0001 : 4'b1000;
										assign node3153 = (inp[10]) ? node3199 : node3154;
											assign node3154 = (inp[1]) ? node3182 : node3155;
												assign node3155 = (inp[12]) ? node3169 : node3156;
													assign node3156 = (inp[13]) ? node3164 : node3157;
														assign node3157 = (inp[14]) ? 4'b0000 : node3158;
															assign node3158 = (inp[15]) ? 4'b0000 : node3159;
																assign node3159 = (inp[7]) ? 4'b0000 : 4'b0100;
														assign node3164 = (inp[14]) ? 4'b0100 : node3165;
															assign node3165 = (inp[15]) ? 4'b0000 : 4'b1001;
													assign node3169 = (inp[13]) ? node3175 : node3170;
														assign node3170 = (inp[7]) ? 4'b1000 : node3171;
															assign node3171 = (inp[15]) ? 4'b1100 : 4'b1000;
														assign node3175 = (inp[7]) ? 4'b1000 : node3176;
															assign node3176 = (inp[15]) ? 4'b1000 : node3177;
																assign node3177 = (inp[14]) ? 4'b0000 : 4'b0001;
												assign node3182 = (inp[15]) ? node3194 : node3183;
													assign node3183 = (inp[7]) ? node3189 : node3184;
														assign node3184 = (inp[13]) ? node3186 : 4'b0100;
															assign node3186 = (inp[14]) ? 4'b1001 : 4'b0000;
														assign node3189 = (inp[13]) ? node3191 : 4'b0000;
															assign node3191 = (inp[14]) ? 4'b0100 : 4'b0000;
													assign node3194 = (inp[13]) ? 4'b0000 : node3195;
														assign node3195 = (inp[7]) ? 4'b1000 : 4'b0000;
											assign node3199 = (inp[1]) ? node3225 : node3200;
												assign node3200 = (inp[12]) ? node3210 : node3201;
													assign node3201 = (inp[13]) ? node3207 : node3202;
														assign node3202 = (inp[7]) ? 4'b0101 : node3203;
															assign node3203 = (inp[14]) ? 4'b1000 : 4'b1100;
														assign node3207 = (inp[15]) ? 4'b1000 : 4'b0000;
													assign node3210 = (inp[7]) ? node3220 : node3211;
														assign node3211 = (inp[13]) ? node3215 : node3212;
															assign node3212 = (inp[15]) ? 4'b0000 : 4'b0100;
															assign node3215 = (inp[14]) ? 4'b0000 : node3216;
																assign node3216 = (inp[15]) ? 4'b0000 : 4'b0001;
														assign node3220 = (inp[15]) ? 4'b1001 : node3221;
															assign node3221 = (inp[14]) ? 4'b0000 : 4'b0001;
												assign node3225 = (inp[13]) ? node3239 : node3226;
													assign node3226 = (inp[12]) ? node3234 : node3227;
														assign node3227 = (inp[7]) ? 4'b1000 : node3228;
															assign node3228 = (inp[15]) ? 4'b1000 : node3229;
																assign node3229 = (inp[14]) ? 4'b0001 : 4'b0000;
														assign node3234 = (inp[7]) ? 4'b0101 : node3235;
															assign node3235 = (inp[15]) ? 4'b1000 : 4'b1100;
													assign node3239 = (inp[12]) ? 4'b1000 : node3240;
														assign node3240 = (inp[14]) ? node3242 : 4'b1000;
															assign node3242 = (inp[15]) ? 4'b1000 : 4'b1001;
									assign node3246 = (inp[1]) ? node3318 : node3247;
										assign node3247 = (inp[15]) ? node3287 : node3248;
											assign node3248 = (inp[10]) ? node3262 : node3249;
												assign node3249 = (inp[13]) ? node3257 : node3250;
													assign node3250 = (inp[0]) ? node3254 : node3251;
														assign node3251 = (inp[12]) ? 4'b0000 : 4'b1000;
														assign node3254 = (inp[7]) ? 4'b0001 : 4'b1001;
													assign node3257 = (inp[12]) ? node3259 : 4'b1001;
														assign node3259 = (inp[14]) ? 4'b1001 : 4'b0001;
												assign node3262 = (inp[13]) ? node3272 : node3263;
													assign node3263 = (inp[0]) ? node3269 : node3264;
														assign node3264 = (inp[7]) ? 4'b1000 : node3265;
															assign node3265 = (inp[12]) ? 4'b1100 : 4'b0001;
														assign node3269 = (inp[12]) ? 4'b0001 : 4'b1001;
													assign node3272 = (inp[7]) ? node3280 : node3273;
														assign node3273 = (inp[12]) ? node3277 : node3274;
															assign node3274 = (inp[0]) ? 4'b1000 : 4'b0000;
															assign node3277 = (inp[0]) ? 4'b0000 : 4'b1000;
														assign node3280 = (inp[12]) ? node3284 : node3281;
															assign node3281 = (inp[0]) ? 4'b1000 : 4'b0000;
															assign node3284 = (inp[0]) ? 4'b0000 : 4'b1001;
											assign node3287 = (inp[12]) ? node3303 : node3288;
												assign node3288 = (inp[10]) ? node3298 : node3289;
													assign node3289 = (inp[13]) ? 4'b0001 : node3290;
														assign node3290 = (inp[7]) ? node3294 : node3291;
															assign node3291 = (inp[0]) ? 4'b0001 : 4'b0101;
															assign node3294 = (inp[0]) ? 4'b0100 : 4'b0001;
													assign node3298 = (inp[0]) ? 4'b1001 : node3299;
														assign node3299 = (inp[13]) ? 4'b0001 : 4'b1000;
												assign node3303 = (inp[13]) ? node3311 : node3304;
													assign node3304 = (inp[7]) ? node3306 : 4'b1000;
														assign node3306 = (inp[0]) ? 4'b1000 : node3307;
															assign node3307 = (inp[10]) ? 4'b0101 : 4'b0001;
													assign node3311 = (inp[0]) ? node3315 : node3312;
														assign node3312 = (inp[10]) ? 4'b0100 : 4'b1000;
														assign node3315 = (inp[10]) ? 4'b0001 : 4'b0100;
										assign node3318 = (inp[10]) ? node3348 : node3319;
											assign node3319 = (inp[13]) ? node3339 : node3320;
												assign node3320 = (inp[12]) ? node3328 : node3321;
													assign node3321 = (inp[15]) ? node3325 : node3322;
														assign node3322 = (inp[7]) ? 4'b0001 : 4'b0101;
														assign node3325 = (inp[7]) ? 4'b1001 : 4'b0001;
													assign node3328 = (inp[0]) ? node3334 : node3329;
														assign node3329 = (inp[15]) ? node3331 : 4'b1001;
															assign node3331 = (inp[7]) ? 4'b1001 : 4'b1101;
														assign node3334 = (inp[15]) ? 4'b1001 : node3335;
															assign node3335 = (inp[14]) ? 4'b0001 : 4'b0101;
												assign node3339 = (inp[15]) ? node3341 : 4'b0001;
													assign node3341 = (inp[0]) ? 4'b0001 : node3342;
														assign node3342 = (inp[12]) ? 4'b0001 : node3343;
															assign node3343 = (inp[7]) ? 4'b1001 : 4'b0001;
											assign node3348 = (inp[13]) ? 4'b1001 : node3349;
												assign node3349 = (inp[0]) ? node3355 : node3350;
													assign node3350 = (inp[15]) ? 4'b0001 : node3351;
														assign node3351 = (inp[7]) ? 4'b0101 : 4'b1001;
													assign node3355 = (inp[7]) ? node3359 : node3356;
														assign node3356 = (inp[15]) ? 4'b1001 : 4'b0001;
														assign node3359 = (inp[15]) ? 4'b0101 : 4'b1001;
								assign node3363 = (inp[0]) ? node3517 : node3364;
									assign node3364 = (inp[1]) ? node3440 : node3365;
										assign node3365 = (inp[11]) ? node3411 : node3366;
											assign node3366 = (inp[12]) ? node3390 : node3367;
												assign node3367 = (inp[15]) ? node3375 : node3368;
													assign node3368 = (inp[13]) ? node3370 : 4'b0001;
														assign node3370 = (inp[14]) ? 4'b0101 : node3371;
															assign node3371 = (inp[10]) ? 4'b0000 : 4'b0101;
													assign node3375 = (inp[14]) ? node3385 : node3376;
														assign node3376 = (inp[10]) ? node3382 : node3377;
															assign node3377 = (inp[13]) ? node3379 : 4'b0001;
																assign node3379 = (inp[7]) ? 4'b1001 : 4'b0001;
															assign node3382 = (inp[13]) ? 4'b0001 : 4'b1001;
														assign node3385 = (inp[10]) ? 4'b0001 : node3386;
															assign node3386 = (inp[13]) ? 4'b1000 : 4'b0000;
												assign node3390 = (inp[7]) ? node3400 : node3391;
													assign node3391 = (inp[10]) ? node3395 : node3392;
														assign node3392 = (inp[15]) ? 4'b1001 : 4'b1101;
														assign node3395 = (inp[14]) ? 4'b1001 : node3396;
															assign node3396 = (inp[13]) ? 4'b1000 : 4'b1001;
													assign node3400 = (inp[15]) ? node3404 : node3401;
														assign node3401 = (inp[13]) ? 4'b1001 : 4'b1100;
														assign node3404 = (inp[10]) ? node3408 : node3405;
															assign node3405 = (inp[14]) ? 4'b0000 : 4'b0001;
															assign node3408 = (inp[14]) ? 4'b0100 : 4'b0101;
											assign node3411 = (inp[7]) ? node3425 : node3412;
												assign node3412 = (inp[15]) ? node3420 : node3413;
													assign node3413 = (inp[13]) ? node3415 : 4'b0001;
														assign node3415 = (inp[10]) ? 4'b0000 : node3416;
															assign node3416 = (inp[12]) ? 4'b0101 : 4'b0000;
													assign node3420 = (inp[13]) ? 4'b0001 : node3421;
														assign node3421 = (inp[10]) ? 4'b0100 : 4'b0000;
												assign node3425 = (inp[13]) ? node3433 : node3426;
													assign node3426 = (inp[15]) ? node3428 : 4'b0100;
														assign node3428 = (inp[10]) ? node3430 : 4'b0000;
															assign node3430 = (inp[12]) ? 4'b1000 : 4'b0000;
													assign node3433 = (inp[10]) ? node3437 : node3434;
														assign node3434 = (inp[15]) ? 4'b1000 : 4'b0001;
														assign node3437 = (inp[15]) ? 4'b0001 : 4'b0000;
										assign node3440 = (inp[12]) ? node3478 : node3441;
											assign node3441 = (inp[15]) ? node3459 : node3442;
												assign node3442 = (inp[10]) ? node3452 : node3443;
													assign node3443 = (inp[7]) ? node3447 : node3444;
														assign node3444 = (inp[13]) ? 4'b0001 : 4'b1001;
														assign node3447 = (inp[13]) ? 4'b1001 : node3448;
															assign node3448 = (inp[11]) ? 4'b1101 : 4'b0101;
													assign node3452 = (inp[11]) ? 4'b1001 : node3453;
														assign node3453 = (inp[13]) ? node3455 : 4'b1001;
															assign node3455 = (inp[14]) ? 4'b1000 : 4'b1001;
												assign node3459 = (inp[14]) ? node3471 : node3460;
													assign node3460 = (inp[11]) ? node3468 : node3461;
														assign node3461 = (inp[7]) ? 4'b0100 : node3462;
															assign node3462 = (inp[13]) ? 4'b1001 : node3463;
																assign node3463 = (inp[10]) ? 4'b0100 : 4'b1000;
														assign node3468 = (inp[10]) ? 4'b0101 : 4'b1001;
													assign node3471 = (inp[13]) ? 4'b1001 : node3472;
														assign node3472 = (inp[11]) ? node3474 : 4'b0001;
															assign node3474 = (inp[10]) ? 4'b0001 : 4'b1001;
											assign node3478 = (inp[11]) ? node3508 : node3479;
												assign node3479 = (inp[13]) ? node3497 : node3480;
													assign node3480 = (inp[14]) ? node3488 : node3481;
														assign node3481 = (inp[10]) ? 4'b0100 : node3482;
															assign node3482 = (inp[7]) ? 4'b0100 : node3483;
																assign node3483 = (inp[15]) ? 4'b0000 : 4'b0001;
														assign node3488 = (inp[15]) ? node3494 : node3489;
															assign node3489 = (inp[10]) ? 4'b0001 : node3490;
																assign node3490 = (inp[7]) ? 4'b0101 : 4'b0001;
															assign node3494 = (inp[10]) ? 4'b1001 : 4'b0001;
													assign node3497 = (inp[14]) ? node3505 : node3498;
														assign node3498 = (inp[10]) ? 4'b0001 : node3499;
															assign node3499 = (inp[7]) ? node3501 : 4'b0001;
																assign node3501 = (inp[15]) ? 4'b1000 : 4'b0001;
														assign node3505 = (inp[15]) ? 4'b0001 : 4'b0000;
												assign node3508 = (inp[13]) ? 4'b1001 : node3509;
													assign node3509 = (inp[10]) ? node3513 : node3510;
														assign node3510 = (inp[15]) ? 4'b0001 : 4'b0101;
														assign node3513 = (inp[7]) ? 4'b1001 : 4'b0101;
									assign node3517 = (inp[15]) ? 4'b1001 : node3518;
										assign node3518 = (inp[13]) ? node3542 : node3519;
											assign node3519 = (inp[12]) ? node3531 : node3520;
												assign node3520 = (inp[1]) ? node3526 : node3521;
													assign node3521 = (inp[11]) ? 4'b0000 : node3522;
														assign node3522 = (inp[10]) ? 4'b0001 : 4'b0000;
													assign node3526 = (inp[14]) ? node3528 : 4'b0001;
														assign node3528 = (inp[11]) ? 4'b0001 : 4'b0000;
												assign node3531 = (inp[10]) ? node3537 : node3532;
													assign node3532 = (inp[7]) ? 4'b1101 : node3533;
														assign node3533 = (inp[14]) ? 4'b1000 : 4'b1001;
													assign node3537 = (inp[14]) ? 4'b0000 : node3538;
														assign node3538 = (inp[1]) ? 4'b0001 : 4'b0000;
											assign node3542 = (inp[12]) ? node3556 : node3543;
												assign node3543 = (inp[1]) ? node3551 : node3544;
													assign node3544 = (inp[14]) ? node3546 : 4'b1000;
														assign node3546 = (inp[11]) ? 4'b1000 : node3547;
															assign node3547 = (inp[10]) ? 4'b1001 : 4'b0001;
													assign node3551 = (inp[11]) ? 4'b1001 : node3552;
														assign node3552 = (inp[14]) ? 4'b1000 : 4'b1001;
												assign node3556 = (inp[10]) ? node3562 : node3557;
													assign node3557 = (inp[7]) ? 4'b0001 : node3558;
														assign node3558 = (inp[1]) ? 4'b0001 : 4'b0000;
													assign node3562 = (inp[11]) ? 4'b1000 : node3563;
														assign node3563 = (inp[1]) ? node3565 : 4'b0001;
															assign node3565 = (inp[14]) ? 4'b1000 : 4'b1001;
						assign node3570 = (inp[4]) ? node4172 : node3571;
							assign node3571 = (inp[11]) ? node3939 : node3572;
								assign node3572 = (inp[0]) ? node3770 : node3573;
									assign node3573 = (inp[7]) ? node3677 : node3574;
										assign node3574 = (inp[12]) ? node3632 : node3575;
											assign node3575 = (inp[14]) ? node3607 : node3576;
												assign node3576 = (inp[1]) ? node3586 : node3577;
													assign node3577 = (inp[10]) ? node3583 : node3578;
														assign node3578 = (inp[2]) ? 4'b0000 : node3579;
															assign node3579 = (inp[13]) ? 4'b0000 : 4'b0001;
														assign node3583 = (inp[2]) ? 4'b0000 : 4'b1000;
													assign node3586 = (inp[2]) ? node3596 : node3587;
														assign node3587 = (inp[13]) ? node3593 : node3588;
															assign node3588 = (inp[10]) ? 4'b0001 : node3589;
																assign node3589 = (inp[15]) ? 4'b0000 : 4'b0001;
															assign node3593 = (inp[15]) ? 4'b0001 : 4'b0000;
														assign node3596 = (inp[15]) ? node3600 : node3597;
															assign node3597 = (inp[13]) ? 4'b0001 : 4'b0000;
															assign node3600 = (inp[13]) ? node3604 : node3601;
																assign node3601 = (inp[10]) ? 4'b1000 : 4'b1001;
																assign node3604 = (inp[10]) ? 4'b0001 : 4'b1000;
												assign node3607 = (inp[1]) ? node3619 : node3608;
													assign node3608 = (inp[10]) ? 4'b0001 : node3609;
														assign node3609 = (inp[13]) ? 4'b0000 : node3610;
															assign node3610 = (inp[15]) ? node3614 : node3611;
																assign node3611 = (inp[2]) ? 4'b0000 : 4'b0001;
																assign node3614 = (inp[2]) ? 4'b0001 : 4'b0000;
													assign node3619 = (inp[10]) ? node3623 : node3620;
														assign node3620 = (inp[13]) ? 4'b0000 : 4'b1000;
														assign node3623 = (inp[13]) ? node3627 : node3624;
															assign node3624 = (inp[15]) ? 4'b0001 : 4'b0000;
															assign node3627 = (inp[2]) ? node3629 : 4'b0000;
																assign node3629 = (inp[15]) ? 4'b0000 : 4'b0001;
											assign node3632 = (inp[10]) ? node3656 : node3633;
												assign node3633 = (inp[1]) ? node3647 : node3634;
													assign node3634 = (inp[14]) ? 4'b0000 : node3635;
														assign node3635 = (inp[15]) ? node3641 : node3636;
															assign node3636 = (inp[13]) ? node3638 : 4'b0000;
																assign node3638 = (inp[2]) ? 4'b0001 : 4'b0000;
															assign node3641 = (inp[13]) ? node3643 : 4'b0001;
																assign node3643 = (inp[2]) ? 4'b0000 : 4'b1000;
													assign node3647 = (inp[14]) ? 4'b1000 : node3648;
														assign node3648 = (inp[2]) ? node3652 : node3649;
															assign node3649 = (inp[13]) ? 4'b1000 : 4'b0000;
															assign node3652 = (inp[15]) ? 4'b1001 : 4'b0001;
												assign node3656 = (inp[15]) ? node3664 : node3657;
													assign node3657 = (inp[13]) ? 4'b0000 : node3658;
														assign node3658 = (inp[2]) ? 4'b1000 : node3659;
															assign node3659 = (inp[1]) ? 4'b0000 : 4'b1000;
													assign node3664 = (inp[2]) ? node3668 : node3665;
														assign node3665 = (inp[13]) ? 4'b1000 : 4'b0001;
														assign node3668 = (inp[1]) ? node3672 : node3669;
															assign node3669 = (inp[14]) ? 4'b0001 : 4'b0000;
															assign node3672 = (inp[13]) ? node3674 : 4'b0000;
																assign node3674 = (inp[14]) ? 4'b0000 : 4'b0001;
										assign node3677 = (inp[12]) ? node3721 : node3678;
											assign node3678 = (inp[15]) ? node3704 : node3679;
												assign node3679 = (inp[13]) ? node3691 : node3680;
													assign node3680 = (inp[2]) ? node3688 : node3681;
														assign node3681 = (inp[10]) ? 4'b1001 : node3682;
															assign node3682 = (inp[1]) ? 4'b0001 : node3683;
																assign node3683 = (inp[14]) ? 4'b0000 : 4'b0001;
														assign node3688 = (inp[1]) ? 4'b0000 : 4'b0001;
													assign node3691 = (inp[10]) ? node3699 : node3692;
														assign node3692 = (inp[14]) ? 4'b1000 : node3693;
															assign node3693 = (inp[2]) ? node3695 : 4'b1000;
																assign node3695 = (inp[1]) ? 4'b0001 : 4'b1001;
														assign node3699 = (inp[1]) ? 4'b0000 : node3700;
															assign node3700 = (inp[14]) ? 4'b0001 : 4'b0000;
												assign node3704 = (inp[2]) ? node3716 : node3705;
													assign node3705 = (inp[1]) ? node3711 : node3706;
														assign node3706 = (inp[13]) ? node3708 : 4'b0000;
															assign node3708 = (inp[14]) ? 4'b0001 : 4'b0000;
														assign node3711 = (inp[13]) ? 4'b0001 : node3712;
															assign node3712 = (inp[14]) ? 4'b0001 : 4'b0000;
													assign node3716 = (inp[13]) ? node3718 : 4'b0001;
														assign node3718 = (inp[1]) ? 4'b0001 : 4'b0000;
											assign node3721 = (inp[2]) ? node3741 : node3722;
												assign node3722 = (inp[10]) ? node3734 : node3723;
													assign node3723 = (inp[1]) ? node3729 : node3724;
														assign node3724 = (inp[14]) ? node3726 : 4'b0001;
															assign node3726 = (inp[15]) ? 4'b0001 : 4'b0000;
														assign node3729 = (inp[13]) ? 4'b1001 : node3730;
															assign node3730 = (inp[15]) ? 4'b0000 : 4'b0001;
													assign node3734 = (inp[14]) ? node3736 : 4'b1001;
														assign node3736 = (inp[15]) ? 4'b1000 : node3737;
															assign node3737 = (inp[1]) ? 4'b1000 : 4'b0001;
												assign node3741 = (inp[10]) ? node3757 : node3742;
													assign node3742 = (inp[13]) ? node3750 : node3743;
														assign node3743 = (inp[1]) ? 4'b0001 : node3744;
															assign node3744 = (inp[14]) ? 4'b1001 : node3745;
																assign node3745 = (inp[15]) ? 4'b1001 : 4'b0000;
														assign node3750 = (inp[15]) ? node3754 : node3751;
															assign node3751 = (inp[1]) ? 4'b0001 : 4'b1000;
															assign node3754 = (inp[1]) ? 4'b1000 : 4'b0000;
													assign node3757 = (inp[13]) ? node3763 : node3758;
														assign node3758 = (inp[1]) ? 4'b0000 : node3759;
															assign node3759 = (inp[15]) ? 4'b0000 : 4'b1000;
														assign node3763 = (inp[14]) ? node3765 : 4'b0001;
															assign node3765 = (inp[15]) ? 4'b0000 : node3766;
																assign node3766 = (inp[1]) ? 4'b0000 : 4'b0001;
									assign node3770 = (inp[15]) ? node3858 : node3771;
										assign node3771 = (inp[1]) ? node3819 : node3772;
											assign node3772 = (inp[12]) ? node3798 : node3773;
												assign node3773 = (inp[7]) ? node3785 : node3774;
													assign node3774 = (inp[2]) ? node3780 : node3775;
														assign node3775 = (inp[13]) ? node3777 : 4'b0001;
															assign node3777 = (inp[10]) ? 4'b1000 : 4'b1001;
														assign node3780 = (inp[13]) ? 4'b0000 : node3781;
															assign node3781 = (inp[14]) ? 4'b1000 : 4'b0000;
													assign node3785 = (inp[2]) ? node3793 : node3786;
														assign node3786 = (inp[14]) ? node3788 : 4'b0001;
															assign node3788 = (inp[10]) ? 4'b0001 : node3789;
																assign node3789 = (inp[13]) ? 4'b0001 : 4'b0000;
														assign node3793 = (inp[14]) ? 4'b0001 : node3794;
															assign node3794 = (inp[13]) ? 4'b1000 : 4'b0000;
												assign node3798 = (inp[2]) ? node3812 : node3799;
													assign node3799 = (inp[7]) ? node3805 : node3800;
														assign node3800 = (inp[14]) ? node3802 : 4'b1000;
															assign node3802 = (inp[13]) ? 4'b0001 : 4'b1000;
														assign node3805 = (inp[10]) ? node3807 : 4'b1001;
															assign node3807 = (inp[13]) ? node3809 : 4'b1000;
																assign node3809 = (inp[14]) ? 4'b1001 : 4'b1000;
													assign node3812 = (inp[13]) ? 4'b0001 : node3813;
														assign node3813 = (inp[14]) ? 4'b1001 : node3814;
															assign node3814 = (inp[10]) ? 4'b0000 : 4'b1000;
											assign node3819 = (inp[13]) ? node3853 : node3820;
												assign node3820 = (inp[2]) ? node3838 : node3821;
													assign node3821 = (inp[12]) ? node3835 : node3822;
														assign node3822 = (inp[7]) ? node3828 : node3823;
															assign node3823 = (inp[10]) ? node3825 : 4'b1001;
																assign node3825 = (inp[14]) ? 4'b0000 : 4'b0001;
															assign node3828 = (inp[14]) ? node3832 : node3829;
																assign node3829 = (inp[10]) ? 4'b1001 : 4'b1000;
																assign node3832 = (inp[10]) ? 4'b1001 : 4'b0001;
														assign node3835 = (inp[7]) ? 4'b0000 : 4'b0001;
													assign node3838 = (inp[14]) ? node3846 : node3839;
														assign node3839 = (inp[7]) ? node3841 : 4'b0000;
															assign node3841 = (inp[10]) ? 4'b0001 : node3842;
																assign node3842 = (inp[12]) ? 4'b1001 : 4'b0001;
														assign node3846 = (inp[7]) ? node3850 : node3847;
															assign node3847 = (inp[10]) ? 4'b1000 : 4'b0000;
															assign node3850 = (inp[10]) ? 4'b0000 : 4'b1000;
												assign node3853 = (inp[10]) ? node3855 : 4'b0000;
													assign node3855 = (inp[12]) ? 4'b0000 : 4'b1000;
										assign node3858 = (inp[2]) ? node3920 : node3859;
											assign node3859 = (inp[13]) ? node3887 : node3860;
												assign node3860 = (inp[7]) ? node3876 : node3861;
													assign node3861 = (inp[14]) ? node3871 : node3862;
														assign node3862 = (inp[10]) ? 4'b0000 : node3863;
															assign node3863 = (inp[12]) ? node3867 : node3864;
																assign node3864 = (inp[1]) ? 4'b1000 : 4'b0001;
																assign node3867 = (inp[1]) ? 4'b0000 : 4'b1000;
														assign node3871 = (inp[10]) ? node3873 : 4'b0001;
															assign node3873 = (inp[12]) ? 4'b1001 : 4'b1000;
													assign node3876 = (inp[10]) ? node3882 : node3877;
														assign node3877 = (inp[1]) ? 4'b0000 : node3878;
															assign node3878 = (inp[12]) ? 4'b1000 : 4'b0000;
														assign node3882 = (inp[12]) ? node3884 : 4'b1000;
															assign node3884 = (inp[1]) ? 4'b1000 : 4'b0000;
												assign node3887 = (inp[1]) ? node3907 : node3888;
													assign node3888 = (inp[10]) ? node3898 : node3889;
														assign node3889 = (inp[14]) ? node3895 : node3890;
															assign node3890 = (inp[7]) ? node3892 : 4'b0001;
																assign node3892 = (inp[12]) ? 4'b0001 : 4'b1001;
															assign node3895 = (inp[12]) ? 4'b0000 : 4'b1000;
														assign node3898 = (inp[12]) ? node3904 : node3899;
															assign node3899 = (inp[7]) ? 4'b0001 : node3900;
																assign node3900 = (inp[14]) ? 4'b0001 : 4'b0000;
															assign node3904 = (inp[7]) ? 4'b0001 : 4'b1001;
													assign node3907 = (inp[12]) ? node3913 : node3908;
														assign node3908 = (inp[14]) ? 4'b1001 : node3909;
															assign node3909 = (inp[7]) ? 4'b0000 : 4'b1001;
														assign node3913 = (inp[7]) ? node3917 : node3914;
															assign node3914 = (inp[14]) ? 4'b0000 : 4'b0001;
															assign node3917 = (inp[14]) ? 4'b1001 : 4'b1000;
											assign node3920 = (inp[7]) ? 4'b1001 : node3921;
												assign node3921 = (inp[10]) ? node3931 : node3922;
													assign node3922 = (inp[13]) ? node3926 : node3923;
														assign node3923 = (inp[12]) ? 4'b1001 : 4'b0001;
														assign node3926 = (inp[12]) ? node3928 : 4'b1000;
															assign node3928 = (inp[1]) ? 4'b0001 : 4'b0000;
													assign node3931 = (inp[13]) ? node3935 : node3932;
														assign node3932 = (inp[14]) ? 4'b0000 : 4'b0001;
														assign node3935 = (inp[12]) ? 4'b0001 : 4'b1000;
								assign node3939 = (inp[1]) ? node4075 : node3940;
									assign node3940 = (inp[0]) ? node4018 : node3941;
										assign node3941 = (inp[12]) ? node3983 : node3942;
											assign node3942 = (inp[13]) ? node3960 : node3943;
												assign node3943 = (inp[10]) ? node3949 : node3944;
													assign node3944 = (inp[15]) ? node3946 : 4'b1000;
														assign node3946 = (inp[7]) ? 4'b1001 : 4'b1000;
													assign node3949 = (inp[7]) ? node3955 : node3950;
														assign node3950 = (inp[15]) ? node3952 : 4'b1000;
															assign node3952 = (inp[2]) ? 4'b0001 : 4'b1001;
														assign node3955 = (inp[15]) ? 4'b1000 : node3956;
															assign node3956 = (inp[2]) ? 4'b0001 : 4'b0000;
												assign node3960 = (inp[7]) ? node3970 : node3961;
													assign node3961 = (inp[10]) ? node3967 : node3962;
														assign node3962 = (inp[14]) ? 4'b1000 : node3963;
															assign node3963 = (inp[2]) ? 4'b0000 : 4'b0001;
														assign node3967 = (inp[2]) ? 4'b1001 : 4'b0001;
													assign node3970 = (inp[10]) ? node3976 : node3971;
														assign node3971 = (inp[15]) ? node3973 : 4'b0001;
															assign node3973 = (inp[2]) ? 4'b1001 : 4'b1000;
														assign node3976 = (inp[15]) ? node3980 : node3977;
															assign node3977 = (inp[2]) ? 4'b1000 : 4'b0000;
															assign node3980 = (inp[2]) ? 4'b0000 : 4'b1000;
											assign node3983 = (inp[7]) ? node3999 : node3984;
												assign node3984 = (inp[13]) ? node3994 : node3985;
													assign node3985 = (inp[10]) ? node3991 : node3986;
														assign node3986 = (inp[15]) ? 4'b0000 : node3987;
															assign node3987 = (inp[2]) ? 4'b0001 : 4'b1001;
														assign node3991 = (inp[15]) ? 4'b1001 : 4'b0000;
													assign node3994 = (inp[10]) ? 4'b0001 : node3995;
														assign node3995 = (inp[2]) ? 4'b1001 : 4'b0000;
												assign node3999 = (inp[15]) ? node4011 : node4000;
													assign node4000 = (inp[2]) ? node4006 : node4001;
														assign node4001 = (inp[10]) ? 4'b0000 : node4002;
															assign node4002 = (inp[13]) ? 4'b1001 : 4'b1000;
														assign node4006 = (inp[10]) ? node4008 : 4'b0000;
															assign node4008 = (inp[13]) ? 4'b1000 : 4'b1001;
													assign node4011 = (inp[10]) ? node4015 : node4012;
														assign node4012 = (inp[2]) ? 4'b0001 : 4'b0000;
														assign node4015 = (inp[2]) ? 4'b1000 : 4'b0000;
										assign node4018 = (inp[2]) ? node4048 : node4019;
											assign node4019 = (inp[13]) ? node4031 : node4020;
												assign node4020 = (inp[15]) ? node4022 : 4'b0001;
													assign node4022 = (inp[12]) ? node4024 : 4'b0000;
														assign node4024 = (inp[7]) ? node4028 : node4025;
															assign node4025 = (inp[10]) ? 4'b1000 : 4'b0000;
															assign node4028 = (inp[10]) ? 4'b0001 : 4'b1001;
												assign node4031 = (inp[12]) ? node4035 : node4032;
													assign node4032 = (inp[15]) ? 4'b0001 : 4'b0000;
													assign node4035 = (inp[7]) ? node4041 : node4036;
														assign node4036 = (inp[15]) ? 4'b0000 : node4037;
															assign node4037 = (inp[10]) ? 4'b1001 : 4'b1000;
														assign node4041 = (inp[10]) ? node4045 : node4042;
															assign node4042 = (inp[15]) ? 4'b1000 : 4'b0001;
															assign node4045 = (inp[15]) ? 4'b0001 : 4'b0000;
											assign node4048 = (inp[13]) ? node4062 : node4049;
												assign node4049 = (inp[10]) ? node4055 : node4050;
													assign node4050 = (inp[15]) ? 4'b1001 : node4051;
														assign node4051 = (inp[12]) ? 4'b1000 : 4'b0000;
													assign node4055 = (inp[14]) ? 4'b0000 : node4056;
														assign node4056 = (inp[12]) ? node4058 : 4'b1001;
															assign node4058 = (inp[15]) ? 4'b0000 : 4'b0001;
												assign node4062 = (inp[7]) ? node4068 : node4063;
													assign node4063 = (inp[10]) ? 4'b1000 : node4064;
														assign node4064 = (inp[12]) ? 4'b0000 : 4'b0001;
													assign node4068 = (inp[15]) ? 4'b1001 : node4069;
														assign node4069 = (inp[12]) ? 4'b0001 : node4070;
															assign node4070 = (inp[10]) ? 4'b1001 : 4'b0001;
									assign node4075 = (inp[13]) ? node4139 : node4076;
										assign node4076 = (inp[0]) ? node4110 : node4077;
											assign node4077 = (inp[2]) ? node4097 : node4078;
												assign node4078 = (inp[7]) ? node4088 : node4079;
													assign node4079 = (inp[15]) ? node4085 : node4080;
														assign node4080 = (inp[12]) ? 4'b1001 : node4081;
															assign node4081 = (inp[10]) ? 4'b1001 : 4'b0001;
														assign node4085 = (inp[10]) ? 4'b0001 : 4'b1001;
													assign node4088 = (inp[15]) ? node4092 : node4089;
														assign node4089 = (inp[10]) ? 4'b0001 : 4'b1001;
														assign node4092 = (inp[10]) ? 4'b1001 : node4093;
															assign node4093 = (inp[12]) ? 4'b0001 : 4'b1001;
												assign node4097 = (inp[15]) ? node4099 : 4'b0001;
													assign node4099 = (inp[7]) ? node4105 : node4100;
														assign node4100 = (inp[10]) ? 4'b1001 : node4101;
															assign node4101 = (inp[12]) ? 4'b1001 : 4'b0001;
														assign node4105 = (inp[12]) ? node4107 : 4'b0001;
															assign node4107 = (inp[10]) ? 4'b0001 : 4'b1001;
											assign node4110 = (inp[7]) ? node4126 : node4111;
												assign node4111 = (inp[14]) ? node4117 : node4112;
													assign node4112 = (inp[15]) ? node4114 : 4'b1001;
														assign node4114 = (inp[10]) ? 4'b0001 : 4'b1001;
													assign node4117 = (inp[15]) ? 4'b0001 : node4118;
														assign node4118 = (inp[10]) ? node4122 : node4119;
															assign node4119 = (inp[2]) ? 4'b0001 : 4'b1001;
															assign node4122 = (inp[2]) ? 4'b1001 : 4'b0001;
												assign node4126 = (inp[14]) ? node4134 : node4127;
													assign node4127 = (inp[12]) ? 4'b0001 : node4128;
														assign node4128 = (inp[2]) ? 4'b1001 : node4129;
															assign node4129 = (inp[15]) ? 4'b0001 : 4'b1001;
													assign node4134 = (inp[15]) ? 4'b1001 : node4135;
														assign node4135 = (inp[2]) ? 4'b0001 : 4'b1001;
										assign node4139 = (inp[10]) ? 4'b1001 : node4140;
											assign node4140 = (inp[15]) ? node4154 : node4141;
												assign node4141 = (inp[0]) ? node4147 : node4142;
													assign node4142 = (inp[7]) ? node4144 : 4'b1001;
														assign node4144 = (inp[2]) ? 4'b1001 : 4'b0001;
													assign node4147 = (inp[7]) ? node4149 : 4'b0001;
														assign node4149 = (inp[2]) ? 4'b0001 : node4150;
															assign node4150 = (inp[12]) ? 4'b0001 : 4'b1001;
												assign node4154 = (inp[0]) ? node4160 : node4155;
													assign node4155 = (inp[12]) ? node4157 : 4'b0001;
														assign node4157 = (inp[7]) ? 4'b0001 : 4'b1001;
													assign node4160 = (inp[14]) ? node4162 : 4'b1001;
														assign node4162 = (inp[2]) ? node4166 : node4163;
															assign node4163 = (inp[7]) ? 4'b0001 : 4'b1001;
															assign node4166 = (inp[7]) ? 4'b1001 : node4167;
																assign node4167 = (inp[12]) ? 4'b0001 : 4'b1001;
							assign node4172 = (inp[13]) ? node4504 : node4173;
								assign node4173 = (inp[1]) ? node4359 : node4174;
									assign node4174 = (inp[15]) ? node4260 : node4175;
										assign node4175 = (inp[0]) ? node4229 : node4176;
											assign node4176 = (inp[11]) ? node4206 : node4177;
												assign node4177 = (inp[12]) ? node4187 : node4178;
													assign node4178 = (inp[14]) ? 4'b1000 : node4179;
														assign node4179 = (inp[2]) ? 4'b1001 : node4180;
															assign node4180 = (inp[7]) ? node4182 : 4'b0000;
																assign node4182 = (inp[10]) ? 4'b1000 : 4'b1001;
													assign node4187 = (inp[7]) ? node4197 : node4188;
														assign node4188 = (inp[14]) ? node4194 : node4189;
															assign node4189 = (inp[10]) ? 4'b0000 : node4190;
																assign node4190 = (inp[2]) ? 4'b0001 : 4'b1001;
															assign node4194 = (inp[2]) ? 4'b1001 : 4'b1000;
														assign node4197 = (inp[10]) ? node4201 : node4198;
															assign node4198 = (inp[14]) ? 4'b0000 : 4'b0001;
															assign node4201 = (inp[14]) ? 4'b0001 : node4202;
																assign node4202 = (inp[2]) ? 4'b0001 : 4'b0000;
												assign node4206 = (inp[10]) ? node4220 : node4207;
													assign node4207 = (inp[12]) ? node4215 : node4208;
														assign node4208 = (inp[14]) ? node4210 : 4'b0001;
															assign node4210 = (inp[2]) ? 4'b0001 : node4211;
																assign node4211 = (inp[7]) ? 4'b0000 : 4'b0001;
														assign node4215 = (inp[2]) ? node4217 : 4'b1000;
															assign node4217 = (inp[7]) ? 4'b0001 : 4'b0000;
													assign node4220 = (inp[2]) ? node4224 : node4221;
														assign node4221 = (inp[12]) ? 4'b0000 : 4'b1000;
														assign node4224 = (inp[12]) ? node4226 : 4'b0000;
															assign node4226 = (inp[7]) ? 4'b0000 : 4'b0001;
											assign node4229 = (inp[10]) ? node4245 : node4230;
												assign node4230 = (inp[7]) ? node4240 : node4231;
													assign node4231 = (inp[12]) ? node4235 : node4232;
														assign node4232 = (inp[2]) ? 4'b0001 : 4'b0000;
														assign node4235 = (inp[14]) ? node4237 : 4'b1001;
															assign node4237 = (inp[2]) ? 4'b0001 : 4'b1001;
													assign node4240 = (inp[2]) ? 4'b0000 : node4241;
														assign node4241 = (inp[11]) ? 4'b1000 : 4'b0001;
												assign node4245 = (inp[7]) ? node4255 : node4246;
													assign node4246 = (inp[2]) ? node4252 : node4247;
														assign node4247 = (inp[11]) ? 4'b0001 : node4248;
															assign node4248 = (inp[12]) ? 4'b0001 : 4'b0000;
														assign node4252 = (inp[14]) ? 4'b0001 : 4'b1000;
													assign node4255 = (inp[2]) ? 4'b0001 : node4256;
														assign node4256 = (inp[12]) ? 4'b0001 : 4'b0000;
										assign node4260 = (inp[14]) ? node4306 : node4261;
											assign node4261 = (inp[2]) ? node4279 : node4262;
												assign node4262 = (inp[0]) ? node4270 : node4263;
													assign node4263 = (inp[7]) ? 4'b0001 : node4264;
														assign node4264 = (inp[10]) ? node4266 : 4'b1000;
															assign node4266 = (inp[11]) ? 4'b1000 : 4'b1001;
													assign node4270 = (inp[11]) ? node4272 : 4'b0001;
														assign node4272 = (inp[12]) ? 4'b0000 : node4273;
															assign node4273 = (inp[7]) ? 4'b1000 : node4274;
																assign node4274 = (inp[10]) ? 4'b0000 : 4'b1001;
												assign node4279 = (inp[11]) ? node4299 : node4280;
													assign node4280 = (inp[7]) ? node4292 : node4281;
														assign node4281 = (inp[0]) ? node4287 : node4282;
															assign node4282 = (inp[12]) ? 4'b0000 : node4283;
																assign node4283 = (inp[10]) ? 4'b0000 : 4'b1000;
															assign node4287 = (inp[10]) ? 4'b1000 : node4288;
																assign node4288 = (inp[12]) ? 4'b1000 : 4'b0000;
														assign node4292 = (inp[12]) ? node4294 : 4'b0000;
															assign node4294 = (inp[10]) ? node4296 : 4'b1001;
																assign node4296 = (inp[0]) ? 4'b0000 : 4'b0001;
													assign node4299 = (inp[7]) ? node4301 : 4'b0001;
														assign node4301 = (inp[12]) ? 4'b1000 : node4302;
															assign node4302 = (inp[0]) ? 4'b0000 : 4'b0001;
											assign node4306 = (inp[2]) ? node4328 : node4307;
												assign node4307 = (inp[0]) ? node4319 : node4308;
													assign node4308 = (inp[12]) ? node4316 : node4309;
														assign node4309 = (inp[10]) ? node4311 : 4'b1000;
															assign node4311 = (inp[11]) ? 4'b0001 : node4312;
																assign node4312 = (inp[7]) ? 4'b1000 : 4'b0001;
														assign node4316 = (inp[7]) ? 4'b0001 : 4'b1000;
													assign node4319 = (inp[7]) ? node4323 : node4320;
														assign node4320 = (inp[11]) ? 4'b0001 : 4'b0000;
														assign node4323 = (inp[12]) ? node4325 : 4'b1000;
															assign node4325 = (inp[11]) ? 4'b0000 : 4'b1000;
												assign node4328 = (inp[11]) ? node4344 : node4329;
													assign node4329 = (inp[7]) ? node4335 : node4330;
														assign node4330 = (inp[0]) ? node4332 : 4'b0000;
															assign node4332 = (inp[12]) ? 4'b1001 : 4'b1000;
														assign node4335 = (inp[10]) ? node4339 : node4336;
															assign node4336 = (inp[0]) ? 4'b1001 : 4'b0001;
															assign node4339 = (inp[12]) ? 4'b0001 : node4340;
																assign node4340 = (inp[0]) ? 4'b0001 : 4'b1001;
													assign node4344 = (inp[10]) ? node4352 : node4345;
														assign node4345 = (inp[12]) ? node4347 : 4'b0001;
															assign node4347 = (inp[7]) ? node4349 : 4'b0000;
																assign node4349 = (inp[0]) ? 4'b1001 : 4'b1000;
														assign node4352 = (inp[0]) ? node4354 : 4'b1000;
															assign node4354 = (inp[12]) ? node4356 : 4'b0000;
																assign node4356 = (inp[7]) ? 4'b0000 : 4'b0001;
									assign node4359 = (inp[11]) ? node4461 : node4360;
										assign node4360 = (inp[10]) ? node4406 : node4361;
											assign node4361 = (inp[15]) ? node4387 : node4362;
												assign node4362 = (inp[12]) ? node4376 : node4363;
													assign node4363 = (inp[7]) ? node4371 : node4364;
														assign node4364 = (inp[2]) ? 4'b1001 : node4365;
															assign node4365 = (inp[0]) ? node4367 : 4'b1000;
																assign node4367 = (inp[14]) ? 4'b1000 : 4'b1001;
														assign node4371 = (inp[2]) ? 4'b1000 : node4372;
															assign node4372 = (inp[0]) ? 4'b0001 : 4'b0000;
													assign node4376 = (inp[2]) ? 4'b0001 : node4377;
														assign node4377 = (inp[7]) ? node4383 : node4378;
															assign node4378 = (inp[14]) ? node4380 : 4'b0001;
																assign node4380 = (inp[0]) ? 4'b0000 : 4'b0001;
															assign node4383 = (inp[0]) ? 4'b0001 : 4'b0000;
												assign node4387 = (inp[12]) ? node4399 : node4388;
													assign node4388 = (inp[14]) ? node4394 : node4389;
														assign node4389 = (inp[0]) ? node4391 : 4'b0001;
															assign node4391 = (inp[2]) ? 4'b0001 : 4'b0000;
														assign node4394 = (inp[0]) ? 4'b0000 : node4395;
															assign node4395 = (inp[7]) ? 4'b1000 : 4'b0000;
													assign node4399 = (inp[0]) ? node4403 : node4400;
														assign node4400 = (inp[7]) ? 4'b1000 : 4'b1001;
														assign node4403 = (inp[14]) ? 4'b1000 : 4'b0000;
											assign node4406 = (inp[14]) ? node4434 : node4407;
												assign node4407 = (inp[15]) ? node4413 : node4408;
													assign node4408 = (inp[2]) ? 4'b0000 : node4409;
														assign node4409 = (inp[12]) ? 4'b1000 : 4'b0000;
													assign node4413 = (inp[12]) ? node4429 : node4414;
														assign node4414 = (inp[2]) ? node4422 : node4415;
															assign node4415 = (inp[7]) ? node4419 : node4416;
																assign node4416 = (inp[0]) ? 4'b0000 : 4'b0001;
																assign node4419 = (inp[0]) ? 4'b0001 : 4'b0000;
															assign node4422 = (inp[7]) ? node4426 : node4423;
																assign node4423 = (inp[0]) ? 4'b0000 : 4'b0001;
																assign node4426 = (inp[0]) ? 4'b0001 : 4'b1000;
														assign node4429 = (inp[7]) ? node4431 : 4'b0000;
															assign node4431 = (inp[0]) ? 4'b0001 : 4'b0000;
												assign node4434 = (inp[15]) ? node4446 : node4435;
													assign node4435 = (inp[7]) ? node4441 : node4436;
														assign node4436 = (inp[0]) ? node4438 : 4'b0001;
															assign node4438 = (inp[12]) ? 4'b0000 : 4'b1000;
														assign node4441 = (inp[0]) ? 4'b0001 : node4442;
															assign node4442 = (inp[2]) ? 4'b0001 : 4'b0000;
													assign node4446 = (inp[7]) ? node4454 : node4447;
														assign node4447 = (inp[0]) ? node4451 : node4448;
															assign node4448 = (inp[2]) ? 4'b0000 : 4'b0001;
															assign node4451 = (inp[2]) ? 4'b0001 : 4'b0000;
														assign node4454 = (inp[0]) ? node4458 : node4455;
															assign node4455 = (inp[12]) ? 4'b0000 : 4'b1000;
															assign node4458 = (inp[2]) ? 4'b0000 : 4'b0001;
										assign node4461 = (inp[10]) ? 4'b0001 : node4462;
											assign node4462 = (inp[7]) ? node4482 : node4463;
												assign node4463 = (inp[15]) ? node4471 : node4464;
													assign node4464 = (inp[0]) ? 4'b0001 : node4465;
														assign node4465 = (inp[12]) ? node4467 : 4'b1001;
															assign node4467 = (inp[14]) ? 4'b0001 : 4'b1001;
													assign node4471 = (inp[0]) ? node4477 : node4472;
														assign node4472 = (inp[2]) ? node4474 : 4'b0001;
															assign node4474 = (inp[12]) ? 4'b1001 : 4'b0001;
														assign node4477 = (inp[2]) ? 4'b0001 : node4478;
															assign node4478 = (inp[12]) ? 4'b0001 : 4'b1001;
												assign node4482 = (inp[2]) ? node4496 : node4483;
													assign node4483 = (inp[0]) ? node4491 : node4484;
														assign node4484 = (inp[15]) ? node4488 : node4485;
															assign node4485 = (inp[12]) ? 4'b0001 : 4'b1001;
															assign node4488 = (inp[12]) ? 4'b1001 : 4'b0001;
														assign node4491 = (inp[12]) ? node4493 : 4'b0001;
															assign node4493 = (inp[15]) ? 4'b0001 : 4'b1001;
													assign node4496 = (inp[0]) ? 4'b1001 : node4497;
														assign node4497 = (inp[15]) ? node4499 : 4'b0001;
															assign node4499 = (inp[14]) ? 4'b1001 : 4'b0001;
								assign node4504 = (inp[10]) ? node4622 : node4505;
									assign node4505 = (inp[1]) ? node4589 : node4506;
										assign node4506 = (inp[11]) ? node4550 : node4507;
											assign node4507 = (inp[15]) ? node4525 : node4508;
												assign node4508 = (inp[12]) ? node4514 : node4509;
													assign node4509 = (inp[2]) ? 4'b0001 : node4510;
														assign node4510 = (inp[0]) ? 4'b0001 : 4'b0000;
													assign node4514 = (inp[2]) ? node4520 : node4515;
														assign node4515 = (inp[7]) ? 4'b0001 : node4516;
															assign node4516 = (inp[0]) ? 4'b0000 : 4'b0001;
														assign node4520 = (inp[14]) ? 4'b0000 : node4521;
															assign node4521 = (inp[0]) ? 4'b0001 : 4'b0000;
												assign node4525 = (inp[12]) ? node4537 : node4526;
													assign node4526 = (inp[7]) ? node4532 : node4527;
														assign node4527 = (inp[14]) ? 4'b0001 : node4528;
															assign node4528 = (inp[0]) ? 4'b0000 : 4'b0001;
														assign node4532 = (inp[14]) ? 4'b0000 : node4533;
															assign node4533 = (inp[0]) ? 4'b0001 : 4'b0000;
													assign node4537 = (inp[2]) ? node4543 : node4538;
														assign node4538 = (inp[7]) ? 4'b0000 : node4539;
															assign node4539 = (inp[0]) ? 4'b0001 : 4'b0000;
														assign node4543 = (inp[7]) ? node4545 : 4'b0000;
															assign node4545 = (inp[14]) ? 4'b0001 : node4546;
																assign node4546 = (inp[0]) ? 4'b0000 : 4'b0001;
											assign node4550 = (inp[12]) ? node4568 : node4551;
												assign node4551 = (inp[15]) ? node4563 : node4552;
													assign node4552 = (inp[2]) ? 4'b0000 : node4553;
														assign node4553 = (inp[14]) ? node4555 : 4'b0000;
															assign node4555 = (inp[7]) ? node4559 : node4556;
																assign node4556 = (inp[0]) ? 4'b0000 : 4'b0001;
																assign node4559 = (inp[0]) ? 4'b0001 : 4'b0000;
													assign node4563 = (inp[2]) ? node4565 : 4'b0000;
														assign node4565 = (inp[14]) ? 4'b0000 : 4'b0001;
												assign node4568 = (inp[2]) ? node4580 : node4569;
													assign node4569 = (inp[15]) ? node4575 : node4570;
														assign node4570 = (inp[0]) ? node4572 : 4'b0000;
															assign node4572 = (inp[7]) ? 4'b0000 : 4'b0001;
														assign node4575 = (inp[7]) ? node4577 : 4'b0001;
															assign node4577 = (inp[0]) ? 4'b0001 : 4'b0000;
													assign node4580 = (inp[15]) ? node4584 : node4581;
														assign node4581 = (inp[0]) ? 4'b0000 : 4'b0001;
														assign node4584 = (inp[0]) ? node4586 : 4'b0000;
															assign node4586 = (inp[7]) ? 4'b0000 : 4'b0001;
										assign node4589 = (inp[11]) ? 4'b0001 : node4590;
											assign node4590 = (inp[14]) ? node4604 : node4591;
												assign node4591 = (inp[0]) ? node4599 : node4592;
													assign node4592 = (inp[15]) ? node4594 : 4'b0000;
														assign node4594 = (inp[12]) ? node4596 : 4'b0001;
															assign node4596 = (inp[7]) ? 4'b0001 : 4'b0000;
													assign node4599 = (inp[15]) ? 4'b0000 : node4600;
														assign node4600 = (inp[12]) ? 4'b0001 : 4'b0000;
												assign node4604 = (inp[7]) ? node4614 : node4605;
													assign node4605 = (inp[2]) ? 4'b0001 : node4606;
														assign node4606 = (inp[0]) ? node4610 : node4607;
															assign node4607 = (inp[15]) ? 4'b0001 : 4'b0000;
															assign node4610 = (inp[15]) ? 4'b0000 : 4'b0001;
													assign node4614 = (inp[0]) ? node4616 : 4'b0001;
														assign node4616 = (inp[2]) ? node4618 : 4'b0001;
															assign node4618 = (inp[15]) ? 4'b0000 : 4'b0001;
									assign node4622 = (inp[11]) ? 4'b0000 : node4623;
										assign node4623 = (inp[1]) ? 4'b0000 : node4624;
											assign node4624 = (inp[2]) ? node4642 : node4625;
												assign node4625 = (inp[12]) ? node4635 : node4626;
													assign node4626 = (inp[14]) ? node4628 : 4'b0000;
														assign node4628 = (inp[15]) ? node4632 : node4629;
															assign node4629 = (inp[0]) ? 4'b0001 : 4'b0000;
															assign node4632 = (inp[0]) ? 4'b0000 : 4'b0001;
													assign node4635 = (inp[14]) ? 4'b0000 : node4636;
														assign node4636 = (inp[0]) ? 4'b0000 : node4637;
															assign node4637 = (inp[15]) ? 4'b0000 : 4'b0001;
												assign node4642 = (inp[15]) ? node4654 : node4643;
													assign node4643 = (inp[14]) ? 4'b0000 : node4644;
														assign node4644 = (inp[7]) ? 4'b0000 : node4645;
															assign node4645 = (inp[0]) ? node4649 : node4646;
																assign node4646 = (inp[12]) ? 4'b0000 : 4'b0001;
																assign node4649 = (inp[12]) ? 4'b0001 : 4'b0000;
													assign node4654 = (inp[12]) ? node4658 : node4655;
														assign node4655 = (inp[14]) ? 4'b0001 : 4'b0000;
														assign node4658 = (inp[14]) ? 4'b0000 : node4659;
															assign node4659 = (inp[7]) ? 4'b0001 : node4660;
																assign node4660 = (inp[0]) ? 4'b0000 : 4'b0001;
			assign node4667 = (inp[15]) ? node7255 : node4668;
				assign node4668 = (inp[6]) ? node5370 : node4669;
					assign node4669 = (inp[0]) ? 4'b0101 : node4670;
						assign node4670 = (inp[5]) ? node4878 : node4671;
							assign node4671 = (inp[2]) ? 4'b0111 : node4672;
								assign node4672 = (inp[3]) ? node4754 : node4673;
									assign node4673 = (inp[7]) ? node4729 : node4674;
										assign node4674 = (inp[4]) ? node4694 : node4675;
											assign node4675 = (inp[13]) ? node4677 : 4'b0111;
												assign node4677 = (inp[12]) ? node4683 : node4678;
													assign node4678 = (inp[14]) ? 4'b0000 : node4679;
														assign node4679 = (inp[1]) ? 4'b0001 : 4'b0000;
													assign node4683 = (inp[10]) ? node4685 : 4'b0111;
														assign node4685 = (inp[14]) ? node4687 : 4'b0000;
															assign node4687 = (inp[1]) ? node4691 : node4688;
																assign node4688 = (inp[11]) ? 4'b0000 : 4'b0111;
																assign node4691 = (inp[11]) ? 4'b0001 : 4'b0000;
											assign node4694 = (inp[1]) ? node4716 : node4695;
												assign node4695 = (inp[11]) ? node4707 : node4696;
													assign node4696 = (inp[14]) ? node4698 : 4'b1000;
														assign node4698 = (inp[12]) ? node4704 : node4699;
															assign node4699 = (inp[13]) ? 4'b0001 : node4700;
																assign node4700 = (inp[10]) ? 4'b1001 : 4'b0001;
															assign node4704 = (inp[13]) ? 4'b1001 : 4'b0001;
													assign node4707 = (inp[10]) ? 4'b1000 : node4708;
														assign node4708 = (inp[14]) ? 4'b0000 : node4709;
															assign node4709 = (inp[13]) ? 4'b1000 : node4710;
																assign node4710 = (inp[12]) ? 4'b0000 : 4'b1000;
												assign node4716 = (inp[13]) ? node4722 : node4717;
													assign node4717 = (inp[12]) ? node4719 : 4'b1001;
														assign node4719 = (inp[10]) ? 4'b1001 : 4'b0001;
													assign node4722 = (inp[10]) ? 4'b0001 : node4723;
														assign node4723 = (inp[12]) ? 4'b1001 : node4724;
															assign node4724 = (inp[11]) ? 4'b0001 : 4'b0000;
										assign node4729 = (inp[13]) ? node4731 : 4'b0111;
											assign node4731 = (inp[4]) ? node4733 : 4'b0111;
												assign node4733 = (inp[12]) ? node4749 : node4734;
													assign node4734 = (inp[14]) ? node4736 : 4'b0000;
														assign node4736 = (inp[10]) ? node4742 : node4737;
															assign node4737 = (inp[1]) ? 4'b0000 : node4738;
																assign node4738 = (inp[11]) ? 4'b0000 : 4'b0111;
															assign node4742 = (inp[1]) ? node4746 : node4743;
																assign node4743 = (inp[11]) ? 4'b0000 : 4'b0001;
																assign node4746 = (inp[11]) ? 4'b0001 : 4'b0000;
													assign node4749 = (inp[10]) ? node4751 : 4'b0111;
														assign node4751 = (inp[1]) ? 4'b0001 : 4'b0000;
									assign node4754 = (inp[13]) ? node4812 : node4755;
										assign node4755 = (inp[1]) ? node4783 : node4756;
											assign node4756 = (inp[14]) ? node4766 : node4757;
												assign node4757 = (inp[4]) ? node4763 : node4758;
													assign node4758 = (inp[10]) ? 4'b1000 : node4759;
														assign node4759 = (inp[12]) ? 4'b0000 : 4'b1000;
													assign node4763 = (inp[7]) ? 4'b1000 : 4'b1100;
												assign node4766 = (inp[11]) ? node4770 : node4767;
													assign node4767 = (inp[7]) ? 4'b0001 : 4'b0101;
													assign node4770 = (inp[12]) ? node4776 : node4771;
														assign node4771 = (inp[4]) ? node4773 : 4'b1000;
															assign node4773 = (inp[7]) ? 4'b1000 : 4'b1100;
														assign node4776 = (inp[10]) ? node4780 : node4777;
															assign node4777 = (inp[7]) ? 4'b0000 : 4'b0100;
															assign node4780 = (inp[4]) ? 4'b1100 : 4'b1000;
											assign node4783 = (inp[4]) ? node4797 : node4784;
												assign node4784 = (inp[12]) ? node4790 : node4785;
													assign node4785 = (inp[11]) ? 4'b1001 : node4786;
														assign node4786 = (inp[14]) ? 4'b1000 : 4'b1001;
													assign node4790 = (inp[10]) ? 4'b1001 : node4791;
														assign node4791 = (inp[7]) ? node4793 : 4'b0001;
															assign node4793 = (inp[14]) ? 4'b0000 : 4'b0001;
												assign node4797 = (inp[7]) ? node4807 : node4798;
													assign node4798 = (inp[14]) ? node4804 : node4799;
														assign node4799 = (inp[12]) ? node4801 : 4'b1101;
															assign node4801 = (inp[10]) ? 4'b1101 : 4'b0101;
														assign node4804 = (inp[11]) ? 4'b1101 : 4'b1100;
													assign node4807 = (inp[12]) ? node4809 : 4'b1001;
														assign node4809 = (inp[10]) ? 4'b1001 : 4'b0001;
										assign node4812 = (inp[10]) ? node4844 : node4813;
											assign node4813 = (inp[12]) ? node4831 : node4814;
												assign node4814 = (inp[4]) ? node4826 : node4815;
													assign node4815 = (inp[7]) ? node4821 : node4816;
														assign node4816 = (inp[11]) ? 4'b0100 : node4817;
															assign node4817 = (inp[14]) ? 4'b1001 : 4'b0100;
														assign node4821 = (inp[1]) ? node4823 : 4'b0000;
															assign node4823 = (inp[11]) ? 4'b0001 : 4'b0000;
													assign node4826 = (inp[11]) ? node4828 : 4'b0100;
														assign node4828 = (inp[1]) ? 4'b0101 : 4'b0100;
												assign node4831 = (inp[1]) ? node4839 : node4832;
													assign node4832 = (inp[4]) ? node4836 : node4833;
														assign node4833 = (inp[14]) ? 4'b1001 : 4'b1000;
														assign node4836 = (inp[7]) ? 4'b1000 : 4'b1100;
													assign node4839 = (inp[11]) ? 4'b1001 : node4840;
														assign node4840 = (inp[4]) ? 4'b1001 : 4'b1000;
											assign node4844 = (inp[7]) ? node4856 : node4845;
												assign node4845 = (inp[1]) ? node4851 : node4846;
													assign node4846 = (inp[11]) ? 4'b0100 : node4847;
														assign node4847 = (inp[4]) ? 4'b0100 : 4'b0101;
													assign node4851 = (inp[11]) ? 4'b0101 : node4852;
														assign node4852 = (inp[14]) ? 4'b0100 : 4'b0101;
												assign node4856 = (inp[4]) ? node4866 : node4857;
													assign node4857 = (inp[12]) ? node4859 : 4'b0001;
														assign node4859 = (inp[11]) ? 4'b0000 : node4860;
															assign node4860 = (inp[1]) ? node4862 : 4'b1001;
																assign node4862 = (inp[14]) ? 4'b0000 : 4'b0001;
													assign node4866 = (inp[11]) ? 4'b0100 : node4867;
														assign node4867 = (inp[12]) ? 4'b0100 : node4868;
															assign node4868 = (inp[1]) ? node4872 : node4869;
																assign node4869 = (inp[14]) ? 4'b0101 : 4'b0100;
																assign node4872 = (inp[14]) ? 4'b0100 : 4'b0101;
							assign node4878 = (inp[1]) ? node5110 : node4879;
								assign node4879 = (inp[2]) ? node5005 : node4880;
									assign node4880 = (inp[14]) ? node4924 : node4881;
										assign node4881 = (inp[13]) ? node4907 : node4882;
											assign node4882 = (inp[10]) ? node4896 : node4883;
												assign node4883 = (inp[12]) ? node4889 : node4884;
													assign node4884 = (inp[3]) ? node4886 : 4'b1100;
														assign node4886 = (inp[4]) ? 4'b1100 : 4'b1000;
													assign node4889 = (inp[4]) ? node4891 : 4'b0100;
														assign node4891 = (inp[7]) ? 4'b0000 : node4892;
															assign node4892 = (inp[3]) ? 4'b0100 : 4'b0000;
												assign node4896 = (inp[3]) ? node4902 : node4897;
													assign node4897 = (inp[7]) ? 4'b1100 : node4898;
														assign node4898 = (inp[4]) ? 4'b1000 : 4'b1100;
													assign node4902 = (inp[7]) ? 4'b1000 : node4903;
														assign node4903 = (inp[4]) ? 4'b1100 : 4'b1000;
											assign node4907 = (inp[10]) ? node4915 : node4908;
												assign node4908 = (inp[12]) ? node4912 : node4909;
													assign node4909 = (inp[3]) ? 4'b0100 : 4'b0000;
													assign node4912 = (inp[3]) ? 4'b1000 : 4'b1100;
												assign node4915 = (inp[3]) ? node4921 : node4916;
													assign node4916 = (inp[7]) ? node4918 : 4'b0000;
														assign node4918 = (inp[4]) ? 4'b0000 : 4'b0100;
													assign node4921 = (inp[7]) ? 4'b0000 : 4'b0100;
										assign node4924 = (inp[11]) ? node4960 : node4925;
											assign node4925 = (inp[13]) ? node4941 : node4926;
												assign node4926 = (inp[10]) ? node4936 : node4927;
													assign node4927 = (inp[4]) ? node4931 : node4928;
														assign node4928 = (inp[3]) ? 4'b0001 : 4'b0101;
														assign node4931 = (inp[3]) ? 4'b0101 : node4932;
															assign node4932 = (inp[7]) ? 4'b0101 : 4'b0001;
													assign node4936 = (inp[12]) ? 4'b0001 : node4937;
														assign node4937 = (inp[4]) ? 4'b1001 : 4'b1101;
												assign node4941 = (inp[10]) ? node4949 : node4942;
													assign node4942 = (inp[7]) ? 4'b1001 : node4943;
														assign node4943 = (inp[12]) ? 4'b1101 : node4944;
															assign node4944 = (inp[4]) ? 4'b1101 : 4'b1001;
													assign node4949 = (inp[12]) ? node4955 : node4950;
														assign node4950 = (inp[3]) ? 4'b0101 : node4951;
															assign node4951 = (inp[7]) ? 4'b0101 : 4'b0001;
														assign node4955 = (inp[4]) ? 4'b1001 : node4956;
															assign node4956 = (inp[3]) ? 4'b1001 : 4'b1101;
											assign node4960 = (inp[10]) ? node4986 : node4961;
												assign node4961 = (inp[3]) ? node4975 : node4962;
													assign node4962 = (inp[7]) ? node4972 : node4963;
														assign node4963 = (inp[4]) ? node4967 : node4964;
															assign node4964 = (inp[12]) ? 4'b0100 : 4'b1100;
															assign node4967 = (inp[12]) ? node4969 : 4'b0000;
																assign node4969 = (inp[13]) ? 4'b1000 : 4'b0000;
														assign node4972 = (inp[13]) ? 4'b1100 : 4'b0100;
													assign node4975 = (inp[7]) ? node4979 : node4976;
														assign node4976 = (inp[4]) ? 4'b1100 : 4'b1000;
														assign node4979 = (inp[4]) ? 4'b1000 : node4980;
															assign node4980 = (inp[12]) ? node4982 : 4'b1000;
																assign node4982 = (inp[13]) ? 4'b1000 : 4'b0000;
												assign node4986 = (inp[13]) ? node5000 : node4987;
													assign node4987 = (inp[12]) ? 4'b1100 : node4988;
														assign node4988 = (inp[3]) ? node4994 : node4989;
															assign node4989 = (inp[4]) ? node4991 : 4'b1100;
																assign node4991 = (inp[7]) ? 4'b1100 : 4'b1000;
															assign node4994 = (inp[4]) ? node4996 : 4'b1000;
																assign node4996 = (inp[7]) ? 4'b1000 : 4'b1100;
													assign node5000 = (inp[3]) ? 4'b0100 : node5001;
														assign node5001 = (inp[4]) ? 4'b0000 : 4'b0100;
									assign node5005 = (inp[3]) ? node5045 : node5006;
										assign node5006 = (inp[7]) ? node5034 : node5007;
											assign node5007 = (inp[4]) ? node5017 : node5008;
												assign node5008 = (inp[13]) ? node5010 : 4'b0111;
													assign node5010 = (inp[10]) ? 4'b0000 : node5011;
														assign node5011 = (inp[12]) ? 4'b0111 : node5012;
															assign node5012 = (inp[14]) ? 4'b0111 : 4'b0000;
												assign node5017 = (inp[10]) ? node5027 : node5018;
													assign node5018 = (inp[11]) ? node5022 : node5019;
														assign node5019 = (inp[14]) ? 4'b0001 : 4'b0000;
														assign node5022 = (inp[13]) ? 4'b0000 : node5023;
															assign node5023 = (inp[12]) ? 4'b0000 : 4'b1000;
													assign node5027 = (inp[11]) ? node5031 : node5028;
														assign node5028 = (inp[14]) ? 4'b1001 : 4'b1000;
														assign node5031 = (inp[13]) ? 4'b0000 : 4'b1000;
											assign node5034 = (inp[13]) ? node5036 : 4'b0111;
												assign node5036 = (inp[4]) ? node5038 : 4'b0111;
													assign node5038 = (inp[12]) ? node5040 : 4'b0000;
														assign node5040 = (inp[10]) ? node5042 : 4'b0111;
															assign node5042 = (inp[14]) ? 4'b0111 : 4'b0000;
										assign node5045 = (inp[14]) ? node5073 : node5046;
											assign node5046 = (inp[13]) ? node5060 : node5047;
												assign node5047 = (inp[7]) ? node5055 : node5048;
													assign node5048 = (inp[4]) ? node5052 : node5049;
														assign node5049 = (inp[10]) ? 4'b1000 : 4'b0000;
														assign node5052 = (inp[12]) ? 4'b0100 : 4'b1100;
													assign node5055 = (inp[4]) ? 4'b1000 : node5056;
														assign node5056 = (inp[12]) ? 4'b0000 : 4'b1000;
												assign node5060 = (inp[7]) ? node5066 : node5061;
													assign node5061 = (inp[12]) ? node5063 : 4'b0100;
														assign node5063 = (inp[10]) ? 4'b0100 : 4'b1000;
													assign node5066 = (inp[4]) ? 4'b0100 : node5067;
														assign node5067 = (inp[12]) ? node5069 : 4'b0000;
															assign node5069 = (inp[10]) ? 4'b0000 : 4'b1000;
											assign node5073 = (inp[11]) ? node5095 : node5074;
												assign node5074 = (inp[4]) ? node5084 : node5075;
													assign node5075 = (inp[12]) ? 4'b0001 : node5076;
														assign node5076 = (inp[13]) ? node5080 : node5077;
															assign node5077 = (inp[10]) ? 4'b1001 : 4'b0001;
															assign node5080 = (inp[10]) ? 4'b0001 : 4'b1001;
													assign node5084 = (inp[7]) ? node5090 : node5085;
														assign node5085 = (inp[13]) ? node5087 : 4'b0101;
															assign node5087 = (inp[10]) ? 4'b0101 : 4'b1101;
														assign node5090 = (inp[13]) ? 4'b0101 : node5091;
															assign node5091 = (inp[10]) ? 4'b1001 : 4'b0001;
												assign node5095 = (inp[13]) ? node5107 : node5096;
													assign node5096 = (inp[12]) ? node5102 : node5097;
														assign node5097 = (inp[7]) ? 4'b1000 : node5098;
															assign node5098 = (inp[4]) ? 4'b1100 : 4'b1000;
														assign node5102 = (inp[10]) ? 4'b1000 : node5103;
															assign node5103 = (inp[4]) ? 4'b0100 : 4'b0000;
													assign node5107 = (inp[4]) ? 4'b0100 : 4'b0000;
								assign node5110 = (inp[14]) ? node5196 : node5111;
									assign node5111 = (inp[13]) ? node5151 : node5112;
										assign node5112 = (inp[3]) ? node5134 : node5113;
											assign node5113 = (inp[2]) ? node5127 : node5114;
												assign node5114 = (inp[4]) ? node5120 : node5115;
													assign node5115 = (inp[12]) ? node5117 : 4'b1101;
														assign node5117 = (inp[10]) ? 4'b1101 : 4'b0101;
													assign node5120 = (inp[7]) ? 4'b1101 : node5121;
														assign node5121 = (inp[12]) ? node5123 : 4'b1001;
															assign node5123 = (inp[10]) ? 4'b1001 : 4'b0001;
												assign node5127 = (inp[4]) ? node5129 : 4'b0111;
													assign node5129 = (inp[7]) ? 4'b0111 : node5130;
														assign node5130 = (inp[12]) ? 4'b0001 : 4'b1001;
											assign node5134 = (inp[10]) ? node5146 : node5135;
												assign node5135 = (inp[12]) ? node5141 : node5136;
													assign node5136 = (inp[4]) ? node5138 : 4'b1001;
														assign node5138 = (inp[7]) ? 4'b1001 : 4'b1101;
													assign node5141 = (inp[4]) ? node5143 : 4'b0001;
														assign node5143 = (inp[7]) ? 4'b0001 : 4'b0101;
												assign node5146 = (inp[4]) ? node5148 : 4'b1001;
													assign node5148 = (inp[7]) ? 4'b1001 : 4'b1101;
										assign node5151 = (inp[12]) ? node5165 : node5152;
											assign node5152 = (inp[3]) ? node5160 : node5153;
												assign node5153 = (inp[4]) ? 4'b0001 : node5154;
													assign node5154 = (inp[7]) ? node5156 : 4'b0001;
														assign node5156 = (inp[2]) ? 4'b0111 : 4'b0101;
												assign node5160 = (inp[7]) ? node5162 : 4'b0101;
													assign node5162 = (inp[4]) ? 4'b0101 : 4'b0001;
											assign node5165 = (inp[10]) ? node5185 : node5166;
												assign node5166 = (inp[11]) ? node5176 : node5167;
													assign node5167 = (inp[4]) ? node5169 : 4'b1101;
														assign node5169 = (inp[3]) ? node5173 : node5170;
															assign node5170 = (inp[7]) ? 4'b1101 : 4'b1001;
															assign node5173 = (inp[7]) ? 4'b1001 : 4'b1101;
													assign node5176 = (inp[3]) ? node5182 : node5177;
														assign node5177 = (inp[7]) ? node5179 : 4'b1001;
															assign node5179 = (inp[4]) ? 4'b0111 : 4'b1101;
														assign node5182 = (inp[7]) ? 4'b1001 : 4'b1101;
												assign node5185 = (inp[3]) ? node5191 : node5186;
													assign node5186 = (inp[7]) ? node5188 : 4'b0001;
														assign node5188 = (inp[4]) ? 4'b0001 : 4'b0111;
													assign node5191 = (inp[4]) ? 4'b0101 : node5192;
														assign node5192 = (inp[7]) ? 4'b0001 : 4'b0101;
									assign node5196 = (inp[11]) ? node5282 : node5197;
										assign node5197 = (inp[2]) ? node5235 : node5198;
											assign node5198 = (inp[13]) ? node5216 : node5199;
												assign node5199 = (inp[12]) ? node5205 : node5200;
													assign node5200 = (inp[3]) ? node5202 : 4'b1100;
														assign node5202 = (inp[4]) ? 4'b1100 : 4'b1000;
													assign node5205 = (inp[10]) ? node5213 : node5206;
														assign node5206 = (inp[3]) ? 4'b0000 : node5207;
															assign node5207 = (inp[4]) ? node5209 : 4'b0100;
																assign node5209 = (inp[7]) ? 4'b0100 : 4'b0000;
														assign node5213 = (inp[7]) ? 4'b1100 : 4'b1000;
												assign node5216 = (inp[12]) ? node5222 : node5217;
													assign node5217 = (inp[3]) ? 4'b0100 : node5218;
														assign node5218 = (inp[4]) ? 4'b0000 : 4'b0100;
													assign node5222 = (inp[10]) ? node5226 : node5223;
														assign node5223 = (inp[3]) ? 4'b1000 : 4'b1100;
														assign node5226 = (inp[7]) ? node5228 : 4'b0100;
															assign node5228 = (inp[3]) ? node5232 : node5229;
																assign node5229 = (inp[4]) ? 4'b0000 : 4'b0100;
																assign node5232 = (inp[4]) ? 4'b0100 : 4'b0000;
											assign node5235 = (inp[3]) ? node5261 : node5236;
												assign node5236 = (inp[4]) ? node5244 : node5237;
													assign node5237 = (inp[7]) ? 4'b0111 : node5238;
														assign node5238 = (inp[12]) ? 4'b0111 : node5239;
															assign node5239 = (inp[13]) ? 4'b0000 : 4'b0111;
													assign node5244 = (inp[7]) ? node5254 : node5245;
														assign node5245 = (inp[12]) ? node5247 : 4'b1000;
															assign node5247 = (inp[10]) ? node5251 : node5248;
																assign node5248 = (inp[13]) ? 4'b1000 : 4'b0000;
																assign node5251 = (inp[13]) ? 4'b0000 : 4'b1000;
														assign node5254 = (inp[13]) ? node5256 : 4'b0111;
															assign node5256 = (inp[10]) ? 4'b0000 : node5257;
																assign node5257 = (inp[12]) ? 4'b0111 : 4'b0000;
												assign node5261 = (inp[13]) ? node5273 : node5262;
													assign node5262 = (inp[12]) ? node5270 : node5263;
														assign node5263 = (inp[10]) ? node5265 : 4'b1000;
															assign node5265 = (inp[7]) ? 4'b1000 : node5266;
																assign node5266 = (inp[4]) ? 4'b1100 : 4'b1000;
														assign node5270 = (inp[4]) ? 4'b1000 : 4'b0000;
													assign node5273 = (inp[7]) ? node5275 : 4'b0100;
														assign node5275 = (inp[10]) ? node5279 : node5276;
															assign node5276 = (inp[4]) ? 4'b1000 : 4'b0000;
															assign node5279 = (inp[4]) ? 4'b0100 : 4'b0000;
										assign node5282 = (inp[2]) ? node5336 : node5283;
											assign node5283 = (inp[3]) ? node5309 : node5284;
												assign node5284 = (inp[4]) ? node5302 : node5285;
													assign node5285 = (inp[12]) ? node5289 : node5286;
														assign node5286 = (inp[13]) ? 4'b0101 : 4'b1101;
														assign node5289 = (inp[7]) ? node5295 : node5290;
															assign node5290 = (inp[10]) ? 4'b0001 : node5291;
																assign node5291 = (inp[13]) ? 4'b1101 : 4'b0101;
															assign node5295 = (inp[13]) ? node5299 : node5296;
																assign node5296 = (inp[10]) ? 4'b1101 : 4'b0101;
																assign node5299 = (inp[10]) ? 4'b0101 : 4'b1101;
													assign node5302 = (inp[12]) ? node5304 : 4'b0001;
														assign node5304 = (inp[7]) ? 4'b1101 : node5305;
															assign node5305 = (inp[13]) ? 4'b1001 : 4'b0001;
												assign node5309 = (inp[7]) ? node5325 : node5310;
													assign node5310 = (inp[13]) ? node5318 : node5311;
														assign node5311 = (inp[4]) ? 4'b1101 : node5312;
															assign node5312 = (inp[10]) ? 4'b1001 : node5313;
																assign node5313 = (inp[12]) ? 4'b0001 : 4'b1001;
														assign node5318 = (inp[12]) ? node5320 : 4'b0101;
															assign node5320 = (inp[10]) ? 4'b0101 : node5321;
																assign node5321 = (inp[4]) ? 4'b1101 : 4'b1001;
													assign node5325 = (inp[10]) ? node5333 : node5326;
														assign node5326 = (inp[13]) ? node5330 : node5327;
															assign node5327 = (inp[4]) ? 4'b0001 : 4'b1001;
															assign node5330 = (inp[12]) ? 4'b1001 : 4'b0001;
														assign node5333 = (inp[13]) ? 4'b0001 : 4'b1001;
											assign node5336 = (inp[3]) ? node5352 : node5337;
												assign node5337 = (inp[7]) ? node5347 : node5338;
													assign node5338 = (inp[4]) ? node5342 : node5339;
														assign node5339 = (inp[13]) ? 4'b0001 : 4'b0111;
														assign node5342 = (inp[10]) ? 4'b1001 : node5343;
															assign node5343 = (inp[13]) ? 4'b1001 : 4'b0001;
													assign node5347 = (inp[13]) ? node5349 : 4'b0111;
														assign node5349 = (inp[4]) ? 4'b0001 : 4'b0111;
												assign node5352 = (inp[4]) ? node5366 : node5353;
													assign node5353 = (inp[13]) ? node5359 : node5354;
														assign node5354 = (inp[10]) ? 4'b1001 : node5355;
															assign node5355 = (inp[12]) ? 4'b0001 : 4'b1001;
														assign node5359 = (inp[7]) ? node5361 : 4'b0101;
															assign node5361 = (inp[10]) ? 4'b0001 : node5362;
																assign node5362 = (inp[12]) ? 4'b1001 : 4'b0001;
													assign node5366 = (inp[13]) ? 4'b0101 : 4'b1101;
					assign node5370 = (inp[5]) ? node6186 : node5371;
						assign node5371 = (inp[0]) ? node5953 : node5372;
							assign node5372 = (inp[11]) ? node5700 : node5373;
								assign node5373 = (inp[10]) ? node5545 : node5374;
									assign node5374 = (inp[4]) ? node5456 : node5375;
										assign node5375 = (inp[3]) ? node5415 : node5376;
											assign node5376 = (inp[13]) ? node5388 : node5377;
												assign node5377 = (inp[12]) ? node5383 : node5378;
													assign node5378 = (inp[2]) ? node5380 : 4'b1100;
														assign node5380 = (inp[14]) ? 4'b1100 : 4'b1101;
													assign node5383 = (inp[14]) ? node5385 : 4'b0100;
														assign node5385 = (inp[1]) ? 4'b0100 : 4'b0101;
												assign node5388 = (inp[2]) ? node5400 : node5389;
													assign node5389 = (inp[7]) ? node5391 : 4'b1000;
														assign node5391 = (inp[12]) ? node5395 : node5392;
															assign node5392 = (inp[14]) ? 4'b1101 : 4'b0100;
															assign node5395 = (inp[14]) ? 4'b1100 : node5396;
																assign node5396 = (inp[1]) ? 4'b1101 : 4'b1100;
													assign node5400 = (inp[12]) ? node5408 : node5401;
														assign node5401 = (inp[1]) ? node5403 : 4'b1101;
															assign node5403 = (inp[14]) ? 4'b0100 : node5404;
																assign node5404 = (inp[7]) ? 4'b0101 : 4'b0001;
														assign node5408 = (inp[1]) ? node5412 : node5409;
															assign node5409 = (inp[14]) ? 4'b1101 : 4'b1100;
															assign node5412 = (inp[14]) ? 4'b1100 : 4'b1101;
											assign node5415 = (inp[2]) ? node5431 : node5416;
												assign node5416 = (inp[1]) ? node5426 : node5417;
													assign node5417 = (inp[12]) ? node5421 : node5418;
														assign node5418 = (inp[13]) ? 4'b1000 : 4'b1100;
														assign node5421 = (inp[13]) ? node5423 : 4'b0100;
															assign node5423 = (inp[7]) ? 4'b0100 : 4'b0000;
													assign node5426 = (inp[13]) ? node5428 : 4'b1100;
														assign node5428 = (inp[7]) ? 4'b1100 : 4'b1000;
												assign node5431 = (inp[13]) ? node5443 : node5432;
													assign node5432 = (inp[12]) ? node5438 : node5433;
														assign node5433 = (inp[1]) ? 4'b1000 : node5434;
															assign node5434 = (inp[14]) ? 4'b0001 : 4'b1000;
														assign node5438 = (inp[1]) ? 4'b0001 : node5439;
															assign node5439 = (inp[14]) ? 4'b0001 : 4'b0000;
													assign node5443 = (inp[7]) ? node5449 : node5444;
														assign node5444 = (inp[12]) ? node5446 : 4'b1000;
															assign node5446 = (inp[1]) ? 4'b1000 : 4'b0000;
														assign node5449 = (inp[12]) ? node5453 : node5450;
															assign node5450 = (inp[14]) ? 4'b0000 : 4'b0001;
															assign node5453 = (inp[1]) ? 4'b1000 : 4'b1001;
										assign node5456 = (inp[1]) ? node5504 : node5457;
											assign node5457 = (inp[13]) ? node5475 : node5458;
												assign node5458 = (inp[12]) ? node5466 : node5459;
													assign node5459 = (inp[2]) ? 4'b1100 : node5460;
														assign node5460 = (inp[14]) ? 4'b1000 : node5461;
															assign node5461 = (inp[7]) ? 4'b1000 : 4'b1001;
													assign node5466 = (inp[7]) ? node5472 : node5467;
														assign node5467 = (inp[14]) ? 4'b0000 : node5468;
															assign node5468 = (inp[2]) ? 4'b0000 : 4'b0001;
														assign node5472 = (inp[2]) ? 4'b0100 : 4'b0000;
												assign node5475 = (inp[3]) ? node5491 : node5476;
													assign node5476 = (inp[14]) ? node5486 : node5477;
														assign node5477 = (inp[2]) ? node5481 : node5478;
															assign node5478 = (inp[12]) ? 4'b0100 : 4'b1100;
															assign node5481 = (inp[12]) ? node5483 : 4'b0000;
																assign node5483 = (inp[7]) ? 4'b1100 : 4'b1000;
														assign node5486 = (inp[2]) ? node5488 : 4'b0100;
															assign node5488 = (inp[7]) ? 4'b1101 : 4'b1001;
													assign node5491 = (inp[2]) ? node5501 : node5492;
														assign node5492 = (inp[12]) ? node5498 : node5493;
															assign node5493 = (inp[14]) ? 4'b0100 : node5494;
																assign node5494 = (inp[7]) ? 4'b0001 : 4'b0101;
															assign node5498 = (inp[14]) ? 4'b1000 : 4'b1001;
														assign node5501 = (inp[7]) ? 4'b0000 : 4'b0100;
											assign node5504 = (inp[13]) ? node5524 : node5505;
												assign node5505 = (inp[7]) ? node5515 : node5506;
													assign node5506 = (inp[12]) ? node5510 : node5507;
														assign node5507 = (inp[2]) ? 4'b1000 : 4'b0000;
														assign node5510 = (inp[2]) ? node5512 : 4'b1000;
															assign node5512 = (inp[3]) ? 4'b1000 : 4'b0000;
													assign node5515 = (inp[3]) ? node5519 : node5516;
														assign node5516 = (inp[14]) ? 4'b1100 : 4'b1000;
														assign node5519 = (inp[2]) ? 4'b1000 : node5520;
															assign node5520 = (inp[14]) ? 4'b1000 : 4'b0000;
												assign node5524 = (inp[7]) ? node5532 : node5525;
													assign node5525 = (inp[2]) ? node5527 : 4'b1100;
														assign node5527 = (inp[3]) ? 4'b1100 : node5528;
															assign node5528 = (inp[12]) ? 4'b1001 : 4'b0001;
													assign node5532 = (inp[2]) ? node5538 : node5533;
														assign node5533 = (inp[3]) ? node5535 : 4'b1000;
															assign node5535 = (inp[12]) ? 4'b0000 : 4'b1000;
														assign node5538 = (inp[12]) ? node5542 : node5539;
															assign node5539 = (inp[3]) ? 4'b1000 : 4'b0000;
															assign node5542 = (inp[3]) ? 4'b1000 : 4'b1100;
									assign node5545 = (inp[12]) ? node5613 : node5546;
										assign node5546 = (inp[4]) ? node5580 : node5547;
											assign node5547 = (inp[13]) ? node5561 : node5548;
												assign node5548 = (inp[7]) ? node5554 : node5549;
													assign node5549 = (inp[2]) ? node5551 : 4'b0000;
														assign node5551 = (inp[14]) ? 4'b1100 : 4'b0000;
													assign node5554 = (inp[2]) ? node5558 : node5555;
														assign node5555 = (inp[3]) ? 4'b0100 : 4'b1100;
														assign node5558 = (inp[3]) ? 4'b1000 : 4'b1101;
												assign node5561 = (inp[7]) ? node5575 : node5562;
													assign node5562 = (inp[14]) ? node5564 : 4'b0001;
														assign node5564 = (inp[2]) ? node5570 : node5565;
															assign node5565 = (inp[3]) ? node5567 : 4'b0000;
																assign node5567 = (inp[1]) ? 4'b0001 : 4'b0000;
															assign node5570 = (inp[1]) ? 4'b0000 : node5571;
																assign node5571 = (inp[3]) ? 4'b0000 : 4'b0001;
													assign node5575 = (inp[2]) ? node5577 : 4'b0000;
														assign node5577 = (inp[14]) ? 4'b0000 : 4'b0100;
											assign node5580 = (inp[13]) ? node5598 : node5581;
												assign node5581 = (inp[3]) ? node5589 : node5582;
													assign node5582 = (inp[2]) ? node5584 : 4'b0100;
														assign node5584 = (inp[7]) ? node5586 : 4'b1000;
															assign node5586 = (inp[14]) ? 4'b1100 : 4'b1101;
													assign node5589 = (inp[2]) ? node5595 : node5590;
														assign node5590 = (inp[1]) ? 4'b1000 : node5591;
															assign node5591 = (inp[14]) ? 4'b0000 : 4'b0001;
														assign node5595 = (inp[7]) ? 4'b0000 : 4'b0100;
												assign node5598 = (inp[3]) ? node5606 : node5599;
													assign node5599 = (inp[2]) ? node5601 : 4'b0100;
														assign node5601 = (inp[1]) ? node5603 : 4'b0000;
															assign node5603 = (inp[14]) ? 4'b0000 : 4'b0001;
													assign node5606 = (inp[2]) ? 4'b0100 : node5607;
														assign node5607 = (inp[1]) ? node5609 : 4'b1100;
															assign node5609 = (inp[14]) ? 4'b0101 : 4'b0100;
										assign node5613 = (inp[1]) ? node5653 : node5614;
											assign node5614 = (inp[4]) ? node5630 : node5615;
												assign node5615 = (inp[14]) ? node5625 : node5616;
													assign node5616 = (inp[3]) ? node5618 : 4'b1100;
														assign node5618 = (inp[2]) ? 4'b1000 : node5619;
															assign node5619 = (inp[7]) ? 4'b1100 : node5620;
																assign node5620 = (inp[13]) ? 4'b1000 : 4'b1100;
													assign node5625 = (inp[3]) ? 4'b1100 : node5626;
														assign node5626 = (inp[2]) ? 4'b0101 : 4'b1101;
												assign node5630 = (inp[13]) ? node5640 : node5631;
													assign node5631 = (inp[14]) ? node5635 : node5632;
														assign node5632 = (inp[3]) ? 4'b0001 : 4'b1000;
														assign node5635 = (inp[3]) ? node5637 : 4'b0001;
															assign node5637 = (inp[2]) ? 4'b1000 : 4'b0000;
													assign node5640 = (inp[3]) ? node5650 : node5641;
														assign node5641 = (inp[14]) ? node5645 : node5642;
															assign node5642 = (inp[2]) ? 4'b0000 : 4'b1000;
															assign node5645 = (inp[2]) ? node5647 : 4'b1000;
																assign node5647 = (inp[7]) ? 4'b1101 : 4'b1001;
														assign node5650 = (inp[7]) ? 4'b1000 : 4'b1100;
											assign node5653 = (inp[13]) ? node5681 : node5654;
												assign node5654 = (inp[3]) ? node5670 : node5655;
													assign node5655 = (inp[2]) ? node5665 : node5656;
														assign node5656 = (inp[7]) ? node5660 : node5657;
															assign node5657 = (inp[4]) ? 4'b0100 : 4'b0000;
															assign node5660 = (inp[4]) ? 4'b0000 : node5661;
																assign node5661 = (inp[14]) ? 4'b1100 : 4'b1101;
														assign node5665 = (inp[7]) ? 4'b1100 : node5666;
															assign node5666 = (inp[14]) ? 4'b1000 : 4'b1001;
													assign node5670 = (inp[2]) ? node5676 : node5671;
														assign node5671 = (inp[14]) ? node5673 : 4'b1000;
															assign node5673 = (inp[7]) ? 4'b0100 : 4'b0000;
														assign node5676 = (inp[7]) ? 4'b0000 : node5677;
															assign node5677 = (inp[4]) ? 4'b0100 : 4'b0000;
												assign node5681 = (inp[4]) ? node5691 : node5682;
													assign node5682 = (inp[2]) ? node5684 : 4'b0000;
														assign node5684 = (inp[7]) ? node5688 : node5685;
															assign node5685 = (inp[3]) ? 4'b0000 : 4'b0001;
															assign node5688 = (inp[14]) ? 4'b0100 : 4'b0101;
													assign node5691 = (inp[3]) ? node5695 : node5692;
														assign node5692 = (inp[2]) ? 4'b0001 : 4'b0100;
														assign node5695 = (inp[2]) ? 4'b0100 : node5696;
															assign node5696 = (inp[7]) ? 4'b1001 : 4'b1101;
								assign node5700 = (inp[1]) ? node5848 : node5701;
									assign node5701 = (inp[2]) ? node5781 : node5702;
										assign node5702 = (inp[4]) ? node5728 : node5703;
											assign node5703 = (inp[13]) ? node5717 : node5704;
												assign node5704 = (inp[3]) ? node5712 : node5705;
													assign node5705 = (inp[10]) ? node5707 : 4'b1100;
														assign node5707 = (inp[12]) ? 4'b1100 : node5708;
															assign node5708 = (inp[14]) ? 4'b0001 : 4'b1100;
													assign node5712 = (inp[12]) ? node5714 : 4'b1101;
														assign node5714 = (inp[10]) ? 4'b1101 : 4'b0101;
												assign node5717 = (inp[7]) ? node5725 : node5718;
													assign node5718 = (inp[12]) ? node5722 : node5719;
														assign node5719 = (inp[3]) ? 4'b0000 : 4'b0001;
														assign node5722 = (inp[10]) ? 4'b1001 : 4'b0001;
													assign node5725 = (inp[3]) ? 4'b1101 : 4'b0100;
											assign node5728 = (inp[3]) ? node5758 : node5729;
												assign node5729 = (inp[7]) ? node5739 : node5730;
													assign node5730 = (inp[13]) ? node5734 : node5731;
														assign node5731 = (inp[12]) ? 4'b0001 : 4'b0101;
														assign node5734 = (inp[12]) ? 4'b1101 : node5735;
															assign node5735 = (inp[10]) ? 4'b0101 : 4'b1101;
													assign node5739 = (inp[14]) ? node5745 : node5740;
														assign node5740 = (inp[12]) ? 4'b0001 : node5741;
															assign node5741 = (inp[10]) ? 4'b0001 : 4'b1001;
														assign node5745 = (inp[13]) ? node5753 : node5746;
															assign node5746 = (inp[12]) ? node5750 : node5747;
																assign node5747 = (inp[10]) ? 4'b0001 : 4'b1001;
																assign node5750 = (inp[10]) ? 4'b1001 : 4'b0001;
															assign node5753 = (inp[10]) ? node5755 : 4'b1001;
																assign node5755 = (inp[12]) ? 4'b1001 : 4'b0101;
												assign node5758 = (inp[13]) ? node5770 : node5759;
													assign node5759 = (inp[12]) ? node5763 : node5760;
														assign node5760 = (inp[10]) ? 4'b1000 : 4'b1001;
														assign node5763 = (inp[7]) ? node5767 : node5764;
															assign node5764 = (inp[10]) ? 4'b0000 : 4'b1000;
															assign node5767 = (inp[10]) ? 4'b0000 : 4'b0001;
													assign node5770 = (inp[12]) ? node5776 : node5771;
														assign node5771 = (inp[7]) ? node5773 : 4'b0100;
															assign node5773 = (inp[10]) ? 4'b0100 : 4'b0000;
														assign node5776 = (inp[7]) ? node5778 : 4'b1100;
															assign node5778 = (inp[14]) ? 4'b0000 : 4'b1000;
										assign node5781 = (inp[3]) ? node5807 : node5782;
											assign node5782 = (inp[7]) ? node5796 : node5783;
												assign node5783 = (inp[13]) ? node5789 : node5784;
													assign node5784 = (inp[10]) ? 4'b1000 : node5785;
														assign node5785 = (inp[12]) ? 4'b0000 : 4'b1000;
													assign node5789 = (inp[12]) ? node5791 : 4'b0000;
														assign node5791 = (inp[10]) ? 4'b0000 : node5792;
															assign node5792 = (inp[4]) ? 4'b1000 : 4'b1100;
												assign node5796 = (inp[13]) ? node5798 : 4'b1100;
													assign node5798 = (inp[10]) ? node5804 : node5799;
														assign node5799 = (inp[12]) ? 4'b1100 : node5800;
															assign node5800 = (inp[4]) ? 4'b0000 : 4'b0100;
														assign node5804 = (inp[4]) ? 4'b0000 : 4'b0100;
											assign node5807 = (inp[4]) ? node5825 : node5808;
												assign node5808 = (inp[7]) ? node5820 : node5809;
													assign node5809 = (inp[12]) ? node5813 : node5810;
														assign node5810 = (inp[10]) ? 4'b0001 : 4'b1001;
														assign node5813 = (inp[13]) ? node5817 : node5814;
															assign node5814 = (inp[10]) ? 4'b1000 : 4'b0000;
															assign node5817 = (inp[10]) ? 4'b1001 : 4'b0001;
													assign node5820 = (inp[12]) ? node5822 : 4'b1000;
														assign node5822 = (inp[13]) ? 4'b1000 : 4'b0000;
												assign node5825 = (inp[13]) ? node5835 : node5826;
													assign node5826 = (inp[12]) ? node5832 : node5827;
														assign node5827 = (inp[10]) ? node5829 : 4'b1001;
															assign node5829 = (inp[7]) ? 4'b0001 : 4'b0101;
														assign node5832 = (inp[10]) ? 4'b1001 : 4'b0001;
													assign node5835 = (inp[7]) ? node5845 : node5836;
														assign node5836 = (inp[14]) ? 4'b1101 : node5837;
															assign node5837 = (inp[12]) ? node5841 : node5838;
																assign node5838 = (inp[10]) ? 4'b0101 : 4'b1101;
																assign node5841 = (inp[10]) ? 4'b1101 : 4'b0101;
														assign node5845 = (inp[12]) ? 4'b0001 : 4'b1001;
									assign node5848 = (inp[10]) ? node5910 : node5849;
										assign node5849 = (inp[4]) ? node5879 : node5850;
											assign node5850 = (inp[2]) ? node5862 : node5851;
												assign node5851 = (inp[7]) ? node5855 : node5852;
													assign node5852 = (inp[13]) ? 4'b1001 : 4'b1101;
													assign node5855 = (inp[3]) ? 4'b1101 : node5856;
														assign node5856 = (inp[13]) ? 4'b0101 : node5857;
															assign node5857 = (inp[12]) ? 4'b0101 : 4'b1101;
												assign node5862 = (inp[3]) ? node5870 : node5863;
													assign node5863 = (inp[14]) ? node5865 : 4'b1101;
														assign node5865 = (inp[12]) ? node5867 : 4'b0001;
															assign node5867 = (inp[13]) ? 4'b1101 : 4'b0101;
													assign node5870 = (inp[12]) ? node5876 : node5871;
														assign node5871 = (inp[13]) ? node5873 : 4'b1001;
															assign node5873 = (inp[7]) ? 4'b0001 : 4'b1001;
														assign node5876 = (inp[13]) ? 4'b1001 : 4'b0001;
											assign node5879 = (inp[13]) ? node5895 : node5880;
												assign node5880 = (inp[2]) ? node5886 : node5881;
													assign node5881 = (inp[12]) ? 4'b1001 : node5882;
														assign node5882 = (inp[3]) ? 4'b0001 : 4'b1001;
													assign node5886 = (inp[7]) ? node5892 : node5887;
														assign node5887 = (inp[12]) ? node5889 : 4'b1001;
															assign node5889 = (inp[3]) ? 4'b1001 : 4'b0001;
														assign node5892 = (inp[3]) ? 4'b1001 : 4'b1101;
												assign node5895 = (inp[7]) ? node5903 : node5896;
													assign node5896 = (inp[2]) ? node5898 : 4'b1101;
														assign node5898 = (inp[3]) ? 4'b1101 : node5899;
															assign node5899 = (inp[12]) ? 4'b1001 : 4'b0001;
													assign node5903 = (inp[2]) ? node5907 : node5904;
														assign node5904 = (inp[3]) ? 4'b0001 : 4'b1001;
														assign node5907 = (inp[3]) ? 4'b1001 : 4'b1101;
										assign node5910 = (inp[13]) ? node5940 : node5911;
											assign node5911 = (inp[7]) ? node5927 : node5912;
												assign node5912 = (inp[4]) ? node5914 : 4'b0001;
													assign node5914 = (inp[12]) ? node5918 : node5915;
														assign node5915 = (inp[2]) ? 4'b1001 : 4'b0101;
														assign node5918 = (inp[14]) ? 4'b0101 : node5919;
															assign node5919 = (inp[3]) ? node5923 : node5920;
																assign node5920 = (inp[2]) ? 4'b1001 : 4'b0101;
																assign node5923 = (inp[2]) ? 4'b0101 : 4'b1001;
												assign node5927 = (inp[4]) ? node5933 : node5928;
													assign node5928 = (inp[3]) ? node5930 : 4'b1101;
														assign node5930 = (inp[2]) ? 4'b1001 : 4'b0101;
													assign node5933 = (inp[2]) ? node5937 : node5934;
														assign node5934 = (inp[3]) ? 4'b1001 : 4'b0001;
														assign node5937 = (inp[3]) ? 4'b0001 : 4'b1101;
											assign node5940 = (inp[4]) ? node5948 : node5941;
												assign node5941 = (inp[7]) ? node5943 : 4'b0001;
													assign node5943 = (inp[3]) ? 4'b0001 : node5944;
														assign node5944 = (inp[2]) ? 4'b0101 : 4'b0001;
												assign node5948 = (inp[2]) ? node5950 : 4'b0101;
													assign node5950 = (inp[3]) ? 4'b0101 : 4'b0001;
							assign node5953 = (inp[2]) ? 4'b0101 : node5954;
								assign node5954 = (inp[3]) ? node6044 : node5955;
									assign node5955 = (inp[7]) ? node6019 : node5956;
										assign node5956 = (inp[4]) ? node5978 : node5957;
											assign node5957 = (inp[13]) ? node5959 : 4'b0101;
												assign node5959 = (inp[10]) ? node5969 : node5960;
													assign node5960 = (inp[12]) ? 4'b0101 : node5961;
														assign node5961 = (inp[14]) ? node5965 : node5962;
															assign node5962 = (inp[1]) ? 4'b0001 : 4'b0000;
															assign node5965 = (inp[11]) ? 4'b0001 : 4'b0101;
													assign node5969 = (inp[1]) ? node5975 : node5970;
														assign node5970 = (inp[14]) ? node5972 : 4'b0000;
															assign node5972 = (inp[11]) ? 4'b0000 : 4'b0001;
														assign node5975 = (inp[11]) ? 4'b0001 : 4'b0000;
											assign node5978 = (inp[1]) ? node6004 : node5979;
												assign node5979 = (inp[14]) ? node5989 : node5980;
													assign node5980 = (inp[13]) ? node5986 : node5981;
														assign node5981 = (inp[10]) ? 4'b1000 : node5982;
															assign node5982 = (inp[12]) ? 4'b0000 : 4'b1000;
														assign node5986 = (inp[12]) ? 4'b1000 : 4'b0000;
													assign node5989 = (inp[11]) ? node5997 : node5990;
														assign node5990 = (inp[10]) ? node5992 : 4'b1001;
															assign node5992 = (inp[13]) ? node5994 : 4'b0001;
																assign node5994 = (inp[12]) ? 4'b1001 : 4'b0001;
														assign node5997 = (inp[12]) ? node5999 : 4'b1000;
															assign node5999 = (inp[13]) ? node6001 : 4'b0000;
																assign node6001 = (inp[10]) ? 4'b0000 : 4'b1000;
												assign node6004 = (inp[13]) ? node6010 : node6005;
													assign node6005 = (inp[12]) ? node6007 : 4'b1001;
														assign node6007 = (inp[10]) ? 4'b1001 : 4'b0001;
													assign node6010 = (inp[11]) ? 4'b0001 : node6011;
														assign node6011 = (inp[10]) ? node6015 : node6012;
															assign node6012 = (inp[14]) ? 4'b1000 : 4'b1001;
															assign node6015 = (inp[14]) ? 4'b0000 : 4'b0001;
										assign node6019 = (inp[4]) ? node6021 : 4'b0101;
											assign node6021 = (inp[13]) ? node6023 : 4'b0101;
												assign node6023 = (inp[10]) ? node6031 : node6024;
													assign node6024 = (inp[12]) ? 4'b0101 : node6025;
														assign node6025 = (inp[1]) ? 4'b0001 : node6026;
															assign node6026 = (inp[11]) ? 4'b0000 : 4'b0101;
													assign node6031 = (inp[1]) ? node6039 : node6032;
														assign node6032 = (inp[14]) ? node6034 : 4'b0000;
															assign node6034 = (inp[11]) ? 4'b0000 : node6035;
																assign node6035 = (inp[12]) ? 4'b0101 : 4'b0001;
														assign node6039 = (inp[14]) ? node6041 : 4'b0001;
															assign node6041 = (inp[11]) ? 4'b0001 : 4'b0000;
									assign node6044 = (inp[7]) ? node6116 : node6045;
										assign node6045 = (inp[4]) ? node6085 : node6046;
											assign node6046 = (inp[13]) ? node6072 : node6047;
												assign node6047 = (inp[10]) ? node6063 : node6048;
													assign node6048 = (inp[12]) ? node6054 : node6049;
														assign node6049 = (inp[11]) ? 4'b1000 : node6050;
															assign node6050 = (inp[14]) ? 4'b0001 : 4'b1001;
														assign node6054 = (inp[11]) ? 4'b0001 : node6055;
															assign node6055 = (inp[14]) ? node6059 : node6056;
																assign node6056 = (inp[1]) ? 4'b0001 : 4'b0000;
																assign node6059 = (inp[1]) ? 4'b0000 : 4'b0001;
													assign node6063 = (inp[1]) ? node6067 : node6064;
														assign node6064 = (inp[12]) ? 4'b0001 : 4'b1001;
														assign node6067 = (inp[14]) ? node6069 : 4'b1001;
															assign node6069 = (inp[11]) ? 4'b1001 : 4'b1000;
												assign node6072 = (inp[11]) ? node6082 : node6073;
													assign node6073 = (inp[1]) ? node6077 : node6074;
														assign node6074 = (inp[14]) ? 4'b1001 : 4'b0100;
														assign node6077 = (inp[14]) ? 4'b0100 : node6078;
															assign node6078 = (inp[12]) ? 4'b1001 : 4'b0101;
													assign node6082 = (inp[1]) ? 4'b0101 : 4'b0100;
											assign node6085 = (inp[1]) ? node6101 : node6086;
												assign node6086 = (inp[14]) ? node6092 : node6087;
													assign node6087 = (inp[13]) ? node6089 : 4'b1100;
														assign node6089 = (inp[12]) ? 4'b1100 : 4'b0100;
													assign node6092 = (inp[11]) ? node6098 : node6093;
														assign node6093 = (inp[13]) ? node6095 : 4'b0101;
															assign node6095 = (inp[10]) ? 4'b0101 : 4'b1101;
														assign node6098 = (inp[12]) ? 4'b1100 : 4'b0100;
												assign node6101 = (inp[11]) ? node6111 : node6102;
													assign node6102 = (inp[14]) ? node6106 : node6103;
														assign node6103 = (inp[12]) ? 4'b0101 : 4'b1101;
														assign node6106 = (inp[13]) ? node6108 : 4'b1100;
															assign node6108 = (inp[10]) ? 4'b0100 : 4'b1100;
													assign node6111 = (inp[13]) ? 4'b0101 : node6112;
														assign node6112 = (inp[10]) ? 4'b1101 : 4'b0101;
										assign node6116 = (inp[13]) ? node6150 : node6117;
											assign node6117 = (inp[12]) ? node6131 : node6118;
												assign node6118 = (inp[1]) ? node6126 : node6119;
													assign node6119 = (inp[14]) ? node6121 : 4'b1000;
														assign node6121 = (inp[11]) ? 4'b1000 : node6122;
															assign node6122 = (inp[10]) ? 4'b1001 : 4'b0001;
													assign node6126 = (inp[14]) ? node6128 : 4'b1001;
														assign node6128 = (inp[11]) ? 4'b1001 : 4'b1000;
												assign node6131 = (inp[10]) ? node6141 : node6132;
													assign node6132 = (inp[4]) ? 4'b0001 : node6133;
														assign node6133 = (inp[1]) ? node6137 : node6134;
															assign node6134 = (inp[14]) ? 4'b0001 : 4'b0000;
															assign node6137 = (inp[14]) ? 4'b0000 : 4'b0001;
													assign node6141 = (inp[1]) ? node6147 : node6142;
														assign node6142 = (inp[11]) ? 4'b1000 : node6143;
															assign node6143 = (inp[14]) ? 4'b0001 : 4'b1000;
														assign node6147 = (inp[14]) ? 4'b1000 : 4'b1001;
											assign node6150 = (inp[12]) ? node6166 : node6151;
												assign node6151 = (inp[4]) ? node6159 : node6152;
													assign node6152 = (inp[1]) ? 4'b0001 : node6153;
														assign node6153 = (inp[14]) ? node6155 : 4'b0000;
															assign node6155 = (inp[10]) ? 4'b0001 : 4'b1001;
													assign node6159 = (inp[1]) ? 4'b0101 : node6160;
														assign node6160 = (inp[11]) ? 4'b0100 : node6161;
															assign node6161 = (inp[10]) ? 4'b0101 : 4'b0100;
												assign node6166 = (inp[10]) ? node6176 : node6167;
													assign node6167 = (inp[14]) ? node6169 : 4'b1001;
														assign node6169 = (inp[11]) ? node6173 : node6170;
															assign node6170 = (inp[1]) ? 4'b1000 : 4'b1001;
															assign node6173 = (inp[1]) ? 4'b1001 : 4'b1000;
													assign node6176 = (inp[4]) ? 4'b0100 : node6177;
														assign node6177 = (inp[1]) ? node6181 : node6178;
															assign node6178 = (inp[11]) ? 4'b0000 : 4'b1001;
															assign node6181 = (inp[14]) ? 4'b0000 : 4'b0001;
						assign node6186 = (inp[3]) ? node6708 : node6187;
							assign node6187 = (inp[4]) ? node6453 : node6188;
								assign node6188 = (inp[13]) ? node6326 : node6189;
									assign node6189 = (inp[7]) ? node6255 : node6190;
										assign node6190 = (inp[10]) ? node6226 : node6191;
											assign node6191 = (inp[1]) ? node6207 : node6192;
												assign node6192 = (inp[2]) ? node6202 : node6193;
													assign node6193 = (inp[11]) ? node6197 : node6194;
														assign node6194 = (inp[0]) ? 4'b0100 : 4'b0101;
														assign node6197 = (inp[0]) ? node6199 : 4'b1100;
															assign node6199 = (inp[12]) ? 4'b0100 : 4'b1100;
													assign node6202 = (inp[0]) ? 4'b0101 : node6203;
														assign node6203 = (inp[11]) ? 4'b0101 : 4'b0100;
												assign node6207 = (inp[11]) ? node6219 : node6208;
													assign node6208 = (inp[12]) ? 4'b1100 : node6209;
														assign node6209 = (inp[0]) ? node6215 : node6210;
															assign node6210 = (inp[2]) ? node6212 : 4'b0001;
																assign node6212 = (inp[14]) ? 4'b1100 : 4'b0000;
															assign node6215 = (inp[2]) ? 4'b0101 : 4'b1101;
													assign node6219 = (inp[2]) ? node6223 : node6220;
														assign node6220 = (inp[0]) ? 4'b0101 : 4'b0001;
														assign node6223 = (inp[12]) ? 4'b1101 : 4'b0001;
											assign node6226 = (inp[0]) ? node6246 : node6227;
												assign node6227 = (inp[11]) ? node6239 : node6228;
													assign node6228 = (inp[12]) ? node6232 : node6229;
														assign node6229 = (inp[14]) ? 4'b1001 : 4'b0001;
														assign node6232 = (inp[2]) ? node6234 : 4'b0001;
															assign node6234 = (inp[1]) ? 4'b0001 : node6235;
																assign node6235 = (inp[14]) ? 4'b0000 : 4'b0001;
													assign node6239 = (inp[1]) ? node6243 : node6240;
														assign node6240 = (inp[2]) ? 4'b1000 : 4'b1001;
														assign node6243 = (inp[2]) ? 4'b1001 : 4'b0001;
												assign node6246 = (inp[2]) ? 4'b0101 : node6247;
													assign node6247 = (inp[11]) ? node6249 : 4'b0000;
														assign node6249 = (inp[1]) ? 4'b0001 : node6250;
															assign node6250 = (inp[12]) ? 4'b1100 : 4'b0001;
										assign node6255 = (inp[2]) ? node6305 : node6256;
											assign node6256 = (inp[1]) ? node6282 : node6257;
												assign node6257 = (inp[11]) ? node6275 : node6258;
													assign node6258 = (inp[12]) ? node6268 : node6259;
														assign node6259 = (inp[10]) ? node6265 : node6260;
															assign node6260 = (inp[0]) ? node6262 : 4'b1100;
																assign node6262 = (inp[14]) ? 4'b0101 : 4'b1100;
															assign node6265 = (inp[0]) ? 4'b1100 : 4'b0101;
														assign node6268 = (inp[0]) ? node6270 : 4'b0101;
															assign node6270 = (inp[14]) ? 4'b0101 : node6271;
																assign node6271 = (inp[10]) ? 4'b1100 : 4'b0100;
													assign node6275 = (inp[10]) ? node6279 : node6276;
														assign node6276 = (inp[0]) ? 4'b0100 : 4'b1100;
														assign node6279 = (inp[0]) ? 4'b1100 : 4'b0100;
												assign node6282 = (inp[0]) ? node6298 : node6283;
													assign node6283 = (inp[14]) ? node6293 : node6284;
														assign node6284 = (inp[11]) ? node6290 : node6285;
															assign node6285 = (inp[12]) ? 4'b1100 : node6286;
																assign node6286 = (inp[10]) ? 4'b0001 : 4'b0100;
															assign node6290 = (inp[12]) ? 4'b0001 : 4'b0101;
														assign node6293 = (inp[12]) ? node6295 : 4'b0101;
															assign node6295 = (inp[10]) ? 4'b0101 : 4'b1101;
													assign node6298 = (inp[12]) ? 4'b0101 : node6299;
														assign node6299 = (inp[11]) ? 4'b1101 : node6300;
															assign node6300 = (inp[14]) ? 4'b1100 : 4'b1101;
											assign node6305 = (inp[0]) ? 4'b0101 : node6306;
												assign node6306 = (inp[11]) ? node6318 : node6307;
													assign node6307 = (inp[1]) ? node6315 : node6308;
														assign node6308 = (inp[14]) ? node6310 : 4'b0100;
															assign node6310 = (inp[12]) ? node6312 : 4'b1100;
																assign node6312 = (inp[10]) ? 4'b1100 : 4'b0100;
														assign node6315 = (inp[10]) ? 4'b0100 : 4'b1100;
													assign node6318 = (inp[10]) ? 4'b0101 : node6319;
														assign node6319 = (inp[1]) ? 4'b1101 : node6320;
															assign node6320 = (inp[12]) ? 4'b0101 : 4'b1101;
									assign node6326 = (inp[0]) ? node6384 : node6327;
										assign node6327 = (inp[1]) ? node6351 : node6328;
											assign node6328 = (inp[2]) ? node6338 : node6329;
												assign node6329 = (inp[10]) ? node6335 : node6330;
													assign node6330 = (inp[11]) ? 4'b1001 : node6331;
														assign node6331 = (inp[12]) ? 4'b0001 : 4'b1001;
													assign node6335 = (inp[7]) ? 4'b1001 : 4'b1101;
												assign node6338 = (inp[11]) ? node6346 : node6339;
													assign node6339 = (inp[14]) ? 4'b1000 : node6340;
														assign node6340 = (inp[10]) ? 4'b1001 : node6341;
															assign node6341 = (inp[7]) ? 4'b0001 : 4'b1001;
													assign node6346 = (inp[10]) ? node6348 : 4'b0000;
														assign node6348 = (inp[14]) ? 4'b0100 : 4'b1000;
											assign node6351 = (inp[2]) ? node6369 : node6352;
												assign node6352 = (inp[12]) ? node6358 : node6353;
													assign node6353 = (inp[11]) ? node6355 : 4'b0101;
														assign node6355 = (inp[14]) ? 4'b0101 : 4'b0001;
													assign node6358 = (inp[11]) ? node6364 : node6359;
														assign node6359 = (inp[7]) ? 4'b1001 : node6360;
															assign node6360 = (inp[10]) ? 4'b1101 : 4'b1001;
														assign node6364 = (inp[7]) ? node6366 : 4'b0101;
															assign node6366 = (inp[10]) ? 4'b0101 : 4'b0001;
												assign node6369 = (inp[11]) ? node6377 : node6370;
													assign node6370 = (inp[14]) ? node6374 : node6371;
														assign node6371 = (inp[7]) ? 4'b0000 : 4'b1000;
														assign node6374 = (inp[12]) ? 4'b1001 : 4'b0001;
													assign node6377 = (inp[10]) ? node6381 : node6378;
														assign node6378 = (inp[12]) ? 4'b0001 : 4'b1001;
														assign node6381 = (inp[7]) ? 4'b0001 : 4'b0101;
										assign node6384 = (inp[7]) ? node6428 : node6385;
											assign node6385 = (inp[2]) ? node6411 : node6386;
												assign node6386 = (inp[11]) ? node6402 : node6387;
													assign node6387 = (inp[14]) ? node6395 : node6388;
														assign node6388 = (inp[1]) ? 4'b0000 : node6389;
															assign node6389 = (inp[12]) ? node6391 : 4'b0000;
																assign node6391 = (inp[10]) ? 4'b1000 : 4'b0000;
														assign node6395 = (inp[10]) ? node6397 : 4'b1000;
															assign node6397 = (inp[1]) ? 4'b0000 : node6398;
																assign node6398 = (inp[12]) ? 4'b1000 : 4'b0000;
													assign node6402 = (inp[1]) ? node6408 : node6403;
														assign node6403 = (inp[12]) ? node6405 : 4'b0001;
															assign node6405 = (inp[10]) ? 4'b1001 : 4'b0001;
														assign node6408 = (inp[10]) ? 4'b0001 : 4'b1001;
												assign node6411 = (inp[12]) ? node6421 : node6412;
													assign node6412 = (inp[11]) ? 4'b0001 : node6413;
														assign node6413 = (inp[10]) ? node6415 : 4'b0000;
															assign node6415 = (inp[1]) ? 4'b0001 : node6416;
																assign node6416 = (inp[14]) ? 4'b0001 : 4'b0000;
													assign node6421 = (inp[10]) ? node6423 : 4'b0101;
														assign node6423 = (inp[11]) ? 4'b0000 : node6424;
															assign node6424 = (inp[1]) ? 4'b0000 : 4'b0101;
											assign node6428 = (inp[2]) ? 4'b0101 : node6429;
												assign node6429 = (inp[10]) ? node6441 : node6430;
													assign node6430 = (inp[12]) ? node6438 : node6431;
														assign node6431 = (inp[14]) ? node6433 : 4'b0100;
															assign node6433 = (inp[1]) ? 4'b0100 : node6434;
																assign node6434 = (inp[11]) ? 4'b0100 : 4'b1101;
														assign node6438 = (inp[11]) ? 4'b1101 : 4'b1100;
													assign node6441 = (inp[1]) ? node6449 : node6442;
														assign node6442 = (inp[12]) ? node6444 : 4'b0001;
															assign node6444 = (inp[11]) ? 4'b0100 : node6445;
																assign node6445 = (inp[14]) ? 4'b1101 : 4'b0100;
														assign node6449 = (inp[11]) ? 4'b0001 : 4'b0000;
								assign node6453 = (inp[11]) ? node6605 : node6454;
									assign node6454 = (inp[2]) ? node6542 : node6455;
										assign node6455 = (inp[10]) ? node6487 : node6456;
											assign node6456 = (inp[0]) ? node6472 : node6457;
												assign node6457 = (inp[13]) ? node6467 : node6458;
													assign node6458 = (inp[1]) ? node6464 : node6459;
														assign node6459 = (inp[7]) ? node6461 : 4'b1001;
															assign node6461 = (inp[12]) ? 4'b0101 : 4'b1101;
														assign node6464 = (inp[14]) ? 4'b0000 : 4'b0001;
													assign node6467 = (inp[7]) ? node6469 : 4'b1000;
														assign node6469 = (inp[12]) ? 4'b0000 : 4'b1000;
												assign node6472 = (inp[1]) ? node6482 : node6473;
													assign node6473 = (inp[12]) ? node6477 : node6474;
														assign node6474 = (inp[13]) ? 4'b0001 : 4'b1000;
														assign node6477 = (inp[13]) ? node6479 : 4'b0000;
															assign node6479 = (inp[7]) ? 4'b0000 : 4'b0100;
													assign node6482 = (inp[13]) ? node6484 : 4'b1000;
														assign node6484 = (inp[7]) ? 4'b1000 : 4'b0001;
											assign node6487 = (inp[12]) ? node6517 : node6488;
												assign node6488 = (inp[0]) ? node6508 : node6489;
													assign node6489 = (inp[13]) ? node6501 : node6490;
														assign node6490 = (inp[14]) ? node6498 : node6491;
															assign node6491 = (inp[1]) ? node6495 : node6492;
																assign node6492 = (inp[7]) ? 4'b0000 : 4'b0100;
																assign node6495 = (inp[7]) ? 4'b1001 : 4'b0000;
															assign node6498 = (inp[7]) ? 4'b1000 : 4'b1001;
														assign node6501 = (inp[7]) ? 4'b0100 : node6502;
															assign node6502 = (inp[14]) ? 4'b0000 : node6503;
																assign node6503 = (inp[1]) ? 4'b0000 : 4'b0001;
													assign node6508 = (inp[13]) ? node6512 : node6509;
														assign node6509 = (inp[7]) ? 4'b0000 : 4'b0100;
														assign node6512 = (inp[1]) ? 4'b0001 : node6513;
															assign node6513 = (inp[7]) ? 4'b0100 : 4'b1000;
												assign node6517 = (inp[7]) ? node6531 : node6518;
													assign node6518 = (inp[14]) ? node6524 : node6519;
														assign node6519 = (inp[13]) ? node6521 : 4'b1000;
															assign node6521 = (inp[1]) ? 4'b1000 : 4'b0100;
														assign node6524 = (inp[1]) ? node6528 : node6525;
															assign node6525 = (inp[0]) ? 4'b1000 : 4'b1001;
															assign node6528 = (inp[13]) ? 4'b1001 : 4'b0100;
													assign node6531 = (inp[0]) ? node6537 : node6532;
														assign node6532 = (inp[13]) ? node6534 : 4'b0001;
															assign node6534 = (inp[1]) ? 4'b1000 : 4'b0000;
														assign node6537 = (inp[1]) ? node6539 : 4'b1000;
															assign node6539 = (inp[13]) ? 4'b0100 : 4'b0000;
										assign node6542 = (inp[13]) ? node6574 : node6543;
											assign node6543 = (inp[7]) ? node6557 : node6544;
												assign node6544 = (inp[0]) ? node6552 : node6545;
													assign node6545 = (inp[10]) ? 4'b0001 : node6546;
														assign node6546 = (inp[12]) ? node6548 : 4'b0001;
															assign node6548 = (inp[14]) ? 4'b1101 : 4'b1100;
													assign node6552 = (inp[10]) ? 4'b1000 : node6553;
														assign node6553 = (inp[1]) ? 4'b0001 : 4'b1000;
												assign node6557 = (inp[0]) ? 4'b0101 : node6558;
													assign node6558 = (inp[10]) ? node6568 : node6559;
														assign node6559 = (inp[12]) ? node6563 : node6560;
															assign node6560 = (inp[14]) ? 4'b1000 : 4'b0100;
															assign node6563 = (inp[1]) ? node6565 : 4'b0001;
																assign node6565 = (inp[14]) ? 4'b1001 : 4'b1000;
														assign node6568 = (inp[14]) ? node6570 : 4'b1100;
															assign node6570 = (inp[1]) ? 4'b0101 : 4'b0100;
											assign node6574 = (inp[0]) ? node6592 : node6575;
												assign node6575 = (inp[10]) ? node6585 : node6576;
													assign node6576 = (inp[12]) ? node6582 : node6577;
														assign node6577 = (inp[1]) ? node6579 : 4'b1001;
															assign node6579 = (inp[7]) ? 4'b0001 : 4'b0101;
														assign node6582 = (inp[1]) ? 4'b1001 : 4'b0001;
													assign node6585 = (inp[14]) ? node6589 : node6586;
														assign node6586 = (inp[7]) ? 4'b1001 : 4'b1000;
														assign node6589 = (inp[1]) ? 4'b1000 : 4'b0001;
												assign node6592 = (inp[10]) ? node6600 : node6593;
													assign node6593 = (inp[7]) ? 4'b0101 : node6594;
														assign node6594 = (inp[12]) ? node6596 : 4'b0000;
															assign node6596 = (inp[14]) ? 4'b1001 : 4'b1000;
													assign node6600 = (inp[12]) ? 4'b0000 : node6601;
														assign node6601 = (inp[1]) ? 4'b0000 : 4'b0001;
									assign node6605 = (inp[1]) ? node6675 : node6606;
										assign node6606 = (inp[13]) ? node6642 : node6607;
											assign node6607 = (inp[0]) ? node6625 : node6608;
												assign node6608 = (inp[2]) ? node6616 : node6609;
													assign node6609 = (inp[12]) ? node6611 : 4'b0000;
														assign node6611 = (inp[10]) ? node6613 : 4'b1101;
															assign node6613 = (inp[7]) ? 4'b0000 : 4'b0100;
													assign node6616 = (inp[7]) ? node6620 : node6617;
														assign node6617 = (inp[10]) ? 4'b1001 : 4'b1100;
														assign node6620 = (inp[10]) ? node6622 : 4'b1000;
															assign node6622 = (inp[14]) ? 4'b1100 : 4'b0100;
												assign node6625 = (inp[2]) ? node6637 : node6626;
													assign node6626 = (inp[7]) ? node6630 : node6627;
														assign node6627 = (inp[12]) ? 4'b0001 : 4'b0101;
														assign node6630 = (inp[10]) ? node6634 : node6631;
															assign node6631 = (inp[12]) ? 4'b0001 : 4'b1001;
															assign node6634 = (inp[12]) ? 4'b1001 : 4'b0001;
													assign node6637 = (inp[7]) ? 4'b0101 : node6638;
														assign node6638 = (inp[14]) ? 4'b1000 : 4'b0000;
											assign node6642 = (inp[0]) ? node6656 : node6643;
												assign node6643 = (inp[2]) ? node6651 : node6644;
													assign node6644 = (inp[10]) ? node6648 : node6645;
														assign node6645 = (inp[12]) ? 4'b1001 : 4'b0001;
														assign node6648 = (inp[12]) ? 4'b0000 : 4'b1000;
													assign node6651 = (inp[10]) ? node6653 : 4'b1001;
														assign node6653 = (inp[7]) ? 4'b1001 : 4'b1000;
												assign node6656 = (inp[7]) ? node6668 : node6657;
													assign node6657 = (inp[12]) ? node6659 : 4'b0000;
														assign node6659 = (inp[14]) ? 4'b1000 : node6660;
															assign node6660 = (inp[10]) ? node6664 : node6661;
																assign node6661 = (inp[2]) ? 4'b1000 : 4'b0000;
																assign node6664 = (inp[2]) ? 4'b0000 : 4'b1000;
													assign node6668 = (inp[10]) ? node6670 : 4'b0001;
														assign node6670 = (inp[2]) ? 4'b0000 : node6671;
															assign node6671 = (inp[14]) ? 4'b0000 : 4'b1001;
										assign node6675 = (inp[10]) ? node6697 : node6676;
											assign node6676 = (inp[2]) ? node6686 : node6677;
												assign node6677 = (inp[12]) ? node6679 : 4'b1001;
													assign node6679 = (inp[0]) ? node6683 : node6680;
														assign node6680 = (inp[13]) ? 4'b1001 : 4'b0001;
														assign node6683 = (inp[7]) ? 4'b1001 : 4'b0001;
												assign node6686 = (inp[7]) ? node6690 : node6687;
													assign node6687 = (inp[0]) ? 4'b1001 : 4'b0001;
													assign node6690 = (inp[13]) ? 4'b0001 : node6691;
														assign node6691 = (inp[12]) ? node6693 : 4'b0101;
															assign node6693 = (inp[0]) ? 4'b0101 : 4'b1001;
											assign node6697 = (inp[13]) ? 4'b0001 : node6698;
												assign node6698 = (inp[2]) ? node6704 : node6699;
													assign node6699 = (inp[0]) ? 4'b0001 : node6700;
														assign node6700 = (inp[7]) ? 4'b1001 : 4'b0001;
													assign node6704 = (inp[7]) ? 4'b0101 : 4'b1001;
							assign node6708 = (inp[4]) ? node6988 : node6709;
								assign node6709 = (inp[1]) ? node6859 : node6710;
									assign node6710 = (inp[2]) ? node6778 : node6711;
										assign node6711 = (inp[11]) ? node6747 : node6712;
											assign node6712 = (inp[10]) ? node6728 : node6713;
												assign node6713 = (inp[13]) ? node6719 : node6714;
													assign node6714 = (inp[14]) ? 4'b1000 : node6715;
														assign node6715 = (inp[0]) ? 4'b0001 : 4'b1001;
													assign node6719 = (inp[7]) ? node6723 : node6720;
														assign node6720 = (inp[12]) ? 4'b1000 : 4'b0000;
														assign node6723 = (inp[0]) ? 4'b1001 : node6724;
															assign node6724 = (inp[12]) ? 4'b0001 : 4'b0000;
												assign node6728 = (inp[0]) ? node6740 : node6729;
													assign node6729 = (inp[12]) ? node6733 : node6730;
														assign node6730 = (inp[14]) ? 4'b0001 : 4'b0000;
														assign node6733 = (inp[7]) ? node6737 : node6734;
															assign node6734 = (inp[13]) ? 4'b1001 : 4'b0000;
															assign node6737 = (inp[13]) ? 4'b0000 : 4'b1001;
													assign node6740 = (inp[13]) ? node6744 : node6741;
														assign node6741 = (inp[14]) ? 4'b0000 : 4'b0001;
														assign node6744 = (inp[7]) ? 4'b1000 : 4'b0000;
											assign node6747 = (inp[10]) ? node6761 : node6748;
												assign node6748 = (inp[0]) ? node6752 : node6749;
													assign node6749 = (inp[14]) ? 4'b0000 : 4'b0001;
													assign node6752 = (inp[7]) ? node6758 : node6753;
														assign node6753 = (inp[12]) ? node6755 : 4'b1000;
															assign node6755 = (inp[13]) ? 4'b0000 : 4'b1000;
														assign node6758 = (inp[13]) ? 4'b1001 : 4'b1000;
												assign node6761 = (inp[7]) ? node6769 : node6762;
													assign node6762 = (inp[0]) ? node6764 : 4'b1000;
														assign node6764 = (inp[13]) ? node6766 : 4'b1001;
															assign node6766 = (inp[12]) ? 4'b0001 : 4'b1001;
													assign node6769 = (inp[0]) ? node6773 : node6770;
														assign node6770 = (inp[13]) ? 4'b1001 : 4'b0001;
														assign node6773 = (inp[13]) ? 4'b1000 : node6774;
															assign node6774 = (inp[14]) ? 4'b1000 : 4'b0000;
										assign node6778 = (inp[7]) ? node6814 : node6779;
											assign node6779 = (inp[10]) ? node6799 : node6780;
												assign node6780 = (inp[13]) ? node6794 : node6781;
													assign node6781 = (inp[14]) ? node6789 : node6782;
														assign node6782 = (inp[12]) ? 4'b0000 : node6783;
															assign node6783 = (inp[0]) ? 4'b1000 : node6784;
																assign node6784 = (inp[11]) ? 4'b0001 : 4'b1000;
														assign node6789 = (inp[0]) ? 4'b0001 : node6790;
															assign node6790 = (inp[12]) ? 4'b0001 : 4'b1001;
													assign node6794 = (inp[11]) ? 4'b0001 : node6795;
														assign node6795 = (inp[14]) ? 4'b0000 : 4'b0001;
												assign node6799 = (inp[11]) ? node6801 : 4'b0000;
													assign node6801 = (inp[0]) ? node6807 : node6802;
														assign node6802 = (inp[12]) ? node6804 : 4'b0001;
															assign node6804 = (inp[13]) ? 4'b0000 : 4'b0001;
														assign node6807 = (inp[14]) ? node6811 : node6808;
															assign node6808 = (inp[12]) ? 4'b1000 : 4'b0000;
															assign node6811 = (inp[12]) ? 4'b1001 : 4'b0001;
											assign node6814 = (inp[11]) ? node6838 : node6815;
												assign node6815 = (inp[14]) ? node6827 : node6816;
													assign node6816 = (inp[13]) ? node6822 : node6817;
														assign node6817 = (inp[10]) ? node6819 : 4'b1000;
															assign node6819 = (inp[0]) ? 4'b1000 : 4'b0000;
														assign node6822 = (inp[10]) ? 4'b1001 : node6823;
															assign node6823 = (inp[0]) ? 4'b0000 : 4'b0001;
													assign node6827 = (inp[13]) ? 4'b1001 : node6828;
														assign node6828 = (inp[12]) ? node6834 : node6829;
															assign node6829 = (inp[0]) ? node6831 : 4'b1001;
																assign node6831 = (inp[10]) ? 4'b1001 : 4'b0001;
															assign node6834 = (inp[10]) ? 4'b0000 : 4'b0001;
												assign node6838 = (inp[10]) ? node6852 : node6839;
													assign node6839 = (inp[13]) ? node6845 : node6840;
														assign node6840 = (inp[12]) ? node6842 : 4'b0000;
															assign node6842 = (inp[0]) ? 4'b0000 : 4'b1000;
														assign node6845 = (inp[14]) ? 4'b1000 : node6846;
															assign node6846 = (inp[12]) ? 4'b1000 : node6847;
																assign node6847 = (inp[0]) ? 4'b0000 : 4'b1000;
													assign node6852 = (inp[13]) ? 4'b0000 : node6853;
														assign node6853 = (inp[12]) ? 4'b0001 : node6854;
															assign node6854 = (inp[0]) ? 4'b1000 : 4'b1001;
									assign node6859 = (inp[11]) ? node6943 : node6860;
										assign node6860 = (inp[10]) ? node6900 : node6861;
											assign node6861 = (inp[7]) ? node6877 : node6862;
												assign node6862 = (inp[0]) ? node6870 : node6863;
													assign node6863 = (inp[14]) ? 4'b1001 : node6864;
														assign node6864 = (inp[13]) ? 4'b1001 : node6865;
															assign node6865 = (inp[12]) ? 4'b1001 : 4'b1000;
													assign node6870 = (inp[14]) ? 4'b1000 : node6871;
														assign node6871 = (inp[13]) ? 4'b1000 : node6872;
															assign node6872 = (inp[12]) ? 4'b0001 : 4'b1001;
												assign node6877 = (inp[13]) ? node6887 : node6878;
													assign node6878 = (inp[0]) ? node6882 : node6879;
														assign node6879 = (inp[12]) ? 4'b0001 : 4'b1001;
														assign node6882 = (inp[14]) ? node6884 : 4'b1000;
															assign node6884 = (inp[12]) ? 4'b0000 : 4'b1000;
													assign node6887 = (inp[12]) ? node6895 : node6888;
														assign node6888 = (inp[0]) ? node6890 : 4'b0000;
															assign node6890 = (inp[14]) ? node6892 : 4'b0001;
																assign node6892 = (inp[2]) ? 4'b0000 : 4'b0001;
														assign node6895 = (inp[0]) ? 4'b1001 : node6896;
															assign node6896 = (inp[2]) ? 4'b1001 : 4'b0000;
											assign node6900 = (inp[14]) ? node6920 : node6901;
												assign node6901 = (inp[7]) ? node6909 : node6902;
													assign node6902 = (inp[2]) ? node6904 : 4'b0001;
														assign node6904 = (inp[0]) ? 4'b0000 : node6905;
															assign node6905 = (inp[12]) ? 4'b0000 : 4'b1000;
													assign node6909 = (inp[12]) ? 4'b1001 : node6910;
														assign node6910 = (inp[2]) ? node6912 : 4'b1001;
															assign node6912 = (inp[13]) ? node6916 : node6913;
																assign node6913 = (inp[0]) ? 4'b1001 : 4'b0000;
																assign node6916 = (inp[0]) ? 4'b0000 : 4'b1001;
												assign node6920 = (inp[12]) ? node6930 : node6921;
													assign node6921 = (inp[0]) ? node6925 : node6922;
														assign node6922 = (inp[13]) ? 4'b1000 : 4'b0000;
														assign node6925 = (inp[13]) ? 4'b0000 : node6926;
															assign node6926 = (inp[7]) ? 4'b1000 : 4'b0000;
													assign node6930 = (inp[13]) ? node6938 : node6931;
														assign node6931 = (inp[0]) ? 4'b0001 : node6932;
															assign node6932 = (inp[7]) ? node6934 : 4'b0001;
																assign node6934 = (inp[2]) ? 4'b1000 : 4'b0000;
														assign node6938 = (inp[7]) ? 4'b0000 : node6939;
															assign node6939 = (inp[0]) ? 4'b1000 : 4'b0000;
										assign node6943 = (inp[13]) ? node6973 : node6944;
											assign node6944 = (inp[2]) ? node6958 : node6945;
												assign node6945 = (inp[7]) ? node6947 : 4'b0001;
													assign node6947 = (inp[12]) ? node6951 : node6948;
														assign node6948 = (inp[10]) ? 4'b1001 : 4'b0001;
														assign node6951 = (inp[14]) ? node6953 : 4'b1001;
															assign node6953 = (inp[10]) ? 4'b0001 : node6954;
																assign node6954 = (inp[0]) ? 4'b1001 : 4'b0001;
												assign node6958 = (inp[12]) ? node6964 : node6959;
													assign node6959 = (inp[10]) ? node6961 : 4'b1001;
														assign node6961 = (inp[7]) ? 4'b0001 : 4'b1001;
													assign node6964 = (inp[7]) ? node6968 : node6965;
														assign node6965 = (inp[0]) ? 4'b0001 : 4'b1001;
														assign node6968 = (inp[10]) ? node6970 : 4'b0001;
															assign node6970 = (inp[0]) ? 4'b1001 : 4'b0001;
											assign node6973 = (inp[10]) ? 4'b0001 : node6974;
												assign node6974 = (inp[0]) ? node6980 : node6975;
													assign node6975 = (inp[14]) ? node6977 : 4'b0001;
														assign node6977 = (inp[7]) ? 4'b1001 : 4'b0001;
													assign node6980 = (inp[7]) ? 4'b0001 : node6981;
														assign node6981 = (inp[12]) ? 4'b1001 : node6982;
															assign node6982 = (inp[2]) ? 4'b1001 : 4'b0001;
								assign node6988 = (inp[13]) ? node7154 : node6989;
									assign node6989 = (inp[1]) ? node7085 : node6990;
										assign node6990 = (inp[10]) ? node7028 : node6991;
											assign node6991 = (inp[14]) ? node7011 : node6992;
												assign node6992 = (inp[7]) ? node7002 : node6993;
													assign node6993 = (inp[11]) ? 4'b0000 : node6994;
														assign node6994 = (inp[2]) ? node6996 : 4'b1001;
															assign node6996 = (inp[0]) ? 4'b0001 : node6997;
																assign node6997 = (inp[12]) ? 4'b1001 : 4'b0001;
													assign node7002 = (inp[12]) ? node7008 : node7003;
														assign node7003 = (inp[0]) ? node7005 : 4'b0001;
															assign node7005 = (inp[11]) ? 4'b1001 : 4'b1000;
														assign node7008 = (inp[0]) ? 4'b0000 : 4'b1000;
												assign node7011 = (inp[11]) ? node7023 : node7012;
													assign node7012 = (inp[0]) ? node7018 : node7013;
														assign node7013 = (inp[7]) ? 4'b0000 : node7014;
															assign node7014 = (inp[12]) ? 4'b1000 : 4'b0001;
														assign node7018 = (inp[2]) ? node7020 : 4'b1000;
															assign node7020 = (inp[12]) ? 4'b0000 : 4'b1000;
													assign node7023 = (inp[12]) ? node7025 : 4'b1000;
														assign node7025 = (inp[7]) ? 4'b0001 : 4'b1001;
											assign node7028 = (inp[0]) ? node7050 : node7029;
												assign node7029 = (inp[11]) ? node7039 : node7030;
													assign node7030 = (inp[12]) ? node7036 : node7031;
														assign node7031 = (inp[2]) ? node7033 : 4'b0000;
															assign node7033 = (inp[14]) ? 4'b0000 : 4'b0001;
														assign node7036 = (inp[2]) ? 4'b1000 : 4'b0000;
													assign node7039 = (inp[7]) ? node7045 : node7040;
														assign node7040 = (inp[2]) ? node7042 : 4'b0001;
															assign node7042 = (inp[12]) ? 4'b1000 : 4'b0001;
														assign node7045 = (inp[2]) ? 4'b0001 : node7046;
															assign node7046 = (inp[12]) ? 4'b0001 : 4'b0000;
												assign node7050 = (inp[11]) ? node7070 : node7051;
													assign node7051 = (inp[2]) ? node7061 : node7052;
														assign node7052 = (inp[7]) ? node7056 : node7053;
															assign node7053 = (inp[12]) ? 4'b0000 : 4'b1000;
															assign node7056 = (inp[12]) ? 4'b1001 : node7057;
																assign node7057 = (inp[14]) ? 4'b0001 : 4'b0000;
														assign node7061 = (inp[12]) ? node7067 : node7062;
															assign node7062 = (inp[14]) ? 4'b1001 : node7063;
																assign node7063 = (inp[7]) ? 4'b0001 : 4'b0000;
															assign node7067 = (inp[7]) ? 4'b0000 : 4'b0001;
													assign node7070 = (inp[2]) ? node7080 : node7071;
														assign node7071 = (inp[14]) ? 4'b1000 : node7072;
															assign node7072 = (inp[7]) ? node7076 : node7073;
																assign node7073 = (inp[12]) ? 4'b0000 : 4'b1000;
																assign node7076 = (inp[12]) ? 4'b1000 : 4'b0001;
														assign node7080 = (inp[12]) ? 4'b0000 : node7081;
															assign node7081 = (inp[7]) ? 4'b1000 : 4'b0000;
										assign node7085 = (inp[11]) ? node7127 : node7086;
											assign node7086 = (inp[10]) ? node7112 : node7087;
												assign node7087 = (inp[7]) ? node7093 : node7088;
													assign node7088 = (inp[12]) ? 4'b1000 : node7089;
														assign node7089 = (inp[2]) ? 4'b0001 : 4'b0000;
													assign node7093 = (inp[12]) ? node7103 : node7094;
														assign node7094 = (inp[2]) ? node7100 : node7095;
															assign node7095 = (inp[14]) ? node7097 : 4'b1000;
																assign node7097 = (inp[0]) ? 4'b1001 : 4'b1000;
															assign node7100 = (inp[0]) ? 4'b1000 : 4'b1001;
														assign node7103 = (inp[14]) ? node7105 : 4'b0001;
															assign node7105 = (inp[2]) ? node7109 : node7106;
																assign node7106 = (inp[0]) ? 4'b0001 : 4'b0000;
																assign node7109 = (inp[0]) ? 4'b1000 : 4'b0001;
												assign node7112 = (inp[7]) ? node7122 : node7113;
													assign node7113 = (inp[12]) ? node7117 : node7114;
														assign node7114 = (inp[0]) ? 4'b0000 : 4'b0001;
														assign node7117 = (inp[14]) ? 4'b0000 : node7118;
															assign node7118 = (inp[0]) ? 4'b0001 : 4'b0000;
													assign node7122 = (inp[0]) ? node7124 : 4'b0000;
														assign node7124 = (inp[2]) ? 4'b0001 : 4'b0000;
											assign node7127 = (inp[10]) ? 4'b0001 : node7128;
												assign node7128 = (inp[14]) ? node7140 : node7129;
													assign node7129 = (inp[12]) ? 4'b0001 : node7130;
														assign node7130 = (inp[7]) ? node7134 : node7131;
															assign node7131 = (inp[0]) ? 4'b1001 : 4'b0001;
															assign node7134 = (inp[2]) ? node7136 : 4'b0001;
																assign node7136 = (inp[0]) ? 4'b0001 : 4'b1001;
													assign node7140 = (inp[12]) ? node7146 : node7141;
														assign node7141 = (inp[2]) ? 4'b0001 : node7142;
															assign node7142 = (inp[0]) ? 4'b1001 : 4'b0001;
														assign node7146 = (inp[2]) ? 4'b1001 : node7147;
															assign node7147 = (inp[7]) ? node7149 : 4'b0001;
																assign node7149 = (inp[0]) ? 4'b0001 : 4'b1001;
									assign node7154 = (inp[10]) ? node7224 : node7155;
										assign node7155 = (inp[11]) ? node7203 : node7156;
											assign node7156 = (inp[1]) ? node7192 : node7157;
												assign node7157 = (inp[12]) ? node7177 : node7158;
													assign node7158 = (inp[2]) ? node7168 : node7159;
														assign node7159 = (inp[14]) ? node7163 : node7160;
															assign node7160 = (inp[0]) ? 4'b0000 : 4'b0001;
															assign node7163 = (inp[7]) ? 4'b0001 : node7164;
																assign node7164 = (inp[0]) ? 4'b0001 : 4'b0000;
														assign node7168 = (inp[0]) ? node7170 : 4'b0000;
															assign node7170 = (inp[7]) ? node7174 : node7171;
																assign node7171 = (inp[14]) ? 4'b0000 : 4'b0001;
																assign node7174 = (inp[14]) ? 4'b0001 : 4'b0000;
													assign node7177 = (inp[2]) ? node7179 : 4'b0000;
														assign node7179 = (inp[0]) ? node7185 : node7180;
															assign node7180 = (inp[7]) ? node7182 : 4'b0000;
																assign node7182 = (inp[14]) ? 4'b0000 : 4'b0001;
															assign node7185 = (inp[7]) ? node7189 : node7186;
																assign node7186 = (inp[14]) ? 4'b0000 : 4'b0001;
																assign node7189 = (inp[14]) ? 4'b0001 : 4'b0000;
												assign node7192 = (inp[0]) ? 4'b0000 : node7193;
													assign node7193 = (inp[14]) ? 4'b0000 : node7194;
														assign node7194 = (inp[7]) ? node7198 : node7195;
															assign node7195 = (inp[2]) ? 4'b0000 : 4'b0001;
															assign node7198 = (inp[2]) ? 4'b0001 : 4'b0000;
											assign node7203 = (inp[1]) ? 4'b0001 : node7204;
												assign node7204 = (inp[12]) ? node7210 : node7205;
													assign node7205 = (inp[0]) ? 4'b0000 : node7206;
														assign node7206 = (inp[14]) ? 4'b0001 : 4'b0000;
													assign node7210 = (inp[14]) ? node7216 : node7211;
														assign node7211 = (inp[7]) ? node7213 : 4'b0001;
															assign node7213 = (inp[0]) ? 4'b0001 : 4'b0000;
														assign node7216 = (inp[2]) ? 4'b0000 : node7217;
															assign node7217 = (inp[7]) ? node7219 : 4'b0000;
																assign node7219 = (inp[0]) ? 4'b0001 : 4'b0000;
										assign node7224 = (inp[11]) ? 4'b0000 : node7225;
											assign node7225 = (inp[1]) ? 4'b0000 : node7226;
												assign node7226 = (inp[7]) ? node7238 : node7227;
													assign node7227 = (inp[0]) ? node7229 : 4'b0000;
														assign node7229 = (inp[14]) ? node7233 : node7230;
															assign node7230 = (inp[2]) ? 4'b0000 : 4'b0001;
															assign node7233 = (inp[2]) ? node7235 : 4'b0000;
																assign node7235 = (inp[12]) ? 4'b0001 : 4'b0000;
													assign node7238 = (inp[14]) ? node7248 : node7239;
														assign node7239 = (inp[12]) ? node7241 : 4'b0000;
															assign node7241 = (inp[2]) ? node7245 : node7242;
																assign node7242 = (inp[0]) ? 4'b0000 : 4'b0001;
																assign node7245 = (inp[0]) ? 4'b0001 : 4'b0000;
														assign node7248 = (inp[12]) ? node7250 : 4'b0001;
															assign node7250 = (inp[2]) ? 4'b0000 : 4'b0001;
				assign node7255 = (inp[0]) ? node8851 : node7256;
					assign node7256 = (inp[6]) ? node7702 : node7257;
						assign node7257 = (inp[5]) ? node7355 : node7258;
							assign node7258 = (inp[3]) ? node7260 : 4'b0011;
								assign node7260 = (inp[2]) ? 4'b0011 : node7261;
									assign node7261 = (inp[7]) ? node7333 : node7262;
										assign node7262 = (inp[4]) ? node7282 : node7263;
											assign node7263 = (inp[13]) ? node7265 : 4'b0011;
												assign node7265 = (inp[12]) ? node7271 : node7266;
													assign node7266 = (inp[1]) ? node7268 : 4'b0000;
														assign node7268 = (inp[11]) ? 4'b0001 : 4'b0000;
													assign node7271 = (inp[10]) ? node7273 : 4'b0011;
														assign node7273 = (inp[1]) ? node7277 : node7274;
															assign node7274 = (inp[14]) ? 4'b0011 : 4'b0000;
															assign node7277 = (inp[14]) ? node7279 : 4'b0001;
																assign node7279 = (inp[11]) ? 4'b0001 : 4'b0000;
											assign node7282 = (inp[1]) ? node7308 : node7283;
												assign node7283 = (inp[14]) ? node7295 : node7284;
													assign node7284 = (inp[13]) ? node7290 : node7285;
														assign node7285 = (inp[12]) ? node7287 : 4'b1000;
															assign node7287 = (inp[10]) ? 4'b1000 : 4'b0000;
														assign node7290 = (inp[10]) ? 4'b0000 : node7291;
															assign node7291 = (inp[12]) ? 4'b1000 : 4'b0000;
													assign node7295 = (inp[11]) ? node7303 : node7296;
														assign node7296 = (inp[13]) ? node7298 : 4'b0001;
															assign node7298 = (inp[10]) ? node7300 : 4'b1001;
																assign node7300 = (inp[12]) ? 4'b1001 : 4'b0001;
														assign node7303 = (inp[10]) ? 4'b0000 : node7304;
															assign node7304 = (inp[13]) ? 4'b1000 : 4'b0000;
												assign node7308 = (inp[13]) ? node7322 : node7309;
													assign node7309 = (inp[14]) ? node7315 : node7310;
														assign node7310 = (inp[10]) ? 4'b1001 : node7311;
															assign node7311 = (inp[12]) ? 4'b0001 : 4'b1001;
														assign node7315 = (inp[11]) ? node7319 : node7316;
															assign node7316 = (inp[10]) ? 4'b1000 : 4'b0000;
															assign node7319 = (inp[10]) ? 4'b1001 : 4'b0001;
													assign node7322 = (inp[10]) ? node7328 : node7323;
														assign node7323 = (inp[12]) ? 4'b1001 : node7324;
															assign node7324 = (inp[11]) ? 4'b0001 : 4'b0000;
														assign node7328 = (inp[11]) ? 4'b0001 : node7329;
															assign node7329 = (inp[14]) ? 4'b0000 : 4'b0001;
										assign node7333 = (inp[13]) ? node7335 : 4'b0011;
											assign node7335 = (inp[4]) ? node7337 : 4'b0011;
												assign node7337 = (inp[1]) ? node7349 : node7338;
													assign node7338 = (inp[14]) ? node7344 : node7339;
														assign node7339 = (inp[10]) ? 4'b0000 : node7340;
															assign node7340 = (inp[11]) ? 4'b0000 : 4'b0011;
														assign node7344 = (inp[12]) ? 4'b0011 : node7345;
															assign node7345 = (inp[11]) ? 4'b0000 : 4'b0011;
													assign node7349 = (inp[12]) ? node7351 : 4'b0001;
														assign node7351 = (inp[11]) ? 4'b0001 : 4'b0000;
							assign node7355 = (inp[2]) ? node7611 : node7356;
								assign node7356 = (inp[1]) ? node7474 : node7357;
									assign node7357 = (inp[14]) ? node7413 : node7358;
										assign node7358 = (inp[13]) ? node7386 : node7359;
											assign node7359 = (inp[3]) ? node7373 : node7360;
												assign node7360 = (inp[7]) ? node7368 : node7361;
													assign node7361 = (inp[4]) ? node7363 : 4'b1000;
														assign node7363 = (inp[10]) ? 4'b1100 : node7364;
															assign node7364 = (inp[12]) ? 4'b0100 : 4'b1100;
													assign node7368 = (inp[12]) ? node7370 : 4'b1000;
														assign node7370 = (inp[10]) ? 4'b1000 : 4'b0000;
												assign node7373 = (inp[7]) ? node7381 : node7374;
													assign node7374 = (inp[4]) ? 4'b1000 : node7375;
														assign node7375 = (inp[12]) ? node7377 : 4'b1100;
															assign node7377 = (inp[11]) ? 4'b0100 : 4'b1100;
													assign node7381 = (inp[12]) ? node7383 : 4'b1100;
														assign node7383 = (inp[10]) ? 4'b1100 : 4'b0100;
											assign node7386 = (inp[12]) ? node7398 : node7387;
												assign node7387 = (inp[3]) ? node7393 : node7388;
													assign node7388 = (inp[4]) ? 4'b0100 : node7389;
														assign node7389 = (inp[7]) ? 4'b0000 : 4'b0100;
													assign node7393 = (inp[7]) ? node7395 : 4'b0000;
														assign node7395 = (inp[4]) ? 4'b0000 : 4'b0100;
												assign node7398 = (inp[10]) ? node7402 : node7399;
													assign node7399 = (inp[3]) ? 4'b1100 : 4'b1000;
													assign node7402 = (inp[3]) ? node7408 : node7403;
														assign node7403 = (inp[4]) ? 4'b0100 : node7404;
															assign node7404 = (inp[7]) ? 4'b0000 : 4'b0100;
														assign node7408 = (inp[7]) ? node7410 : 4'b0000;
															assign node7410 = (inp[4]) ? 4'b0000 : 4'b0100;
										assign node7413 = (inp[11]) ? node7451 : node7414;
											assign node7414 = (inp[13]) ? node7438 : node7415;
												assign node7415 = (inp[12]) ? node7429 : node7416;
													assign node7416 = (inp[10]) ? node7424 : node7417;
														assign node7417 = (inp[4]) ? node7419 : 4'b0001;
															assign node7419 = (inp[7]) ? 4'b0101 : node7420;
																assign node7420 = (inp[3]) ? 4'b0001 : 4'b0101;
														assign node7424 = (inp[3]) ? node7426 : 4'b1001;
															assign node7426 = (inp[4]) ? 4'b1001 : 4'b1101;
													assign node7429 = (inp[7]) ? 4'b0101 : node7430;
														assign node7430 = (inp[4]) ? node7434 : node7431;
															assign node7431 = (inp[3]) ? 4'b0101 : 4'b0001;
															assign node7434 = (inp[3]) ? 4'b0001 : 4'b0101;
												assign node7438 = (inp[3]) ? node7446 : node7439;
													assign node7439 = (inp[10]) ? node7441 : 4'b1001;
														assign node7441 = (inp[4]) ? 4'b0101 : node7442;
															assign node7442 = (inp[12]) ? 4'b1001 : 4'b0001;
													assign node7446 = (inp[10]) ? node7448 : 4'b1101;
														assign node7448 = (inp[12]) ? 4'b1101 : 4'b0001;
											assign node7451 = (inp[13]) ? node7465 : node7452;
												assign node7452 = (inp[3]) ? node7460 : node7453;
													assign node7453 = (inp[12]) ? 4'b0100 : node7454;
														assign node7454 = (inp[7]) ? 4'b1000 : node7455;
															assign node7455 = (inp[4]) ? 4'b1100 : 4'b1000;
													assign node7460 = (inp[4]) ? node7462 : 4'b1100;
														assign node7462 = (inp[7]) ? 4'b1100 : 4'b1000;
												assign node7465 = (inp[7]) ? 4'b0100 : node7466;
													assign node7466 = (inp[10]) ? 4'b0000 : node7467;
														assign node7467 = (inp[4]) ? 4'b0100 : node7468;
															assign node7468 = (inp[3]) ? 4'b1100 : 4'b1000;
									assign node7474 = (inp[11]) ? node7544 : node7475;
										assign node7475 = (inp[14]) ? node7507 : node7476;
											assign node7476 = (inp[13]) ? node7486 : node7477;
												assign node7477 = (inp[10]) ? 4'b1101 : node7478;
													assign node7478 = (inp[12]) ? node7482 : node7479;
														assign node7479 = (inp[3]) ? 4'b1101 : 4'b1001;
														assign node7482 = (inp[3]) ? 4'b0101 : 4'b0001;
												assign node7486 = (inp[12]) ? node7496 : node7487;
													assign node7487 = (inp[3]) ? node7493 : node7488;
														assign node7488 = (inp[7]) ? node7490 : 4'b0101;
															assign node7490 = (inp[4]) ? 4'b0101 : 4'b0001;
														assign node7493 = (inp[4]) ? 4'b0001 : 4'b0101;
													assign node7496 = (inp[10]) ? node7500 : node7497;
														assign node7497 = (inp[7]) ? 4'b1001 : 4'b1101;
														assign node7500 = (inp[4]) ? 4'b0001 : node7501;
															assign node7501 = (inp[7]) ? node7503 : 4'b0101;
																assign node7503 = (inp[3]) ? 4'b0101 : 4'b0001;
											assign node7507 = (inp[13]) ? node7519 : node7508;
												assign node7508 = (inp[3]) ? node7510 : 4'b1000;
													assign node7510 = (inp[4]) ? node7516 : node7511;
														assign node7511 = (inp[10]) ? 4'b1100 : node7512;
															assign node7512 = (inp[12]) ? 4'b0100 : 4'b1100;
														assign node7516 = (inp[7]) ? 4'b1100 : 4'b1000;
												assign node7519 = (inp[12]) ? node7529 : node7520;
													assign node7520 = (inp[10]) ? 4'b0100 : node7521;
														assign node7521 = (inp[7]) ? node7523 : 4'b0000;
															assign node7523 = (inp[4]) ? 4'b0100 : node7524;
																assign node7524 = (inp[3]) ? 4'b0100 : 4'b0000;
													assign node7529 = (inp[10]) ? node7541 : node7530;
														assign node7530 = (inp[3]) ? node7536 : node7531;
															assign node7531 = (inp[4]) ? node7533 : 4'b1000;
																assign node7533 = (inp[7]) ? 4'b1000 : 4'b1100;
															assign node7536 = (inp[4]) ? node7538 : 4'b1100;
																assign node7538 = (inp[7]) ? 4'b1100 : 4'b1000;
														assign node7541 = (inp[3]) ? 4'b0000 : 4'b0100;
										assign node7544 = (inp[13]) ? node7580 : node7545;
											assign node7545 = (inp[12]) ? node7557 : node7546;
												assign node7546 = (inp[3]) ? node7552 : node7547;
													assign node7547 = (inp[7]) ? 4'b1001 : node7548;
														assign node7548 = (inp[4]) ? 4'b1101 : 4'b1001;
													assign node7552 = (inp[7]) ? 4'b1101 : node7553;
														assign node7553 = (inp[4]) ? 4'b1001 : 4'b1101;
												assign node7557 = (inp[10]) ? node7569 : node7558;
													assign node7558 = (inp[3]) ? node7564 : node7559;
														assign node7559 = (inp[4]) ? node7561 : 4'b0001;
															assign node7561 = (inp[7]) ? 4'b0001 : 4'b0101;
														assign node7564 = (inp[7]) ? 4'b0101 : node7565;
															assign node7565 = (inp[14]) ? 4'b0001 : 4'b0101;
													assign node7569 = (inp[14]) ? 4'b1001 : node7570;
														assign node7570 = (inp[3]) ? node7574 : node7571;
															assign node7571 = (inp[7]) ? 4'b1001 : 4'b1101;
															assign node7574 = (inp[4]) ? node7576 : 4'b1101;
																assign node7576 = (inp[7]) ? 4'b1101 : 4'b1001;
											assign node7580 = (inp[12]) ? node7588 : node7581;
												assign node7581 = (inp[3]) ? node7583 : 4'b0101;
													assign node7583 = (inp[4]) ? 4'b0001 : node7584;
														assign node7584 = (inp[7]) ? 4'b0101 : 4'b0001;
												assign node7588 = (inp[10]) ? node7602 : node7589;
													assign node7589 = (inp[14]) ? node7597 : node7590;
														assign node7590 = (inp[7]) ? 4'b1001 : node7591;
															assign node7591 = (inp[3]) ? node7593 : 4'b1101;
																assign node7593 = (inp[4]) ? 4'b1001 : 4'b1101;
														assign node7597 = (inp[7]) ? 4'b1101 : node7598;
															assign node7598 = (inp[4]) ? 4'b1001 : 4'b1101;
													assign node7602 = (inp[3]) ? node7606 : node7603;
														assign node7603 = (inp[4]) ? 4'b0101 : 4'b0001;
														assign node7606 = (inp[4]) ? 4'b0001 : node7607;
															assign node7607 = (inp[14]) ? 4'b0001 : 4'b0101;
								assign node7611 = (inp[3]) ? node7613 : 4'b0011;
									assign node7613 = (inp[7]) ? node7687 : node7614;
										assign node7614 = (inp[4]) ? node7642 : node7615;
											assign node7615 = (inp[13]) ? node7617 : 4'b0011;
												assign node7617 = (inp[12]) ? node7629 : node7618;
													assign node7618 = (inp[1]) ? node7624 : node7619;
														assign node7619 = (inp[14]) ? node7621 : 4'b0000;
															assign node7621 = (inp[11]) ? 4'b0000 : 4'b0001;
														assign node7624 = (inp[11]) ? 4'b0001 : node7625;
															assign node7625 = (inp[14]) ? 4'b0000 : 4'b0001;
													assign node7629 = (inp[10]) ? node7631 : 4'b0011;
														assign node7631 = (inp[1]) ? node7637 : node7632;
															assign node7632 = (inp[14]) ? node7634 : 4'b0000;
																assign node7634 = (inp[11]) ? 4'b0000 : 4'b0011;
															assign node7637 = (inp[11]) ? 4'b0001 : node7638;
																assign node7638 = (inp[14]) ? 4'b0000 : 4'b0001;
											assign node7642 = (inp[1]) ? node7662 : node7643;
												assign node7643 = (inp[14]) ? node7655 : node7644;
													assign node7644 = (inp[13]) ? node7650 : node7645;
														assign node7645 = (inp[10]) ? 4'b1000 : node7646;
															assign node7646 = (inp[12]) ? 4'b0000 : 4'b1000;
														assign node7650 = (inp[10]) ? 4'b0000 : node7651;
															assign node7651 = (inp[12]) ? 4'b1000 : 4'b0000;
													assign node7655 = (inp[11]) ? node7657 : 4'b0001;
														assign node7657 = (inp[13]) ? 4'b1000 : node7658;
															assign node7658 = (inp[12]) ? 4'b0000 : 4'b1000;
												assign node7662 = (inp[11]) ? node7676 : node7663;
													assign node7663 = (inp[14]) ? node7669 : node7664;
														assign node7664 = (inp[13]) ? node7666 : 4'b1001;
															assign node7666 = (inp[10]) ? 4'b0001 : 4'b1001;
														assign node7669 = (inp[12]) ? node7671 : 4'b1000;
															assign node7671 = (inp[10]) ? 4'b0000 : node7672;
																assign node7672 = (inp[13]) ? 4'b1000 : 4'b0000;
													assign node7676 = (inp[13]) ? node7682 : node7677;
														assign node7677 = (inp[12]) ? node7679 : 4'b1001;
															assign node7679 = (inp[10]) ? 4'b1001 : 4'b0001;
														assign node7682 = (inp[10]) ? 4'b0001 : node7683;
															assign node7683 = (inp[12]) ? 4'b1001 : 4'b0001;
										assign node7687 = (inp[4]) ? node7689 : 4'b0011;
											assign node7689 = (inp[13]) ? node7691 : 4'b0011;
												assign node7691 = (inp[12]) ? node7693 : 4'b0000;
													assign node7693 = (inp[10]) ? node7695 : 4'b0011;
														assign node7695 = (inp[1]) ? node7699 : node7696;
															assign node7696 = (inp[14]) ? 4'b0011 : 4'b0000;
															assign node7699 = (inp[14]) ? 4'b0000 : 4'b0001;
						assign node7702 = (inp[5]) ? node8258 : node7703;
							assign node7703 = (inp[1]) ? node8007 : node7704;
								assign node7704 = (inp[14]) ? node7846 : node7705;
									assign node7705 = (inp[13]) ? node7767 : node7706;
										assign node7706 = (inp[3]) ? node7732 : node7707;
											assign node7707 = (inp[4]) ? node7715 : node7708;
												assign node7708 = (inp[11]) ? 4'b1000 : node7709;
													assign node7709 = (inp[12]) ? node7711 : 4'b1000;
														assign node7711 = (inp[10]) ? 4'b1000 : 4'b0000;
												assign node7715 = (inp[7]) ? node7727 : node7716;
													assign node7716 = (inp[2]) ? node7722 : node7717;
														assign node7717 = (inp[10]) ? 4'b0000 : node7718;
															assign node7718 = (inp[12]) ? 4'b0100 : 4'b1100;
														assign node7722 = (inp[10]) ? 4'b1100 : node7723;
															assign node7723 = (inp[11]) ? 4'b1100 : 4'b0100;
													assign node7727 = (inp[12]) ? node7729 : 4'b1000;
														assign node7729 = (inp[10]) ? 4'b1000 : 4'b0000;
											assign node7732 = (inp[2]) ? node7758 : node7733;
												assign node7733 = (inp[11]) ? node7749 : node7734;
													assign node7734 = (inp[4]) ? node7744 : node7735;
														assign node7735 = (inp[7]) ? 4'b1000 : node7736;
															assign node7736 = (inp[12]) ? node7740 : node7737;
																assign node7737 = (inp[10]) ? 4'b0100 : 4'b1000;
																assign node7740 = (inp[10]) ? 4'b1000 : 4'b0000;
														assign node7744 = (inp[10]) ? node7746 : 4'b0100;
															assign node7746 = (inp[12]) ? 4'b1100 : 4'b0100;
													assign node7749 = (inp[4]) ? 4'b1101 : node7750;
														assign node7750 = (inp[10]) ? node7754 : node7751;
															assign node7751 = (inp[12]) ? 4'b0001 : 4'b1001;
															assign node7754 = (inp[7]) ? 4'b0001 : 4'b0101;
												assign node7758 = (inp[7]) ? node7762 : node7759;
													assign node7759 = (inp[4]) ? 4'b1000 : 4'b1100;
													assign node7762 = (inp[12]) ? node7764 : 4'b1100;
														assign node7764 = (inp[10]) ? 4'b1100 : 4'b0100;
										assign node7767 = (inp[12]) ? node7805 : node7768;
											assign node7768 = (inp[4]) ? node7788 : node7769;
												assign node7769 = (inp[2]) ? node7781 : node7770;
													assign node7770 = (inp[10]) ? node7774 : node7771;
														assign node7771 = (inp[7]) ? 4'b1000 : 4'b1100;
														assign node7774 = (inp[7]) ? 4'b0000 : node7775;
															assign node7775 = (inp[3]) ? node7777 : 4'b0100;
																assign node7777 = (inp[11]) ? 4'b0101 : 4'b0100;
													assign node7781 = (inp[3]) ? node7785 : node7782;
														assign node7782 = (inp[7]) ? 4'b0000 : 4'b0100;
														assign node7785 = (inp[7]) ? 4'b0100 : 4'b0000;
												assign node7788 = (inp[3]) ? node7796 : node7789;
													assign node7789 = (inp[2]) ? 4'b0100 : node7790;
														assign node7790 = (inp[11]) ? 4'b0001 : node7791;
															assign node7791 = (inp[10]) ? 4'b0000 : 4'b0100;
													assign node7796 = (inp[11]) ? node7800 : node7797;
														assign node7797 = (inp[7]) ? 4'b0000 : 4'b1001;
														assign node7800 = (inp[7]) ? 4'b1101 : node7801;
															assign node7801 = (inp[2]) ? 4'b1001 : 4'b0000;
											assign node7805 = (inp[2]) ? node7827 : node7806;
												assign node7806 = (inp[11]) ? node7812 : node7807;
													assign node7807 = (inp[3]) ? node7809 : 4'b1000;
														assign node7809 = (inp[4]) ? 4'b0000 : 4'b1000;
													assign node7812 = (inp[3]) ? node7820 : node7813;
														assign node7813 = (inp[7]) ? node7817 : node7814;
															assign node7814 = (inp[4]) ? 4'b0001 : 4'b0100;
															assign node7817 = (inp[10]) ? 4'b0000 : 4'b1000;
														assign node7820 = (inp[10]) ? node7824 : node7821;
															assign node7821 = (inp[4]) ? 4'b0101 : 4'b0001;
															assign node7824 = (inp[4]) ? 4'b1000 : 4'b1101;
												assign node7827 = (inp[10]) ? node7835 : node7828;
													assign node7828 = (inp[3]) ? 4'b1100 : node7829;
														assign node7829 = (inp[4]) ? node7831 : 4'b1000;
															assign node7831 = (inp[7]) ? 4'b1000 : 4'b1100;
													assign node7835 = (inp[3]) ? node7839 : node7836;
														assign node7836 = (inp[4]) ? 4'b0100 : 4'b0000;
														assign node7839 = (inp[7]) ? node7843 : node7840;
															assign node7840 = (inp[11]) ? 4'b1001 : 4'b1000;
															assign node7843 = (inp[4]) ? 4'b0000 : 4'b0100;
									assign node7846 = (inp[11]) ? node7928 : node7847;
										assign node7847 = (inp[3]) ? node7877 : node7848;
											assign node7848 = (inp[13]) ? node7860 : node7849;
												assign node7849 = (inp[10]) ? node7855 : node7850;
													assign node7850 = (inp[7]) ? 4'b0001 : node7851;
														assign node7851 = (inp[4]) ? 4'b0101 : 4'b0001;
													assign node7855 = (inp[12]) ? 4'b0001 : node7856;
														assign node7856 = (inp[4]) ? 4'b1101 : 4'b1001;
												assign node7860 = (inp[10]) ? node7868 : node7861;
													assign node7861 = (inp[4]) ? node7863 : 4'b1001;
														assign node7863 = (inp[12]) ? node7865 : 4'b1000;
															assign node7865 = (inp[7]) ? 4'b1001 : 4'b1101;
													assign node7868 = (inp[12]) ? 4'b1001 : node7869;
														assign node7869 = (inp[2]) ? node7873 : node7870;
															assign node7870 = (inp[4]) ? 4'b0000 : 4'b0101;
															assign node7873 = (inp[7]) ? 4'b0001 : 4'b0101;
											assign node7877 = (inp[2]) ? node7901 : node7878;
												assign node7878 = (inp[13]) ? node7890 : node7879;
													assign node7879 = (inp[4]) ? node7885 : node7880;
														assign node7880 = (inp[10]) ? 4'b1000 : node7881;
															assign node7881 = (inp[12]) ? 4'b0000 : 4'b1000;
														assign node7885 = (inp[12]) ? 4'b1100 : node7886;
															assign node7886 = (inp[10]) ? 4'b0000 : 4'b1100;
													assign node7890 = (inp[7]) ? node7894 : node7891;
														assign node7891 = (inp[4]) ? 4'b0000 : 4'b0100;
														assign node7894 = (inp[4]) ? node7898 : node7895;
															assign node7895 = (inp[10]) ? 4'b1000 : 4'b0000;
															assign node7898 = (inp[12]) ? 4'b0100 : 4'b1100;
												assign node7901 = (inp[4]) ? node7917 : node7902;
													assign node7902 = (inp[7]) ? node7910 : node7903;
														assign node7903 = (inp[10]) ? node7905 : 4'b1101;
															assign node7905 = (inp[13]) ? node7907 : 4'b1101;
																assign node7907 = (inp[12]) ? 4'b1101 : 4'b0001;
														assign node7910 = (inp[13]) ? node7912 : 4'b0101;
															assign node7912 = (inp[10]) ? node7914 : 4'b1101;
																assign node7914 = (inp[12]) ? 4'b1101 : 4'b0101;
													assign node7917 = (inp[7]) ? node7923 : node7918;
														assign node7918 = (inp[10]) ? 4'b0000 : node7919;
															assign node7919 = (inp[12]) ? 4'b0000 : 4'b0001;
														assign node7923 = (inp[13]) ? node7925 : 4'b0101;
															assign node7925 = (inp[10]) ? 4'b0000 : 4'b1101;
										assign node7928 = (inp[3]) ? node7962 : node7929;
											assign node7929 = (inp[13]) ? node7943 : node7930;
												assign node7930 = (inp[10]) ? node7938 : node7931;
													assign node7931 = (inp[12]) ? node7935 : node7932;
														assign node7932 = (inp[4]) ? 4'b1100 : 4'b1000;
														assign node7935 = (inp[7]) ? 4'b0000 : 4'b0100;
													assign node7938 = (inp[7]) ? 4'b1000 : node7939;
														assign node7939 = (inp[4]) ? 4'b1100 : 4'b1000;
												assign node7943 = (inp[10]) ? node7957 : node7944;
													assign node7944 = (inp[12]) ? node7952 : node7945;
														assign node7945 = (inp[2]) ? node7949 : node7946;
															assign node7946 = (inp[4]) ? 4'b1001 : 4'b0100;
															assign node7949 = (inp[4]) ? 4'b0100 : 4'b0000;
														assign node7952 = (inp[4]) ? node7954 : 4'b1000;
															assign node7954 = (inp[7]) ? 4'b1000 : 4'b1100;
													assign node7957 = (inp[7]) ? 4'b0100 : node7958;
														assign node7958 = (inp[4]) ? 4'b0001 : 4'b0100;
											assign node7962 = (inp[2]) ? node7988 : node7963;
												assign node7963 = (inp[4]) ? node7977 : node7964;
													assign node7964 = (inp[12]) ? node7974 : node7965;
														assign node7965 = (inp[10]) ? node7969 : node7966;
															assign node7966 = (inp[13]) ? 4'b1101 : 4'b1001;
															assign node7969 = (inp[7]) ? node7971 : 4'b0101;
																assign node7971 = (inp[13]) ? 4'b0101 : 4'b0001;
														assign node7974 = (inp[10]) ? 4'b1001 : 4'b0001;
													assign node7977 = (inp[10]) ? node7985 : node7978;
														assign node7978 = (inp[7]) ? node7982 : node7979;
															assign node7979 = (inp[13]) ? 4'b0000 : 4'b1101;
															assign node7982 = (inp[12]) ? 4'b0101 : 4'b1101;
														assign node7985 = (inp[12]) ? 4'b1000 : 4'b0000;
												assign node7988 = (inp[4]) ? node7996 : node7989;
													assign node7989 = (inp[13]) ? node7991 : 4'b1100;
														assign node7991 = (inp[7]) ? node7993 : 4'b0000;
															assign node7993 = (inp[12]) ? 4'b1100 : 4'b0100;
													assign node7996 = (inp[13]) ? node8002 : node7997;
														assign node7997 = (inp[7]) ? 4'b1100 : node7998;
															assign node7998 = (inp[10]) ? 4'b0001 : 4'b0000;
														assign node8002 = (inp[10]) ? node8004 : 4'b0001;
															assign node8004 = (inp[12]) ? 4'b1001 : 4'b0001;
								assign node8007 = (inp[11]) ? node8159 : node8008;
									assign node8008 = (inp[14]) ? node8094 : node8009;
										assign node8009 = (inp[3]) ? node8055 : node8010;
											assign node8010 = (inp[7]) ? node8040 : node8011;
												assign node8011 = (inp[2]) ? node8021 : node8012;
													assign node8012 = (inp[4]) ? node8014 : 4'b0101;
														assign node8014 = (inp[12]) ? node8018 : node8015;
															assign node8015 = (inp[13]) ? 4'b1000 : 4'b0000;
															assign node8018 = (inp[13]) ? 4'b0000 : 4'b0101;
													assign node8021 = (inp[4]) ? node8031 : node8022;
														assign node8022 = (inp[10]) ? node8028 : node8023;
															assign node8023 = (inp[13]) ? 4'b1001 : node8024;
																assign node8024 = (inp[12]) ? 4'b0001 : 4'b1001;
															assign node8028 = (inp[13]) ? 4'b0101 : 4'b1001;
														assign node8031 = (inp[12]) ? node8035 : node8032;
															assign node8032 = (inp[10]) ? 4'b1101 : 4'b0101;
															assign node8035 = (inp[10]) ? 4'b0101 : node8036;
																assign node8036 = (inp[13]) ? 4'b1101 : 4'b0101;
												assign node8040 = (inp[13]) ? node8046 : node8041;
													assign node8041 = (inp[10]) ? 4'b1001 : node8042;
														assign node8042 = (inp[12]) ? 4'b0001 : 4'b1001;
													assign node8046 = (inp[12]) ? node8052 : node8047;
														assign node8047 = (inp[10]) ? node8049 : 4'b0101;
															assign node8049 = (inp[2]) ? 4'b0101 : 4'b0000;
														assign node8052 = (inp[10]) ? 4'b0001 : 4'b1001;
											assign node8055 = (inp[10]) ? node8077 : node8056;
												assign node8056 = (inp[2]) ? node8066 : node8057;
													assign node8057 = (inp[4]) ? node8063 : node8058;
														assign node8058 = (inp[7]) ? 4'b1000 : node8059;
															assign node8059 = (inp[13]) ? 4'b1100 : 4'b1000;
														assign node8063 = (inp[7]) ? 4'b1100 : 4'b1000;
													assign node8066 = (inp[4]) ? node8074 : node8067;
														assign node8067 = (inp[13]) ? node8071 : node8068;
															assign node8068 = (inp[12]) ? 4'b0101 : 4'b1101;
															assign node8071 = (inp[12]) ? 4'b1101 : 4'b0101;
														assign node8074 = (inp[7]) ? 4'b1101 : 4'b1000;
												assign node8077 = (inp[4]) ? node8089 : node8078;
													assign node8078 = (inp[2]) ? node8084 : node8079;
														assign node8079 = (inp[7]) ? node8081 : 4'b0100;
															assign node8081 = (inp[13]) ? 4'b0100 : 4'b0000;
														assign node8084 = (inp[12]) ? 4'b1101 : node8085;
															assign node8085 = (inp[7]) ? 4'b0101 : 4'b0001;
													assign node8089 = (inp[7]) ? node8091 : 4'b0000;
														assign node8091 = (inp[13]) ? 4'b0000 : 4'b0100;
										assign node8094 = (inp[13]) ? node8128 : node8095;
											assign node8095 = (inp[3]) ? node8107 : node8096;
												assign node8096 = (inp[10]) ? 4'b1000 : node8097;
													assign node8097 = (inp[12]) ? node8103 : node8098;
														assign node8098 = (inp[7]) ? 4'b1000 : node8099;
															assign node8099 = (inp[4]) ? 4'b1100 : 4'b1000;
														assign node8103 = (inp[7]) ? 4'b0000 : 4'b0100;
												assign node8107 = (inp[10]) ? node8119 : node8108;
													assign node8108 = (inp[2]) ? node8112 : node8109;
														assign node8109 = (inp[4]) ? 4'b1100 : 4'b1000;
														assign node8112 = (inp[12]) ? 4'b0100 : node8113;
															assign node8113 = (inp[7]) ? 4'b1100 : node8114;
																assign node8114 = (inp[4]) ? 4'b1000 : 4'b1100;
													assign node8119 = (inp[2]) ? node8123 : node8120;
														assign node8120 = (inp[4]) ? 4'b0100 : 4'b0000;
														assign node8123 = (inp[12]) ? 4'b1100 : node8124;
															assign node8124 = (inp[7]) ? 4'b1100 : 4'b0000;
											assign node8128 = (inp[10]) ? node8142 : node8129;
												assign node8129 = (inp[4]) ? 4'b0001 : node8130;
													assign node8130 = (inp[12]) ? node8138 : node8131;
														assign node8131 = (inp[2]) ? node8133 : 4'b1000;
															assign node8133 = (inp[3]) ? node8135 : 4'b0000;
																assign node8135 = (inp[7]) ? 4'b0100 : 4'b0000;
														assign node8138 = (inp[3]) ? 4'b1100 : 4'b1000;
												assign node8142 = (inp[4]) ? node8148 : node8143;
													assign node8143 = (inp[7]) ? node8145 : 4'b0100;
														assign node8145 = (inp[3]) ? 4'b0100 : 4'b0000;
													assign node8148 = (inp[3]) ? node8152 : node8149;
														assign node8149 = (inp[2]) ? 4'b0100 : 4'b0000;
														assign node8152 = (inp[2]) ? 4'b0000 : node8153;
															assign node8153 = (inp[7]) ? 4'b0000 : node8154;
																assign node8154 = (inp[12]) ? 4'b1001 : 4'b0001;
									assign node8159 = (inp[13]) ? node8201 : node8160;
										assign node8160 = (inp[3]) ? node8176 : node8161;
											assign node8161 = (inp[10]) ? node8169 : node8162;
												assign node8162 = (inp[4]) ? node8166 : node8163;
													assign node8163 = (inp[12]) ? 4'b0001 : 4'b1001;
													assign node8166 = (inp[12]) ? 4'b0101 : 4'b1101;
												assign node8169 = (inp[7]) ? 4'b1001 : node8170;
													assign node8170 = (inp[4]) ? node8172 : 4'b1001;
														assign node8172 = (inp[12]) ? 4'b1101 : 4'b0001;
											assign node8176 = (inp[10]) ? node8188 : node8177;
												assign node8177 = (inp[2]) ? node8181 : node8178;
													assign node8178 = (inp[4]) ? 4'b1101 : 4'b1001;
													assign node8181 = (inp[12]) ? 4'b0101 : node8182;
														assign node8182 = (inp[7]) ? 4'b1101 : node8183;
															assign node8183 = (inp[4]) ? 4'b1001 : 4'b1101;
												assign node8188 = (inp[2]) ? node8196 : node8189;
													assign node8189 = (inp[7]) ? node8193 : node8190;
														assign node8190 = (inp[4]) ? 4'b0001 : 4'b0101;
														assign node8193 = (inp[4]) ? 4'b0101 : 4'b0001;
													assign node8196 = (inp[4]) ? node8198 : 4'b1101;
														assign node8198 = (inp[7]) ? 4'b1101 : 4'b0001;
										assign node8201 = (inp[10]) ? node8235 : node8202;
											assign node8202 = (inp[12]) ? node8224 : node8203;
												assign node8203 = (inp[3]) ? node8213 : node8204;
													assign node8204 = (inp[7]) ? node8210 : node8205;
														assign node8205 = (inp[4]) ? node8207 : 4'b0101;
															assign node8207 = (inp[2]) ? 4'b0101 : 4'b1001;
														assign node8210 = (inp[4]) ? 4'b0101 : 4'b0001;
													assign node8213 = (inp[2]) ? node8221 : node8214;
														assign node8214 = (inp[14]) ? node8216 : 4'b1101;
															assign node8216 = (inp[7]) ? 4'b1001 : node8217;
																assign node8217 = (inp[4]) ? 4'b1001 : 4'b1101;
														assign node8221 = (inp[14]) ? 4'b0001 : 4'b0101;
												assign node8224 = (inp[4]) ? node8226 : 4'b1001;
													assign node8226 = (inp[3]) ? node8230 : node8227;
														assign node8227 = (inp[7]) ? 4'b1001 : 4'b1101;
														assign node8230 = (inp[7]) ? 4'b1101 : node8231;
															assign node8231 = (inp[2]) ? 4'b1001 : 4'b0001;
											assign node8235 = (inp[4]) ? node8253 : node8236;
												assign node8236 = (inp[14]) ? 4'b0101 : node8237;
													assign node8237 = (inp[2]) ? node8239 : 4'b0101;
														assign node8239 = (inp[12]) ? node8245 : node8240;
															assign node8240 = (inp[3]) ? node8242 : 4'b0001;
																assign node8242 = (inp[7]) ? 4'b0101 : 4'b0001;
															assign node8245 = (inp[3]) ? node8249 : node8246;
																assign node8246 = (inp[7]) ? 4'b0001 : 4'b0101;
																assign node8249 = (inp[7]) ? 4'b0101 : 4'b0001;
												assign node8253 = (inp[3]) ? 4'b0001 : node8254;
													assign node8254 = (inp[2]) ? 4'b0101 : 4'b0001;
							assign node8258 = (inp[3]) ? node8566 : node8259;
								assign node8259 = (inp[11]) ? node8413 : node8260;
									assign node8260 = (inp[2]) ? node8340 : node8261;
										assign node8261 = (inp[4]) ? node8299 : node8262;
											assign node8262 = (inp[13]) ? node8278 : node8263;
												assign node8263 = (inp[1]) ? node8269 : node8264;
													assign node8264 = (inp[7]) ? 4'b0000 : node8265;
														assign node8265 = (inp[12]) ? 4'b0000 : 4'b1000;
													assign node8269 = (inp[14]) ? node8275 : node8270;
														assign node8270 = (inp[12]) ? 4'b1000 : node8271;
															assign node8271 = (inp[10]) ? 4'b1100 : 4'b0100;
														assign node8275 = (inp[10]) ? 4'b1101 : 4'b1001;
												assign node8278 = (inp[10]) ? node8288 : node8279;
													assign node8279 = (inp[7]) ? node8285 : node8280;
														assign node8280 = (inp[1]) ? node8282 : 4'b0101;
															assign node8282 = (inp[12]) ? 4'b0101 : 4'b0001;
														assign node8285 = (inp[1]) ? 4'b1100 : 4'b0101;
													assign node8288 = (inp[1]) ? node8294 : node8289;
														assign node8289 = (inp[7]) ? node8291 : 4'b1001;
															assign node8291 = (inp[14]) ? 4'b1100 : 4'b1101;
														assign node8294 = (inp[12]) ? node8296 : 4'b0001;
															assign node8296 = (inp[7]) ? 4'b1101 : 4'b1001;
											assign node8299 = (inp[10]) ? node8313 : node8300;
												assign node8300 = (inp[1]) ? node8306 : node8301;
													assign node8301 = (inp[12]) ? node8303 : 4'b0001;
														assign node8303 = (inp[13]) ? 4'b1001 : 4'b0001;
													assign node8306 = (inp[13]) ? node8310 : node8307;
														assign node8307 = (inp[12]) ? 4'b1001 : 4'b0001;
														assign node8310 = (inp[14]) ? 4'b1000 : 4'b1001;
												assign node8313 = (inp[13]) ? node8329 : node8314;
													assign node8314 = (inp[14]) ? node8324 : node8315;
														assign node8315 = (inp[1]) ? node8317 : 4'b1001;
															assign node8317 = (inp[12]) ? node8321 : node8318;
																assign node8318 = (inp[7]) ? 4'b0101 : 4'b1001;
																assign node8321 = (inp[7]) ? 4'b1001 : 4'b0001;
														assign node8324 = (inp[1]) ? node8326 : 4'b0101;
															assign node8326 = (inp[12]) ? 4'b0000 : 4'b1000;
													assign node8329 = (inp[7]) ? node8331 : 4'b0000;
														assign node8331 = (inp[1]) ? node8335 : node8332;
															assign node8332 = (inp[14]) ? 4'b0001 : 4'b1000;
															assign node8335 = (inp[12]) ? node8337 : 4'b0000;
																assign node8337 = (inp[14]) ? 4'b1000 : 4'b1001;
										assign node8340 = (inp[4]) ? node8370 : node8341;
											assign node8341 = (inp[10]) ? node8355 : node8342;
												assign node8342 = (inp[7]) ? node8350 : node8343;
													assign node8343 = (inp[13]) ? node8345 : 4'b1000;
														assign node8345 = (inp[12]) ? node8347 : 4'b1100;
															assign node8347 = (inp[14]) ? 4'b0100 : 4'b1100;
													assign node8350 = (inp[12]) ? node8352 : 4'b1000;
														assign node8352 = (inp[1]) ? 4'b1000 : 4'b0000;
												assign node8355 = (inp[13]) ? node8361 : node8356;
													assign node8356 = (inp[1]) ? node8358 : 4'b1000;
														assign node8358 = (inp[7]) ? 4'b0000 : 4'b0100;
													assign node8361 = (inp[7]) ? 4'b0100 : node8362;
														assign node8362 = (inp[14]) ? node8364 : 4'b0000;
															assign node8364 = (inp[1]) ? node8366 : 4'b0100;
																assign node8366 = (inp[12]) ? 4'b0100 : 4'b0001;
											assign node8370 = (inp[7]) ? node8392 : node8371;
												assign node8371 = (inp[13]) ? node8383 : node8372;
													assign node8372 = (inp[1]) ? node8378 : node8373;
														assign node8373 = (inp[14]) ? 4'b0000 : node8374;
															assign node8374 = (inp[12]) ? 4'b0001 : 4'b1001;
														assign node8378 = (inp[14]) ? 4'b1001 : node8379;
															assign node8379 = (inp[12]) ? 4'b1000 : 4'b0000;
													assign node8383 = (inp[12]) ? node8385 : 4'b0001;
														assign node8385 = (inp[10]) ? 4'b1001 : node8386;
															assign node8386 = (inp[1]) ? 4'b0100 : node8387;
																assign node8387 = (inp[14]) ? 4'b1000 : 4'b1001;
												assign node8392 = (inp[1]) ? node8402 : node8393;
													assign node8393 = (inp[13]) ? node8399 : node8394;
														assign node8394 = (inp[10]) ? node8396 : 4'b0100;
															assign node8396 = (inp[12]) ? 4'b0000 : 4'b0001;
														assign node8399 = (inp[10]) ? 4'b1001 : 4'b0001;
													assign node8402 = (inp[13]) ? 4'b0100 : node8403;
														assign node8403 = (inp[10]) ? node8409 : node8404;
															assign node8404 = (inp[14]) ? 4'b1100 : node8405;
																assign node8405 = (inp[12]) ? 4'b1100 : 4'b0000;
															assign node8409 = (inp[14]) ? 4'b1001 : 4'b1000;
									assign node8413 = (inp[1]) ? node8503 : node8414;
										assign node8414 = (inp[13]) ? node8468 : node8415;
											assign node8415 = (inp[12]) ? node8441 : node8416;
												assign node8416 = (inp[10]) ? node8432 : node8417;
													assign node8417 = (inp[7]) ? node8425 : node8418;
														assign node8418 = (inp[2]) ? node8422 : node8419;
															assign node8419 = (inp[4]) ? 4'b1001 : 4'b1000;
															assign node8422 = (inp[4]) ? 4'b1000 : 4'b1001;
														assign node8425 = (inp[2]) ? node8429 : node8426;
															assign node8426 = (inp[4]) ? 4'b1001 : 4'b1000;
															assign node8429 = (inp[4]) ? 4'b1101 : 4'b1001;
													assign node8432 = (inp[14]) ? node8438 : node8433;
														assign node8433 = (inp[7]) ? 4'b1000 : node8434;
															assign node8434 = (inp[4]) ? 4'b1000 : 4'b1100;
														assign node8438 = (inp[7]) ? 4'b1001 : 4'b1000;
												assign node8441 = (inp[7]) ? node8455 : node8442;
													assign node8442 = (inp[10]) ? node8450 : node8443;
														assign node8443 = (inp[2]) ? node8447 : node8444;
															assign node8444 = (inp[4]) ? 4'b1001 : 4'b1000;
															assign node8447 = (inp[4]) ? 4'b1000 : 4'b0001;
														assign node8450 = (inp[2]) ? node8452 : 4'b0100;
															assign node8452 = (inp[4]) ? 4'b0000 : 4'b1001;
													assign node8455 = (inp[14]) ? node8459 : node8456;
														assign node8456 = (inp[10]) ? 4'b1001 : 4'b1000;
														assign node8459 = (inp[2]) ? node8463 : node8460;
															assign node8460 = (inp[10]) ? 4'b0000 : 4'b1001;
															assign node8463 = (inp[10]) ? 4'b1001 : node8464;
																assign node8464 = (inp[4]) ? 4'b0101 : 4'b0001;
											assign node8468 = (inp[10]) ? node8484 : node8469;
												assign node8469 = (inp[2]) ? node8473 : node8470;
													assign node8470 = (inp[4]) ? 4'b0000 : 4'b0100;
													assign node8473 = (inp[4]) ? node8481 : node8474;
														assign node8474 = (inp[7]) ? node8478 : node8475;
															assign node8475 = (inp[12]) ? 4'b0101 : 4'b1101;
															assign node8478 = (inp[12]) ? 4'b0001 : 4'b1001;
														assign node8481 = (inp[7]) ? 4'b0000 : 4'b0100;
												assign node8484 = (inp[7]) ? node8496 : node8485;
													assign node8485 = (inp[2]) ? node8491 : node8486;
														assign node8486 = (inp[12]) ? node8488 : 4'b1001;
															assign node8488 = (inp[4]) ? 4'b0001 : 4'b1001;
														assign node8491 = (inp[12]) ? 4'b1101 : node8492;
															assign node8492 = (inp[14]) ? 4'b1001 : 4'b0000;
													assign node8496 = (inp[12]) ? node8500 : node8497;
														assign node8497 = (inp[2]) ? 4'b0101 : 4'b0100;
														assign node8500 = (inp[2]) ? 4'b1001 : 4'b1000;
										assign node8503 = (inp[13]) ? node8537 : node8504;
											assign node8504 = (inp[7]) ? node8522 : node8505;
												assign node8505 = (inp[12]) ? node8515 : node8506;
													assign node8506 = (inp[4]) ? node8512 : node8507;
														assign node8507 = (inp[10]) ? 4'b0101 : node8508;
															assign node8508 = (inp[2]) ? 4'b1001 : 4'b0101;
														assign node8512 = (inp[10]) ? 4'b1001 : 4'b0101;
													assign node8515 = (inp[2]) ? 4'b1001 : node8516;
														assign node8516 = (inp[10]) ? 4'b1001 : node8517;
															assign node8517 = (inp[4]) ? 4'b0101 : 4'b1001;
												assign node8522 = (inp[2]) ? node8528 : node8523;
													assign node8523 = (inp[10]) ? 4'b0101 : node8524;
														assign node8524 = (inp[4]) ? 4'b0001 : 4'b1001;
													assign node8528 = (inp[10]) ? node8534 : node8529;
														assign node8529 = (inp[4]) ? node8531 : 4'b1001;
															assign node8531 = (inp[12]) ? 4'b1101 : 4'b0001;
														assign node8534 = (inp[4]) ? 4'b1001 : 4'b0001;
											assign node8537 = (inp[10]) ? node8557 : node8538;
												assign node8538 = (inp[7]) ? node8544 : node8539;
													assign node8539 = (inp[4]) ? node8541 : 4'b1101;
														assign node8541 = (inp[2]) ? 4'b0001 : 4'b0101;
													assign node8544 = (inp[14]) ? node8550 : node8545;
														assign node8545 = (inp[12]) ? 4'b0101 : node8546;
															assign node8546 = (inp[2]) ? 4'b1001 : 4'b0001;
														assign node8550 = (inp[4]) ? node8552 : 4'b1001;
															assign node8552 = (inp[12]) ? node8554 : 4'b1001;
																assign node8554 = (inp[2]) ? 4'b0001 : 4'b1001;
												assign node8557 = (inp[14]) ? node8559 : 4'b0001;
													assign node8559 = (inp[7]) ? node8561 : 4'b0001;
														assign node8561 = (inp[2]) ? node8563 : 4'b0001;
															assign node8563 = (inp[4]) ? 4'b0001 : 4'b0101;
								assign node8566 = (inp[4]) ? node8716 : node8567;
									assign node8567 = (inp[11]) ? node8653 : node8568;
										assign node8568 = (inp[2]) ? node8624 : node8569;
											assign node8569 = (inp[12]) ? node8597 : node8570;
												assign node8570 = (inp[10]) ? node8586 : node8571;
													assign node8571 = (inp[13]) ? node8577 : node8572;
														assign node8572 = (inp[14]) ? node8574 : 4'b1000;
															assign node8574 = (inp[1]) ? 4'b1001 : 4'b1000;
														assign node8577 = (inp[1]) ? node8583 : node8578;
															assign node8578 = (inp[14]) ? 4'b0001 : node8579;
																assign node8579 = (inp[7]) ? 4'b1001 : 4'b1000;
															assign node8583 = (inp[7]) ? 4'b1000 : 4'b0000;
													assign node8586 = (inp[1]) ? node8592 : node8587;
														assign node8587 = (inp[14]) ? 4'b1000 : node8588;
															assign node8588 = (inp[13]) ? 4'b1000 : 4'b1001;
														assign node8592 = (inp[7]) ? node8594 : 4'b1001;
															assign node8594 = (inp[13]) ? 4'b1001 : 4'b0001;
												assign node8597 = (inp[10]) ? node8607 : node8598;
													assign node8598 = (inp[1]) ? 4'b0000 : node8599;
														assign node8599 = (inp[13]) ? node8601 : 4'b1000;
															assign node8601 = (inp[7]) ? 4'b1001 : node8602;
																assign node8602 = (inp[14]) ? 4'b0001 : 4'b0000;
													assign node8607 = (inp[1]) ? node8615 : node8608;
														assign node8608 = (inp[14]) ? 4'b0000 : node8609;
															assign node8609 = (inp[13]) ? node8611 : 4'b0001;
																assign node8611 = (inp[7]) ? 4'b0000 : 4'b0001;
														assign node8615 = (inp[14]) ? node8619 : node8616;
															assign node8616 = (inp[13]) ? 4'b1000 : 4'b0000;
															assign node8619 = (inp[7]) ? 4'b0001 : node8620;
																assign node8620 = (inp[13]) ? 4'b0001 : 4'b1001;
											assign node8624 = (inp[12]) ? node8640 : node8625;
												assign node8625 = (inp[1]) ? node8631 : node8626;
													assign node8626 = (inp[14]) ? 4'b0000 : node8627;
														assign node8627 = (inp[13]) ? 4'b0001 : 4'b0000;
													assign node8631 = (inp[14]) ? 4'b0001 : node8632;
														assign node8632 = (inp[10]) ? node8634 : 4'b1000;
															assign node8634 = (inp[13]) ? 4'b0000 : node8635;
																assign node8635 = (inp[7]) ? 4'b1001 : 4'b0000;
												assign node8640 = (inp[10]) ? node8650 : node8641;
													assign node8641 = (inp[13]) ? node8645 : node8642;
														assign node8642 = (inp[14]) ? 4'b1001 : 4'b0001;
														assign node8645 = (inp[7]) ? 4'b0000 : node8646;
															assign node8646 = (inp[1]) ? 4'b0000 : 4'b1000;
													assign node8650 = (inp[13]) ? 4'b1001 : 4'b1000;
										assign node8653 = (inp[1]) ? node8689 : node8654;
											assign node8654 = (inp[12]) ? node8668 : node8655;
												assign node8655 = (inp[2]) ? node8661 : node8656;
													assign node8656 = (inp[14]) ? node8658 : 4'b0000;
														assign node8658 = (inp[13]) ? 4'b0000 : 4'b0001;
													assign node8661 = (inp[13]) ? 4'b0001 : node8662;
														assign node8662 = (inp[10]) ? 4'b0000 : node8663;
															assign node8663 = (inp[7]) ? 4'b1001 : 4'b0000;
												assign node8668 = (inp[10]) ? node8678 : node8669;
													assign node8669 = (inp[2]) ? 4'b1001 : node8670;
														assign node8670 = (inp[7]) ? node8674 : node8671;
															assign node8671 = (inp[13]) ? 4'b1000 : 4'b0000;
															assign node8674 = (inp[13]) ? 4'b0001 : 4'b1001;
													assign node8678 = (inp[2]) ? node8684 : node8679;
														assign node8679 = (inp[13]) ? node8681 : 4'b0001;
															assign node8681 = (inp[7]) ? 4'b1001 : 4'b1000;
														assign node8684 = (inp[7]) ? 4'b0000 : node8685;
															assign node8685 = (inp[14]) ? 4'b0001 : 4'b0000;
											assign node8689 = (inp[10]) ? node8709 : node8690;
												assign node8690 = (inp[14]) ? node8700 : node8691;
													assign node8691 = (inp[12]) ? node8695 : node8692;
														assign node8692 = (inp[2]) ? 4'b1001 : 4'b0001;
														assign node8695 = (inp[2]) ? node8697 : 4'b1001;
															assign node8697 = (inp[13]) ? 4'b1001 : 4'b0001;
													assign node8700 = (inp[13]) ? node8706 : node8701;
														assign node8701 = (inp[12]) ? node8703 : 4'b0001;
															assign node8703 = (inp[2]) ? 4'b0001 : 4'b1001;
														assign node8706 = (inp[12]) ? 4'b0001 : 4'b1001;
												assign node8709 = (inp[7]) ? node8711 : 4'b0001;
													assign node8711 = (inp[2]) ? node8713 : 4'b0001;
														assign node8713 = (inp[13]) ? 4'b0001 : 4'b1001;
									assign node8716 = (inp[13]) ? node8802 : node8717;
										assign node8717 = (inp[1]) ? node8769 : node8718;
											assign node8718 = (inp[7]) ? node8742 : node8719;
												assign node8719 = (inp[2]) ? node8727 : node8720;
													assign node8720 = (inp[10]) ? node8722 : 4'b0000;
														assign node8722 = (inp[14]) ? 4'b0000 : node8723;
															assign node8723 = (inp[11]) ? 4'b0000 : 4'b0001;
													assign node8727 = (inp[14]) ? node8733 : node8728;
														assign node8728 = (inp[11]) ? node8730 : 4'b1000;
															assign node8730 = (inp[12]) ? 4'b0001 : 4'b0000;
														assign node8733 = (inp[12]) ? node8737 : node8734;
															assign node8734 = (inp[10]) ? 4'b0001 : 4'b0000;
															assign node8737 = (inp[10]) ? 4'b0001 : node8738;
																assign node8738 = (inp[11]) ? 4'b0001 : 4'b1001;
												assign node8742 = (inp[11]) ? node8758 : node8743;
													assign node8743 = (inp[12]) ? node8751 : node8744;
														assign node8744 = (inp[14]) ? node8746 : 4'b0000;
															assign node8746 = (inp[2]) ? 4'b0001 : node8747;
																assign node8747 = (inp[10]) ? 4'b0000 : 4'b0001;
														assign node8751 = (inp[14]) ? node8755 : node8752;
															assign node8752 = (inp[2]) ? 4'b1001 : 4'b1000;
															assign node8755 = (inp[2]) ? 4'b1000 : 4'b0001;
													assign node8758 = (inp[2]) ? node8764 : node8759;
														assign node8759 = (inp[10]) ? 4'b1000 : node8760;
															assign node8760 = (inp[12]) ? 4'b1000 : 4'b0001;
														assign node8764 = (inp[12]) ? 4'b0000 : node8765;
															assign node8765 = (inp[10]) ? 4'b0000 : 4'b1000;
											assign node8769 = (inp[11]) ? node8785 : node8770;
												assign node8770 = (inp[7]) ? node8776 : node8771;
													assign node8771 = (inp[2]) ? 4'b0001 : node8772;
														assign node8772 = (inp[14]) ? 4'b0001 : 4'b0000;
													assign node8776 = (inp[2]) ? node8780 : node8777;
														assign node8777 = (inp[10]) ? 4'b0000 : 4'b0001;
														assign node8780 = (inp[12]) ? 4'b0000 : node8781;
															assign node8781 = (inp[14]) ? 4'b1000 : 4'b0000;
												assign node8785 = (inp[10]) ? 4'b0001 : node8786;
													assign node8786 = (inp[14]) ? node8794 : node8787;
														assign node8787 = (inp[12]) ? node8789 : 4'b0001;
															assign node8789 = (inp[7]) ? node8791 : 4'b0001;
																assign node8791 = (inp[2]) ? 4'b1001 : 4'b0001;
														assign node8794 = (inp[7]) ? node8796 : 4'b1001;
															assign node8796 = (inp[12]) ? node8798 : 4'b0001;
																assign node8798 = (inp[2]) ? 4'b1001 : 4'b0001;
										assign node8802 = (inp[10]) ? node8832 : node8803;
											assign node8803 = (inp[11]) ? node8819 : node8804;
												assign node8804 = (inp[7]) ? node8812 : node8805;
													assign node8805 = (inp[12]) ? node8807 : 4'b0000;
														assign node8807 = (inp[1]) ? node8809 : 4'b0000;
															assign node8809 = (inp[14]) ? 4'b0000 : 4'b0001;
													assign node8812 = (inp[12]) ? 4'b0000 : node8813;
														assign node8813 = (inp[14]) ? node8815 : 4'b0001;
															assign node8815 = (inp[2]) ? 4'b0000 : 4'b0001;
												assign node8819 = (inp[1]) ? 4'b0001 : node8820;
													assign node8820 = (inp[12]) ? node8826 : node8821;
														assign node8821 = (inp[2]) ? node8823 : 4'b0000;
															assign node8823 = (inp[7]) ? 4'b0001 : 4'b0000;
														assign node8826 = (inp[2]) ? node8828 : 4'b0001;
															assign node8828 = (inp[7]) ? 4'b0000 : 4'b0001;
											assign node8832 = (inp[11]) ? 4'b0000 : node8833;
												assign node8833 = (inp[1]) ? 4'b0000 : node8834;
													assign node8834 = (inp[14]) ? node8842 : node8835;
														assign node8835 = (inp[12]) ? node8839 : node8836;
															assign node8836 = (inp[7]) ? 4'b0000 : 4'b0001;
															assign node8839 = (inp[7]) ? 4'b0001 : 4'b0000;
														assign node8842 = (inp[12]) ? node8846 : node8843;
															assign node8843 = (inp[7]) ? 4'b0001 : 4'b0000;
															assign node8846 = (inp[7]) ? 4'b0000 : 4'b0001;
					assign node8851 = (inp[6]) ? node8853 : 4'b0001;
						assign node8853 = (inp[5]) ? node8927 : node8854;
							assign node8854 = (inp[3]) ? node8856 : 4'b0001;
								assign node8856 = (inp[2]) ? 4'b0001 : node8857;
									assign node8857 = (inp[7]) ? node8909 : node8858;
										assign node8858 = (inp[4]) ? node8876 : node8859;
											assign node8859 = (inp[13]) ? node8861 : 4'b0001;
												assign node8861 = (inp[14]) ? node8867 : node8862;
													assign node8862 = (inp[1]) ? 4'b0001 : node8863;
														assign node8863 = (inp[10]) ? 4'b0000 : 4'b0001;
													assign node8867 = (inp[11]) ? 4'b0000 : node8868;
														assign node8868 = (inp[1]) ? node8870 : 4'b0001;
															assign node8870 = (inp[10]) ? 4'b0000 : node8871;
																assign node8871 = (inp[12]) ? 4'b0001 : 4'b0000;
											assign node8876 = (inp[1]) ? node8896 : node8877;
												assign node8877 = (inp[11]) ? node8887 : node8878;
													assign node8878 = (inp[14]) ? node8882 : node8879;
														assign node8879 = (inp[13]) ? 4'b0000 : 4'b1000;
														assign node8882 = (inp[13]) ? 4'b1001 : node8883;
															assign node8883 = (inp[12]) ? 4'b0001 : 4'b1001;
													assign node8887 = (inp[14]) ? 4'b0000 : node8888;
														assign node8888 = (inp[13]) ? node8892 : node8889;
															assign node8889 = (inp[12]) ? 4'b0000 : 4'b1000;
															assign node8892 = (inp[12]) ? 4'b1000 : 4'b0000;
												assign node8896 = (inp[11]) ? node8902 : node8897;
													assign node8897 = (inp[14]) ? 4'b0000 : node8898;
														assign node8898 = (inp[12]) ? 4'b1001 : 4'b0001;
													assign node8902 = (inp[10]) ? node8906 : node8903;
														assign node8903 = (inp[13]) ? 4'b1001 : 4'b0001;
														assign node8906 = (inp[13]) ? 4'b0001 : 4'b1001;
										assign node8909 = (inp[13]) ? node8911 : 4'b0001;
											assign node8911 = (inp[12]) ? 4'b0001 : node8912;
												assign node8912 = (inp[4]) ? node8914 : 4'b0001;
													assign node8914 = (inp[11]) ? 4'b0001 : node8915;
														assign node8915 = (inp[10]) ? node8917 : 4'b0000;
															assign node8917 = (inp[1]) ? node8921 : node8918;
																assign node8918 = (inp[14]) ? 4'b0001 : 4'b0000;
																assign node8921 = (inp[14]) ? 4'b0000 : 4'b0001;
							assign node8927 = (inp[2]) ? node9237 : node8928;
								assign node8928 = (inp[13]) ? node9090 : node8929;
									assign node8929 = (inp[11]) ? node9027 : node8930;
										assign node8930 = (inp[12]) ? node8978 : node8931;
											assign node8931 = (inp[10]) ? node8959 : node8932;
												assign node8932 = (inp[3]) ? node8946 : node8933;
													assign node8933 = (inp[4]) ? node8941 : node8934;
														assign node8934 = (inp[14]) ? node8938 : node8935;
															assign node8935 = (inp[1]) ? 4'b1001 : 4'b1000;
															assign node8938 = (inp[1]) ? 4'b1000 : 4'b0001;
														assign node8941 = (inp[7]) ? node8943 : 4'b1100;
															assign node8943 = (inp[1]) ? 4'b1000 : 4'b0001;
													assign node8946 = (inp[4]) ? node8952 : node8947;
														assign node8947 = (inp[7]) ? 4'b1000 : node8948;
															assign node8948 = (inp[14]) ? 4'b1000 : 4'b0000;
														assign node8952 = (inp[1]) ? 4'b1000 : node8953;
															assign node8953 = (inp[14]) ? 4'b1001 : node8954;
																assign node8954 = (inp[7]) ? 4'b1001 : 4'b1000;
												assign node8959 = (inp[4]) ? node8967 : node8960;
													assign node8960 = (inp[3]) ? node8962 : 4'b1001;
														assign node8962 = (inp[7]) ? 4'b0000 : node8963;
															assign node8963 = (inp[14]) ? 4'b1001 : 4'b1000;
													assign node8967 = (inp[7]) ? node8975 : node8968;
														assign node8968 = (inp[14]) ? node8970 : 4'b1001;
															assign node8970 = (inp[3]) ? node8972 : 4'b0000;
																assign node8972 = (inp[1]) ? 4'b0000 : 4'b1000;
														assign node8975 = (inp[1]) ? 4'b0001 : 4'b0000;
											assign node8978 = (inp[3]) ? node9008 : node8979;
												assign node8979 = (inp[7]) ? node8995 : node8980;
													assign node8980 = (inp[4]) ? node8986 : node8981;
														assign node8981 = (inp[1]) ? node8983 : 4'b0001;
															assign node8983 = (inp[14]) ? 4'b0000 : 4'b0001;
														assign node8986 = (inp[14]) ? node8992 : node8987;
															assign node8987 = (inp[1]) ? 4'b0000 : node8988;
																assign node8988 = (inp[10]) ? 4'b1100 : 4'b0100;
															assign node8992 = (inp[1]) ? 4'b0100 : 4'b0101;
													assign node8995 = (inp[10]) ? node9003 : node8996;
														assign node8996 = (inp[14]) ? node9000 : node8997;
															assign node8997 = (inp[1]) ? 4'b0001 : 4'b0000;
															assign node9000 = (inp[1]) ? 4'b0000 : 4'b0001;
														assign node9003 = (inp[1]) ? node9005 : 4'b0001;
															assign node9005 = (inp[14]) ? 4'b1000 : 4'b1001;
												assign node9008 = (inp[4]) ? node9020 : node9009;
													assign node9009 = (inp[1]) ? node9015 : node9010;
														assign node9010 = (inp[10]) ? node9012 : 4'b0000;
															assign node9012 = (inp[7]) ? 4'b1000 : 4'b0000;
														assign node9015 = (inp[10]) ? node9017 : 4'b1000;
															assign node9017 = (inp[7]) ? 4'b0000 : 4'b1000;
													assign node9020 = (inp[1]) ? 4'b0000 : node9021;
														assign node9021 = (inp[14]) ? 4'b0001 : node9022;
															assign node9022 = (inp[10]) ? 4'b0001 : 4'b1000;
										assign node9027 = (inp[1]) ? node9067 : node9028;
											assign node9028 = (inp[3]) ? node9048 : node9029;
												assign node9029 = (inp[10]) ? node9037 : node9030;
													assign node9030 = (inp[12]) ? 4'b0000 : node9031;
														assign node9031 = (inp[4]) ? node9033 : 4'b1000;
															assign node9033 = (inp[7]) ? 4'b1000 : 4'b1100;
													assign node9037 = (inp[12]) ? node9043 : node9038;
														assign node9038 = (inp[4]) ? node9040 : 4'b1000;
															assign node9040 = (inp[14]) ? 4'b0001 : 4'b1000;
														assign node9043 = (inp[7]) ? 4'b1000 : node9044;
															assign node9044 = (inp[4]) ? 4'b1100 : 4'b1000;
												assign node9048 = (inp[7]) ? node9060 : node9049;
													assign node9049 = (inp[10]) ? node9055 : node9050;
														assign node9050 = (inp[14]) ? node9052 : 4'b0001;
															assign node9052 = (inp[12]) ? 4'b1000 : 4'b0001;
														assign node9055 = (inp[12]) ? node9057 : 4'b1000;
															assign node9057 = (inp[4]) ? 4'b0001 : 4'b0000;
													assign node9060 = (inp[14]) ? node9062 : 4'b1001;
														assign node9062 = (inp[4]) ? node9064 : 4'b0001;
															assign node9064 = (inp[10]) ? 4'b0001 : 4'b1001;
											assign node9067 = (inp[4]) ? node9075 : node9068;
												assign node9068 = (inp[10]) ? 4'b1001 : node9069;
													assign node9069 = (inp[3]) ? 4'b1001 : node9070;
														assign node9070 = (inp[12]) ? 4'b0001 : 4'b1001;
												assign node9075 = (inp[10]) ? node9085 : node9076;
													assign node9076 = (inp[3]) ? node9080 : node9077;
														assign node9077 = (inp[14]) ? 4'b0101 : 4'b1101;
														assign node9080 = (inp[12]) ? 4'b1001 : node9081;
															assign node9081 = (inp[7]) ? 4'b1001 : 4'b0001;
													assign node9085 = (inp[12]) ? node9087 : 4'b0001;
														assign node9087 = (inp[7]) ? 4'b1001 : 4'b0001;
									assign node9090 = (inp[3]) ? node9168 : node9091;
										assign node9091 = (inp[10]) ? node9129 : node9092;
											assign node9092 = (inp[12]) ? node9116 : node9093;
												assign node9093 = (inp[14]) ? node9107 : node9094;
													assign node9094 = (inp[1]) ? node9096 : 4'b0100;
														assign node9096 = (inp[11]) ? node9102 : node9097;
															assign node9097 = (inp[4]) ? 4'b0101 : node9098;
																assign node9098 = (inp[7]) ? 4'b0001 : 4'b0101;
															assign node9102 = (inp[4]) ? 4'b1001 : node9103;
																assign node9103 = (inp[7]) ? 4'b0001 : 4'b0101;
													assign node9107 = (inp[7]) ? node9111 : node9108;
														assign node9108 = (inp[11]) ? 4'b1001 : 4'b1000;
														assign node9111 = (inp[4]) ? node9113 : 4'b1001;
															assign node9113 = (inp[1]) ? 4'b0101 : 4'b0100;
												assign node9116 = (inp[1]) ? node9124 : node9117;
													assign node9117 = (inp[14]) ? node9121 : node9118;
														assign node9118 = (inp[4]) ? 4'b0000 : 4'b1000;
														assign node9121 = (inp[7]) ? 4'b1001 : 4'b0001;
													assign node9124 = (inp[11]) ? 4'b1001 : node9125;
														assign node9125 = (inp[14]) ? 4'b1000 : 4'b1001;
											assign node9129 = (inp[11]) ? node9153 : node9130;
												assign node9130 = (inp[12]) ? node9142 : node9131;
													assign node9131 = (inp[4]) ? 4'b0000 : node9132;
														assign node9132 = (inp[7]) ? node9136 : node9133;
															assign node9133 = (inp[14]) ? 4'b0101 : 4'b0100;
															assign node9136 = (inp[14]) ? node9138 : 4'b0001;
																assign node9138 = (inp[1]) ? 4'b0000 : 4'b0001;
													assign node9142 = (inp[1]) ? node9150 : node9143;
														assign node9143 = (inp[14]) ? node9145 : 4'b1000;
															assign node9145 = (inp[7]) ? 4'b1001 : node9146;
																assign node9146 = (inp[4]) ? 4'b1000 : 4'b1001;
														assign node9150 = (inp[7]) ? 4'b0001 : 4'b0000;
												assign node9153 = (inp[1]) ? node9163 : node9154;
													assign node9154 = (inp[4]) ? node9158 : node9155;
														assign node9155 = (inp[7]) ? 4'b0000 : 4'b0100;
														assign node9158 = (inp[12]) ? node9160 : 4'b0001;
															assign node9160 = (inp[7]) ? 4'b0100 : 4'b1001;
													assign node9163 = (inp[7]) ? 4'b0001 : node9164;
														assign node9164 = (inp[4]) ? 4'b0001 : 4'b0101;
										assign node9168 = (inp[4]) ? node9208 : node9169;
											assign node9169 = (inp[10]) ? node9187 : node9170;
												assign node9170 = (inp[1]) ? node9180 : node9171;
													assign node9171 = (inp[11]) ? 4'b0000 : node9172;
														assign node9172 = (inp[14]) ? 4'b0000 : node9173;
															assign node9173 = (inp[7]) ? node9175 : 4'b1001;
																assign node9175 = (inp[12]) ? 4'b0000 : 4'b0001;
													assign node9180 = (inp[14]) ? 4'b0001 : node9181;
														assign node9181 = (inp[11]) ? 4'b0001 : node9182;
															assign node9182 = (inp[12]) ? 4'b0000 : 4'b0001;
												assign node9187 = (inp[1]) ? node9201 : node9188;
													assign node9188 = (inp[7]) ? node9194 : node9189;
														assign node9189 = (inp[12]) ? node9191 : 4'b1001;
															assign node9191 = (inp[11]) ? 4'b1001 : 4'b0001;
														assign node9194 = (inp[11]) ? node9198 : node9195;
															assign node9195 = (inp[14]) ? 4'b1000 : 4'b1001;
															assign node9198 = (inp[12]) ? 4'b1000 : 4'b0000;
													assign node9201 = (inp[11]) ? 4'b0001 : node9202;
														assign node9202 = (inp[7]) ? 4'b0000 : node9203;
															assign node9203 = (inp[12]) ? 4'b1001 : 4'b0000;
											assign node9208 = (inp[10]) ? node9224 : node9209;
												assign node9209 = (inp[1]) ? node9219 : node9210;
													assign node9210 = (inp[7]) ? 4'b0000 : node9211;
														assign node9211 = (inp[12]) ? node9213 : 4'b0001;
															assign node9213 = (inp[14]) ? 4'b0000 : node9214;
																assign node9214 = (inp[11]) ? 4'b0000 : 4'b0001;
													assign node9219 = (inp[11]) ? 4'b0001 : node9220;
														assign node9220 = (inp[7]) ? 4'b0000 : 4'b0001;
												assign node9224 = (inp[1]) ? 4'b0000 : node9225;
													assign node9225 = (inp[11]) ? 4'b0000 : node9226;
														assign node9226 = (inp[12]) ? 4'b0001 : node9227;
															assign node9227 = (inp[7]) ? node9231 : node9228;
																assign node9228 = (inp[14]) ? 4'b0001 : 4'b0000;
																assign node9231 = (inp[14]) ? 4'b0000 : 4'b0001;
								assign node9237 = (inp[3]) ? node9239 : 4'b0001;
									assign node9239 = (inp[4]) ? node9257 : node9240;
										assign node9240 = (inp[7]) ? 4'b0001 : node9241;
											assign node9241 = (inp[13]) ? node9243 : 4'b0001;
												assign node9243 = (inp[12]) ? node9251 : node9244;
													assign node9244 = (inp[1]) ? node9248 : node9245;
														assign node9245 = (inp[11]) ? 4'b0000 : 4'b0001;
														assign node9248 = (inp[10]) ? 4'b0001 : 4'b0000;
													assign node9251 = (inp[10]) ? node9253 : 4'b0001;
														assign node9253 = (inp[1]) ? 4'b0001 : 4'b0000;
										assign node9257 = (inp[13]) ? node9279 : node9258;
											assign node9258 = (inp[7]) ? 4'b0001 : node9259;
												assign node9259 = (inp[11]) ? node9269 : node9260;
													assign node9260 = (inp[10]) ? node9264 : node9261;
														assign node9261 = (inp[12]) ? 4'b0001 : 4'b1000;
														assign node9264 = (inp[1]) ? 4'b0000 : node9265;
															assign node9265 = (inp[14]) ? 4'b0000 : 4'b1000;
													assign node9269 = (inp[1]) ? node9273 : node9270;
														assign node9270 = (inp[12]) ? 4'b1000 : 4'b0001;
														assign node9273 = (inp[10]) ? 4'b0001 : node9274;
															assign node9274 = (inp[12]) ? 4'b0001 : 4'b1001;
											assign node9279 = (inp[10]) ? node9299 : node9280;
												assign node9280 = (inp[12]) ? node9292 : node9281;
													assign node9281 = (inp[7]) ? node9285 : node9282;
														assign node9282 = (inp[14]) ? 4'b0000 : 4'b0001;
														assign node9285 = (inp[11]) ? 4'b0000 : node9286;
															assign node9286 = (inp[1]) ? 4'b0000 : node9287;
																assign node9287 = (inp[14]) ? 4'b0001 : 4'b0000;
													assign node9292 = (inp[7]) ? 4'b0001 : node9293;
														assign node9293 = (inp[1]) ? node9295 : 4'b0000;
															assign node9295 = (inp[14]) ? 4'b0001 : 4'b0000;
												assign node9299 = (inp[11]) ? 4'b0000 : node9300;
													assign node9300 = (inp[14]) ? 4'b0000 : node9301;
														assign node9301 = (inp[12]) ? 4'b0000 : 4'b0001;
		assign node9306 = (inp[9]) ? node14048 : node9307;
			assign node9307 = (inp[15]) ? node11965 : node9308;
				assign node9308 = (inp[6]) ? node9942 : node9309;
					assign node9309 = (inp[0]) ? 4'b1100 : node9310;
						assign node9310 = (inp[5]) ? node9540 : node9311;
							assign node9311 = (inp[2]) ? 4'b1110 : node9312;
								assign node9312 = (inp[3]) ? node9418 : node9313;
									assign node9313 = (inp[7]) ? node9383 : node9314;
										assign node9314 = (inp[1]) ? node9344 : node9315;
											assign node9315 = (inp[13]) ? node9327 : node9316;
												assign node9316 = (inp[4]) ? node9324 : node9317;
													assign node9317 = (inp[14]) ? node9319 : 4'b1110;
														assign node9319 = (inp[12]) ? 4'b1110 : node9320;
															assign node9320 = (inp[11]) ? 4'b0001 : 4'b0000;
													assign node9324 = (inp[10]) ? 4'b0001 : 4'b1001;
												assign node9327 = (inp[12]) ? node9339 : node9328;
													assign node9328 = (inp[10]) ? node9334 : node9329;
														assign node9329 = (inp[14]) ? node9331 : 4'b0001;
															assign node9331 = (inp[11]) ? 4'b0001 : 4'b0000;
														assign node9334 = (inp[11]) ? 4'b1001 : node9335;
															assign node9335 = (inp[14]) ? 4'b1000 : 4'b1001;
													assign node9339 = (inp[14]) ? node9341 : 4'b0001;
														assign node9341 = (inp[11]) ? 4'b0001 : 4'b0000;
											assign node9344 = (inp[4]) ? node9358 : node9345;
												assign node9345 = (inp[13]) ? 4'b1000 : node9346;
													assign node9346 = (inp[10]) ? node9348 : 4'b1110;
														assign node9348 = (inp[12]) ? node9352 : node9349;
															assign node9349 = (inp[11]) ? 4'b0000 : 4'b0001;
															assign node9352 = (inp[11]) ? 4'b0000 : node9353;
																assign node9353 = (inp[14]) ? 4'b1110 : 4'b0000;
												assign node9358 = (inp[14]) ? node9368 : node9359;
													assign node9359 = (inp[10]) ? 4'b0000 : node9360;
														assign node9360 = (inp[12]) ? node9364 : node9361;
															assign node9361 = (inp[13]) ? 4'b1000 : 4'b0000;
															assign node9364 = (inp[13]) ? 4'b0000 : 4'b1000;
													assign node9368 = (inp[11]) ? node9376 : node9369;
														assign node9369 = (inp[13]) ? 4'b0001 : node9370;
															assign node9370 = (inp[10]) ? node9372 : 4'b1001;
																assign node9372 = (inp[12]) ? 4'b1001 : 4'b0001;
														assign node9376 = (inp[13]) ? node9380 : node9377;
															assign node9377 = (inp[10]) ? 4'b0000 : 4'b1000;
															assign node9380 = (inp[10]) ? 4'b1000 : 4'b0000;
										assign node9383 = (inp[4]) ? node9385 : 4'b1110;
											assign node9385 = (inp[13]) ? node9399 : node9386;
												assign node9386 = (inp[1]) ? node9388 : 4'b1110;
													assign node9388 = (inp[12]) ? node9392 : node9389;
														assign node9389 = (inp[11]) ? 4'b0000 : 4'b0001;
														assign node9392 = (inp[10]) ? node9394 : 4'b1110;
															assign node9394 = (inp[11]) ? 4'b0000 : node9395;
																assign node9395 = (inp[14]) ? 4'b1110 : 4'b0000;
												assign node9399 = (inp[1]) ? node9409 : node9400;
													assign node9400 = (inp[12]) ? node9404 : node9401;
														assign node9401 = (inp[14]) ? 4'b1000 : 4'b1001;
														assign node9404 = (inp[11]) ? 4'b0001 : node9405;
															assign node9405 = (inp[14]) ? 4'b0000 : 4'b0001;
													assign node9409 = (inp[14]) ? node9411 : 4'b1000;
														assign node9411 = (inp[11]) ? node9415 : node9412;
															assign node9412 = (inp[10]) ? 4'b1001 : 4'b0001;
															assign node9415 = (inp[10]) ? 4'b1000 : 4'b0000;
									assign node9418 = (inp[4]) ? node9488 : node9419;
										assign node9419 = (inp[7]) ? node9451 : node9420;
											assign node9420 = (inp[13]) ? node9434 : node9421;
												assign node9421 = (inp[12]) ? node9429 : node9422;
													assign node9422 = (inp[10]) ? 4'b0100 : node9423;
														assign node9423 = (inp[11]) ? node9425 : 4'b1001;
															assign node9425 = (inp[1]) ? 4'b0100 : 4'b1001;
													assign node9429 = (inp[1]) ? node9431 : 4'b1001;
														assign node9431 = (inp[14]) ? 4'b1001 : 4'b1000;
												assign node9434 = (inp[1]) ? node9440 : node9435;
													assign node9435 = (inp[10]) ? node9437 : 4'b0101;
														assign node9437 = (inp[12]) ? 4'b0101 : 4'b1101;
													assign node9440 = (inp[12]) ? node9446 : node9441;
														assign node9441 = (inp[11]) ? 4'b1100 : node9442;
															assign node9442 = (inp[14]) ? 4'b0101 : 4'b1100;
														assign node9446 = (inp[14]) ? 4'b0101 : node9447;
															assign node9447 = (inp[10]) ? 4'b1100 : 4'b0100;
											assign node9451 = (inp[1]) ? node9471 : node9452;
												assign node9452 = (inp[11]) ? node9462 : node9453;
													assign node9453 = (inp[14]) ? node9457 : node9454;
														assign node9454 = (inp[13]) ? 4'b0001 : 4'b1001;
														assign node9457 = (inp[12]) ? 4'b1000 : node9458;
															assign node9458 = (inp[13]) ? 4'b1000 : 4'b0000;
													assign node9462 = (inp[13]) ? node9466 : node9463;
														assign node9463 = (inp[10]) ? 4'b0001 : 4'b1001;
														assign node9466 = (inp[12]) ? 4'b0001 : node9467;
															assign node9467 = (inp[10]) ? 4'b1001 : 4'b0001;
												assign node9471 = (inp[14]) ? node9479 : node9472;
													assign node9472 = (inp[13]) ? 4'b1000 : node9473;
														assign node9473 = (inp[12]) ? node9475 : 4'b0000;
															assign node9475 = (inp[10]) ? 4'b0000 : 4'b1000;
													assign node9479 = (inp[11]) ? node9485 : node9480;
														assign node9480 = (inp[13]) ? 4'b0001 : node9481;
															assign node9481 = (inp[12]) ? 4'b1001 : 4'b0001;
														assign node9485 = (inp[13]) ? 4'b1000 : 4'b0000;
										assign node9488 = (inp[1]) ? node9514 : node9489;
											assign node9489 = (inp[13]) ? node9505 : node9490;
												assign node9490 = (inp[7]) ? 4'b1001 : node9491;
													assign node9491 = (inp[11]) ? node9499 : node9492;
														assign node9492 = (inp[14]) ? node9494 : 4'b1101;
															assign node9494 = (inp[12]) ? 4'b1100 : node9495;
																assign node9495 = (inp[10]) ? 4'b0100 : 4'b1100;
														assign node9499 = (inp[10]) ? node9501 : 4'b1101;
															assign node9501 = (inp[12]) ? 4'b1101 : 4'b0101;
												assign node9505 = (inp[10]) ? node9511 : node9506;
													assign node9506 = (inp[14]) ? node9508 : 4'b0101;
														assign node9508 = (inp[11]) ? 4'b0101 : 4'b0100;
													assign node9511 = (inp[12]) ? 4'b0101 : 4'b1101;
											assign node9514 = (inp[14]) ? node9528 : node9515;
												assign node9515 = (inp[13]) ? node9523 : node9516;
													assign node9516 = (inp[10]) ? 4'b0100 : node9517;
														assign node9517 = (inp[12]) ? node9519 : 4'b0100;
															assign node9519 = (inp[7]) ? 4'b1000 : 4'b1100;
													assign node9523 = (inp[10]) ? 4'b1100 : node9524;
														assign node9524 = (inp[12]) ? 4'b0100 : 4'b1100;
												assign node9528 = (inp[11]) ? 4'b1100 : node9529;
													assign node9529 = (inp[13]) ? node9535 : node9530;
														assign node9530 = (inp[7]) ? 4'b1001 : node9531;
															assign node9531 = (inp[12]) ? 4'b1101 : 4'b0101;
														assign node9535 = (inp[12]) ? 4'b0101 : 4'b1101;
							assign node9540 = (inp[1]) ? node9756 : node9541;
								assign node9541 = (inp[13]) ? node9661 : node9542;
									assign node9542 = (inp[14]) ? node9586 : node9543;
										assign node9543 = (inp[10]) ? node9559 : node9544;
											assign node9544 = (inp[3]) ? node9554 : node9545;
												assign node9545 = (inp[4]) ? node9549 : node9546;
													assign node9546 = (inp[2]) ? 4'b1110 : 4'b1101;
													assign node9549 = (inp[7]) ? node9551 : 4'b1001;
														assign node9551 = (inp[2]) ? 4'b1110 : 4'b1101;
												assign node9554 = (inp[4]) ? node9556 : 4'b1001;
													assign node9556 = (inp[7]) ? 4'b1001 : 4'b1101;
											assign node9559 = (inp[12]) ? node9573 : node9560;
												assign node9560 = (inp[3]) ? node9568 : node9561;
													assign node9561 = (inp[7]) ? node9563 : 4'b0001;
														assign node9563 = (inp[4]) ? 4'b0001 : node9564;
															assign node9564 = (inp[2]) ? 4'b1110 : 4'b0101;
													assign node9568 = (inp[7]) ? node9570 : 4'b0101;
														assign node9570 = (inp[4]) ? 4'b0101 : 4'b0001;
												assign node9573 = (inp[3]) ? node9581 : node9574;
													assign node9574 = (inp[7]) ? node9578 : node9575;
														assign node9575 = (inp[4]) ? 4'b1001 : 4'b1101;
														assign node9578 = (inp[2]) ? 4'b1110 : 4'b1101;
													assign node9581 = (inp[4]) ? node9583 : 4'b1001;
														assign node9583 = (inp[2]) ? 4'b1001 : 4'b1101;
										assign node9586 = (inp[11]) ? node9628 : node9587;
											assign node9587 = (inp[12]) ? node9607 : node9588;
												assign node9588 = (inp[10]) ? node9596 : node9589;
													assign node9589 = (inp[3]) ? 4'b1000 : node9590;
														assign node9590 = (inp[2]) ? 4'b1110 : node9591;
															assign node9591 = (inp[4]) ? 4'b1000 : 4'b1100;
													assign node9596 = (inp[2]) ? node9598 : 4'b0000;
														assign node9598 = (inp[3]) ? node9602 : node9599;
															assign node9599 = (inp[7]) ? 4'b1110 : 4'b0000;
															assign node9602 = (inp[7]) ? node9604 : 4'b0100;
																assign node9604 = (inp[4]) ? 4'b0100 : 4'b0000;
												assign node9607 = (inp[2]) ? node9619 : node9608;
													assign node9608 = (inp[7]) ? 4'b1000 : node9609;
														assign node9609 = (inp[10]) ? node9613 : node9610;
															assign node9610 = (inp[4]) ? 4'b1000 : 4'b1100;
															assign node9613 = (inp[4]) ? 4'b1100 : node9614;
																assign node9614 = (inp[3]) ? 4'b1000 : 4'b1100;
													assign node9619 = (inp[4]) ? node9621 : 4'b1110;
														assign node9621 = (inp[7]) ? node9625 : node9622;
															assign node9622 = (inp[3]) ? 4'b1100 : 4'b1000;
															assign node9625 = (inp[10]) ? 4'b1000 : 4'b1110;
											assign node9628 = (inp[3]) ? node9644 : node9629;
												assign node9629 = (inp[2]) ? node9637 : node9630;
													assign node9630 = (inp[7]) ? 4'b1101 : node9631;
														assign node9631 = (inp[12]) ? node9633 : 4'b0001;
															assign node9633 = (inp[4]) ? 4'b1001 : 4'b1101;
													assign node9637 = (inp[10]) ? node9639 : 4'b1110;
														assign node9639 = (inp[4]) ? node9641 : 4'b1110;
															assign node9641 = (inp[7]) ? 4'b1110 : 4'b1001;
												assign node9644 = (inp[4]) ? node9650 : node9645;
													assign node9645 = (inp[12]) ? 4'b1001 : node9646;
														assign node9646 = (inp[10]) ? 4'b0001 : 4'b1001;
													assign node9650 = (inp[7]) ? node9656 : node9651;
														assign node9651 = (inp[10]) ? node9653 : 4'b1101;
															assign node9653 = (inp[2]) ? 4'b1101 : 4'b0101;
														assign node9656 = (inp[10]) ? node9658 : 4'b1001;
															assign node9658 = (inp[12]) ? 4'b1001 : 4'b0101;
									assign node9661 = (inp[10]) ? node9693 : node9662;
										assign node9662 = (inp[3]) ? node9678 : node9663;
											assign node9663 = (inp[7]) ? node9669 : node9664;
												assign node9664 = (inp[11]) ? 4'b0001 : node9665;
													assign node9665 = (inp[14]) ? 4'b0000 : 4'b0001;
												assign node9669 = (inp[4]) ? 4'b0001 : node9670;
													assign node9670 = (inp[2]) ? 4'b1110 : node9671;
														assign node9671 = (inp[14]) ? node9673 : 4'b0101;
															assign node9673 = (inp[11]) ? 4'b0101 : 4'b0100;
											assign node9678 = (inp[4]) ? node9688 : node9679;
												assign node9679 = (inp[7]) ? node9683 : node9680;
													assign node9680 = (inp[11]) ? 4'b0101 : 4'b0100;
													assign node9683 = (inp[2]) ? 4'b0001 : node9684;
														assign node9684 = (inp[14]) ? 4'b0000 : 4'b0001;
												assign node9688 = (inp[11]) ? 4'b0101 : node9689;
													assign node9689 = (inp[14]) ? 4'b0100 : 4'b0101;
										assign node9693 = (inp[12]) ? node9727 : node9694;
											assign node9694 = (inp[14]) ? node9706 : node9695;
												assign node9695 = (inp[3]) ? 4'b1101 : node9696;
													assign node9696 = (inp[11]) ? node9698 : 4'b1001;
														assign node9698 = (inp[7]) ? node9700 : 4'b1001;
															assign node9700 = (inp[4]) ? 4'b1001 : node9701;
																assign node9701 = (inp[2]) ? 4'b1110 : 4'b1101;
												assign node9706 = (inp[11]) ? node9718 : node9707;
													assign node9707 = (inp[3]) ? node9715 : node9708;
														assign node9708 = (inp[7]) ? node9710 : 4'b1000;
															assign node9710 = (inp[4]) ? 4'b1000 : node9711;
																assign node9711 = (inp[2]) ? 4'b1110 : 4'b1100;
														assign node9715 = (inp[7]) ? 4'b1000 : 4'b1100;
													assign node9718 = (inp[4]) ? node9724 : node9719;
														assign node9719 = (inp[3]) ? 4'b1001 : node9720;
															assign node9720 = (inp[2]) ? 4'b1110 : 4'b1101;
														assign node9724 = (inp[3]) ? 4'b1101 : 4'b1001;
											assign node9727 = (inp[11]) ? node9743 : node9728;
												assign node9728 = (inp[14]) ? node9736 : node9729;
													assign node9729 = (inp[2]) ? node9731 : 4'b0001;
														assign node9731 = (inp[4]) ? node9733 : 4'b1110;
															assign node9733 = (inp[7]) ? 4'b0001 : 4'b0101;
													assign node9736 = (inp[2]) ? node9740 : node9737;
														assign node9737 = (inp[4]) ? 4'b0000 : 4'b0100;
														assign node9740 = (inp[4]) ? 4'b0100 : 4'b1110;
												assign node9743 = (inp[3]) ? node9751 : node9744;
													assign node9744 = (inp[7]) ? node9746 : 4'b0001;
														assign node9746 = (inp[4]) ? 4'b0001 : node9747;
															assign node9747 = (inp[2]) ? 4'b1110 : 4'b0101;
													assign node9751 = (inp[7]) ? node9753 : 4'b0101;
														assign node9753 = (inp[4]) ? 4'b0101 : 4'b0001;
								assign node9756 = (inp[3]) ? node9848 : node9757;
									assign node9757 = (inp[7]) ? node9797 : node9758;
										assign node9758 = (inp[14]) ? node9774 : node9759;
											assign node9759 = (inp[13]) ? node9769 : node9760;
												assign node9760 = (inp[12]) ? node9762 : 4'b0000;
													assign node9762 = (inp[10]) ? 4'b0000 : node9763;
														assign node9763 = (inp[4]) ? 4'b1000 : node9764;
															assign node9764 = (inp[2]) ? 4'b1110 : 4'b1100;
												assign node9769 = (inp[12]) ? node9771 : 4'b1000;
													assign node9771 = (inp[10]) ? 4'b1000 : 4'b0000;
											assign node9774 = (inp[11]) ? node9790 : node9775;
												assign node9775 = (inp[13]) ? node9785 : node9776;
													assign node9776 = (inp[12]) ? node9780 : node9777;
														assign node9777 = (inp[4]) ? 4'b1001 : 4'b0001;
														assign node9780 = (inp[4]) ? 4'b1001 : node9781;
															assign node9781 = (inp[10]) ? 4'b1110 : 4'b1101;
													assign node9785 = (inp[12]) ? 4'b0001 : node9786;
														assign node9786 = (inp[10]) ? 4'b1001 : 4'b0001;
												assign node9790 = (inp[13]) ? node9792 : 4'b0000;
													assign node9792 = (inp[10]) ? 4'b1000 : node9793;
														assign node9793 = (inp[12]) ? 4'b0000 : 4'b1000;
										assign node9797 = (inp[4]) ? node9817 : node9798;
											assign node9798 = (inp[2]) ? 4'b1110 : node9799;
												assign node9799 = (inp[13]) ? node9807 : node9800;
													assign node9800 = (inp[11]) ? 4'b0100 : node9801;
														assign node9801 = (inp[14]) ? node9803 : 4'b0100;
															assign node9803 = (inp[10]) ? 4'b0101 : 4'b1101;
													assign node9807 = (inp[12]) ? node9813 : node9808;
														assign node9808 = (inp[11]) ? 4'b1100 : node9809;
															assign node9809 = (inp[10]) ? 4'b1101 : 4'b1100;
														assign node9813 = (inp[10]) ? 4'b1100 : 4'b0100;
											assign node9817 = (inp[13]) ? node9831 : node9818;
												assign node9818 = (inp[10]) ? node9826 : node9819;
													assign node9819 = (inp[11]) ? node9821 : 4'b1110;
														assign node9821 = (inp[14]) ? 4'b0000 : node9822;
															assign node9822 = (inp[2]) ? 4'b1110 : 4'b1100;
													assign node9826 = (inp[14]) ? node9828 : 4'b0000;
														assign node9828 = (inp[2]) ? 4'b0000 : 4'b1101;
												assign node9831 = (inp[14]) ? node9837 : node9832;
													assign node9832 = (inp[12]) ? node9834 : 4'b1000;
														assign node9834 = (inp[10]) ? 4'b1000 : 4'b0000;
													assign node9837 = (inp[11]) ? node9843 : node9838;
														assign node9838 = (inp[12]) ? 4'b0001 : node9839;
															assign node9839 = (inp[10]) ? 4'b1001 : 4'b0001;
														assign node9843 = (inp[12]) ? node9845 : 4'b1000;
															assign node9845 = (inp[10]) ? 4'b1000 : 4'b0000;
									assign node9848 = (inp[14]) ? node9886 : node9849;
										assign node9849 = (inp[7]) ? node9863 : node9850;
											assign node9850 = (inp[13]) ? node9858 : node9851;
												assign node9851 = (inp[12]) ? node9853 : 4'b0100;
													assign node9853 = (inp[10]) ? 4'b0100 : node9854;
														assign node9854 = (inp[4]) ? 4'b1100 : 4'b1000;
												assign node9858 = (inp[12]) ? node9860 : 4'b1100;
													assign node9860 = (inp[10]) ? 4'b1100 : 4'b0100;
											assign node9863 = (inp[4]) ? node9877 : node9864;
												assign node9864 = (inp[2]) ? 4'b0000 : node9865;
													assign node9865 = (inp[13]) ? node9871 : node9866;
														assign node9866 = (inp[10]) ? 4'b0000 : node9867;
															assign node9867 = (inp[12]) ? 4'b1000 : 4'b0000;
														assign node9871 = (inp[12]) ? node9873 : 4'b1000;
															assign node9873 = (inp[11]) ? 4'b0000 : 4'b1000;
												assign node9877 = (inp[12]) ? node9881 : node9878;
													assign node9878 = (inp[13]) ? 4'b1100 : 4'b0100;
													assign node9881 = (inp[13]) ? node9883 : 4'b1000;
														assign node9883 = (inp[10]) ? 4'b1100 : 4'b0100;
										assign node9886 = (inp[11]) ? node9912 : node9887;
											assign node9887 = (inp[13]) ? node9903 : node9888;
												assign node9888 = (inp[7]) ? node9898 : node9889;
													assign node9889 = (inp[12]) ? node9895 : node9890;
														assign node9890 = (inp[10]) ? 4'b0101 : node9891;
															assign node9891 = (inp[4]) ? 4'b1101 : 4'b1001;
														assign node9895 = (inp[4]) ? 4'b1101 : 4'b1001;
													assign node9898 = (inp[10]) ? node9900 : 4'b1001;
														assign node9900 = (inp[12]) ? 4'b1001 : 4'b0001;
												assign node9903 = (inp[12]) ? node9907 : node9904;
													assign node9904 = (inp[10]) ? 4'b1101 : 4'b0101;
													assign node9907 = (inp[7]) ? node9909 : 4'b0101;
														assign node9909 = (inp[4]) ? 4'b0101 : 4'b0001;
											assign node9912 = (inp[4]) ? node9928 : node9913;
												assign node9913 = (inp[7]) ? node9923 : node9914;
													assign node9914 = (inp[12]) ? node9916 : 4'b0100;
														assign node9916 = (inp[10]) ? node9920 : node9917;
															assign node9917 = (inp[13]) ? 4'b0100 : 4'b1000;
															assign node9920 = (inp[13]) ? 4'b1100 : 4'b0100;
													assign node9923 = (inp[12]) ? 4'b0000 : node9924;
														assign node9924 = (inp[13]) ? 4'b1000 : 4'b0000;
												assign node9928 = (inp[13]) ? node9936 : node9929;
													assign node9929 = (inp[10]) ? 4'b0100 : node9930;
														assign node9930 = (inp[12]) ? node9932 : 4'b0100;
															assign node9932 = (inp[2]) ? 4'b1000 : 4'b1100;
													assign node9936 = (inp[12]) ? node9938 : 4'b1100;
														assign node9938 = (inp[10]) ? 4'b1100 : 4'b0100;
					assign node9942 = (inp[5]) ? node10776 : node9943;
						assign node9943 = (inp[0]) ? node10519 : node9944;
							assign node9944 = (inp[11]) ? node10244 : node9945;
								assign node9945 = (inp[10]) ? node10095 : node9946;
									assign node9946 = (inp[13]) ? node10014 : node9947;
										assign node9947 = (inp[4]) ? node9985 : node9948;
											assign node9948 = (inp[2]) ? node9962 : node9949;
												assign node9949 = (inp[1]) ? node9955 : node9950;
													assign node9950 = (inp[3]) ? 4'b1101 : node9951;
														assign node9951 = (inp[14]) ? 4'b1100 : 4'b1101;
													assign node9955 = (inp[12]) ? 4'b1101 : node9956;
														assign node9956 = (inp[7]) ? node9958 : 4'b0001;
															assign node9958 = (inp[3]) ? 4'b0101 : 4'b1101;
												assign node9962 = (inp[3]) ? node9974 : node9963;
													assign node9963 = (inp[7]) ? node9969 : node9964;
														assign node9964 = (inp[1]) ? 4'b1101 : node9965;
															assign node9965 = (inp[14]) ? 4'b1100 : 4'b1101;
														assign node9969 = (inp[1]) ? 4'b1100 : node9970;
															assign node9970 = (inp[14]) ? 4'b1100 : 4'b1101;
													assign node9974 = (inp[12]) ? node9980 : node9975;
														assign node9975 = (inp[14]) ? node9977 : 4'b0000;
															assign node9977 = (inp[1]) ? 4'b1001 : 4'b1000;
														assign node9980 = (inp[14]) ? 4'b1001 : node9981;
															assign node9981 = (inp[1]) ? 4'b1000 : 4'b1001;
											assign node9985 = (inp[1]) ? node9997 : node9986;
												assign node9986 = (inp[3]) ? node9992 : node9987;
													assign node9987 = (inp[2]) ? node9989 : 4'b1001;
														assign node9989 = (inp[14]) ? 4'b1000 : 4'b1101;
													assign node9992 = (inp[14]) ? 4'b1001 : node9993;
														assign node9993 = (inp[12]) ? 4'b1001 : 4'b0000;
												assign node9997 = (inp[2]) ? node10005 : node9998;
													assign node9998 = (inp[3]) ? node10002 : node9999;
														assign node9999 = (inp[12]) ? 4'b1001 : 4'b0001;
														assign node10002 = (inp[14]) ? 4'b0000 : 4'b0001;
													assign node10005 = (inp[12]) ? 4'b1001 : node10006;
														assign node10006 = (inp[14]) ? node10010 : node10007;
															assign node10007 = (inp[7]) ? 4'b0001 : 4'b0101;
															assign node10010 = (inp[7]) ? 4'b1101 : 4'b1001;
										assign node10014 = (inp[2]) ? node10052 : node10015;
											assign node10015 = (inp[4]) ? node10031 : node10016;
												assign node10016 = (inp[7]) ? node10022 : node10017;
													assign node10017 = (inp[12]) ? 4'b1001 : node10018;
														assign node10018 = (inp[1]) ? 4'b0001 : 4'b1001;
													assign node10022 = (inp[3]) ? node10026 : node10023;
														assign node10023 = (inp[12]) ? 4'b0101 : 4'b0001;
														assign node10026 = (inp[1]) ? node10028 : 4'b1101;
															assign node10028 = (inp[12]) ? 4'b1101 : 4'b0001;
												assign node10031 = (inp[7]) ? node10045 : node10032;
													assign node10032 = (inp[3]) ? node10038 : node10033;
														assign node10033 = (inp[12]) ? 4'b1101 : node10034;
															assign node10034 = (inp[1]) ? 4'b0101 : 4'b1101;
														assign node10038 = (inp[12]) ? node10040 : 4'b1100;
															assign node10040 = (inp[1]) ? node10042 : 4'b0101;
																assign node10042 = (inp[14]) ? 4'b1100 : 4'b1101;
													assign node10045 = (inp[3]) ? 4'b0001 : node10046;
														assign node10046 = (inp[1]) ? node10048 : 4'b1001;
															assign node10048 = (inp[12]) ? 4'b1001 : 4'b0101;
											assign node10052 = (inp[3]) ? node10082 : node10053;
												assign node10053 = (inp[7]) ? node10065 : node10054;
													assign node10054 = (inp[12]) ? node10060 : node10055;
														assign node10055 = (inp[1]) ? 4'b0001 : node10056;
															assign node10056 = (inp[14]) ? 4'b0000 : 4'b0001;
														assign node10060 = (inp[1]) ? 4'b0000 : node10061;
															assign node10061 = (inp[14]) ? 4'b0000 : 4'b0001;
													assign node10065 = (inp[4]) ? node10075 : node10066;
														assign node10066 = (inp[12]) ? node10068 : 4'b0101;
															assign node10068 = (inp[1]) ? node10072 : node10069;
																assign node10069 = (inp[14]) ? 4'b0100 : 4'b0101;
																assign node10072 = (inp[14]) ? 4'b0101 : 4'b0100;
														assign node10075 = (inp[1]) ? node10079 : node10076;
															assign node10076 = (inp[14]) ? 4'b0000 : 4'b0001;
															assign node10079 = (inp[14]) ? 4'b0001 : 4'b0000;
												assign node10082 = (inp[4]) ? node10088 : node10083;
													assign node10083 = (inp[7]) ? node10085 : 4'b1001;
														assign node10085 = (inp[14]) ? 4'b0000 : 4'b0001;
													assign node10088 = (inp[7]) ? node10090 : 4'b1101;
														assign node10090 = (inp[12]) ? 4'b1001 : node10091;
															assign node10091 = (inp[1]) ? 4'b0101 : 4'b1001;
									assign node10095 = (inp[4]) ? node10161 : node10096;
										assign node10096 = (inp[3]) ? node10136 : node10097;
											assign node10097 = (inp[2]) ? node10107 : node10098;
												assign node10098 = (inp[12]) ? 4'b0001 : node10099;
													assign node10099 = (inp[1]) ? 4'b1001 : node10100;
														assign node10100 = (inp[14]) ? node10102 : 4'b0001;
															assign node10102 = (inp[13]) ? 4'b0001 : 4'b0100;
												assign node10107 = (inp[7]) ? node10123 : node10108;
													assign node10108 = (inp[12]) ? node10116 : node10109;
														assign node10109 = (inp[13]) ? node10113 : node10110;
															assign node10110 = (inp[1]) ? 4'b0000 : 4'b0001;
															assign node10113 = (inp[1]) ? 4'b1000 : 4'b1001;
														assign node10116 = (inp[13]) ? 4'b1000 : node10117;
															assign node10117 = (inp[14]) ? node10119 : 4'b1101;
																assign node10119 = (inp[1]) ? 4'b1101 : 4'b1100;
													assign node10123 = (inp[1]) ? node10127 : node10124;
														assign node10124 = (inp[14]) ? 4'b1100 : 4'b1101;
														assign node10127 = (inp[14]) ? node10131 : node10128;
															assign node10128 = (inp[12]) ? 4'b0100 : 4'b1100;
															assign node10131 = (inp[13]) ? node10133 : 4'b1101;
																assign node10133 = (inp[12]) ? 4'b0101 : 4'b1101;
											assign node10136 = (inp[1]) ? node10146 : node10137;
												assign node10137 = (inp[7]) ? node10139 : 4'b0001;
													assign node10139 = (inp[2]) ? node10141 : 4'b0101;
														assign node10141 = (inp[13]) ? 4'b0001 : node10142;
															assign node10142 = (inp[14]) ? 4'b0000 : 4'b0001;
												assign node10146 = (inp[12]) ? node10154 : node10147;
													assign node10147 = (inp[13]) ? 4'b1001 : node10148;
														assign node10148 = (inp[14]) ? node10150 : 4'b0000;
															assign node10150 = (inp[2]) ? 4'b1001 : 4'b1101;
													assign node10154 = (inp[14]) ? node10156 : 4'b0001;
														assign node10156 = (inp[2]) ? 4'b0001 : node10157;
															assign node10157 = (inp[13]) ? 4'b0000 : 4'b0001;
										assign node10161 = (inp[13]) ? node10209 : node10162;
											assign node10162 = (inp[7]) ? node10190 : node10163;
												assign node10163 = (inp[2]) ? node10175 : node10164;
													assign node10164 = (inp[3]) ? node10170 : node10165;
														assign node10165 = (inp[12]) ? 4'b0101 : node10166;
															assign node10166 = (inp[1]) ? 4'b1101 : 4'b0101;
														assign node10170 = (inp[12]) ? 4'b1001 : node10171;
															assign node10171 = (inp[14]) ? 4'b0100 : 4'b0101;
													assign node10175 = (inp[3]) ? node10185 : node10176;
														assign node10176 = (inp[12]) ? node10182 : node10177;
															assign node10177 = (inp[1]) ? 4'b0001 : node10178;
																assign node10178 = (inp[14]) ? 4'b0000 : 4'b0001;
															assign node10182 = (inp[14]) ? 4'b1000 : 4'b0000;
														assign node10185 = (inp[12]) ? 4'b0101 : node10186;
															assign node10186 = (inp[14]) ? 4'b0101 : 4'b1101;
												assign node10190 = (inp[2]) ? node10200 : node10191;
													assign node10191 = (inp[3]) ? node10195 : node10192;
														assign node10192 = (inp[14]) ? 4'b0001 : 4'b1001;
														assign node10195 = (inp[14]) ? 4'b1001 : node10196;
															assign node10196 = (inp[1]) ? 4'b1001 : 4'b1000;
													assign node10200 = (inp[3]) ? 4'b0001 : node10201;
														assign node10201 = (inp[14]) ? node10205 : node10202;
															assign node10202 = (inp[1]) ? 4'b0000 : 4'b0001;
															assign node10205 = (inp[1]) ? 4'b1101 : 4'b1100;
											assign node10209 = (inp[12]) ? node10225 : node10210;
												assign node10210 = (inp[1]) ? node10216 : node10211;
													assign node10211 = (inp[14]) ? 4'b0101 : node10212;
														assign node10212 = (inp[3]) ? 4'b0101 : 4'b1001;
													assign node10216 = (inp[3]) ? node10220 : node10217;
														assign node10217 = (inp[2]) ? 4'b1001 : 4'b1101;
														assign node10220 = (inp[14]) ? node10222 : 4'b1101;
															assign node10222 = (inp[2]) ? 4'b1101 : 4'b1100;
												assign node10225 = (inp[2]) ? node10237 : node10226;
													assign node10226 = (inp[3]) ? node10228 : 4'b0101;
														assign node10228 = (inp[14]) ? node10232 : node10229;
															assign node10229 = (inp[1]) ? 4'b0101 : 4'b0100;
															assign node10232 = (inp[1]) ? 4'b0100 : node10233;
																assign node10233 = (inp[7]) ? 4'b1001 : 4'b1101;
													assign node10237 = (inp[3]) ? 4'b0101 : node10238;
														assign node10238 = (inp[1]) ? 4'b0001 : node10239;
															assign node10239 = (inp[14]) ? 4'b0000 : 4'b0001;
								assign node10244 = (inp[1]) ? node10402 : node10245;
									assign node10245 = (inp[13]) ? node10317 : node10246;
										assign node10246 = (inp[3]) ? node10276 : node10247;
											assign node10247 = (inp[2]) ? node10263 : node10248;
												assign node10248 = (inp[4]) ? node10254 : node10249;
													assign node10249 = (inp[7]) ? node10251 : 4'b0000;
														assign node10251 = (inp[12]) ? 4'b1101 : 4'b0101;
													assign node10254 = (inp[7]) ? 4'b1000 : node10255;
														assign node10255 = (inp[10]) ? node10259 : node10256;
															assign node10256 = (inp[12]) ? 4'b1000 : 4'b0100;
															assign node10259 = (inp[12]) ? 4'b0100 : 4'b1100;
												assign node10263 = (inp[10]) ? node10269 : node10264;
													assign node10264 = (inp[4]) ? node10266 : 4'b1101;
														assign node10266 = (inp[7]) ? 4'b1101 : 4'b1001;
													assign node10269 = (inp[12]) ? node10271 : 4'b0001;
														assign node10271 = (inp[4]) ? node10273 : 4'b1101;
															assign node10273 = (inp[7]) ? 4'b1101 : 4'b1001;
											assign node10276 = (inp[4]) ? node10300 : node10277;
												assign node10277 = (inp[2]) ? node10289 : node10278;
													assign node10278 = (inp[7]) ? node10286 : node10279;
														assign node10279 = (inp[10]) ? node10283 : node10280;
															assign node10280 = (inp[12]) ? 4'b1100 : 4'b0000;
															assign node10283 = (inp[12]) ? 4'b0000 : 4'b1000;
														assign node10286 = (inp[12]) ? 4'b0100 : 4'b1100;
													assign node10289 = (inp[7]) ? node10297 : node10290;
														assign node10290 = (inp[12]) ? node10294 : node10291;
															assign node10291 = (inp[10]) ? 4'b1000 : 4'b0000;
															assign node10294 = (inp[10]) ? 4'b0000 : 4'b1001;
														assign node10297 = (inp[10]) ? 4'b0001 : 4'b1001;
												assign node10300 = (inp[2]) ? node10308 : node10301;
													assign node10301 = (inp[10]) ? 4'b1001 : node10302;
														assign node10302 = (inp[12]) ? node10304 : 4'b0001;
															assign node10304 = (inp[7]) ? 4'b1000 : 4'b1001;
													assign node10308 = (inp[7]) ? node10314 : node10309;
														assign node10309 = (inp[10]) ? node10311 : 4'b0100;
															assign node10311 = (inp[12]) ? 4'b0100 : 4'b1100;
														assign node10314 = (inp[10]) ? 4'b1000 : 4'b0000;
										assign node10317 = (inp[4]) ? node10363 : node10318;
											assign node10318 = (inp[2]) ? node10344 : node10319;
												assign node10319 = (inp[14]) ? node10333 : node10320;
													assign node10320 = (inp[3]) ? node10330 : node10321;
														assign node10321 = (inp[7]) ? 4'b0000 : node10322;
															assign node10322 = (inp[10]) ? node10326 : node10323;
																assign node10323 = (inp[12]) ? 4'b1000 : 4'b0000;
																assign node10326 = (inp[12]) ? 4'b0000 : 4'b1000;
														assign node10330 = (inp[10]) ? 4'b0001 : 4'b0000;
													assign node10333 = (inp[10]) ? node10337 : node10334;
														assign node10334 = (inp[7]) ? 4'b1100 : 4'b1000;
														assign node10337 = (inp[12]) ? 4'b0000 : node10338;
															assign node10338 = (inp[7]) ? 4'b1000 : node10339;
																assign node10339 = (inp[3]) ? 4'b0001 : 4'b1000;
												assign node10344 = (inp[3]) ? node10354 : node10345;
													assign node10345 = (inp[7]) ? node10349 : node10346;
														assign node10346 = (inp[10]) ? 4'b1001 : 4'b0001;
														assign node10349 = (inp[12]) ? 4'b0101 : node10350;
															assign node10350 = (inp[10]) ? 4'b1101 : 4'b0101;
													assign node10354 = (inp[7]) ? node10360 : node10355;
														assign node10355 = (inp[10]) ? 4'b0000 : node10356;
															assign node10356 = (inp[12]) ? 4'b1000 : 4'b0000;
														assign node10360 = (inp[12]) ? 4'b0001 : 4'b0000;
											assign node10363 = (inp[12]) ? node10383 : node10364;
												assign node10364 = (inp[10]) ? node10376 : node10365;
													assign node10365 = (inp[7]) ? node10371 : node10366;
														assign node10366 = (inp[2]) ? 4'b0100 : node10367;
															assign node10367 = (inp[3]) ? 4'b1101 : 4'b0100;
														assign node10371 = (inp[2]) ? node10373 : 4'b1001;
															assign node10373 = (inp[3]) ? 4'b0100 : 4'b0001;
													assign node10376 = (inp[3]) ? node10380 : node10377;
														assign node10377 = (inp[2]) ? 4'b1001 : 4'b1100;
														assign node10380 = (inp[2]) ? 4'b1100 : 4'b0101;
												assign node10383 = (inp[10]) ? node10391 : node10384;
													assign node10384 = (inp[7]) ? 4'b0001 : node10385;
														assign node10385 = (inp[2]) ? node10387 : 4'b1100;
															assign node10387 = (inp[3]) ? 4'b1100 : 4'b0001;
													assign node10391 = (inp[14]) ? node10397 : node10392;
														assign node10392 = (inp[2]) ? 4'b0001 : node10393;
															assign node10393 = (inp[3]) ? 4'b0101 : 4'b0100;
														assign node10397 = (inp[3]) ? node10399 : 4'b0100;
															assign node10399 = (inp[2]) ? 4'b0100 : 4'b0101;
									assign node10402 = (inp[10]) ? node10474 : node10403;
										assign node10403 = (inp[4]) ? node10427 : node10404;
											assign node10404 = (inp[2]) ? node10410 : node10405;
												assign node10405 = (inp[7]) ? node10407 : 4'b0000;
													assign node10407 = (inp[13]) ? 4'b0000 : 4'b1100;
												assign node10410 = (inp[3]) ? node10422 : node10411;
													assign node10411 = (inp[7]) ? node10419 : node10412;
														assign node10412 = (inp[14]) ? 4'b1000 : node10413;
															assign node10413 = (inp[12]) ? node10415 : 4'b0000;
																assign node10415 = (inp[13]) ? 4'b0000 : 4'b1100;
														assign node10419 = (inp[12]) ? 4'b0100 : 4'b1100;
													assign node10422 = (inp[13]) ? 4'b0000 : node10423;
														assign node10423 = (inp[7]) ? 4'b1000 : 4'b0000;
											assign node10427 = (inp[7]) ? node10455 : node10428;
												assign node10428 = (inp[14]) ? node10438 : node10429;
													assign node10429 = (inp[12]) ? node10431 : 4'b0100;
														assign node10431 = (inp[3]) ? node10435 : node10432;
															assign node10432 = (inp[2]) ? 4'b0000 : 4'b0100;
															assign node10435 = (inp[2]) ? 4'b0100 : 4'b0000;
													assign node10438 = (inp[2]) ? node10448 : node10439;
														assign node10439 = (inp[3]) ? node10441 : 4'b0100;
															assign node10441 = (inp[13]) ? node10445 : node10442;
																assign node10442 = (inp[12]) ? 4'b0000 : 4'b1000;
																assign node10445 = (inp[12]) ? 4'b1100 : 4'b0100;
														assign node10448 = (inp[3]) ? 4'b0100 : node10449;
															assign node10449 = (inp[13]) ? node10451 : 4'b1000;
																assign node10451 = (inp[12]) ? 4'b0000 : 4'b1000;
												assign node10455 = (inp[13]) ? node10463 : node10456;
													assign node10456 = (inp[3]) ? 4'b0000 : node10457;
														assign node10457 = (inp[14]) ? 4'b0000 : node10458;
															assign node10458 = (inp[2]) ? 4'b1100 : 4'b0000;
													assign node10463 = (inp[3]) ? node10469 : node10464;
														assign node10464 = (inp[2]) ? node10466 : 4'b0100;
															assign node10466 = (inp[12]) ? 4'b0000 : 4'b1000;
														assign node10469 = (inp[2]) ? 4'b0100 : node10470;
															assign node10470 = (inp[12]) ? 4'b1000 : 4'b0100;
										assign node10474 = (inp[13]) ? node10506 : node10475;
											assign node10475 = (inp[2]) ? node10497 : node10476;
												assign node10476 = (inp[12]) ? node10484 : node10477;
													assign node10477 = (inp[14]) ? node10479 : 4'b0100;
														assign node10479 = (inp[3]) ? node10481 : 4'b1000;
															assign node10481 = (inp[7]) ? 4'b0000 : 4'b0100;
													assign node10484 = (inp[7]) ? node10490 : node10485;
														assign node10485 = (inp[4]) ? node10487 : 4'b1000;
															assign node10487 = (inp[3]) ? 4'b0100 : 4'b1100;
														assign node10490 = (inp[4]) ? node10494 : node10491;
															assign node10491 = (inp[3]) ? 4'b1100 : 4'b0100;
															assign node10494 = (inp[3]) ? 4'b0000 : 4'b1000;
												assign node10497 = (inp[3]) ? node10501 : node10498;
													assign node10498 = (inp[7]) ? 4'b0100 : 4'b0000;
													assign node10501 = (inp[4]) ? 4'b1000 : node10502;
														assign node10502 = (inp[7]) ? 4'b0000 : 4'b1000;
											assign node10506 = (inp[4]) ? node10514 : node10507;
												assign node10507 = (inp[7]) ? node10509 : 4'b1000;
													assign node10509 = (inp[2]) ? node10511 : 4'b1000;
														assign node10511 = (inp[12]) ? 4'b1100 : 4'b1000;
												assign node10514 = (inp[2]) ? node10516 : 4'b1100;
													assign node10516 = (inp[3]) ? 4'b1100 : 4'b1000;
							assign node10519 = (inp[2]) ? 4'b1100 : node10520;
								assign node10520 = (inp[3]) ? node10634 : node10521;
									assign node10521 = (inp[4]) ? node10551 : node10522;
										assign node10522 = (inp[7]) ? 4'b1100 : node10523;
											assign node10523 = (inp[13]) ? node10535 : node10524;
												assign node10524 = (inp[10]) ? node10530 : node10525;
													assign node10525 = (inp[1]) ? node10527 : 4'b1100;
														assign node10527 = (inp[12]) ? 4'b1100 : 4'b0000;
													assign node10530 = (inp[12]) ? node10532 : 4'b0001;
														assign node10532 = (inp[14]) ? 4'b1100 : 4'b0000;
												assign node10535 = (inp[12]) ? node10541 : node10536;
													assign node10536 = (inp[1]) ? 4'b1000 : node10537;
														assign node10537 = (inp[10]) ? 4'b1001 : 4'b0001;
													assign node10541 = (inp[10]) ? node10547 : node10542;
														assign node10542 = (inp[14]) ? node10544 : 4'b0000;
															assign node10544 = (inp[1]) ? 4'b0001 : 4'b0000;
														assign node10547 = (inp[14]) ? 4'b0000 : 4'b0001;
										assign node10551 = (inp[13]) ? node10603 : node10552;
											assign node10552 = (inp[7]) ? node10588 : node10553;
												assign node10553 = (inp[12]) ? node10573 : node10554;
													assign node10554 = (inp[10]) ? node10564 : node10555;
														assign node10555 = (inp[14]) ? node10557 : 4'b0000;
															assign node10557 = (inp[11]) ? node10561 : node10558;
																assign node10558 = (inp[1]) ? 4'b1001 : 4'b1000;
																assign node10561 = (inp[1]) ? 4'b0000 : 4'b1001;
														assign node10564 = (inp[14]) ? node10568 : node10565;
															assign node10565 = (inp[1]) ? 4'b0000 : 4'b0001;
															assign node10568 = (inp[1]) ? node10570 : 4'b0000;
																assign node10570 = (inp[11]) ? 4'b0000 : 4'b0001;
													assign node10573 = (inp[11]) ? node10583 : node10574;
														assign node10574 = (inp[10]) ? node10578 : node10575;
															assign node10575 = (inp[14]) ? 4'b1001 : 4'b1000;
															assign node10578 = (inp[1]) ? 4'b1001 : node10579;
																assign node10579 = (inp[14]) ? 4'b1000 : 4'b1001;
														assign node10583 = (inp[10]) ? 4'b0000 : node10584;
															assign node10584 = (inp[1]) ? 4'b1000 : 4'b1001;
												assign node10588 = (inp[12]) ? node10596 : node10589;
													assign node10589 = (inp[10]) ? node10591 : 4'b1100;
														assign node10591 = (inp[1]) ? node10593 : 4'b0001;
															assign node10593 = (inp[14]) ? 4'b0001 : 4'b0000;
													assign node10596 = (inp[1]) ? node10598 : 4'b1100;
														assign node10598 = (inp[14]) ? node10600 : 4'b1100;
															assign node10600 = (inp[11]) ? 4'b0000 : 4'b1100;
											assign node10603 = (inp[10]) ? node10619 : node10604;
												assign node10604 = (inp[1]) ? node10610 : node10605;
													assign node10605 = (inp[11]) ? 4'b0001 : node10606;
														assign node10606 = (inp[14]) ? 4'b0000 : 4'b0001;
													assign node10610 = (inp[14]) ? node10614 : node10611;
														assign node10611 = (inp[12]) ? 4'b0000 : 4'b1000;
														assign node10614 = (inp[11]) ? node10616 : 4'b0001;
															assign node10616 = (inp[12]) ? 4'b0000 : 4'b1000;
												assign node10619 = (inp[1]) ? node10629 : node10620;
													assign node10620 = (inp[12]) ? node10626 : node10621;
														assign node10621 = (inp[11]) ? 4'b1001 : node10622;
															assign node10622 = (inp[14]) ? 4'b1000 : 4'b1001;
														assign node10626 = (inp[11]) ? 4'b0001 : 4'b0000;
													assign node10629 = (inp[14]) ? node10631 : 4'b1000;
														assign node10631 = (inp[12]) ? 4'b0001 : 4'b1001;
									assign node10634 = (inp[4]) ? node10714 : node10635;
										assign node10635 = (inp[7]) ? node10679 : node10636;
											assign node10636 = (inp[13]) ? node10660 : node10637;
												assign node10637 = (inp[12]) ? node10651 : node10638;
													assign node10638 = (inp[1]) ? node10646 : node10639;
														assign node10639 = (inp[10]) ? node10643 : node10640;
															assign node10640 = (inp[11]) ? 4'b1001 : 4'b1000;
															assign node10643 = (inp[11]) ? 4'b0101 : 4'b0100;
														assign node10646 = (inp[11]) ? 4'b0100 : node10647;
															assign node10647 = (inp[10]) ? 4'b0101 : 4'b0100;
													assign node10651 = (inp[10]) ? node10653 : 4'b1000;
														assign node10653 = (inp[11]) ? 4'b1001 : node10654;
															assign node10654 = (inp[14]) ? node10656 : 4'b0100;
																assign node10656 = (inp[1]) ? 4'b1001 : 4'b1000;
												assign node10660 = (inp[12]) ? node10674 : node10661;
													assign node10661 = (inp[11]) ? node10671 : node10662;
														assign node10662 = (inp[10]) ? 4'b1100 : node10663;
															assign node10663 = (inp[1]) ? node10667 : node10664;
																assign node10664 = (inp[14]) ? 4'b0100 : 4'b0101;
																assign node10667 = (inp[14]) ? 4'b0101 : 4'b1100;
														assign node10671 = (inp[1]) ? 4'b1100 : 4'b1101;
													assign node10674 = (inp[1]) ? node10676 : 4'b0101;
														assign node10676 = (inp[14]) ? 4'b0101 : 4'b1100;
											assign node10679 = (inp[1]) ? node10697 : node10680;
												assign node10680 = (inp[11]) ? node10690 : node10681;
													assign node10681 = (inp[10]) ? node10683 : 4'b0000;
														assign node10683 = (inp[13]) ? node10687 : node10684;
															assign node10684 = (inp[12]) ? 4'b1000 : 4'b0000;
															assign node10687 = (inp[12]) ? 4'b0000 : 4'b1000;
													assign node10690 = (inp[13]) ? node10692 : 4'b1001;
														assign node10692 = (inp[10]) ? node10694 : 4'b0001;
															assign node10694 = (inp[12]) ? 4'b0001 : 4'b1001;
												assign node10697 = (inp[14]) ? node10709 : node10698;
													assign node10698 = (inp[13]) ? node10704 : node10699;
														assign node10699 = (inp[10]) ? 4'b0000 : node10700;
															assign node10700 = (inp[12]) ? 4'b1000 : 4'b0000;
														assign node10704 = (inp[10]) ? 4'b1000 : node10705;
															assign node10705 = (inp[12]) ? 4'b0000 : 4'b1000;
													assign node10709 = (inp[13]) ? 4'b0001 : node10710;
														assign node10710 = (inp[11]) ? 4'b1000 : 4'b1001;
										assign node10714 = (inp[1]) ? node10742 : node10715;
											assign node10715 = (inp[11]) ? node10729 : node10716;
												assign node10716 = (inp[14]) ? node10724 : node10717;
													assign node10717 = (inp[12]) ? 4'b0101 : node10718;
														assign node10718 = (inp[13]) ? 4'b1101 : node10719;
															assign node10719 = (inp[10]) ? 4'b0101 : 4'b1101;
													assign node10724 = (inp[10]) ? node10726 : 4'b0100;
														assign node10726 = (inp[13]) ? 4'b1100 : 4'b0100;
												assign node10729 = (inp[13]) ? node10737 : node10730;
													assign node10730 = (inp[10]) ? node10734 : node10731;
														assign node10731 = (inp[7]) ? 4'b1001 : 4'b1101;
														assign node10734 = (inp[14]) ? 4'b1101 : 4'b0101;
													assign node10737 = (inp[12]) ? 4'b0101 : node10738;
														assign node10738 = (inp[10]) ? 4'b1101 : 4'b0101;
											assign node10742 = (inp[11]) ? node10762 : node10743;
												assign node10743 = (inp[14]) ? node10751 : node10744;
													assign node10744 = (inp[10]) ? 4'b0100 : node10745;
														assign node10745 = (inp[12]) ? node10747 : 4'b0100;
															assign node10747 = (inp[7]) ? 4'b1000 : 4'b1100;
													assign node10751 = (inp[13]) ? node10757 : node10752;
														assign node10752 = (inp[10]) ? node10754 : 4'b1001;
															assign node10754 = (inp[12]) ? 4'b1101 : 4'b0101;
														assign node10757 = (inp[12]) ? 4'b0101 : node10758;
															assign node10758 = (inp[7]) ? 4'b0101 : 4'b1101;
												assign node10762 = (inp[13]) ? node10770 : node10763;
													assign node10763 = (inp[12]) ? node10765 : 4'b0100;
														assign node10765 = (inp[10]) ? 4'b0100 : node10766;
															assign node10766 = (inp[7]) ? 4'b1000 : 4'b1100;
													assign node10770 = (inp[10]) ? 4'b1100 : node10771;
														assign node10771 = (inp[12]) ? 4'b0100 : 4'b1100;
						assign node10776 = (inp[3]) ? node11396 : node10777;
							assign node10777 = (inp[1]) ? node11105 : node10778;
								assign node10778 = (inp[13]) ? node10932 : node10779;
									assign node10779 = (inp[4]) ? node10855 : node10780;
										assign node10780 = (inp[7]) ? node10828 : node10781;
											assign node10781 = (inp[10]) ? node10805 : node10782;
												assign node10782 = (inp[11]) ? node10794 : node10783;
													assign node10783 = (inp[0]) ? node10789 : node10784;
														assign node10784 = (inp[14]) ? 4'b1101 : node10785;
															assign node10785 = (inp[2]) ? 4'b1101 : 4'b1100;
														assign node10789 = (inp[2]) ? 4'b1100 : node10790;
															assign node10790 = (inp[14]) ? 4'b1100 : 4'b1101;
													assign node10794 = (inp[0]) ? node10802 : node10795;
														assign node10795 = (inp[12]) ? node10799 : node10796;
															assign node10796 = (inp[2]) ? 4'b0001 : 4'b0000;
															assign node10799 = (inp[2]) ? 4'b1100 : 4'b0000;
														assign node10802 = (inp[2]) ? 4'b1100 : 4'b1101;
												assign node10805 = (inp[2]) ? node10813 : node10806;
													assign node10806 = (inp[12]) ? node10810 : node10807;
														assign node10807 = (inp[11]) ? 4'b1000 : 4'b0000;
														assign node10810 = (inp[14]) ? 4'b0001 : 4'b0000;
													assign node10813 = (inp[12]) ? node10823 : node10814;
														assign node10814 = (inp[0]) ? node10818 : node10815;
															assign node10815 = (inp[11]) ? 4'b1001 : 4'b1000;
															assign node10818 = (inp[14]) ? node10820 : 4'b0001;
																assign node10820 = (inp[11]) ? 4'b0001 : 4'b0000;
														assign node10823 = (inp[0]) ? 4'b1100 : node10824;
															assign node10824 = (inp[14]) ? 4'b1001 : 4'b1000;
											assign node10828 = (inp[0]) ? node10848 : node10829;
												assign node10829 = (inp[10]) ? node10841 : node10830;
													assign node10830 = (inp[14]) ? node10838 : node10831;
														assign node10831 = (inp[12]) ? 4'b1101 : node10832;
															assign node10832 = (inp[2]) ? 4'b1101 : node10833;
																assign node10833 = (inp[11]) ? 4'b0101 : 4'b0100;
														assign node10838 = (inp[12]) ? 4'b1100 : 4'b0100;
													assign node10841 = (inp[2]) ? node10843 : 4'b0000;
														assign node10843 = (inp[11]) ? node10845 : 4'b0101;
															assign node10845 = (inp[14]) ? 4'b0100 : 4'b1100;
												assign node10848 = (inp[2]) ? 4'b1100 : node10849;
													assign node10849 = (inp[10]) ? 4'b0101 : node10850;
														assign node10850 = (inp[14]) ? 4'b1100 : 4'b1101;
										assign node10855 = (inp[2]) ? node10897 : node10856;
											assign node10856 = (inp[7]) ? node10878 : node10857;
												assign node10857 = (inp[10]) ? node10869 : node10858;
													assign node10858 = (inp[0]) ? node10864 : node10859;
														assign node10859 = (inp[11]) ? 4'b0001 : node10860;
															assign node10860 = (inp[14]) ? 4'b1000 : 4'b0001;
														assign node10864 = (inp[11]) ? node10866 : 4'b1001;
															assign node10866 = (inp[12]) ? 4'b1000 : 4'b0100;
													assign node10869 = (inp[11]) ? node10871 : 4'b0101;
														assign node10871 = (inp[12]) ? node10875 : node10872;
															assign node10872 = (inp[0]) ? 4'b1100 : 4'b0000;
															assign node10875 = (inp[0]) ? 4'b0100 : 4'b0101;
												assign node10878 = (inp[11]) ? node10886 : node10879;
													assign node10879 = (inp[0]) ? node10883 : node10880;
														assign node10880 = (inp[12]) ? 4'b1100 : 4'b0000;
														assign node10883 = (inp[10]) ? 4'b0001 : 4'b1001;
													assign node10886 = (inp[0]) ? node10892 : node10887;
														assign node10887 = (inp[12]) ? 4'b0001 : node10888;
															assign node10888 = (inp[10]) ? 4'b1001 : 4'b0001;
														assign node10892 = (inp[12]) ? 4'b0000 : node10893;
															assign node10893 = (inp[10]) ? 4'b1000 : 4'b0000;
											assign node10897 = (inp[12]) ? node10915 : node10898;
												assign node10898 = (inp[10]) ? node10910 : node10899;
													assign node10899 = (inp[0]) ? node10907 : node10900;
														assign node10900 = (inp[7]) ? node10902 : 4'b0000;
															assign node10902 = (inp[14]) ? 4'b1001 : node10903;
																assign node10903 = (inp[11]) ? 4'b0101 : 4'b0100;
														assign node10907 = (inp[7]) ? 4'b1100 : 4'b1001;
													assign node10910 = (inp[0]) ? node10912 : 4'b0000;
														assign node10912 = (inp[11]) ? 4'b0001 : 4'b0000;
												assign node10915 = (inp[7]) ? node10925 : node10916;
													assign node10916 = (inp[0]) ? node10922 : node10917;
														assign node10917 = (inp[10]) ? 4'b0000 : node10918;
															assign node10918 = (inp[14]) ? 4'b1101 : 4'b1100;
														assign node10922 = (inp[14]) ? 4'b1000 : 4'b1001;
													assign node10925 = (inp[0]) ? 4'b1100 : node10926;
														assign node10926 = (inp[14]) ? 4'b1001 : node10927;
															assign node10927 = (inp[10]) ? 4'b1100 : 4'b1000;
									assign node10932 = (inp[0]) ? node11024 : node10933;
										assign node10933 = (inp[11]) ? node10985 : node10934;
											assign node10934 = (inp[12]) ? node10958 : node10935;
												assign node10935 = (inp[4]) ? node10945 : node10936;
													assign node10936 = (inp[2]) ? node10938 : 4'b0100;
														assign node10938 = (inp[14]) ? node10942 : node10939;
															assign node10939 = (inp[7]) ? 4'b0000 : 4'b1000;
															assign node10942 = (inp[10]) ? 4'b0101 : 4'b0001;
													assign node10945 = (inp[2]) ? node10953 : node10946;
														assign node10946 = (inp[10]) ? node10948 : 4'b0001;
															assign node10948 = (inp[14]) ? node10950 : 4'b1000;
																assign node10950 = (inp[7]) ? 4'b1001 : 4'b0001;
														assign node10953 = (inp[10]) ? 4'b1000 : node10954;
															assign node10954 = (inp[7]) ? 4'b0000 : 4'b0100;
												assign node10958 = (inp[7]) ? node10980 : node10959;
													assign node10959 = (inp[14]) ? node10971 : node10960;
														assign node10960 = (inp[10]) ? node10968 : node10961;
															assign node10961 = (inp[2]) ? node10965 : node10962;
																assign node10962 = (inp[4]) ? 4'b1001 : 4'b1000;
																assign node10965 = (inp[4]) ? 4'b1000 : 4'b0000;
															assign node10968 = (inp[2]) ? 4'b0100 : 4'b1100;
														assign node10971 = (inp[10]) ? node10975 : node10972;
															assign node10972 = (inp[2]) ? 4'b0001 : 4'b1001;
															assign node10975 = (inp[2]) ? node10977 : 4'b0001;
																assign node10977 = (inp[4]) ? 4'b1000 : 4'b1001;
													assign node10980 = (inp[4]) ? node10982 : 4'b1000;
														assign node10982 = (inp[14]) ? 4'b0100 : 4'b1000;
											assign node10985 = (inp[2]) ? node11005 : node10986;
												assign node10986 = (inp[4]) ? node10996 : node10987;
													assign node10987 = (inp[7]) ? node10993 : node10988;
														assign node10988 = (inp[12]) ? 4'b0100 : node10989;
															assign node10989 = (inp[10]) ? 4'b0001 : 4'b0100;
														assign node10993 = (inp[10]) ? 4'b0100 : 4'b0000;
													assign node10996 = (inp[10]) ? node11000 : node10997;
														assign node10997 = (inp[12]) ? 4'b0000 : 4'b1000;
														assign node11000 = (inp[7]) ? node11002 : 4'b1001;
															assign node11002 = (inp[14]) ? 4'b1000 : 4'b0100;
												assign node11005 = (inp[4]) ? node11013 : node11006;
													assign node11006 = (inp[10]) ? node11010 : node11007;
														assign node11007 = (inp[12]) ? 4'b0001 : 4'b1001;
														assign node11010 = (inp[7]) ? 4'b0001 : 4'b0101;
													assign node11013 = (inp[12]) ? node11019 : node11014;
														assign node11014 = (inp[10]) ? 4'b0001 : node11015;
															assign node11015 = (inp[7]) ? 4'b0000 : 4'b0100;
														assign node11019 = (inp[10]) ? 4'b0100 : node11020;
															assign node11020 = (inp[7]) ? 4'b0000 : 4'b0100;
										assign node11024 = (inp[12]) ? node11064 : node11025;
											assign node11025 = (inp[10]) ? node11049 : node11026;
												assign node11026 = (inp[7]) ? node11038 : node11027;
													assign node11027 = (inp[2]) ? node11033 : node11028;
														assign node11028 = (inp[11]) ? 4'b0000 : node11029;
															assign node11029 = (inp[4]) ? 4'b1000 : 4'b1001;
														assign node11033 = (inp[14]) ? node11035 : 4'b0001;
															assign node11035 = (inp[4]) ? 4'b0000 : 4'b0001;
													assign node11038 = (inp[4]) ? node11046 : node11039;
														assign node11039 = (inp[2]) ? 4'b1100 : node11040;
															assign node11040 = (inp[14]) ? node11042 : 4'b0101;
																assign node11042 = (inp[11]) ? 4'b0000 : 4'b0100;
														assign node11046 = (inp[2]) ? 4'b0001 : 4'b1001;
												assign node11049 = (inp[2]) ? node11055 : node11050;
													assign node11050 = (inp[11]) ? node11052 : 4'b0001;
														assign node11052 = (inp[4]) ? 4'b0001 : 4'b1000;
													assign node11055 = (inp[4]) ? node11059 : node11056;
														assign node11056 = (inp[7]) ? 4'b1100 : 4'b1001;
														assign node11059 = (inp[11]) ? 4'b1001 : node11060;
															assign node11060 = (inp[14]) ? 4'b1000 : 4'b1001;
											assign node11064 = (inp[10]) ? node11086 : node11065;
												assign node11065 = (inp[2]) ? node11079 : node11066;
													assign node11066 = (inp[4]) ? node11072 : node11067;
														assign node11067 = (inp[7]) ? 4'b0101 : node11068;
															assign node11068 = (inp[11]) ? 4'b1000 : 4'b1001;
														assign node11072 = (inp[7]) ? node11076 : node11073;
															assign node11073 = (inp[11]) ? 4'b0001 : 4'b0000;
															assign node11076 = (inp[11]) ? 4'b1000 : 4'b1001;
													assign node11079 = (inp[7]) ? node11083 : node11080;
														assign node11080 = (inp[14]) ? 4'b0000 : 4'b0001;
														assign node11083 = (inp[4]) ? 4'b0000 : 4'b1100;
												assign node11086 = (inp[2]) ? 4'b0001 : node11087;
													assign node11087 = (inp[7]) ? node11097 : node11088;
														assign node11088 = (inp[14]) ? node11092 : node11089;
															assign node11089 = (inp[11]) ? 4'b0001 : 4'b0000;
															assign node11092 = (inp[4]) ? node11094 : 4'b0001;
																assign node11094 = (inp[11]) ? 4'b0001 : 4'b1001;
														assign node11097 = (inp[11]) ? node11101 : node11098;
															assign node11098 = (inp[4]) ? 4'b0000 : 4'b0001;
															assign node11101 = (inp[4]) ? 4'b0001 : 4'b0000;
								assign node11105 = (inp[11]) ? node11279 : node11106;
									assign node11106 = (inp[4]) ? node11194 : node11107;
										assign node11107 = (inp[7]) ? node11165 : node11108;
											assign node11108 = (inp[0]) ? node11146 : node11109;
												assign node11109 = (inp[14]) ? node11123 : node11110;
													assign node11110 = (inp[2]) ? node11114 : node11111;
														assign node11111 = (inp[12]) ? 4'b0000 : 4'b1000;
														assign node11114 = (inp[13]) ? node11120 : node11115;
															assign node11115 = (inp[10]) ? node11117 : 4'b0001;
																assign node11117 = (inp[12]) ? 4'b1001 : 4'b0001;
															assign node11120 = (inp[10]) ? 4'b1101 : 4'b1001;
													assign node11123 = (inp[12]) ? node11133 : node11124;
														assign node11124 = (inp[10]) ? node11130 : node11125;
															assign node11125 = (inp[13]) ? 4'b1000 : node11126;
																assign node11126 = (inp[2]) ? 4'b0000 : 4'b1000;
															assign node11130 = (inp[13]) ? 4'b1100 : 4'b1000;
														assign node11133 = (inp[2]) ? node11139 : node11134;
															assign node11134 = (inp[10]) ? 4'b0001 : node11135;
																assign node11135 = (inp[13]) ? 4'b0100 : 4'b0000;
															assign node11139 = (inp[10]) ? node11143 : node11140;
																assign node11140 = (inp[13]) ? 4'b1000 : 4'b0000;
																assign node11143 = (inp[13]) ? 4'b0100 : 4'b1000;
												assign node11146 = (inp[2]) ? node11154 : node11147;
													assign node11147 = (inp[12]) ? node11151 : node11148;
														assign node11148 = (inp[10]) ? 4'b1001 : 4'b0001;
														assign node11151 = (inp[10]) ? 4'b0001 : 4'b1101;
													assign node11154 = (inp[14]) ? node11160 : node11155;
														assign node11155 = (inp[12]) ? 4'b0000 : node11156;
															assign node11156 = (inp[13]) ? 4'b1000 : 4'b0000;
														assign node11160 = (inp[12]) ? 4'b0001 : node11161;
															assign node11161 = (inp[13]) ? 4'b1001 : 4'b0001;
											assign node11165 = (inp[2]) ? node11189 : node11166;
												assign node11166 = (inp[0]) ? node11178 : node11167;
													assign node11167 = (inp[12]) ? node11173 : node11168;
														assign node11168 = (inp[13]) ? node11170 : 4'b0100;
															assign node11170 = (inp[10]) ? 4'b1100 : 4'b1000;
														assign node11173 = (inp[10]) ? 4'b0100 : node11174;
															assign node11174 = (inp[13]) ? 4'b0000 : 4'b0100;
													assign node11178 = (inp[13]) ? node11184 : node11179;
														assign node11179 = (inp[14]) ? node11181 : 4'b0100;
															assign node11181 = (inp[10]) ? 4'b0101 : 4'b1101;
														assign node11184 = (inp[14]) ? 4'b0001 : node11185;
															assign node11185 = (inp[10]) ? 4'b1001 : 4'b0001;
												assign node11189 = (inp[0]) ? 4'b1100 : node11190;
													assign node11190 = (inp[14]) ? 4'b1000 : 4'b1001;
										assign node11194 = (inp[2]) ? node11244 : node11195;
											assign node11195 = (inp[10]) ? node11223 : node11196;
												assign node11196 = (inp[12]) ? node11210 : node11197;
													assign node11197 = (inp[0]) ? node11203 : node11198;
														assign node11198 = (inp[14]) ? 4'b1001 : node11199;
															assign node11199 = (inp[13]) ? 4'b1001 : 4'b1000;
														assign node11203 = (inp[14]) ? 4'b0001 : node11204;
															assign node11204 = (inp[13]) ? node11206 : 4'b0101;
																assign node11206 = (inp[7]) ? 4'b0101 : 4'b1001;
													assign node11210 = (inp[7]) ? 4'b1001 : node11211;
														assign node11211 = (inp[14]) ? node11217 : node11212;
															assign node11212 = (inp[0]) ? 4'b1001 : node11213;
																assign node11213 = (inp[13]) ? 4'b1001 : 4'b1000;
															assign node11217 = (inp[0]) ? node11219 : 4'b1001;
																assign node11219 = (inp[13]) ? 4'b1000 : 4'b1001;
												assign node11223 = (inp[14]) ? node11229 : node11224;
													assign node11224 = (inp[12]) ? 4'b0001 : node11225;
														assign node11225 = (inp[13]) ? 4'b1001 : 4'b0001;
													assign node11229 = (inp[13]) ? node11241 : node11230;
														assign node11230 = (inp[7]) ? node11236 : node11231;
															assign node11231 = (inp[12]) ? 4'b0101 : node11232;
																assign node11232 = (inp[0]) ? 4'b0000 : 4'b0001;
															assign node11236 = (inp[12]) ? node11238 : 4'b1001;
																assign node11238 = (inp[0]) ? 4'b0001 : 4'b1001;
														assign node11241 = (inp[12]) ? 4'b0000 : 4'b1000;
											assign node11244 = (inp[14]) ? node11260 : node11245;
												assign node11245 = (inp[13]) ? node11255 : node11246;
													assign node11246 = (inp[10]) ? 4'b0000 : node11247;
														assign node11247 = (inp[7]) ? node11251 : node11248;
															assign node11248 = (inp[12]) ? 4'b0000 : 4'b1000;
															assign node11251 = (inp[0]) ? 4'b1100 : 4'b0101;
													assign node11255 = (inp[12]) ? node11257 : 4'b1000;
														assign node11257 = (inp[0]) ? 4'b1000 : 4'b0000;
												assign node11260 = (inp[0]) ? node11268 : node11261;
													assign node11261 = (inp[13]) ? node11263 : 4'b1000;
														assign node11263 = (inp[10]) ? 4'b0001 : node11264;
															assign node11264 = (inp[12]) ? 4'b0000 : 4'b1000;
													assign node11268 = (inp[10]) ? node11274 : node11269;
														assign node11269 = (inp[13]) ? 4'b0001 : node11270;
															assign node11270 = (inp[7]) ? 4'b1100 : 4'b1001;
														assign node11274 = (inp[13]) ? node11276 : 4'b0001;
															assign node11276 = (inp[12]) ? 4'b0001 : 4'b1001;
									assign node11279 = (inp[10]) ? node11349 : node11280;
										assign node11280 = (inp[2]) ? node11308 : node11281;
											assign node11281 = (inp[0]) ? node11295 : node11282;
												assign node11282 = (inp[4]) ? node11290 : node11283;
													assign node11283 = (inp[12]) ? node11287 : node11284;
														assign node11284 = (inp[14]) ? 4'b1100 : 4'b1000;
														assign node11287 = (inp[13]) ? 4'b1100 : 4'b0100;
													assign node11290 = (inp[12]) ? 4'b1000 : node11291;
														assign node11291 = (inp[13]) ? 4'b0000 : 4'b0100;
												assign node11295 = (inp[13]) ? 4'b0000 : node11296;
													assign node11296 = (inp[14]) ? node11302 : node11297;
														assign node11297 = (inp[4]) ? 4'b0100 : node11298;
															assign node11298 = (inp[7]) ? 4'b0100 : 4'b0000;
														assign node11302 = (inp[4]) ? 4'b0000 : node11303;
															assign node11303 = (inp[7]) ? 4'b0100 : 4'b0000;
											assign node11308 = (inp[7]) ? node11334 : node11309;
												assign node11309 = (inp[4]) ? node11323 : node11310;
													assign node11310 = (inp[14]) ? node11316 : node11311;
														assign node11311 = (inp[12]) ? 4'b0000 : node11312;
															assign node11312 = (inp[0]) ? 4'b1000 : 4'b0100;
														assign node11316 = (inp[0]) ? node11318 : 4'b1000;
															assign node11318 = (inp[13]) ? 4'b0000 : node11319;
																assign node11319 = (inp[12]) ? 4'b1100 : 4'b0000;
													assign node11323 = (inp[0]) ? node11329 : node11324;
														assign node11324 = (inp[14]) ? node11326 : 4'b1000;
															assign node11326 = (inp[13]) ? 4'b0000 : 4'b1000;
														assign node11329 = (inp[13]) ? node11331 : 4'b0000;
															assign node11331 = (inp[12]) ? 4'b0000 : 4'b1000;
												assign node11334 = (inp[12]) ? node11344 : node11335;
													assign node11335 = (inp[4]) ? node11339 : node11336;
														assign node11336 = (inp[0]) ? 4'b1100 : 4'b0000;
														assign node11339 = (inp[13]) ? 4'b1000 : node11340;
															assign node11340 = (inp[0]) ? 4'b0000 : 4'b1100;
													assign node11344 = (inp[14]) ? node11346 : 4'b0000;
														assign node11346 = (inp[0]) ? 4'b1100 : 4'b0100;
										assign node11349 = (inp[13]) ? node11383 : node11350;
											assign node11350 = (inp[0]) ? node11374 : node11351;
												assign node11351 = (inp[12]) ? node11369 : node11352;
													assign node11352 = (inp[14]) ? node11358 : node11353;
														assign node11353 = (inp[2]) ? node11355 : 4'b0100;
															assign node11355 = (inp[4]) ? 4'b1000 : 4'b0000;
														assign node11358 = (inp[7]) ? node11364 : node11359;
															assign node11359 = (inp[4]) ? 4'b1000 : node11360;
																assign node11360 = (inp[2]) ? 4'b0000 : 4'b1000;
															assign node11364 = (inp[2]) ? 4'b1000 : node11365;
																assign node11365 = (inp[4]) ? 4'b0100 : 4'b1000;
													assign node11369 = (inp[2]) ? node11371 : 4'b1000;
														assign node11371 = (inp[4]) ? 4'b1000 : 4'b0000;
												assign node11374 = (inp[2]) ? 4'b0000 : node11375;
													assign node11375 = (inp[4]) ? node11379 : node11376;
														assign node11376 = (inp[7]) ? 4'b0100 : 4'b1000;
														assign node11379 = (inp[7]) ? 4'b1000 : 4'b0000;
											assign node11383 = (inp[4]) ? 4'b1000 : node11384;
												assign node11384 = (inp[0]) ? node11390 : node11385;
													assign node11385 = (inp[2]) ? 4'b1100 : node11386;
														assign node11386 = (inp[7]) ? 4'b1100 : 4'b1000;
													assign node11390 = (inp[7]) ? node11392 : 4'b1000;
														assign node11392 = (inp[2]) ? 4'b1100 : 4'b1000;
							assign node11396 = (inp[4]) ? node11708 : node11397;
								assign node11397 = (inp[11]) ? node11591 : node11398;
									assign node11398 = (inp[2]) ? node11492 : node11399;
										assign node11399 = (inp[13]) ? node11449 : node11400;
											assign node11400 = (inp[10]) ? node11416 : node11401;
												assign node11401 = (inp[7]) ? node11403 : 4'b0000;
													assign node11403 = (inp[0]) ? node11409 : node11404;
														assign node11404 = (inp[14]) ? node11406 : 4'b0000;
															assign node11406 = (inp[1]) ? 4'b0000 : 4'b0001;
														assign node11409 = (inp[1]) ? node11413 : node11410;
															assign node11410 = (inp[14]) ? 4'b1001 : 4'b1000;
															assign node11413 = (inp[14]) ? 4'b0000 : 4'b0001;
												assign node11416 = (inp[0]) ? node11430 : node11417;
													assign node11417 = (inp[7]) ? 4'b1000 : node11418;
														assign node11418 = (inp[12]) ? node11424 : node11419;
															assign node11419 = (inp[14]) ? 4'b1000 : node11420;
																assign node11420 = (inp[1]) ? 4'b0001 : 4'b1001;
															assign node11424 = (inp[14]) ? node11426 : 4'b1000;
																assign node11426 = (inp[1]) ? 4'b0001 : 4'b0000;
													assign node11430 = (inp[14]) ? node11440 : node11431;
														assign node11431 = (inp[12]) ? node11437 : node11432;
															assign node11432 = (inp[7]) ? node11434 : 4'b0000;
																assign node11434 = (inp[1]) ? 4'b1000 : 4'b0000;
															assign node11437 = (inp[1]) ? 4'b0000 : 4'b1000;
														assign node11440 = (inp[7]) ? node11444 : node11441;
															assign node11441 = (inp[12]) ? 4'b1000 : 4'b0000;
															assign node11444 = (inp[1]) ? 4'b0000 : node11445;
																assign node11445 = (inp[12]) ? 4'b0001 : 4'b0000;
											assign node11449 = (inp[1]) ? node11467 : node11450;
												assign node11450 = (inp[0]) ? node11460 : node11451;
													assign node11451 = (inp[10]) ? node11453 : 4'b0001;
														assign node11453 = (inp[14]) ? node11457 : node11454;
															assign node11454 = (inp[7]) ? 4'b0000 : 4'b0001;
															assign node11457 = (inp[7]) ? 4'b1000 : 4'b0000;
													assign node11460 = (inp[12]) ? node11462 : 4'b1001;
														assign node11462 = (inp[7]) ? 4'b1000 : node11463;
															assign node11463 = (inp[10]) ? 4'b0001 : 4'b0000;
												assign node11467 = (inp[12]) ? node11479 : node11468;
													assign node11468 = (inp[14]) ? node11474 : node11469;
														assign node11469 = (inp[10]) ? 4'b0001 : node11470;
															assign node11470 = (inp[0]) ? 4'b0000 : 4'b0001;
														assign node11474 = (inp[10]) ? 4'b0000 : node11475;
															assign node11475 = (inp[0]) ? 4'b0001 : 4'b0000;
													assign node11479 = (inp[7]) ? node11487 : node11480;
														assign node11480 = (inp[14]) ? node11482 : 4'b0000;
															assign node11482 = (inp[0]) ? node11484 : 4'b0000;
																assign node11484 = (inp[10]) ? 4'b0000 : 4'b1001;
														assign node11487 = (inp[14]) ? 4'b0001 : node11488;
															assign node11488 = (inp[10]) ? 4'b1000 : 4'b0001;
										assign node11492 = (inp[12]) ? node11542 : node11493;
											assign node11493 = (inp[14]) ? node11515 : node11494;
												assign node11494 = (inp[10]) ? node11506 : node11495;
													assign node11495 = (inp[0]) ? node11499 : node11496;
														assign node11496 = (inp[13]) ? 4'b0000 : 4'b0001;
														assign node11499 = (inp[1]) ? 4'b0001 : node11500;
															assign node11500 = (inp[7]) ? node11502 : 4'b1001;
																assign node11502 = (inp[13]) ? 4'b0001 : 4'b1001;
													assign node11506 = (inp[0]) ? node11508 : 4'b0001;
														assign node11508 = (inp[1]) ? 4'b0000 : node11509;
															assign node11509 = (inp[7]) ? 4'b0001 : node11510;
																assign node11510 = (inp[13]) ? 4'b0000 : 4'b0001;
												assign node11515 = (inp[1]) ? node11529 : node11516;
													assign node11516 = (inp[7]) ? node11522 : node11517;
														assign node11517 = (inp[13]) ? 4'b0000 : node11518;
															assign node11518 = (inp[0]) ? 4'b0001 : 4'b1001;
														assign node11522 = (inp[10]) ? 4'b0000 : node11523;
															assign node11523 = (inp[0]) ? 4'b0000 : node11524;
																assign node11524 = (inp[13]) ? 4'b1001 : 4'b0000;
													assign node11529 = (inp[7]) ? node11535 : node11530;
														assign node11530 = (inp[10]) ? node11532 : 4'b0001;
															assign node11532 = (inp[13]) ? 4'b1000 : 4'b1001;
														assign node11535 = (inp[10]) ? node11539 : node11536;
															assign node11536 = (inp[0]) ? 4'b0001 : 4'b1001;
															assign node11539 = (inp[0]) ? 4'b1001 : 4'b0001;
											assign node11542 = (inp[10]) ? node11568 : node11543;
												assign node11543 = (inp[13]) ? node11555 : node11544;
													assign node11544 = (inp[7]) ? node11546 : 4'b1001;
														assign node11546 = (inp[0]) ? node11548 : 4'b1000;
															assign node11548 = (inp[14]) ? node11552 : node11549;
																assign node11549 = (inp[1]) ? 4'b1000 : 4'b1001;
																assign node11552 = (inp[1]) ? 4'b1001 : 4'b1000;
													assign node11555 = (inp[0]) ? node11563 : node11556;
														assign node11556 = (inp[1]) ? 4'b0000 : node11557;
															assign node11557 = (inp[14]) ? node11559 : 4'b1000;
																assign node11559 = (inp[7]) ? 4'b0001 : 4'b0000;
														assign node11563 = (inp[7]) ? node11565 : 4'b1001;
															assign node11565 = (inp[1]) ? 4'b0000 : 4'b0001;
												assign node11568 = (inp[0]) ? node11580 : node11569;
													assign node11569 = (inp[1]) ? node11575 : node11570;
														assign node11570 = (inp[13]) ? node11572 : 4'b0001;
															assign node11572 = (inp[7]) ? 4'b0000 : 4'b1001;
														assign node11575 = (inp[13]) ? 4'b1001 : node11576;
															assign node11576 = (inp[14]) ? 4'b1000 : 4'b1001;
													assign node11580 = (inp[7]) ? node11584 : node11581;
														assign node11581 = (inp[13]) ? 4'b0000 : 4'b0001;
														assign node11584 = (inp[13]) ? 4'b0001 : node11585;
															assign node11585 = (inp[14]) ? node11587 : 4'b0000;
																assign node11587 = (inp[1]) ? 4'b1001 : 4'b1000;
									assign node11591 = (inp[1]) ? node11665 : node11592;
										assign node11592 = (inp[7]) ? node11614 : node11593;
											assign node11593 = (inp[13]) ? node11611 : node11594;
												assign node11594 = (inp[0]) ? node11602 : node11595;
													assign node11595 = (inp[10]) ? 4'b0001 : node11596;
														assign node11596 = (inp[2]) ? node11598 : 4'b1000;
															assign node11598 = (inp[14]) ? 4'b0000 : 4'b1000;
													assign node11602 = (inp[2]) ? node11604 : 4'b0000;
														assign node11604 = (inp[14]) ? node11606 : 4'b0000;
															assign node11606 = (inp[10]) ? node11608 : 4'b1001;
																assign node11608 = (inp[12]) ? 4'b0000 : 4'b1000;
												assign node11611 = (inp[2]) ? 4'b1000 : 4'b1001;
											assign node11614 = (inp[10]) ? node11636 : node11615;
												assign node11615 = (inp[13]) ? node11623 : node11616;
													assign node11616 = (inp[0]) ? node11618 : 4'b0001;
														assign node11618 = (inp[2]) ? 4'b1001 : node11619;
															assign node11619 = (inp[12]) ? 4'b1001 : 4'b0001;
													assign node11623 = (inp[2]) ? node11629 : node11624;
														assign node11624 = (inp[12]) ? node11626 : 4'b0000;
															assign node11626 = (inp[0]) ? 4'b0000 : 4'b1000;
														assign node11629 = (inp[12]) ? node11633 : node11630;
															assign node11630 = (inp[14]) ? 4'b0001 : 4'b0000;
															assign node11633 = (inp[0]) ? 4'b0001 : 4'b1001;
												assign node11636 = (inp[12]) ? node11654 : node11637;
													assign node11637 = (inp[13]) ? node11647 : node11638;
														assign node11638 = (inp[14]) ? node11640 : 4'b0000;
															assign node11640 = (inp[2]) ? node11644 : node11641;
																assign node11641 = (inp[0]) ? 4'b0000 : 4'b0001;
																assign node11644 = (inp[0]) ? 4'b0001 : 4'b0000;
														assign node11647 = (inp[2]) ? node11651 : node11648;
															assign node11648 = (inp[0]) ? 4'b0000 : 4'b0001;
															assign node11651 = (inp[0]) ? 4'b1000 : 4'b1001;
													assign node11654 = (inp[13]) ? node11658 : node11655;
														assign node11655 = (inp[0]) ? 4'b0000 : 4'b1000;
														assign node11658 = (inp[0]) ? node11662 : node11659;
															assign node11659 = (inp[2]) ? 4'b0001 : 4'b0000;
															assign node11662 = (inp[2]) ? 4'b0000 : 4'b1001;
										assign node11665 = (inp[13]) ? node11691 : node11666;
											assign node11666 = (inp[0]) ? node11676 : node11667;
												assign node11667 = (inp[7]) ? 4'b0000 : node11668;
													assign node11668 = (inp[2]) ? 4'b0000 : node11669;
														assign node11669 = (inp[12]) ? 4'b1000 : node11670;
															assign node11670 = (inp[10]) ? 4'b1000 : 4'b0000;
												assign node11676 = (inp[2]) ? node11686 : node11677;
													assign node11677 = (inp[7]) ? node11681 : node11678;
														assign node11678 = (inp[10]) ? 4'b0000 : 4'b1000;
														assign node11681 = (inp[10]) ? 4'b1000 : node11682;
															assign node11682 = (inp[12]) ? 4'b0000 : 4'b1000;
													assign node11686 = (inp[7]) ? 4'b0000 : node11687;
														assign node11687 = (inp[10]) ? 4'b1000 : 4'b0000;
											assign node11691 = (inp[10]) ? 4'b1000 : node11692;
												assign node11692 = (inp[0]) ? node11700 : node11693;
													assign node11693 = (inp[14]) ? 4'b1000 : node11694;
														assign node11694 = (inp[12]) ? node11696 : 4'b1000;
															assign node11696 = (inp[2]) ? 4'b0000 : 4'b1000;
													assign node11700 = (inp[7]) ? node11702 : 4'b0000;
														assign node11702 = (inp[12]) ? 4'b0000 : node11703;
															assign node11703 = (inp[2]) ? 4'b0000 : 4'b1000;
								assign node11708 = (inp[13]) ? node11864 : node11709;
									assign node11709 = (inp[10]) ? node11803 : node11710;
										assign node11710 = (inp[12]) ? node11756 : node11711;
											assign node11711 = (inp[0]) ? node11735 : node11712;
												assign node11712 = (inp[1]) ? node11726 : node11713;
													assign node11713 = (inp[14]) ? node11719 : node11714;
														assign node11714 = (inp[11]) ? node11716 : 4'b1000;
															assign node11716 = (inp[7]) ? 4'b1000 : 4'b0000;
														assign node11719 = (inp[2]) ? node11721 : 4'b1001;
															assign node11721 = (inp[11]) ? 4'b0001 : node11722;
																assign node11722 = (inp[7]) ? 4'b0001 : 4'b1000;
													assign node11726 = (inp[11]) ? node11730 : node11727;
														assign node11727 = (inp[2]) ? 4'b0000 : 4'b0001;
														assign node11730 = (inp[7]) ? node11732 : 4'b0000;
															assign node11732 = (inp[2]) ? 4'b0000 : 4'b1000;
												assign node11735 = (inp[2]) ? node11745 : node11736;
													assign node11736 = (inp[7]) ? 4'b0000 : node11737;
														assign node11737 = (inp[11]) ? 4'b1000 : node11738;
															assign node11738 = (inp[14]) ? 4'b0001 : node11739;
																assign node11739 = (inp[1]) ? 4'b1000 : 4'b0000;
													assign node11745 = (inp[7]) ? node11747 : 4'b0000;
														assign node11747 = (inp[11]) ? node11753 : node11748;
															assign node11748 = (inp[1]) ? node11750 : 4'b0000;
																assign node11750 = (inp[14]) ? 4'b0000 : 4'b0001;
															assign node11753 = (inp[14]) ? 4'b0001 : 4'b1000;
											assign node11756 = (inp[1]) ? node11784 : node11757;
												assign node11757 = (inp[14]) ? node11771 : node11758;
													assign node11758 = (inp[2]) ? node11766 : node11759;
														assign node11759 = (inp[7]) ? node11761 : 4'b1000;
															assign node11761 = (inp[0]) ? node11763 : 4'b1000;
																assign node11763 = (inp[11]) ? 4'b0001 : 4'b0000;
														assign node11766 = (inp[0]) ? 4'b1001 : node11767;
															assign node11767 = (inp[11]) ? 4'b0001 : 4'b0000;
													assign node11771 = (inp[11]) ? node11777 : node11772;
														assign node11772 = (inp[2]) ? node11774 : 4'b1000;
															assign node11774 = (inp[0]) ? 4'b1001 : 4'b0001;
														assign node11777 = (inp[2]) ? node11781 : node11778;
															assign node11778 = (inp[7]) ? 4'b0001 : 4'b1001;
															assign node11781 = (inp[7]) ? 4'b1000 : 4'b0001;
												assign node11784 = (inp[0]) ? node11794 : node11785;
													assign node11785 = (inp[7]) ? node11789 : node11786;
														assign node11786 = (inp[2]) ? 4'b0000 : 4'b1000;
														assign node11789 = (inp[2]) ? 4'b1000 : node11790;
															assign node11790 = (inp[14]) ? 4'b1001 : 4'b1000;
													assign node11794 = (inp[11]) ? node11796 : 4'b0000;
														assign node11796 = (inp[14]) ? node11798 : 4'b1000;
															assign node11798 = (inp[7]) ? node11800 : 4'b0000;
																assign node11800 = (inp[2]) ? 4'b0000 : 4'b1000;
										assign node11803 = (inp[11]) ? node11847 : node11804;
											assign node11804 = (inp[12]) ? node11820 : node11805;
												assign node11805 = (inp[7]) ? node11807 : 4'b0001;
													assign node11807 = (inp[0]) ? node11815 : node11808;
														assign node11808 = (inp[1]) ? 4'b0001 : node11809;
															assign node11809 = (inp[2]) ? 4'b0001 : node11810;
																assign node11810 = (inp[14]) ? 4'b0000 : 4'b0001;
														assign node11815 = (inp[1]) ? 4'b0000 : node11816;
															assign node11816 = (inp[2]) ? 4'b0000 : 4'b1001;
												assign node11820 = (inp[0]) ? node11834 : node11821;
													assign node11821 = (inp[7]) ? node11829 : node11822;
														assign node11822 = (inp[2]) ? node11826 : node11823;
															assign node11823 = (inp[14]) ? 4'b0000 : 4'b0001;
															assign node11826 = (inp[1]) ? 4'b0000 : 4'b1000;
														assign node11829 = (inp[2]) ? 4'b0001 : node11830;
															assign node11830 = (inp[1]) ? 4'b1000 : 4'b0000;
													assign node11834 = (inp[14]) ? node11840 : node11835;
														assign node11835 = (inp[2]) ? 4'b0001 : node11836;
															assign node11836 = (inp[1]) ? 4'b0000 : 4'b0001;
														assign node11840 = (inp[2]) ? node11842 : 4'b0000;
															assign node11842 = (inp[1]) ? 4'b0000 : node11843;
																assign node11843 = (inp[7]) ? 4'b0001 : 4'b0000;
											assign node11847 = (inp[1]) ? 4'b0000 : node11848;
												assign node11848 = (inp[0]) ? node11856 : node11849;
													assign node11849 = (inp[2]) ? node11851 : 4'b0001;
														assign node11851 = (inp[7]) ? 4'b1000 : node11852;
															assign node11852 = (inp[12]) ? 4'b0000 : 4'b1000;
													assign node11856 = (inp[12]) ? node11858 : 4'b0000;
														assign node11858 = (inp[2]) ? node11860 : 4'b0000;
															assign node11860 = (inp[7]) ? 4'b0000 : 4'b0001;
									assign node11864 = (inp[10]) ? node11932 : node11865;
										assign node11865 = (inp[11]) ? node11909 : node11866;
											assign node11866 = (inp[0]) ? node11886 : node11867;
												assign node11867 = (inp[1]) ? node11881 : node11868;
													assign node11868 = (inp[7]) ? node11876 : node11869;
														assign node11869 = (inp[2]) ? 4'b0001 : node11870;
															assign node11870 = (inp[12]) ? node11872 : 4'b0000;
																assign node11872 = (inp[14]) ? 4'b0001 : 4'b0000;
														assign node11876 = (inp[2]) ? 4'b0000 : node11877;
															assign node11877 = (inp[14]) ? 4'b0000 : 4'b0001;
													assign node11881 = (inp[7]) ? 4'b0001 : node11882;
														assign node11882 = (inp[2]) ? 4'b0000 : 4'b0001;
												assign node11886 = (inp[1]) ? node11902 : node11887;
													assign node11887 = (inp[2]) ? 4'b0001 : node11888;
														assign node11888 = (inp[12]) ? node11894 : node11889;
															assign node11889 = (inp[14]) ? node11891 : 4'b0001;
																assign node11891 = (inp[7]) ? 4'b0001 : 4'b0000;
															assign node11894 = (inp[7]) ? node11898 : node11895;
																assign node11895 = (inp[14]) ? 4'b0000 : 4'b0001;
																assign node11898 = (inp[14]) ? 4'b0001 : 4'b0000;
													assign node11902 = (inp[2]) ? 4'b0000 : node11903;
														assign node11903 = (inp[7]) ? node11905 : 4'b0000;
															assign node11905 = (inp[14]) ? 4'b0001 : 4'b0000;
											assign node11909 = (inp[1]) ? 4'b0000 : node11910;
												assign node11910 = (inp[0]) ? node11918 : node11911;
													assign node11911 = (inp[7]) ? node11913 : 4'b0001;
														assign node11913 = (inp[12]) ? 4'b0000 : node11914;
															assign node11914 = (inp[14]) ? 4'b0001 : 4'b0000;
													assign node11918 = (inp[12]) ? node11924 : node11919;
														assign node11919 = (inp[7]) ? node11921 : 4'b0000;
															assign node11921 = (inp[2]) ? 4'b0001 : 4'b0000;
														assign node11924 = (inp[2]) ? node11928 : node11925;
															assign node11925 = (inp[7]) ? 4'b0001 : 4'b0000;
															assign node11928 = (inp[7]) ? 4'b0000 : 4'b0001;
										assign node11932 = (inp[1]) ? 4'b0000 : node11933;
											assign node11933 = (inp[11]) ? 4'b0000 : node11934;
												assign node11934 = (inp[7]) ? node11944 : node11935;
													assign node11935 = (inp[2]) ? node11937 : 4'b0000;
														assign node11937 = (inp[0]) ? 4'b0000 : node11938;
															assign node11938 = (inp[12]) ? node11940 : 4'b0000;
																assign node11940 = (inp[14]) ? 4'b0000 : 4'b0001;
													assign node11944 = (inp[0]) ? node11954 : node11945;
														assign node11945 = (inp[2]) ? 4'b0001 : node11946;
															assign node11946 = (inp[14]) ? node11950 : node11947;
																assign node11947 = (inp[12]) ? 4'b0001 : 4'b0000;
																assign node11950 = (inp[12]) ? 4'b0000 : 4'b0001;
														assign node11954 = (inp[12]) ? node11956 : 4'b0000;
															assign node11956 = (inp[14]) ? node11960 : node11957;
																assign node11957 = (inp[2]) ? 4'b0001 : 4'b0000;
																assign node11960 = (inp[2]) ? 4'b0000 : 4'b0001;
				assign node11965 = (inp[0]) ? node13567 : node11966;
					assign node11966 = (inp[6]) ? node12428 : node11967;
						assign node11967 = (inp[5]) ? node12065 : node11968;
							assign node11968 = (inp[3]) ? node11970 : 4'b1010;
								assign node11970 = (inp[2]) ? 4'b1010 : node11971;
									assign node11971 = (inp[7]) ? node12029 : node11972;
										assign node11972 = (inp[1]) ? node11994 : node11973;
											assign node11973 = (inp[13]) ? node11985 : node11974;
												assign node11974 = (inp[12]) ? node11982 : node11975;
													assign node11975 = (inp[10]) ? node11977 : 4'b1001;
														assign node11977 = (inp[14]) ? node11979 : 4'b0001;
															assign node11979 = (inp[11]) ? 4'b0001 : 4'b0000;
													assign node11982 = (inp[4]) ? 4'b1001 : 4'b1010;
												assign node11985 = (inp[10]) ? node11987 : 4'b0001;
													assign node11987 = (inp[12]) ? 4'b0001 : node11988;
														assign node11988 = (inp[14]) ? node11990 : 4'b1001;
															assign node11990 = (inp[11]) ? 4'b1001 : 4'b1000;
											assign node11994 = (inp[11]) ? node12018 : node11995;
												assign node11995 = (inp[14]) ? node12007 : node11996;
													assign node11996 = (inp[13]) ? node12002 : node11997;
														assign node11997 = (inp[12]) ? node11999 : 4'b0000;
															assign node11999 = (inp[4]) ? 4'b1000 : 4'b1010;
														assign node12002 = (inp[12]) ? node12004 : 4'b1000;
															assign node12004 = (inp[10]) ? 4'b1000 : 4'b0000;
													assign node12007 = (inp[4]) ? 4'b1001 : node12008;
														assign node12008 = (inp[13]) ? node12014 : node12009;
															assign node12009 = (inp[12]) ? 4'b1010 : node12010;
																assign node12010 = (inp[10]) ? 4'b0001 : 4'b1010;
															assign node12014 = (inp[12]) ? 4'b0001 : 4'b1001;
												assign node12018 = (inp[13]) ? node12026 : node12019;
													assign node12019 = (inp[12]) ? node12021 : 4'b0000;
														assign node12021 = (inp[4]) ? node12023 : 4'b1010;
															assign node12023 = (inp[10]) ? 4'b0000 : 4'b1000;
													assign node12026 = (inp[12]) ? 4'b0000 : 4'b1000;
										assign node12029 = (inp[4]) ? node12031 : 4'b1010;
											assign node12031 = (inp[13]) ? node12041 : node12032;
												assign node12032 = (inp[10]) ? node12034 : 4'b1010;
													assign node12034 = (inp[12]) ? 4'b1010 : node12035;
														assign node12035 = (inp[1]) ? 4'b0000 : node12036;
															assign node12036 = (inp[11]) ? 4'b0001 : 4'b0000;
												assign node12041 = (inp[10]) ? node12047 : node12042;
													assign node12042 = (inp[1]) ? node12044 : 4'b0001;
														assign node12044 = (inp[14]) ? 4'b0001 : 4'b1000;
													assign node12047 = (inp[12]) ? node12057 : node12048;
														assign node12048 = (inp[14]) ? node12050 : 4'b1001;
															assign node12050 = (inp[11]) ? node12054 : node12051;
																assign node12051 = (inp[1]) ? 4'b1001 : 4'b1000;
																assign node12054 = (inp[1]) ? 4'b1000 : 4'b1001;
														assign node12057 = (inp[14]) ? node12059 : 4'b1000;
															assign node12059 = (inp[11]) ? 4'b0001 : node12060;
																assign node12060 = (inp[1]) ? 4'b0001 : 4'b0000;
							assign node12065 = (inp[2]) ? node12333 : node12066;
								assign node12066 = (inp[1]) ? node12196 : node12067;
									assign node12067 = (inp[11]) ? node12141 : node12068;
										assign node12068 = (inp[14]) ? node12104 : node12069;
											assign node12069 = (inp[13]) ? node12085 : node12070;
												assign node12070 = (inp[10]) ? node12078 : node12071;
													assign node12071 = (inp[3]) ? node12073 : 4'b1001;
														assign node12073 = (inp[7]) ? 4'b1101 : node12074;
															assign node12074 = (inp[4]) ? 4'b1001 : 4'b1101;
													assign node12078 = (inp[12]) ? 4'b1101 : node12079;
														assign node12079 = (inp[3]) ? 4'b0001 : node12080;
															assign node12080 = (inp[4]) ? 4'b0101 : 4'b0001;
												assign node12085 = (inp[12]) ? node12095 : node12086;
													assign node12086 = (inp[10]) ? node12088 : 4'b0101;
														assign node12088 = (inp[3]) ? node12092 : node12089;
															assign node12089 = (inp[7]) ? 4'b1001 : 4'b1101;
															assign node12092 = (inp[7]) ? 4'b1101 : 4'b1001;
													assign node12095 = (inp[4]) ? 4'b0101 : node12096;
														assign node12096 = (inp[10]) ? node12098 : 4'b0001;
															assign node12098 = (inp[3]) ? 4'b0101 : node12099;
																assign node12099 = (inp[7]) ? 4'b0001 : 4'b0101;
											assign node12104 = (inp[13]) ? node12120 : node12105;
												assign node12105 = (inp[3]) ? node12113 : node12106;
													assign node12106 = (inp[7]) ? 4'b1000 : node12107;
														assign node12107 = (inp[10]) ? 4'b0100 : node12108;
															assign node12108 = (inp[4]) ? 4'b1100 : 4'b1000;
													assign node12113 = (inp[7]) ? node12117 : node12114;
														assign node12114 = (inp[4]) ? 4'b1000 : 4'b1100;
														assign node12117 = (inp[12]) ? 4'b1100 : 4'b0100;
												assign node12120 = (inp[3]) ? node12130 : node12121;
													assign node12121 = (inp[4]) ? node12125 : node12122;
														assign node12122 = (inp[7]) ? 4'b0000 : 4'b0100;
														assign node12125 = (inp[12]) ? 4'b0100 : node12126;
															assign node12126 = (inp[10]) ? 4'b1100 : 4'b0100;
													assign node12130 = (inp[4]) ? node12136 : node12131;
														assign node12131 = (inp[7]) ? node12133 : 4'b0000;
															assign node12133 = (inp[12]) ? 4'b0100 : 4'b1100;
														assign node12136 = (inp[12]) ? 4'b0000 : node12137;
															assign node12137 = (inp[10]) ? 4'b1000 : 4'b0000;
										assign node12141 = (inp[13]) ? node12171 : node12142;
											assign node12142 = (inp[10]) ? node12154 : node12143;
												assign node12143 = (inp[3]) ? node12149 : node12144;
													assign node12144 = (inp[4]) ? node12146 : 4'b1001;
														assign node12146 = (inp[14]) ? 4'b1101 : 4'b1001;
													assign node12149 = (inp[7]) ? 4'b1101 : node12150;
														assign node12150 = (inp[4]) ? 4'b1001 : 4'b1101;
												assign node12154 = (inp[12]) ? node12166 : node12155;
													assign node12155 = (inp[3]) ? node12161 : node12156;
														assign node12156 = (inp[7]) ? node12158 : 4'b0101;
															assign node12158 = (inp[4]) ? 4'b0101 : 4'b0001;
														assign node12161 = (inp[7]) ? node12163 : 4'b0001;
															assign node12163 = (inp[4]) ? 4'b0001 : 4'b0101;
													assign node12166 = (inp[3]) ? node12168 : 4'b1001;
														assign node12168 = (inp[4]) ? 4'b1001 : 4'b1101;
											assign node12171 = (inp[10]) ? node12179 : node12172;
												assign node12172 = (inp[3]) ? node12174 : 4'b0101;
													assign node12174 = (inp[4]) ? 4'b0001 : node12175;
														assign node12175 = (inp[7]) ? 4'b0101 : 4'b0001;
												assign node12179 = (inp[12]) ? node12185 : node12180;
													assign node12180 = (inp[7]) ? 4'b1101 : node12181;
														assign node12181 = (inp[3]) ? 4'b1001 : 4'b1101;
													assign node12185 = (inp[14]) ? node12187 : 4'b0101;
														assign node12187 = (inp[7]) ? node12189 : 4'b0001;
															assign node12189 = (inp[4]) ? node12193 : node12190;
																assign node12190 = (inp[3]) ? 4'b0101 : 4'b0001;
																assign node12193 = (inp[3]) ? 4'b0001 : 4'b0101;
									assign node12196 = (inp[11]) ? node12276 : node12197;
										assign node12197 = (inp[14]) ? node12235 : node12198;
											assign node12198 = (inp[13]) ? node12218 : node12199;
												assign node12199 = (inp[12]) ? node12211 : node12200;
													assign node12200 = (inp[7]) ? node12202 : 4'b0100;
														assign node12202 = (inp[10]) ? node12206 : node12203;
															assign node12203 = (inp[3]) ? 4'b0100 : 4'b0000;
															assign node12206 = (inp[4]) ? node12208 : 4'b0000;
																assign node12208 = (inp[3]) ? 4'b0000 : 4'b0100;
													assign node12211 = (inp[10]) ? node12215 : node12212;
														assign node12212 = (inp[3]) ? 4'b1100 : 4'b1000;
														assign node12215 = (inp[4]) ? 4'b0100 : 4'b0000;
												assign node12218 = (inp[10]) ? node12228 : node12219;
													assign node12219 = (inp[12]) ? node12223 : node12220;
														assign node12220 = (inp[7]) ? 4'b1000 : 4'b1100;
														assign node12223 = (inp[3]) ? node12225 : 4'b0100;
															assign node12225 = (inp[4]) ? 4'b0000 : 4'b0100;
													assign node12228 = (inp[4]) ? node12232 : node12229;
														assign node12229 = (inp[3]) ? 4'b1100 : 4'b1000;
														assign node12232 = (inp[3]) ? 4'b1000 : 4'b1100;
											assign node12235 = (inp[13]) ? node12257 : node12236;
												assign node12236 = (inp[10]) ? node12248 : node12237;
													assign node12237 = (inp[3]) ? node12243 : node12238;
														assign node12238 = (inp[4]) ? node12240 : 4'b1001;
															assign node12240 = (inp[7]) ? 4'b1001 : 4'b1101;
														assign node12243 = (inp[7]) ? 4'b1101 : node12244;
															assign node12244 = (inp[4]) ? 4'b1001 : 4'b1101;
													assign node12248 = (inp[12]) ? 4'b1101 : node12249;
														assign node12249 = (inp[3]) ? node12251 : 4'b0101;
															assign node12251 = (inp[4]) ? 4'b0001 : node12252;
																assign node12252 = (inp[7]) ? 4'b0101 : 4'b0001;
												assign node12257 = (inp[10]) ? node12263 : node12258;
													assign node12258 = (inp[7]) ? 4'b0001 : node12259;
														assign node12259 = (inp[3]) ? 4'b0001 : 4'b0101;
													assign node12263 = (inp[12]) ? node12273 : node12264;
														assign node12264 = (inp[7]) ? node12266 : 4'b1101;
															assign node12266 = (inp[3]) ? node12270 : node12267;
																assign node12267 = (inp[4]) ? 4'b1101 : 4'b1001;
																assign node12270 = (inp[4]) ? 4'b1001 : 4'b1101;
														assign node12273 = (inp[4]) ? 4'b0001 : 4'b0101;
										assign node12276 = (inp[13]) ? node12308 : node12277;
											assign node12277 = (inp[12]) ? node12293 : node12278;
												assign node12278 = (inp[14]) ? node12288 : node12279;
													assign node12279 = (inp[3]) ? node12285 : node12280;
														assign node12280 = (inp[4]) ? 4'b0100 : node12281;
															assign node12281 = (inp[7]) ? 4'b0000 : 4'b0100;
														assign node12285 = (inp[4]) ? 4'b0000 : 4'b0100;
													assign node12288 = (inp[7]) ? 4'b0000 : node12289;
														assign node12289 = (inp[3]) ? 4'b0000 : 4'b0100;
												assign node12293 = (inp[10]) ? node12301 : node12294;
													assign node12294 = (inp[3]) ? node12298 : node12295;
														assign node12295 = (inp[7]) ? 4'b1000 : 4'b1100;
														assign node12298 = (inp[4]) ? 4'b1000 : 4'b1100;
													assign node12301 = (inp[3]) ? node12303 : 4'b0100;
														assign node12303 = (inp[4]) ? 4'b0000 : node12304;
															assign node12304 = (inp[14]) ? 4'b0000 : 4'b0100;
											assign node12308 = (inp[3]) ? node12320 : node12309;
												assign node12309 = (inp[7]) ? node12315 : node12310;
													assign node12310 = (inp[12]) ? node12312 : 4'b1100;
														assign node12312 = (inp[10]) ? 4'b1100 : 4'b0100;
													assign node12315 = (inp[4]) ? 4'b1100 : node12316;
														assign node12316 = (inp[10]) ? 4'b1000 : 4'b0000;
												assign node12320 = (inp[7]) ? node12326 : node12321;
													assign node12321 = (inp[10]) ? 4'b1000 : node12322;
														assign node12322 = (inp[12]) ? 4'b0000 : 4'b1000;
													assign node12326 = (inp[10]) ? node12330 : node12327;
														assign node12327 = (inp[4]) ? 4'b0000 : 4'b0100;
														assign node12330 = (inp[4]) ? 4'b1000 : 4'b1100;
								assign node12333 = (inp[3]) ? node12335 : 4'b1010;
									assign node12335 = (inp[4]) ? node12367 : node12336;
										assign node12336 = (inp[7]) ? 4'b1010 : node12337;
											assign node12337 = (inp[10]) ? node12347 : node12338;
												assign node12338 = (inp[13]) ? 4'b0000 : node12339;
													assign node12339 = (inp[12]) ? 4'b1010 : node12340;
														assign node12340 = (inp[14]) ? 4'b1010 : node12341;
															assign node12341 = (inp[1]) ? 4'b0000 : 4'b1010;
												assign node12347 = (inp[13]) ? node12355 : node12348;
													assign node12348 = (inp[12]) ? node12352 : node12349;
														assign node12349 = (inp[11]) ? 4'b0000 : 4'b0001;
														assign node12352 = (inp[1]) ? 4'b0000 : 4'b1010;
													assign node12355 = (inp[12]) ? node12359 : node12356;
														assign node12356 = (inp[1]) ? 4'b1000 : 4'b1001;
														assign node12359 = (inp[1]) ? node12363 : node12360;
															assign node12360 = (inp[14]) ? 4'b0000 : 4'b0001;
															assign node12363 = (inp[14]) ? 4'b0001 : 4'b1000;
										assign node12367 = (inp[13]) ? node12401 : node12368;
											assign node12368 = (inp[7]) ? node12392 : node12369;
												assign node12369 = (inp[1]) ? node12383 : node12370;
													assign node12370 = (inp[11]) ? node12378 : node12371;
														assign node12371 = (inp[14]) ? node12373 : 4'b1001;
															assign node12373 = (inp[12]) ? 4'b1000 : node12374;
																assign node12374 = (inp[10]) ? 4'b0000 : 4'b1000;
														assign node12378 = (inp[10]) ? node12380 : 4'b1001;
															assign node12380 = (inp[12]) ? 4'b1001 : 4'b0001;
													assign node12383 = (inp[10]) ? 4'b0000 : node12384;
														assign node12384 = (inp[14]) ? node12388 : node12385;
															assign node12385 = (inp[12]) ? 4'b1000 : 4'b0000;
															assign node12388 = (inp[11]) ? 4'b1000 : 4'b1001;
												assign node12392 = (inp[10]) ? node12394 : 4'b1010;
													assign node12394 = (inp[1]) ? node12398 : node12395;
														assign node12395 = (inp[12]) ? 4'b1010 : 4'b0001;
														assign node12398 = (inp[11]) ? 4'b0000 : 4'b0001;
											assign node12401 = (inp[1]) ? node12411 : node12402;
												assign node12402 = (inp[10]) ? node12408 : node12403;
													assign node12403 = (inp[14]) ? node12405 : 4'b0001;
														assign node12405 = (inp[11]) ? 4'b0001 : 4'b0000;
													assign node12408 = (inp[12]) ? 4'b0001 : 4'b1001;
												assign node12411 = (inp[14]) ? node12417 : node12412;
													assign node12412 = (inp[12]) ? node12414 : 4'b1000;
														assign node12414 = (inp[10]) ? 4'b1000 : 4'b0000;
													assign node12417 = (inp[11]) ? node12423 : node12418;
														assign node12418 = (inp[12]) ? 4'b0001 : node12419;
															assign node12419 = (inp[10]) ? 4'b1001 : 4'b0001;
														assign node12423 = (inp[12]) ? node12425 : 4'b1000;
															assign node12425 = (inp[10]) ? 4'b1000 : 4'b0000;
						assign node12428 = (inp[5]) ? node13014 : node12429;
							assign node12429 = (inp[11]) ? node12773 : node12430;
								assign node12430 = (inp[3]) ? node12604 : node12431;
									assign node12431 = (inp[7]) ? node12523 : node12432;
										assign node12432 = (inp[2]) ? node12476 : node12433;
											assign node12433 = (inp[4]) ? node12461 : node12434;
												assign node12434 = (inp[13]) ? node12448 : node12435;
													assign node12435 = (inp[14]) ? node12441 : node12436;
														assign node12436 = (inp[1]) ? 4'b0100 : node12437;
															assign node12437 = (inp[10]) ? 4'b0101 : 4'b1001;
														assign node12441 = (inp[1]) ? node12443 : 4'b1000;
															assign node12443 = (inp[10]) ? node12445 : 4'b1001;
																assign node12445 = (inp[12]) ? 4'b1001 : 4'b0101;
													assign node12448 = (inp[10]) ? node12458 : node12449;
														assign node12449 = (inp[12]) ? node12451 : 4'b0100;
															assign node12451 = (inp[14]) ? node12455 : node12452;
																assign node12452 = (inp[1]) ? 4'b0100 : 4'b0101;
																assign node12455 = (inp[1]) ? 4'b0101 : 4'b0100;
														assign node12458 = (inp[12]) ? 4'b0100 : 4'b1101;
												assign node12461 = (inp[10]) ? node12471 : node12462;
													assign node12462 = (inp[13]) ? 4'b1001 : node12463;
														assign node12463 = (inp[1]) ? node12467 : node12464;
															assign node12464 = (inp[14]) ? 4'b1100 : 4'b1101;
															assign node12467 = (inp[12]) ? 4'b1101 : 4'b0001;
													assign node12471 = (inp[1]) ? node12473 : 4'b0001;
														assign node12473 = (inp[13]) ? 4'b1001 : 4'b0001;
											assign node12476 = (inp[13]) ? node12500 : node12477;
												assign node12477 = (inp[14]) ? node12487 : node12478;
													assign node12478 = (inp[1]) ? node12482 : node12479;
														assign node12479 = (inp[4]) ? 4'b1101 : 4'b0101;
														assign node12482 = (inp[4]) ? node12484 : 4'b0100;
															assign node12484 = (inp[10]) ? 4'b0100 : 4'b1100;
													assign node12487 = (inp[1]) ? node12495 : node12488;
														assign node12488 = (inp[12]) ? node12492 : node12489;
															assign node12489 = (inp[10]) ? 4'b0100 : 4'b1000;
															assign node12492 = (inp[10]) ? 4'b1000 : 4'b1100;
														assign node12495 = (inp[4]) ? node12497 : 4'b1001;
															assign node12497 = (inp[10]) ? 4'b0101 : 4'b1101;
												assign node12500 = (inp[12]) ? node12514 : node12501;
													assign node12501 = (inp[10]) ? node12509 : node12502;
														assign node12502 = (inp[4]) ? 4'b1100 : node12503;
															assign node12503 = (inp[14]) ? node12505 : 4'b0101;
																assign node12505 = (inp[1]) ? 4'b0101 : 4'b0100;
														assign node12509 = (inp[1]) ? 4'b1100 : node12510;
															assign node12510 = (inp[14]) ? 4'b1100 : 4'b1101;
													assign node12514 = (inp[1]) ? node12518 : node12515;
														assign node12515 = (inp[14]) ? 4'b0100 : 4'b0101;
														assign node12518 = (inp[14]) ? 4'b0101 : node12519;
															assign node12519 = (inp[10]) ? 4'b1100 : 4'b0100;
										assign node12523 = (inp[4]) ? node12555 : node12524;
											assign node12524 = (inp[1]) ? node12542 : node12525;
												assign node12525 = (inp[14]) ? node12535 : node12526;
													assign node12526 = (inp[10]) ? node12528 : 4'b1001;
														assign node12528 = (inp[2]) ? 4'b0001 : node12529;
															assign node12529 = (inp[12]) ? 4'b1001 : node12530;
																assign node12530 = (inp[13]) ? 4'b1001 : 4'b0001;
													assign node12535 = (inp[13]) ? node12537 : 4'b1000;
														assign node12537 = (inp[10]) ? node12539 : 4'b0000;
															assign node12539 = (inp[12]) ? 4'b0000 : 4'b1000;
												assign node12542 = (inp[14]) ? node12548 : node12543;
													assign node12543 = (inp[13]) ? node12545 : 4'b0000;
														assign node12545 = (inp[12]) ? 4'b0000 : 4'b1000;
													assign node12548 = (inp[13]) ? node12550 : 4'b1001;
														assign node12550 = (inp[12]) ? 4'b0001 : node12551;
															assign node12551 = (inp[10]) ? 4'b1001 : 4'b0001;
											assign node12555 = (inp[13]) ? node12575 : node12556;
												assign node12556 = (inp[10]) ? node12564 : node12557;
													assign node12557 = (inp[14]) ? node12561 : node12558;
														assign node12558 = (inp[1]) ? 4'b1000 : 4'b1001;
														assign node12561 = (inp[1]) ? 4'b1001 : 4'b1000;
													assign node12564 = (inp[12]) ? node12570 : node12565;
														assign node12565 = (inp[1]) ? node12567 : 4'b0101;
															assign node12567 = (inp[14]) ? 4'b0101 : 4'b0100;
														assign node12570 = (inp[1]) ? 4'b0100 : node12571;
															assign node12571 = (inp[14]) ? 4'b1000 : 4'b1001;
												assign node12575 = (inp[2]) ? node12589 : node12576;
													assign node12576 = (inp[10]) ? node12586 : node12577;
														assign node12577 = (inp[14]) ? 4'b0100 : node12578;
															assign node12578 = (inp[12]) ? node12582 : node12579;
																assign node12579 = (inp[1]) ? 4'b0001 : 4'b0101;
																assign node12582 = (inp[1]) ? 4'b0100 : 4'b0101;
														assign node12586 = (inp[14]) ? 4'b1001 : 4'b0001;
													assign node12589 = (inp[12]) ? node12601 : node12590;
														assign node12590 = (inp[10]) ? node12594 : node12591;
															assign node12591 = (inp[14]) ? 4'b0100 : 4'b0101;
															assign node12594 = (inp[1]) ? node12598 : node12595;
																assign node12595 = (inp[14]) ? 4'b1100 : 4'b1101;
																assign node12598 = (inp[14]) ? 4'b1101 : 4'b1100;
														assign node12601 = (inp[14]) ? 4'b0100 : 4'b0101;
									assign node12604 = (inp[7]) ? node12684 : node12605;
										assign node12605 = (inp[4]) ? node12639 : node12606;
											assign node12606 = (inp[2]) ? node12624 : node12607;
												assign node12607 = (inp[10]) ? node12619 : node12608;
													assign node12608 = (inp[13]) ? node12614 : node12609;
														assign node12609 = (inp[12]) ? 4'b1001 : node12610;
															assign node12610 = (inp[1]) ? 4'b0101 : 4'b1001;
														assign node12614 = (inp[12]) ? 4'b1101 : node12615;
															assign node12615 = (inp[1]) ? 4'b0101 : 4'b1101;
													assign node12619 = (inp[1]) ? node12621 : 4'b0101;
														assign node12621 = (inp[13]) ? 4'b0101 : 4'b1101;
												assign node12624 = (inp[14]) ? node12632 : node12625;
													assign node12625 = (inp[1]) ? node12627 : 4'b0001;
														assign node12627 = (inp[13]) ? node12629 : 4'b0000;
															assign node12629 = (inp[10]) ? 4'b1000 : 4'b0000;
													assign node12632 = (inp[13]) ? node12636 : node12633;
														assign node12633 = (inp[1]) ? 4'b1101 : 4'b1100;
														assign node12636 = (inp[12]) ? 4'b0000 : 4'b1000;
											assign node12639 = (inp[10]) ? node12663 : node12640;
												assign node12640 = (inp[12]) ? node12656 : node12641;
													assign node12641 = (inp[1]) ? node12649 : node12642;
														assign node12642 = (inp[14]) ? node12646 : node12643;
															assign node12643 = (inp[2]) ? 4'b1001 : 4'b1000;
															assign node12646 = (inp[13]) ? 4'b0001 : 4'b1000;
														assign node12649 = (inp[13]) ? node12651 : 4'b0001;
															assign node12651 = (inp[14]) ? 4'b1000 : node12652;
																assign node12652 = (inp[2]) ? 4'b0001 : 4'b1001;
													assign node12656 = (inp[13]) ? node12660 : node12657;
														assign node12657 = (inp[2]) ? 4'b1001 : 4'b1101;
														assign node12660 = (inp[1]) ? 4'b1001 : 4'b0001;
												assign node12663 = (inp[2]) ? node12679 : node12664;
													assign node12664 = (inp[13]) ? node12672 : node12665;
														assign node12665 = (inp[14]) ? node12667 : 4'b0001;
															assign node12667 = (inp[12]) ? 4'b0001 : node12668;
																assign node12668 = (inp[1]) ? 4'b0000 : 4'b0001;
														assign node12672 = (inp[12]) ? node12674 : 4'b1000;
															assign node12674 = (inp[14]) ? 4'b0000 : node12675;
																assign node12675 = (inp[1]) ? 4'b0001 : 4'b0000;
													assign node12679 = (inp[1]) ? node12681 : 4'b0001;
														assign node12681 = (inp[12]) ? 4'b0001 : 4'b1001;
										assign node12684 = (inp[2]) ? node12726 : node12685;
											assign node12685 = (inp[10]) ? node12699 : node12686;
												assign node12686 = (inp[4]) ? node12694 : node12687;
													assign node12687 = (inp[12]) ? 4'b1001 : node12688;
														assign node12688 = (inp[14]) ? node12690 : 4'b0101;
															assign node12690 = (inp[13]) ? 4'b1001 : 4'b0001;
													assign node12694 = (inp[1]) ? node12696 : 4'b1101;
														assign node12696 = (inp[12]) ? 4'b1101 : 4'b0101;
												assign node12699 = (inp[12]) ? node12711 : node12700;
													assign node12700 = (inp[1]) ? node12704 : node12701;
														assign node12701 = (inp[4]) ? 4'b0000 : 4'b0101;
														assign node12704 = (inp[13]) ? node12708 : node12705;
															assign node12705 = (inp[4]) ? 4'b1101 : 4'b1001;
															assign node12708 = (inp[4]) ? 4'b1001 : 4'b1101;
													assign node12711 = (inp[1]) ? node12721 : node12712;
														assign node12712 = (inp[14]) ? node12716 : node12713;
															assign node12713 = (inp[13]) ? 4'b0000 : 4'b0101;
															assign node12716 = (inp[4]) ? 4'b0001 : node12717;
																assign node12717 = (inp[13]) ? 4'b0101 : 4'b0001;
														assign node12721 = (inp[4]) ? 4'b0101 : node12722;
															assign node12722 = (inp[13]) ? 4'b0101 : 4'b0001;
											assign node12726 = (inp[4]) ? node12758 : node12727;
												assign node12727 = (inp[12]) ? node12747 : node12728;
													assign node12728 = (inp[13]) ? node12738 : node12729;
														assign node12729 = (inp[10]) ? node12733 : node12730;
															assign node12730 = (inp[1]) ? 4'b1101 : 4'b1100;
															assign node12733 = (inp[1]) ? node12735 : 4'b0100;
																assign node12735 = (inp[14]) ? 4'b0101 : 4'b0100;
														assign node12738 = (inp[10]) ? node12740 : 4'b1100;
															assign node12740 = (inp[14]) ? node12744 : node12741;
																assign node12741 = (inp[1]) ? 4'b1100 : 4'b1101;
																assign node12744 = (inp[1]) ? 4'b1101 : 4'b1100;
													assign node12747 = (inp[13]) ? node12755 : node12748;
														assign node12748 = (inp[14]) ? node12752 : node12749;
															assign node12749 = (inp[1]) ? 4'b0100 : 4'b1101;
															assign node12752 = (inp[1]) ? 4'b1101 : 4'b1100;
														assign node12755 = (inp[10]) ? 4'b0101 : 4'b0100;
												assign node12758 = (inp[13]) ? node12766 : node12759;
													assign node12759 = (inp[12]) ? 4'b1101 : node12760;
														assign node12760 = (inp[10]) ? 4'b0000 : node12761;
															assign node12761 = (inp[14]) ? 4'b1100 : 4'b1101;
													assign node12766 = (inp[1]) ? 4'b0001 : node12767;
														assign node12767 = (inp[10]) ? 4'b0001 : node12768;
															assign node12768 = (inp[14]) ? 4'b0000 : 4'b0001;
								assign node12773 = (inp[1]) ? node12893 : node12774;
									assign node12774 = (inp[3]) ? node12830 : node12775;
										assign node12775 = (inp[7]) ? node12809 : node12776;
											assign node12776 = (inp[2]) ? node12792 : node12777;
												assign node12777 = (inp[4]) ? node12785 : node12778;
													assign node12778 = (inp[13]) ? node12782 : node12779;
														assign node12779 = (inp[12]) ? 4'b1001 : 4'b0101;
														assign node12782 = (inp[12]) ? 4'b0101 : 4'b1101;
													assign node12785 = (inp[10]) ? node12789 : node12786;
														assign node12786 = (inp[12]) ? 4'b1000 : 4'b0000;
														assign node12789 = (inp[12]) ? 4'b0000 : 4'b1000;
												assign node12792 = (inp[4]) ? node12800 : node12793;
													assign node12793 = (inp[12]) ? 4'b0101 : node12794;
														assign node12794 = (inp[14]) ? 4'b0101 : node12795;
															assign node12795 = (inp[13]) ? 4'b1101 : 4'b0101;
													assign node12800 = (inp[13]) ? node12806 : node12801;
														assign node12801 = (inp[10]) ? node12803 : 4'b1101;
															assign node12803 = (inp[12]) ? 4'b1101 : 4'b0101;
														assign node12806 = (inp[10]) ? 4'b1101 : 4'b0101;
											assign node12809 = (inp[13]) ? node12817 : node12810;
												assign node12810 = (inp[12]) ? 4'b1001 : node12811;
													assign node12811 = (inp[10]) ? node12813 : 4'b1001;
														assign node12813 = (inp[4]) ? 4'b0101 : 4'b0001;
												assign node12817 = (inp[4]) ? node12823 : node12818;
													assign node12818 = (inp[10]) ? node12820 : 4'b0001;
														assign node12820 = (inp[12]) ? 4'b0001 : 4'b1001;
													assign node12823 = (inp[2]) ? 4'b0101 : node12824;
														assign node12824 = (inp[12]) ? node12826 : 4'b0000;
															assign node12826 = (inp[10]) ? 4'b0000 : 4'b0101;
										assign node12830 = (inp[13]) ? node12860 : node12831;
											assign node12831 = (inp[2]) ? node12851 : node12832;
												assign node12832 = (inp[4]) ? node12838 : node12833;
													assign node12833 = (inp[7]) ? 4'b1000 : node12834;
														assign node12834 = (inp[12]) ? 4'b1000 : 4'b0100;
													assign node12838 = (inp[7]) ? node12846 : node12839;
														assign node12839 = (inp[14]) ? 4'b0000 : node12840;
															assign node12840 = (inp[10]) ? node12842 : 4'b1100;
																assign node12842 = (inp[12]) ? 4'b0000 : 4'b1000;
														assign node12846 = (inp[12]) ? node12848 : 4'b0100;
															assign node12848 = (inp[10]) ? 4'b0100 : 4'b1100;
												assign node12851 = (inp[12]) ? 4'b1101 : node12852;
													assign node12852 = (inp[7]) ? node12856 : node12853;
														assign node12853 = (inp[10]) ? 4'b1000 : 4'b0000;
														assign node12856 = (inp[10]) ? 4'b0101 : 4'b1101;
											assign node12860 = (inp[4]) ? node12878 : node12861;
												assign node12861 = (inp[2]) ? node12869 : node12862;
													assign node12862 = (inp[12]) ? node12864 : 4'b0100;
														assign node12864 = (inp[10]) ? 4'b0100 : node12865;
															assign node12865 = (inp[7]) ? 4'b1000 : 4'b1100;
													assign node12869 = (inp[7]) ? node12875 : node12870;
														assign node12870 = (inp[10]) ? node12872 : 4'b0001;
															assign node12872 = (inp[12]) ? 4'b0001 : 4'b1001;
														assign node12875 = (inp[10]) ? 4'b1101 : 4'b0101;
												assign node12878 = (inp[2]) ? node12884 : node12879;
													assign node12879 = (inp[10]) ? 4'b0001 : node12880;
														assign node12880 = (inp[7]) ? 4'b0000 : 4'b1001;
													assign node12884 = (inp[12]) ? node12888 : node12885;
														assign node12885 = (inp[10]) ? 4'b1000 : 4'b0000;
														assign node12888 = (inp[10]) ? 4'b0000 : node12889;
															assign node12889 = (inp[7]) ? 4'b0001 : 4'b1000;
									assign node12893 = (inp[13]) ? node12955 : node12894;
										assign node12894 = (inp[12]) ? node12920 : node12895;
											assign node12895 = (inp[7]) ? node12909 : node12896;
												assign node12896 = (inp[3]) ? node12902 : node12897;
													assign node12897 = (inp[14]) ? node12899 : 4'b0100;
														assign node12899 = (inp[2]) ? 4'b0100 : 4'b0000;
													assign node12902 = (inp[10]) ? 4'b1100 : node12903;
														assign node12903 = (inp[2]) ? 4'b0000 : node12904;
															assign node12904 = (inp[4]) ? 4'b0000 : 4'b0100;
												assign node12909 = (inp[4]) ? node12915 : node12910;
													assign node12910 = (inp[3]) ? node12912 : 4'b0000;
														assign node12912 = (inp[2]) ? 4'b0100 : 4'b1000;
													assign node12915 = (inp[10]) ? node12917 : 4'b0100;
														assign node12917 = (inp[3]) ? 4'b0000 : 4'b0100;
											assign node12920 = (inp[10]) ? node12940 : node12921;
												assign node12921 = (inp[3]) ? node12931 : node12922;
													assign node12922 = (inp[2]) ? node12928 : node12923;
														assign node12923 = (inp[14]) ? node12925 : 4'b1000;
															assign node12925 = (inp[7]) ? 4'b1000 : 4'b0000;
														assign node12928 = (inp[7]) ? 4'b1000 : 4'b1100;
													assign node12931 = (inp[2]) ? 4'b1100 : node12932;
														assign node12932 = (inp[4]) ? node12936 : node12933;
															assign node12933 = (inp[7]) ? 4'b0000 : 4'b0100;
															assign node12936 = (inp[7]) ? 4'b0100 : 4'b0000;
												assign node12940 = (inp[4]) ? node12946 : node12941;
													assign node12941 = (inp[3]) ? 4'b0100 : node12942;
														assign node12942 = (inp[7]) ? 4'b0000 : 4'b0100;
													assign node12946 = (inp[7]) ? node12952 : node12947;
														assign node12947 = (inp[14]) ? 4'b1000 : node12948;
															assign node12948 = (inp[3]) ? 4'b1000 : 4'b0100;
														assign node12952 = (inp[3]) ? 4'b1100 : 4'b0100;
										assign node12955 = (inp[10]) ? node12997 : node12956;
											assign node12956 = (inp[12]) ? node12978 : node12957;
												assign node12957 = (inp[4]) ? node12973 : node12958;
													assign node12958 = (inp[14]) ? node12966 : node12959;
														assign node12959 = (inp[3]) ? node12963 : node12960;
															assign node12960 = (inp[7]) ? 4'b1000 : 4'b1100;
															assign node12963 = (inp[7]) ? 4'b1100 : 4'b1000;
														assign node12966 = (inp[2]) ? node12970 : node12967;
															assign node12967 = (inp[7]) ? 4'b0100 : 4'b1100;
															assign node12970 = (inp[3]) ? 4'b1100 : 4'b1000;
													assign node12973 = (inp[2]) ? node12975 : 4'b0000;
														assign node12975 = (inp[3]) ? 4'b0000 : 4'b1100;
												assign node12978 = (inp[14]) ? node12992 : node12979;
													assign node12979 = (inp[7]) ? node12985 : node12980;
														assign node12980 = (inp[3]) ? 4'b0000 : node12981;
															assign node12981 = (inp[2]) ? 4'b0100 : 4'b0000;
														assign node12985 = (inp[3]) ? 4'b0100 : node12986;
															assign node12986 = (inp[2]) ? node12988 : 4'b0000;
																assign node12988 = (inp[4]) ? 4'b0100 : 4'b0000;
													assign node12992 = (inp[7]) ? 4'b0000 : node12993;
														assign node12993 = (inp[3]) ? 4'b0000 : 4'b0100;
											assign node12997 = (inp[2]) ? node13003 : node12998;
												assign node12998 = (inp[4]) ? 4'b1000 : node12999;
													assign node12999 = (inp[12]) ? 4'b1100 : 4'b1000;
												assign node13003 = (inp[3]) ? node13009 : node13004;
													assign node13004 = (inp[4]) ? 4'b1100 : node13005;
														assign node13005 = (inp[7]) ? 4'b1000 : 4'b1100;
													assign node13009 = (inp[4]) ? 4'b1000 : node13010;
														assign node13010 = (inp[7]) ? 4'b1100 : 4'b1000;
							assign node13014 = (inp[3]) ? node13310 : node13015;
								assign node13015 = (inp[4]) ? node13165 : node13016;
									assign node13016 = (inp[11]) ? node13096 : node13017;
										assign node13017 = (inp[2]) ? node13067 : node13018;
											assign node13018 = (inp[13]) ? node13046 : node13019;
												assign node13019 = (inp[7]) ? node13031 : node13020;
													assign node13020 = (inp[12]) ? node13022 : 4'b0100;
														assign node13022 = (inp[10]) ? node13028 : node13023;
															assign node13023 = (inp[1]) ? 4'b0100 : node13024;
																assign node13024 = (inp[14]) ? 4'b1001 : 4'b1000;
															assign node13028 = (inp[14]) ? 4'b0101 : 4'b1101;
													assign node13031 = (inp[1]) ? node13037 : node13032;
														assign node13032 = (inp[10]) ? node13034 : 4'b1001;
															assign node13034 = (inp[12]) ? 4'b0001 : 4'b1001;
														assign node13037 = (inp[14]) ? node13043 : node13038;
															assign node13038 = (inp[12]) ? node13040 : 4'b0101;
																assign node13040 = (inp[10]) ? 4'b1001 : 4'b0001;
															assign node13043 = (inp[12]) ? 4'b1000 : 4'b0000;
												assign node13046 = (inp[12]) ? node13060 : node13047;
													assign node13047 = (inp[1]) ? node13053 : node13048;
														assign node13048 = (inp[7]) ? node13050 : 4'b0000;
															assign node13050 = (inp[10]) ? 4'b0000 : 4'b1100;
														assign node13053 = (inp[10]) ? 4'b1000 : node13054;
															assign node13054 = (inp[14]) ? node13056 : 4'b1101;
																assign node13056 = (inp[7]) ? 4'b1100 : 4'b1000;
													assign node13060 = (inp[1]) ? 4'b0000 : node13061;
														assign node13061 = (inp[14]) ? 4'b0101 : node13062;
															assign node13062 = (inp[7]) ? 4'b0100 : 4'b1000;
											assign node13067 = (inp[10]) ? node13081 : node13068;
												assign node13068 = (inp[12]) ? node13076 : node13069;
													assign node13069 = (inp[1]) ? 4'b0101 : node13070;
														assign node13070 = (inp[7]) ? 4'b1001 : node13071;
															assign node13071 = (inp[13]) ? 4'b1101 : 4'b1001;
													assign node13076 = (inp[13]) ? node13078 : 4'b1001;
														assign node13078 = (inp[7]) ? 4'b1001 : 4'b1101;
												assign node13081 = (inp[12]) ? 4'b0101 : node13082;
													assign node13082 = (inp[1]) ? node13090 : node13083;
														assign node13083 = (inp[14]) ? 4'b0001 : node13084;
															assign node13084 = (inp[13]) ? node13086 : 4'b0101;
																assign node13086 = (inp[7]) ? 4'b0101 : 4'b0000;
														assign node13090 = (inp[13]) ? 4'b1000 : node13091;
															assign node13091 = (inp[7]) ? 4'b1001 : 4'b1101;
										assign node13096 = (inp[1]) ? node13136 : node13097;
											assign node13097 = (inp[2]) ? node13111 : node13098;
												assign node13098 = (inp[13]) ? node13106 : node13099;
													assign node13099 = (inp[12]) ? 4'b1001 : node13100;
														assign node13100 = (inp[7]) ? 4'b0001 : node13101;
															assign node13101 = (inp[10]) ? 4'b1101 : 4'b0101;
													assign node13106 = (inp[10]) ? 4'b0000 : node13107;
														assign node13107 = (inp[7]) ? 4'b1101 : 4'b0000;
												assign node13111 = (inp[13]) ? node13129 : node13112;
													assign node13112 = (inp[7]) ? node13124 : node13113;
														assign node13113 = (inp[14]) ? node13119 : node13114;
															assign node13114 = (inp[12]) ? 4'b0100 : node13115;
																assign node13115 = (inp[10]) ? 4'b1100 : 4'b0100;
															assign node13119 = (inp[10]) ? 4'b0100 : node13120;
																assign node13120 = (inp[12]) ? 4'b1000 : 4'b0100;
														assign node13124 = (inp[14]) ? node13126 : 4'b0000;
															assign node13126 = (inp[12]) ? 4'b1000 : 4'b0000;
													assign node13129 = (inp[10]) ? node13131 : 4'b1100;
														assign node13131 = (inp[7]) ? node13133 : 4'b0001;
															assign node13133 = (inp[12]) ? 4'b0100 : 4'b1100;
											assign node13136 = (inp[10]) ? node13154 : node13137;
												assign node13137 = (inp[2]) ? node13151 : node13138;
													assign node13138 = (inp[12]) ? node13146 : node13139;
														assign node13139 = (inp[7]) ? node13143 : node13140;
															assign node13140 = (inp[13]) ? 4'b1000 : 4'b1100;
															assign node13143 = (inp[13]) ? 4'b0100 : 4'b1000;
														assign node13146 = (inp[13]) ? 4'b1100 : node13147;
															assign node13147 = (inp[7]) ? 4'b0000 : 4'b0100;
													assign node13151 = (inp[13]) ? 4'b0100 : 4'b0000;
												assign node13154 = (inp[13]) ? node13160 : node13155;
													assign node13155 = (inp[2]) ? node13157 : 4'b0100;
														assign node13157 = (inp[7]) ? 4'b1000 : 4'b1100;
													assign node13160 = (inp[2]) ? node13162 : 4'b1000;
														assign node13162 = (inp[7]) ? 4'b1100 : 4'b1000;
									assign node13165 = (inp[1]) ? node13241 : node13166;
										assign node13166 = (inp[2]) ? node13208 : node13167;
											assign node13167 = (inp[13]) ? node13189 : node13168;
												assign node13168 = (inp[12]) ? node13178 : node13169;
													assign node13169 = (inp[7]) ? node13175 : node13170;
														assign node13170 = (inp[10]) ? node13172 : 4'b0100;
															assign node13172 = (inp[14]) ? 4'b0000 : 4'b1001;
														assign node13175 = (inp[10]) ? 4'b0100 : 4'b0000;
													assign node13178 = (inp[7]) ? node13184 : node13179;
														assign node13179 = (inp[14]) ? node13181 : 4'b0001;
															assign node13181 = (inp[11]) ? 4'b0001 : 4'b0000;
														assign node13184 = (inp[11]) ? node13186 : 4'b1000;
															assign node13186 = (inp[14]) ? 4'b0100 : 4'b0000;
												assign node13189 = (inp[14]) ? node13199 : node13190;
													assign node13190 = (inp[11]) ? node13194 : node13191;
														assign node13191 = (inp[12]) ? 4'b0001 : 4'b1001;
														assign node13194 = (inp[10]) ? node13196 : 4'b1001;
															assign node13196 = (inp[12]) ? 4'b1001 : 4'b0000;
													assign node13199 = (inp[11]) ? node13205 : node13200;
														assign node13200 = (inp[12]) ? node13202 : 4'b1000;
															assign node13202 = (inp[10]) ? 4'b0001 : 4'b0000;
														assign node13205 = (inp[10]) ? 4'b1000 : 4'b1001;
											assign node13208 = (inp[13]) ? node13228 : node13209;
												assign node13209 = (inp[11]) ? node13223 : node13210;
													assign node13210 = (inp[14]) ? node13218 : node13211;
														assign node13211 = (inp[12]) ? node13215 : node13212;
															assign node13212 = (inp[10]) ? 4'b1000 : 4'b0000;
															assign node13215 = (inp[7]) ? 4'b1101 : 4'b1000;
														assign node13218 = (inp[12]) ? node13220 : 4'b1001;
															assign node13220 = (inp[10]) ? 4'b0001 : 4'b1001;
													assign node13223 = (inp[10]) ? 4'b1001 : node13224;
														assign node13224 = (inp[12]) ? 4'b1001 : 4'b0001;
												assign node13228 = (inp[10]) ? node13232 : node13229;
													assign node13229 = (inp[7]) ? 4'b0001 : 4'b0100;
													assign node13232 = (inp[11]) ? 4'b0000 : node13233;
														assign node13233 = (inp[14]) ? 4'b1001 : node13234;
															assign node13234 = (inp[7]) ? 4'b0100 : node13235;
																assign node13235 = (inp[12]) ? 4'b1000 : 4'b0000;
										assign node13241 = (inp[11]) ? node13281 : node13242;
											assign node13242 = (inp[2]) ? node13264 : node13243;
												assign node13243 = (inp[13]) ? node13257 : node13244;
													assign node13244 = (inp[12]) ? node13252 : node13245;
														assign node13245 = (inp[10]) ? node13249 : node13246;
															assign node13246 = (inp[7]) ? 4'b1000 : 4'b1100;
															assign node13249 = (inp[7]) ? 4'b1100 : 4'b1001;
														assign node13252 = (inp[14]) ? node13254 : 4'b0100;
															assign node13254 = (inp[7]) ? 4'b0100 : 4'b1001;
													assign node13257 = (inp[10]) ? 4'b0001 : node13258;
														assign node13258 = (inp[14]) ? 4'b1001 : node13259;
															assign node13259 = (inp[7]) ? 4'b0000 : 4'b0100;
												assign node13264 = (inp[14]) ? node13274 : node13265;
													assign node13265 = (inp[13]) ? node13267 : 4'b0001;
														assign node13267 = (inp[12]) ? 4'b0000 : node13268;
															assign node13268 = (inp[7]) ? node13270 : 4'b1000;
																assign node13270 = (inp[10]) ? 4'b1000 : 4'b1001;
													assign node13274 = (inp[10]) ? node13276 : 4'b0000;
														assign node13276 = (inp[13]) ? 4'b0000 : node13277;
															assign node13277 = (inp[12]) ? 4'b1000 : 4'b0000;
											assign node13281 = (inp[13]) ? node13297 : node13282;
												assign node13282 = (inp[7]) ? node13290 : node13283;
													assign node13283 = (inp[10]) ? 4'b0100 : node13284;
														assign node13284 = (inp[2]) ? 4'b0000 : node13285;
															assign node13285 = (inp[12]) ? 4'b1100 : 4'b0000;
													assign node13290 = (inp[10]) ? 4'b0000 : node13291;
														assign node13291 = (inp[2]) ? node13293 : 4'b1000;
															assign node13293 = (inp[12]) ? 4'b0000 : 4'b1000;
												assign node13297 = (inp[10]) ? 4'b1000 : node13298;
													assign node13298 = (inp[2]) ? node13304 : node13299;
														assign node13299 = (inp[12]) ? 4'b0000 : node13300;
															assign node13300 = (inp[7]) ? 4'b1000 : 4'b0000;
														assign node13304 = (inp[12]) ? 4'b1000 : node13305;
															assign node13305 = (inp[7]) ? 4'b0100 : 4'b1000;
								assign node13310 = (inp[4]) ? node13460 : node13311;
									assign node13311 = (inp[1]) ? node13395 : node13312;
										assign node13312 = (inp[7]) ? node13360 : node13313;
											assign node13313 = (inp[10]) ? node13339 : node13314;
												assign node13314 = (inp[11]) ? node13330 : node13315;
													assign node13315 = (inp[12]) ? node13323 : node13316;
														assign node13316 = (inp[13]) ? node13318 : 4'b0000;
															assign node13318 = (inp[2]) ? 4'b0001 : node13319;
																assign node13319 = (inp[14]) ? 4'b1000 : 4'b1001;
														assign node13323 = (inp[13]) ? node13327 : node13324;
															assign node13324 = (inp[2]) ? 4'b1000 : 4'b1001;
															assign node13327 = (inp[14]) ? 4'b1000 : 4'b1001;
													assign node13330 = (inp[2]) ? node13334 : node13331;
														assign node13331 = (inp[13]) ? 4'b0000 : 4'b1001;
														assign node13334 = (inp[13]) ? node13336 : 4'b0001;
															assign node13336 = (inp[12]) ? 4'b0000 : 4'b0001;
												assign node13339 = (inp[11]) ? node13353 : node13340;
													assign node13340 = (inp[12]) ? node13348 : node13341;
														assign node13341 = (inp[2]) ? node13345 : node13342;
															assign node13342 = (inp[14]) ? 4'b1001 : 4'b0000;
															assign node13345 = (inp[13]) ? 4'b0000 : 4'b0001;
														assign node13348 = (inp[14]) ? 4'b0000 : node13349;
															assign node13349 = (inp[2]) ? 4'b0001 : 4'b0000;
													assign node13353 = (inp[2]) ? node13357 : node13354;
														assign node13354 = (inp[13]) ? 4'b0000 : 4'b1000;
														assign node13357 = (inp[13]) ? 4'b1000 : 4'b0000;
											assign node13360 = (inp[10]) ? node13380 : node13361;
												assign node13361 = (inp[13]) ? node13371 : node13362;
													assign node13362 = (inp[2]) ? node13366 : node13363;
														assign node13363 = (inp[11]) ? 4'b1000 : 4'b1001;
														assign node13366 = (inp[11]) ? 4'b0000 : node13367;
															assign node13367 = (inp[12]) ? 4'b1000 : 4'b0000;
													assign node13371 = (inp[12]) ? 4'b0000 : node13372;
														assign node13372 = (inp[2]) ? node13376 : node13373;
															assign node13373 = (inp[11]) ? 4'b0001 : 4'b0000;
															assign node13376 = (inp[11]) ? 4'b1000 : 4'b0001;
												assign node13380 = (inp[13]) ? node13388 : node13381;
													assign node13381 = (inp[11]) ? 4'b0001 : node13382;
														assign node13382 = (inp[14]) ? 4'b0000 : node13383;
															assign node13383 = (inp[2]) ? 4'b0001 : 4'b0000;
													assign node13388 = (inp[2]) ? node13392 : node13389;
														assign node13389 = (inp[11]) ? 4'b0001 : 4'b1001;
														assign node13392 = (inp[11]) ? 4'b1001 : 4'b0001;
										assign node13395 = (inp[11]) ? node13431 : node13396;
											assign node13396 = (inp[10]) ? node13422 : node13397;
												assign node13397 = (inp[13]) ? node13409 : node13398;
													assign node13398 = (inp[14]) ? node13402 : node13399;
														assign node13399 = (inp[2]) ? 4'b1000 : 4'b1001;
														assign node13402 = (inp[12]) ? node13406 : node13403;
															assign node13403 = (inp[2]) ? 4'b1000 : 4'b0000;
															assign node13406 = (inp[2]) ? 4'b0000 : 4'b1001;
													assign node13409 = (inp[12]) ? node13417 : node13410;
														assign node13410 = (inp[7]) ? node13412 : 4'b1001;
															assign node13412 = (inp[2]) ? 4'b1001 : node13413;
																assign node13413 = (inp[14]) ? 4'b1001 : 4'b0000;
														assign node13417 = (inp[7]) ? 4'b1001 : node13418;
															assign node13418 = (inp[14]) ? 4'b0000 : 4'b0001;
												assign node13422 = (inp[2]) ? node13428 : node13423;
													assign node13423 = (inp[14]) ? node13425 : 4'b0000;
														assign node13425 = (inp[13]) ? 4'b1000 : 4'b0000;
													assign node13428 = (inp[12]) ? 4'b0000 : 4'b0001;
											assign node13431 = (inp[7]) ? node13447 : node13432;
												assign node13432 = (inp[2]) ? node13442 : node13433;
													assign node13433 = (inp[12]) ? 4'b0000 : node13434;
														assign node13434 = (inp[10]) ? node13438 : node13435;
															assign node13435 = (inp[13]) ? 4'b0000 : 4'b1000;
															assign node13438 = (inp[13]) ? 4'b1000 : 4'b0000;
													assign node13442 = (inp[10]) ? 4'b1000 : node13443;
														assign node13443 = (inp[12]) ? 4'b1000 : 4'b0000;
												assign node13447 = (inp[2]) ? node13453 : node13448;
													assign node13448 = (inp[12]) ? node13450 : 4'b1000;
														assign node13450 = (inp[10]) ? 4'b1000 : 4'b0000;
													assign node13453 = (inp[10]) ? node13457 : node13454;
														assign node13454 = (inp[12]) ? 4'b1000 : 4'b0000;
														assign node13457 = (inp[13]) ? 4'b1000 : 4'b0000;
									assign node13460 = (inp[13]) ? node13534 : node13461;
										assign node13461 = (inp[1]) ? node13507 : node13462;
											assign node13462 = (inp[7]) ? node13480 : node13463;
												assign node13463 = (inp[2]) ? node13467 : node13464;
													assign node13464 = (inp[12]) ? 4'b0001 : 4'b1001;
													assign node13467 = (inp[12]) ? node13469 : 4'b0001;
														assign node13469 = (inp[14]) ? node13475 : node13470;
															assign node13470 = (inp[10]) ? node13472 : 4'b1000;
																assign node13472 = (inp[11]) ? 4'b0001 : 4'b1001;
															assign node13475 = (inp[10]) ? 4'b1000 : node13476;
																assign node13476 = (inp[11]) ? 4'b1000 : 4'b0001;
												assign node13480 = (inp[10]) ? node13490 : node13481;
													assign node13481 = (inp[14]) ? node13487 : node13482;
														assign node13482 = (inp[11]) ? 4'b0000 : node13483;
															assign node13483 = (inp[2]) ? 4'b0001 : 4'b1001;
														assign node13487 = (inp[12]) ? 4'b1001 : 4'b1000;
													assign node13490 = (inp[14]) ? node13498 : node13491;
														assign node13491 = (inp[2]) ? node13495 : node13492;
															assign node13492 = (inp[12]) ? 4'b0000 : 4'b0001;
															assign node13495 = (inp[11]) ? 4'b0001 : 4'b1000;
														assign node13498 = (inp[11]) ? node13502 : node13499;
															assign node13499 = (inp[2]) ? 4'b0000 : 4'b0001;
															assign node13502 = (inp[2]) ? node13504 : 4'b0000;
																assign node13504 = (inp[12]) ? 4'b0001 : 4'b0000;
											assign node13507 = (inp[10]) ? node13525 : node13508;
												assign node13508 = (inp[14]) ? node13514 : node13509;
													assign node13509 = (inp[12]) ? node13511 : 4'b0000;
														assign node13511 = (inp[2]) ? 4'b1001 : 4'b1000;
													assign node13514 = (inp[12]) ? node13516 : 4'b1000;
														assign node13516 = (inp[2]) ? 4'b1000 : node13517;
															assign node13517 = (inp[7]) ? node13521 : node13518;
																assign node13518 = (inp[11]) ? 4'b0000 : 4'b1000;
																assign node13521 = (inp[11]) ? 4'b1000 : 4'b0000;
												assign node13525 = (inp[11]) ? 4'b0000 : node13526;
													assign node13526 = (inp[7]) ? node13528 : 4'b0000;
														assign node13528 = (inp[2]) ? node13530 : 4'b0001;
															assign node13530 = (inp[14]) ? 4'b0000 : 4'b0001;
										assign node13534 = (inp[1]) ? node13556 : node13535;
											assign node13535 = (inp[7]) ? node13547 : node13536;
												assign node13536 = (inp[11]) ? 4'b0000 : node13537;
													assign node13537 = (inp[14]) ? node13539 : 4'b0000;
														assign node13539 = (inp[10]) ? node13543 : node13540;
															assign node13540 = (inp[12]) ? 4'b0000 : 4'b0001;
															assign node13543 = (inp[12]) ? 4'b0001 : 4'b0000;
												assign node13547 = (inp[11]) ? node13553 : node13548;
													assign node13548 = (inp[10]) ? node13550 : 4'b0000;
														assign node13550 = (inp[14]) ? 4'b0001 : 4'b0000;
													assign node13553 = (inp[10]) ? 4'b0000 : 4'b0001;
											assign node13556 = (inp[10]) ? 4'b0000 : node13557;
												assign node13557 = (inp[11]) ? 4'b0000 : node13558;
													assign node13558 = (inp[7]) ? 4'b0000 : node13559;
														assign node13559 = (inp[14]) ? node13561 : 4'b0001;
															assign node13561 = (inp[12]) ? 4'b0001 : 4'b0000;
					assign node13567 = (inp[6]) ? node13569 : 4'b1000;
						assign node13569 = (inp[5]) ? node13673 : node13570;
							assign node13570 = (inp[3]) ? node13572 : 4'b1000;
								assign node13572 = (inp[2]) ? 4'b1000 : node13573;
									assign node13573 = (inp[1]) ? node13615 : node13574;
										assign node13574 = (inp[4]) ? node13588 : node13575;
											assign node13575 = (inp[7]) ? 4'b1000 : node13576;
												assign node13576 = (inp[13]) ? node13582 : node13577;
													assign node13577 = (inp[10]) ? node13579 : 4'b1000;
														assign node13579 = (inp[12]) ? 4'b1000 : 4'b0001;
													assign node13582 = (inp[11]) ? 4'b0001 : node13583;
														assign node13583 = (inp[12]) ? 4'b0000 : 4'b0001;
											assign node13588 = (inp[13]) ? node13604 : node13589;
												assign node13589 = (inp[11]) ? node13597 : node13590;
													assign node13590 = (inp[14]) ? node13592 : 4'b0001;
														assign node13592 = (inp[12]) ? 4'b1000 : node13593;
															assign node13593 = (inp[10]) ? 4'b0000 : 4'b1000;
													assign node13597 = (inp[7]) ? 4'b1000 : node13598;
														assign node13598 = (inp[12]) ? 4'b1001 : node13599;
															assign node13599 = (inp[10]) ? 4'b0001 : 4'b1001;
												assign node13604 = (inp[10]) ? node13610 : node13605;
													assign node13605 = (inp[14]) ? node13607 : 4'b0001;
														assign node13607 = (inp[11]) ? 4'b0001 : 4'b0000;
													assign node13610 = (inp[12]) ? node13612 : 4'b1001;
														assign node13612 = (inp[14]) ? 4'b0000 : 4'b0001;
										assign node13615 = (inp[14]) ? node13637 : node13616;
											assign node13616 = (inp[13]) ? node13628 : node13617;
												assign node13617 = (inp[10]) ? node13623 : node13618;
													assign node13618 = (inp[7]) ? 4'b1000 : node13619;
														assign node13619 = (inp[4]) ? 4'b1000 : 4'b0000;
													assign node13623 = (inp[4]) ? 4'b0000 : node13624;
														assign node13624 = (inp[7]) ? 4'b1000 : 4'b0000;
												assign node13628 = (inp[10]) ? 4'b1000 : node13629;
													assign node13629 = (inp[12]) ? node13631 : 4'b1000;
														assign node13631 = (inp[4]) ? 4'b0000 : node13632;
															assign node13632 = (inp[7]) ? 4'b1000 : 4'b0000;
											assign node13637 = (inp[11]) ? node13657 : node13638;
												assign node13638 = (inp[4]) ? node13648 : node13639;
													assign node13639 = (inp[7]) ? 4'b1000 : node13640;
														assign node13640 = (inp[13]) ? 4'b0001 : node13641;
															assign node13641 = (inp[12]) ? 4'b1000 : node13642;
																assign node13642 = (inp[10]) ? 4'b0001 : 4'b1000;
													assign node13648 = (inp[12]) ? 4'b1001 : node13649;
														assign node13649 = (inp[10]) ? node13653 : node13650;
															assign node13650 = (inp[13]) ? 4'b0001 : 4'b1000;
															assign node13653 = (inp[13]) ? 4'b1001 : 4'b0001;
												assign node13657 = (inp[12]) ? node13663 : node13658;
													assign node13658 = (inp[13]) ? 4'b1000 : node13659;
														assign node13659 = (inp[7]) ? 4'b1000 : 4'b0000;
													assign node13663 = (inp[4]) ? node13665 : 4'b1000;
														assign node13665 = (inp[10]) ? node13669 : node13666;
															assign node13666 = (inp[13]) ? 4'b0000 : 4'b1000;
															assign node13669 = (inp[13]) ? 4'b1000 : 4'b0000;
							assign node13673 = (inp[2]) ? node13957 : node13674;
								assign node13674 = (inp[3]) ? node13838 : node13675;
									assign node13675 = (inp[1]) ? node13759 : node13676;
										assign node13676 = (inp[13]) ? node13728 : node13677;
											assign node13677 = (inp[10]) ? node13701 : node13678;
												assign node13678 = (inp[14]) ? node13690 : node13679;
													assign node13679 = (inp[11]) ? node13685 : node13680;
														assign node13680 = (inp[7]) ? 4'b1001 : node13681;
															assign node13681 = (inp[4]) ? 4'b1101 : 4'b1001;
														assign node13685 = (inp[4]) ? node13687 : 4'b1001;
															assign node13687 = (inp[7]) ? 4'b1001 : 4'b0000;
													assign node13690 = (inp[11]) ? node13696 : node13691;
														assign node13691 = (inp[7]) ? 4'b1000 : node13692;
															assign node13692 = (inp[4]) ? 4'b1100 : 4'b1000;
														assign node13696 = (inp[7]) ? 4'b1001 : node13697;
															assign node13697 = (inp[4]) ? 4'b0000 : 4'b1001;
												assign node13701 = (inp[12]) ? node13719 : node13702;
													assign node13702 = (inp[4]) ? node13710 : node13703;
														assign node13703 = (inp[7]) ? node13705 : 4'b0101;
															assign node13705 = (inp[14]) ? node13707 : 4'b0001;
																assign node13707 = (inp[11]) ? 4'b0001 : 4'b0000;
														assign node13710 = (inp[7]) ? node13714 : node13711;
															assign node13711 = (inp[11]) ? 4'b1000 : 4'b0001;
															assign node13714 = (inp[11]) ? 4'b0101 : node13715;
																assign node13715 = (inp[14]) ? 4'b0100 : 4'b0101;
													assign node13719 = (inp[4]) ? node13725 : node13720;
														assign node13720 = (inp[11]) ? 4'b1001 : node13721;
															assign node13721 = (inp[14]) ? 4'b1000 : 4'b1001;
														assign node13725 = (inp[11]) ? 4'b1001 : 4'b0001;
											assign node13728 = (inp[4]) ? node13740 : node13729;
												assign node13729 = (inp[7]) ? node13733 : node13730;
													assign node13730 = (inp[12]) ? 4'b0101 : 4'b1101;
													assign node13733 = (inp[12]) ? node13737 : node13734;
														assign node13734 = (inp[10]) ? 4'b1001 : 4'b0001;
														assign node13737 = (inp[11]) ? 4'b0001 : 4'b0000;
												assign node13740 = (inp[11]) ? node13750 : node13741;
													assign node13741 = (inp[7]) ? node13745 : node13742;
														assign node13742 = (inp[10]) ? 4'b0001 : 4'b1001;
														assign node13745 = (inp[12]) ? node13747 : 4'b0100;
															assign node13747 = (inp[10]) ? 4'b0001 : 4'b0101;
													assign node13750 = (inp[12]) ? node13754 : node13751;
														assign node13751 = (inp[10]) ? 4'b1000 : 4'b0000;
														assign node13754 = (inp[10]) ? 4'b0000 : node13755;
															assign node13755 = (inp[7]) ? 4'b0101 : 4'b1000;
										assign node13759 = (inp[11]) ? node13805 : node13760;
											assign node13760 = (inp[14]) ? node13782 : node13761;
												assign node13761 = (inp[4]) ? node13771 : node13762;
													assign node13762 = (inp[7]) ? node13768 : node13763;
														assign node13763 = (inp[12]) ? 4'b0100 : node13764;
															assign node13764 = (inp[13]) ? 4'b1100 : 4'b0100;
														assign node13768 = (inp[13]) ? 4'b1000 : 4'b0000;
													assign node13771 = (inp[10]) ? node13779 : node13772;
														assign node13772 = (inp[12]) ? node13774 : 4'b0001;
															assign node13774 = (inp[13]) ? 4'b0100 : node13775;
																assign node13775 = (inp[7]) ? 4'b1000 : 4'b1100;
														assign node13779 = (inp[12]) ? 4'b0001 : 4'b1001;
												assign node13782 = (inp[13]) ? node13790 : node13783;
													assign node13783 = (inp[12]) ? 4'b1001 : node13784;
														assign node13784 = (inp[10]) ? node13786 : 4'b1001;
															assign node13786 = (inp[4]) ? 4'b0101 : 4'b0001;
													assign node13790 = (inp[4]) ? node13798 : node13791;
														assign node13791 = (inp[7]) ? 4'b0001 : node13792;
															assign node13792 = (inp[12]) ? 4'b0101 : node13793;
																assign node13793 = (inp[10]) ? 4'b1101 : 4'b0101;
														assign node13798 = (inp[7]) ? node13800 : 4'b1001;
															assign node13800 = (inp[10]) ? node13802 : 4'b0101;
																assign node13802 = (inp[12]) ? 4'b0001 : 4'b1001;
											assign node13805 = (inp[4]) ? node13825 : node13806;
												assign node13806 = (inp[7]) ? node13818 : node13807;
													assign node13807 = (inp[13]) ? node13813 : node13808;
														assign node13808 = (inp[10]) ? 4'b0100 : node13809;
															assign node13809 = (inp[12]) ? 4'b1000 : 4'b0100;
														assign node13813 = (inp[10]) ? 4'b1100 : node13814;
															assign node13814 = (inp[12]) ? 4'b0100 : 4'b1100;
													assign node13818 = (inp[13]) ? node13820 : 4'b0000;
														assign node13820 = (inp[14]) ? node13822 : 4'b1000;
															assign node13822 = (inp[12]) ? 4'b0000 : 4'b1000;
												assign node13825 = (inp[10]) ? node13833 : node13826;
													assign node13826 = (inp[13]) ? 4'b0000 : node13827;
														assign node13827 = (inp[12]) ? 4'b1000 : node13828;
															assign node13828 = (inp[14]) ? 4'b0000 : 4'b0100;
													assign node13833 = (inp[7]) ? node13835 : 4'b1000;
														assign node13835 = (inp[13]) ? 4'b1000 : 4'b0100;
									assign node13838 = (inp[11]) ? node13916 : node13839;
										assign node13839 = (inp[10]) ? node13881 : node13840;
											assign node13840 = (inp[13]) ? node13858 : node13841;
												assign node13841 = (inp[1]) ? node13849 : node13842;
													assign node13842 = (inp[4]) ? node13844 : 4'b1001;
														assign node13844 = (inp[12]) ? node13846 : 4'b0001;
															assign node13846 = (inp[14]) ? 4'b1000 : 4'b1001;
													assign node13849 = (inp[4]) ? node13851 : 4'b0001;
														assign node13851 = (inp[12]) ? node13855 : node13852;
															assign node13852 = (inp[14]) ? 4'b1001 : 4'b1000;
															assign node13855 = (inp[14]) ? 4'b0001 : 4'b1001;
												assign node13858 = (inp[4]) ? node13868 : node13859;
													assign node13859 = (inp[1]) ? node13863 : node13860;
														assign node13860 = (inp[12]) ? 4'b0001 : 4'b0000;
														assign node13863 = (inp[7]) ? node13865 : 4'b1000;
															assign node13865 = (inp[12]) ? 4'b1000 : 4'b1001;
													assign node13868 = (inp[7]) ? node13876 : node13869;
														assign node13869 = (inp[12]) ? node13871 : 4'b0001;
															assign node13871 = (inp[14]) ? node13873 : 4'b0000;
																assign node13873 = (inp[1]) ? 4'b0001 : 4'b0000;
														assign node13876 = (inp[12]) ? 4'b0001 : node13877;
															assign node13877 = (inp[14]) ? 4'b0000 : 4'b0001;
											assign node13881 = (inp[4]) ? node13899 : node13882;
												assign node13882 = (inp[13]) ? node13890 : node13883;
													assign node13883 = (inp[7]) ? 4'b0001 : node13884;
														assign node13884 = (inp[1]) ? node13886 : 4'b1001;
															assign node13886 = (inp[12]) ? 4'b1001 : 4'b0000;
													assign node13890 = (inp[12]) ? 4'b1000 : node13891;
														assign node13891 = (inp[1]) ? node13893 : 4'b0000;
															assign node13893 = (inp[7]) ? 4'b1000 : node13894;
																assign node13894 = (inp[14]) ? 4'b0001 : 4'b1000;
												assign node13899 = (inp[13]) ? node13911 : node13900;
													assign node13900 = (inp[7]) ? node13904 : node13901;
														assign node13901 = (inp[1]) ? 4'b0001 : 4'b0000;
														assign node13904 = (inp[1]) ? 4'b0000 : node13905;
															assign node13905 = (inp[14]) ? 4'b1001 : node13906;
																assign node13906 = (inp[12]) ? 4'b0001 : 4'b0000;
													assign node13911 = (inp[12]) ? 4'b0000 : node13912;
														assign node13912 = (inp[1]) ? 4'b0000 : 4'b0001;
										assign node13916 = (inp[4]) ? node13944 : node13917;
											assign node13917 = (inp[1]) ? node13931 : node13918;
												assign node13918 = (inp[13]) ? node13924 : node13919;
													assign node13919 = (inp[14]) ? node13921 : 4'b1001;
														assign node13921 = (inp[12]) ? 4'b0000 : 4'b1000;
													assign node13924 = (inp[12]) ? 4'b0000 : node13925;
														assign node13925 = (inp[7]) ? 4'b1001 : node13926;
															assign node13926 = (inp[10]) ? 4'b0001 : 4'b0000;
												assign node13931 = (inp[13]) ? node13937 : node13932;
													assign node13932 = (inp[10]) ? 4'b0000 : node13933;
														assign node13933 = (inp[7]) ? 4'b0000 : 4'b1000;
													assign node13937 = (inp[7]) ? node13939 : 4'b1000;
														assign node13939 = (inp[10]) ? 4'b1000 : node13940;
															assign node13940 = (inp[12]) ? 4'b1000 : 4'b0000;
											assign node13944 = (inp[13]) ? 4'b0000 : node13945;
												assign node13945 = (inp[7]) ? node13953 : node13946;
													assign node13946 = (inp[12]) ? node13948 : 4'b1000;
														assign node13948 = (inp[14]) ? 4'b0000 : node13949;
															assign node13949 = (inp[1]) ? 4'b0000 : 4'b1000;
													assign node13953 = (inp[1]) ? 4'b0000 : 4'b0001;
								assign node13957 = (inp[3]) ? node13959 : 4'b1000;
									assign node13959 = (inp[4]) ? node14001 : node13960;
										assign node13960 = (inp[7]) ? 4'b1000 : node13961;
											assign node13961 = (inp[13]) ? node13977 : node13962;
												assign node13962 = (inp[12]) ? node13972 : node13963;
													assign node13963 = (inp[10]) ? node13967 : node13964;
														assign node13964 = (inp[1]) ? 4'b0000 : 4'b1000;
														assign node13967 = (inp[14]) ? 4'b0001 : node13968;
															assign node13968 = (inp[1]) ? 4'b0000 : 4'b0001;
													assign node13972 = (inp[1]) ? node13974 : 4'b1000;
														assign node13974 = (inp[14]) ? 4'b1000 : 4'b0000;
												assign node13977 = (inp[12]) ? node13991 : node13978;
													assign node13978 = (inp[14]) ? node13982 : node13979;
														assign node13979 = (inp[1]) ? 4'b1000 : 4'b1001;
														assign node13982 = (inp[10]) ? node13986 : node13983;
															assign node13983 = (inp[11]) ? 4'b1000 : 4'b0001;
															assign node13986 = (inp[11]) ? 4'b1001 : node13987;
																assign node13987 = (inp[1]) ? 4'b1001 : 4'b1000;
													assign node13991 = (inp[14]) ? node13993 : 4'b0001;
														assign node13993 = (inp[1]) ? node13997 : node13994;
															assign node13994 = (inp[11]) ? 4'b0001 : 4'b0000;
															assign node13997 = (inp[11]) ? 4'b0000 : 4'b0001;
										assign node14001 = (inp[13]) ? node14035 : node14002;
											assign node14002 = (inp[7]) ? node14022 : node14003;
												assign node14003 = (inp[11]) ? node14013 : node14004;
													assign node14004 = (inp[10]) ? 4'b0001 : node14005;
														assign node14005 = (inp[12]) ? 4'b1000 : node14006;
															assign node14006 = (inp[1]) ? 4'b0001 : node14007;
																assign node14007 = (inp[14]) ? 4'b1000 : 4'b1001;
													assign node14013 = (inp[1]) ? 4'b0000 : node14014;
														assign node14014 = (inp[12]) ? node14018 : node14015;
															assign node14015 = (inp[10]) ? 4'b1000 : 4'b0000;
															assign node14018 = (inp[10]) ? 4'b0000 : 4'b1001;
												assign node14022 = (inp[12]) ? 4'b1000 : node14023;
													assign node14023 = (inp[10]) ? node14027 : node14024;
														assign node14024 = (inp[1]) ? 4'b0000 : 4'b1000;
														assign node14027 = (inp[1]) ? 4'b0000 : node14028;
															assign node14028 = (inp[14]) ? node14030 : 4'b0001;
																assign node14030 = (inp[11]) ? 4'b0001 : 4'b0000;
											assign node14035 = (inp[10]) ? 4'b0000 : node14036;
												assign node14036 = (inp[11]) ? node14042 : node14037;
													assign node14037 = (inp[7]) ? 4'b0001 : node14038;
														assign node14038 = (inp[1]) ? 4'b0000 : 4'b0001;
													assign node14042 = (inp[12]) ? node14044 : 4'b0000;
														assign node14044 = (inp[1]) ? 4'b0000 : 4'b0001;
			assign node14048 = (inp[15]) ? node16498 : node14049;
				assign node14049 = (inp[6]) ? node14665 : node14050;
					assign node14050 = (inp[0]) ? 4'b0100 : node14051;
						assign node14051 = (inp[2]) ? node14445 : node14052;
							assign node14052 = (inp[3]) ? node14254 : node14053;
								assign node14053 = (inp[5]) ? node14129 : node14054;
									assign node14054 = (inp[4]) ? node14070 : node14055;
										assign node14055 = (inp[7]) ? 4'b0110 : node14056;
											assign node14056 = (inp[13]) ? node14058 : 4'b0110;
												assign node14058 = (inp[12]) ? node14064 : node14059;
													assign node14059 = (inp[1]) ? 4'b0000 : node14060;
														assign node14060 = (inp[10]) ? 4'b0001 : 4'b0110;
													assign node14064 = (inp[10]) ? node14066 : 4'b0110;
														assign node14066 = (inp[14]) ? 4'b0110 : 4'b0000;
										assign node14070 = (inp[7]) ? node14114 : node14071;
											assign node14071 = (inp[1]) ? node14089 : node14072;
												assign node14072 = (inp[13]) ? node14086 : node14073;
													assign node14073 = (inp[11]) ? node14081 : node14074;
														assign node14074 = (inp[14]) ? node14076 : 4'b0001;
															assign node14076 = (inp[10]) ? node14078 : 4'b0000;
																assign node14078 = (inp[12]) ? 4'b0000 : 4'b1000;
														assign node14081 = (inp[12]) ? 4'b0001 : node14082;
															assign node14082 = (inp[10]) ? 4'b1001 : 4'b0001;
													assign node14086 = (inp[12]) ? 4'b1001 : 4'b1000;
												assign node14089 = (inp[11]) ? node14103 : node14090;
													assign node14090 = (inp[14]) ? node14098 : node14091;
														assign node14091 = (inp[12]) ? node14093 : 4'b1000;
															assign node14093 = (inp[10]) ? 4'b0000 : node14094;
																assign node14094 = (inp[13]) ? 4'b1000 : 4'b0000;
														assign node14098 = (inp[10]) ? 4'b1001 : node14099;
															assign node14099 = (inp[13]) ? 4'b1001 : 4'b0001;
													assign node14103 = (inp[10]) ? node14111 : node14104;
														assign node14104 = (inp[14]) ? 4'b1000 : node14105;
															assign node14105 = (inp[12]) ? node14107 : 4'b1000;
																assign node14107 = (inp[13]) ? 4'b1000 : 4'b0000;
														assign node14111 = (inp[13]) ? 4'b0000 : 4'b1000;
											assign node14114 = (inp[12]) ? 4'b0110 : node14115;
												assign node14115 = (inp[13]) ? node14117 : 4'b0110;
													assign node14117 = (inp[10]) ? node14121 : node14118;
														assign node14118 = (inp[11]) ? 4'b0000 : 4'b0110;
														assign node14121 = (inp[1]) ? node14125 : node14122;
															assign node14122 = (inp[11]) ? 4'b0001 : 4'b0000;
															assign node14125 = (inp[11]) ? 4'b0000 : 4'b0001;
									assign node14129 = (inp[1]) ? node14197 : node14130;
										assign node14130 = (inp[13]) ? node14166 : node14131;
											assign node14131 = (inp[14]) ? node14145 : node14132;
												assign node14132 = (inp[4]) ? node14138 : node14133;
													assign node14133 = (inp[12]) ? 4'b0101 : node14134;
														assign node14134 = (inp[10]) ? 4'b1101 : 4'b0101;
													assign node14138 = (inp[7]) ? 4'b0101 : node14139;
														assign node14139 = (inp[10]) ? node14141 : 4'b0001;
															assign node14141 = (inp[12]) ? 4'b0001 : 4'b1001;
												assign node14145 = (inp[11]) ? node14157 : node14146;
													assign node14146 = (inp[4]) ? node14152 : node14147;
														assign node14147 = (inp[12]) ? 4'b0100 : node14148;
															assign node14148 = (inp[10]) ? 4'b1100 : 4'b0100;
														assign node14152 = (inp[7]) ? node14154 : 4'b0000;
															assign node14154 = (inp[10]) ? 4'b1100 : 4'b0100;
													assign node14157 = (inp[12]) ? node14161 : node14158;
														assign node14158 = (inp[10]) ? 4'b1101 : 4'b0101;
														assign node14161 = (inp[10]) ? 4'b0101 : node14162;
															assign node14162 = (inp[4]) ? 4'b0001 : 4'b0101;
											assign node14166 = (inp[4]) ? node14176 : node14167;
												assign node14167 = (inp[14]) ? node14169 : 4'b1101;
													assign node14169 = (inp[11]) ? node14171 : 4'b1100;
														assign node14171 = (inp[7]) ? node14173 : 4'b1101;
															assign node14173 = (inp[10]) ? 4'b0101 : 4'b1101;
												assign node14176 = (inp[7]) ? node14184 : node14177;
													assign node14177 = (inp[12]) ? 4'b1001 : node14178;
														assign node14178 = (inp[10]) ? 4'b0001 : node14179;
															assign node14179 = (inp[11]) ? 4'b1001 : 4'b1000;
													assign node14184 = (inp[12]) ? node14190 : node14185;
														assign node14185 = (inp[10]) ? 4'b0001 : node14186;
															assign node14186 = (inp[11]) ? 4'b1101 : 4'b1100;
														assign node14190 = (inp[10]) ? node14192 : 4'b1100;
															assign node14192 = (inp[14]) ? node14194 : 4'b1101;
																assign node14194 = (inp[11]) ? 4'b1101 : 4'b1100;
										assign node14197 = (inp[13]) ? node14225 : node14198;
											assign node14198 = (inp[10]) ? node14214 : node14199;
												assign node14199 = (inp[12]) ? node14209 : node14200;
													assign node14200 = (inp[7]) ? 4'b1100 : node14201;
														assign node14201 = (inp[14]) ? node14203 : 4'b1100;
															assign node14203 = (inp[11]) ? 4'b1000 : node14204;
																assign node14204 = (inp[4]) ? 4'b0001 : 4'b0101;
													assign node14209 = (inp[11]) ? 4'b0100 : node14210;
														assign node14210 = (inp[14]) ? 4'b0101 : 4'b0100;
												assign node14214 = (inp[11]) ? node14220 : node14215;
													assign node14215 = (inp[14]) ? node14217 : 4'b1100;
														assign node14217 = (inp[12]) ? 4'b0101 : 4'b1101;
													assign node14220 = (inp[7]) ? 4'b1100 : node14221;
														assign node14221 = (inp[14]) ? 4'b1100 : 4'b1000;
											assign node14225 = (inp[7]) ? node14231 : node14226;
												assign node14226 = (inp[11]) ? 4'b0000 : node14227;
													assign node14227 = (inp[14]) ? 4'b1001 : 4'b0000;
												assign node14231 = (inp[4]) ? node14245 : node14232;
													assign node14232 = (inp[12]) ? node14238 : node14233;
														assign node14233 = (inp[10]) ? node14235 : 4'b0100;
															assign node14235 = (inp[11]) ? 4'b0100 : 4'b0101;
														assign node14238 = (inp[10]) ? 4'b0100 : node14239;
															assign node14239 = (inp[14]) ? node14241 : 4'b1100;
																assign node14241 = (inp[11]) ? 4'b1100 : 4'b1101;
													assign node14245 = (inp[12]) ? node14251 : node14246;
														assign node14246 = (inp[14]) ? node14248 : 4'b0000;
															assign node14248 = (inp[11]) ? 4'b0000 : 4'b0001;
														assign node14251 = (inp[10]) ? 4'b0000 : 4'b1100;
								assign node14254 = (inp[4]) ? node14338 : node14255;
									assign node14255 = (inp[1]) ? node14295 : node14256;
										assign node14256 = (inp[11]) ? node14284 : node14257;
											assign node14257 = (inp[14]) ? node14271 : node14258;
												assign node14258 = (inp[13]) ? node14264 : node14259;
													assign node14259 = (inp[10]) ? node14261 : 4'b0001;
														assign node14261 = (inp[12]) ? 4'b0001 : 4'b1001;
													assign node14264 = (inp[10]) ? node14266 : 4'b1001;
														assign node14266 = (inp[7]) ? node14268 : 4'b0101;
															assign node14268 = (inp[12]) ? 4'b1001 : 4'b0001;
												assign node14271 = (inp[13]) ? node14277 : node14272;
													assign node14272 = (inp[12]) ? 4'b0000 : node14273;
														assign node14273 = (inp[10]) ? 4'b1000 : 4'b0000;
													assign node14277 = (inp[10]) ? node14279 : 4'b1000;
														assign node14279 = (inp[12]) ? 4'b1000 : node14280;
															assign node14280 = (inp[7]) ? 4'b0000 : 4'b0100;
											assign node14284 = (inp[13]) ? node14290 : node14285;
												assign node14285 = (inp[10]) ? node14287 : 4'b0001;
													assign node14287 = (inp[12]) ? 4'b0001 : 4'b1001;
												assign node14290 = (inp[10]) ? node14292 : 4'b1001;
													assign node14292 = (inp[12]) ? 4'b1001 : 4'b0001;
										assign node14295 = (inp[11]) ? node14321 : node14296;
											assign node14296 = (inp[14]) ? node14310 : node14297;
												assign node14297 = (inp[13]) ? node14303 : node14298;
													assign node14298 = (inp[12]) ? node14300 : 4'b1000;
														assign node14300 = (inp[10]) ? 4'b1000 : 4'b0000;
													assign node14303 = (inp[10]) ? node14307 : node14304;
														assign node14304 = (inp[12]) ? 4'b1000 : 4'b0100;
														assign node14307 = (inp[7]) ? 4'b0000 : 4'b0100;
												assign node14310 = (inp[13]) ? node14314 : node14311;
													assign node14311 = (inp[10]) ? 4'b1001 : 4'b0001;
													assign node14314 = (inp[10]) ? node14316 : 4'b1001;
														assign node14316 = (inp[12]) ? 4'b1001 : node14317;
															assign node14317 = (inp[7]) ? 4'b0001 : 4'b0101;
											assign node14321 = (inp[13]) ? node14327 : node14322;
												assign node14322 = (inp[12]) ? node14324 : 4'b1000;
													assign node14324 = (inp[10]) ? 4'b1000 : 4'b0000;
												assign node14327 = (inp[7]) ? node14333 : node14328;
													assign node14328 = (inp[12]) ? node14330 : 4'b0100;
														assign node14330 = (inp[10]) ? 4'b0100 : 4'b1000;
													assign node14333 = (inp[10]) ? 4'b0000 : node14334;
														assign node14334 = (inp[12]) ? 4'b1000 : 4'b0000;
									assign node14338 = (inp[7]) ? node14388 : node14339;
										assign node14339 = (inp[1]) ? node14365 : node14340;
											assign node14340 = (inp[14]) ? node14350 : node14341;
												assign node14341 = (inp[13]) ? node14347 : node14342;
													assign node14342 = (inp[10]) ? node14344 : 4'b0101;
														assign node14344 = (inp[12]) ? 4'b0101 : 4'b1101;
													assign node14347 = (inp[10]) ? 4'b0101 : 4'b1101;
												assign node14350 = (inp[11]) ? node14358 : node14351;
													assign node14351 = (inp[13]) ? node14355 : node14352;
														assign node14352 = (inp[10]) ? 4'b1100 : 4'b0100;
														assign node14355 = (inp[10]) ? 4'b0100 : 4'b1100;
													assign node14358 = (inp[13]) ? 4'b1101 : node14359;
														assign node14359 = (inp[5]) ? 4'b0101 : node14360;
															assign node14360 = (inp[12]) ? 4'b0101 : 4'b1101;
											assign node14365 = (inp[14]) ? node14377 : node14366;
												assign node14366 = (inp[13]) ? node14372 : node14367;
													assign node14367 = (inp[10]) ? 4'b1100 : node14368;
														assign node14368 = (inp[12]) ? 4'b0100 : 4'b1100;
													assign node14372 = (inp[12]) ? node14374 : 4'b0100;
														assign node14374 = (inp[10]) ? 4'b0100 : 4'b1100;
												assign node14377 = (inp[11]) ? node14385 : node14378;
													assign node14378 = (inp[13]) ? 4'b1101 : node14379;
														assign node14379 = (inp[10]) ? node14381 : 4'b0101;
															assign node14381 = (inp[12]) ? 4'b0101 : 4'b1101;
													assign node14385 = (inp[12]) ? 4'b1100 : 4'b0100;
										assign node14388 = (inp[1]) ? node14412 : node14389;
											assign node14389 = (inp[13]) ? node14401 : node14390;
												assign node14390 = (inp[12]) ? node14396 : node14391;
													assign node14391 = (inp[10]) ? 4'b1001 : node14392;
														assign node14392 = (inp[14]) ? 4'b0000 : 4'b0001;
													assign node14396 = (inp[11]) ? 4'b0001 : node14397;
														assign node14397 = (inp[14]) ? 4'b0000 : 4'b0001;
												assign node14401 = (inp[12]) ? node14407 : node14402;
													assign node14402 = (inp[10]) ? 4'b0101 : node14403;
														assign node14403 = (inp[11]) ? 4'b1001 : 4'b1000;
													assign node14407 = (inp[5]) ? 4'b1001 : node14408;
														assign node14408 = (inp[14]) ? 4'b1000 : 4'b1001;
											assign node14412 = (inp[14]) ? node14424 : node14413;
												assign node14413 = (inp[13]) ? node14419 : node14414;
													assign node14414 = (inp[10]) ? 4'b1000 : node14415;
														assign node14415 = (inp[12]) ? 4'b0000 : 4'b1000;
													assign node14419 = (inp[12]) ? node14421 : 4'b0100;
														assign node14421 = (inp[10]) ? 4'b0100 : 4'b1000;
												assign node14424 = (inp[11]) ? node14436 : node14425;
													assign node14425 = (inp[13]) ? node14431 : node14426;
														assign node14426 = (inp[10]) ? node14428 : 4'b0001;
															assign node14428 = (inp[12]) ? 4'b0001 : 4'b1001;
														assign node14431 = (inp[10]) ? node14433 : 4'b1001;
															assign node14433 = (inp[12]) ? 4'b1001 : 4'b0101;
													assign node14436 = (inp[12]) ? node14440 : node14437;
														assign node14437 = (inp[13]) ? 4'b0100 : 4'b1000;
														assign node14440 = (inp[13]) ? 4'b1000 : node14441;
															assign node14441 = (inp[10]) ? 4'b1000 : 4'b0000;
							assign node14445 = (inp[5]) ? node14447 : 4'b0110;
								assign node14447 = (inp[3]) ? node14523 : node14448;
									assign node14448 = (inp[4]) ? node14462 : node14449;
										assign node14449 = (inp[13]) ? node14451 : 4'b0110;
											assign node14451 = (inp[7]) ? 4'b0110 : node14452;
												assign node14452 = (inp[10]) ? node14454 : 4'b0110;
													assign node14454 = (inp[12]) ? node14456 : 4'b0001;
														assign node14456 = (inp[14]) ? 4'b0110 : node14457;
															assign node14457 = (inp[1]) ? 4'b0000 : 4'b0110;
										assign node14462 = (inp[7]) ? node14502 : node14463;
											assign node14463 = (inp[1]) ? node14485 : node14464;
												assign node14464 = (inp[14]) ? node14474 : node14465;
													assign node14465 = (inp[10]) ? node14467 : 4'b1001;
														assign node14467 = (inp[12]) ? node14471 : node14468;
															assign node14468 = (inp[13]) ? 4'b0001 : 4'b1001;
															assign node14471 = (inp[13]) ? 4'b1001 : 4'b0001;
													assign node14474 = (inp[11]) ? node14480 : node14475;
														assign node14475 = (inp[13]) ? node14477 : 4'b0000;
															assign node14477 = (inp[10]) ? 4'b0000 : 4'b1000;
														assign node14480 = (inp[10]) ? 4'b1001 : node14481;
															assign node14481 = (inp[13]) ? 4'b1001 : 4'b0001;
												assign node14485 = (inp[14]) ? node14489 : node14486;
													assign node14486 = (inp[13]) ? 4'b0000 : 4'b1000;
													assign node14489 = (inp[11]) ? 4'b1000 : node14490;
														assign node14490 = (inp[13]) ? node14496 : node14491;
															assign node14491 = (inp[12]) ? 4'b0001 : node14492;
																assign node14492 = (inp[10]) ? 4'b1001 : 4'b0001;
															assign node14496 = (inp[10]) ? node14498 : 4'b1001;
																assign node14498 = (inp[12]) ? 4'b1001 : 4'b0001;
											assign node14502 = (inp[13]) ? node14504 : 4'b0110;
												assign node14504 = (inp[10]) ? node14510 : node14505;
													assign node14505 = (inp[12]) ? 4'b0110 : node14506;
														assign node14506 = (inp[14]) ? 4'b0110 : 4'b0000;
													assign node14510 = (inp[12]) ? node14518 : node14511;
														assign node14511 = (inp[1]) ? 4'b0000 : node14512;
															assign node14512 = (inp[14]) ? node14514 : 4'b0001;
																assign node14514 = (inp[11]) ? 4'b0001 : 4'b0000;
														assign node14518 = (inp[1]) ? node14520 : 4'b0110;
															assign node14520 = (inp[11]) ? 4'b0000 : 4'b0110;
									assign node14523 = (inp[4]) ? node14589 : node14524;
										assign node14524 = (inp[1]) ? node14554 : node14525;
											assign node14525 = (inp[11]) ? node14543 : node14526;
												assign node14526 = (inp[14]) ? node14536 : node14527;
													assign node14527 = (inp[10]) ? node14529 : 4'b1001;
														assign node14529 = (inp[7]) ? node14531 : 4'b1001;
															assign node14531 = (inp[12]) ? 4'b0001 : node14532;
																assign node14532 = (inp[13]) ? 4'b0001 : 4'b1001;
													assign node14536 = (inp[13]) ? 4'b1000 : node14537;
														assign node14537 = (inp[10]) ? node14539 : 4'b0000;
															assign node14539 = (inp[12]) ? 4'b0000 : 4'b1000;
												assign node14543 = (inp[13]) ? node14549 : node14544;
													assign node14544 = (inp[12]) ? 4'b0001 : node14545;
														assign node14545 = (inp[7]) ? 4'b0001 : 4'b1001;
													assign node14549 = (inp[12]) ? 4'b1001 : node14550;
														assign node14550 = (inp[7]) ? 4'b0001 : 4'b0101;
											assign node14554 = (inp[11]) ? node14578 : node14555;
												assign node14555 = (inp[14]) ? node14569 : node14556;
													assign node14556 = (inp[7]) ? node14564 : node14557;
														assign node14557 = (inp[12]) ? node14559 : 4'b0100;
															assign node14559 = (inp[10]) ? 4'b0100 : node14560;
																assign node14560 = (inp[13]) ? 4'b1000 : 4'b0000;
														assign node14564 = (inp[12]) ? 4'b0000 : node14565;
															assign node14565 = (inp[13]) ? 4'b0000 : 4'b1000;
													assign node14569 = (inp[13]) ? node14575 : node14570;
														assign node14570 = (inp[12]) ? 4'b0001 : node14571;
															assign node14571 = (inp[10]) ? 4'b1001 : 4'b0001;
														assign node14575 = (inp[10]) ? 4'b0101 : 4'b1001;
												assign node14578 = (inp[13]) ? node14584 : node14579;
													assign node14579 = (inp[10]) ? 4'b1000 : node14580;
														assign node14580 = (inp[12]) ? 4'b0000 : 4'b1000;
													assign node14584 = (inp[10]) ? node14586 : 4'b1000;
														assign node14586 = (inp[7]) ? 4'b0000 : 4'b0100;
										assign node14589 = (inp[7]) ? node14629 : node14590;
											assign node14590 = (inp[13]) ? node14614 : node14591;
												assign node14591 = (inp[10]) ? node14603 : node14592;
													assign node14592 = (inp[1]) ? node14596 : node14593;
														assign node14593 = (inp[14]) ? 4'b0100 : 4'b0101;
														assign node14596 = (inp[14]) ? node14600 : node14597;
															assign node14597 = (inp[12]) ? 4'b0100 : 4'b1100;
															assign node14600 = (inp[11]) ? 4'b0100 : 4'b0101;
													assign node14603 = (inp[1]) ? node14611 : node14604;
														assign node14604 = (inp[12]) ? node14608 : node14605;
															assign node14605 = (inp[14]) ? 4'b1100 : 4'b1101;
															assign node14608 = (inp[11]) ? 4'b0101 : 4'b0100;
														assign node14611 = (inp[12]) ? 4'b1100 : 4'b1101;
												assign node14614 = (inp[10]) ? node14622 : node14615;
													assign node14615 = (inp[12]) ? 4'b1100 : node14616;
														assign node14616 = (inp[1]) ? 4'b1101 : node14617;
															assign node14617 = (inp[14]) ? 4'b1100 : 4'b1101;
													assign node14622 = (inp[12]) ? 4'b1101 : node14623;
														assign node14623 = (inp[11]) ? 4'b0101 : node14624;
															assign node14624 = (inp[14]) ? 4'b0101 : 4'b0100;
											assign node14629 = (inp[1]) ? node14645 : node14630;
												assign node14630 = (inp[13]) ? node14640 : node14631;
													assign node14631 = (inp[10]) ? node14633 : 4'b0001;
														assign node14633 = (inp[12]) ? node14637 : node14634;
															assign node14634 = (inp[14]) ? 4'b1000 : 4'b1001;
															assign node14637 = (inp[11]) ? 4'b0001 : 4'b0000;
													assign node14640 = (inp[10]) ? node14642 : 4'b1001;
														assign node14642 = (inp[12]) ? 4'b1001 : 4'b0101;
												assign node14645 = (inp[11]) ? node14655 : node14646;
													assign node14646 = (inp[14]) ? node14648 : 4'b0100;
														assign node14648 = (inp[10]) ? node14652 : node14649;
															assign node14649 = (inp[13]) ? 4'b1001 : 4'b0001;
															assign node14652 = (inp[13]) ? 4'b0101 : 4'b1001;
													assign node14655 = (inp[13]) ? node14659 : node14656;
														assign node14656 = (inp[10]) ? 4'b1000 : 4'b0000;
														assign node14659 = (inp[14]) ? node14661 : 4'b0100;
															assign node14661 = (inp[12]) ? 4'b1000 : 4'b0100;
					assign node14665 = (inp[5]) ? node15435 : node14666;
						assign node14666 = (inp[0]) ? node15206 : node14667;
							assign node14667 = (inp[11]) ? node14953 : node14668;
								assign node14668 = (inp[3]) ? node14808 : node14669;
									assign node14669 = (inp[4]) ? node14733 : node14670;
										assign node14670 = (inp[13]) ? node14696 : node14671;
											assign node14671 = (inp[10]) ? node14681 : node14672;
												assign node14672 = (inp[1]) ? node14676 : node14673;
													assign node14673 = (inp[14]) ? 4'b0100 : 4'b0101;
													assign node14676 = (inp[14]) ? 4'b0101 : node14677;
														assign node14677 = (inp[12]) ? 4'b0100 : 4'b1100;
												assign node14681 = (inp[2]) ? node14693 : node14682;
													assign node14682 = (inp[12]) ? node14688 : node14683;
														assign node14683 = (inp[1]) ? 4'b0001 : node14684;
															assign node14684 = (inp[14]) ? 4'b1100 : 4'b1101;
														assign node14688 = (inp[1]) ? node14690 : 4'b0101;
															assign node14690 = (inp[14]) ? 4'b0101 : 4'b1100;
													assign node14693 = (inp[12]) ? 4'b0101 : 4'b1101;
											assign node14696 = (inp[7]) ? node14712 : node14697;
												assign node14697 = (inp[2]) ? node14705 : node14698;
													assign node14698 = (inp[14]) ? 4'b1001 : node14699;
														assign node14699 = (inp[12]) ? node14701 : 4'b0001;
															assign node14701 = (inp[10]) ? 4'b1001 : 4'b0001;
													assign node14705 = (inp[14]) ? node14709 : node14706;
														assign node14706 = (inp[1]) ? 4'b0000 : 4'b1101;
														assign node14709 = (inp[1]) ? 4'b1101 : 4'b1100;
												assign node14712 = (inp[12]) ? node14724 : node14713;
													assign node14713 = (inp[10]) ? node14719 : node14714;
														assign node14714 = (inp[1]) ? 4'b0100 : node14715;
															assign node14715 = (inp[14]) ? 4'b1100 : 4'b1101;
														assign node14719 = (inp[1]) ? node14721 : 4'b0100;
															assign node14721 = (inp[14]) ? 4'b0101 : 4'b0100;
													assign node14724 = (inp[14]) ? node14730 : node14725;
														assign node14725 = (inp[1]) ? node14727 : 4'b1101;
															assign node14727 = (inp[10]) ? 4'b0100 : 4'b1100;
														assign node14730 = (inp[1]) ? 4'b1101 : 4'b1100;
										assign node14733 = (inp[2]) ? node14765 : node14734;
											assign node14734 = (inp[7]) ? node14754 : node14735;
												assign node14735 = (inp[13]) ? node14743 : node14736;
													assign node14736 = (inp[10]) ? node14738 : 4'b0001;
														assign node14738 = (inp[1]) ? node14740 : 4'b1001;
															assign node14740 = (inp[12]) ? 4'b1001 : 4'b0101;
													assign node14743 = (inp[10]) ? node14749 : node14744;
														assign node14744 = (inp[1]) ? node14746 : 4'b0101;
															assign node14746 = (inp[12]) ? 4'b0101 : 4'b1101;
														assign node14749 = (inp[12]) ? 4'b1101 : node14750;
															assign node14750 = (inp[1]) ? 4'b0101 : 4'b1101;
												assign node14754 = (inp[10]) ? node14760 : node14755;
													assign node14755 = (inp[12]) ? 4'b0001 : node14756;
														assign node14756 = (inp[1]) ? 4'b1001 : 4'b0001;
													assign node14760 = (inp[1]) ? node14762 : 4'b1001;
														assign node14762 = (inp[12]) ? 4'b1001 : 4'b0101;
											assign node14765 = (inp[7]) ? node14783 : node14766;
												assign node14766 = (inp[12]) ? node14780 : node14767;
													assign node14767 = (inp[10]) ? node14771 : node14768;
														assign node14768 = (inp[14]) ? 4'b1000 : 4'b1001;
														assign node14771 = (inp[13]) ? node14773 : 4'b1000;
															assign node14773 = (inp[14]) ? node14777 : node14774;
																assign node14774 = (inp[1]) ? 4'b0000 : 4'b0001;
																assign node14777 = (inp[1]) ? 4'b0001 : 4'b0000;
													assign node14780 = (inp[13]) ? 4'b1001 : 4'b0001;
												assign node14783 = (inp[13]) ? node14799 : node14784;
													assign node14784 = (inp[10]) ? node14796 : node14785;
														assign node14785 = (inp[12]) ? node14791 : node14786;
															assign node14786 = (inp[1]) ? 4'b0101 : node14787;
																assign node14787 = (inp[14]) ? 4'b0100 : 4'b0101;
															assign node14791 = (inp[1]) ? node14793 : 4'b0100;
																assign node14793 = (inp[14]) ? 4'b0101 : 4'b0100;
														assign node14796 = (inp[14]) ? 4'b0101 : 4'b1100;
													assign node14799 = (inp[12]) ? node14803 : node14800;
														assign node14800 = (inp[10]) ? 4'b0001 : 4'b0000;
														assign node14803 = (inp[1]) ? node14805 : 4'b1100;
															assign node14805 = (inp[14]) ? 4'b1101 : 4'b1100;
									assign node14808 = (inp[2]) ? node14888 : node14809;
										assign node14809 = (inp[4]) ? node14841 : node14810;
											assign node14810 = (inp[13]) ? node14824 : node14811;
												assign node14811 = (inp[10]) ? node14817 : node14812;
													assign node14812 = (inp[1]) ? node14814 : 4'b0101;
														assign node14814 = (inp[12]) ? 4'b0101 : 4'b1101;
													assign node14817 = (inp[14]) ? 4'b1101 : node14818;
														assign node14818 = (inp[1]) ? node14820 : 4'b1101;
															assign node14820 = (inp[12]) ? 4'b1101 : 4'b0101;
												assign node14824 = (inp[7]) ? node14832 : node14825;
													assign node14825 = (inp[10]) ? node14827 : 4'b0001;
														assign node14827 = (inp[1]) ? node14829 : 4'b1001;
															assign node14829 = (inp[12]) ? 4'b1001 : 4'b0001;
													assign node14832 = (inp[10]) ? node14838 : node14833;
														assign node14833 = (inp[12]) ? 4'b0101 : node14834;
															assign node14834 = (inp[1]) ? 4'b1101 : 4'b0101;
														assign node14838 = (inp[12]) ? 4'b1101 : 4'b0001;
											assign node14841 = (inp[7]) ? node14863 : node14842;
												assign node14842 = (inp[13]) ? node14854 : node14843;
													assign node14843 = (inp[1]) ? node14847 : node14844;
														assign node14844 = (inp[14]) ? 4'b0001 : 4'b1000;
														assign node14847 = (inp[14]) ? 4'b1000 : node14848;
															assign node14848 = (inp[12]) ? node14850 : 4'b1001;
																assign node14850 = (inp[10]) ? 4'b0001 : 4'b1001;
													assign node14854 = (inp[1]) ? node14858 : node14855;
														assign node14855 = (inp[10]) ? 4'b0101 : 4'b1001;
														assign node14858 = (inp[12]) ? node14860 : 4'b0101;
															assign node14860 = (inp[10]) ? 4'b1101 : 4'b0101;
												assign node14863 = (inp[1]) ? node14871 : node14864;
													assign node14864 = (inp[14]) ? 4'b0001 : node14865;
														assign node14865 = (inp[13]) ? node14867 : 4'b0000;
															assign node14867 = (inp[12]) ? 4'b1000 : 4'b0000;
													assign node14871 = (inp[14]) ? node14881 : node14872;
														assign node14872 = (inp[10]) ? node14874 : 4'b0001;
															assign node14874 = (inp[13]) ? node14878 : node14875;
																assign node14875 = (inp[12]) ? 4'b0001 : 4'b1001;
																assign node14878 = (inp[12]) ? 4'b1001 : 4'b0101;
														assign node14881 = (inp[13]) ? node14885 : node14882;
															assign node14882 = (inp[12]) ? 4'b0001 : 4'b1001;
															assign node14885 = (inp[10]) ? 4'b1000 : 4'b0000;
										assign node14888 = (inp[4]) ? node14936 : node14889;
											assign node14889 = (inp[13]) ? node14913 : node14890;
												assign node14890 = (inp[10]) ? node14904 : node14891;
													assign node14891 = (inp[12]) ? node14897 : node14892;
														assign node14892 = (inp[1]) ? 4'b0001 : node14893;
															assign node14893 = (inp[14]) ? 4'b0000 : 4'b0001;
														assign node14897 = (inp[1]) ? node14901 : node14898;
															assign node14898 = (inp[14]) ? 4'b0000 : 4'b0001;
															assign node14901 = (inp[14]) ? 4'b0001 : 4'b0000;
													assign node14904 = (inp[7]) ? node14906 : 4'b0001;
														assign node14906 = (inp[14]) ? 4'b1000 : node14907;
															assign node14907 = (inp[1]) ? 4'b1000 : node14908;
																assign node14908 = (inp[12]) ? 4'b0001 : 4'b1001;
												assign node14913 = (inp[7]) ? node14921 : node14914;
													assign node14914 = (inp[10]) ? 4'b1001 : node14915;
														assign node14915 = (inp[12]) ? 4'b0001 : node14916;
															assign node14916 = (inp[1]) ? 4'b1001 : 4'b0001;
													assign node14921 = (inp[12]) ? node14931 : node14922;
														assign node14922 = (inp[10]) ? node14926 : node14923;
															assign node14923 = (inp[14]) ? 4'b1001 : 4'b0000;
															assign node14926 = (inp[14]) ? node14928 : 4'b0001;
																assign node14928 = (inp[1]) ? 4'b0001 : 4'b0000;
														assign node14931 = (inp[10]) ? 4'b1000 : node14932;
															assign node14932 = (inp[1]) ? 4'b1000 : 4'b1001;
											assign node14936 = (inp[10]) ? node14946 : node14937;
												assign node14937 = (inp[1]) ? node14943 : node14938;
													assign node14938 = (inp[14]) ? node14940 : 4'b0001;
														assign node14940 = (inp[13]) ? 4'b0101 : 4'b0001;
													assign node14943 = (inp[12]) ? 4'b0001 : 4'b1001;
												assign node14946 = (inp[12]) ? 4'b1001 : node14947;
													assign node14947 = (inp[14]) ? node14949 : 4'b0101;
														assign node14949 = (inp[7]) ? 4'b1001 : 4'b1101;
								assign node14953 = (inp[1]) ? node15087 : node14954;
									assign node14954 = (inp[3]) ? node15016 : node14955;
										assign node14955 = (inp[2]) ? node14989 : node14956;
											assign node14956 = (inp[4]) ? node14968 : node14957;
												assign node14957 = (inp[13]) ? node14959 : 4'b0101;
													assign node14959 = (inp[12]) ? node14963 : node14960;
														assign node14960 = (inp[7]) ? 4'b0000 : 4'b1000;
														assign node14963 = (inp[7]) ? 4'b1101 : node14964;
															assign node14964 = (inp[10]) ? 4'b1000 : 4'b0000;
												assign node14968 = (inp[13]) ? node14976 : node14969;
													assign node14969 = (inp[14]) ? node14971 : 4'b0000;
														assign node14971 = (inp[12]) ? node14973 : 4'b1000;
															assign node14973 = (inp[10]) ? 4'b1000 : 4'b0000;
													assign node14976 = (inp[7]) ? node14984 : node14977;
														assign node14977 = (inp[10]) ? node14981 : node14978;
															assign node14978 = (inp[14]) ? 4'b0100 : 4'b1100;
															assign node14981 = (inp[12]) ? 4'b1100 : 4'b0100;
														assign node14984 = (inp[12]) ? 4'b1000 : node14985;
															assign node14985 = (inp[10]) ? 4'b0100 : 4'b1000;
											assign node14989 = (inp[4]) ? node15001 : node14990;
												assign node14990 = (inp[13]) ? node14994 : node14991;
													assign node14991 = (inp[12]) ? 4'b0101 : 4'b1101;
													assign node14994 = (inp[12]) ? 4'b1101 : node14995;
														assign node14995 = (inp[10]) ? node14997 : 4'b1101;
															assign node14997 = (inp[7]) ? 4'b0101 : 4'b0001;
												assign node15001 = (inp[7]) ? node15007 : node15002;
													assign node15002 = (inp[12]) ? node15004 : 4'b0001;
														assign node15004 = (inp[13]) ? 4'b1001 : 4'b0001;
													assign node15007 = (inp[10]) ? node15011 : node15008;
														assign node15008 = (inp[13]) ? 4'b1101 : 4'b0101;
														assign node15011 = (inp[12]) ? node15013 : 4'b0001;
															assign node15013 = (inp[13]) ? 4'b1101 : 4'b0101;
										assign node15016 = (inp[2]) ? node15052 : node15017;
											assign node15017 = (inp[4]) ? node15035 : node15018;
												assign node15018 = (inp[10]) ? node15026 : node15019;
													assign node15019 = (inp[12]) ? node15021 : 4'b1100;
														assign node15021 = (inp[7]) ? 4'b0100 : node15022;
															assign node15022 = (inp[14]) ? 4'b0000 : 4'b0100;
													assign node15026 = (inp[12]) ? node15032 : node15027;
														assign node15027 = (inp[7]) ? node15029 : 4'b0000;
															assign node15029 = (inp[13]) ? 4'b0000 : 4'b0100;
														assign node15032 = (inp[7]) ? 4'b1100 : 4'b1000;
												assign node15035 = (inp[13]) ? node15043 : node15036;
													assign node15036 = (inp[10]) ? 4'b0001 : node15037;
														assign node15037 = (inp[7]) ? node15039 : 4'b1001;
															assign node15039 = (inp[12]) ? 4'b0000 : 4'b1000;
													assign node15043 = (inp[12]) ? 4'b1001 : node15044;
														assign node15044 = (inp[10]) ? node15048 : node15045;
															assign node15045 = (inp[7]) ? 4'b0001 : 4'b0101;
															assign node15048 = (inp[14]) ? 4'b1001 : 4'b1101;
											assign node15052 = (inp[4]) ? node15072 : node15053;
												assign node15053 = (inp[7]) ? node15065 : node15054;
													assign node15054 = (inp[13]) ? node15058 : node15055;
														assign node15055 = (inp[10]) ? 4'b0000 : 4'b0001;
														assign node15058 = (inp[10]) ? node15062 : node15059;
															assign node15059 = (inp[12]) ? 4'b0000 : 4'b1000;
															assign node15062 = (inp[12]) ? 4'b1000 : 4'b0000;
													assign node15065 = (inp[13]) ? node15067 : 4'b0001;
														assign node15067 = (inp[12]) ? 4'b1001 : node15068;
															assign node15068 = (inp[10]) ? 4'b0000 : 4'b1001;
												assign node15072 = (inp[7]) ? node15080 : node15073;
													assign node15073 = (inp[10]) ? node15075 : 4'b1000;
														assign node15075 = (inp[12]) ? node15077 : 4'b0100;
															assign node15077 = (inp[13]) ? 4'b1100 : 4'b1000;
													assign node15080 = (inp[10]) ? node15084 : node15081;
														assign node15081 = (inp[12]) ? 4'b0000 : 4'b1000;
														assign node15084 = (inp[12]) ? 4'b1000 : 4'b0000;
									assign node15087 = (inp[10]) ? node15157 : node15088;
										assign node15088 = (inp[3]) ? node15120 : node15089;
											assign node15089 = (inp[4]) ? node15101 : node15090;
												assign node15090 = (inp[13]) ? node15094 : node15091;
													assign node15091 = (inp[12]) ? 4'b0100 : 4'b1100;
													assign node15094 = (inp[12]) ? node15098 : node15095;
														assign node15095 = (inp[2]) ? 4'b0000 : 4'b1000;
														assign node15098 = (inp[2]) ? 4'b1100 : 4'b1000;
												assign node15101 = (inp[2]) ? node15107 : node15102;
													assign node15102 = (inp[7]) ? 4'b1000 : node15103;
														assign node15103 = (inp[13]) ? 4'b1100 : 4'b1000;
													assign node15107 = (inp[7]) ? node15115 : node15108;
														assign node15108 = (inp[13]) ? node15112 : node15109;
															assign node15109 = (inp[14]) ? 4'b1000 : 4'b0000;
															assign node15112 = (inp[12]) ? 4'b1000 : 4'b0000;
														assign node15115 = (inp[12]) ? 4'b1100 : node15116;
															assign node15116 = (inp[13]) ? 4'b0000 : 4'b1100;
											assign node15120 = (inp[7]) ? node15138 : node15121;
												assign node15121 = (inp[13]) ? node15131 : node15122;
													assign node15122 = (inp[4]) ? node15126 : node15123;
														assign node15123 = (inp[2]) ? 4'b0000 : 4'b1100;
														assign node15126 = (inp[12]) ? 4'b1000 : node15127;
															assign node15127 = (inp[2]) ? 4'b1000 : 4'b0000;
													assign node15131 = (inp[4]) ? node15133 : 4'b1000;
														assign node15133 = (inp[12]) ? node15135 : 4'b1100;
															assign node15135 = (inp[2]) ? 4'b1100 : 4'b0100;
												assign node15138 = (inp[2]) ? node15146 : node15139;
													assign node15139 = (inp[4]) ? node15141 : 4'b1100;
														assign node15141 = (inp[12]) ? node15143 : 4'b0000;
															assign node15143 = (inp[13]) ? 4'b0000 : 4'b1000;
													assign node15146 = (inp[4]) ? 4'b1000 : node15147;
														assign node15147 = (inp[14]) ? node15149 : 4'b0000;
															assign node15149 = (inp[13]) ? node15153 : node15150;
																assign node15150 = (inp[12]) ? 4'b0000 : 4'b1000;
																assign node15153 = (inp[12]) ? 4'b1000 : 4'b0000;
										assign node15157 = (inp[13]) ? node15193 : node15158;
											assign node15158 = (inp[4]) ? node15170 : node15159;
												assign node15159 = (inp[3]) ? node15165 : node15160;
													assign node15160 = (inp[2]) ? 4'b1100 : node15161;
														assign node15161 = (inp[7]) ? 4'b1100 : 4'b0000;
													assign node15165 = (inp[2]) ? node15167 : 4'b0100;
														assign node15167 = (inp[7]) ? 4'b1000 : 4'b0000;
												assign node15170 = (inp[7]) ? node15188 : node15171;
													assign node15171 = (inp[12]) ? node15183 : node15172;
														assign node15172 = (inp[14]) ? node15178 : node15173;
															assign node15173 = (inp[3]) ? node15175 : 4'b1000;
																assign node15175 = (inp[2]) ? 4'b0100 : 4'b1000;
															assign node15178 = (inp[3]) ? 4'b1000 : node15179;
																assign node15179 = (inp[2]) ? 4'b1000 : 4'b0100;
														assign node15183 = (inp[3]) ? 4'b0100 : node15184;
															assign node15184 = (inp[2]) ? 4'b1000 : 4'b0100;
													assign node15188 = (inp[3]) ? node15190 : 4'b0000;
														assign node15190 = (inp[2]) ? 4'b0000 : 4'b1000;
											assign node15193 = (inp[4]) ? node15201 : node15194;
												assign node15194 = (inp[7]) ? node15196 : 4'b0000;
													assign node15196 = (inp[2]) ? node15198 : 4'b0000;
														assign node15198 = (inp[3]) ? 4'b0000 : 4'b0100;
												assign node15201 = (inp[3]) ? 4'b0100 : node15202;
													assign node15202 = (inp[2]) ? 4'b0000 : 4'b0100;
							assign node15206 = (inp[2]) ? 4'b0100 : node15207;
								assign node15207 = (inp[3]) ? node15275 : node15208;
									assign node15208 = (inp[4]) ? node15222 : node15209;
										assign node15209 = (inp[7]) ? 4'b0100 : node15210;
											assign node15210 = (inp[1]) ? node15212 : 4'b0100;
												assign node15212 = (inp[13]) ? node15214 : 4'b0100;
													assign node15214 = (inp[12]) ? 4'b0100 : node15215;
														assign node15215 = (inp[14]) ? node15217 : 4'b0000;
															assign node15217 = (inp[10]) ? 4'b0001 : 4'b0100;
										assign node15222 = (inp[7]) ? node15258 : node15223;
											assign node15223 = (inp[1]) ? node15241 : node15224;
												assign node15224 = (inp[13]) ? node15234 : node15225;
													assign node15225 = (inp[12]) ? node15229 : node15226;
														assign node15226 = (inp[14]) ? 4'b0001 : 4'b1001;
														assign node15229 = (inp[14]) ? node15231 : 4'b0001;
															assign node15231 = (inp[11]) ? 4'b0001 : 4'b0000;
													assign node15234 = (inp[10]) ? node15238 : node15235;
														assign node15235 = (inp[14]) ? 4'b1000 : 4'b1001;
														assign node15238 = (inp[12]) ? 4'b1001 : 4'b0001;
												assign node15241 = (inp[13]) ? node15247 : node15242;
													assign node15242 = (inp[12]) ? node15244 : 4'b1000;
														assign node15244 = (inp[11]) ? 4'b1000 : 4'b0001;
													assign node15247 = (inp[11]) ? 4'b0000 : node15248;
														assign node15248 = (inp[14]) ? node15254 : node15249;
															assign node15249 = (inp[12]) ? node15251 : 4'b0000;
																assign node15251 = (inp[10]) ? 4'b0000 : 4'b1000;
															assign node15254 = (inp[12]) ? 4'b1001 : 4'b0001;
											assign node15258 = (inp[13]) ? node15260 : 4'b0100;
												assign node15260 = (inp[1]) ? node15266 : node15261;
													assign node15261 = (inp[10]) ? node15263 : 4'b0100;
														assign node15263 = (inp[12]) ? 4'b0100 : 4'b0001;
													assign node15266 = (inp[12]) ? node15270 : node15267;
														assign node15267 = (inp[10]) ? 4'b0001 : 4'b0000;
														assign node15270 = (inp[11]) ? node15272 : 4'b0100;
															assign node15272 = (inp[10]) ? 4'b0000 : 4'b0100;
									assign node15275 = (inp[7]) ? node15361 : node15276;
										assign node15276 = (inp[4]) ? node15318 : node15277;
											assign node15277 = (inp[1]) ? node15293 : node15278;
												assign node15278 = (inp[13]) ? node15288 : node15279;
													assign node15279 = (inp[10]) ? node15281 : 4'b0001;
														assign node15281 = (inp[12]) ? node15285 : node15282;
															assign node15282 = (inp[14]) ? 4'b1000 : 4'b1001;
															assign node15285 = (inp[11]) ? 4'b0001 : 4'b0000;
													assign node15288 = (inp[12]) ? 4'b1001 : node15289;
														assign node15289 = (inp[10]) ? 4'b0101 : 4'b1001;
												assign node15293 = (inp[11]) ? node15307 : node15294;
													assign node15294 = (inp[14]) ? node15302 : node15295;
														assign node15295 = (inp[13]) ? node15297 : 4'b1000;
															assign node15297 = (inp[10]) ? 4'b0100 : node15298;
																assign node15298 = (inp[12]) ? 4'b1000 : 4'b0100;
														assign node15302 = (inp[12]) ? node15304 : 4'b0101;
															assign node15304 = (inp[13]) ? 4'b1001 : 4'b0001;
													assign node15307 = (inp[10]) ? 4'b1000 : node15308;
														assign node15308 = (inp[14]) ? node15314 : node15309;
															assign node15309 = (inp[12]) ? node15311 : 4'b1000;
																assign node15311 = (inp[13]) ? 4'b1000 : 4'b0000;
															assign node15314 = (inp[12]) ? 4'b1000 : 4'b0100;
											assign node15318 = (inp[1]) ? node15342 : node15319;
												assign node15319 = (inp[11]) ? node15333 : node15320;
													assign node15320 = (inp[14]) ? node15324 : node15321;
														assign node15321 = (inp[10]) ? 4'b1101 : 4'b0101;
														assign node15324 = (inp[13]) ? node15328 : node15325;
															assign node15325 = (inp[12]) ? 4'b0100 : 4'b1100;
															assign node15328 = (inp[12]) ? 4'b1100 : node15329;
																assign node15329 = (inp[10]) ? 4'b0100 : 4'b1100;
													assign node15333 = (inp[13]) ? node15339 : node15334;
														assign node15334 = (inp[10]) ? node15336 : 4'b0101;
															assign node15336 = (inp[12]) ? 4'b0101 : 4'b1101;
														assign node15339 = (inp[10]) ? 4'b0101 : 4'b1101;
												assign node15342 = (inp[14]) ? node15352 : node15343;
													assign node15343 = (inp[10]) ? node15349 : node15344;
														assign node15344 = (inp[13]) ? 4'b1100 : node15345;
															assign node15345 = (inp[12]) ? 4'b0100 : 4'b1100;
														assign node15349 = (inp[13]) ? 4'b0100 : 4'b1100;
													assign node15352 = (inp[11]) ? node15356 : node15353;
														assign node15353 = (inp[13]) ? 4'b1101 : 4'b0101;
														assign node15356 = (inp[13]) ? 4'b0100 : node15357;
															assign node15357 = (inp[10]) ? 4'b1100 : 4'b0100;
										assign node15361 = (inp[1]) ? node15395 : node15362;
											assign node15362 = (inp[11]) ? node15382 : node15363;
												assign node15363 = (inp[14]) ? node15373 : node15364;
													assign node15364 = (inp[10]) ? node15366 : 4'b0001;
														assign node15366 = (inp[4]) ? 4'b0001 : node15367;
															assign node15367 = (inp[13]) ? node15369 : 4'b1001;
																assign node15369 = (inp[12]) ? 4'b1001 : 4'b0001;
													assign node15373 = (inp[13]) ? node15379 : node15374;
														assign node15374 = (inp[10]) ? node15376 : 4'b0000;
															assign node15376 = (inp[12]) ? 4'b0000 : 4'b1000;
														assign node15379 = (inp[12]) ? 4'b1000 : 4'b0000;
												assign node15382 = (inp[13]) ? node15388 : node15383;
													assign node15383 = (inp[10]) ? node15385 : 4'b0001;
														assign node15385 = (inp[12]) ? 4'b0001 : 4'b1001;
													assign node15388 = (inp[10]) ? node15390 : 4'b1001;
														assign node15390 = (inp[12]) ? 4'b1001 : node15391;
															assign node15391 = (inp[4]) ? 4'b0101 : 4'b0001;
											assign node15395 = (inp[11]) ? node15417 : node15396;
												assign node15396 = (inp[14]) ? node15406 : node15397;
													assign node15397 = (inp[10]) ? 4'b1000 : node15398;
														assign node15398 = (inp[13]) ? node15402 : node15399;
															assign node15399 = (inp[12]) ? 4'b0000 : 4'b1000;
															assign node15402 = (inp[12]) ? 4'b1000 : 4'b0000;
													assign node15406 = (inp[13]) ? node15412 : node15407;
														assign node15407 = (inp[4]) ? 4'b0001 : node15408;
															assign node15408 = (inp[10]) ? 4'b1001 : 4'b0001;
														assign node15412 = (inp[4]) ? 4'b1001 : node15413;
															assign node15413 = (inp[12]) ? 4'b1001 : 4'b0001;
												assign node15417 = (inp[13]) ? node15423 : node15418;
													assign node15418 = (inp[12]) ? node15420 : 4'b1000;
														assign node15420 = (inp[10]) ? 4'b1000 : 4'b0000;
													assign node15423 = (inp[4]) ? node15429 : node15424;
														assign node15424 = (inp[12]) ? node15426 : 4'b0000;
															assign node15426 = (inp[10]) ? 4'b0000 : 4'b1000;
														assign node15429 = (inp[12]) ? node15431 : 4'b0100;
															assign node15431 = (inp[10]) ? 4'b0100 : 4'b1000;
						assign node15435 = (inp[3]) ? node15969 : node15436;
							assign node15436 = (inp[4]) ? node15672 : node15437;
								assign node15437 = (inp[13]) ? node15553 : node15438;
									assign node15438 = (inp[0]) ? node15518 : node15439;
										assign node15439 = (inp[7]) ? node15483 : node15440;
											assign node15440 = (inp[10]) ? node15462 : node15441;
												assign node15441 = (inp[11]) ? node15453 : node15442;
													assign node15442 = (inp[2]) ? 4'b0101 : node15443;
														assign node15443 = (inp[1]) ? node15449 : node15444;
															assign node15444 = (inp[14]) ? 4'b0101 : node15445;
																assign node15445 = (inp[12]) ? 4'b0100 : 4'b1100;
															assign node15449 = (inp[12]) ? 4'b1101 : 4'b0000;
													assign node15453 = (inp[12]) ? node15457 : node15454;
														assign node15454 = (inp[2]) ? 4'b1100 : 4'b1101;
														assign node15457 = (inp[2]) ? node15459 : 4'b0000;
															assign node15459 = (inp[1]) ? 4'b1100 : 4'b0100;
												assign node15462 = (inp[1]) ? node15468 : node15463;
													assign node15463 = (inp[2]) ? 4'b0001 : node15464;
														assign node15464 = (inp[11]) ? 4'b1000 : 4'b0000;
													assign node15468 = (inp[2]) ? node15474 : node15469;
														assign node15469 = (inp[11]) ? 4'b0000 : node15470;
															assign node15470 = (inp[12]) ? 4'b1000 : 4'b0000;
														assign node15474 = (inp[14]) ? node15478 : node15475;
															assign node15475 = (inp[11]) ? 4'b1000 : 4'b1001;
															assign node15478 = (inp[11]) ? 4'b1000 : node15479;
																assign node15479 = (inp[12]) ? 4'b0000 : 4'b1000;
											assign node15483 = (inp[12]) ? node15505 : node15484;
												assign node15484 = (inp[10]) ? node15496 : node15485;
													assign node15485 = (inp[11]) ? node15493 : node15486;
														assign node15486 = (inp[2]) ? 4'b0101 : node15487;
															assign node15487 = (inp[14]) ? node15489 : 4'b1100;
																assign node15489 = (inp[1]) ? 4'b1100 : 4'b0101;
														assign node15493 = (inp[2]) ? 4'b1100 : 4'b1101;
													assign node15496 = (inp[2]) ? node15500 : node15497;
														assign node15497 = (inp[1]) ? 4'b0000 : 4'b0100;
														assign node15500 = (inp[11]) ? 4'b0100 : node15501;
															assign node15501 = (inp[1]) ? 4'b0101 : 4'b1101;
												assign node15505 = (inp[11]) ? node15515 : node15506;
													assign node15506 = (inp[2]) ? node15512 : node15507;
														assign node15507 = (inp[10]) ? 4'b1101 : node15508;
															assign node15508 = (inp[14]) ? 4'b1100 : 4'b1101;
														assign node15512 = (inp[10]) ? 4'b1101 : 4'b0101;
													assign node15515 = (inp[2]) ? 4'b1100 : 4'b0101;
										assign node15518 = (inp[2]) ? 4'b0100 : node15519;
											assign node15519 = (inp[1]) ? node15535 : node15520;
												assign node15520 = (inp[14]) ? node15526 : node15521;
													assign node15521 = (inp[12]) ? 4'b0101 : node15522;
														assign node15522 = (inp[10]) ? 4'b1101 : 4'b0101;
													assign node15526 = (inp[11]) ? node15528 : 4'b0100;
														assign node15528 = (inp[7]) ? node15532 : node15529;
															assign node15529 = (inp[10]) ? 4'b0000 : 4'b0101;
															assign node15532 = (inp[12]) ? 4'b0101 : 4'b1101;
												assign node15535 = (inp[14]) ? node15541 : node15536;
													assign node15536 = (inp[7]) ? 4'b1100 : node15537;
														assign node15537 = (inp[11]) ? 4'b0100 : 4'b1100;
													assign node15541 = (inp[11]) ? node15547 : node15542;
														assign node15542 = (inp[10]) ? node15544 : 4'b0101;
															assign node15544 = (inp[7]) ? 4'b1101 : 4'b0101;
														assign node15547 = (inp[10]) ? 4'b1100 : node15548;
															assign node15548 = (inp[12]) ? 4'b0100 : 4'b1100;
									assign node15553 = (inp[2]) ? node15613 : node15554;
										assign node15554 = (inp[0]) ? node15580 : node15555;
											assign node15555 = (inp[1]) ? node15567 : node15556;
												assign node15556 = (inp[12]) ? node15558 : 4'b1000;
													assign node15558 = (inp[11]) ? node15564 : node15559;
														assign node15559 = (inp[10]) ? node15561 : 4'b0000;
															assign node15561 = (inp[7]) ? 4'b0000 : 4'b0100;
														assign node15564 = (inp[7]) ? 4'b1000 : 4'b1100;
												assign node15567 = (inp[11]) ? node15575 : node15568;
													assign node15568 = (inp[12]) ? node15572 : node15569;
														assign node15569 = (inp[14]) ? 4'b0000 : 4'b0100;
														assign node15572 = (inp[10]) ? 4'b1100 : 4'b1000;
													assign node15575 = (inp[7]) ? 4'b0100 : node15576;
														assign node15576 = (inp[10]) ? 4'b0000 : 4'b0100;
											assign node15580 = (inp[7]) ? node15592 : node15581;
												assign node15581 = (inp[11]) ? node15589 : node15582;
													assign node15582 = (inp[10]) ? node15584 : 4'b0001;
														assign node15584 = (inp[12]) ? 4'b1001 : node15585;
															assign node15585 = (inp[1]) ? 4'b0001 : 4'b1001;
													assign node15589 = (inp[10]) ? 4'b0000 : 4'b1000;
												assign node15592 = (inp[10]) ? node15602 : node15593;
													assign node15593 = (inp[14]) ? node15595 : 4'b1101;
														assign node15595 = (inp[11]) ? node15599 : node15596;
															assign node15596 = (inp[1]) ? 4'b1101 : 4'b1100;
															assign node15599 = (inp[1]) ? 4'b1100 : 4'b1101;
													assign node15602 = (inp[12]) ? node15606 : node15603;
														assign node15603 = (inp[11]) ? 4'b0000 : 4'b0001;
														assign node15606 = (inp[1]) ? node15608 : 4'b1101;
															assign node15608 = (inp[11]) ? 4'b0000 : node15609;
																assign node15609 = (inp[14]) ? 4'b1101 : 4'b0100;
										assign node15613 = (inp[0]) ? node15653 : node15614;
											assign node15614 = (inp[1]) ? node15636 : node15615;
												assign node15615 = (inp[10]) ? node15629 : node15616;
													assign node15616 = (inp[14]) ? node15624 : node15617;
														assign node15617 = (inp[11]) ? node15621 : node15618;
															assign node15618 = (inp[12]) ? 4'b1000 : 4'b0000;
															assign node15621 = (inp[12]) ? 4'b0100 : 4'b0001;
														assign node15624 = (inp[12]) ? 4'b1001 : node15625;
															assign node15625 = (inp[11]) ? 4'b0001 : 4'b0101;
													assign node15629 = (inp[11]) ? 4'b1001 : node15630;
														assign node15630 = (inp[14]) ? node15632 : 4'b1000;
															assign node15632 = (inp[12]) ? 4'b0001 : 4'b1001;
												assign node15636 = (inp[11]) ? node15648 : node15637;
													assign node15637 = (inp[12]) ? node15645 : node15638;
														assign node15638 = (inp[14]) ? node15642 : node15639;
															assign node15639 = (inp[7]) ? 4'b0001 : 4'b0101;
															assign node15642 = (inp[7]) ? 4'b0000 : 4'b0100;
														assign node15645 = (inp[14]) ? 4'b1000 : 4'b1001;
													assign node15648 = (inp[7]) ? 4'b0000 : node15649;
														assign node15649 = (inp[10]) ? 4'b0100 : 4'b0000;
											assign node15653 = (inp[7]) ? 4'b0100 : node15654;
												assign node15654 = (inp[12]) ? node15662 : node15655;
													assign node15655 = (inp[1]) ? 4'b0000 : node15656;
														assign node15656 = (inp[11]) ? 4'b0001 : node15657;
															assign node15657 = (inp[10]) ? 4'b0000 : 4'b0100;
													assign node15662 = (inp[14]) ? 4'b0100 : node15663;
														assign node15663 = (inp[11]) ? node15665 : 4'b0000;
															assign node15665 = (inp[10]) ? node15667 : 4'b0100;
																assign node15667 = (inp[1]) ? 4'b0000 : 4'b0100;
								assign node15672 = (inp[2]) ? node15810 : node15673;
									assign node15673 = (inp[11]) ? node15753 : node15674;
										assign node15674 = (inp[10]) ? node15714 : node15675;
											assign node15675 = (inp[13]) ? node15693 : node15676;
												assign node15676 = (inp[0]) ? node15688 : node15677;
													assign node15677 = (inp[7]) ? node15681 : node15678;
														assign node15678 = (inp[12]) ? 4'b0000 : 4'b1000;
														assign node15681 = (inp[12]) ? node15683 : 4'b1100;
															assign node15683 = (inp[14]) ? 4'b1100 : node15684;
																assign node15684 = (inp[1]) ? 4'b0000 : 4'b0100;
													assign node15688 = (inp[12]) ? 4'b0001 : node15689;
														assign node15689 = (inp[1]) ? 4'b1001 : 4'b0001;
												assign node15693 = (inp[7]) ? node15703 : node15694;
													assign node15694 = (inp[0]) ? node15696 : 4'b0001;
														assign node15696 = (inp[12]) ? 4'b0101 : node15697;
															assign node15697 = (inp[1]) ? 4'b0000 : node15698;
																assign node15698 = (inp[14]) ? 4'b0101 : 4'b0000;
													assign node15703 = (inp[0]) ? node15709 : node15704;
														assign node15704 = (inp[12]) ? 4'b1001 : node15705;
															assign node15705 = (inp[1]) ? 4'b0001 : 4'b0101;
														assign node15709 = (inp[1]) ? node15711 : 4'b0001;
															assign node15711 = (inp[12]) ? 4'b0001 : 4'b1001;
											assign node15714 = (inp[7]) ? node15734 : node15715;
												assign node15715 = (inp[12]) ? node15727 : node15716;
													assign node15716 = (inp[0]) ? node15724 : node15717;
														assign node15717 = (inp[13]) ? 4'b0101 : node15718;
															assign node15718 = (inp[1]) ? 4'b1100 : node15719;
																assign node15719 = (inp[14]) ? 4'b1000 : 4'b1001;
														assign node15724 = (inp[13]) ? 4'b0000 : 4'b0101;
													assign node15727 = (inp[14]) ? 4'b0001 : node15728;
														assign node15728 = (inp[1]) ? 4'b1001 : node15729;
															assign node15729 = (inp[0]) ? 4'b1000 : 4'b1001;
												assign node15734 = (inp[13]) ? node15748 : node15735;
													assign node15735 = (inp[1]) ? node15741 : node15736;
														assign node15736 = (inp[14]) ? node15738 : 4'b1001;
															assign node15738 = (inp[0]) ? 4'b1001 : 4'b1000;
														assign node15741 = (inp[0]) ? 4'b0001 : node15742;
															assign node15742 = (inp[12]) ? node15744 : 4'b1000;
																assign node15744 = (inp[14]) ? 4'b0001 : 4'b0000;
													assign node15748 = (inp[12]) ? 4'b1001 : node15749;
														assign node15749 = (inp[1]) ? 4'b1001 : 4'b0001;
										assign node15753 = (inp[10]) ? node15773 : node15754;
											assign node15754 = (inp[1]) ? 4'b1000 : node15755;
												assign node15755 = (inp[7]) ? node15763 : node15756;
													assign node15756 = (inp[12]) ? node15760 : node15757;
														assign node15757 = (inp[0]) ? 4'b0001 : 4'b1001;
														assign node15760 = (inp[13]) ? 4'b1000 : 4'b0000;
													assign node15763 = (inp[12]) ? 4'b0000 : node15764;
														assign node15764 = (inp[13]) ? node15768 : node15765;
															assign node15765 = (inp[0]) ? 4'b1000 : 4'b1100;
															assign node15768 = (inp[0]) ? 4'b1000 : 4'b0000;
											assign node15773 = (inp[1]) ? node15801 : node15774;
												assign node15774 = (inp[12]) ? node15790 : node15775;
													assign node15775 = (inp[0]) ? node15783 : node15776;
														assign node15776 = (inp[13]) ? node15780 : node15777;
															assign node15777 = (inp[7]) ? 4'b0001 : 4'b0101;
															assign node15780 = (inp[7]) ? 4'b1000 : 4'b0001;
														assign node15783 = (inp[13]) ? node15787 : node15784;
															assign node15784 = (inp[7]) ? 4'b0000 : 4'b0100;
															assign node15787 = (inp[7]) ? 4'b0100 : 4'b1001;
													assign node15790 = (inp[0]) ? node15796 : node15791;
														assign node15791 = (inp[13]) ? node15793 : 4'b1001;
															assign node15793 = (inp[14]) ? 4'b0000 : 4'b0001;
														assign node15796 = (inp[7]) ? 4'b1000 : node15797;
															assign node15797 = (inp[13]) ? 4'b1001 : 4'b1000;
												assign node15801 = (inp[13]) ? 4'b0000 : node15802;
													assign node15802 = (inp[7]) ? node15806 : node15803;
														assign node15803 = (inp[0]) ? 4'b0100 : 4'b0000;
														assign node15806 = (inp[0]) ? 4'b0000 : 4'b1000;
									assign node15810 = (inp[7]) ? node15916 : node15811;
										assign node15811 = (inp[1]) ? node15865 : node15812;
											assign node15812 = (inp[11]) ? node15844 : node15813;
												assign node15813 = (inp[14]) ? node15831 : node15814;
													assign node15814 = (inp[0]) ? node15824 : node15815;
														assign node15815 = (inp[12]) ? 4'b0000 : node15816;
															assign node15816 = (inp[13]) ? node15820 : node15817;
																assign node15817 = (inp[10]) ? 4'b1000 : 4'b1100;
																assign node15820 = (inp[10]) ? 4'b0001 : 4'b1000;
														assign node15824 = (inp[13]) ? node15828 : node15825;
															assign node15825 = (inp[12]) ? 4'b0001 : 4'b1001;
															assign node15828 = (inp[12]) ? 4'b1001 : 4'b0001;
													assign node15831 = (inp[0]) ? node15835 : node15832;
														assign node15832 = (inp[12]) ? 4'b0000 : 4'b0101;
														assign node15835 = (inp[13]) ? node15841 : node15836;
															assign node15836 = (inp[12]) ? 4'b0000 : node15837;
																assign node15837 = (inp[10]) ? 4'b1000 : 4'b0000;
															assign node15841 = (inp[12]) ? 4'b1000 : 4'b0000;
												assign node15844 = (inp[13]) ? node15852 : node15845;
													assign node15845 = (inp[0]) ? 4'b0001 : node15846;
														assign node15846 = (inp[10]) ? 4'b1000 : node15847;
															assign node15847 = (inp[12]) ? 4'b0101 : 4'b1101;
													assign node15852 = (inp[10]) ? node15856 : node15853;
														assign node15853 = (inp[0]) ? 4'b1001 : 4'b1000;
														assign node15856 = (inp[14]) ? node15858 : 4'b0001;
															assign node15858 = (inp[0]) ? node15862 : node15859;
																assign node15859 = (inp[12]) ? 4'b0001 : 4'b1001;
																assign node15862 = (inp[12]) ? 4'b1001 : 4'b0001;
											assign node15865 = (inp[11]) ? node15899 : node15866;
												assign node15866 = (inp[14]) ? node15884 : node15867;
													assign node15867 = (inp[12]) ? node15875 : node15868;
														assign node15868 = (inp[13]) ? node15872 : node15869;
															assign node15869 = (inp[0]) ? 4'b1000 : 4'b0000;
															assign node15872 = (inp[0]) ? 4'b0000 : 4'b0100;
														assign node15875 = (inp[13]) ? node15879 : node15876;
															assign node15876 = (inp[10]) ? 4'b1000 : 4'b1101;
															assign node15879 = (inp[0]) ? node15881 : 4'b1000;
																assign node15881 = (inp[10]) ? 4'b0000 : 4'b1000;
													assign node15884 = (inp[0]) ? node15890 : node15885;
														assign node15885 = (inp[10]) ? node15887 : 4'b0100;
															assign node15887 = (inp[13]) ? 4'b1001 : 4'b1000;
														assign node15890 = (inp[13]) ? node15894 : node15891;
															assign node15891 = (inp[10]) ? 4'b1001 : 4'b0001;
															assign node15894 = (inp[12]) ? 4'b1001 : node15895;
																assign node15895 = (inp[10]) ? 4'b0001 : 4'b1001;
												assign node15899 = (inp[0]) ? node15905 : node15900;
													assign node15900 = (inp[10]) ? 4'b0000 : node15901;
														assign node15901 = (inp[14]) ? 4'b0000 : 4'b0100;
													assign node15905 = (inp[13]) ? node15911 : node15906;
														assign node15906 = (inp[10]) ? 4'b1000 : node15907;
															assign node15907 = (inp[12]) ? 4'b0000 : 4'b1000;
														assign node15911 = (inp[10]) ? 4'b0000 : node15912;
															assign node15912 = (inp[12]) ? 4'b1000 : 4'b0000;
										assign node15916 = (inp[0]) ? node15952 : node15917;
											assign node15917 = (inp[13]) ? node15939 : node15918;
												assign node15918 = (inp[1]) ? node15928 : node15919;
													assign node15919 = (inp[14]) ? node15925 : node15920;
														assign node15920 = (inp[10]) ? 4'b0100 : node15921;
															assign node15921 = (inp[11]) ? 4'b0001 : 4'b0000;
														assign node15925 = (inp[10]) ? 4'b1001 : 4'b0001;
													assign node15928 = (inp[10]) ? node15934 : node15929;
														assign node15929 = (inp[11]) ? node15931 : 4'b1000;
															assign node15931 = (inp[14]) ? 4'b0100 : 4'b1000;
														assign node15934 = (inp[11]) ? 4'b0000 : node15935;
															assign node15935 = (inp[12]) ? 4'b0101 : 4'b0000;
												assign node15939 = (inp[1]) ? node15945 : node15940;
													assign node15940 = (inp[12]) ? node15942 : 4'b1000;
														assign node15942 = (inp[11]) ? 4'b1000 : 4'b0000;
													assign node15945 = (inp[12]) ? 4'b1000 : node15946;
														assign node15946 = (inp[14]) ? node15948 : 4'b0000;
															assign node15948 = (inp[11]) ? 4'b0000 : 4'b0100;
											assign node15952 = (inp[13]) ? node15954 : 4'b0100;
												assign node15954 = (inp[12]) ? node15962 : node15955;
													assign node15955 = (inp[10]) ? node15959 : node15956;
														assign node15956 = (inp[11]) ? 4'b0000 : 4'b0100;
														assign node15959 = (inp[11]) ? 4'b0001 : 4'b0000;
													assign node15962 = (inp[10]) ? node15964 : 4'b0100;
														assign node15964 = (inp[1]) ? node15966 : 4'b0100;
															assign node15966 = (inp[11]) ? 4'b0000 : 4'b0100;
							assign node15969 = (inp[4]) ? node16257 : node15970;
								assign node15970 = (inp[11]) ? node16146 : node15971;
									assign node15971 = (inp[1]) ? node16055 : node15972;
										assign node15972 = (inp[0]) ? node16010 : node15973;
											assign node15973 = (inp[10]) ? node15993 : node15974;
												assign node15974 = (inp[12]) ? node15984 : node15975;
													assign node15975 = (inp[2]) ? node15979 : node15976;
														assign node15976 = (inp[14]) ? 4'b1001 : 4'b1000;
														assign node15979 = (inp[13]) ? 4'b0000 : node15980;
															assign node15980 = (inp[14]) ? 4'b1000 : 4'b1001;
													assign node15984 = (inp[13]) ? node15990 : node15985;
														assign node15985 = (inp[2]) ? node15987 : 4'b0001;
															assign node15987 = (inp[14]) ? 4'b0000 : 4'b0001;
														assign node15990 = (inp[7]) ? 4'b0000 : 4'b1001;
												assign node15993 = (inp[12]) ? node16001 : node15994;
													assign node15994 = (inp[13]) ? node15998 : node15995;
														assign node15995 = (inp[2]) ? 4'b0001 : 4'b0000;
														assign node15998 = (inp[2]) ? 4'b1000 : 4'b0000;
													assign node16001 = (inp[2]) ? node16003 : 4'b1000;
														assign node16003 = (inp[7]) ? 4'b1000 : node16004;
															assign node16004 = (inp[13]) ? node16006 : 4'b1001;
																assign node16006 = (inp[14]) ? 4'b0000 : 4'b0001;
											assign node16010 = (inp[10]) ? node16030 : node16011;
												assign node16011 = (inp[7]) ? node16023 : node16012;
													assign node16012 = (inp[2]) ? node16018 : node16013;
														assign node16013 = (inp[13]) ? 4'b0000 : node16014;
															assign node16014 = (inp[12]) ? 4'b0000 : 4'b0001;
														assign node16018 = (inp[14]) ? node16020 : 4'b0001;
															assign node16020 = (inp[13]) ? 4'b0001 : 4'b0000;
													assign node16023 = (inp[12]) ? node16025 : 4'b1000;
														assign node16025 = (inp[14]) ? node16027 : 4'b0000;
															assign node16027 = (inp[2]) ? 4'b0000 : 4'b0001;
												assign node16030 = (inp[2]) ? node16044 : node16031;
													assign node16031 = (inp[13]) ? node16039 : node16032;
														assign node16032 = (inp[7]) ? node16036 : node16033;
															assign node16033 = (inp[14]) ? 4'b0000 : 4'b1000;
															assign node16036 = (inp[12]) ? 4'b1001 : 4'b0001;
														assign node16039 = (inp[14]) ? node16041 : 4'b0001;
															assign node16041 = (inp[7]) ? 4'b0000 : 4'b0001;
													assign node16044 = (inp[14]) ? node16048 : node16045;
														assign node16045 = (inp[7]) ? 4'b0001 : 4'b1001;
														assign node16048 = (inp[13]) ? node16052 : node16049;
															assign node16049 = (inp[12]) ? 4'b0000 : 4'b1000;
															assign node16052 = (inp[7]) ? 4'b1000 : 4'b1001;
										assign node16055 = (inp[13]) ? node16101 : node16056;
											assign node16056 = (inp[2]) ? node16084 : node16057;
												assign node16057 = (inp[10]) ? node16071 : node16058;
													assign node16058 = (inp[14]) ? node16068 : node16059;
														assign node16059 = (inp[7]) ? node16063 : node16060;
															assign node16060 = (inp[12]) ? 4'b1001 : 4'b0000;
															assign node16063 = (inp[0]) ? 4'b1001 : node16064;
																assign node16064 = (inp[12]) ? 4'b0001 : 4'b1001;
														assign node16068 = (inp[12]) ? 4'b0000 : 4'b1000;
													assign node16071 = (inp[12]) ? node16075 : node16072;
														assign node16072 = (inp[0]) ? 4'b0000 : 4'b0001;
														assign node16075 = (inp[0]) ? node16079 : node16076;
															assign node16076 = (inp[14]) ? 4'b1000 : 4'b0000;
															assign node16079 = (inp[7]) ? node16081 : 4'b1000;
																assign node16081 = (inp[14]) ? 4'b0000 : 4'b0001;
												assign node16084 = (inp[14]) ? node16094 : node16085;
													assign node16085 = (inp[0]) ? node16087 : 4'b0001;
														assign node16087 = (inp[12]) ? 4'b0000 : node16088;
															assign node16088 = (inp[7]) ? 4'b1000 : node16089;
																assign node16089 = (inp[10]) ? 4'b0001 : 4'b1000;
													assign node16094 = (inp[0]) ? 4'b0001 : node16095;
														assign node16095 = (inp[7]) ? node16097 : 4'b0000;
															assign node16097 = (inp[10]) ? 4'b1001 : 4'b0001;
											assign node16101 = (inp[10]) ? node16121 : node16102;
												assign node16102 = (inp[7]) ? node16112 : node16103;
													assign node16103 = (inp[0]) ? node16109 : node16104;
														assign node16104 = (inp[14]) ? 4'b1000 : node16105;
															assign node16105 = (inp[2]) ? 4'b1000 : 4'b1001;
														assign node16109 = (inp[12]) ? 4'b0001 : 4'b1001;
													assign node16112 = (inp[12]) ? node16116 : node16113;
														assign node16113 = (inp[0]) ? 4'b0000 : 4'b0001;
														assign node16116 = (inp[0]) ? node16118 : 4'b1001;
															assign node16118 = (inp[2]) ? 4'b1001 : 4'b1000;
												assign node16121 = (inp[14]) ? node16135 : node16122;
													assign node16122 = (inp[7]) ? node16130 : node16123;
														assign node16123 = (inp[12]) ? 4'b1001 : node16124;
															assign node16124 = (inp[0]) ? 4'b0001 : node16125;
																assign node16125 = (inp[2]) ? 4'b1001 : 4'b0001;
														assign node16130 = (inp[0]) ? 4'b0000 : node16131;
															assign node16131 = (inp[2]) ? 4'b1000 : 4'b0000;
													assign node16135 = (inp[0]) ? node16141 : node16136;
														assign node16136 = (inp[2]) ? node16138 : 4'b0001;
															assign node16138 = (inp[12]) ? 4'b0001 : 4'b1001;
														assign node16141 = (inp[2]) ? node16143 : 4'b1001;
															assign node16143 = (inp[7]) ? 4'b0001 : 4'b0000;
									assign node16146 = (inp[1]) ? node16216 : node16147;
										assign node16147 = (inp[12]) ? node16187 : node16148;
											assign node16148 = (inp[7]) ? node16164 : node16149;
												assign node16149 = (inp[2]) ? node16159 : node16150;
													assign node16150 = (inp[10]) ? node16156 : node16151;
														assign node16151 = (inp[13]) ? 4'b0001 : node16152;
															assign node16152 = (inp[0]) ? 4'b1001 : 4'b0000;
														assign node16156 = (inp[0]) ? 4'b1000 : 4'b1001;
													assign node16159 = (inp[13]) ? node16161 : 4'b0000;
														assign node16161 = (inp[14]) ? 4'b0000 : 4'b1000;
												assign node16164 = (inp[10]) ? node16172 : node16165;
													assign node16165 = (inp[2]) ? 4'b1001 : node16166;
														assign node16166 = (inp[13]) ? 4'b1000 : node16167;
															assign node16167 = (inp[0]) ? 4'b1001 : 4'b0001;
													assign node16172 = (inp[0]) ? node16180 : node16173;
														assign node16173 = (inp[2]) ? node16177 : node16174;
															assign node16174 = (inp[13]) ? 4'b1000 : 4'b0000;
															assign node16177 = (inp[13]) ? 4'b0001 : 4'b1000;
														assign node16180 = (inp[2]) ? node16184 : node16181;
															assign node16181 = (inp[13]) ? 4'b1001 : 4'b0001;
															assign node16184 = (inp[13]) ? 4'b0000 : 4'b1001;
											assign node16187 = (inp[13]) ? node16199 : node16188;
												assign node16188 = (inp[7]) ? node16196 : node16189;
													assign node16189 = (inp[10]) ? node16193 : node16190;
														assign node16190 = (inp[0]) ? 4'b0001 : 4'b1001;
														assign node16193 = (inp[2]) ? 4'b0000 : 4'b1000;
													assign node16196 = (inp[0]) ? 4'b0001 : 4'b0000;
												assign node16199 = (inp[7]) ? node16207 : node16200;
													assign node16200 = (inp[10]) ? node16202 : 4'b0000;
														assign node16202 = (inp[0]) ? node16204 : 4'b1001;
															assign node16204 = (inp[2]) ? 4'b1000 : 4'b0000;
													assign node16207 = (inp[2]) ? 4'b1001 : node16208;
														assign node16208 = (inp[0]) ? node16212 : node16209;
															assign node16209 = (inp[10]) ? 4'b1000 : 4'b0000;
															assign node16212 = (inp[10]) ? 4'b0001 : 4'b1000;
										assign node16216 = (inp[13]) ? node16244 : node16217;
											assign node16217 = (inp[12]) ? node16233 : node16218;
												assign node16218 = (inp[2]) ? node16224 : node16219;
													assign node16219 = (inp[10]) ? node16221 : 4'b0000;
														assign node16221 = (inp[0]) ? 4'b0000 : 4'b1000;
													assign node16224 = (inp[10]) ? node16226 : 4'b1000;
														assign node16226 = (inp[7]) ? node16230 : node16227;
															assign node16227 = (inp[0]) ? 4'b0000 : 4'b1000;
															assign node16230 = (inp[0]) ? 4'b1000 : 4'b0000;
												assign node16233 = (inp[0]) ? 4'b0000 : node16234;
													assign node16234 = (inp[7]) ? node16238 : node16235;
														assign node16235 = (inp[2]) ? 4'b1000 : 4'b0000;
														assign node16238 = (inp[10]) ? node16240 : 4'b0000;
															assign node16240 = (inp[2]) ? 4'b0000 : 4'b1000;
											assign node16244 = (inp[10]) ? 4'b0000 : node16245;
												assign node16245 = (inp[0]) ? node16253 : node16246;
													assign node16246 = (inp[2]) ? 4'b0000 : node16247;
														assign node16247 = (inp[7]) ? node16249 : 4'b0000;
															assign node16249 = (inp[12]) ? 4'b0000 : 4'b1000;
													assign node16253 = (inp[7]) ? 4'b0000 : 4'b1000;
								assign node16257 = (inp[13]) ? node16425 : node16258;
									assign node16258 = (inp[11]) ? node16352 : node16259;
										assign node16259 = (inp[7]) ? node16305 : node16260;
											assign node16260 = (inp[2]) ? node16284 : node16261;
												assign node16261 = (inp[10]) ? node16275 : node16262;
													assign node16262 = (inp[0]) ? node16268 : node16263;
														assign node16263 = (inp[1]) ? node16265 : 4'b0000;
															assign node16265 = (inp[12]) ? 4'b0001 : 4'b1001;
														assign node16268 = (inp[1]) ? node16272 : node16269;
															assign node16269 = (inp[14]) ? 4'b1001 : 4'b1000;
															assign node16272 = (inp[14]) ? 4'b1000 : 4'b0000;
													assign node16275 = (inp[1]) ? node16281 : node16276;
														assign node16276 = (inp[12]) ? node16278 : 4'b0001;
															assign node16278 = (inp[14]) ? 4'b0001 : 4'b1001;
														assign node16281 = (inp[0]) ? 4'b0000 : 4'b0001;
												assign node16284 = (inp[14]) ? node16294 : node16285;
													assign node16285 = (inp[10]) ? node16291 : node16286;
														assign node16286 = (inp[0]) ? 4'b0000 : node16287;
															assign node16287 = (inp[1]) ? 4'b1000 : 4'b0000;
														assign node16291 = (inp[1]) ? 4'b0000 : 4'b1000;
													assign node16294 = (inp[10]) ? node16300 : node16295;
														assign node16295 = (inp[12]) ? node16297 : 4'b0000;
															assign node16297 = (inp[1]) ? 4'b0001 : 4'b1001;
														assign node16300 = (inp[12]) ? 4'b0000 : node16301;
															assign node16301 = (inp[0]) ? 4'b0001 : 4'b0000;
											assign node16305 = (inp[0]) ? node16325 : node16306;
												assign node16306 = (inp[14]) ? node16320 : node16307;
													assign node16307 = (inp[2]) ? node16311 : node16308;
														assign node16308 = (inp[12]) ? 4'b0000 : 4'b1000;
														assign node16311 = (inp[12]) ? node16315 : node16312;
															assign node16312 = (inp[1]) ? 4'b0001 : 4'b0000;
															assign node16315 = (inp[1]) ? 4'b1000 : node16316;
																assign node16316 = (inp[10]) ? 4'b0001 : 4'b1001;
													assign node16320 = (inp[10]) ? 4'b0001 : node16321;
														assign node16321 = (inp[2]) ? 4'b0000 : 4'b0001;
												assign node16325 = (inp[10]) ? node16337 : node16326;
													assign node16326 = (inp[12]) ? 4'b0001 : node16327;
														assign node16327 = (inp[1]) ? node16331 : node16328;
															assign node16328 = (inp[2]) ? 4'b0001 : 4'b1001;
															assign node16331 = (inp[14]) ? node16333 : 4'b1001;
																assign node16333 = (inp[2]) ? 4'b1001 : 4'b1000;
													assign node16337 = (inp[12]) ? node16347 : node16338;
														assign node16338 = (inp[1]) ? 4'b0000 : node16339;
															assign node16339 = (inp[2]) ? node16343 : node16340;
																assign node16340 = (inp[14]) ? 4'b0000 : 4'b0001;
																assign node16343 = (inp[14]) ? 4'b0001 : 4'b0000;
														assign node16347 = (inp[1]) ? 4'b0001 : node16348;
															assign node16348 = (inp[2]) ? 4'b1001 : 4'b1000;
										assign node16352 = (inp[1]) ? node16398 : node16353;
											assign node16353 = (inp[2]) ? node16371 : node16354;
												assign node16354 = (inp[0]) ? node16364 : node16355;
													assign node16355 = (inp[7]) ? node16359 : node16356;
														assign node16356 = (inp[10]) ? 4'b0000 : 4'b0001;
														assign node16359 = (inp[10]) ? node16361 : 4'b0000;
															assign node16361 = (inp[14]) ? 4'b1000 : 4'b0000;
													assign node16364 = (inp[12]) ? node16366 : 4'b0001;
														assign node16366 = (inp[10]) ? 4'b0001 : node16367;
															assign node16367 = (inp[7]) ? 4'b1000 : 4'b0000;
												assign node16371 = (inp[10]) ? node16387 : node16372;
													assign node16372 = (inp[12]) ? node16382 : node16373;
														assign node16373 = (inp[14]) ? node16375 : 4'b1000;
															assign node16375 = (inp[7]) ? node16379 : node16376;
																assign node16376 = (inp[0]) ? 4'b1001 : 4'b1000;
																assign node16379 = (inp[0]) ? 4'b1000 : 4'b1001;
														assign node16382 = (inp[7]) ? node16384 : 4'b1000;
															assign node16384 = (inp[0]) ? 4'b0000 : 4'b0001;
													assign node16387 = (inp[0]) ? node16393 : node16388;
														assign node16388 = (inp[12]) ? node16390 : 4'b0000;
															assign node16390 = (inp[7]) ? 4'b0000 : 4'b0001;
														assign node16393 = (inp[12]) ? node16395 : 4'b0001;
															assign node16395 = (inp[14]) ? 4'b1000 : 4'b0001;
											assign node16398 = (inp[10]) ? 4'b0000 : node16399;
												assign node16399 = (inp[12]) ? node16413 : node16400;
													assign node16400 = (inp[14]) ? node16406 : node16401;
														assign node16401 = (inp[0]) ? node16403 : 4'b1000;
															assign node16403 = (inp[7]) ? 4'b0000 : 4'b1000;
														assign node16406 = (inp[2]) ? 4'b0000 : node16407;
															assign node16407 = (inp[7]) ? 4'b0000 : node16408;
																assign node16408 = (inp[0]) ? 4'b1000 : 4'b0000;
													assign node16413 = (inp[7]) ? node16415 : 4'b0000;
														assign node16415 = (inp[14]) ? 4'b1000 : node16416;
															assign node16416 = (inp[2]) ? node16420 : node16417;
																assign node16417 = (inp[0]) ? 4'b0000 : 4'b1000;
																assign node16420 = (inp[0]) ? 4'b1000 : 4'b0000;
									assign node16425 = (inp[11]) ? node16477 : node16426;
										assign node16426 = (inp[10]) ? node16454 : node16427;
											assign node16427 = (inp[14]) ? node16437 : node16428;
												assign node16428 = (inp[0]) ? node16430 : 4'b0000;
													assign node16430 = (inp[1]) ? node16432 : 4'b0000;
														assign node16432 = (inp[2]) ? node16434 : 4'b0001;
															assign node16434 = (inp[7]) ? 4'b0001 : 4'b0000;
												assign node16437 = (inp[7]) ? node16447 : node16438;
													assign node16438 = (inp[0]) ? node16442 : node16439;
														assign node16439 = (inp[2]) ? 4'b0000 : 4'b0001;
														assign node16442 = (inp[2]) ? 4'b0001 : node16443;
															assign node16443 = (inp[1]) ? 4'b0001 : 4'b0000;
													assign node16447 = (inp[0]) ? 4'b0000 : node16448;
														assign node16448 = (inp[12]) ? node16450 : 4'b0001;
															assign node16450 = (inp[2]) ? 4'b0001 : 4'b0000;
											assign node16454 = (inp[1]) ? 4'b0000 : node16455;
												assign node16455 = (inp[7]) ? node16461 : node16456;
													assign node16456 = (inp[0]) ? node16458 : 4'b0000;
														assign node16458 = (inp[2]) ? 4'b0000 : 4'b0001;
													assign node16461 = (inp[0]) ? node16467 : node16462;
														assign node16462 = (inp[12]) ? node16464 : 4'b0001;
															assign node16464 = (inp[2]) ? 4'b0000 : 4'b0001;
														assign node16467 = (inp[2]) ? node16473 : node16468;
															assign node16468 = (inp[12]) ? 4'b0000 : node16469;
																assign node16469 = (inp[14]) ? 4'b0000 : 4'b0001;
															assign node16473 = (inp[14]) ? 4'b0001 : 4'b0000;
										assign node16477 = (inp[1]) ? 4'b0000 : node16478;
											assign node16478 = (inp[10]) ? 4'b0000 : node16479;
												assign node16479 = (inp[7]) ? node16487 : node16480;
													assign node16480 = (inp[2]) ? node16484 : node16481;
														assign node16481 = (inp[12]) ? 4'b0000 : 4'b0001;
														assign node16484 = (inp[0]) ? 4'b0000 : 4'b0001;
													assign node16487 = (inp[2]) ? node16489 : 4'b0000;
														assign node16489 = (inp[12]) ? node16493 : node16490;
															assign node16490 = (inp[0]) ? 4'b0000 : 4'b0001;
															assign node16493 = (inp[14]) ? 4'b0001 : 4'b0000;
				assign node16498 = (inp[0]) ? node18010 : node16499;
					assign node16499 = (inp[6]) ? node16917 : node16500;
						assign node16500 = (inp[5]) ? node16586 : node16501;
							assign node16501 = (inp[2]) ? 4'b0010 : node16502;
								assign node16502 = (inp[3]) ? node16504 : 4'b0010;
									assign node16504 = (inp[7]) ? node16568 : node16505;
										assign node16505 = (inp[4]) ? node16523 : node16506;
											assign node16506 = (inp[13]) ? node16508 : 4'b0010;
												assign node16508 = (inp[10]) ? node16518 : node16509;
													assign node16509 = (inp[12]) ? 4'b0010 : node16510;
														assign node16510 = (inp[1]) ? node16512 : 4'b0010;
															assign node16512 = (inp[14]) ? node16514 : 4'b0000;
																assign node16514 = (inp[11]) ? 4'b0000 : 4'b0010;
													assign node16518 = (inp[1]) ? 4'b0000 : node16519;
														assign node16519 = (inp[12]) ? 4'b0010 : 4'b0000;
											assign node16523 = (inp[1]) ? node16545 : node16524;
												assign node16524 = (inp[14]) ? node16532 : node16525;
													assign node16525 = (inp[10]) ? node16529 : node16526;
														assign node16526 = (inp[13]) ? 4'b1001 : 4'b0001;
														assign node16529 = (inp[13]) ? 4'b0001 : 4'b1001;
													assign node16532 = (inp[11]) ? node16542 : node16533;
														assign node16533 = (inp[13]) ? node16539 : node16534;
															assign node16534 = (inp[12]) ? 4'b0000 : node16535;
																assign node16535 = (inp[10]) ? 4'b1000 : 4'b0000;
															assign node16539 = (inp[12]) ? 4'b1000 : 4'b0000;
														assign node16542 = (inp[13]) ? 4'b1001 : 4'b0001;
												assign node16545 = (inp[14]) ? node16557 : node16546;
													assign node16546 = (inp[13]) ? node16552 : node16547;
														assign node16547 = (inp[12]) ? node16549 : 4'b1000;
															assign node16549 = (inp[10]) ? 4'b1000 : 4'b0000;
														assign node16552 = (inp[12]) ? node16554 : 4'b0000;
															assign node16554 = (inp[10]) ? 4'b0000 : 4'b1000;
													assign node16557 = (inp[11]) ? 4'b0000 : node16558;
														assign node16558 = (inp[12]) ? 4'b0001 : node16559;
															assign node16559 = (inp[13]) ? node16563 : node16560;
																assign node16560 = (inp[10]) ? 4'b1001 : 4'b0001;
																assign node16563 = (inp[10]) ? 4'b0001 : 4'b1001;
										assign node16568 = (inp[1]) ? node16570 : 4'b0010;
											assign node16570 = (inp[13]) ? node16572 : 4'b0010;
												assign node16572 = (inp[4]) ? node16574 : 4'b0010;
													assign node16574 = (inp[12]) ? node16580 : node16575;
														assign node16575 = (inp[11]) ? 4'b0000 : node16576;
															assign node16576 = (inp[14]) ? 4'b0010 : 4'b0000;
														assign node16580 = (inp[10]) ? node16582 : 4'b0010;
															assign node16582 = (inp[14]) ? 4'b0010 : 4'b0000;
							assign node16586 = (inp[2]) ? node16834 : node16587;
								assign node16587 = (inp[1]) ? node16711 : node16588;
									assign node16588 = (inp[13]) ? node16644 : node16589;
										assign node16589 = (inp[14]) ? node16617 : node16590;
											assign node16590 = (inp[10]) ? node16602 : node16591;
												assign node16591 = (inp[3]) ? node16597 : node16592;
													assign node16592 = (inp[7]) ? 4'b0001 : node16593;
														assign node16593 = (inp[4]) ? 4'b0101 : 4'b0001;
													assign node16597 = (inp[7]) ? 4'b0101 : node16598;
														assign node16598 = (inp[4]) ? 4'b0001 : 4'b0101;
												assign node16602 = (inp[12]) ? node16610 : node16603;
													assign node16603 = (inp[4]) ? node16605 : 4'b1101;
														assign node16605 = (inp[11]) ? node16607 : 4'b1001;
															assign node16607 = (inp[3]) ? 4'b1001 : 4'b1101;
													assign node16610 = (inp[11]) ? 4'b0001 : node16611;
														assign node16611 = (inp[3]) ? node16613 : 4'b0101;
															assign node16613 = (inp[7]) ? 4'b0101 : 4'b0001;
											assign node16617 = (inp[11]) ? node16635 : node16618;
												assign node16618 = (inp[10]) ? node16628 : node16619;
													assign node16619 = (inp[3]) ? node16625 : node16620;
														assign node16620 = (inp[4]) ? node16622 : 4'b0000;
															assign node16622 = (inp[7]) ? 4'b0000 : 4'b0100;
														assign node16625 = (inp[7]) ? 4'b0100 : 4'b0000;
													assign node16628 = (inp[12]) ? 4'b0100 : node16629;
														assign node16629 = (inp[4]) ? 4'b1100 : node16630;
															assign node16630 = (inp[3]) ? 4'b1100 : 4'b1000;
												assign node16635 = (inp[3]) ? node16639 : node16636;
													assign node16636 = (inp[7]) ? 4'b0001 : 4'b0101;
													assign node16639 = (inp[10]) ? node16641 : 4'b0101;
														assign node16641 = (inp[4]) ? 4'b0001 : 4'b1101;
										assign node16644 = (inp[12]) ? node16686 : node16645;
											assign node16645 = (inp[10]) ? node16665 : node16646;
												assign node16646 = (inp[14]) ? node16658 : node16647;
													assign node16647 = (inp[11]) ? node16653 : node16648;
														assign node16648 = (inp[3]) ? 4'b1101 : node16649;
															assign node16649 = (inp[4]) ? 4'b1101 : 4'b1001;
														assign node16653 = (inp[3]) ? node16655 : 4'b1001;
															assign node16655 = (inp[4]) ? 4'b1001 : 4'b1101;
													assign node16658 = (inp[11]) ? 4'b1001 : node16659;
														assign node16659 = (inp[3]) ? 4'b1100 : node16660;
															assign node16660 = (inp[4]) ? 4'b1100 : 4'b1000;
												assign node16665 = (inp[3]) ? node16675 : node16666;
													assign node16666 = (inp[7]) ? node16672 : node16667;
														assign node16667 = (inp[14]) ? node16669 : 4'b0101;
															assign node16669 = (inp[11]) ? 4'b0101 : 4'b0100;
														assign node16672 = (inp[4]) ? 4'b0101 : 4'b0001;
													assign node16675 = (inp[4]) ? 4'b0001 : node16676;
														assign node16676 = (inp[7]) ? node16680 : node16677;
															assign node16677 = (inp[14]) ? 4'b0000 : 4'b0001;
															assign node16680 = (inp[11]) ? 4'b0101 : node16681;
																assign node16681 = (inp[14]) ? 4'b0100 : 4'b0101;
											assign node16686 = (inp[3]) ? node16696 : node16687;
												assign node16687 = (inp[4]) ? node16693 : node16688;
													assign node16688 = (inp[11]) ? 4'b1001 : node16689;
														assign node16689 = (inp[14]) ? 4'b1000 : 4'b1001;
													assign node16693 = (inp[7]) ? 4'b1001 : 4'b1101;
												assign node16696 = (inp[11]) ? node16706 : node16697;
													assign node16697 = (inp[14]) ? node16701 : node16698;
														assign node16698 = (inp[7]) ? 4'b1101 : 4'b1001;
														assign node16701 = (inp[7]) ? 4'b1100 : node16702;
															assign node16702 = (inp[10]) ? 4'b1000 : 4'b1100;
													assign node16706 = (inp[4]) ? node16708 : 4'b1101;
														assign node16708 = (inp[7]) ? 4'b1101 : 4'b1001;
									assign node16711 = (inp[14]) ? node16769 : node16712;
										assign node16712 = (inp[13]) ? node16744 : node16713;
											assign node16713 = (inp[12]) ? node16725 : node16714;
												assign node16714 = (inp[3]) ? node16720 : node16715;
													assign node16715 = (inp[7]) ? 4'b1000 : node16716;
														assign node16716 = (inp[4]) ? 4'b1100 : 4'b1000;
													assign node16720 = (inp[4]) ? node16722 : 4'b1100;
														assign node16722 = (inp[7]) ? 4'b1100 : 4'b1000;
												assign node16725 = (inp[10]) ? node16737 : node16726;
													assign node16726 = (inp[3]) ? node16732 : node16727;
														assign node16727 = (inp[4]) ? node16729 : 4'b0000;
															assign node16729 = (inp[7]) ? 4'b0000 : 4'b0100;
														assign node16732 = (inp[4]) ? node16734 : 4'b0100;
															assign node16734 = (inp[7]) ? 4'b0100 : 4'b0000;
													assign node16737 = (inp[7]) ? 4'b1000 : node16738;
														assign node16738 = (inp[11]) ? 4'b1100 : node16739;
															assign node16739 = (inp[4]) ? 4'b1000 : 4'b1100;
											assign node16744 = (inp[12]) ? node16756 : node16745;
												assign node16745 = (inp[3]) ? node16751 : node16746;
													assign node16746 = (inp[4]) ? 4'b0100 : node16747;
														assign node16747 = (inp[7]) ? 4'b0000 : 4'b0100;
													assign node16751 = (inp[10]) ? 4'b0000 : node16752;
														assign node16752 = (inp[7]) ? 4'b0100 : 4'b0000;
												assign node16756 = (inp[10]) ? node16762 : node16757;
													assign node16757 = (inp[3]) ? node16759 : 4'b1000;
														assign node16759 = (inp[7]) ? 4'b1100 : 4'b1000;
													assign node16762 = (inp[3]) ? 4'b0000 : node16763;
														assign node16763 = (inp[4]) ? 4'b0100 : node16764;
															assign node16764 = (inp[7]) ? 4'b0000 : 4'b0100;
										assign node16769 = (inp[11]) ? node16805 : node16770;
											assign node16770 = (inp[13]) ? node16792 : node16771;
												assign node16771 = (inp[10]) ? node16783 : node16772;
													assign node16772 = (inp[3]) ? node16778 : node16773;
														assign node16773 = (inp[4]) ? node16775 : 4'b0001;
															assign node16775 = (inp[7]) ? 4'b0001 : 4'b0101;
														assign node16778 = (inp[12]) ? 4'b0101 : node16779;
															assign node16779 = (inp[4]) ? 4'b0001 : 4'b0101;
													assign node16783 = (inp[12]) ? node16787 : node16784;
														assign node16784 = (inp[7]) ? 4'b1001 : 4'b1101;
														assign node16787 = (inp[7]) ? 4'b0101 : node16788;
															assign node16788 = (inp[3]) ? 4'b0001 : 4'b0101;
												assign node16792 = (inp[3]) ? node16794 : 4'b1001;
													assign node16794 = (inp[7]) ? node16800 : node16795;
														assign node16795 = (inp[4]) ? node16797 : 4'b1101;
															assign node16797 = (inp[12]) ? 4'b1001 : 4'b0001;
														assign node16800 = (inp[12]) ? 4'b1101 : node16801;
															assign node16801 = (inp[4]) ? 4'b1101 : 4'b0101;
											assign node16805 = (inp[13]) ? node16819 : node16806;
												assign node16806 = (inp[3]) ? node16810 : node16807;
													assign node16807 = (inp[10]) ? 4'b1000 : 4'b0000;
													assign node16810 = (inp[7]) ? node16814 : node16811;
														assign node16811 = (inp[4]) ? 4'b1000 : 4'b1100;
														assign node16814 = (inp[12]) ? node16816 : 4'b1100;
															assign node16816 = (inp[4]) ? 4'b0100 : 4'b1100;
												assign node16819 = (inp[12]) ? node16827 : node16820;
													assign node16820 = (inp[10]) ? 4'b0100 : node16821;
														assign node16821 = (inp[7]) ? node16823 : 4'b0000;
															assign node16823 = (inp[3]) ? 4'b0100 : 4'b0000;
													assign node16827 = (inp[10]) ? 4'b0000 : node16828;
														assign node16828 = (inp[4]) ? node16830 : 4'b1000;
															assign node16830 = (inp[7]) ? 4'b1000 : 4'b1100;
								assign node16834 = (inp[3]) ? node16836 : 4'b0010;
									assign node16836 = (inp[4]) ? node16856 : node16837;
										assign node16837 = (inp[7]) ? 4'b0010 : node16838;
											assign node16838 = (inp[13]) ? node16840 : 4'b0010;
												assign node16840 = (inp[12]) ? node16850 : node16841;
													assign node16841 = (inp[10]) ? node16845 : node16842;
														assign node16842 = (inp[11]) ? 4'b0000 : 4'b0010;
														assign node16845 = (inp[14]) ? 4'b0000 : node16846;
															assign node16846 = (inp[11]) ? 4'b0001 : 4'b0000;
													assign node16850 = (inp[1]) ? node16852 : 4'b0010;
														assign node16852 = (inp[10]) ? 4'b0000 : 4'b0010;
										assign node16856 = (inp[7]) ? node16898 : node16857;
											assign node16857 = (inp[1]) ? node16881 : node16858;
												assign node16858 = (inp[11]) ? node16872 : node16859;
													assign node16859 = (inp[14]) ? node16863 : node16860;
														assign node16860 = (inp[13]) ? 4'b1001 : 4'b0001;
														assign node16863 = (inp[13]) ? node16869 : node16864;
															assign node16864 = (inp[10]) ? node16866 : 4'b0000;
																assign node16866 = (inp[12]) ? 4'b0000 : 4'b1000;
															assign node16869 = (inp[10]) ? 4'b0000 : 4'b1000;
													assign node16872 = (inp[13]) ? node16878 : node16873;
														assign node16873 = (inp[12]) ? 4'b0001 : node16874;
															assign node16874 = (inp[10]) ? 4'b1001 : 4'b0001;
														assign node16878 = (inp[12]) ? 4'b1001 : 4'b0001;
												assign node16881 = (inp[13]) ? node16889 : node16882;
													assign node16882 = (inp[14]) ? node16884 : 4'b1000;
														assign node16884 = (inp[11]) ? 4'b1000 : node16885;
															assign node16885 = (inp[12]) ? 4'b0001 : 4'b1001;
													assign node16889 = (inp[12]) ? node16891 : 4'b0000;
														assign node16891 = (inp[10]) ? 4'b0000 : node16892;
															assign node16892 = (inp[14]) ? node16894 : 4'b1000;
																assign node16894 = (inp[11]) ? 4'b1000 : 4'b1001;
											assign node16898 = (inp[13]) ? node16900 : 4'b0010;
												assign node16900 = (inp[12]) ? node16910 : node16901;
													assign node16901 = (inp[11]) ? 4'b0001 : node16902;
														assign node16902 = (inp[1]) ? node16906 : node16903;
															assign node16903 = (inp[14]) ? 4'b0000 : 4'b0001;
															assign node16906 = (inp[14]) ? 4'b0001 : 4'b0000;
													assign node16910 = (inp[14]) ? 4'b0010 : node16911;
														assign node16911 = (inp[10]) ? node16913 : 4'b0010;
															assign node16913 = (inp[1]) ? 4'b0000 : 4'b0010;
						assign node16917 = (inp[5]) ? node17429 : node16918;
							assign node16918 = (inp[1]) ? node17172 : node16919;
								assign node16919 = (inp[3]) ? node17017 : node16920;
									assign node16920 = (inp[11]) ? node16978 : node16921;
										assign node16921 = (inp[14]) ? node16947 : node16922;
											assign node16922 = (inp[4]) ? node16934 : node16923;
												assign node16923 = (inp[13]) ? node16929 : node16924;
													assign node16924 = (inp[12]) ? 4'b0001 : node16925;
														assign node16925 = (inp[10]) ? 4'b1001 : 4'b0001;
													assign node16929 = (inp[12]) ? 4'b1001 : node16930;
														assign node16930 = (inp[10]) ? 4'b0001 : 4'b1001;
												assign node16934 = (inp[7]) ? 4'b1001 : node16935;
													assign node16935 = (inp[10]) ? node16937 : 4'b0101;
														assign node16937 = (inp[12]) ? node16941 : node16938;
															assign node16938 = (inp[2]) ? 4'b0101 : 4'b1101;
															assign node16941 = (inp[13]) ? node16943 : 4'b0101;
																assign node16943 = (inp[2]) ? 4'b1101 : 4'b1001;
											assign node16947 = (inp[4]) ? node16959 : node16948;
												assign node16948 = (inp[13]) ? node16954 : node16949;
													assign node16949 = (inp[10]) ? node16951 : 4'b0000;
														assign node16951 = (inp[12]) ? 4'b0000 : 4'b1000;
													assign node16954 = (inp[10]) ? node16956 : 4'b1000;
														assign node16956 = (inp[2]) ? 4'b0000 : 4'b1000;
												assign node16959 = (inp[7]) ? node16971 : node16960;
													assign node16960 = (inp[13]) ? node16966 : node16961;
														assign node16961 = (inp[10]) ? node16963 : 4'b0100;
															assign node16963 = (inp[12]) ? 4'b0100 : 4'b1100;
														assign node16966 = (inp[2]) ? node16968 : 4'b1001;
															assign node16968 = (inp[12]) ? 4'b1100 : 4'b0100;
													assign node16971 = (inp[10]) ? node16975 : node16972;
														assign node16972 = (inp[13]) ? 4'b1000 : 4'b0000;
														assign node16975 = (inp[13]) ? 4'b0100 : 4'b1000;
										assign node16978 = (inp[7]) ? node17006 : node16979;
											assign node16979 = (inp[4]) ? node16989 : node16980;
												assign node16980 = (inp[13]) ? node16986 : node16981;
													assign node16981 = (inp[10]) ? node16983 : 4'b0001;
														assign node16983 = (inp[12]) ? 4'b0001 : 4'b1001;
													assign node16986 = (inp[10]) ? 4'b0101 : 4'b1001;
												assign node16989 = (inp[13]) ? node16995 : node16990;
													assign node16990 = (inp[12]) ? 4'b0101 : node16991;
														assign node16991 = (inp[10]) ? 4'b1101 : 4'b0101;
													assign node16995 = (inp[2]) ? node17003 : node16996;
														assign node16996 = (inp[10]) ? node17000 : node16997;
															assign node16997 = (inp[12]) ? 4'b0000 : 4'b1000;
															assign node17000 = (inp[12]) ? 4'b1000 : 4'b0000;
														assign node17003 = (inp[12]) ? 4'b1101 : 4'b0101;
											assign node17006 = (inp[13]) ? node17012 : node17007;
												assign node17007 = (inp[10]) ? node17009 : 4'b0001;
													assign node17009 = (inp[12]) ? 4'b0001 : 4'b1001;
												assign node17012 = (inp[10]) ? node17014 : 4'b1001;
													assign node17014 = (inp[12]) ? 4'b1001 : 4'b0001;
									assign node17017 = (inp[10]) ? node17085 : node17018;
										assign node17018 = (inp[13]) ? node17056 : node17019;
											assign node17019 = (inp[14]) ? node17033 : node17020;
												assign node17020 = (inp[2]) ? node17028 : node17021;
													assign node17021 = (inp[4]) ? node17025 : node17022;
														assign node17022 = (inp[11]) ? 4'b0000 : 4'b0001;
														assign node17025 = (inp[11]) ? 4'b0100 : 4'b0101;
													assign node17028 = (inp[7]) ? 4'b0101 : node17029;
														assign node17029 = (inp[4]) ? 4'b0001 : 4'b0101;
												assign node17033 = (inp[12]) ? node17049 : node17034;
													assign node17034 = (inp[2]) ? node17040 : node17035;
														assign node17035 = (inp[11]) ? 4'b1100 : node17036;
															assign node17036 = (inp[7]) ? 4'b0001 : 4'b0101;
														assign node17040 = (inp[11]) ? node17044 : node17041;
															assign node17041 = (inp[4]) ? 4'b0000 : 4'b0100;
															assign node17044 = (inp[4]) ? node17046 : 4'b0101;
																assign node17046 = (inp[7]) ? 4'b0101 : 4'b0001;
													assign node17049 = (inp[11]) ? 4'b0000 : node17050;
														assign node17050 = (inp[2]) ? 4'b0100 : node17051;
															assign node17051 = (inp[7]) ? 4'b0101 : 4'b0001;
											assign node17056 = (inp[4]) ? node17066 : node17057;
												assign node17057 = (inp[2]) ? node17061 : node17058;
													assign node17058 = (inp[12]) ? 4'b0100 : 4'b1100;
													assign node17061 = (inp[11]) ? 4'b1101 : node17062;
														assign node17062 = (inp[7]) ? 4'b1100 : 4'b1101;
												assign node17066 = (inp[7]) ? node17076 : node17067;
													assign node17067 = (inp[11]) ? node17073 : node17068;
														assign node17068 = (inp[12]) ? 4'b0001 : node17069;
															assign node17069 = (inp[2]) ? 4'b0001 : 4'b0000;
														assign node17073 = (inp[12]) ? 4'b0000 : 4'b0001;
													assign node17076 = (inp[2]) ? node17082 : node17077;
														assign node17077 = (inp[11]) ? node17079 : 4'b0101;
															assign node17079 = (inp[12]) ? 4'b0100 : 4'b1100;
														assign node17082 = (inp[14]) ? 4'b1100 : 4'b1101;
										assign node17085 = (inp[11]) ? node17135 : node17086;
											assign node17086 = (inp[2]) ? node17096 : node17087;
												assign node17087 = (inp[4]) ? node17091 : node17088;
													assign node17088 = (inp[7]) ? 4'b1001 : 4'b1101;
													assign node17091 = (inp[13]) ? node17093 : 4'b1101;
														assign node17093 = (inp[7]) ? 4'b1101 : 4'b0001;
												assign node17096 = (inp[14]) ? node17114 : node17097;
													assign node17097 = (inp[7]) ? node17107 : node17098;
														assign node17098 = (inp[4]) ? node17104 : node17099;
															assign node17099 = (inp[13]) ? 4'b0001 : node17100;
																assign node17100 = (inp[12]) ? 4'b0101 : 4'b1101;
															assign node17104 = (inp[12]) ? 4'b0001 : 4'b1001;
														assign node17107 = (inp[12]) ? node17111 : node17108;
															assign node17108 = (inp[13]) ? 4'b0101 : 4'b1101;
															assign node17111 = (inp[13]) ? 4'b1101 : 4'b0101;
													assign node17114 = (inp[7]) ? node17122 : node17115;
														assign node17115 = (inp[4]) ? node17119 : node17116;
															assign node17116 = (inp[12]) ? 4'b1100 : 4'b0000;
															assign node17119 = (inp[13]) ? 4'b1001 : 4'b1000;
														assign node17122 = (inp[4]) ? node17130 : node17123;
															assign node17123 = (inp[12]) ? node17127 : node17124;
																assign node17124 = (inp[13]) ? 4'b0100 : 4'b1100;
																assign node17127 = (inp[13]) ? 4'b1100 : 4'b0100;
															assign node17130 = (inp[13]) ? 4'b0000 : node17131;
																assign node17131 = (inp[12]) ? 4'b0100 : 4'b1100;
											assign node17135 = (inp[12]) ? node17153 : node17136;
												assign node17136 = (inp[4]) ? node17144 : node17137;
													assign node17137 = (inp[2]) ? node17141 : node17138;
														assign node17138 = (inp[7]) ? 4'b0000 : 4'b0100;
														assign node17141 = (inp[13]) ? 4'b0001 : 4'b1101;
													assign node17144 = (inp[2]) ? 4'b0000 : node17145;
														assign node17145 = (inp[13]) ? node17149 : node17146;
															assign node17146 = (inp[7]) ? 4'b0100 : 4'b0000;
															assign node17149 = (inp[7]) ? 4'b0000 : 4'b1001;
												assign node17153 = (inp[2]) ? node17161 : node17154;
													assign node17154 = (inp[4]) ? 4'b1100 : node17155;
														assign node17155 = (inp[13]) ? node17157 : 4'b1000;
															assign node17157 = (inp[7]) ? 4'b1000 : 4'b1100;
													assign node17161 = (inp[13]) ? node17167 : node17162;
														assign node17162 = (inp[4]) ? node17164 : 4'b0101;
															assign node17164 = (inp[14]) ? 4'b0101 : 4'b0001;
														assign node17167 = (inp[4]) ? node17169 : 4'b1101;
															assign node17169 = (inp[7]) ? 4'b1101 : 4'b1000;
								assign node17172 = (inp[11]) ? node17316 : node17173;
									assign node17173 = (inp[14]) ? node17247 : node17174;
										assign node17174 = (inp[3]) ? node17210 : node17175;
											assign node17175 = (inp[7]) ? node17197 : node17176;
												assign node17176 = (inp[12]) ? node17186 : node17177;
													assign node17177 = (inp[4]) ? node17179 : 4'b0100;
														assign node17179 = (inp[2]) ? node17183 : node17180;
															assign node17180 = (inp[10]) ? 4'b0001 : 4'b1001;
															assign node17183 = (inp[10]) ? 4'b0100 : 4'b1100;
													assign node17186 = (inp[4]) ? node17192 : node17187;
														assign node17187 = (inp[10]) ? node17189 : 4'b1000;
															assign node17189 = (inp[13]) ? 4'b0100 : 4'b1000;
														assign node17192 = (inp[10]) ? 4'b1100 : node17193;
															assign node17193 = (inp[13]) ? 4'b1100 : 4'b0100;
												assign node17197 = (inp[13]) ? node17203 : node17198;
													assign node17198 = (inp[12]) ? node17200 : 4'b1000;
														assign node17200 = (inp[10]) ? 4'b1000 : 4'b0000;
													assign node17203 = (inp[12]) ? node17207 : node17204;
														assign node17204 = (inp[10]) ? 4'b0000 : 4'b0100;
														assign node17207 = (inp[10]) ? 4'b0100 : 4'b1000;
											assign node17210 = (inp[2]) ? node17230 : node17211;
												assign node17211 = (inp[7]) ? node17219 : node17212;
													assign node17212 = (inp[13]) ? node17214 : 4'b1101;
														assign node17214 = (inp[12]) ? node17216 : 4'b0001;
															assign node17216 = (inp[10]) ? 4'b1101 : 4'b0101;
													assign node17219 = (inp[4]) ? 4'b1101 : node17220;
														assign node17220 = (inp[13]) ? node17222 : 4'b0001;
															assign node17222 = (inp[10]) ? node17226 : node17223;
																assign node17223 = (inp[12]) ? 4'b0001 : 4'b1001;
																assign node17226 = (inp[12]) ? 4'b1001 : 4'b0101;
												assign node17230 = (inp[13]) ? node17238 : node17231;
													assign node17231 = (inp[10]) ? 4'b1100 : node17232;
														assign node17232 = (inp[7]) ? 4'b1100 : node17233;
															assign node17233 = (inp[4]) ? 4'b0000 : 4'b0100;
													assign node17238 = (inp[7]) ? node17242 : node17239;
														assign node17239 = (inp[4]) ? 4'b1001 : 4'b0000;
														assign node17242 = (inp[12]) ? node17244 : 4'b0000;
															assign node17244 = (inp[4]) ? 4'b1100 : 4'b0100;
										assign node17247 = (inp[13]) ? node17279 : node17248;
											assign node17248 = (inp[3]) ? node17264 : node17249;
												assign node17249 = (inp[10]) ? node17255 : node17250;
													assign node17250 = (inp[7]) ? 4'b0001 : node17251;
														assign node17251 = (inp[4]) ? 4'b0101 : 4'b0001;
													assign node17255 = (inp[12]) ? 4'b0001 : node17256;
														assign node17256 = (inp[2]) ? node17260 : node17257;
															assign node17257 = (inp[7]) ? 4'b1001 : 4'b0001;
															assign node17260 = (inp[4]) ? 4'b1101 : 4'b1001;
												assign node17264 = (inp[2]) ? node17270 : node17265;
													assign node17265 = (inp[4]) ? 4'b1101 : node17266;
														assign node17266 = (inp[12]) ? 4'b0001 : 4'b1001;
													assign node17270 = (inp[7]) ? node17274 : node17271;
														assign node17271 = (inp[4]) ? 4'b0001 : 4'b0101;
														assign node17274 = (inp[10]) ? node17276 : 4'b0101;
															assign node17276 = (inp[12]) ? 4'b0101 : 4'b1101;
											assign node17279 = (inp[2]) ? node17297 : node17280;
												assign node17280 = (inp[3]) ? node17286 : node17281;
													assign node17281 = (inp[7]) ? 4'b1001 : node17282;
														assign node17282 = (inp[4]) ? 4'b1001 : 4'b0101;
													assign node17286 = (inp[4]) ? node17290 : node17287;
														assign node17287 = (inp[7]) ? 4'b1001 : 4'b1101;
														assign node17290 = (inp[12]) ? 4'b1000 : node17291;
															assign node17291 = (inp[7]) ? node17293 : 4'b0000;
																assign node17293 = (inp[10]) ? 4'b0000 : 4'b1101;
												assign node17297 = (inp[10]) ? node17307 : node17298;
													assign node17298 = (inp[3]) ? node17304 : node17299;
														assign node17299 = (inp[4]) ? node17301 : 4'b1001;
															assign node17301 = (inp[7]) ? 4'b1001 : 4'b1101;
														assign node17304 = (inp[7]) ? 4'b1101 : 4'b0001;
													assign node17307 = (inp[12]) ? node17313 : node17308;
														assign node17308 = (inp[3]) ? 4'b0001 : node17309;
															assign node17309 = (inp[4]) ? 4'b0101 : 4'b0001;
														assign node17313 = (inp[3]) ? 4'b1101 : 4'b1001;
									assign node17316 = (inp[10]) ? node17386 : node17317;
										assign node17317 = (inp[3]) ? node17353 : node17318;
											assign node17318 = (inp[7]) ? node17334 : node17319;
												assign node17319 = (inp[4]) ? node17327 : node17320;
													assign node17320 = (inp[13]) ? node17324 : node17321;
														assign node17321 = (inp[12]) ? 4'b0000 : 4'b1000;
														assign node17324 = (inp[12]) ? 4'b1000 : 4'b0100;
													assign node17327 = (inp[13]) ? node17329 : 4'b0100;
														assign node17329 = (inp[2]) ? node17331 : 4'b1000;
															assign node17331 = (inp[14]) ? 4'b0100 : 4'b1100;
												assign node17334 = (inp[2]) ? node17344 : node17335;
													assign node17335 = (inp[13]) ? node17339 : node17336;
														assign node17336 = (inp[12]) ? 4'b0000 : 4'b1000;
														assign node17339 = (inp[12]) ? 4'b1000 : node17340;
															assign node17340 = (inp[4]) ? 4'b0100 : 4'b0000;
													assign node17344 = (inp[13]) ? node17348 : node17345;
														assign node17345 = (inp[12]) ? 4'b0000 : 4'b1000;
														assign node17348 = (inp[12]) ? 4'b1000 : node17349;
															assign node17349 = (inp[4]) ? 4'b0100 : 4'b0000;
											assign node17353 = (inp[7]) ? node17373 : node17354;
												assign node17354 = (inp[4]) ? node17364 : node17355;
													assign node17355 = (inp[14]) ? 4'b1100 : node17356;
														assign node17356 = (inp[2]) ? node17358 : 4'b1000;
															assign node17358 = (inp[12]) ? 4'b1100 : node17359;
																assign node17359 = (inp[13]) ? 4'b0000 : 4'b1100;
													assign node17364 = (inp[13]) ? node17370 : node17365;
														assign node17365 = (inp[2]) ? node17367 : 4'b1100;
															assign node17367 = (inp[12]) ? 4'b0000 : 4'b1000;
														assign node17370 = (inp[2]) ? 4'b1000 : 4'b0000;
												assign node17373 = (inp[4]) ? node17379 : node17374;
													assign node17374 = (inp[2]) ? node17376 : 4'b1000;
														assign node17376 = (inp[13]) ? 4'b1100 : 4'b0100;
													assign node17379 = (inp[2]) ? node17381 : 4'b1100;
														assign node17381 = (inp[13]) ? node17383 : 4'b1100;
															assign node17383 = (inp[12]) ? 4'b1100 : 4'b0000;
										assign node17386 = (inp[13]) ? node17414 : node17387;
											assign node17387 = (inp[3]) ? node17399 : node17388;
												assign node17388 = (inp[2]) ? node17394 : node17389;
													assign node17389 = (inp[7]) ? 4'b1000 : node17390;
														assign node17390 = (inp[4]) ? 4'b0000 : 4'b1000;
													assign node17394 = (inp[4]) ? node17396 : 4'b1000;
														assign node17396 = (inp[7]) ? 4'b1000 : 4'b1100;
												assign node17399 = (inp[2]) ? node17409 : node17400;
													assign node17400 = (inp[14]) ? node17402 : 4'b0000;
														assign node17402 = (inp[7]) ? node17406 : node17403;
															assign node17403 = (inp[4]) ? 4'b0000 : 4'b0100;
															assign node17406 = (inp[4]) ? 4'b0100 : 4'b0000;
													assign node17409 = (inp[4]) ? node17411 : 4'b1100;
														assign node17411 = (inp[14]) ? 4'b1100 : 4'b0000;
											assign node17414 = (inp[4]) ? node17424 : node17415;
												assign node17415 = (inp[7]) ? node17421 : node17416;
													assign node17416 = (inp[2]) ? node17418 : 4'b0100;
														assign node17418 = (inp[14]) ? 4'b0000 : 4'b0100;
													assign node17421 = (inp[3]) ? 4'b0100 : 4'b0000;
												assign node17424 = (inp[3]) ? 4'b0000 : node17425;
													assign node17425 = (inp[2]) ? 4'b0100 : 4'b0000;
							assign node17429 = (inp[3]) ? node17757 : node17430;
								assign node17430 = (inp[1]) ? node17604 : node17431;
									assign node17431 = (inp[14]) ? node17515 : node17432;
										assign node17432 = (inp[13]) ? node17472 : node17433;
											assign node17433 = (inp[2]) ? node17455 : node17434;
												assign node17434 = (inp[11]) ? node17442 : node17435;
													assign node17435 = (inp[10]) ? node17439 : node17436;
														assign node17436 = (inp[12]) ? 4'b0000 : 4'b1000;
														assign node17439 = (inp[7]) ? 4'b0000 : 4'b0100;
													assign node17442 = (inp[4]) ? node17450 : node17443;
														assign node17443 = (inp[10]) ? node17447 : node17444;
															assign node17444 = (inp[12]) ? 4'b0001 : 4'b1001;
															assign node17447 = (inp[7]) ? 4'b0001 : 4'b0101;
														assign node17450 = (inp[7]) ? 4'b1000 : node17451;
															assign node17451 = (inp[12]) ? 4'b1000 : 4'b0001;
												assign node17455 = (inp[4]) ? node17461 : node17456;
													assign node17456 = (inp[10]) ? 4'b1001 : node17457;
														assign node17457 = (inp[11]) ? 4'b0000 : 4'b0001;
													assign node17461 = (inp[10]) ? node17469 : node17462;
														assign node17462 = (inp[7]) ? node17466 : node17463;
															assign node17463 = (inp[11]) ? 4'b0001 : 4'b0000;
															assign node17466 = (inp[12]) ? 4'b0100 : 4'b0101;
														assign node17469 = (inp[11]) ? 4'b0001 : 4'b0000;
											assign node17472 = (inp[4]) ? node17500 : node17473;
												assign node17473 = (inp[12]) ? node17485 : node17474;
													assign node17474 = (inp[7]) ? node17480 : node17475;
														assign node17475 = (inp[2]) ? node17477 : 4'b1000;
															assign node17477 = (inp[11]) ? 4'b0100 : 4'b0101;
														assign node17480 = (inp[2]) ? 4'b1000 : node17481;
															assign node17481 = (inp[10]) ? 4'b1100 : 4'b0100;
													assign node17485 = (inp[10]) ? node17491 : node17486;
														assign node17486 = (inp[2]) ? 4'b0001 : node17487;
															assign node17487 = (inp[11]) ? 4'b1001 : 4'b1000;
														assign node17491 = (inp[7]) ? node17495 : node17492;
															assign node17492 = (inp[2]) ? 4'b1101 : 4'b0000;
															assign node17495 = (inp[2]) ? 4'b1000 : node17496;
																assign node17496 = (inp[11]) ? 4'b1101 : 4'b1100;
												assign node17500 = (inp[2]) ? node17506 : node17501;
													assign node17501 = (inp[7]) ? 4'b0001 : node17502;
														assign node17502 = (inp[11]) ? 4'b1000 : 4'b0001;
													assign node17506 = (inp[11]) ? node17508 : 4'b1000;
														assign node17508 = (inp[10]) ? node17512 : node17509;
															assign node17509 = (inp[12]) ? 4'b1001 : 4'b0101;
															assign node17512 = (inp[7]) ? 4'b1001 : 4'b1000;
										assign node17515 = (inp[4]) ? node17569 : node17516;
											assign node17516 = (inp[11]) ? node17538 : node17517;
												assign node17517 = (inp[7]) ? node17529 : node17518;
													assign node17518 = (inp[13]) ? node17524 : node17519;
														assign node17519 = (inp[10]) ? node17521 : 4'b0001;
															assign node17521 = (inp[12]) ? 4'b1001 : 4'b0101;
														assign node17524 = (inp[10]) ? 4'b1101 : node17525;
															assign node17525 = (inp[2]) ? 4'b0101 : 4'b1101;
													assign node17529 = (inp[2]) ? node17535 : node17530;
														assign node17530 = (inp[10]) ? node17532 : 4'b1001;
															assign node17532 = (inp[13]) ? 4'b0101 : 4'b0001;
														assign node17535 = (inp[10]) ? 4'b1001 : 4'b0001;
												assign node17538 = (inp[2]) ? node17550 : node17539;
													assign node17539 = (inp[13]) ? node17547 : node17540;
														assign node17540 = (inp[10]) ? node17544 : node17541;
															assign node17541 = (inp[12]) ? 4'b0001 : 4'b1001;
															assign node17544 = (inp[7]) ? 4'b0001 : 4'b0101;
														assign node17547 = (inp[10]) ? 4'b1000 : 4'b0101;
													assign node17550 = (inp[13]) ? node17558 : node17551;
														assign node17551 = (inp[7]) ? 4'b0000 : node17552;
															assign node17552 = (inp[12]) ? node17554 : 4'b1000;
																assign node17554 = (inp[10]) ? 4'b1000 : 4'b0000;
														assign node17558 = (inp[7]) ? node17564 : node17559;
															assign node17559 = (inp[10]) ? node17561 : 4'b1100;
																assign node17561 = (inp[12]) ? 4'b1100 : 4'b0100;
															assign node17564 = (inp[12]) ? 4'b1000 : node17565;
																assign node17565 = (inp[10]) ? 4'b0100 : 4'b1000;
											assign node17569 = (inp[2]) ? node17581 : node17570;
												assign node17570 = (inp[13]) ? node17576 : node17571;
													assign node17571 = (inp[12]) ? node17573 : 4'b1000;
														assign node17573 = (inp[7]) ? 4'b1000 : 4'b1100;
													assign node17576 = (inp[11]) ? 4'b0001 : node17577;
														assign node17577 = (inp[7]) ? 4'b0000 : 4'b0001;
												assign node17581 = (inp[13]) ? node17591 : node17582;
													assign node17582 = (inp[7]) ? node17584 : 4'b0001;
														assign node17584 = (inp[11]) ? 4'b0001 : node17585;
															assign node17585 = (inp[12]) ? 4'b1101 : node17586;
																assign node17586 = (inp[10]) ? 4'b0001 : 4'b0101;
													assign node17591 = (inp[7]) ? node17599 : node17592;
														assign node17592 = (inp[10]) ? node17596 : node17593;
															assign node17593 = (inp[11]) ? 4'b0101 : 4'b1001;
															assign node17596 = (inp[12]) ? 4'b0000 : 4'b1000;
														assign node17599 = (inp[11]) ? 4'b1001 : node17600;
															assign node17600 = (inp[12]) ? 4'b0001 : 4'b1001;
									assign node17604 = (inp[11]) ? node17704 : node17605;
										assign node17605 = (inp[2]) ? node17653 : node17606;
											assign node17606 = (inp[13]) ? node17630 : node17607;
												assign node17607 = (inp[4]) ? node17619 : node17608;
													assign node17608 = (inp[14]) ? node17612 : node17609;
														assign node17609 = (inp[10]) ? 4'b0001 : 4'b1001;
														assign node17612 = (inp[12]) ? node17614 : 4'b1000;
															assign node17614 = (inp[7]) ? node17616 : 4'b0100;
																assign node17616 = (inp[10]) ? 4'b0000 : 4'b1000;
													assign node17619 = (inp[12]) ? node17627 : node17620;
														assign node17620 = (inp[14]) ? 4'b0100 : node17621;
															assign node17621 = (inp[10]) ? 4'b1000 : node17622;
																assign node17622 = (inp[7]) ? 4'b0000 : 4'b0100;
														assign node17627 = (inp[7]) ? 4'b1000 : 4'b0001;
												assign node17630 = (inp[4]) ? node17642 : node17631;
													assign node17631 = (inp[10]) ? node17639 : node17632;
														assign node17632 = (inp[7]) ? node17636 : node17633;
															assign node17633 = (inp[12]) ? 4'b0100 : 4'b0000;
															assign node17636 = (inp[14]) ? 4'b0100 : 4'b0101;
														assign node17639 = (inp[7]) ? 4'b0000 : 4'b1000;
													assign node17642 = (inp[14]) ? node17648 : node17643;
														assign node17643 = (inp[12]) ? 4'b1000 : node17644;
															assign node17644 = (inp[7]) ? 4'b0100 : 4'b1001;
														assign node17648 = (inp[10]) ? 4'b1001 : node17649;
															assign node17649 = (inp[12]) ? 4'b0001 : 4'b1001;
											assign node17653 = (inp[4]) ? node17679 : node17654;
												assign node17654 = (inp[13]) ? node17664 : node17655;
													assign node17655 = (inp[14]) ? node17659 : node17656;
														assign node17656 = (inp[12]) ? 4'b0001 : 4'b1001;
														assign node17659 = (inp[10]) ? node17661 : 4'b1001;
															assign node17661 = (inp[12]) ? 4'b1001 : 4'b0001;
													assign node17664 = (inp[10]) ? node17672 : node17665;
														assign node17665 = (inp[12]) ? node17669 : node17666;
															assign node17666 = (inp[7]) ? 4'b1001 : 4'b1101;
															assign node17669 = (inp[7]) ? 4'b0001 : 4'b0101;
														assign node17672 = (inp[12]) ? 4'b1001 : node17673;
															assign node17673 = (inp[7]) ? 4'b0101 : node17674;
																assign node17674 = (inp[14]) ? 4'b0000 : 4'b0001;
												assign node17679 = (inp[14]) ? node17687 : node17680;
													assign node17680 = (inp[13]) ? node17684 : node17681;
														assign node17681 = (inp[7]) ? 4'b1101 : 4'b1001;
														assign node17684 = (inp[7]) ? 4'b0001 : 4'b0101;
													assign node17687 = (inp[10]) ? node17695 : node17688;
														assign node17688 = (inp[13]) ? node17690 : 4'b0101;
															assign node17690 = (inp[7]) ? 4'b0000 : node17691;
																assign node17691 = (inp[12]) ? 4'b0100 : 4'b0000;
														assign node17695 = (inp[7]) ? node17697 : 4'b0000;
															assign node17697 = (inp[12]) ? node17701 : node17698;
																assign node17698 = (inp[13]) ? 4'b0000 : 4'b1000;
																assign node17701 = (inp[13]) ? 4'b1000 : 4'b0000;
										assign node17704 = (inp[13]) ? node17732 : node17705;
											assign node17705 = (inp[10]) ? node17721 : node17706;
												assign node17706 = (inp[4]) ? node17714 : node17707;
													assign node17707 = (inp[2]) ? 4'b1000 : node17708;
														assign node17708 = (inp[14]) ? node17710 : 4'b1000;
															assign node17710 = (inp[7]) ? 4'b0000 : 4'b0100;
													assign node17714 = (inp[7]) ? node17718 : node17715;
														assign node17715 = (inp[2]) ? 4'b0000 : 4'b0100;
														assign node17718 = (inp[2]) ? 4'b1100 : 4'b0000;
												assign node17721 = (inp[4]) ? node17727 : node17722;
													assign node17722 = (inp[7]) ? 4'b1000 : node17723;
														assign node17723 = (inp[2]) ? 4'b0100 : 4'b1100;
													assign node17727 = (inp[7]) ? node17729 : 4'b1000;
														assign node17729 = (inp[2]) ? 4'b1000 : 4'b0100;
											assign node17732 = (inp[10]) ? node17750 : node17733;
												assign node17733 = (inp[4]) ? node17741 : node17734;
													assign node17734 = (inp[2]) ? node17738 : node17735;
														assign node17735 = (inp[7]) ? 4'b0100 : 4'b0000;
														assign node17738 = (inp[7]) ? 4'b1000 : 4'b1100;
													assign node17741 = (inp[12]) ? node17747 : node17742;
														assign node17742 = (inp[2]) ? 4'b0000 : node17743;
															assign node17743 = (inp[7]) ? 4'b0000 : 4'b0100;
														assign node17747 = (inp[2]) ? 4'b0000 : 4'b1000;
												assign node17750 = (inp[7]) ? node17752 : 4'b0000;
													assign node17752 = (inp[2]) ? node17754 : 4'b0000;
														assign node17754 = (inp[4]) ? 4'b0000 : 4'b0100;
								assign node17757 = (inp[4]) ? node17901 : node17758;
									assign node17758 = (inp[11]) ? node17834 : node17759;
										assign node17759 = (inp[12]) ? node17787 : node17760;
											assign node17760 = (inp[1]) ? node17772 : node17761;
												assign node17761 = (inp[13]) ? node17769 : node17762;
													assign node17762 = (inp[14]) ? 4'b1000 : node17763;
														assign node17763 = (inp[7]) ? 4'b1001 : node17764;
															assign node17764 = (inp[2]) ? 4'b1001 : 4'b1000;
													assign node17769 = (inp[10]) ? 4'b0000 : 4'b1001;
												assign node17772 = (inp[10]) ? node17782 : node17773;
													assign node17773 = (inp[13]) ? 4'b0001 : node17774;
														assign node17774 = (inp[7]) ? node17778 : node17775;
															assign node17775 = (inp[2]) ? 4'b0001 : 4'b1000;
															assign node17778 = (inp[2]) ? 4'b0000 : 4'b0001;
													assign node17782 = (inp[7]) ? node17784 : 4'b1000;
														assign node17784 = (inp[13]) ? 4'b1001 : 4'b0001;
											assign node17787 = (inp[2]) ? node17807 : node17788;
												assign node17788 = (inp[10]) ? node17794 : node17789;
													assign node17789 = (inp[1]) ? node17791 : 4'b0001;
														assign node17791 = (inp[14]) ? 4'b0000 : 4'b0001;
													assign node17794 = (inp[7]) ? node17800 : node17795;
														assign node17795 = (inp[1]) ? node17797 : 4'b0000;
															assign node17797 = (inp[13]) ? 4'b0000 : 4'b1000;
														assign node17800 = (inp[1]) ? node17804 : node17801;
															assign node17801 = (inp[13]) ? 4'b0001 : 4'b0000;
															assign node17804 = (inp[14]) ? 4'b0000 : 4'b0001;
												assign node17807 = (inp[13]) ? node17825 : node17808;
													assign node17808 = (inp[10]) ? node17816 : node17809;
														assign node17809 = (inp[1]) ? node17811 : 4'b0000;
															assign node17811 = (inp[14]) ? 4'b1000 : node17812;
																assign node17812 = (inp[7]) ? 4'b1000 : 4'b0000;
														assign node17816 = (inp[7]) ? 4'b0000 : node17817;
															assign node17817 = (inp[1]) ? node17821 : node17818;
																assign node17818 = (inp[14]) ? 4'b1000 : 4'b1001;
																assign node17821 = (inp[14]) ? 4'b0001 : 4'b0000;
													assign node17825 = (inp[10]) ? node17831 : node17826;
														assign node17826 = (inp[1]) ? 4'b0001 : node17827;
															assign node17827 = (inp[7]) ? 4'b1000 : 4'b0001;
														assign node17831 = (inp[1]) ? 4'b1000 : 4'b1001;
										assign node17834 = (inp[1]) ? node17876 : node17835;
											assign node17835 = (inp[2]) ? node17863 : node17836;
												assign node17836 = (inp[12]) ? node17846 : node17837;
													assign node17837 = (inp[13]) ? 4'b1001 : node17838;
														assign node17838 = (inp[10]) ? node17842 : node17839;
															assign node17839 = (inp[7]) ? 4'b0000 : 4'b0001;
															assign node17842 = (inp[14]) ? 4'b0000 : 4'b1001;
													assign node17846 = (inp[14]) ? node17852 : node17847;
														assign node17847 = (inp[10]) ? 4'b1001 : node17848;
															assign node17848 = (inp[13]) ? 4'b1001 : 4'b1000;
														assign node17852 = (inp[10]) ? node17858 : node17853;
															assign node17853 = (inp[7]) ? 4'b0000 : node17854;
																assign node17854 = (inp[13]) ? 4'b1001 : 4'b1000;
															assign node17858 = (inp[7]) ? node17860 : 4'b0000;
																assign node17860 = (inp[13]) ? 4'b1000 : 4'b1001;
												assign node17863 = (inp[13]) ? node17867 : node17864;
													assign node17864 = (inp[10]) ? 4'b0001 : 4'b1000;
													assign node17867 = (inp[7]) ? node17873 : node17868;
														assign node17868 = (inp[10]) ? 4'b0000 : node17869;
															assign node17869 = (inp[12]) ? 4'b1000 : 4'b0000;
														assign node17873 = (inp[14]) ? 4'b0001 : 4'b0000;
											assign node17876 = (inp[10]) ? node17894 : node17877;
												assign node17877 = (inp[13]) ? node17885 : node17878;
													assign node17878 = (inp[12]) ? node17882 : node17879;
														assign node17879 = (inp[2]) ? 4'b1000 : 4'b0000;
														assign node17882 = (inp[2]) ? 4'b0000 : 4'b1000;
													assign node17885 = (inp[7]) ? node17889 : node17886;
														assign node17886 = (inp[12]) ? 4'b0000 : 4'b1000;
														assign node17889 = (inp[12]) ? 4'b1000 : node17890;
															assign node17890 = (inp[14]) ? 4'b1000 : 4'b0000;
												assign node17894 = (inp[13]) ? 4'b0000 : node17895;
													assign node17895 = (inp[7]) ? node17897 : 4'b0000;
														assign node17897 = (inp[2]) ? 4'b1000 : 4'b0000;
									assign node17901 = (inp[13]) ? node17977 : node17902;
										assign node17902 = (inp[1]) ? node17948 : node17903;
											assign node17903 = (inp[2]) ? node17931 : node17904;
												assign node17904 = (inp[12]) ? node17916 : node17905;
													assign node17905 = (inp[7]) ? node17911 : node17906;
														assign node17906 = (inp[11]) ? 4'b0001 : node17907;
															assign node17907 = (inp[14]) ? 4'b0001 : 4'b0000;
														assign node17911 = (inp[10]) ? node17913 : 4'b0000;
															assign node17913 = (inp[14]) ? 4'b1000 : 4'b1001;
													assign node17916 = (inp[10]) ? node17924 : node17917;
														assign node17917 = (inp[7]) ? node17921 : node17918;
															assign node17918 = (inp[14]) ? 4'b1000 : 4'b1001;
															assign node17921 = (inp[11]) ? 4'b1001 : 4'b1000;
														assign node17924 = (inp[7]) ? node17928 : node17925;
															assign node17925 = (inp[11]) ? 4'b1000 : 4'b1001;
															assign node17928 = (inp[14]) ? 4'b0000 : 4'b0001;
												assign node17931 = (inp[12]) ? node17945 : node17932;
													assign node17932 = (inp[10]) ? node17938 : node17933;
														assign node17933 = (inp[14]) ? 4'b1000 : node17934;
															assign node17934 = (inp[7]) ? 4'b1000 : 4'b1001;
														assign node17938 = (inp[7]) ? node17942 : node17939;
															assign node17939 = (inp[11]) ? 4'b1000 : 4'b0000;
															assign node17942 = (inp[14]) ? 4'b0000 : 4'b0001;
													assign node17945 = (inp[11]) ? 4'b0000 : 4'b0001;
											assign node17948 = (inp[11]) ? node17966 : node17949;
												assign node17949 = (inp[7]) ? node17957 : node17950;
													assign node17950 = (inp[14]) ? 4'b0000 : node17951;
														assign node17951 = (inp[12]) ? node17953 : 4'b0001;
															assign node17953 = (inp[10]) ? 4'b0001 : 4'b0000;
													assign node17957 = (inp[12]) ? node17963 : node17958;
														assign node17958 = (inp[2]) ? 4'b0001 : node17959;
															assign node17959 = (inp[10]) ? 4'b1000 : 4'b0000;
														assign node17963 = (inp[10]) ? 4'b0001 : 4'b1001;
												assign node17966 = (inp[10]) ? 4'b0000 : node17967;
													assign node17967 = (inp[14]) ? 4'b0000 : node17968;
														assign node17968 = (inp[12]) ? node17972 : node17969;
															assign node17969 = (inp[7]) ? 4'b0000 : 4'b1000;
															assign node17972 = (inp[2]) ? 4'b1000 : 4'b0000;
										assign node17977 = (inp[11]) ? node18001 : node17978;
											assign node17978 = (inp[2]) ? node17992 : node17979;
												assign node17979 = (inp[1]) ? node17987 : node17980;
													assign node17980 = (inp[7]) ? 4'b0000 : node17981;
														assign node17981 = (inp[10]) ? node17983 : 4'b0001;
															assign node17983 = (inp[14]) ? 4'b0000 : 4'b0001;
													assign node17987 = (inp[10]) ? 4'b0000 : node17988;
														assign node17988 = (inp[7]) ? 4'b0001 : 4'b0000;
												assign node17992 = (inp[12]) ? 4'b0000 : node17993;
													assign node17993 = (inp[14]) ? 4'b0000 : node17994;
														assign node17994 = (inp[1]) ? node17996 : 4'b0000;
															assign node17996 = (inp[7]) ? 4'b0001 : 4'b0000;
											assign node18001 = (inp[1]) ? 4'b0000 : node18002;
												assign node18002 = (inp[10]) ? 4'b0000 : node18003;
													assign node18003 = (inp[7]) ? node18005 : 4'b0000;
														assign node18005 = (inp[12]) ? 4'b0001 : 4'b0000;
					assign node18010 = (inp[6]) ? node18012 : 4'b0000;
						assign node18012 = (inp[2]) ? node18342 : node18013;
							assign node18013 = (inp[5]) ? node18063 : node18014;
								assign node18014 = (inp[3]) ? node18016 : 4'b0000;
									assign node18016 = (inp[7]) ? 4'b0000 : node18017;
										assign node18017 = (inp[4]) ? node18027 : node18018;
											assign node18018 = (inp[13]) ? node18020 : 4'b0000;
												assign node18020 = (inp[12]) ? 4'b0000 : node18021;
													assign node18021 = (inp[11]) ? 4'b0000 : node18022;
														assign node18022 = (inp[10]) ? 4'b0001 : 4'b0000;
											assign node18027 = (inp[1]) ? node18047 : node18028;
												assign node18028 = (inp[11]) ? node18040 : node18029;
													assign node18029 = (inp[14]) ? node18031 : 4'b0001;
														assign node18031 = (inp[13]) ? node18037 : node18032;
															assign node18032 = (inp[12]) ? 4'b0000 : node18033;
																assign node18033 = (inp[10]) ? 4'b1000 : 4'b0000;
															assign node18037 = (inp[12]) ? 4'b1000 : 4'b0000;
													assign node18040 = (inp[13]) ? node18042 : 4'b0001;
														assign node18042 = (inp[10]) ? node18044 : 4'b1001;
															assign node18044 = (inp[12]) ? 4'b1001 : 4'b0001;
												assign node18047 = (inp[14]) ? node18057 : node18048;
													assign node18048 = (inp[12]) ? node18052 : node18049;
														assign node18049 = (inp[13]) ? 4'b0000 : 4'b1000;
														assign node18052 = (inp[13]) ? 4'b1000 : node18053;
															assign node18053 = (inp[10]) ? 4'b1000 : 4'b0000;
													assign node18057 = (inp[11]) ? node18059 : 4'b0001;
														assign node18059 = (inp[13]) ? 4'b0000 : 4'b1000;
								assign node18063 = (inp[1]) ? node18217 : node18064;
									assign node18064 = (inp[4]) ? node18134 : node18065;
										assign node18065 = (inp[13]) ? node18097 : node18066;
											assign node18066 = (inp[10]) ? node18080 : node18067;
												assign node18067 = (inp[7]) ? node18069 : 4'b0001;
													assign node18069 = (inp[12]) ? node18073 : node18070;
														assign node18070 = (inp[11]) ? 4'b1000 : 4'b0001;
														assign node18073 = (inp[11]) ? 4'b0001 : node18074;
															assign node18074 = (inp[3]) ? 4'b0001 : node18075;
																assign node18075 = (inp[14]) ? 4'b0000 : 4'b0001;
												assign node18080 = (inp[7]) ? node18090 : node18081;
													assign node18081 = (inp[12]) ? node18085 : node18082;
														assign node18082 = (inp[3]) ? 4'b0001 : 4'b1001;
														assign node18085 = (inp[14]) ? 4'b0000 : node18086;
															assign node18086 = (inp[3]) ? 4'b0000 : 4'b0001;
													assign node18090 = (inp[11]) ? node18094 : node18091;
														assign node18091 = (inp[3]) ? 4'b1001 : 4'b1000;
														assign node18094 = (inp[12]) ? 4'b0001 : 4'b1001;
											assign node18097 = (inp[12]) ? node18117 : node18098;
												assign node18098 = (inp[10]) ? node18106 : node18099;
													assign node18099 = (inp[3]) ? 4'b0001 : node18100;
														assign node18100 = (inp[11]) ? 4'b1001 : node18101;
															assign node18101 = (inp[14]) ? 4'b1000 : 4'b1001;
													assign node18106 = (inp[3]) ? node18114 : node18107;
														assign node18107 = (inp[7]) ? node18111 : node18108;
															assign node18108 = (inp[14]) ? 4'b0100 : 4'b0101;
															assign node18111 = (inp[14]) ? 4'b0000 : 4'b0001;
														assign node18114 = (inp[7]) ? 4'b1001 : 4'b1000;
												assign node18117 = (inp[3]) ? node18123 : node18118;
													assign node18118 = (inp[11]) ? 4'b1001 : node18119;
														assign node18119 = (inp[14]) ? 4'b1000 : 4'b1001;
													assign node18123 = (inp[7]) ? node18127 : node18124;
														assign node18124 = (inp[14]) ? 4'b1001 : 4'b1000;
														assign node18127 = (inp[10]) ? node18129 : 4'b0000;
															assign node18129 = (inp[14]) ? 4'b0001 : node18130;
																assign node18130 = (inp[11]) ? 4'b1001 : 4'b1000;
										assign node18134 = (inp[3]) ? node18178 : node18135;
											assign node18135 = (inp[14]) ? node18151 : node18136;
												assign node18136 = (inp[13]) ? node18142 : node18137;
													assign node18137 = (inp[12]) ? 4'b0101 : node18138;
														assign node18138 = (inp[7]) ? 4'b0001 : 4'b0000;
													assign node18142 = (inp[11]) ? 4'b1001 : node18143;
														assign node18143 = (inp[12]) ? 4'b0001 : node18144;
															assign node18144 = (inp[7]) ? node18146 : 4'b1001;
																assign node18146 = (inp[10]) ? 4'b0101 : 4'b1001;
												assign node18151 = (inp[11]) ? node18169 : node18152;
													assign node18152 = (inp[7]) ? node18160 : node18153;
														assign node18153 = (inp[13]) ? node18157 : node18154;
															assign node18154 = (inp[12]) ? 4'b0100 : 4'b1100;
															assign node18157 = (inp[10]) ? 4'b1001 : 4'b0001;
														assign node18160 = (inp[13]) ? node18164 : node18161;
															assign node18161 = (inp[12]) ? 4'b0000 : 4'b1000;
															assign node18164 = (inp[10]) ? node18166 : 4'b1000;
																assign node18166 = (inp[12]) ? 4'b1000 : 4'b0100;
													assign node18169 = (inp[13]) ? 4'b0000 : node18170;
														assign node18170 = (inp[7]) ? node18172 : 4'b0000;
															assign node18172 = (inp[12]) ? 4'b0001 : node18173;
																assign node18173 = (inp[10]) ? 4'b1001 : 4'b0001;
											assign node18178 = (inp[13]) ? node18202 : node18179;
												assign node18179 = (inp[10]) ? node18191 : node18180;
													assign node18180 = (inp[7]) ? node18188 : node18181;
														assign node18181 = (inp[12]) ? node18185 : node18182;
															assign node18182 = (inp[11]) ? 4'b0000 : 4'b1000;
															assign node18185 = (inp[11]) ? 4'b1001 : 4'b0001;
														assign node18188 = (inp[12]) ? 4'b0000 : 4'b1000;
													assign node18191 = (inp[11]) ? node18199 : node18192;
														assign node18192 = (inp[12]) ? 4'b1000 : node18193;
															assign node18193 = (inp[7]) ? 4'b0001 : node18194;
																assign node18194 = (inp[14]) ? 4'b0001 : 4'b1000;
														assign node18199 = (inp[7]) ? 4'b1000 : 4'b0000;
												assign node18202 = (inp[10]) ? node18210 : node18203;
													assign node18203 = (inp[11]) ? 4'b0001 : node18204;
														assign node18204 = (inp[7]) ? 4'b0000 : node18205;
															assign node18205 = (inp[12]) ? 4'b0001 : 4'b0000;
													assign node18210 = (inp[7]) ? node18212 : 4'b0000;
														assign node18212 = (inp[11]) ? 4'b0000 : node18213;
															assign node18213 = (inp[12]) ? 4'b0001 : 4'b0000;
									assign node18217 = (inp[11]) ? node18291 : node18218;
										assign node18218 = (inp[14]) ? node18256 : node18219;
											assign node18219 = (inp[3]) ? node18241 : node18220;
												assign node18220 = (inp[13]) ? node18230 : node18221;
													assign node18221 = (inp[12]) ? node18223 : 4'b1000;
														assign node18223 = (inp[10]) ? 4'b1100 : node18224;
															assign node18224 = (inp[4]) ? node18226 : 4'b0000;
																assign node18226 = (inp[7]) ? 4'b0000 : 4'b0100;
													assign node18230 = (inp[4]) ? node18234 : node18231;
														assign node18231 = (inp[7]) ? 4'b0000 : 4'b0100;
														assign node18234 = (inp[7]) ? node18236 : 4'b1001;
															assign node18236 = (inp[12]) ? 4'b1000 : node18237;
																assign node18237 = (inp[10]) ? 4'b0001 : 4'b0100;
												assign node18241 = (inp[12]) ? node18247 : node18242;
													assign node18242 = (inp[13]) ? 4'b0000 : node18243;
														assign node18243 = (inp[10]) ? 4'b0001 : 4'b0000;
													assign node18247 = (inp[4]) ? 4'b0000 : node18248;
														assign node18248 = (inp[13]) ? node18250 : 4'b0001;
															assign node18250 = (inp[10]) ? node18252 : 4'b0001;
																assign node18252 = (inp[7]) ? 4'b1001 : 4'b1000;
											assign node18256 = (inp[3]) ? node18272 : node18257;
												assign node18257 = (inp[13]) ? node18265 : node18258;
													assign node18258 = (inp[7]) ? node18262 : node18259;
														assign node18259 = (inp[4]) ? 4'b0101 : 4'b0001;
														assign node18262 = (inp[12]) ? 4'b0001 : 4'b1001;
													assign node18265 = (inp[4]) ? node18267 : 4'b1001;
														assign node18267 = (inp[7]) ? 4'b0001 : node18268;
															assign node18268 = (inp[10]) ? 4'b1001 : 4'b0001;
												assign node18272 = (inp[13]) ? node18280 : node18273;
													assign node18273 = (inp[10]) ? node18277 : node18274;
														assign node18274 = (inp[12]) ? 4'b0001 : 4'b1001;
														assign node18277 = (inp[7]) ? 4'b0001 : 4'b1000;
													assign node18280 = (inp[7]) ? node18288 : node18281;
														assign node18281 = (inp[10]) ? node18283 : 4'b0000;
															assign node18283 = (inp[4]) ? 4'b0000 : node18284;
																assign node18284 = (inp[12]) ? 4'b1000 : 4'b0000;
														assign node18288 = (inp[4]) ? 4'b0001 : 4'b0000;
										assign node18291 = (inp[13]) ? node18323 : node18292;
											assign node18292 = (inp[4]) ? node18308 : node18293;
												assign node18293 = (inp[10]) ? node18303 : node18294;
													assign node18294 = (inp[12]) ? node18300 : node18295;
														assign node18295 = (inp[3]) ? node18297 : 4'b1000;
															assign node18297 = (inp[7]) ? 4'b1000 : 4'b0000;
														assign node18300 = (inp[3]) ? 4'b1000 : 4'b0000;
													assign node18303 = (inp[3]) ? node18305 : 4'b1000;
														assign node18305 = (inp[7]) ? 4'b0000 : 4'b1000;
												assign node18308 = (inp[3]) ? node18314 : node18309;
													assign node18309 = (inp[7]) ? 4'b1000 : node18310;
														assign node18310 = (inp[12]) ? 4'b0100 : 4'b1100;
													assign node18314 = (inp[10]) ? 4'b0000 : node18315;
														assign node18315 = (inp[7]) ? node18319 : node18316;
															assign node18316 = (inp[12]) ? 4'b1000 : 4'b0000;
															assign node18319 = (inp[12]) ? 4'b0000 : 4'b1000;
											assign node18323 = (inp[10]) ? node18335 : node18324;
												assign node18324 = (inp[3]) ? node18328 : node18325;
													assign node18325 = (inp[12]) ? 4'b1000 : 4'b0100;
													assign node18328 = (inp[7]) ? node18330 : 4'b0000;
														assign node18330 = (inp[4]) ? 4'b0000 : node18331;
															assign node18331 = (inp[12]) ? 4'b0000 : 4'b1000;
												assign node18335 = (inp[7]) ? 4'b0000 : node18336;
													assign node18336 = (inp[3]) ? 4'b0000 : node18337;
														assign node18337 = (inp[4]) ? 4'b0000 : 4'b0100;
							assign node18342 = (inp[5]) ? node18344 : 4'b0000;
								assign node18344 = (inp[3]) ? node18346 : 4'b0000;
									assign node18346 = (inp[7]) ? node18390 : node18347;
										assign node18347 = (inp[4]) ? node18359 : node18348;
											assign node18348 = (inp[10]) ? node18350 : 4'b0000;
												assign node18350 = (inp[13]) ? node18352 : 4'b0000;
													assign node18352 = (inp[1]) ? node18354 : 4'b0001;
														assign node18354 = (inp[14]) ? node18356 : 4'b0000;
															assign node18356 = (inp[11]) ? 4'b0000 : 4'b0001;
											assign node18359 = (inp[13]) ? node18379 : node18360;
												assign node18360 = (inp[1]) ? node18372 : node18361;
													assign node18361 = (inp[11]) ? node18367 : node18362;
														assign node18362 = (inp[12]) ? 4'b0001 : node18363;
															assign node18363 = (inp[10]) ? 4'b1001 : 4'b0001;
														assign node18367 = (inp[12]) ? 4'b0001 : node18368;
															assign node18368 = (inp[10]) ? 4'b0000 : 4'b0001;
													assign node18372 = (inp[10]) ? node18376 : node18373;
														assign node18373 = (inp[12]) ? 4'b0000 : 4'b1000;
														assign node18376 = (inp[11]) ? 4'b0000 : 4'b0001;
												assign node18379 = (inp[1]) ? 4'b0000 : node18380;
													assign node18380 = (inp[11]) ? 4'b0000 : node18381;
														assign node18381 = (inp[10]) ? node18385 : node18382;
															assign node18382 = (inp[14]) ? 4'b0001 : 4'b0000;
															assign node18385 = (inp[14]) ? 4'b0000 : 4'b0001;
										assign node18390 = (inp[1]) ? 4'b0000 : node18391;
											assign node18391 = (inp[10]) ? node18393 : 4'b0000;
												assign node18393 = (inp[13]) ? node18395 : 4'b0000;
													assign node18395 = (inp[11]) ? 4'b0000 : node18396;
														assign node18396 = (inp[4]) ? node18398 : 4'b0000;
															assign node18398 = (inp[14]) ? 4'b0000 : 4'b0001;

endmodule