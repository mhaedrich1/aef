module dtc_split5_bm39 (
	input  wire [14-1:0] inp,
	output wire [14-1:0] outp
);

	wire [14-1:0] node1;
	wire [14-1:0] node3;
	wire [14-1:0] node4;
	wire [14-1:0] node5;
	wire [14-1:0] node6;
	wire [14-1:0] node7;
	wire [14-1:0] node8;
	wire [14-1:0] node9;
	wire [14-1:0] node11;
	wire [14-1:0] node12;
	wire [14-1:0] node13;
	wire [14-1:0] node14;
	wire [14-1:0] node17;
	wire [14-1:0] node20;
	wire [14-1:0] node21;
	wire [14-1:0] node24;
	wire [14-1:0] node27;
	wire [14-1:0] node28;
	wire [14-1:0] node29;
	wire [14-1:0] node32;
	wire [14-1:0] node35;
	wire [14-1:0] node36;
	wire [14-1:0] node39;
	wire [14-1:0] node42;
	wire [14-1:0] node43;
	wire [14-1:0] node44;
	wire [14-1:0] node45;
	wire [14-1:0] node46;
	wire [14-1:0] node50;
	wire [14-1:0] node53;
	wire [14-1:0] node54;
	wire [14-1:0] node57;
	wire [14-1:0] node58;
	wire [14-1:0] node62;
	wire [14-1:0] node63;
	wire [14-1:0] node65;
	wire [14-1:0] node67;
	wire [14-1:0] node70;
	wire [14-1:0] node71;
	wire [14-1:0] node72;
	wire [14-1:0] node76;
	wire [14-1:0] node78;
	wire [14-1:0] node81;
	wire [14-1:0] node82;
	wire [14-1:0] node83;
	wire [14-1:0] node84;
	wire [14-1:0] node85;
	wire [14-1:0] node88;
	wire [14-1:0] node91;
	wire [14-1:0] node92;
	wire [14-1:0] node94;
	wire [14-1:0] node97;
	wire [14-1:0] node98;
	wire [14-1:0] node101;
	wire [14-1:0] node104;
	wire [14-1:0] node105;
	wire [14-1:0] node106;
	wire [14-1:0] node107;
	wire [14-1:0] node110;
	wire [14-1:0] node113;
	wire [14-1:0] node116;
	wire [14-1:0] node117;
	wire [14-1:0] node118;
	wire [14-1:0] node122;
	wire [14-1:0] node124;
	wire [14-1:0] node127;
	wire [14-1:0] node128;
	wire [14-1:0] node129;
	wire [14-1:0] node130;
	wire [14-1:0] node131;
	wire [14-1:0] node135;
	wire [14-1:0] node136;
	wire [14-1:0] node139;
	wire [14-1:0] node142;
	wire [14-1:0] node143;
	wire [14-1:0] node145;
	wire [14-1:0] node149;
	wire [14-1:0] node150;
	wire [14-1:0] node151;
	wire [14-1:0] node153;
	wire [14-1:0] node157;
	wire [14-1:0] node158;
	wire [14-1:0] node159;
	wire [14-1:0] node163;
	wire [14-1:0] node165;
	wire [14-1:0] node168;
	wire [14-1:0] node169;
	wire [14-1:0] node170;
	wire [14-1:0] node171;
	wire [14-1:0] node172;
	wire [14-1:0] node174;
	wire [14-1:0] node177;
	wire [14-1:0] node178;
	wire [14-1:0] node180;
	wire [14-1:0] node183;
	wire [14-1:0] node184;
	wire [14-1:0] node187;
	wire [14-1:0] node190;
	wire [14-1:0] node191;
	wire [14-1:0] node192;
	wire [14-1:0] node193;
	wire [14-1:0] node196;
	wire [14-1:0] node199;
	wire [14-1:0] node200;
	wire [14-1:0] node203;
	wire [14-1:0] node206;
	wire [14-1:0] node207;
	wire [14-1:0] node209;
	wire [14-1:0] node212;
	wire [14-1:0] node213;
	wire [14-1:0] node217;
	wire [14-1:0] node218;
	wire [14-1:0] node219;
	wire [14-1:0] node220;
	wire [14-1:0] node223;
	wire [14-1:0] node224;
	wire [14-1:0] node228;
	wire [14-1:0] node229;
	wire [14-1:0] node231;
	wire [14-1:0] node234;
	wire [14-1:0] node237;
	wire [14-1:0] node239;
	wire [14-1:0] node241;
	wire [14-1:0] node242;
	wire [14-1:0] node245;
	wire [14-1:0] node248;
	wire [14-1:0] node249;
	wire [14-1:0] node250;
	wire [14-1:0] node252;
	wire [14-1:0] node253;
	wire [14-1:0] node254;
	wire [14-1:0] node258;
	wire [14-1:0] node259;
	wire [14-1:0] node263;
	wire [14-1:0] node264;
	wire [14-1:0] node265;
	wire [14-1:0] node266;
	wire [14-1:0] node269;
	wire [14-1:0] node272;
	wire [14-1:0] node273;
	wire [14-1:0] node279;
	wire [14-1:0] node280;
	wire [14-1:0] node281;
	wire [14-1:0] node282;
	wire [14-1:0] node283;
	wire [14-1:0] node284;
	wire [14-1:0] node285;
	wire [14-1:0] node286;
	wire [14-1:0] node290;
	wire [14-1:0] node291;
	wire [14-1:0] node294;
	wire [14-1:0] node297;
	wire [14-1:0] node298;
	wire [14-1:0] node299;
	wire [14-1:0] node302;
	wire [14-1:0] node306;
	wire [14-1:0] node307;
	wire [14-1:0] node308;
	wire [14-1:0] node311;
	wire [14-1:0] node312;
	wire [14-1:0] node316;
	wire [14-1:0] node317;
	wire [14-1:0] node318;
	wire [14-1:0] node322;
	wire [14-1:0] node324;
	wire [14-1:0] node327;
	wire [14-1:0] node328;
	wire [14-1:0] node329;
	wire [14-1:0] node330;
	wire [14-1:0] node333;
	wire [14-1:0] node334;
	wire [14-1:0] node337;
	wire [14-1:0] node340;
	wire [14-1:0] node341;
	wire [14-1:0] node343;
	wire [14-1:0] node347;
	wire [14-1:0] node348;
	wire [14-1:0] node349;
	wire [14-1:0] node350;
	wire [14-1:0] node353;
	wire [14-1:0] node356;
	wire [14-1:0] node359;
	wire [14-1:0] node360;
	wire [14-1:0] node361;
	wire [14-1:0] node366;
	wire [14-1:0] node367;
	wire [14-1:0] node368;
	wire [14-1:0] node369;
	wire [14-1:0] node370;
	wire [14-1:0] node371;
	wire [14-1:0] node374;
	wire [14-1:0] node378;
	wire [14-1:0] node379;
	wire [14-1:0] node380;
	wire [14-1:0] node385;
	wire [14-1:0] node386;
	wire [14-1:0] node387;
	wire [14-1:0] node388;
	wire [14-1:0] node392;
	wire [14-1:0] node393;
	wire [14-1:0] node397;
	wire [14-1:0] node398;
	wire [14-1:0] node399;
	wire [14-1:0] node402;
	wire [14-1:0] node405;
	wire [14-1:0] node408;
	wire [14-1:0] node409;
	wire [14-1:0] node410;
	wire [14-1:0] node411;
	wire [14-1:0] node415;
	wire [14-1:0] node416;
	wire [14-1:0] node417;
	wire [14-1:0] node421;
	wire [14-1:0] node422;
	wire [14-1:0] node425;
	wire [14-1:0] node428;
	wire [14-1:0] node429;
	wire [14-1:0] node430;
	wire [14-1:0] node432;
	wire [14-1:0] node437;
	wire [14-1:0] node439;
	wire [14-1:0] node440;
	wire [14-1:0] node441;
	wire [14-1:0] node442;
	wire [14-1:0] node443;
	wire [14-1:0] node444;
	wire [14-1:0] node452;
	wire [14-1:0] node453;
	wire [14-1:0] node454;
	wire [14-1:0] node455;
	wire [14-1:0] node456;
	wire [14-1:0] node457;
	wire [14-1:0] node458;
	wire [14-1:0] node461;
	wire [14-1:0] node462;
	wire [14-1:0] node465;
	wire [14-1:0] node466;
	wire [14-1:0] node470;
	wire [14-1:0] node471;
	wire [14-1:0] node472;
	wire [14-1:0] node475;
	wire [14-1:0] node477;
	wire [14-1:0] node480;
	wire [14-1:0] node481;
	wire [14-1:0] node483;
	wire [14-1:0] node486;
	wire [14-1:0] node487;
	wire [14-1:0] node491;
	wire [14-1:0] node492;
	wire [14-1:0] node493;
	wire [14-1:0] node494;
	wire [14-1:0] node497;
	wire [14-1:0] node498;
	wire [14-1:0] node501;
	wire [14-1:0] node504;
	wire [14-1:0] node505;
	wire [14-1:0] node506;
	wire [14-1:0] node510;
	wire [14-1:0] node513;
	wire [14-1:0] node514;
	wire [14-1:0] node515;
	wire [14-1:0] node519;
	wire [14-1:0] node520;
	wire [14-1:0] node521;
	wire [14-1:0] node525;
	wire [14-1:0] node527;
	wire [14-1:0] node530;
	wire [14-1:0] node531;
	wire [14-1:0] node532;
	wire [14-1:0] node533;
	wire [14-1:0] node534;
	wire [14-1:0] node536;
	wire [14-1:0] node539;
	wire [14-1:0] node540;
	wire [14-1:0] node543;
	wire [14-1:0] node546;
	wire [14-1:0] node547;
	wire [14-1:0] node548;
	wire [14-1:0] node551;
	wire [14-1:0] node555;
	wire [14-1:0] node556;
	wire [14-1:0] node557;
	wire [14-1:0] node558;
	wire [14-1:0] node561;
	wire [14-1:0] node564;
	wire [14-1:0] node565;
	wire [14-1:0] node568;
	wire [14-1:0] node571;
	wire [14-1:0] node572;
	wire [14-1:0] node573;
	wire [14-1:0] node576;
	wire [14-1:0] node579;
	wire [14-1:0] node583;
	wire [14-1:0] node584;
	wire [14-1:0] node585;
	wire [14-1:0] node586;
	wire [14-1:0] node587;
	wire [14-1:0] node592;
	wire [14-1:0] node593;
	wire [14-1:0] node594;
	wire [14-1:0] node595;
	wire [14-1:0] node598;
	wire [14-1:0] node601;
	wire [14-1:0] node602;
	wire [14-1:0] node603;
	wire [14-1:0] node606;
	wire [14-1:0] node609;
	wire [14-1:0] node610;
	wire [14-1:0] node613;
	wire [14-1:0] node616;
	wire [14-1:0] node617;
	wire [14-1:0] node618;
	wire [14-1:0] node619;
	wire [14-1:0] node623;
	wire [14-1:0] node625;
	wire [14-1:0] node629;
	wire [14-1:0] node631;
	wire [14-1:0] node633;
	wire [14-1:0] node635;
	wire [14-1:0] node639;
	wire [14-1:0] node640;
	wire [14-1:0] node641;
	wire [14-1:0] node642;
	wire [14-1:0] node643;
	wire [14-1:0] node644;
	wire [14-1:0] node645;
	wire [14-1:0] node646;
	wire [14-1:0] node648;
	wire [14-1:0] node649;
	wire [14-1:0] node652;
	wire [14-1:0] node655;
	wire [14-1:0] node656;
	wire [14-1:0] node658;
	wire [14-1:0] node661;
	wire [14-1:0] node662;
	wire [14-1:0] node666;
	wire [14-1:0] node667;
	wire [14-1:0] node668;
	wire [14-1:0] node669;
	wire [14-1:0] node672;
	wire [14-1:0] node675;
	wire [14-1:0] node676;
	wire [14-1:0] node680;
	wire [14-1:0] node681;
	wire [14-1:0] node682;
	wire [14-1:0] node686;
	wire [14-1:0] node687;
	wire [14-1:0] node690;
	wire [14-1:0] node693;
	wire [14-1:0] node694;
	wire [14-1:0] node695;
	wire [14-1:0] node696;
	wire [14-1:0] node697;
	wire [14-1:0] node701;
	wire [14-1:0] node702;
	wire [14-1:0] node705;
	wire [14-1:0] node708;
	wire [14-1:0] node709;
	wire [14-1:0] node711;
	wire [14-1:0] node715;
	wire [14-1:0] node716;
	wire [14-1:0] node717;
	wire [14-1:0] node720;
	wire [14-1:0] node721;
	wire [14-1:0] node724;
	wire [14-1:0] node728;
	wire [14-1:0] node729;
	wire [14-1:0] node730;
	wire [14-1:0] node731;
	wire [14-1:0] node732;
	wire [14-1:0] node733;
	wire [14-1:0] node736;
	wire [14-1:0] node739;
	wire [14-1:0] node742;
	wire [14-1:0] node743;
	wire [14-1:0] node744;
	wire [14-1:0] node748;
	wire [14-1:0] node751;
	wire [14-1:0] node752;
	wire [14-1:0] node755;
	wire [14-1:0] node756;
	wire [14-1:0] node757;
	wire [14-1:0] node760;
	wire [14-1:0] node763;
	wire [14-1:0] node765;
	wire [14-1:0] node768;
	wire [14-1:0] node769;
	wire [14-1:0] node770;
	wire [14-1:0] node772;
	wire [14-1:0] node773;
	wire [14-1:0] node776;
	wire [14-1:0] node779;
	wire [14-1:0] node780;
	wire [14-1:0] node782;
	wire [14-1:0] node787;
	wire [14-1:0] node788;
	wire [14-1:0] node789;
	wire [14-1:0] node790;
	wire [14-1:0] node791;
	wire [14-1:0] node792;
	wire [14-1:0] node793;
	wire [14-1:0] node796;
	wire [14-1:0] node799;
	wire [14-1:0] node802;
	wire [14-1:0] node803;
	wire [14-1:0] node805;
	wire [14-1:0] node808;
	wire [14-1:0] node809;
	wire [14-1:0] node812;
	wire [14-1:0] node815;
	wire [14-1:0] node816;
	wire [14-1:0] node817;
	wire [14-1:0] node820;
	wire [14-1:0] node823;
	wire [14-1:0] node824;
	wire [14-1:0] node825;
	wire [14-1:0] node828;
	wire [14-1:0] node831;
	wire [14-1:0] node832;
	wire [14-1:0] node835;
	wire [14-1:0] node838;
	wire [14-1:0] node840;
	wire [14-1:0] node841;
	wire [14-1:0] node842;
	wire [14-1:0] node843;
	wire [14-1:0] node850;
	wire [14-1:0] node851;
	wire [14-1:0] node853;
	wire [14-1:0] node854;
	wire [14-1:0] node855;
	wire [14-1:0] node856;
	wire [14-1:0] node857;
	wire [14-1:0] node858;
	wire [14-1:0] node861;
	wire [14-1:0] node864;
	wire [14-1:0] node866;
	wire [14-1:0] node869;
	wire [14-1:0] node870;
	wire [14-1:0] node873;
	wire [14-1:0] node874;
	wire [14-1:0] node877;
	wire [14-1:0] node880;
	wire [14-1:0] node881;
	wire [14-1:0] node882;
	wire [14-1:0] node884;
	wire [14-1:0] node887;
	wire [14-1:0] node891;
	wire [14-1:0] node892;
	wire [14-1:0] node893;
	wire [14-1:0] node894;
	wire [14-1:0] node896;
	wire [14-1:0] node899;
	wire [14-1:0] node902;
	wire [14-1:0] node904;
	wire [14-1:0] node907;
	wire [14-1:0] node908;
	wire [14-1:0] node909;
	wire [14-1:0] node915;
	wire [14-1:0] node916;
	wire [14-1:0] node917;
	wire [14-1:0] node918;
	wire [14-1:0] node919;
	wire [14-1:0] node920;
	wire [14-1:0] node921;
	wire [14-1:0] node922;
	wire [14-1:0] node925;
	wire [14-1:0] node926;
	wire [14-1:0] node936;
	wire [14-1:0] node937;
	wire [14-1:0] node938;
	wire [14-1:0] node939;
	wire [14-1:0] node940;
	wire [14-1:0] node941;
	wire [14-1:0] node942;
	wire [14-1:0] node943;
	wire [14-1:0] node944;
	wire [14-1:0] node946;
	wire [14-1:0] node947;
	wire [14-1:0] node949;
	wire [14-1:0] node952;
	wire [14-1:0] node953;
	wire [14-1:0] node957;
	wire [14-1:0] node958;
	wire [14-1:0] node959;
	wire [14-1:0] node961;
	wire [14-1:0] node964;
	wire [14-1:0] node966;
	wire [14-1:0] node969;
	wire [14-1:0] node970;
	wire [14-1:0] node971;
	wire [14-1:0] node974;
	wire [14-1:0] node977;
	wire [14-1:0] node979;
	wire [14-1:0] node982;
	wire [14-1:0] node983;
	wire [14-1:0] node984;
	wire [14-1:0] node985;
	wire [14-1:0] node988;
	wire [14-1:0] node990;
	wire [14-1:0] node993;
	wire [14-1:0] node994;
	wire [14-1:0] node997;
	wire [14-1:0] node999;
	wire [14-1:0] node1002;
	wire [14-1:0] node1003;
	wire [14-1:0] node1004;
	wire [14-1:0] node1006;
	wire [14-1:0] node1009;
	wire [14-1:0] node1010;
	wire [14-1:0] node1013;
	wire [14-1:0] node1016;
	wire [14-1:0] node1017;
	wire [14-1:0] node1018;
	wire [14-1:0] node1021;
	wire [14-1:0] node1024;
	wire [14-1:0] node1026;
	wire [14-1:0] node1029;
	wire [14-1:0] node1030;
	wire [14-1:0] node1031;
	wire [14-1:0] node1032;
	wire [14-1:0] node1034;
	wire [14-1:0] node1035;
	wire [14-1:0] node1038;
	wire [14-1:0] node1041;
	wire [14-1:0] node1042;
	wire [14-1:0] node1043;
	wire [14-1:0] node1046;
	wire [14-1:0] node1049;
	wire [14-1:0] node1052;
	wire [14-1:0] node1053;
	wire [14-1:0] node1054;
	wire [14-1:0] node1056;
	wire [14-1:0] node1059;
	wire [14-1:0] node1060;
	wire [14-1:0] node1063;
	wire [14-1:0] node1067;
	wire [14-1:0] node1068;
	wire [14-1:0] node1069;
	wire [14-1:0] node1070;
	wire [14-1:0] node1071;
	wire [14-1:0] node1074;
	wire [14-1:0] node1077;
	wire [14-1:0] node1078;
	wire [14-1:0] node1081;
	wire [14-1:0] node1084;
	wire [14-1:0] node1085;
	wire [14-1:0] node1086;
	wire [14-1:0] node1090;
	wire [14-1:0] node1092;
	wire [14-1:0] node1095;
	wire [14-1:0] node1096;
	wire [14-1:0] node1098;
	wire [14-1:0] node1099;
	wire [14-1:0] node1102;
	wire [14-1:0] node1105;
	wire [14-1:0] node1106;
	wire [14-1:0] node1107;
	wire [14-1:0] node1110;
	wire [14-1:0] node1113;
	wire [14-1:0] node1114;
	wire [14-1:0] node1118;
	wire [14-1:0] node1119;
	wire [14-1:0] node1120;
	wire [14-1:0] node1121;
	wire [14-1:0] node1122;
	wire [14-1:0] node1123;
	wire [14-1:0] node1126;
	wire [14-1:0] node1127;
	wire [14-1:0] node1130;
	wire [14-1:0] node1133;
	wire [14-1:0] node1134;
	wire [14-1:0] node1137;
	wire [14-1:0] node1140;
	wire [14-1:0] node1141;
	wire [14-1:0] node1142;
	wire [14-1:0] node1145;
	wire [14-1:0] node1146;
	wire [14-1:0] node1149;
	wire [14-1:0] node1152;
	wire [14-1:0] node1153;
	wire [14-1:0] node1154;
	wire [14-1:0] node1157;
	wire [14-1:0] node1160;
	wire [14-1:0] node1161;
	wire [14-1:0] node1164;
	wire [14-1:0] node1167;
	wire [14-1:0] node1168;
	wire [14-1:0] node1169;
	wire [14-1:0] node1170;
	wire [14-1:0] node1172;
	wire [14-1:0] node1175;
	wire [14-1:0] node1176;
	wire [14-1:0] node1180;
	wire [14-1:0] node1181;
	wire [14-1:0] node1183;
	wire [14-1:0] node1186;
	wire [14-1:0] node1187;
	wire [14-1:0] node1190;
	wire [14-1:0] node1195;
	wire [14-1:0] node1196;
	wire [14-1:0] node1197;
	wire [14-1:0] node1198;
	wire [14-1:0] node1199;
	wire [14-1:0] node1200;
	wire [14-1:0] node1202;
	wire [14-1:0] node1206;
	wire [14-1:0] node1207;
	wire [14-1:0] node1208;
	wire [14-1:0] node1211;
	wire [14-1:0] node1214;
	wire [14-1:0] node1215;
	wire [14-1:0] node1218;
	wire [14-1:0] node1221;
	wire [14-1:0] node1222;
	wire [14-1:0] node1223;
	wire [14-1:0] node1225;
	wire [14-1:0] node1228;
	wire [14-1:0] node1229;
	wire [14-1:0] node1233;
	wire [14-1:0] node1234;
	wire [14-1:0] node1235;
	wire [14-1:0] node1238;
	wire [14-1:0] node1241;
	wire [14-1:0] node1242;
	wire [14-1:0] node1245;
	wire [14-1:0] node1248;
	wire [14-1:0] node1249;
	wire [14-1:0] node1250;
	wire [14-1:0] node1251;
	wire [14-1:0] node1253;
	wire [14-1:0] node1256;
	wire [14-1:0] node1257;
	wire [14-1:0] node1260;
	wire [14-1:0] node1263;
	wire [14-1:0] node1264;
	wire [14-1:0] node1265;
	wire [14-1:0] node1268;
	wire [14-1:0] node1271;
	wire [14-1:0] node1272;
	wire [14-1:0] node1275;
	wire [14-1:0] node1278;
	wire [14-1:0] node1279;
	wire [14-1:0] node1280;
	wire [14-1:0] node1282;
	wire [14-1:0] node1285;
	wire [14-1:0] node1286;
	wire [14-1:0] node1289;
	wire [14-1:0] node1292;
	wire [14-1:0] node1293;
	wire [14-1:0] node1294;
	wire [14-1:0] node1297;
	wire [14-1:0] node1300;
	wire [14-1:0] node1301;
	wire [14-1:0] node1304;
	wire [14-1:0] node1307;
	wire [14-1:0] node1308;
	wire [14-1:0] node1309;
	wire [14-1:0] node1310;
	wire [14-1:0] node1312;
	wire [14-1:0] node1313;
	wire [14-1:0] node1316;
	wire [14-1:0] node1319;
	wire [14-1:0] node1320;
	wire [14-1:0] node1321;
	wire [14-1:0] node1325;
	wire [14-1:0] node1326;
	wire [14-1:0] node1330;
	wire [14-1:0] node1331;
	wire [14-1:0] node1332;
	wire [14-1:0] node1333;
	wire [14-1:0] node1336;
	wire [14-1:0] node1339;
	wire [14-1:0] node1340;
	wire [14-1:0] node1343;
	wire [14-1:0] node1346;
	wire [14-1:0] node1347;
	wire [14-1:0] node1348;
	wire [14-1:0] node1351;
	wire [14-1:0] node1354;
	wire [14-1:0] node1355;
	wire [14-1:0] node1358;
	wire [14-1:0] node1362;
	wire [14-1:0] node1363;
	wire [14-1:0] node1364;
	wire [14-1:0] node1365;
	wire [14-1:0] node1366;
	wire [14-1:0] node1367;
	wire [14-1:0] node1368;
	wire [14-1:0] node1369;
	wire [14-1:0] node1372;
	wire [14-1:0] node1374;
	wire [14-1:0] node1377;
	wire [14-1:0] node1378;
	wire [14-1:0] node1381;
	wire [14-1:0] node1382;
	wire [14-1:0] node1385;
	wire [14-1:0] node1388;
	wire [14-1:0] node1389;
	wire [14-1:0] node1390;
	wire [14-1:0] node1392;
	wire [14-1:0] node1395;
	wire [14-1:0] node1396;
	wire [14-1:0] node1399;
	wire [14-1:0] node1402;
	wire [14-1:0] node1403;
	wire [14-1:0] node1404;
	wire [14-1:0] node1407;
	wire [14-1:0] node1410;
	wire [14-1:0] node1412;
	wire [14-1:0] node1415;
	wire [14-1:0] node1416;
	wire [14-1:0] node1417;
	wire [14-1:0] node1418;
	wire [14-1:0] node1419;
	wire [14-1:0] node1422;
	wire [14-1:0] node1425;
	wire [14-1:0] node1427;
	wire [14-1:0] node1430;
	wire [14-1:0] node1431;
	wire [14-1:0] node1433;
	wire [14-1:0] node1436;
	wire [14-1:0] node1438;
	wire [14-1:0] node1442;
	wire [14-1:0] node1443;
	wire [14-1:0] node1444;
	wire [14-1:0] node1445;
	wire [14-1:0] node1447;
	wire [14-1:0] node1450;
	wire [14-1:0] node1451;
	wire [14-1:0] node1454;
	wire [14-1:0] node1457;
	wire [14-1:0] node1458;
	wire [14-1:0] node1459;
	wire [14-1:0] node1462;
	wire [14-1:0] node1465;
	wire [14-1:0] node1466;
	wire [14-1:0] node1469;
	wire [14-1:0] node1472;
	wire [14-1:0] node1473;
	wire [14-1:0] node1474;
	wire [14-1:0] node1475;
	wire [14-1:0] node1478;
	wire [14-1:0] node1481;
	wire [14-1:0] node1483;
	wire [14-1:0] node1486;
	wire [14-1:0] node1487;
	wire [14-1:0] node1488;
	wire [14-1:0] node1491;
	wire [14-1:0] node1494;
	wire [14-1:0] node1495;
	wire [14-1:0] node1498;
	wire [14-1:0] node1501;
	wire [14-1:0] node1502;
	wire [14-1:0] node1503;
	wire [14-1:0] node1504;
	wire [14-1:0] node1505;
	wire [14-1:0] node1506;
	wire [14-1:0] node1508;
	wire [14-1:0] node1511;
	wire [14-1:0] node1512;
	wire [14-1:0] node1516;
	wire [14-1:0] node1517;
	wire [14-1:0] node1518;
	wire [14-1:0] node1521;
	wire [14-1:0] node1524;
	wire [14-1:0] node1525;
	wire [14-1:0] node1528;
	wire [14-1:0] node1531;
	wire [14-1:0] node1532;
	wire [14-1:0] node1533;
	wire [14-1:0] node1534;
	wire [14-1:0] node1538;
	wire [14-1:0] node1539;
	wire [14-1:0] node1542;
	wire [14-1:0] node1545;
	wire [14-1:0] node1546;
	wire [14-1:0] node1547;
	wire [14-1:0] node1550;
	wire [14-1:0] node1553;
	wire [14-1:0] node1554;
	wire [14-1:0] node1557;
	wire [14-1:0] node1560;
	wire [14-1:0] node1561;
	wire [14-1:0] node1563;
	wire [14-1:0] node1564;
	wire [14-1:0] node1565;
	wire [14-1:0] node1568;
	wire [14-1:0] node1571;
	wire [14-1:0] node1572;
	wire [14-1:0] node1577;
	wire [14-1:0] node1579;
	wire [14-1:0] node1580;
	wire [14-1:0] node1581;
	wire [14-1:0] node1582;
	wire [14-1:0] node1588;
	wire [14-1:0] node1589;
	wire [14-1:0] node1590;
	wire [14-1:0] node1591;
	wire [14-1:0] node1592;
	wire [14-1:0] node1593;
	wire [14-1:0] node1594;
	wire [14-1:0] node1597;
	wire [14-1:0] node1598;
	wire [14-1:0] node1605;
	wire [14-1:0] node1606;
	wire [14-1:0] node1607;
	wire [14-1:0] node1608;
	wire [14-1:0] node1609;
	wire [14-1:0] node1610;
	wire [14-1:0] node1613;
	wire [14-1:0] node1616;
	wire [14-1:0] node1617;
	wire [14-1:0] node1620;
	wire [14-1:0] node1623;
	wire [14-1:0] node1624;
	wire [14-1:0] node1627;
	wire [14-1:0] node1628;
	wire [14-1:0] node1631;
	wire [14-1:0] node1634;
	wire [14-1:0] node1635;
	wire [14-1:0] node1636;
	wire [14-1:0] node1638;
	wire [14-1:0] node1641;
	wire [14-1:0] node1645;
	wire [14-1:0] node1646;
	wire [14-1:0] node1648;
	wire [14-1:0] node1650;
	wire [14-1:0] node1651;
	wire [14-1:0] node1656;
	wire [14-1:0] node1657;
	wire [14-1:0] node1658;
	wire [14-1:0] node1660;
	wire [14-1:0] node1662;
	wire [14-1:0] node1663;
	wire [14-1:0] node1669;
	wire [14-1:0] node1670;
	wire [14-1:0] node1671;
	wire [14-1:0] node1672;
	wire [14-1:0] node1673;
	wire [14-1:0] node1674;
	wire [14-1:0] node1675;
	wire [14-1:0] node1676;
	wire [14-1:0] node1677;
	wire [14-1:0] node1679;
	wire [14-1:0] node1683;
	wire [14-1:0] node1684;
	wire [14-1:0] node1685;
	wire [14-1:0] node1688;
	wire [14-1:0] node1691;
	wire [14-1:0] node1693;
	wire [14-1:0] node1696;
	wire [14-1:0] node1697;
	wire [14-1:0] node1698;
	wire [14-1:0] node1701;
	wire [14-1:0] node1702;
	wire [14-1:0] node1705;
	wire [14-1:0] node1708;
	wire [14-1:0] node1709;
	wire [14-1:0] node1710;
	wire [14-1:0] node1713;
	wire [14-1:0] node1716;
	wire [14-1:0] node1718;
	wire [14-1:0] node1721;
	wire [14-1:0] node1722;
	wire [14-1:0] node1723;
	wire [14-1:0] node1724;
	wire [14-1:0] node1727;
	wire [14-1:0] node1729;
	wire [14-1:0] node1732;
	wire [14-1:0] node1733;
	wire [14-1:0] node1734;
	wire [14-1:0] node1737;
	wire [14-1:0] node1740;
	wire [14-1:0] node1742;
	wire [14-1:0] node1745;
	wire [14-1:0] node1746;
	wire [14-1:0] node1748;
	wire [14-1:0] node1751;
	wire [14-1:0] node1752;
	wire [14-1:0] node1753;
	wire [14-1:0] node1756;
	wire [14-1:0] node1759;
	wire [14-1:0] node1761;
	wire [14-1:0] node1764;
	wire [14-1:0] node1765;
	wire [14-1:0] node1766;
	wire [14-1:0] node1767;
	wire [14-1:0] node1768;
	wire [14-1:0] node1769;
	wire [14-1:0] node1773;
	wire [14-1:0] node1774;
	wire [14-1:0] node1780;
	wire [14-1:0] node1781;
	wire [14-1:0] node1782;
	wire [14-1:0] node1783;
	wire [14-1:0] node1784;
	wire [14-1:0] node1787;
	wire [14-1:0] node1790;
	wire [14-1:0] node1791;
	wire [14-1:0] node1794;
	wire [14-1:0] node1797;
	wire [14-1:0] node1798;
	wire [14-1:0] node1800;
	wire [14-1:0] node1803;
	wire [14-1:0] node1804;
	wire [14-1:0] node1808;
	wire [14-1:0] node1809;
	wire [14-1:0] node1810;
	wire [14-1:0] node1811;
	wire [14-1:0] node1814;
	wire [14-1:0] node1817;
	wire [14-1:0] node1820;
	wire [14-1:0] node1822;
	wire [14-1:0] node1823;
	wire [14-1:0] node1826;
	wire [14-1:0] node1829;
	wire [14-1:0] node1830;
	wire [14-1:0] node1831;
	wire [14-1:0] node1832;
	wire [14-1:0] node1833;
	wire [14-1:0] node1834;
	wire [14-1:0] node1835;
	wire [14-1:0] node1838;
	wire [14-1:0] node1841;
	wire [14-1:0] node1844;
	wire [14-1:0] node1846;
	wire [14-1:0] node1848;
	wire [14-1:0] node1851;
	wire [14-1:0] node1852;
	wire [14-1:0] node1853;
	wire [14-1:0] node1854;
	wire [14-1:0] node1857;
	wire [14-1:0] node1862;
	wire [14-1:0] node1863;
	wire [14-1:0] node1864;
	wire [14-1:0] node1865;
	wire [14-1:0] node1868;
	wire [14-1:0] node1871;
	wire [14-1:0] node1872;
	wire [14-1:0] node1876;
	wire [14-1:0] node1877;
	wire [14-1:0] node1878;
	wire [14-1:0] node1881;
	wire [14-1:0] node1885;
	wire [14-1:0] node1886;
	wire [14-1:0] node1887;
	wire [14-1:0] node1888;
	wire [14-1:0] node1889;
	wire [14-1:0] node1890;
	wire [14-1:0] node1893;
	wire [14-1:0] node1896;
	wire [14-1:0] node1897;
	wire [14-1:0] node1900;
	wire [14-1:0] node1903;
	wire [14-1:0] node1904;
	wire [14-1:0] node1905;
	wire [14-1:0] node1908;
	wire [14-1:0] node1912;
	wire [14-1:0] node1914;
	wire [14-1:0] node1915;
	wire [14-1:0] node1920;
	wire [14-1:0] node1921;
	wire [14-1:0] node1922;
	wire [14-1:0] node1923;
	wire [14-1:0] node1924;
	wire [14-1:0] node1925;
	wire [14-1:0] node1926;
	wire [14-1:0] node1928;
	wire [14-1:0] node1936;
	wire [14-1:0] node1937;
	wire [14-1:0] node1938;
	wire [14-1:0] node1939;
	wire [14-1:0] node1940;
	wire [14-1:0] node1942;
	wire [14-1:0] node1945;
	wire [14-1:0] node1947;
	wire [14-1:0] node1950;
	wire [14-1:0] node1951;
	wire [14-1:0] node1952;
	wire [14-1:0] node1955;
	wire [14-1:0] node1958;
	wire [14-1:0] node1959;
	wire [14-1:0] node1962;
	wire [14-1:0] node1965;
	wire [14-1:0] node1966;
	wire [14-1:0] node1967;
	wire [14-1:0] node1968;
	wire [14-1:0] node1972;
	wire [14-1:0] node1973;
	wire [14-1:0] node1978;
	wire [14-1:0] node1979;
	wire [14-1:0] node1980;
	wire [14-1:0] node1981;
	wire [14-1:0] node1982;
	wire [14-1:0] node1985;
	wire [14-1:0] node1988;
	wire [14-1:0] node1989;
	wire [14-1:0] node1995;
	wire [14-1:0] node1996;
	wire [14-1:0] node1997;
	wire [14-1:0] node1998;
	wire [14-1:0] node1999;
	wire [14-1:0] node2001;
	wire [14-1:0] node2002;
	wire [14-1:0] node2004;
	wire [14-1:0] node2005;
	wire [14-1:0] node2010;
	wire [14-1:0] node2011;
	wire [14-1:0] node2012;
	wire [14-1:0] node2013;
	wire [14-1:0] node2016;
	wire [14-1:0] node2019;
	wire [14-1:0] node2020;
	wire [14-1:0] node2021;
	wire [14-1:0] node2024;
	wire [14-1:0] node2027;
	wire [14-1:0] node2029;
	wire [14-1:0] node2032;
	wire [14-1:0] node2033;
	wire [14-1:0] node2034;
	wire [14-1:0] node2036;
	wire [14-1:0] node2039;
	wire [14-1:0] node2041;
	wire [14-1:0] node2045;
	wire [14-1:0] node2046;
	wire [14-1:0] node2047;
	wire [14-1:0] node2048;
	wire [14-1:0] node2049;
	wire [14-1:0] node2050;
	wire [14-1:0] node2053;
	wire [14-1:0] node2056;
	wire [14-1:0] node2059;
	wire [14-1:0] node2060;
	wire [14-1:0] node2063;
	wire [14-1:0] node2064;
	wire [14-1:0] node2068;
	wire [14-1:0] node2069;
	wire [14-1:0] node2070;
	wire [14-1:0] node2071;
	wire [14-1:0] node2074;
	wire [14-1:0] node2077;
	wire [14-1:0] node2078;
	wire [14-1:0] node2081;
	wire [14-1:0] node2084;
	wire [14-1:0] node2085;
	wire [14-1:0] node2086;
	wire [14-1:0] node2091;
	wire [14-1:0] node2092;
	wire [14-1:0] node2093;
	wire [14-1:0] node2094;
	wire [14-1:0] node2095;
	wire [14-1:0] node2098;
	wire [14-1:0] node2102;
	wire [14-1:0] node2103;
	wire [14-1:0] node2104;
	wire [14-1:0] node2108;
	wire [14-1:0] node2110;
	wire [14-1:0] node2114;
	wire [14-1:0] node2115;
	wire [14-1:0] node2116;
	wire [14-1:0] node2117;
	wire [14-1:0] node2119;
	wire [14-1:0] node2120;
	wire [14-1:0] node2123;
	wire [14-1:0] node2126;
	wire [14-1:0] node2128;
	wire [14-1:0] node2129;
	wire [14-1:0] node2134;
	wire [14-1:0] node2135;
	wire [14-1:0] node2137;
	wire [14-1:0] node2139;
	wire [14-1:0] node2144;
	wire [14-1:0] node2145;
	wire [14-1:0] node2146;
	wire [14-1:0] node2147;
	wire [14-1:0] node2148;
	wire [14-1:0] node2149;
	wire [14-1:0] node2150;
	wire [14-1:0] node2151;
	wire [14-1:0] node2152;
	wire [14-1:0] node2153;
	wire [14-1:0] node2154;
	wire [14-1:0] node2157;
	wire [14-1:0] node2160;
	wire [14-1:0] node2161;
	wire [14-1:0] node2164;
	wire [14-1:0] node2167;
	wire [14-1:0] node2168;
	wire [14-1:0] node2170;
	wire [14-1:0] node2173;
	wire [14-1:0] node2174;
	wire [14-1:0] node2177;
	wire [14-1:0] node2180;
	wire [14-1:0] node2181;
	wire [14-1:0] node2182;
	wire [14-1:0] node2183;
	wire [14-1:0] node2186;
	wire [14-1:0] node2189;
	wire [14-1:0] node2190;
	wire [14-1:0] node2193;
	wire [14-1:0] node2196;
	wire [14-1:0] node2197;
	wire [14-1:0] node2198;
	wire [14-1:0] node2202;
	wire [14-1:0] node2203;
	wire [14-1:0] node2206;
	wire [14-1:0] node2209;
	wire [14-1:0] node2210;
	wire [14-1:0] node2211;
	wire [14-1:0] node2212;
	wire [14-1:0] node2214;
	wire [14-1:0] node2217;
	wire [14-1:0] node2218;
	wire [14-1:0] node2221;
	wire [14-1:0] node2224;
	wire [14-1:0] node2226;
	wire [14-1:0] node2227;
	wire [14-1:0] node2231;
	wire [14-1:0] node2233;
	wire [14-1:0] node2234;
	wire [14-1:0] node2238;
	wire [14-1:0] node2239;
	wire [14-1:0] node2240;
	wire [14-1:0] node2241;
	wire [14-1:0] node2242;
	wire [14-1:0] node2244;
	wire [14-1:0] node2247;
	wire [14-1:0] node2248;
	wire [14-1:0] node2251;
	wire [14-1:0] node2254;
	wire [14-1:0] node2255;
	wire [14-1:0] node2257;
	wire [14-1:0] node2260;
	wire [14-1:0] node2262;
	wire [14-1:0] node2265;
	wire [14-1:0] node2266;
	wire [14-1:0] node2267;
	wire [14-1:0] node2268;
	wire [14-1:0] node2272;
	wire [14-1:0] node2273;
	wire [14-1:0] node2277;
	wire [14-1:0] node2278;
	wire [14-1:0] node2279;
	wire [14-1:0] node2285;
	wire [14-1:0] node2286;
	wire [14-1:0] node2287;
	wire [14-1:0] node2288;
	wire [14-1:0] node2289;
	wire [14-1:0] node2290;
	wire [14-1:0] node2292;
	wire [14-1:0] node2295;
	wire [14-1:0] node2298;
	wire [14-1:0] node2299;
	wire [14-1:0] node2301;
	wire [14-1:0] node2304;
	wire [14-1:0] node2307;
	wire [14-1:0] node2308;
	wire [14-1:0] node2309;
	wire [14-1:0] node2312;
	wire [14-1:0] node2315;
	wire [14-1:0] node2316;
	wire [14-1:0] node2320;
	wire [14-1:0] node2321;
	wire [14-1:0] node2322;
	wire [14-1:0] node2325;
	wire [14-1:0] node2326;
	wire [14-1:0] node2329;
	wire [14-1:0] node2333;
	wire [14-1:0] node2334;
	wire [14-1:0] node2335;
	wire [14-1:0] node2337;
	wire [14-1:0] node2338;
	wire [14-1:0] node2343;
	wire [14-1:0] node2344;
	wire [14-1:0] node2345;
	wire [14-1:0] node2346;
	wire [14-1:0] node2349;
	wire [14-1:0] node2352;
	wire [14-1:0] node2353;
	wire [14-1:0] node2357;
	wire [14-1:0] node2358;
	wire [14-1:0] node2359;
	wire [14-1:0] node2363;
	wire [14-1:0] node2365;
	wire [14-1:0] node2368;
	wire [14-1:0] node2369;
	wire [14-1:0] node2370;
	wire [14-1:0] node2371;
	wire [14-1:0] node2372;
	wire [14-1:0] node2373;
	wire [14-1:0] node2374;
	wire [14-1:0] node2377;
	wire [14-1:0] node2378;
	wire [14-1:0] node2382;
	wire [14-1:0] node2383;
	wire [14-1:0] node2385;
	wire [14-1:0] node2388;
	wire [14-1:0] node2389;
	wire [14-1:0] node2393;
	wire [14-1:0] node2394;
	wire [14-1:0] node2395;
	wire [14-1:0] node2396;
	wire [14-1:0] node2399;
	wire [14-1:0] node2403;
	wire [14-1:0] node2405;
	wire [14-1:0] node2408;
	wire [14-1:0] node2409;
	wire [14-1:0] node2410;
	wire [14-1:0] node2411;
	wire [14-1:0] node2414;
	wire [14-1:0] node2415;
	wire [14-1:0] node2418;
	wire [14-1:0] node2421;
	wire [14-1:0] node2422;
	wire [14-1:0] node2424;
	wire [14-1:0] node2427;
	wire [14-1:0] node2428;
	wire [14-1:0] node2433;
	wire [14-1:0] node2434;
	wire [14-1:0] node2435;
	wire [14-1:0] node2436;
	wire [14-1:0] node2438;
	wire [14-1:0] node2441;
	wire [14-1:0] node2442;
	wire [14-1:0] node2445;
	wire [14-1:0] node2448;
	wire [14-1:0] node2449;
	wire [14-1:0] node2450;
	wire [14-1:0] node2453;
	wire [14-1:0] node2457;
	wire [14-1:0] node2458;
	wire [14-1:0] node2459;
	wire [14-1:0] node2461;
	wire [14-1:0] node2465;
	wire [14-1:0] node2467;
	wire [14-1:0] node2468;
	wire [14-1:0] node2473;
	wire [14-1:0] node2474;
	wire [14-1:0] node2475;
	wire [14-1:0] node2476;
	wire [14-1:0] node2477;
	wire [14-1:0] node2478;
	wire [14-1:0] node2479;
	wire [14-1:0] node2480;
	wire [14-1:0] node2482;
	wire [14-1:0] node2485;
	wire [14-1:0] node2486;
	wire [14-1:0] node2489;
	wire [14-1:0] node2492;
	wire [14-1:0] node2493;
	wire [14-1:0] node2494;
	wire [14-1:0] node2497;
	wire [14-1:0] node2500;
	wire [14-1:0] node2502;
	wire [14-1:0] node2505;
	wire [14-1:0] node2506;
	wire [14-1:0] node2507;
	wire [14-1:0] node2508;
	wire [14-1:0] node2511;
	wire [14-1:0] node2514;
	wire [14-1:0] node2515;
	wire [14-1:0] node2518;
	wire [14-1:0] node2521;
	wire [14-1:0] node2523;
	wire [14-1:0] node2524;
	wire [14-1:0] node2528;
	wire [14-1:0] node2530;
	wire [14-1:0] node2531;
	wire [14-1:0] node2532;
	wire [14-1:0] node2533;
	wire [14-1:0] node2536;
	wire [14-1:0] node2539;
	wire [14-1:0] node2540;
	wire [14-1:0] node2544;
	wire [14-1:0] node2545;
	wire [14-1:0] node2546;
	wire [14-1:0] node2551;
	wire [14-1:0] node2552;
	wire [14-1:0] node2553;
	wire [14-1:0] node2554;
	wire [14-1:0] node2555;
	wire [14-1:0] node2556;
	wire [14-1:0] node2559;
	wire [14-1:0] node2562;
	wire [14-1:0] node2565;
	wire [14-1:0] node2567;
	wire [14-1:0] node2568;
	wire [14-1:0] node2571;
	wire [14-1:0] node2574;
	wire [14-1:0] node2575;
	wire [14-1:0] node2577;
	wire [14-1:0] node2578;
	wire [14-1:0] node2581;
	wire [14-1:0] node2586;
	wire [14-1:0] node2587;
	wire [14-1:0] node2588;
	wire [14-1:0] node2589;
	wire [14-1:0] node2591;
	wire [14-1:0] node2593;
	wire [14-1:0] node2598;
	wire [14-1:0] node2599;
	wire [14-1:0] node2600;
	wire [14-1:0] node2601;
	wire [14-1:0] node2602;
	wire [14-1:0] node2604;
	wire [14-1:0] node2607;
	wire [14-1:0] node2608;
	wire [14-1:0] node2611;
	wire [14-1:0] node2614;
	wire [14-1:0] node2615;
	wire [14-1:0] node2616;
	wire [14-1:0] node2621;
	wire [14-1:0] node2622;
	wire [14-1:0] node2623;
	wire [14-1:0] node2624;
	wire [14-1:0] node2627;
	wire [14-1:0] node2630;
	wire [14-1:0] node2631;
	wire [14-1:0] node2634;
	wire [14-1:0] node2639;
	wire [14-1:0] node2640;
	wire [14-1:0] node2641;
	wire [14-1:0] node2642;
	wire [14-1:0] node2644;
	wire [14-1:0] node2646;
	wire [14-1:0] node2649;
	wire [14-1:0] node2650;
	wire [14-1:0] node2651;
	wire [14-1:0] node2652;
	wire [14-1:0] node2654;
	wire [14-1:0] node2657;
	wire [14-1:0] node2662;
	wire [14-1:0] node2663;
	wire [14-1:0] node2664;
	wire [14-1:0] node2666;
	wire [14-1:0] node2667;
	wire [14-1:0] node2674;
	wire [14-1:0] node2676;
	wire [14-1:0] node2677;
	wire [14-1:0] node2678;
	wire [14-1:0] node2679;
	wire [14-1:0] node2680;
	wire [14-1:0] node2681;
	wire [14-1:0] node2682;
	wire [14-1:0] node2683;
	wire [14-1:0] node2686;
	wire [14-1:0] node2689;
	wire [14-1:0] node2690;
	wire [14-1:0] node2693;
	wire [14-1:0] node2696;
	wire [14-1:0] node2697;
	wire [14-1:0] node2698;
	wire [14-1:0] node2701;
	wire [14-1:0] node2704;
	wire [14-1:0] node2706;
	wire [14-1:0] node2709;
	wire [14-1:0] node2710;
	wire [14-1:0] node2711;
	wire [14-1:0] node2713;
	wire [14-1:0] node2716;
	wire [14-1:0] node2717;
	wire [14-1:0] node2720;
	wire [14-1:0] node2724;
	wire [14-1:0] node2725;
	wire [14-1:0] node2726;
	wire [14-1:0] node2727;
	wire [14-1:0] node2729;
	wire [14-1:0] node2732;
	wire [14-1:0] node2733;
	wire [14-1:0] node2739;
	wire [14-1:0] node2741;
	wire [14-1:0] node2742;
	wire [14-1:0] node2743;
	wire [14-1:0] node2744;
	wire [14-1:0] node2745;
	wire [14-1:0] node2748;
	wire [14-1:0] node2751;
	wire [14-1:0] node2752;
	wire [14-1:0] node2756;
	wire [14-1:0] node2757;
	wire [14-1:0] node2758;
	wire [14-1:0] node2764;
	wire [14-1:0] node2766;
	wire [14-1:0] node2768;
	wire [14-1:0] node2770;
	wire [14-1:0] node2772;
	wire [14-1:0] node2774;
	wire [14-1:0] node2775;

	assign outp = (inp[8]) ? node936 : node1;
		assign node1 = (inp[13]) ? node3 : 14'b00000000000000;
			assign node3 = (inp[0]) ? node639 : node4;
				assign node4 = (inp[10]) ? node452 : node5;
					assign node5 = (inp[6]) ? node279 : node6;
						assign node6 = (inp[4]) ? node168 : node7;
							assign node7 = (inp[3]) ? node81 : node8;
								assign node8 = (inp[1]) ? node42 : node9;
									assign node9 = (inp[9]) ? node11 : 14'b00000000000001;
										assign node11 = (inp[7]) ? node27 : node12;
											assign node12 = (inp[2]) ? node20 : node13;
												assign node13 = (inp[5]) ? node17 : node14;
													assign node14 = (inp[12]) ? 14'b01000000000100 : 14'b00000000000001;
													assign node17 = (inp[12]) ? 14'b01000100000100 : 14'b01000100000110;
												assign node20 = (inp[5]) ? node24 : node21;
													assign node21 = (inp[12]) ? 14'b01100100000100 : 14'b01100100000110;
													assign node24 = (inp[12]) ? 14'b01000100000000 : 14'b01000100000010;
											assign node27 = (inp[2]) ? node35 : node28;
												assign node28 = (inp[12]) ? node32 : node29;
													assign node29 = (inp[5]) ? 14'b01000000000110 : 14'b00000000000010;
													assign node32 = (inp[5]) ? 14'b00000000000001 : 14'b00000000000000;
												assign node35 = (inp[5]) ? node39 : node36;
													assign node36 = (inp[12]) ? 14'b01100000000100 : 14'b01100000000110;
													assign node39 = (inp[11]) ? 14'b00000000000001 : 14'b01000000000000;
									assign node42 = (inp[9]) ? node62 : node43;
										assign node43 = (inp[7]) ? node53 : node44;
											assign node44 = (inp[12]) ? node50 : node45;
												assign node45 = (inp[11]) ? 14'b01010110100010 : node46;
													assign node46 = (inp[5]) ? 14'b01010110100110 : 14'b01110110100110;
												assign node50 = (inp[2]) ? 14'b01110110100100 : 14'b01010010100100;
											assign node53 = (inp[5]) ? node57 : node54;
												assign node54 = (inp[2]) ? 14'b01110010100110 : 14'b00010010100010;
												assign node57 = (inp[2]) ? 14'b00000000000001 : node58;
													assign node58 = (inp[12]) ? 14'b00000000000001 : 14'b01010010100110;
										assign node62 = (inp[12]) ? node70 : node63;
											assign node63 = (inp[7]) ? node65 : 14'b00000000000001;
												assign node65 = (inp[5]) ? node67 : 14'b01110010000110;
													assign node67 = (inp[2]) ? 14'b00000000000001 : 14'b01010010000110;
											assign node70 = (inp[5]) ? node76 : node71;
												assign node71 = (inp[2]) ? 14'b01110010000100 : node72;
													assign node72 = (inp[7]) ? 14'b00010010000000 : 14'b01010010000100;
												assign node76 = (inp[7]) ? node78 : 14'b01010110000100;
													assign node78 = (inp[2]) ? 14'b01010010000000 : 14'b00000000000001;
								assign node81 = (inp[1]) ? node127 : node82;
									assign node82 = (inp[7]) ? node104 : node83;
										assign node83 = (inp[5]) ? node91 : node84;
											assign node84 = (inp[2]) ? node88 : node85;
												assign node85 = (inp[12]) ? 14'b01010010110100 : 14'b00000000000001;
												assign node88 = (inp[12]) ? 14'b01110110010100 : 14'b01110110110110;
											assign node91 = (inp[2]) ? node97 : node92;
												assign node92 = (inp[9]) ? node94 : 14'b01010110110110;
													assign node94 = (inp[12]) ? 14'b01010110010100 : 14'b01010110010110;
												assign node97 = (inp[12]) ? node101 : node98;
													assign node98 = (inp[9]) ? 14'b01010110010010 : 14'b01010110110010;
													assign node101 = (inp[9]) ? 14'b01010110010000 : 14'b01010110110000;
										assign node104 = (inp[5]) ? node116 : node105;
											assign node105 = (inp[2]) ? node113 : node106;
												assign node106 = (inp[9]) ? node110 : node107;
													assign node107 = (inp[12]) ? 14'b00010010110000 : 14'b00010010110010;
													assign node110 = (inp[12]) ? 14'b00010010010000 : 14'b00010010010010;
												assign node113 = (inp[9]) ? 14'b01110010010100 : 14'b01110010110100;
											assign node116 = (inp[12]) ? node122 : node117;
												assign node117 = (inp[2]) ? 14'b00000000000001 : node118;
													assign node118 = (inp[9]) ? 14'b01010010010110 : 14'b01010010110110;
												assign node122 = (inp[2]) ? node124 : 14'b00000000000001;
													assign node124 = (inp[9]) ? 14'b01010010010000 : 14'b01010010110000;
									assign node127 = (inp[9]) ? node149 : node128;
										assign node128 = (inp[2]) ? node142 : node129;
											assign node129 = (inp[7]) ? node135 : node130;
												assign node130 = (inp[5]) ? 14'b01000110100110 : node131;
													assign node131 = (inp[12]) ? 14'b01000010100100 : 14'b00000000000001;
												assign node135 = (inp[12]) ? node139 : node136;
													assign node136 = (inp[5]) ? 14'b01000010100110 : 14'b00000010100010;
													assign node139 = (inp[5]) ? 14'b00000000000001 : 14'b00000010100000;
											assign node142 = (inp[5]) ? 14'b01000010100000 : node143;
												assign node143 = (inp[7]) ? node145 : 14'b01100110100100;
													assign node145 = (inp[12]) ? 14'b01100010100100 : 14'b01100010100110;
										assign node149 = (inp[12]) ? node157 : node150;
											assign node150 = (inp[7]) ? 14'b01000010000110 : node151;
												assign node151 = (inp[5]) ? node153 : 14'b01100110000110;
													assign node153 = (inp[2]) ? 14'b01000110000010 : 14'b01000110000110;
											assign node157 = (inp[7]) ? node163 : node158;
												assign node158 = (inp[2]) ? 14'b01100110000100 : node159;
													assign node159 = (inp[5]) ? 14'b01000110000100 : 14'b01000010000100;
												assign node163 = (inp[2]) ? node165 : 14'b00000010000000;
													assign node165 = (inp[5]) ? 14'b01000010000000 : 14'b01100010000100;
							assign node168 = (inp[2]) ? node248 : node169;
								assign node169 = (inp[5]) ? node217 : node170;
									assign node170 = (inp[3]) ? node190 : node171;
										assign node171 = (inp[1]) ? node177 : node172;
											assign node172 = (inp[9]) ? node174 : 14'b00000000000001;
												assign node174 = (inp[7]) ? 14'b00100000000110 : 14'b00100100000100;
											assign node177 = (inp[9]) ? node183 : node178;
												assign node178 = (inp[12]) ? node180 : 14'b00110110100110;
													assign node180 = (inp[7]) ? 14'b00110010100100 : 14'b00110110100100;
												assign node183 = (inp[12]) ? node187 : node184;
													assign node184 = (inp[11]) ? 14'b00110010000110 : 14'b00110110000110;
													assign node187 = (inp[7]) ? 14'b00110010000100 : 14'b00110110000100;
										assign node190 = (inp[1]) ? node206 : node191;
											assign node191 = (inp[7]) ? node199 : node192;
												assign node192 = (inp[12]) ? node196 : node193;
													assign node193 = (inp[9]) ? 14'b00110110010110 : 14'b00110110110110;
													assign node196 = (inp[9]) ? 14'b00110110010100 : 14'b00110110110100;
												assign node199 = (inp[9]) ? node203 : node200;
													assign node200 = (inp[11]) ? 14'b00110010110100 : 14'b00110010110110;
													assign node203 = (inp[12]) ? 14'b00110010010100 : 14'b00110010010110;
											assign node206 = (inp[12]) ? node212 : node207;
												assign node207 = (inp[9]) ? node209 : 14'b00100110100110;
													assign node209 = (inp[7]) ? 14'b00100010000110 : 14'b00100110000110;
												assign node212 = (inp[7]) ? 14'b00100010000100 : node213;
													assign node213 = (inp[11]) ? 14'b00100110100100 : 14'b00100110000100;
									assign node217 = (inp[12]) ? node237 : node218;
										assign node218 = (inp[3]) ? node228 : node219;
											assign node219 = (inp[1]) ? node223 : node220;
												assign node220 = (inp[9]) ? 14'b00000000000110 : 14'b00000000000001;
												assign node223 = (inp[9]) ? 14'b00010010000110 : node224;
													assign node224 = (inp[7]) ? 14'b00010010100110 : 14'b00010110100110;
											assign node228 = (inp[1]) ? node234 : node229;
												assign node229 = (inp[7]) ? node231 : 14'b00010110110110;
													assign node231 = (inp[9]) ? 14'b00010010010110 : 14'b00010010110110;
												assign node234 = (inp[11]) ? 14'b00000010100110 : 14'b00000110100110;
										assign node237 = (inp[7]) ? node239 : 14'b00000000000001;
											assign node239 = (inp[1]) ? node241 : 14'b00000000000001;
												assign node241 = (inp[3]) ? node245 : node242;
													assign node242 = (inp[9]) ? 14'b00010010000100 : 14'b00010010100100;
													assign node245 = (inp[9]) ? 14'b00000010000100 : 14'b00000010100100;
								assign node248 = (inp[7]) ? 14'b00000000000001 : node249;
									assign node249 = (inp[12]) ? node263 : node250;
										assign node250 = (inp[5]) ? node252 : 14'b00000000000001;
											assign node252 = (inp[3]) ? node258 : node253;
												assign node253 = (inp[1]) ? 14'b01010010100010 : node254;
													assign node254 = (inp[9]) ? 14'b01000000000010 : 14'b00000000000001;
												assign node258 = (inp[1]) ? 14'b01000010000010 : node259;
													assign node259 = (inp[9]) ? 14'b01010010010010 : 14'b01010010110010;
										assign node263 = (inp[5]) ? 14'b00000000000001 : node264;
											assign node264 = (inp[3]) ? node272 : node265;
												assign node265 = (inp[1]) ? node269 : node266;
													assign node266 = (inp[9]) ? 14'b00000100000100 : 14'b00000000000001;
													assign node269 = (inp[9]) ? 14'b00010110000100 : 14'b00010110100100;
												assign node272 = (inp[1]) ? 14'b00000110000100 : node273;
													assign node273 = (inp[11]) ? 14'b00010110110100 : 14'b00010110010100;
						assign node279 = (inp[3]) ? node437 : node280;
							assign node280 = (inp[12]) ? node366 : node281;
								assign node281 = (inp[1]) ? node327 : node282;
									assign node282 = (inp[9]) ? node306 : node283;
										assign node283 = (inp[7]) ? node297 : node284;
											assign node284 = (inp[5]) ? node290 : node285;
												assign node285 = (inp[2]) ? 14'b01110100110110 : node286;
													assign node286 = (inp[4]) ? 14'b00110100110110 : 14'b00000000000001;
												assign node290 = (inp[2]) ? node294 : node291;
													assign node291 = (inp[4]) ? 14'b00010100110110 : 14'b01010100110110;
													assign node294 = (inp[4]) ? 14'b01010000110010 : 14'b01010100110010;
											assign node297 = (inp[2]) ? 14'b00000000000001 : node298;
												assign node298 = (inp[4]) ? node302 : node299;
													assign node299 = (inp[5]) ? 14'b01010000110110 : 14'b00010000110010;
													assign node302 = (inp[5]) ? 14'b00010000110110 : 14'b00110000110110;
										assign node306 = (inp[2]) ? node316 : node307;
											assign node307 = (inp[4]) ? node311 : node308;
												assign node308 = (inp[7]) ? 14'b00010000010010 : 14'b00000000000001;
												assign node311 = (inp[5]) ? 14'b00010100010110 : node312;
													assign node312 = (inp[7]) ? 14'b00110000010110 : 14'b00110100010110;
											assign node316 = (inp[4]) ? node322 : node317;
												assign node317 = (inp[5]) ? 14'b01010100010010 : node318;
													assign node318 = (inp[7]) ? 14'b01110000010110 : 14'b01110100010110;
												assign node322 = (inp[5]) ? node324 : 14'b00000000000001;
													assign node324 = (inp[11]) ? 14'b00000000000001 : 14'b01010000010010;
									assign node327 = (inp[11]) ? node347 : node328;
										assign node328 = (inp[2]) ? node340 : node329;
											assign node329 = (inp[5]) ? node333 : node330;
												assign node330 = (inp[7]) ? 14'b00010000000010 : 14'b00000000000001;
												assign node333 = (inp[4]) ? node337 : node334;
													assign node334 = (inp[7]) ? 14'b01010000000110 : 14'b01010100100110;
													assign node337 = (inp[7]) ? 14'b00010000000110 : 14'b00010100000110;
											assign node340 = (inp[7]) ? 14'b00000000000001 : node341;
												assign node341 = (inp[4]) ? node343 : 14'b01110100100110;
													assign node343 = (inp[5]) ? 14'b01010000000010 : 14'b00000000000001;
										assign node347 = (inp[9]) ? node359 : node348;
											assign node348 = (inp[4]) ? node356 : node349;
												assign node349 = (inp[2]) ? node353 : node350;
													assign node350 = (inp[5]) ? 14'b01010000100110 : 14'b00000000000000;
													assign node353 = (inp[5]) ? 14'b01010100100010 : 14'b01110000100110;
												assign node356 = (inp[5]) ? 14'b00010100100110 : 14'b00110100100110;
											assign node359 = (inp[2]) ? 14'b00000000000001 : node360;
												assign node360 = (inp[4]) ? 14'b00010100000110 : node361;
													assign node361 = (inp[5]) ? 14'b01010000000110 : 14'b00010000000010;
								assign node366 = (inp[4]) ? node408 : node367;
									assign node367 = (inp[2]) ? node385 : node368;
										assign node368 = (inp[7]) ? node378 : node369;
											assign node369 = (inp[5]) ? 14'b01010100000100 : node370;
												assign node370 = (inp[1]) ? node374 : node371;
													assign node371 = (inp[9]) ? 14'b01010000010100 : 14'b01010000110100;
													assign node374 = (inp[9]) ? 14'b01010000000100 : 14'b01010000100100;
											assign node378 = (inp[5]) ? 14'b00000000000001 : node379;
												assign node379 = (inp[1]) ? 14'b00010000000000 : node380;
													assign node380 = (inp[9]) ? 14'b00010000010000 : 14'b00010000110000;
										assign node385 = (inp[5]) ? node397 : node386;
											assign node386 = (inp[7]) ? node392 : node387;
												assign node387 = (inp[9]) ? 14'b01110100000100 : node388;
													assign node388 = (inp[1]) ? 14'b01110100100100 : 14'b01110100110100;
												assign node392 = (inp[9]) ? 14'b01110000010100 : node393;
													assign node393 = (inp[1]) ? 14'b01110000100100 : 14'b01110000110100;
											assign node397 = (inp[1]) ? node405 : node398;
												assign node398 = (inp[7]) ? node402 : node399;
													assign node399 = (inp[9]) ? 14'b01010100010000 : 14'b01010100110000;
													assign node402 = (inp[9]) ? 14'b01010000010000 : 14'b01010000110000;
												assign node405 = (inp[9]) ? 14'b01010000000000 : 14'b01010000100000;
									assign node408 = (inp[2]) ? node428 : node409;
										assign node409 = (inp[7]) ? node415 : node410;
											assign node410 = (inp[5]) ? 14'b00000000000001 : node411;
												assign node411 = (inp[11]) ? 14'b00110100100100 : 14'b00110100000100;
											assign node415 = (inp[1]) ? node421 : node416;
												assign node416 = (inp[9]) ? 14'b00010000010100 : node417;
													assign node417 = (inp[5]) ? 14'b00010000110100 : 14'b00110000110100;
												assign node421 = (inp[9]) ? node425 : node422;
													assign node422 = (inp[5]) ? 14'b00010000100100 : 14'b00110000100100;
													assign node425 = (inp[5]) ? 14'b00010000000100 : 14'b00110000000100;
										assign node428 = (inp[7]) ? 14'b00000000000001 : node429;
											assign node429 = (inp[5]) ? 14'b00000000000001 : node430;
												assign node430 = (inp[1]) ? node432 : 14'b00010100110100;
													assign node432 = (inp[11]) ? 14'b00010100100100 : 14'b00010100000100;
							assign node437 = (inp[2]) ? node439 : 14'b00000000000001;
								assign node439 = (inp[7]) ? 14'b00000000000001 : node440;
									assign node440 = (inp[12]) ? 14'b00000000000001 : node441;
										assign node441 = (inp[9]) ? 14'b00000000000001 : node442;
											assign node442 = (inp[1]) ? 14'b00000000000001 : node443;
												assign node443 = (inp[5]) ? 14'b00000000000001 : node444;
													assign node444 = (inp[4]) ? 14'b10000001001010 : 14'b00000000000001;
					assign node452 = (inp[5]) ? 14'b00000000000001 : node453;
						assign node453 = (inp[2]) ? node583 : node454;
							assign node454 = (inp[6]) ? node530 : node455;
								assign node455 = (inp[4]) ? node491 : node456;
									assign node456 = (inp[1]) ? node470 : node457;
										assign node457 = (inp[3]) ? node461 : node458;
											assign node458 = (inp[9]) ? 14'b01100100000000 : 14'b00000000000001;
											assign node461 = (inp[12]) ? node465 : node462;
												assign node462 = (inp[7]) ? 14'b01110010010010 : 14'b01110110010010;
												assign node465 = (inp[7]) ? 14'b01110010110000 : node466;
													assign node466 = (inp[9]) ? 14'b01110110010000 : 14'b01110110110000;
										assign node470 = (inp[12]) ? node480 : node471;
											assign node471 = (inp[7]) ? node475 : node472;
												assign node472 = (inp[3]) ? 14'b01100110100010 : 14'b01110110100010;
												assign node475 = (inp[9]) ? node477 : 14'b01110010100010;
													assign node477 = (inp[3]) ? 14'b01100010000010 : 14'b01110010000010;
											assign node480 = (inp[7]) ? node486 : node481;
												assign node481 = (inp[9]) ? node483 : 14'b01100110100000;
													assign node483 = (inp[3]) ? 14'b01100110000000 : 14'b01110110000000;
												assign node486 = (inp[3]) ? 14'b01100010100000 : node487;
													assign node487 = (inp[9]) ? 14'b01110010000000 : 14'b01110010100000;
									assign node491 = (inp[7]) ? node513 : node492;
										assign node492 = (inp[12]) ? node504 : node493;
											assign node493 = (inp[9]) ? node497 : node494;
												assign node494 = (inp[1]) ? 14'b00110110100010 : 14'b00110110110010;
												assign node497 = (inp[1]) ? node501 : node498;
													assign node498 = (inp[3]) ? 14'b00110110010010 : 14'b00100100000010;
													assign node501 = (inp[3]) ? 14'b00100110000010 : 14'b00110110000010;
											assign node504 = (inp[1]) ? node510 : node505;
												assign node505 = (inp[3]) ? 14'b00110110010000 : node506;
													assign node506 = (inp[9]) ? 14'b00100100000000 : 14'b00000000000001;
												assign node510 = (inp[3]) ? 14'b00100110100000 : 14'b00110110100000;
										assign node513 = (inp[1]) ? node519 : node514;
											assign node514 = (inp[3]) ? 14'b00110010110000 : node515;
												assign node515 = (inp[9]) ? 14'b00100000000010 : 14'b00000000000001;
											assign node519 = (inp[9]) ? node525 : node520;
												assign node520 = (inp[3]) ? 14'b00100010100000 : node521;
													assign node521 = (inp[11]) ? 14'b00110010100010 : 14'b00110010100000;
												assign node525 = (inp[3]) ? node527 : 14'b00110010000000;
													assign node527 = (inp[11]) ? 14'b00100010000000 : 14'b00100010000010;
								assign node530 = (inp[3]) ? 14'b00000000000001 : node531;
									assign node531 = (inp[7]) ? node555 : node532;
										assign node532 = (inp[1]) ? node546 : node533;
											assign node533 = (inp[12]) ? node539 : node534;
												assign node534 = (inp[9]) ? node536 : 14'b00110100110010;
													assign node536 = (inp[4]) ? 14'b00110100010010 : 14'b01110100010010;
												assign node539 = (inp[4]) ? node543 : node540;
													assign node540 = (inp[9]) ? 14'b01110100010000 : 14'b01110100110000;
													assign node543 = (inp[9]) ? 14'b00110100010000 : 14'b00110100110000;
											assign node546 = (inp[4]) ? 14'b00110100000000 : node547;
												assign node547 = (inp[9]) ? node551 : node548;
													assign node548 = (inp[12]) ? 14'b01110100100000 : 14'b01110100100010;
													assign node551 = (inp[12]) ? 14'b01110100000000 : 14'b01110100000010;
										assign node555 = (inp[12]) ? node571 : node556;
											assign node556 = (inp[9]) ? node564 : node557;
												assign node557 = (inp[1]) ? node561 : node558;
													assign node558 = (inp[4]) ? 14'b00110000110010 : 14'b01110000110010;
													assign node561 = (inp[4]) ? 14'b00110000100010 : 14'b01110000100010;
												assign node564 = (inp[1]) ? node568 : node565;
													assign node565 = (inp[4]) ? 14'b00110000010010 : 14'b01110000010010;
													assign node568 = (inp[4]) ? 14'b00110000000010 : 14'b01110000000010;
											assign node571 = (inp[1]) ? node579 : node572;
												assign node572 = (inp[4]) ? node576 : node573;
													assign node573 = (inp[9]) ? 14'b01110000010000 : 14'b01110000110000;
													assign node576 = (inp[9]) ? 14'b00110000010000 : 14'b00110000110000;
												assign node579 = (inp[4]) ? 14'b00110000100000 : 14'b01110000100000;
							assign node583 = (inp[7]) ? node629 : node584;
								assign node584 = (inp[4]) ? node592 : node585;
									assign node585 = (inp[9]) ? 14'b00000000000001 : node586;
										assign node586 = (inp[1]) ? 14'b00000000000001 : node587;
											assign node587 = (inp[3]) ? 14'b10000001001000 : 14'b00000000000001;
									assign node592 = (inp[6]) ? node616 : node593;
										assign node593 = (inp[1]) ? node601 : node594;
											assign node594 = (inp[3]) ? node598 : node595;
												assign node595 = (inp[9]) ? 14'b00000100000000 : 14'b00000000000001;
												assign node598 = (inp[12]) ? 14'b00010110110000 : 14'b00010110010010;
											assign node601 = (inp[9]) ? node609 : node602;
												assign node602 = (inp[12]) ? node606 : node603;
													assign node603 = (inp[11]) ? 14'b00000110100010 : 14'b00010110100010;
													assign node606 = (inp[3]) ? 14'b00000110100000 : 14'b00010110100000;
												assign node609 = (inp[12]) ? node613 : node610;
													assign node610 = (inp[3]) ? 14'b00000110000010 : 14'b00010110000010;
													assign node613 = (inp[3]) ? 14'b00000110000000 : 14'b00010110000000;
										assign node616 = (inp[3]) ? 14'b00000000000001 : node617;
											assign node617 = (inp[9]) ? node623 : node618;
												assign node618 = (inp[1]) ? 14'b00010100100000 : node619;
													assign node619 = (inp[12]) ? 14'b00010100110000 : 14'b00010100110010;
												assign node623 = (inp[12]) ? node625 : 14'b00010100000010;
													assign node625 = (inp[1]) ? 14'b00010100000000 : 14'b00010100010000;
								assign node629 = (inp[1]) ? node631 : 14'b00000000000001;
									assign node631 = (inp[4]) ? node633 : 14'b00000000000001;
										assign node633 = (inp[6]) ? node635 : 14'b00000000000001;
											assign node635 = (inp[3]) ? 14'b10000000000000 : 14'b00000000000001;
				assign node639 = (inp[1]) ? node915 : node640;
					assign node640 = (inp[3]) ? node850 : node641;
						assign node641 = (inp[10]) ? node787 : node642;
							assign node642 = (inp[4]) ? node728 : node643;
								assign node643 = (inp[7]) ? node693 : node644;
									assign node644 = (inp[5]) ? node666 : node645;
										assign node645 = (inp[2]) ? node655 : node646;
											assign node646 = (inp[12]) ? node648 : 14'b00000000000001;
												assign node648 = (inp[6]) ? node652 : node649;
													assign node649 = (inp[9]) ? 14'b01000010010100 : 14'b01000010110100;
													assign node652 = (inp[11]) ? 14'b01000000010100 : 14'b01000000110100;
											assign node655 = (inp[12]) ? node661 : node656;
												assign node656 = (inp[6]) ? node658 : 14'b01100110010110;
													assign node658 = (inp[9]) ? 14'b01100100010110 : 14'b01100100110110;
												assign node661 = (inp[9]) ? 14'b01100100010100 : node662;
													assign node662 = (inp[6]) ? 14'b01100100110100 : 14'b01100110110100;
										assign node666 = (inp[12]) ? node680 : node667;
											assign node667 = (inp[6]) ? node675 : node668;
												assign node668 = (inp[2]) ? node672 : node669;
													assign node669 = (inp[9]) ? 14'b01000110010110 : 14'b01000110110110;
													assign node672 = (inp[9]) ? 14'b01000110010010 : 14'b01000110110010;
												assign node675 = (inp[9]) ? 14'b01000100010010 : node676;
													assign node676 = (inp[2]) ? 14'b01000100110010 : 14'b01000100110110;
											assign node680 = (inp[9]) ? node686 : node681;
												assign node681 = (inp[2]) ? 14'b01000110110000 : node682;
													assign node682 = (inp[6]) ? 14'b01000100110100 : 14'b01000110110100;
												assign node686 = (inp[2]) ? node690 : node687;
													assign node687 = (inp[6]) ? 14'b01000100010100 : 14'b01000110010100;
													assign node690 = (inp[6]) ? 14'b01000100010000 : 14'b01000110010000;
									assign node693 = (inp[2]) ? node715 : node694;
										assign node694 = (inp[12]) ? node708 : node695;
											assign node695 = (inp[5]) ? node701 : node696;
												assign node696 = (inp[6]) ? 14'b00000000110010 : node697;
													assign node697 = (inp[9]) ? 14'b00000010010010 : 14'b00000010110010;
												assign node701 = (inp[9]) ? node705 : node702;
													assign node702 = (inp[6]) ? 14'b01000000110110 : 14'b01000010110110;
													assign node705 = (inp[6]) ? 14'b01000000010110 : 14'b01000010010110;
											assign node708 = (inp[5]) ? 14'b00000000000001 : node709;
												assign node709 = (inp[9]) ? node711 : 14'b00000010110000;
													assign node711 = (inp[6]) ? 14'b00000000010000 : 14'b00000010010000;
										assign node715 = (inp[5]) ? 14'b00000000000001 : node716;
											assign node716 = (inp[12]) ? node720 : node717;
												assign node717 = (inp[6]) ? 14'b01100000010110 : 14'b01100010010110;
												assign node720 = (inp[6]) ? node724 : node721;
													assign node721 = (inp[9]) ? 14'b01100010010100 : 14'b01100010110100;
													assign node724 = (inp[9]) ? 14'b01100000010100 : 14'b01100000110100;
								assign node728 = (inp[2]) ? node768 : node729;
									assign node729 = (inp[5]) ? node751 : node730;
										assign node730 = (inp[6]) ? node742 : node731;
											assign node731 = (inp[7]) ? node739 : node732;
												assign node732 = (inp[9]) ? node736 : node733;
													assign node733 = (inp[11]) ? 14'b00100110110100 : 14'b00100110110110;
													assign node736 = (inp[12]) ? 14'b00100110010100 : 14'b00100110010110;
												assign node739 = (inp[9]) ? 14'b00100010010100 : 14'b00100010110100;
											assign node742 = (inp[12]) ? node748 : node743;
												assign node743 = (inp[9]) ? 14'b00100000010110 : node744;
													assign node744 = (inp[7]) ? 14'b00100000110110 : 14'b00100100110110;
												assign node748 = (inp[7]) ? 14'b00100000110100 : 14'b00100100110100;
										assign node751 = (inp[7]) ? node755 : node752;
											assign node752 = (inp[12]) ? 14'b00000000000001 : 14'b00000100010110;
											assign node755 = (inp[9]) ? node763 : node756;
												assign node756 = (inp[12]) ? node760 : node757;
													assign node757 = (inp[6]) ? 14'b00000000110110 : 14'b00000010110110;
													assign node760 = (inp[6]) ? 14'b00000000110100 : 14'b00000010110100;
												assign node763 = (inp[12]) ? node765 : 14'b00000000010110;
													assign node765 = (inp[6]) ? 14'b00000000010100 : 14'b00000010010100;
									assign node768 = (inp[7]) ? 14'b00000000000001 : node769;
										assign node769 = (inp[12]) ? node779 : node770;
											assign node770 = (inp[5]) ? node772 : 14'b00000000000001;
												assign node772 = (inp[6]) ? node776 : node773;
													assign node773 = (inp[9]) ? 14'b01000010010010 : 14'b01000010110010;
													assign node776 = (inp[9]) ? 14'b01000000010010 : 14'b01000000110010;
											assign node779 = (inp[5]) ? 14'b00000000000001 : node780;
												assign node780 = (inp[9]) ? node782 : 14'b00000110110100;
													assign node782 = (inp[6]) ? 14'b00000100010100 : 14'b00000110010100;
							assign node787 = (inp[5]) ? 14'b00000000000001 : node788;
								assign node788 = (inp[2]) ? node838 : node789;
									assign node789 = (inp[6]) ? node815 : node790;
										assign node790 = (inp[12]) ? node802 : node791;
											assign node791 = (inp[9]) ? node799 : node792;
												assign node792 = (inp[4]) ? node796 : node793;
													assign node793 = (inp[7]) ? 14'b01100010110010 : 14'b01100110110010;
													assign node796 = (inp[7]) ? 14'b00100010110010 : 14'b00100110110010;
												assign node799 = (inp[7]) ? 14'b01100010010010 : 14'b01100110010010;
											assign node802 = (inp[4]) ? node808 : node803;
												assign node803 = (inp[7]) ? node805 : 14'b01100110110000;
													assign node805 = (inp[9]) ? 14'b01100010010000 : 14'b01100010110000;
												assign node808 = (inp[9]) ? node812 : node809;
													assign node809 = (inp[7]) ? 14'b00100010110000 : 14'b00100110110000;
													assign node812 = (inp[11]) ? 14'b00100110010000 : 14'b00100010010000;
										assign node815 = (inp[12]) ? node823 : node816;
											assign node816 = (inp[9]) ? node820 : node817;
												assign node817 = (inp[4]) ? 14'b00100000110010 : 14'b01100000110010;
												assign node820 = (inp[4]) ? 14'b00100000010010 : 14'b01100000010010;
											assign node823 = (inp[7]) ? node831 : node824;
												assign node824 = (inp[9]) ? node828 : node825;
													assign node825 = (inp[11]) ? 14'b00100100110000 : 14'b01100100110000;
													assign node828 = (inp[4]) ? 14'b00100100010000 : 14'b01100100010000;
												assign node831 = (inp[9]) ? node835 : node832;
													assign node832 = (inp[4]) ? 14'b00100000110000 : 14'b01100000110000;
													assign node835 = (inp[4]) ? 14'b00100000010000 : 14'b01100000010000;
									assign node838 = (inp[4]) ? node840 : 14'b00000000000001;
										assign node840 = (inp[7]) ? 14'b00000000000001 : node841;
											assign node841 = (inp[12]) ? 14'b00000100110000 : node842;
												assign node842 = (inp[9]) ? 14'b00000100010010 : node843;
													assign node843 = (inp[6]) ? 14'b00000100110010 : 14'b00000110110010;
						assign node850 = (inp[9]) ? 14'b00000000000001 : node851;
							assign node851 = (inp[6]) ? node853 : 14'b00000000000001;
								assign node853 = (inp[2]) ? node891 : node854;
									assign node854 = (inp[5]) ? node880 : node855;
										assign node855 = (inp[4]) ? node869 : node856;
											assign node856 = (inp[10]) ? node864 : node857;
												assign node857 = (inp[7]) ? node861 : node858;
													assign node858 = (inp[12]) ? 14'b01000000100100 : 14'b00000000000001;
													assign node861 = (inp[12]) ? 14'b00000000100000 : 14'b00000000100010;
												assign node864 = (inp[7]) ? node866 : 14'b01100100100000;
													assign node866 = (inp[12]) ? 14'b01100000100000 : 14'b01100000100010;
											assign node869 = (inp[10]) ? node873 : node870;
												assign node870 = (inp[12]) ? 14'b00100100100100 : 14'b00100100100110;
												assign node873 = (inp[12]) ? node877 : node874;
													assign node874 = (inp[7]) ? 14'b00100000100010 : 14'b00100100100010;
													assign node877 = (inp[7]) ? 14'b00100000100000 : 14'b00100100100000;
										assign node880 = (inp[10]) ? 14'b00000000000001 : node881;
											assign node881 = (inp[12]) ? node887 : node882;
												assign node882 = (inp[7]) ? node884 : 14'b00000100100110;
													assign node884 = (inp[4]) ? 14'b00000000100110 : 14'b01000000100110;
												assign node887 = (inp[7]) ? 14'b00000000100100 : 14'b00000000000001;
									assign node891 = (inp[7]) ? node907 : node892;
										assign node892 = (inp[10]) ? node902 : node893;
											assign node893 = (inp[4]) ? node899 : node894;
												assign node894 = (inp[5]) ? node896 : 14'b01100100100100;
													assign node896 = (inp[12]) ? 14'b01000100100000 : 14'b01000100100010;
												assign node899 = (inp[12]) ? 14'b00000000000001 : 14'b01000000100010;
											assign node902 = (inp[4]) ? node904 : 14'b00000000000001;
												assign node904 = (inp[12]) ? 14'b00000100100000 : 14'b00000100100010;
										assign node907 = (inp[4]) ? 14'b00000000000001 : node908;
											assign node908 = (inp[10]) ? 14'b00000000000001 : node909;
												assign node909 = (inp[5]) ? 14'b00000000000001 : 14'b01100000100100;
					assign node915 = (inp[7]) ? 14'b00000000000001 : node916;
						assign node916 = (inp[11]) ? 14'b00000000000001 : node917;
							assign node917 = (inp[12]) ? 14'b00000000000001 : node918;
								assign node918 = (inp[6]) ? 14'b00000000000001 : node919;
									assign node919 = (inp[5]) ? 14'b00000000000001 : node920;
										assign node920 = (inp[10]) ? 14'b00000000000001 : node921;
											assign node921 = (inp[3]) ? node925 : node922;
												assign node922 = (inp[2]) ? 14'b10000001000010 : 14'b00000000000001;
												assign node925 = (inp[2]) ? 14'b00000000000001 : node926;
													assign node926 = (inp[4]) ? 14'b00000000000001 : 14'b10000000000010;
		assign node936 = (inp[0]) ? node2144 : node937;
			assign node937 = (inp[3]) ? node1669 : node938;
				assign node938 = (inp[2]) ? node1362 : node939;
					assign node939 = (inp[13]) ? node1195 : node940;
						assign node940 = (inp[10]) ? node1118 : node941;
							assign node941 = (inp[7]) ? node1029 : node942;
								assign node942 = (inp[6]) ? node982 : node943;
									assign node943 = (inp[9]) ? node957 : node944;
										assign node944 = (inp[1]) ? node946 : 14'b00000000000001;
											assign node946 = (inp[4]) ? node952 : node947;
												assign node947 = (inp[12]) ? node949 : 14'b00110010000010;
													assign node949 = (inp[11]) ? 14'b01010010000100 : 14'b01010010000110;
												assign node952 = (inp[11]) ? 14'b00000000000001 : node953;
													assign node953 = (inp[12]) ? 14'b00000000000000 : 14'b01111010000110;
										assign node957 = (inp[4]) ? node969 : node958;
											assign node958 = (inp[1]) ? node964 : node959;
												assign node959 = (inp[12]) ? node961 : 14'b01101100000100;
													assign node961 = (inp[5]) ? 14'b01000100000100 : 14'b01001100000100;
												assign node964 = (inp[12]) ? node966 : 14'b00000000000001;
													assign node966 = (inp[5]) ? 14'b01000000000110 : 14'b01001000000100;
											assign node969 = (inp[11]) ? node977 : node970;
												assign node970 = (inp[12]) ? node974 : node971;
													assign node971 = (inp[1]) ? 14'b01100000000110 : 14'b01100100000110;
													assign node974 = (inp[5]) ? 14'b01000100000010 : 14'b00000000000001;
												assign node977 = (inp[12]) ? node979 : 14'b00000000000001;
													assign node979 = (inp[1]) ? 14'b01000000000000 : 14'b01000100000000;
									assign node982 = (inp[5]) ? node1002 : node983;
										assign node983 = (inp[11]) ? node993 : node984;
											assign node984 = (inp[1]) ? node988 : node985;
												assign node985 = (inp[12]) ? 14'b00000000000001 : 14'b01111100010110;
												assign node988 = (inp[12]) ? node990 : 14'b00000000000001;
													assign node990 = (inp[4]) ? 14'b00000000000001 : 14'b01011000010110;
											assign node993 = (inp[1]) ? node997 : node994;
												assign node994 = (inp[12]) ? 14'b01011100110000 : 14'b00000000000001;
												assign node997 = (inp[9]) ? node999 : 14'b01111000110100;
													assign node999 = (inp[12]) ? 14'b01011000010100 : 14'b01111000010100;
										assign node1002 = (inp[1]) ? node1016 : node1003;
											assign node1003 = (inp[9]) ? node1009 : node1004;
												assign node1004 = (inp[12]) ? node1006 : 14'b01110100110110;
													assign node1006 = (inp[11]) ? 14'b01010100110100 : 14'b01010100110010;
												assign node1009 = (inp[12]) ? node1013 : node1010;
													assign node1010 = (inp[11]) ? 14'b01110100010100 : 14'b00110100010010;
													assign node1013 = (inp[4]) ? 14'b01010100010000 : 14'b01010100010110;
											assign node1016 = (inp[11]) ? node1024 : node1017;
												assign node1017 = (inp[12]) ? node1021 : node1018;
													assign node1018 = (inp[4]) ? 14'b01110000010110 : 14'b00110000010010;
													assign node1021 = (inp[4]) ? 14'b01010000010010 : 14'b01010000010110;
												assign node1024 = (inp[12]) ? node1026 : 14'b00000000000001;
													assign node1026 = (inp[4]) ? 14'b01010000110000 : 14'b01010000010100;
								assign node1029 = (inp[12]) ? node1067 : node1030;
									assign node1030 = (inp[11]) ? node1052 : node1031;
										assign node1031 = (inp[4]) ? node1041 : node1032;
											assign node1032 = (inp[5]) ? node1034 : 14'b00000000000001;
												assign node1034 = (inp[9]) ? node1038 : node1035;
													assign node1035 = (inp[1]) ? 14'b00100000110010 : 14'b00100110110010;
													assign node1038 = (inp[6]) ? 14'b00100100010010 : 14'b00100010010010;
											assign node1041 = (inp[1]) ? node1049 : node1042;
												assign node1042 = (inp[6]) ? node1046 : node1043;
													assign node1043 = (inp[9]) ? 14'b01101110010110 : 14'b01101110110110;
													assign node1046 = (inp[9]) ? 14'b01101100010110 : 14'b01101100110110;
												assign node1049 = (inp[9]) ? 14'b01101010010110 : 14'b01101010110110;
										assign node1052 = (inp[4]) ? 14'b00000000000001 : node1053;
											assign node1053 = (inp[1]) ? node1059 : node1054;
												assign node1054 = (inp[9]) ? node1056 : 14'b01101100110100;
													assign node1056 = (inp[5]) ? 14'b01100100010100 : 14'b01101100010100;
												assign node1059 = (inp[6]) ? node1063 : node1060;
													assign node1060 = (inp[9]) ? 14'b01100010010100 : 14'b01100010110100;
													assign node1063 = (inp[9]) ? 14'b01101000010100 : 14'b01100000110100;
									assign node1067 = (inp[4]) ? node1095 : node1068;
										assign node1068 = (inp[6]) ? node1084 : node1069;
											assign node1069 = (inp[11]) ? node1077 : node1070;
												assign node1070 = (inp[5]) ? node1074 : node1071;
													assign node1071 = (inp[9]) ? 14'b01001010010110 : 14'b01001010110110;
													assign node1074 = (inp[9]) ? 14'b01000010010110 : 14'b01000010110110;
												assign node1077 = (inp[9]) ? node1081 : node1078;
													assign node1078 = (inp[1]) ? 14'b01000010110100 : 14'b01001110110100;
													assign node1081 = (inp[1]) ? 14'b01001010010100 : 14'b01001110010100;
											assign node1084 = (inp[9]) ? node1090 : node1085;
												assign node1085 = (inp[5]) ? 14'b01000100110110 : node1086;
													assign node1086 = (inp[11]) ? 14'b01001000110100 : 14'b01001000110110;
												assign node1090 = (inp[5]) ? node1092 : 14'b01001100010110;
													assign node1092 = (inp[1]) ? 14'b01000000010100 : 14'b01000100010100;
										assign node1095 = (inp[11]) ? node1105 : node1096;
											assign node1096 = (inp[5]) ? node1098 : 14'b00000000000001;
												assign node1098 = (inp[1]) ? node1102 : node1099;
													assign node1099 = (inp[6]) ? 14'b01000100010010 : 14'b01000110110010;
													assign node1102 = (inp[9]) ? 14'b01000010010010 : 14'b01000000110010;
											assign node1105 = (inp[1]) ? node1113 : node1106;
												assign node1106 = (inp[5]) ? node1110 : node1107;
													assign node1107 = (inp[6]) ? 14'b01001100110000 : 14'b01001110010000;
													assign node1110 = (inp[9]) ? 14'b01000110010000 : 14'b01000110110000;
												assign node1113 = (inp[6]) ? 14'b01000000110000 : node1114;
													assign node1114 = (inp[5]) ? 14'b01000010110000 : 14'b01001010110000;
							assign node1118 = (inp[11]) ? 14'b00000000000001 : node1119;
								assign node1119 = (inp[12]) ? node1167 : node1120;
									assign node1120 = (inp[6]) ? node1140 : node1121;
										assign node1121 = (inp[7]) ? node1133 : node1122;
											assign node1122 = (inp[1]) ? node1126 : node1123;
												assign node1123 = (inp[9]) ? 14'b01100100000000 : 14'b00000000000001;
												assign node1126 = (inp[9]) ? node1130 : node1127;
													assign node1127 = (inp[5]) ? 14'b01110010000000 : 14'b01111010000000;
													assign node1130 = (inp[4]) ? 14'b01100000000000 : 14'b01100000000010;
											assign node1133 = (inp[9]) ? node1137 : node1134;
												assign node1134 = (inp[1]) ? 14'b01100010110000 : 14'b01100110110010;
												assign node1137 = (inp[5]) ? 14'b01100110010000 : 14'b01101110010000;
										assign node1140 = (inp[1]) ? node1152 : node1141;
											assign node1141 = (inp[4]) ? node1145 : node1142;
												assign node1142 = (inp[5]) ? 14'b01100100010010 : 14'b01101100010010;
												assign node1145 = (inp[9]) ? node1149 : node1146;
													assign node1146 = (inp[5]) ? 14'b01110100110000 : 14'b01101100110000;
													assign node1149 = (inp[7]) ? 14'b01101100010000 : 14'b01111100010000;
											assign node1152 = (inp[9]) ? node1160 : node1153;
												assign node1153 = (inp[7]) ? node1157 : node1154;
													assign node1154 = (inp[5]) ? 14'b01110000110000 : 14'b01111000110010;
													assign node1157 = (inp[5]) ? 14'b01100000110000 : 14'b01101000110000;
												assign node1160 = (inp[7]) ? node1164 : node1161;
													assign node1161 = (inp[4]) ? 14'b01110000010000 : 14'b01110000010010;
													assign node1164 = (inp[4]) ? 14'b01100000010000 : 14'b01100000010010;
									assign node1167 = (inp[5]) ? 14'b00000000000001 : node1168;
										assign node1168 = (inp[4]) ? node1180 : node1169;
											assign node1169 = (inp[6]) ? node1175 : node1170;
												assign node1170 = (inp[9]) ? node1172 : 14'b00000000000001;
													assign node1172 = (inp[7]) ? 14'b01001110010010 : 14'b01001100000010;
												assign node1175 = (inp[7]) ? 14'b01001000110010 : node1176;
													assign node1176 = (inp[9]) ? 14'b01011000010010 : 14'b01011000110010;
											assign node1180 = (inp[7]) ? node1186 : node1181;
												assign node1181 = (inp[1]) ? node1183 : 14'b00000000000001;
													assign node1183 = (inp[9]) ? 14'b00101000000000 : 14'b00111010000000;
												assign node1186 = (inp[9]) ? node1190 : node1187;
													assign node1187 = (inp[6]) ? 14'b00101000110000 : 14'b00101110110000;
													assign node1190 = (inp[6]) ? 14'b00101100010000 : 14'b00101010010000;
						assign node1195 = (inp[12]) ? node1307 : node1196;
							assign node1196 = (inp[4]) ? node1248 : node1197;
								assign node1197 = (inp[5]) ? node1221 : node1198;
									assign node1198 = (inp[7]) ? node1206 : node1199;
										assign node1199 = (inp[9]) ? 14'b00000000000001 : node1200;
											assign node1200 = (inp[11]) ? node1202 : 14'b00000000000001;
												assign node1202 = (inp[1]) ? 14'b00000000000001 : 14'b10000000001000;
										assign node1206 = (inp[1]) ? node1214 : node1207;
											assign node1207 = (inp[6]) ? node1211 : node1208;
												assign node1208 = (inp[9]) ? 14'b00000000000000 : 14'b00000000000001;
												assign node1211 = (inp[9]) ? 14'b00010000010000 : 14'b00010000110000;
											assign node1214 = (inp[6]) ? node1218 : node1215;
												assign node1215 = (inp[9]) ? 14'b00010010000000 : 14'b00010010100000;
												assign node1218 = (inp[9]) ? 14'b00010000000000 : 14'b00010000100000;
									assign node1221 = (inp[6]) ? node1233 : node1222;
										assign node1222 = (inp[1]) ? node1228 : node1223;
											assign node1223 = (inp[9]) ? node1225 : 14'b00000000000001;
												assign node1225 = (inp[7]) ? 14'b01100000000000 : 14'b01100100000000;
											assign node1228 = (inp[7]) ? 14'b01110010100000 : node1229;
												assign node1229 = (inp[9]) ? 14'b01110110000000 : 14'b01110110100000;
										assign node1233 = (inp[1]) ? node1241 : node1234;
											assign node1234 = (inp[7]) ? node1238 : node1235;
												assign node1235 = (inp[9]) ? 14'b01110100010000 : 14'b01110100110000;
												assign node1238 = (inp[9]) ? 14'b01110000010000 : 14'b01110000110000;
											assign node1241 = (inp[7]) ? node1245 : node1242;
												assign node1242 = (inp[9]) ? 14'b01110100000000 : 14'b01110100100000;
												assign node1245 = (inp[9]) ? 14'b01110000000000 : 14'b01110000100000;
								assign node1248 = (inp[5]) ? node1278 : node1249;
									assign node1249 = (inp[7]) ? node1263 : node1250;
										assign node1250 = (inp[9]) ? node1256 : node1251;
											assign node1251 = (inp[6]) ? node1253 : 14'b00110110100100;
												assign node1253 = (inp[1]) ? 14'b00110100100100 : 14'b00110100110100;
											assign node1256 = (inp[6]) ? node1260 : node1257;
												assign node1257 = (inp[1]) ? 14'b00110110000100 : 14'b00100100000100;
												assign node1260 = (inp[1]) ? 14'b00110100000100 : 14'b00110100010100;
										assign node1263 = (inp[1]) ? node1271 : node1264;
											assign node1264 = (inp[6]) ? node1268 : node1265;
												assign node1265 = (inp[9]) ? 14'b00100000000100 : 14'b00000000000001;
												assign node1268 = (inp[9]) ? 14'b00110000010100 : 14'b00110000110100;
											assign node1271 = (inp[9]) ? node1275 : node1272;
												assign node1272 = (inp[6]) ? 14'b00110000100100 : 14'b00110010100100;
												assign node1275 = (inp[6]) ? 14'b00110000000100 : 14'b00110010000100;
									assign node1278 = (inp[1]) ? node1292 : node1279;
										assign node1279 = (inp[6]) ? node1285 : node1280;
											assign node1280 = (inp[9]) ? node1282 : 14'b00000000000001;
												assign node1282 = (inp[7]) ? 14'b00100000000000 : 14'b00100100000000;
											assign node1285 = (inp[7]) ? node1289 : node1286;
												assign node1286 = (inp[9]) ? 14'b00110100010000 : 14'b00110100110000;
												assign node1289 = (inp[9]) ? 14'b00110000010000 : 14'b00110000110000;
										assign node1292 = (inp[9]) ? node1300 : node1293;
											assign node1293 = (inp[7]) ? node1297 : node1294;
												assign node1294 = (inp[6]) ? 14'b00110100100000 : 14'b00110110100000;
												assign node1297 = (inp[6]) ? 14'b00110000100000 : 14'b00110010100000;
											assign node1300 = (inp[6]) ? node1304 : node1301;
												assign node1301 = (inp[7]) ? 14'b00110010000000 : 14'b00110110000000;
												assign node1304 = (inp[7]) ? 14'b00110000000000 : 14'b00110100000000;
							assign node1307 = (inp[5]) ? 14'b00000000000001 : node1308;
								assign node1308 = (inp[1]) ? node1330 : node1309;
									assign node1309 = (inp[6]) ? node1319 : node1310;
										assign node1310 = (inp[9]) ? node1312 : 14'b00000000000001;
											assign node1312 = (inp[4]) ? node1316 : node1313;
												assign node1313 = (inp[7]) ? 14'b01000000000100 : 14'b01000100000100;
												assign node1316 = (inp[11]) ? 14'b00000100000100 : 14'b00000000000100;
										assign node1319 = (inp[7]) ? node1325 : node1320;
											assign node1320 = (inp[9]) ? 14'b00010100010100 : node1321;
												assign node1321 = (inp[4]) ? 14'b00010100110100 : 14'b01010100110100;
											assign node1325 = (inp[9]) ? 14'b01010000010100 : node1326;
												assign node1326 = (inp[4]) ? 14'b00010000110100 : 14'b01010000110100;
									assign node1330 = (inp[4]) ? node1346 : node1331;
										assign node1331 = (inp[9]) ? node1339 : node1332;
											assign node1332 = (inp[6]) ? node1336 : node1333;
												assign node1333 = (inp[7]) ? 14'b01010010100100 : 14'b01010110100100;
												assign node1336 = (inp[7]) ? 14'b01010000100100 : 14'b01010100100100;
											assign node1339 = (inp[6]) ? node1343 : node1340;
												assign node1340 = (inp[7]) ? 14'b01010010000100 : 14'b01010110000100;
												assign node1343 = (inp[7]) ? 14'b01010000000100 : 14'b01010100000100;
										assign node1346 = (inp[7]) ? node1354 : node1347;
											assign node1347 = (inp[6]) ? node1351 : node1348;
												assign node1348 = (inp[9]) ? 14'b00010110000100 : 14'b00010110100100;
												assign node1351 = (inp[9]) ? 14'b00010100000100 : 14'b00010100100100;
											assign node1354 = (inp[9]) ? node1358 : node1355;
												assign node1355 = (inp[6]) ? 14'b00010000100100 : 14'b00010010100100;
												assign node1358 = (inp[6]) ? 14'b00010000000100 : 14'b00010010000100;
					assign node1362 = (inp[4]) ? node1588 : node1363;
						assign node1363 = (inp[5]) ? node1501 : node1364;
							assign node1364 = (inp[13]) ? node1442 : node1365;
								assign node1365 = (inp[11]) ? node1415 : node1366;
									assign node1366 = (inp[6]) ? node1388 : node1367;
										assign node1367 = (inp[7]) ? node1377 : node1368;
											assign node1368 = (inp[9]) ? node1372 : node1369;
												assign node1369 = (inp[1]) ? 14'b00011010000000 : 14'b00000000000001;
												assign node1372 = (inp[1]) ? node1374 : 14'b00001100000110;
													assign node1374 = (inp[12]) ? 14'b00001000000010 : 14'b00001000000000;
											assign node1377 = (inp[12]) ? node1381 : node1378;
												assign node1378 = (inp[10]) ? 14'b00101010110010 : 14'b00001010110000;
												assign node1381 = (inp[9]) ? node1385 : node1382;
													assign node1382 = (inp[1]) ? 14'b00001010110110 : 14'b00001110110110;
													assign node1385 = (inp[10]) ? 14'b00001010010010 : 14'b00001010010110;
										assign node1388 = (inp[10]) ? node1402 : node1389;
											assign node1389 = (inp[12]) ? node1395 : node1390;
												assign node1390 = (inp[1]) ? node1392 : 14'b00001100010000;
													assign node1392 = (inp[7]) ? 14'b00001000110000 : 14'b00011000110000;
												assign node1395 = (inp[7]) ? node1399 : node1396;
													assign node1396 = (inp[1]) ? 14'b00011000110110 : 14'b00011100110110;
													assign node1399 = (inp[9]) ? 14'b00001000010110 : 14'b00001000110110;
											assign node1402 = (inp[7]) ? node1410 : node1403;
												assign node1403 = (inp[1]) ? node1407 : node1404;
													assign node1404 = (inp[9]) ? 14'b00011100010010 : 14'b00011100110010;
													assign node1407 = (inp[12]) ? 14'b00011000110010 : 14'b00111000010010;
												assign node1410 = (inp[9]) ? node1412 : 14'b00101100110010;
													assign node1412 = (inp[1]) ? 14'b00101000010010 : 14'b00101100010010;
									assign node1415 = (inp[10]) ? 14'b00000000000001 : node1416;
										assign node1416 = (inp[7]) ? node1430 : node1417;
											assign node1417 = (inp[6]) ? node1425 : node1418;
												assign node1418 = (inp[1]) ? node1422 : node1419;
													assign node1419 = (inp[9]) ? 14'b00101100000100 : 14'b00000000000001;
													assign node1422 = (inp[9]) ? 14'b00001000000100 : 14'b00111010000100;
												assign node1425 = (inp[9]) ? node1427 : 14'b00111000110100;
													assign node1427 = (inp[1]) ? 14'b00011000010100 : 14'b00111100010100;
											assign node1430 = (inp[9]) ? node1436 : node1431;
												assign node1431 = (inp[6]) ? node1433 : 14'b00001110110100;
													assign node1433 = (inp[1]) ? 14'b00001000110100 : 14'b00001100110100;
												assign node1436 = (inp[6]) ? node1438 : 14'b00101110010100;
													assign node1438 = (inp[12]) ? 14'b00001100010100 : 14'b00101100010100;
								assign node1442 = (inp[12]) ? node1472 : node1443;
									assign node1443 = (inp[6]) ? node1457 : node1444;
										assign node1444 = (inp[1]) ? node1450 : node1445;
											assign node1445 = (inp[9]) ? node1447 : 14'b00000000000001;
												assign node1447 = (inp[7]) ? 14'b01100000000100 : 14'b01100100000100;
											assign node1450 = (inp[9]) ? node1454 : node1451;
												assign node1451 = (inp[7]) ? 14'b01110010100100 : 14'b01110110100100;
												assign node1454 = (inp[7]) ? 14'b01110010000100 : 14'b01110110000100;
										assign node1457 = (inp[1]) ? node1465 : node1458;
											assign node1458 = (inp[9]) ? node1462 : node1459;
												assign node1459 = (inp[7]) ? 14'b01110000110100 : 14'b01110100110100;
												assign node1462 = (inp[7]) ? 14'b01110000010100 : 14'b01110100010100;
											assign node1465 = (inp[7]) ? node1469 : node1466;
												assign node1466 = (inp[9]) ? 14'b01110100000100 : 14'b01110100100100;
												assign node1469 = (inp[9]) ? 14'b01110000000100 : 14'b01110000100100;
									assign node1472 = (inp[7]) ? node1486 : node1473;
										assign node1473 = (inp[6]) ? node1481 : node1474;
											assign node1474 = (inp[1]) ? node1478 : node1475;
												assign node1475 = (inp[9]) ? 14'b01000100000000 : 14'b00000000000001;
												assign node1478 = (inp[9]) ? 14'b01010110000000 : 14'b01010110100000;
											assign node1481 = (inp[9]) ? node1483 : 14'b01010100110000;
												assign node1483 = (inp[1]) ? 14'b01010100000000 : 14'b01010100010000;
										assign node1486 = (inp[1]) ? node1494 : node1487;
											assign node1487 = (inp[6]) ? node1491 : node1488;
												assign node1488 = (inp[9]) ? 14'b01000000000000 : 14'b00000000000001;
												assign node1491 = (inp[11]) ? 14'b01010000010000 : 14'b01010000110000;
											assign node1494 = (inp[9]) ? node1498 : node1495;
												assign node1495 = (inp[6]) ? 14'b01010000100000 : 14'b01010010100000;
												assign node1498 = (inp[6]) ? 14'b01010000000000 : 14'b01010010000000;
							assign node1501 = (inp[13]) ? node1577 : node1502;
								assign node1502 = (inp[10]) ? node1560 : node1503;
									assign node1503 = (inp[1]) ? node1531 : node1504;
										assign node1504 = (inp[6]) ? node1516 : node1505;
											assign node1505 = (inp[7]) ? node1511 : node1506;
												assign node1506 = (inp[9]) ? node1508 : 14'b00000000000001;
													assign node1508 = (inp[12]) ? 14'b00000100000100 : 14'b00000100000000;
												assign node1511 = (inp[9]) ? 14'b00000110010100 : node1512;
													assign node1512 = (inp[11]) ? 14'b00000110110100 : 14'b00000110110110;
											assign node1516 = (inp[9]) ? node1524 : node1517;
												assign node1517 = (inp[12]) ? node1521 : node1518;
													assign node1518 = (inp[7]) ? 14'b00000100110000 : 14'b00010100110000;
													assign node1521 = (inp[7]) ? 14'b00000100110110 : 14'b00010100110110;
												assign node1524 = (inp[7]) ? node1528 : node1525;
													assign node1525 = (inp[12]) ? 14'b00010100010100 : 14'b00110100010100;
													assign node1528 = (inp[12]) ? 14'b00000100010100 : 14'b00000100010000;
										assign node1531 = (inp[7]) ? node1545 : node1532;
											assign node1532 = (inp[6]) ? node1538 : node1533;
												assign node1533 = (inp[9]) ? 14'b00000000000100 : node1534;
													assign node1534 = (inp[11]) ? 14'b00010010000100 : 14'b00010010000110;
												assign node1538 = (inp[9]) ? node1542 : node1539;
													assign node1539 = (inp[11]) ? 14'b00010000110100 : 14'b00010000110000;
													assign node1542 = (inp[11]) ? 14'b00010000010100 : 14'b00010000010110;
											assign node1545 = (inp[11]) ? node1553 : node1546;
												assign node1546 = (inp[12]) ? node1550 : node1547;
													assign node1547 = (inp[6]) ? 14'b00000000110000 : 14'b00000010010000;
													assign node1550 = (inp[9]) ? 14'b00000010010110 : 14'b00000010110110;
												assign node1553 = (inp[9]) ? node1557 : node1554;
													assign node1554 = (inp[6]) ? 14'b00100000110100 : 14'b00000010110100;
													assign node1557 = (inp[6]) ? 14'b00100000010100 : 14'b00100010010100;
									assign node1560 = (inp[11]) ? 14'b00000000000001 : node1561;
										assign node1561 = (inp[12]) ? node1563 : 14'b00000000000001;
											assign node1563 = (inp[1]) ? node1571 : node1564;
												assign node1564 = (inp[6]) ? node1568 : node1565;
													assign node1565 = (inp[9]) ? 14'b00000100000010 : 14'b00000000000001;
													assign node1568 = (inp[9]) ? 14'b00000100010010 : 14'b00000100110010;
												assign node1571 = (inp[9]) ? 14'b00000000010010 : node1572;
													assign node1572 = (inp[7]) ? 14'b00000000110010 : 14'b00010000110010;
								assign node1577 = (inp[12]) ? node1579 : 14'b00000000000001;
									assign node1579 = (inp[6]) ? 14'b00000000000001 : node1580;
										assign node1580 = (inp[9]) ? 14'b00000000000001 : node1581;
											assign node1581 = (inp[1]) ? 14'b00000000000001 : node1582;
												assign node1582 = (inp[11]) ? 14'b10001000001000 : 14'b00000000000001;
						assign node1588 = (inp[12]) ? node1656 : node1589;
							assign node1589 = (inp[5]) ? node1605 : node1590;
								assign node1590 = (inp[10]) ? 14'b00000000000001 : node1591;
									assign node1591 = (inp[11]) ? 14'b00000000000001 : node1592;
										assign node1592 = (inp[13]) ? 14'b00000000000001 : node1593;
											assign node1593 = (inp[7]) ? node1597 : node1594;
												assign node1594 = (inp[6]) ? 14'b00111000010110 : 14'b00000000000001;
												assign node1597 = (inp[1]) ? 14'b00101010110110 : node1598;
													assign node1598 = (inp[6]) ? 14'b00101100010110 : 14'b00101110010110;
								assign node1605 = (inp[11]) ? node1645 : node1606;
									assign node1606 = (inp[13]) ? node1634 : node1607;
										assign node1607 = (inp[10]) ? node1623 : node1608;
											assign node1608 = (inp[6]) ? node1616 : node1609;
												assign node1609 = (inp[7]) ? node1613 : node1610;
													assign node1610 = (inp[1]) ? 14'b00100000000110 : 14'b00000000000000;
													assign node1613 = (inp[1]) ? 14'b00100010110110 : 14'b00100110110110;
												assign node1616 = (inp[9]) ? node1620 : node1617;
													assign node1617 = (inp[1]) ? 14'b00110000110110 : 14'b00110100110110;
													assign node1620 = (inp[1]) ? 14'b00110000010110 : 14'b00110100010110;
											assign node1623 = (inp[1]) ? node1627 : node1624;
												assign node1624 = (inp[6]) ? 14'b00100100010000 : 14'b00100110010000;
												assign node1627 = (inp[7]) ? node1631 : node1628;
													assign node1628 = (inp[9]) ? 14'b00110000010000 : 14'b00110000110000;
													assign node1631 = (inp[9]) ? 14'b00100000010000 : 14'b00100000110000;
										assign node1634 = (inp[7]) ? 14'b00000000000001 : node1635;
											assign node1635 = (inp[1]) ? node1641 : node1636;
												assign node1636 = (inp[9]) ? node1638 : 14'b00000000000001;
													assign node1638 = (inp[6]) ? 14'b00010100010000 : 14'b00000100000000;
												assign node1641 = (inp[6]) ? 14'b00010100100000 : 14'b00010110100000;
									assign node1645 = (inp[7]) ? 14'b00000000000001 : node1646;
										assign node1646 = (inp[13]) ? node1648 : 14'b00000000000001;
											assign node1648 = (inp[1]) ? node1650 : 14'b00010100010000;
												assign node1650 = (inp[6]) ? 14'b00010100100000 : node1651;
													assign node1651 = (inp[9]) ? 14'b00010110000000 : 14'b00010110100000;
							assign node1656 = (inp[9]) ? 14'b00000000000001 : node1657;
								assign node1657 = (inp[10]) ? 14'b00000000000001 : node1658;
									assign node1658 = (inp[7]) ? node1660 : 14'b00000000000001;
										assign node1660 = (inp[5]) ? node1662 : 14'b00000000000001;
											assign node1662 = (inp[1]) ? 14'b00000000000001 : node1663;
												assign node1663 = (inp[6]) ? 14'b00000000000001 : 14'b10001001000010;
				assign node1669 = (inp[6]) ? node1995 : node1670;
					assign node1670 = (inp[7]) ? node1920 : node1671;
						assign node1671 = (inp[12]) ? node1829 : node1672;
							assign node1672 = (inp[11]) ? node1764 : node1673;
								assign node1673 = (inp[13]) ? node1721 : node1674;
									assign node1674 = (inp[5]) ? node1696 : node1675;
										assign node1675 = (inp[10]) ? node1683 : node1676;
											assign node1676 = (inp[4]) ? 14'b01111110010110 : node1677;
												assign node1677 = (inp[2]) ? node1679 : 14'b00000000000001;
													assign node1679 = (inp[9]) ? 14'b00011110010000 : 14'b00011110110000;
											assign node1683 = (inp[4]) ? node1691 : node1684;
												assign node1684 = (inp[9]) ? node1688 : node1685;
													assign node1685 = (inp[1]) ? 14'b00111010110010 : 14'b00111110110010;
													assign node1688 = (inp[2]) ? 14'b00111110010010 : 14'b01111110010010;
												assign node1691 = (inp[9]) ? node1693 : 14'b00000000000001;
													assign node1693 = (inp[1]) ? 14'b01111010010000 : 14'b01111110010000;
										assign node1696 = (inp[9]) ? node1708 : node1697;
											assign node1697 = (inp[1]) ? node1701 : node1698;
												assign node1698 = (inp[2]) ? 14'b00010110110000 : 14'b01110110110110;
												assign node1701 = (inp[10]) ? node1705 : node1702;
													assign node1702 = (inp[2]) ? 14'b00110010110110 : 14'b00110010110010;
													assign node1705 = (inp[4]) ? 14'b00110010110000 : 14'b01110010110010;
											assign node1708 = (inp[2]) ? node1716 : node1709;
												assign node1709 = (inp[1]) ? node1713 : node1710;
													assign node1710 = (inp[10]) ? 14'b01110110010000 : 14'b00110110010010;
													assign node1713 = (inp[10]) ? 14'b01110010010000 : 14'b01110010010110;
												assign node1716 = (inp[4]) ? node1718 : 14'b00000000000001;
													assign node1718 = (inp[10]) ? 14'b00110010010000 : 14'b00110010010110;
									assign node1721 = (inp[1]) ? node1745 : node1722;
										assign node1722 = (inp[4]) ? node1732 : node1723;
											assign node1723 = (inp[9]) ? node1727 : node1724;
												assign node1724 = (inp[2]) ? 14'b00000000000001 : 14'b01110110110000;
												assign node1727 = (inp[2]) ? node1729 : 14'b00000000000001;
													assign node1729 = (inp[5]) ? 14'b00000000000001 : 14'b01110110010100;
											assign node1732 = (inp[2]) ? node1740 : node1733;
												assign node1733 = (inp[5]) ? node1737 : node1734;
													assign node1734 = (inp[9]) ? 14'b00110110010100 : 14'b00110110110100;
													assign node1737 = (inp[9]) ? 14'b00110110010000 : 14'b00110110110000;
												assign node1740 = (inp[5]) ? node1742 : 14'b00000000000001;
													assign node1742 = (inp[9]) ? 14'b00010110010000 : 14'b00010110110000;
										assign node1745 = (inp[4]) ? node1751 : node1746;
											assign node1746 = (inp[9]) ? node1748 : 14'b00000000000001;
												assign node1748 = (inp[10]) ? 14'b00000000000001 : 14'b01100110000100;
											assign node1751 = (inp[2]) ? node1759 : node1752;
												assign node1752 = (inp[5]) ? node1756 : node1753;
													assign node1753 = (inp[9]) ? 14'b00100110000100 : 14'b00100110100100;
													assign node1756 = (inp[9]) ? 14'b00100110000000 : 14'b00100110100000;
												assign node1759 = (inp[5]) ? node1761 : 14'b00000000000001;
													assign node1761 = (inp[9]) ? 14'b00000110000000 : 14'b00000110100000;
								assign node1764 = (inp[13]) ? node1780 : node1765;
									assign node1765 = (inp[10]) ? 14'b00000000000001 : node1766;
										assign node1766 = (inp[4]) ? 14'b00000000000001 : node1767;
											assign node1767 = (inp[2]) ? node1773 : node1768;
												assign node1768 = (inp[9]) ? 14'b01110110010100 : node1769;
													assign node1769 = (inp[5]) ? 14'b01110010110100 : 14'b01111010110100;
												assign node1773 = (inp[5]) ? 14'b00110010110100 : node1774;
													assign node1774 = (inp[9]) ? 14'b00111010010100 : 14'b00111010110100;
									assign node1780 = (inp[4]) ? node1808 : node1781;
										assign node1781 = (inp[1]) ? node1797 : node1782;
											assign node1782 = (inp[9]) ? node1790 : node1783;
												assign node1783 = (inp[5]) ? node1787 : node1784;
													assign node1784 = (inp[2]) ? 14'b01110110110100 : 14'b00000000000001;
													assign node1787 = (inp[2]) ? 14'b00000000000001 : 14'b01110110110000;
												assign node1790 = (inp[2]) ? node1794 : node1791;
													assign node1791 = (inp[5]) ? 14'b01110110010000 : 14'b00000000000001;
													assign node1794 = (inp[5]) ? 14'b00000000000001 : 14'b01110110010100;
											assign node1797 = (inp[5]) ? node1803 : node1798;
												assign node1798 = (inp[2]) ? node1800 : 14'b00000000000001;
													assign node1800 = (inp[9]) ? 14'b01100110000100 : 14'b01100110100100;
												assign node1803 = (inp[2]) ? 14'b00000000000001 : node1804;
													assign node1804 = (inp[10]) ? 14'b01100110100000 : 14'b01100110000000;
										assign node1808 = (inp[2]) ? node1820 : node1809;
											assign node1809 = (inp[1]) ? node1817 : node1810;
												assign node1810 = (inp[5]) ? node1814 : node1811;
													assign node1811 = (inp[9]) ? 14'b00110110010100 : 14'b00110110110100;
													assign node1814 = (inp[9]) ? 14'b00110110010000 : 14'b00110110110000;
												assign node1817 = (inp[10]) ? 14'b00100110000000 : 14'b00100110000100;
											assign node1820 = (inp[5]) ? node1822 : 14'b00000000000001;
												assign node1822 = (inp[1]) ? node1826 : node1823;
													assign node1823 = (inp[9]) ? 14'b00010110010000 : 14'b00010110110000;
													assign node1826 = (inp[9]) ? 14'b00000110000000 : 14'b00000110100000;
							assign node1829 = (inp[5]) ? node1885 : node1830;
								assign node1830 = (inp[13]) ? node1862 : node1831;
									assign node1831 = (inp[11]) ? node1851 : node1832;
										assign node1832 = (inp[4]) ? node1844 : node1833;
											assign node1833 = (inp[2]) ? node1841 : node1834;
												assign node1834 = (inp[9]) ? node1838 : node1835;
													assign node1835 = (inp[10]) ? 14'b01011010110010 : 14'b01011010110110;
													assign node1838 = (inp[10]) ? 14'b01011010010010 : 14'b01011010010110;
												assign node1841 = (inp[1]) ? 14'b00011010110010 : 14'b00011110110010;
											assign node1844 = (inp[10]) ? node1846 : 14'b00000000000001;
												assign node1846 = (inp[9]) ? node1848 : 14'b00111010110000;
													assign node1848 = (inp[1]) ? 14'b00111010010000 : 14'b00111110010000;
										assign node1851 = (inp[10]) ? 14'b00000000000001 : node1852;
											assign node1852 = (inp[2]) ? 14'b00000000000001 : node1853;
												assign node1853 = (inp[9]) ? node1857 : node1854;
													assign node1854 = (inp[4]) ? 14'b01011110110000 : 14'b01011110110100;
													assign node1857 = (inp[4]) ? 14'b01011110010000 : 14'b01011110010100;
									assign node1862 = (inp[2]) ? node1876 : node1863;
										assign node1863 = (inp[1]) ? node1871 : node1864;
											assign node1864 = (inp[4]) ? node1868 : node1865;
												assign node1865 = (inp[9]) ? 14'b01010110010100 : 14'b01010110110100;
												assign node1868 = (inp[9]) ? 14'b00010110010100 : 14'b00010110110100;
											assign node1871 = (inp[4]) ? 14'b00000110100100 : node1872;
												assign node1872 = (inp[9]) ? 14'b01000110000100 : 14'b01000110100100;
										assign node1876 = (inp[4]) ? 14'b00000000000001 : node1877;
											assign node1877 = (inp[1]) ? node1881 : node1878;
												assign node1878 = (inp[9]) ? 14'b01010110010000 : 14'b01010110110000;
												assign node1881 = (inp[9]) ? 14'b01000110000000 : 14'b01000110100000;
								assign node1885 = (inp[13]) ? 14'b00000000000001 : node1886;
									assign node1886 = (inp[10]) ? node1912 : node1887;
										assign node1887 = (inp[2]) ? node1903 : node1888;
											assign node1888 = (inp[1]) ? node1896 : node1889;
												assign node1889 = (inp[11]) ? node1893 : node1890;
													assign node1890 = (inp[9]) ? 14'b01010110010010 : 14'b01010110110010;
													assign node1893 = (inp[4]) ? 14'b01010110110000 : 14'b01010110110100;
												assign node1896 = (inp[11]) ? node1900 : node1897;
													assign node1897 = (inp[4]) ? 14'b01010010010010 : 14'b01010010010110;
													assign node1900 = (inp[4]) ? 14'b01010010010000 : 14'b01010010010100;
											assign node1903 = (inp[4]) ? 14'b00000000000001 : node1904;
												assign node1904 = (inp[9]) ? node1908 : node1905;
													assign node1905 = (inp[11]) ? 14'b00010110110100 : 14'b00010110110110;
													assign node1908 = (inp[1]) ? 14'b00010010010100 : 14'b00010110010100;
										assign node1912 = (inp[2]) ? node1914 : 14'b00000000000001;
											assign node1914 = (inp[4]) ? 14'b00000000000001 : node1915;
												assign node1915 = (inp[11]) ? 14'b00000000000001 : 14'b00010010110010;
						assign node1920 = (inp[13]) ? node1936 : node1921;
							assign node1921 = (inp[5]) ? 14'b00000000000001 : node1922;
								assign node1922 = (inp[1]) ? 14'b00000000000001 : node1923;
									assign node1923 = (inp[9]) ? 14'b00000000000001 : node1924;
										assign node1924 = (inp[10]) ? 14'b00000000000001 : node1925;
											assign node1925 = (inp[2]) ? 14'b00000000000001 : node1926;
												assign node1926 = (inp[4]) ? node1928 : 14'b00000000000001;
													assign node1928 = (inp[12]) ? 14'b00000000000001 : 14'b10000001000000;
							assign node1936 = (inp[5]) ? node1978 : node1937;
								assign node1937 = (inp[4]) ? node1965 : node1938;
									assign node1938 = (inp[1]) ? node1950 : node1939;
										assign node1939 = (inp[9]) ? node1945 : node1940;
											assign node1940 = (inp[12]) ? node1942 : 14'b00010010110000;
												assign node1942 = (inp[2]) ? 14'b01010010110000 : 14'b01010010110100;
											assign node1945 = (inp[12]) ? node1947 : 14'b01110010010100;
												assign node1947 = (inp[11]) ? 14'b01010010010100 : 14'b01010010010000;
										assign node1950 = (inp[9]) ? node1958 : node1951;
											assign node1951 = (inp[12]) ? node1955 : node1952;
												assign node1952 = (inp[2]) ? 14'b01100010100100 : 14'b00000010100000;
												assign node1955 = (inp[2]) ? 14'b01000010100000 : 14'b01000010100100;
											assign node1958 = (inp[12]) ? node1962 : node1959;
												assign node1959 = (inp[2]) ? 14'b01100010000100 : 14'b00000010000000;
												assign node1962 = (inp[2]) ? 14'b01000010000000 : 14'b01000010000100;
									assign node1965 = (inp[2]) ? 14'b00000000000001 : node1966;
										assign node1966 = (inp[1]) ? node1972 : node1967;
											assign node1967 = (inp[12]) ? 14'b00010010110100 : node1968;
												assign node1968 = (inp[9]) ? 14'b00110010010100 : 14'b00110010110100;
											assign node1972 = (inp[9]) ? 14'b00100010000100 : node1973;
												assign node1973 = (inp[12]) ? 14'b00000010100100 : 14'b00100010100100;
								assign node1978 = (inp[12]) ? 14'b00000000000001 : node1979;
									assign node1979 = (inp[2]) ? 14'b00000000000001 : node1980;
										assign node1980 = (inp[1]) ? node1988 : node1981;
											assign node1981 = (inp[4]) ? node1985 : node1982;
												assign node1982 = (inp[9]) ? 14'b01110010010000 : 14'b01110010110000;
												assign node1985 = (inp[9]) ? 14'b00110010010000 : 14'b00110010110000;
											assign node1988 = (inp[9]) ? 14'b01100010000000 : node1989;
												assign node1989 = (inp[4]) ? 14'b00100010100000 : 14'b01100010100000;
					assign node1995 = (inp[9]) ? 14'b00000000000001 : node1996;
						assign node1996 = (inp[13]) ? node2114 : node1997;
							assign node1997 = (inp[1]) ? node2045 : node1998;
								assign node1998 = (inp[7]) ? node2010 : node1999;
									assign node1999 = (inp[11]) ? node2001 : 14'b00000000000001;
										assign node2001 = (inp[2]) ? 14'b00000000000001 : node2002;
											assign node2002 = (inp[4]) ? node2004 : 14'b00000000000001;
												assign node2004 = (inp[5]) ? 14'b00000000000001 : node2005;
													assign node2005 = (inp[12]) ? 14'b00000000000001 : 14'b10000001001000;
									assign node2010 = (inp[10]) ? node2032 : node2011;
										assign node2011 = (inp[12]) ? node2019 : node2012;
											assign node2012 = (inp[4]) ? node2016 : node2013;
												assign node2013 = (inp[11]) ? 14'b01101100100100 : 14'b00000000000001;
												assign node2016 = (inp[5]) ? 14'b00100100100110 : 14'b01101100100110;
											assign node2019 = (inp[4]) ? node2027 : node2020;
												assign node2020 = (inp[2]) ? node2024 : node2021;
													assign node2021 = (inp[5]) ? 14'b01000100100100 : 14'b01001100100100;
													assign node2024 = (inp[11]) ? 14'b00000100100100 : 14'b00000100100110;
												assign node2027 = (inp[5]) ? node2029 : 14'b00000000000001;
													assign node2029 = (inp[2]) ? 14'b00000000000001 : 14'b01000100100010;
										assign node2032 = (inp[11]) ? 14'b00000000000001 : node2033;
											assign node2033 = (inp[2]) ? node2039 : node2034;
												assign node2034 = (inp[4]) ? node2036 : 14'b01001100100010;
													assign node2036 = (inp[12]) ? 14'b00101100100000 : 14'b01101100100000;
												assign node2039 = (inp[5]) ? node2041 : 14'b00000000000001;
													assign node2041 = (inp[4]) ? 14'b00100100100000 : 14'b00000000000001;
								assign node2045 = (inp[10]) ? node2091 : node2046;
									assign node2046 = (inp[2]) ? node2068 : node2047;
										assign node2047 = (inp[5]) ? node2059 : node2048;
											assign node2048 = (inp[12]) ? node2056 : node2049;
												assign node2049 = (inp[7]) ? node2053 : node2050;
													assign node2050 = (inp[11]) ? 14'b00000000000000 : 14'b01111000100110;
													assign node2053 = (inp[4]) ? 14'b01101000100110 : 14'b00000000000000;
												assign node2056 = (inp[11]) ? 14'b01011000100000 : 14'b00000000000001;
											assign node2059 = (inp[7]) ? node2063 : node2060;
												assign node2060 = (inp[4]) ? 14'b01010000100010 : 14'b01010000100100;
												assign node2063 = (inp[11]) ? 14'b01000000100000 : node2064;
													assign node2064 = (inp[12]) ? 14'b01000000100010 : 14'b01100000100110;
										assign node2068 = (inp[4]) ? node2084 : node2069;
											assign node2069 = (inp[12]) ? node2077 : node2070;
												assign node2070 = (inp[11]) ? node2074 : node2071;
													assign node2071 = (inp[5]) ? 14'b00010000100000 : 14'b00011000100000;
													assign node2074 = (inp[5]) ? 14'b00110000100100 : 14'b00101000100100;
												assign node2077 = (inp[5]) ? node2081 : node2078;
													assign node2078 = (inp[7]) ? 14'b00001000100110 : 14'b00011000100110;
													assign node2081 = (inp[11]) ? 14'b00000000100100 : 14'b00000000100110;
											assign node2084 = (inp[11]) ? 14'b00000000000001 : node2085;
												assign node2085 = (inp[12]) ? 14'b00000000000001 : node2086;
													assign node2086 = (inp[7]) ? 14'b00101000100110 : 14'b00110000100110;
									assign node2091 = (inp[11]) ? 14'b00000000000001 : node2092;
										assign node2092 = (inp[2]) ? node2102 : node2093;
											assign node2093 = (inp[5]) ? 14'b00000000000001 : node2094;
												assign node2094 = (inp[4]) ? node2098 : node2095;
													assign node2095 = (inp[7]) ? 14'b01001000100010 : 14'b01011000100010;
													assign node2098 = (inp[7]) ? 14'b00101000100000 : 14'b00111000100000;
											assign node2102 = (inp[4]) ? node2108 : node2103;
												assign node2103 = (inp[5]) ? 14'b00000000000001 : node2104;
													assign node2104 = (inp[12]) ? 14'b00001000100010 : 14'b00101000100010;
												assign node2108 = (inp[5]) ? node2110 : 14'b00000000000001;
													assign node2110 = (inp[12]) ? 14'b00000000000001 : 14'b00110000100000;
							assign node2114 = (inp[1]) ? node2134 : node2115;
								assign node2115 = (inp[7]) ? 14'b00000000000001 : node2116;
									assign node2116 = (inp[4]) ? node2126 : node2117;
										assign node2117 = (inp[5]) ? node2119 : 14'b00000000000001;
											assign node2119 = (inp[12]) ? node2123 : node2120;
												assign node2120 = (inp[2]) ? 14'b10000001001000 : 14'b00000000000001;
												assign node2123 = (inp[2]) ? 14'b00000000000001 : 14'b10001000000010;
										assign node2126 = (inp[2]) ? node2128 : 14'b00000000000001;
											assign node2128 = (inp[12]) ? 14'b00000000000001 : node2129;
												assign node2129 = (inp[5]) ? 14'b00000000000001 : 14'b10000001001010;
								assign node2134 = (inp[12]) ? 14'b00000000000001 : node2135;
									assign node2135 = (inp[4]) ? node2137 : 14'b00000000000001;
										assign node2137 = (inp[2]) ? node2139 : 14'b00000000000001;
											assign node2139 = (inp[7]) ? 14'b10000000000000 : 14'b00000000000001;
			assign node2144 = (inp[7]) ? node2674 : node2145;
				assign node2145 = (inp[1]) ? node2473 : node2146;
					assign node2146 = (inp[9]) ? node2368 : node2147;
						assign node2147 = (inp[13]) ? node2285 : node2148;
							assign node2148 = (inp[10]) ? node2238 : node2149;
								assign node2149 = (inp[4]) ? node2209 : node2150;
									assign node2150 = (inp[3]) ? node2180 : node2151;
										assign node2151 = (inp[6]) ? node2167 : node2152;
											assign node2152 = (inp[12]) ? node2160 : node2153;
												assign node2153 = (inp[11]) ? node2157 : node2154;
													assign node2154 = (inp[2]) ? 14'b00010110100000 : 14'b00000000000001;
													assign node2157 = (inp[5]) ? 14'b00110110100100 : 14'b00111110100100;
												assign node2160 = (inp[5]) ? node2164 : node2161;
													assign node2161 = (inp[11]) ? 14'b01011110100100 : 14'b01011110100110;
													assign node2164 = (inp[11]) ? 14'b00010110100100 : 14'b00010110100110;
											assign node2167 = (inp[12]) ? node2173 : node2168;
												assign node2168 = (inp[11]) ? node2170 : 14'b00110100100010;
													assign node2170 = (inp[5]) ? 14'b00110100100100 : 14'b01111100100100;
												assign node2173 = (inp[2]) ? node2177 : node2174;
													assign node2174 = (inp[5]) ? 14'b01010100100100 : 14'b01011100100100;
													assign node2177 = (inp[5]) ? 14'b00010100100100 : 14'b00011100100100;
										assign node2180 = (inp[6]) ? node2196 : node2181;
											assign node2181 = (inp[11]) ? node2189 : node2182;
												assign node2182 = (inp[12]) ? node2186 : node2183;
													assign node2183 = (inp[2]) ? 14'b00000110100000 : 14'b00100110100010;
													assign node2186 = (inp[2]) ? 14'b00000110100110 : 14'b01000110100110;
												assign node2189 = (inp[12]) ? node2193 : node2190;
													assign node2190 = (inp[2]) ? 14'b00100110100100 : 14'b01101110100100;
													assign node2193 = (inp[5]) ? 14'b00000110100100 : 14'b00001110100100;
											assign node2196 = (inp[11]) ? node2202 : node2197;
												assign node2197 = (inp[12]) ? 14'b01000110000110 : node2198;
													assign node2198 = (inp[2]) ? 14'b00000110000000 : 14'b00000000000001;
												assign node2202 = (inp[12]) ? node2206 : node2203;
													assign node2203 = (inp[2]) ? 14'b00100110000100 : 14'b01101110000100;
													assign node2206 = (inp[2]) ? 14'b00001110000100 : 14'b01000110000100;
									assign node2209 = (inp[11]) ? node2231 : node2210;
										assign node2210 = (inp[12]) ? node2224 : node2211;
											assign node2211 = (inp[3]) ? node2217 : node2212;
												assign node2212 = (inp[2]) ? node2214 : 14'b01110110100110;
													assign node2214 = (inp[5]) ? 14'b00110100100110 : 14'b00111110100110;
												assign node2217 = (inp[6]) ? node2221 : node2218;
													assign node2218 = (inp[2]) ? 14'b00101110100110 : 14'b01101110100110;
													assign node2221 = (inp[5]) ? 14'b00100110000110 : 14'b00101110000110;
											assign node2224 = (inp[5]) ? node2226 : 14'b00000000000001;
												assign node2226 = (inp[2]) ? 14'b00000000000001 : node2227;
													assign node2227 = (inp[6]) ? 14'b01000110000010 : 14'b01000110100010;
										assign node2231 = (inp[12]) ? node2233 : 14'b00000000000001;
											assign node2233 = (inp[2]) ? 14'b00000000000001 : node2234;
												assign node2234 = (inp[3]) ? 14'b01000110100000 : 14'b01010110100000;
								assign node2238 = (inp[11]) ? 14'b00000000000001 : node2239;
									assign node2239 = (inp[4]) ? node2265 : node2240;
										assign node2240 = (inp[5]) ? node2254 : node2241;
											assign node2241 = (inp[2]) ? node2247 : node2242;
												assign node2242 = (inp[3]) ? node2244 : 14'b01011110100010;
													assign node2244 = (inp[12]) ? 14'b01001110000010 : 14'b01101110000010;
												assign node2247 = (inp[3]) ? node2251 : node2248;
													assign node2248 = (inp[6]) ? 14'b00011100100010 : 14'b00011110100010;
													assign node2251 = (inp[12]) ? 14'b00001110100010 : 14'b00101110100010;
											assign node2254 = (inp[3]) ? node2260 : node2255;
												assign node2255 = (inp[2]) ? node2257 : 14'b01110100100010;
													assign node2257 = (inp[12]) ? 14'b00010110100010 : 14'b00000000000001;
												assign node2260 = (inp[2]) ? node2262 : 14'b00000000000001;
													assign node2262 = (inp[12]) ? 14'b00000110000010 : 14'b00000000000001;
										assign node2265 = (inp[2]) ? node2277 : node2266;
											assign node2266 = (inp[12]) ? node2272 : node2267;
												assign node2267 = (inp[6]) ? 14'b01100110000000 : node2268;
													assign node2268 = (inp[3]) ? 14'b01100110100000 : 14'b01110110100000;
												assign node2272 = (inp[5]) ? 14'b00000000000001 : node2273;
													assign node2273 = (inp[3]) ? 14'b00101110000000 : 14'b00111100100000;
											assign node2277 = (inp[3]) ? 14'b00000000000001 : node2278;
												assign node2278 = (inp[12]) ? 14'b00000000000001 : node2279;
													assign node2279 = (inp[5]) ? 14'b00110100100000 : 14'b00000000000001;
							assign node2285 = (inp[3]) ? node2333 : node2286;
								assign node2286 = (inp[5]) ? node2320 : node2287;
									assign node2287 = (inp[12]) ? node2307 : node2288;
										assign node2288 = (inp[10]) ? node2298 : node2289;
											assign node2289 = (inp[4]) ? node2295 : node2290;
												assign node2290 = (inp[2]) ? node2292 : 14'b00000000000001;
													assign node2292 = (inp[6]) ? 14'b01100100110100 : 14'b01100110110100;
												assign node2295 = (inp[2]) ? 14'b00000000000001 : 14'b00100110110100;
											assign node2298 = (inp[2]) ? node2304 : node2299;
												assign node2299 = (inp[4]) ? node2301 : 14'b00000000000001;
													assign node2301 = (inp[6]) ? 14'b00100100110100 : 14'b00100110110100;
												assign node2304 = (inp[11]) ? 14'b01100100110100 : 14'b01100110110100;
										assign node2307 = (inp[4]) ? node2315 : node2308;
											assign node2308 = (inp[6]) ? node2312 : node2309;
												assign node2309 = (inp[2]) ? 14'b01000110110000 : 14'b01000110110100;
												assign node2312 = (inp[2]) ? 14'b01000100110000 : 14'b01000100110100;
											assign node2315 = (inp[2]) ? 14'b00000000000001 : node2316;
												assign node2316 = (inp[6]) ? 14'b00000100110100 : 14'b00000110110100;
									assign node2320 = (inp[12]) ? 14'b00000000000001 : node2321;
										assign node2321 = (inp[4]) ? node2325 : node2322;
											assign node2322 = (inp[2]) ? 14'b00000000000001 : 14'b01100110110000;
											assign node2325 = (inp[6]) ? node2329 : node2326;
												assign node2326 = (inp[2]) ? 14'b00000110110000 : 14'b00100110110000;
												assign node2329 = (inp[2]) ? 14'b00000100110000 : 14'b00100100110000;
								assign node2333 = (inp[6]) ? node2343 : node2334;
									assign node2334 = (inp[12]) ? 14'b00000000000001 : node2335;
										assign node2335 = (inp[2]) ? node2337 : 14'b00000000000001;
											assign node2337 = (inp[4]) ? 14'b00000000000001 : node2338;
												assign node2338 = (inp[5]) ? 14'b10000001000000 : 14'b00000000000001;
									assign node2343 = (inp[2]) ? node2357 : node2344;
										assign node2344 = (inp[5]) ? node2352 : node2345;
											assign node2345 = (inp[12]) ? node2349 : node2346;
												assign node2346 = (inp[4]) ? 14'b00100100100100 : 14'b00000000000001;
												assign node2349 = (inp[4]) ? 14'b00000100100100 : 14'b01000100100100;
											assign node2352 = (inp[12]) ? 14'b00000000000001 : node2353;
												assign node2353 = (inp[4]) ? 14'b00100100100000 : 14'b01100100100000;
										assign node2357 = (inp[4]) ? node2363 : node2358;
											assign node2358 = (inp[5]) ? 14'b00000000000001 : node2359;
												assign node2359 = (inp[12]) ? 14'b01000100100000 : 14'b01100100100100;
											assign node2363 = (inp[5]) ? node2365 : 14'b00000000000001;
												assign node2365 = (inp[12]) ? 14'b00000000000001 : 14'b00000100100000;
						assign node2368 = (inp[3]) ? 14'b00000000000001 : node2369;
							assign node2369 = (inp[13]) ? node2433 : node2370;
								assign node2370 = (inp[10]) ? node2408 : node2371;
									assign node2371 = (inp[4]) ? node2393 : node2372;
										assign node2372 = (inp[12]) ? node2382 : node2373;
											assign node2373 = (inp[11]) ? node2377 : node2374;
												assign node2374 = (inp[6]) ? 14'b00110100000010 : 14'b00110110000010;
												assign node2377 = (inp[6]) ? 14'b01110100000100 : node2378;
													assign node2378 = (inp[5]) ? 14'b00110110000100 : 14'b00111110000100;
											assign node2382 = (inp[5]) ? node2388 : node2383;
												assign node2383 = (inp[11]) ? node2385 : 14'b00011100000110;
													assign node2385 = (inp[6]) ? 14'b01011100000100 : 14'b01011110000100;
												assign node2388 = (inp[11]) ? 14'b00010100000100 : node2389;
													assign node2389 = (inp[2]) ? 14'b00010100000110 : 14'b01010100000110;
										assign node2393 = (inp[11]) ? node2403 : node2394;
											assign node2394 = (inp[12]) ? 14'b00000000000001 : node2395;
												assign node2395 = (inp[6]) ? node2399 : node2396;
													assign node2396 = (inp[2]) ? 14'b00111110000110 : 14'b01111110000110;
													assign node2399 = (inp[5]) ? 14'b01110100000110 : 14'b01111100000110;
											assign node2403 = (inp[6]) ? node2405 : 14'b00000000000001;
												assign node2405 = (inp[5]) ? 14'b01010100000000 : 14'b00000000000001;
									assign node2408 = (inp[11]) ? 14'b00000000000001 : node2409;
										assign node2409 = (inp[4]) ? node2421 : node2410;
											assign node2410 = (inp[5]) ? node2414 : node2411;
												assign node2411 = (inp[6]) ? 14'b01011100000010 : 14'b00011110000010;
												assign node2414 = (inp[12]) ? node2418 : node2415;
													assign node2415 = (inp[2]) ? 14'b00000000000001 : 14'b01110100000010;
													assign node2418 = (inp[2]) ? 14'b00010110000010 : 14'b00000000000001;
											assign node2421 = (inp[2]) ? node2427 : node2422;
												assign node2422 = (inp[5]) ? node2424 : 14'b00111100000000;
													assign node2424 = (inp[12]) ? 14'b00000000000001 : 14'b01110100000000;
												assign node2427 = (inp[6]) ? 14'b00000000000001 : node2428;
													assign node2428 = (inp[5]) ? 14'b00000000000000 : 14'b00000000000001;
								assign node2433 = (inp[2]) ? node2457 : node2434;
									assign node2434 = (inp[5]) ? node2448 : node2435;
										assign node2435 = (inp[12]) ? node2441 : node2436;
											assign node2436 = (inp[4]) ? node2438 : 14'b00000000000001;
												assign node2438 = (inp[11]) ? 14'b00100110010100 : 14'b00100100010100;
											assign node2441 = (inp[4]) ? node2445 : node2442;
												assign node2442 = (inp[6]) ? 14'b01000100010100 : 14'b01000110010100;
												assign node2445 = (inp[6]) ? 14'b00000100010100 : 14'b00000110010100;
										assign node2448 = (inp[12]) ? 14'b00000000000001 : node2449;
											assign node2449 = (inp[4]) ? node2453 : node2450;
												assign node2450 = (inp[6]) ? 14'b01100100010000 : 14'b01100110010000;
												assign node2453 = (inp[6]) ? 14'b00100100010000 : 14'b00100110010000;
									assign node2457 = (inp[5]) ? node2465 : node2458;
										assign node2458 = (inp[4]) ? 14'b00000000000001 : node2459;
											assign node2459 = (inp[12]) ? node2461 : 14'b01100100010100;
												assign node2461 = (inp[6]) ? 14'b01000100010000 : 14'b01000110010000;
										assign node2465 = (inp[4]) ? node2467 : 14'b00000000000001;
											assign node2467 = (inp[12]) ? 14'b00000000000001 : node2468;
												assign node2468 = (inp[6]) ? 14'b00000100010000 : 14'b00000110010000;
					assign node2473 = (inp[13]) ? node2639 : node2474;
						assign node2474 = (inp[6]) ? node2586 : node2475;
							assign node2475 = (inp[11]) ? node2551 : node2476;
								assign node2476 = (inp[9]) ? node2528 : node2477;
									assign node2477 = (inp[4]) ? node2505 : node2478;
										assign node2478 = (inp[12]) ? node2492 : node2479;
											assign node2479 = (inp[10]) ? node2485 : node2480;
												assign node2480 = (inp[5]) ? node2482 : 14'b00000000000001;
													assign node2482 = (inp[2]) ? 14'b00000010100000 : 14'b00100010100010;
												assign node2485 = (inp[2]) ? node2489 : node2486;
													assign node2486 = (inp[3]) ? 14'b01100010100010 : 14'b01110010100010;
													assign node2489 = (inp[5]) ? 14'b00000000000001 : 14'b00101010100010;
											assign node2492 = (inp[5]) ? node2500 : node2493;
												assign node2493 = (inp[3]) ? node2497 : node2494;
													assign node2494 = (inp[10]) ? 14'b00011010100010 : 14'b00011010100110;
													assign node2497 = (inp[2]) ? 14'b00001010100010 : 14'b01001010100010;
												assign node2500 = (inp[10]) ? node2502 : 14'b01010010100110;
													assign node2502 = (inp[2]) ? 14'b00000010100010 : 14'b00000000000001;
										assign node2505 = (inp[12]) ? node2521 : node2506;
											assign node2506 = (inp[10]) ? node2514 : node2507;
												assign node2507 = (inp[2]) ? node2511 : node2508;
													assign node2508 = (inp[3]) ? 14'b01101010100110 : 14'b01111010100110;
													assign node2511 = (inp[5]) ? 14'b00110010100110 : 14'b00111010100110;
												assign node2514 = (inp[2]) ? node2518 : node2515;
													assign node2515 = (inp[3]) ? 14'b01101010100000 : 14'b01111010100000;
													assign node2518 = (inp[5]) ? 14'b00100010100000 : 14'b00000000000001;
											assign node2521 = (inp[3]) ? node2523 : 14'b00000000000001;
												assign node2523 = (inp[5]) ? 14'b00000000000001 : node2524;
													assign node2524 = (inp[10]) ? 14'b00101010100000 : 14'b00000000000001;
									assign node2528 = (inp[3]) ? node2530 : 14'b00000000000001;
										assign node2530 = (inp[2]) ? node2544 : node2531;
											assign node2531 = (inp[12]) ? node2539 : node2532;
												assign node2532 = (inp[10]) ? node2536 : node2533;
													assign node2533 = (inp[4]) ? 14'b01101010000110 : 14'b00000000000000;
													assign node2536 = (inp[5]) ? 14'b01100010000000 : 14'b01101010000000;
												assign node2539 = (inp[10]) ? 14'b00000000000001 : node2540;
													assign node2540 = (inp[5]) ? 14'b01000010000010 : 14'b01001010000110;
											assign node2544 = (inp[4]) ? 14'b00000000000001 : node2545;
												assign node2545 = (inp[5]) ? 14'b00000000000001 : node2546;
													assign node2546 = (inp[12]) ? 14'b00001010000010 : 14'b00001010000000;
								assign node2551 = (inp[10]) ? 14'b00000000000001 : node2552;
									assign node2552 = (inp[4]) ? node2574 : node2553;
										assign node2553 = (inp[9]) ? node2565 : node2554;
											assign node2554 = (inp[3]) ? node2562 : node2555;
												assign node2555 = (inp[5]) ? node2559 : node2556;
													assign node2556 = (inp[2]) ? 14'b00011010100100 : 14'b01111010100100;
													assign node2559 = (inp[12]) ? 14'b01010010100100 : 14'b00110010100100;
												assign node2562 = (inp[12]) ? 14'b00000010100100 : 14'b00100010100100;
											assign node2565 = (inp[3]) ? node2567 : 14'b00000000000001;
												assign node2567 = (inp[2]) ? node2571 : node2568;
													assign node2568 = (inp[12]) ? 14'b01000010000100 : 14'b01100010000100;
													assign node2571 = (inp[12]) ? 14'b00000010000100 : 14'b00100010000100;
										assign node2574 = (inp[2]) ? 14'b00000000000001 : node2575;
											assign node2575 = (inp[12]) ? node2577 : 14'b00000000000001;
												assign node2577 = (inp[9]) ? node2581 : node2578;
													assign node2578 = (inp[3]) ? 14'b01001010100000 : 14'b01010010100000;
													assign node2581 = (inp[3]) ? 14'b01001010000000 : 14'b00000000000001;
							assign node2586 = (inp[9]) ? node2598 : node2587;
								assign node2587 = (inp[10]) ? 14'b00000000000001 : node2588;
									assign node2588 = (inp[5]) ? 14'b00000000000001 : node2589;
										assign node2589 = (inp[4]) ? node2591 : 14'b00000000000001;
											assign node2591 = (inp[11]) ? node2593 : 14'b00000000000001;
												assign node2593 = (inp[12]) ? 14'b10000000000000 : 14'b00000000000001;
								assign node2598 = (inp[3]) ? 14'b00000000000001 : node2599;
									assign node2599 = (inp[10]) ? node2621 : node2600;
										assign node2600 = (inp[4]) ? node2614 : node2601;
											assign node2601 = (inp[11]) ? node2607 : node2602;
												assign node2602 = (inp[5]) ? node2604 : 14'b00000000000001;
													assign node2604 = (inp[2]) ? 14'b00010000000000 : 14'b00110000000010;
												assign node2607 = (inp[12]) ? node2611 : node2608;
													assign node2608 = (inp[5]) ? 14'b01110000000100 : 14'b00111000000100;
													assign node2611 = (inp[5]) ? 14'b01010000000100 : 14'b01011000000100;
											assign node2614 = (inp[11]) ? 14'b00000000000001 : node2615;
												assign node2615 = (inp[12]) ? 14'b00000000000001 : node2616;
													assign node2616 = (inp[2]) ? 14'b00111000000110 : 14'b01110000000110;
										assign node2621 = (inp[11]) ? 14'b00000000000001 : node2622;
											assign node2622 = (inp[4]) ? node2630 : node2623;
												assign node2623 = (inp[12]) ? node2627 : node2624;
													assign node2624 = (inp[2]) ? 14'b00111000000010 : 14'b01110000000010;
													assign node2627 = (inp[5]) ? 14'b00000000000001 : 14'b00011000000010;
												assign node2630 = (inp[2]) ? node2634 : node2631;
													assign node2631 = (inp[5]) ? 14'b00000000000001 : 14'b00111000000000;
													assign node2634 = (inp[12]) ? 14'b00000000000001 : 14'b00000000000000;
						assign node2639 = (inp[6]) ? 14'b00000000000001 : node2640;
							assign node2640 = (inp[4]) ? node2662 : node2641;
								assign node2641 = (inp[5]) ? node2649 : node2642;
									assign node2642 = (inp[9]) ? node2644 : 14'b00000000000001;
										assign node2644 = (inp[3]) ? node2646 : 14'b00000000000001;
											assign node2646 = (inp[12]) ? 14'b00000000000001 : 14'b10000000000010;
									assign node2649 = (inp[3]) ? 14'b00000000000001 : node2650;
										assign node2650 = (inp[9]) ? 14'b00000000000001 : node2651;
											assign node2651 = (inp[10]) ? node2657 : node2652;
												assign node2652 = (inp[2]) ? node2654 : 14'b00000000000001;
													assign node2654 = (inp[12]) ? 14'b00000000000001 : 14'b10000000001010;
												assign node2657 = (inp[2]) ? 14'b00000000000001 : 14'b10001001001000;
								assign node2662 = (inp[12]) ? 14'b00000000000001 : node2663;
									assign node2663 = (inp[3]) ? 14'b00000000000001 : node2664;
										assign node2664 = (inp[2]) ? node2666 : 14'b00000000000001;
											assign node2666 = (inp[5]) ? 14'b00000000000001 : node2667;
												assign node2667 = (inp[10]) ? 14'b10000001000010 : 14'b00000000000001;
				assign node2674 = (inp[13]) ? node2676 : 14'b00000000000001;
					assign node2676 = (inp[1]) ? node2764 : node2677;
						assign node2677 = (inp[3]) ? node2739 : node2678;
							assign node2678 = (inp[2]) ? node2724 : node2679;
								assign node2679 = (inp[12]) ? node2709 : node2680;
									assign node2680 = (inp[6]) ? node2696 : node2681;
										assign node2681 = (inp[9]) ? node2689 : node2682;
											assign node2682 = (inp[5]) ? node2686 : node2683;
												assign node2683 = (inp[4]) ? 14'b00100010110100 : 14'b00000010110000;
												assign node2686 = (inp[4]) ? 14'b00100010110000 : 14'b01100010110000;
											assign node2689 = (inp[4]) ? node2693 : node2690;
												assign node2690 = (inp[5]) ? 14'b01100010010000 : 14'b00000010010000;
												assign node2693 = (inp[5]) ? 14'b00100010010000 : 14'b00100010010100;
										assign node2696 = (inp[9]) ? node2704 : node2697;
											assign node2697 = (inp[5]) ? node2701 : node2698;
												assign node2698 = (inp[4]) ? 14'b00100000110100 : 14'b00000000110000;
												assign node2701 = (inp[4]) ? 14'b00100000110000 : 14'b01100000110000;
											assign node2704 = (inp[5]) ? node2706 : 14'b00000000010000;
												assign node2706 = (inp[4]) ? 14'b00100000010000 : 14'b01100000010000;
									assign node2709 = (inp[5]) ? 14'b00000000000001 : node2710;
										assign node2710 = (inp[4]) ? node2716 : node2711;
											assign node2711 = (inp[6]) ? node2713 : 14'b01000010110100;
												assign node2713 = (inp[9]) ? 14'b01000000010100 : 14'b01000000110100;
											assign node2716 = (inp[6]) ? node2720 : node2717;
												assign node2717 = (inp[9]) ? 14'b00000010010100 : 14'b00000010110100;
												assign node2720 = (inp[9]) ? 14'b00000000010100 : 14'b00000000110100;
								assign node2724 = (inp[4]) ? 14'b00000000000001 : node2725;
									assign node2725 = (inp[5]) ? 14'b00000000000001 : node2726;
										assign node2726 = (inp[12]) ? node2732 : node2727;
											assign node2727 = (inp[6]) ? node2729 : 14'b01100010110100;
												assign node2729 = (inp[9]) ? 14'b01100000010100 : 14'b01100000110100;
											assign node2732 = (inp[6]) ? 14'b01000000010000 : node2733;
												assign node2733 = (inp[9]) ? 14'b01000010010000 : 14'b01000010110000;
							assign node2739 = (inp[6]) ? node2741 : 14'b00000000000001;
								assign node2741 = (inp[9]) ? 14'b00000000000001 : node2742;
									assign node2742 = (inp[5]) ? node2756 : node2743;
										assign node2743 = (inp[4]) ? node2751 : node2744;
											assign node2744 = (inp[2]) ? node2748 : node2745;
												assign node2745 = (inp[12]) ? 14'b01000000100100 : 14'b00000000100000;
												assign node2748 = (inp[12]) ? 14'b01000000100000 : 14'b01100000100100;
											assign node2751 = (inp[2]) ? 14'b00000000000001 : node2752;
												assign node2752 = (inp[12]) ? 14'b00000000100100 : 14'b00100000100100;
										assign node2756 = (inp[12]) ? 14'b00000000000001 : node2757;
											assign node2757 = (inp[2]) ? 14'b00000000000001 : node2758;
												assign node2758 = (inp[4]) ? 14'b00100000100000 : 14'b01100000100000;
						assign node2764 = (inp[12]) ? node2766 : 14'b00000000000001;
							assign node2766 = (inp[3]) ? node2768 : 14'b00000000000001;
								assign node2768 = (inp[5]) ? node2770 : 14'b00000000000001;
									assign node2770 = (inp[9]) ? node2772 : 14'b00000000000001;
										assign node2772 = (inp[2]) ? node2774 : 14'b00000000000001;
											assign node2774 = (inp[4]) ? 14'b10001001001010 : node2775;
												assign node2775 = (inp[6]) ? 14'b10001001000000 : 14'b10001000000000;

endmodule