module dtc_split75_bm65 (
	input  wire [16-1:0] inp,
	output wire [4-1:0] outp
);

	wire [4-1:0] node1;
	wire [4-1:0] node2;
	wire [4-1:0] node3;
	wire [4-1:0] node4;
	wire [4-1:0] node5;
	wire [4-1:0] node6;
	wire [4-1:0] node7;
	wire [4-1:0] node8;
	wire [4-1:0] node9;
	wire [4-1:0] node10;
	wire [4-1:0] node11;
	wire [4-1:0] node13;
	wire [4-1:0] node14;
	wire [4-1:0] node18;
	wire [4-1:0] node20;
	wire [4-1:0] node23;
	wire [4-1:0] node24;
	wire [4-1:0] node25;
	wire [4-1:0] node26;
	wire [4-1:0] node28;
	wire [4-1:0] node31;
	wire [4-1:0] node33;
	wire [4-1:0] node36;
	wire [4-1:0] node38;
	wire [4-1:0] node41;
	wire [4-1:0] node42;
	wire [4-1:0] node44;
	wire [4-1:0] node45;
	wire [4-1:0] node49;
	wire [4-1:0] node51;
	wire [4-1:0] node54;
	wire [4-1:0] node55;
	wire [4-1:0] node56;
	wire [4-1:0] node57;
	wire [4-1:0] node58;
	wire [4-1:0] node62;
	wire [4-1:0] node64;
	wire [4-1:0] node65;
	wire [4-1:0] node69;
	wire [4-1:0] node71;
	wire [4-1:0] node74;
	wire [4-1:0] node75;
	wire [4-1:0] node76;
	wire [4-1:0] node80;
	wire [4-1:0] node81;
	wire [4-1:0] node83;
	wire [4-1:0] node86;
	wire [4-1:0] node87;
	wire [4-1:0] node91;
	wire [4-1:0] node92;
	wire [4-1:0] node93;
	wire [4-1:0] node94;
	wire [4-1:0] node95;
	wire [4-1:0] node96;
	wire [4-1:0] node97;
	wire [4-1:0] node100;
	wire [4-1:0] node104;
	wire [4-1:0] node105;
	wire [4-1:0] node107;
	wire [4-1:0] node108;
	wire [4-1:0] node112;
	wire [4-1:0] node113;
	wire [4-1:0] node117;
	wire [4-1:0] node118;
	wire [4-1:0] node120;
	wire [4-1:0] node122;
	wire [4-1:0] node125;
	wire [4-1:0] node127;
	wire [4-1:0] node130;
	wire [4-1:0] node131;
	wire [4-1:0] node132;
	wire [4-1:0] node134;
	wire [4-1:0] node137;
	wire [4-1:0] node138;
	wire [4-1:0] node141;
	wire [4-1:0] node144;
	wire [4-1:0] node145;
	wire [4-1:0] node146;
	wire [4-1:0] node147;
	wire [4-1:0] node151;
	wire [4-1:0] node153;
	wire [4-1:0] node156;
	wire [4-1:0] node157;
	wire [4-1:0] node161;
	wire [4-1:0] node162;
	wire [4-1:0] node163;
	wire [4-1:0] node164;
	wire [4-1:0] node165;
	wire [4-1:0] node167;
	wire [4-1:0] node171;
	wire [4-1:0] node172;
	wire [4-1:0] node176;
	wire [4-1:0] node177;
	wire [4-1:0] node178;
	wire [4-1:0] node180;
	wire [4-1:0] node181;
	wire [4-1:0] node185;
	wire [4-1:0] node186;
	wire [4-1:0] node190;
	wire [4-1:0] node191;
	wire [4-1:0] node194;
	wire [4-1:0] node195;
	wire [4-1:0] node196;
	wire [4-1:0] node200;
	wire [4-1:0] node203;
	wire [4-1:0] node204;
	wire [4-1:0] node205;
	wire [4-1:0] node206;
	wire [4-1:0] node208;
	wire [4-1:0] node209;
	wire [4-1:0] node213;
	wire [4-1:0] node216;
	wire [4-1:0] node217;
	wire [4-1:0] node218;
	wire [4-1:0] node220;
	wire [4-1:0] node224;
	wire [4-1:0] node226;
	wire [4-1:0] node229;
	wire [4-1:0] node230;
	wire [4-1:0] node232;
	wire [4-1:0] node233;
	wire [4-1:0] node237;
	wire [4-1:0] node238;
	wire [4-1:0] node242;
	wire [4-1:0] node243;
	wire [4-1:0] node244;
	wire [4-1:0] node245;
	wire [4-1:0] node246;
	wire [4-1:0] node247;
	wire [4-1:0] node248;
	wire [4-1:0] node252;
	wire [4-1:0] node253;
	wire [4-1:0] node257;
	wire [4-1:0] node258;
	wire [4-1:0] node259;
	wire [4-1:0] node261;
	wire [4-1:0] node264;
	wire [4-1:0] node265;
	wire [4-1:0] node269;
	wire [4-1:0] node270;
	wire [4-1:0] node274;
	wire [4-1:0] node275;
	wire [4-1:0] node277;
	wire [4-1:0] node278;
	wire [4-1:0] node282;
	wire [4-1:0] node283;
	wire [4-1:0] node287;
	wire [4-1:0] node288;
	wire [4-1:0] node289;
	wire [4-1:0] node290;
	wire [4-1:0] node292;
	wire [4-1:0] node295;
	wire [4-1:0] node297;
	wire [4-1:0] node298;
	wire [4-1:0] node302;
	wire [4-1:0] node304;
	wire [4-1:0] node307;
	wire [4-1:0] node308;
	wire [4-1:0] node309;
	wire [4-1:0] node311;
	wire [4-1:0] node314;
	wire [4-1:0] node315;
	wire [4-1:0] node319;
	wire [4-1:0] node320;
	wire [4-1:0] node324;
	wire [4-1:0] node325;
	wire [4-1:0] node326;
	wire [4-1:0] node327;
	wire [4-1:0] node328;
	wire [4-1:0] node330;
	wire [4-1:0] node332;
	wire [4-1:0] node333;
	wire [4-1:0] node337;
	wire [4-1:0] node338;
	wire [4-1:0] node339;
	wire [4-1:0] node340;
	wire [4-1:0] node344;
	wire [4-1:0] node345;
	wire [4-1:0] node349;
	wire [4-1:0] node351;
	wire [4-1:0] node354;
	wire [4-1:0] node355;
	wire [4-1:0] node357;
	wire [4-1:0] node358;
	wire [4-1:0] node362;
	wire [4-1:0] node363;
	wire [4-1:0] node367;
	wire [4-1:0] node368;
	wire [4-1:0] node369;
	wire [4-1:0] node370;
	wire [4-1:0] node372;
	wire [4-1:0] node375;
	wire [4-1:0] node378;
	wire [4-1:0] node380;
	wire [4-1:0] node383;
	wire [4-1:0] node384;
	wire [4-1:0] node385;
	wire [4-1:0] node389;
	wire [4-1:0] node390;
	wire [4-1:0] node391;
	wire [4-1:0] node395;
	wire [4-1:0] node396;
	wire [4-1:0] node400;
	wire [4-1:0] node401;
	wire [4-1:0] node402;
	wire [4-1:0] node403;
	wire [4-1:0] node404;
	wire [4-1:0] node406;
	wire [4-1:0] node407;
	wire [4-1:0] node411;
	wire [4-1:0] node413;
	wire [4-1:0] node416;
	wire [4-1:0] node418;
	wire [4-1:0] node419;
	wire [4-1:0] node421;
	wire [4-1:0] node424;
	wire [4-1:0] node427;
	wire [4-1:0] node428;
	wire [4-1:0] node429;
	wire [4-1:0] node431;
	wire [4-1:0] node433;
	wire [4-1:0] node437;
	wire [4-1:0] node438;
	wire [4-1:0] node442;
	wire [4-1:0] node443;
	wire [4-1:0] node444;
	wire [4-1:0] node446;
	wire [4-1:0] node447;
	wire [4-1:0] node451;
	wire [4-1:0] node452;
	wire [4-1:0] node456;
	wire [4-1:0] node457;
	wire [4-1:0] node459;
	wire [4-1:0] node460;
	wire [4-1:0] node463;
	wire [4-1:0] node466;
	wire [4-1:0] node467;
	wire [4-1:0] node469;
	wire [4-1:0] node472;
	wire [4-1:0] node475;
	wire [4-1:0] node477;
	wire [4-1:0] node478;
	wire [4-1:0] node479;
	wire [4-1:0] node480;
	wire [4-1:0] node481;
	wire [4-1:0] node482;
	wire [4-1:0] node483;
	wire [4-1:0] node484;
	wire [4-1:0] node487;
	wire [4-1:0] node491;
	wire [4-1:0] node492;
	wire [4-1:0] node493;
	wire [4-1:0] node497;
	wire [4-1:0] node498;
	wire [4-1:0] node502;
	wire [4-1:0] node503;
	wire [4-1:0] node504;
	wire [4-1:0] node506;
	wire [4-1:0] node509;
	wire [4-1:0] node511;
	wire [4-1:0] node513;
	wire [4-1:0] node516;
	wire [4-1:0] node517;
	wire [4-1:0] node520;
	wire [4-1:0] node521;
	wire [4-1:0] node526;
	wire [4-1:0] node527;
	wire [4-1:0] node528;
	wire [4-1:0] node529;
	wire [4-1:0] node530;
	wire [4-1:0] node533;
	wire [4-1:0] node534;
	wire [4-1:0] node535;
	wire [4-1:0] node539;
	wire [4-1:0] node542;
	wire [4-1:0] node543;
	wire [4-1:0] node544;
	wire [4-1:0] node547;
	wire [4-1:0] node550;
	wire [4-1:0] node552;
	wire [4-1:0] node555;
	wire [4-1:0] node556;
	wire [4-1:0] node558;
	wire [4-1:0] node559;
	wire [4-1:0] node563;
	wire [4-1:0] node564;
	wire [4-1:0] node568;
	wire [4-1:0] node569;
	wire [4-1:0] node570;
	wire [4-1:0] node571;
	wire [4-1:0] node574;
	wire [4-1:0] node577;
	wire [4-1:0] node579;
	wire [4-1:0] node582;
	wire [4-1:0] node583;
	wire [4-1:0] node585;
	wire [4-1:0] node587;
	wire [4-1:0] node590;
	wire [4-1:0] node591;
	wire [4-1:0] node595;
	wire [4-1:0] node596;
	wire [4-1:0] node597;
	wire [4-1:0] node598;
	wire [4-1:0] node599;
	wire [4-1:0] node600;
	wire [4-1:0] node601;
	wire [4-1:0] node602;
	wire [4-1:0] node605;
	wire [4-1:0] node609;
	wire [4-1:0] node610;
	wire [4-1:0] node612;
	wire [4-1:0] node616;
	wire [4-1:0] node617;
	wire [4-1:0] node620;
	wire [4-1:0] node621;
	wire [4-1:0] node625;
	wire [4-1:0] node626;
	wire [4-1:0] node627;
	wire [4-1:0] node629;
	wire [4-1:0] node632;
	wire [4-1:0] node633;
	wire [4-1:0] node636;
	wire [4-1:0] node639;
	wire [4-1:0] node640;
	wire [4-1:0] node641;
	wire [4-1:0] node645;
	wire [4-1:0] node647;
	wire [4-1:0] node650;
	wire [4-1:0] node651;
	wire [4-1:0] node652;
	wire [4-1:0] node653;
	wire [4-1:0] node655;
	wire [4-1:0] node656;
	wire [4-1:0] node660;
	wire [4-1:0] node661;
	wire [4-1:0] node662;
	wire [4-1:0] node667;
	wire [4-1:0] node668;
	wire [4-1:0] node670;
	wire [4-1:0] node673;
	wire [4-1:0] node676;
	wire [4-1:0] node677;
	wire [4-1:0] node678;
	wire [4-1:0] node679;
	wire [4-1:0] node683;
	wire [4-1:0] node684;
	wire [4-1:0] node688;
	wire [4-1:0] node689;
	wire [4-1:0] node690;
	wire [4-1:0] node692;
	wire [4-1:0] node695;
	wire [4-1:0] node696;
	wire [4-1:0] node700;
	wire [4-1:0] node701;
	wire [4-1:0] node705;
	wire [4-1:0] node706;
	wire [4-1:0] node707;
	wire [4-1:0] node708;
	wire [4-1:0] node709;
	wire [4-1:0] node710;
	wire [4-1:0] node711;
	wire [4-1:0] node716;
	wire [4-1:0] node717;
	wire [4-1:0] node721;
	wire [4-1:0] node722;
	wire [4-1:0] node723;
	wire [4-1:0] node726;
	wire [4-1:0] node729;
	wire [4-1:0] node731;
	wire [4-1:0] node734;
	wire [4-1:0] node735;
	wire [4-1:0] node736;
	wire [4-1:0] node738;
	wire [4-1:0] node742;
	wire [4-1:0] node743;
	wire [4-1:0] node747;
	wire [4-1:0] node748;
	wire [4-1:0] node749;
	wire [4-1:0] node750;
	wire [4-1:0] node751;
	wire [4-1:0] node755;
	wire [4-1:0] node757;
	wire [4-1:0] node759;
	wire [4-1:0] node763;
	wire [4-1:0] node764;
	wire [4-1:0] node765;
	wire [4-1:0] node769;
	wire [4-1:0] node771;
	wire [4-1:0] node775;
	wire [4-1:0] node776;
	wire [4-1:0] node777;
	wire [4-1:0] node778;
	wire [4-1:0] node779;
	wire [4-1:0] node780;
	wire [4-1:0] node781;
	wire [4-1:0] node782;
	wire [4-1:0] node783;
	wire [4-1:0] node785;
	wire [4-1:0] node786;
	wire [4-1:0] node789;
	wire [4-1:0] node790;
	wire [4-1:0] node793;
	wire [4-1:0] node797;
	wire [4-1:0] node798;
	wire [4-1:0] node799;
	wire [4-1:0] node801;
	wire [4-1:0] node804;
	wire [4-1:0] node805;
	wire [4-1:0] node806;
	wire [4-1:0] node810;
	wire [4-1:0] node811;
	wire [4-1:0] node814;
	wire [4-1:0] node817;
	wire [4-1:0] node819;
	wire [4-1:0] node820;
	wire [4-1:0] node821;
	wire [4-1:0] node826;
	wire [4-1:0] node827;
	wire [4-1:0] node828;
	wire [4-1:0] node829;
	wire [4-1:0] node831;
	wire [4-1:0] node834;
	wire [4-1:0] node835;
	wire [4-1:0] node836;
	wire [4-1:0] node841;
	wire [4-1:0] node842;
	wire [4-1:0] node843;
	wire [4-1:0] node846;
	wire [4-1:0] node849;
	wire [4-1:0] node850;
	wire [4-1:0] node853;
	wire [4-1:0] node854;
	wire [4-1:0] node858;
	wire [4-1:0] node859;
	wire [4-1:0] node861;
	wire [4-1:0] node862;
	wire [4-1:0] node863;
	wire [4-1:0] node866;
	wire [4-1:0] node869;
	wire [4-1:0] node870;
	wire [4-1:0] node873;
	wire [4-1:0] node876;
	wire [4-1:0] node877;
	wire [4-1:0] node878;
	wire [4-1:0] node881;
	wire [4-1:0] node885;
	wire [4-1:0] node886;
	wire [4-1:0] node887;
	wire [4-1:0] node888;
	wire [4-1:0] node889;
	wire [4-1:0] node893;
	wire [4-1:0] node894;
	wire [4-1:0] node895;
	wire [4-1:0] node897;
	wire [4-1:0] node900;
	wire [4-1:0] node901;
	wire [4-1:0] node905;
	wire [4-1:0] node906;
	wire [4-1:0] node907;
	wire [4-1:0] node911;
	wire [4-1:0] node912;
	wire [4-1:0] node916;
	wire [4-1:0] node917;
	wire [4-1:0] node918;
	wire [4-1:0] node919;
	wire [4-1:0] node920;
	wire [4-1:0] node923;
	wire [4-1:0] node926;
	wire [4-1:0] node927;
	wire [4-1:0] node931;
	wire [4-1:0] node932;
	wire [4-1:0] node935;
	wire [4-1:0] node937;
	wire [4-1:0] node940;
	wire [4-1:0] node941;
	wire [4-1:0] node944;
	wire [4-1:0] node946;
	wire [4-1:0] node949;
	wire [4-1:0] node950;
	wire [4-1:0] node951;
	wire [4-1:0] node952;
	wire [4-1:0] node953;
	wire [4-1:0] node956;
	wire [4-1:0] node957;
	wire [4-1:0] node961;
	wire [4-1:0] node962;
	wire [4-1:0] node963;
	wire [4-1:0] node968;
	wire [4-1:0] node969;
	wire [4-1:0] node971;
	wire [4-1:0] node974;
	wire [4-1:0] node977;
	wire [4-1:0] node978;
	wire [4-1:0] node979;
	wire [4-1:0] node980;
	wire [4-1:0] node983;
	wire [4-1:0] node985;
	wire [4-1:0] node989;
	wire [4-1:0] node990;
	wire [4-1:0] node991;
	wire [4-1:0] node992;
	wire [4-1:0] node996;
	wire [4-1:0] node999;
	wire [4-1:0] node1000;
	wire [4-1:0] node1004;
	wire [4-1:0] node1005;
	wire [4-1:0] node1006;
	wire [4-1:0] node1007;
	wire [4-1:0] node1008;
	wire [4-1:0] node1009;
	wire [4-1:0] node1010;
	wire [4-1:0] node1014;
	wire [4-1:0] node1016;
	wire [4-1:0] node1019;
	wire [4-1:0] node1020;
	wire [4-1:0] node1022;
	wire [4-1:0] node1025;
	wire [4-1:0] node1026;
	wire [4-1:0] node1027;
	wire [4-1:0] node1032;
	wire [4-1:0] node1033;
	wire [4-1:0] node1035;
	wire [4-1:0] node1036;
	wire [4-1:0] node1039;
	wire [4-1:0] node1042;
	wire [4-1:0] node1043;
	wire [4-1:0] node1045;
	wire [4-1:0] node1046;
	wire [4-1:0] node1051;
	wire [4-1:0] node1052;
	wire [4-1:0] node1053;
	wire [4-1:0] node1054;
	wire [4-1:0] node1056;
	wire [4-1:0] node1059;
	wire [4-1:0] node1062;
	wire [4-1:0] node1063;
	wire [4-1:0] node1064;
	wire [4-1:0] node1068;
	wire [4-1:0] node1069;
	wire [4-1:0] node1071;
	wire [4-1:0] node1074;
	wire [4-1:0] node1077;
	wire [4-1:0] node1078;
	wire [4-1:0] node1079;
	wire [4-1:0] node1080;
	wire [4-1:0] node1084;
	wire [4-1:0] node1085;
	wire [4-1:0] node1089;
	wire [4-1:0] node1091;
	wire [4-1:0] node1092;
	wire [4-1:0] node1096;
	wire [4-1:0] node1097;
	wire [4-1:0] node1098;
	wire [4-1:0] node1099;
	wire [4-1:0] node1100;
	wire [4-1:0] node1102;
	wire [4-1:0] node1105;
	wire [4-1:0] node1106;
	wire [4-1:0] node1109;
	wire [4-1:0] node1110;
	wire [4-1:0] node1114;
	wire [4-1:0] node1115;
	wire [4-1:0] node1116;
	wire [4-1:0] node1119;
	wire [4-1:0] node1122;
	wire [4-1:0] node1123;
	wire [4-1:0] node1127;
	wire [4-1:0] node1128;
	wire [4-1:0] node1129;
	wire [4-1:0] node1130;
	wire [4-1:0] node1134;
	wire [4-1:0] node1135;
	wire [4-1:0] node1136;
	wire [4-1:0] node1139;
	wire [4-1:0] node1142;
	wire [4-1:0] node1145;
	wire [4-1:0] node1146;
	wire [4-1:0] node1147;
	wire [4-1:0] node1150;
	wire [4-1:0] node1153;
	wire [4-1:0] node1155;
	wire [4-1:0] node1158;
	wire [4-1:0] node1159;
	wire [4-1:0] node1160;
	wire [4-1:0] node1161;
	wire [4-1:0] node1165;
	wire [4-1:0] node1166;
	wire [4-1:0] node1167;
	wire [4-1:0] node1170;
	wire [4-1:0] node1171;
	wire [4-1:0] node1175;
	wire [4-1:0] node1176;
	wire [4-1:0] node1177;
	wire [4-1:0] node1180;
	wire [4-1:0] node1183;
	wire [4-1:0] node1184;
	wire [4-1:0] node1188;
	wire [4-1:0] node1189;
	wire [4-1:0] node1190;
	wire [4-1:0] node1192;
	wire [4-1:0] node1196;
	wire [4-1:0] node1197;
	wire [4-1:0] node1198;
	wire [4-1:0] node1202;
	wire [4-1:0] node1203;
	wire [4-1:0] node1207;
	wire [4-1:0] node1208;
	wire [4-1:0] node1209;
	wire [4-1:0] node1210;
	wire [4-1:0] node1211;
	wire [4-1:0] node1212;
	wire [4-1:0] node1213;
	wire [4-1:0] node1216;
	wire [4-1:0] node1217;
	wire [4-1:0] node1221;
	wire [4-1:0] node1222;
	wire [4-1:0] node1223;
	wire [4-1:0] node1227;
	wire [4-1:0] node1228;
	wire [4-1:0] node1231;
	wire [4-1:0] node1234;
	wire [4-1:0] node1235;
	wire [4-1:0] node1236;
	wire [4-1:0] node1237;
	wire [4-1:0] node1241;
	wire [4-1:0] node1242;
	wire [4-1:0] node1245;
	wire [4-1:0] node1248;
	wire [4-1:0] node1249;
	wire [4-1:0] node1250;
	wire [4-1:0] node1254;
	wire [4-1:0] node1255;
	wire [4-1:0] node1258;
	wire [4-1:0] node1261;
	wire [4-1:0] node1262;
	wire [4-1:0] node1263;
	wire [4-1:0] node1264;
	wire [4-1:0] node1265;
	wire [4-1:0] node1268;
	wire [4-1:0] node1271;
	wire [4-1:0] node1272;
	wire [4-1:0] node1275;
	wire [4-1:0] node1278;
	wire [4-1:0] node1279;
	wire [4-1:0] node1281;
	wire [4-1:0] node1284;
	wire [4-1:0] node1285;
	wire [4-1:0] node1288;
	wire [4-1:0] node1291;
	wire [4-1:0] node1292;
	wire [4-1:0] node1293;
	wire [4-1:0] node1294;
	wire [4-1:0] node1298;
	wire [4-1:0] node1301;
	wire [4-1:0] node1302;
	wire [4-1:0] node1305;
	wire [4-1:0] node1308;
	wire [4-1:0] node1309;
	wire [4-1:0] node1310;
	wire [4-1:0] node1311;
	wire [4-1:0] node1312;
	wire [4-1:0] node1316;
	wire [4-1:0] node1317;
	wire [4-1:0] node1321;
	wire [4-1:0] node1322;
	wire [4-1:0] node1324;
	wire [4-1:0] node1325;
	wire [4-1:0] node1326;
	wire [4-1:0] node1329;
	wire [4-1:0] node1333;
	wire [4-1:0] node1334;
	wire [4-1:0] node1335;
	wire [4-1:0] node1339;
	wire [4-1:0] node1342;
	wire [4-1:0] node1343;
	wire [4-1:0] node1344;
	wire [4-1:0] node1345;
	wire [4-1:0] node1346;
	wire [4-1:0] node1347;
	wire [4-1:0] node1350;
	wire [4-1:0] node1354;
	wire [4-1:0] node1355;
	wire [4-1:0] node1358;
	wire [4-1:0] node1361;
	wire [4-1:0] node1362;
	wire [4-1:0] node1363;
	wire [4-1:0] node1367;
	wire [4-1:0] node1368;
	wire [4-1:0] node1371;
	wire [4-1:0] node1374;
	wire [4-1:0] node1375;
	wire [4-1:0] node1376;
	wire [4-1:0] node1377;
	wire [4-1:0] node1380;
	wire [4-1:0] node1383;
	wire [4-1:0] node1384;
	wire [4-1:0] node1385;
	wire [4-1:0] node1388;
	wire [4-1:0] node1392;
	wire [4-1:0] node1393;
	wire [4-1:0] node1394;
	wire [4-1:0] node1397;
	wire [4-1:0] node1400;
	wire [4-1:0] node1401;
	wire [4-1:0] node1404;
	wire [4-1:0] node1407;
	wire [4-1:0] node1408;
	wire [4-1:0] node1409;
	wire [4-1:0] node1410;
	wire [4-1:0] node1411;
	wire [4-1:0] node1413;
	wire [4-1:0] node1415;
	wire [4-1:0] node1419;
	wire [4-1:0] node1420;
	wire [4-1:0] node1421;
	wire [4-1:0] node1424;
	wire [4-1:0] node1426;
	wire [4-1:0] node1429;
	wire [4-1:0] node1430;
	wire [4-1:0] node1433;
	wire [4-1:0] node1434;
	wire [4-1:0] node1438;
	wire [4-1:0] node1439;
	wire [4-1:0] node1440;
	wire [4-1:0] node1441;
	wire [4-1:0] node1444;
	wire [4-1:0] node1445;
	wire [4-1:0] node1449;
	wire [4-1:0] node1450;
	wire [4-1:0] node1451;
	wire [4-1:0] node1455;
	wire [4-1:0] node1456;
	wire [4-1:0] node1460;
	wire [4-1:0] node1461;
	wire [4-1:0] node1463;
	wire [4-1:0] node1465;
	wire [4-1:0] node1468;
	wire [4-1:0] node1469;
	wire [4-1:0] node1473;
	wire [4-1:0] node1474;
	wire [4-1:0] node1475;
	wire [4-1:0] node1476;
	wire [4-1:0] node1477;
	wire [4-1:0] node1479;
	wire [4-1:0] node1482;
	wire [4-1:0] node1483;
	wire [4-1:0] node1486;
	wire [4-1:0] node1489;
	wire [4-1:0] node1490;
	wire [4-1:0] node1491;
	wire [4-1:0] node1494;
	wire [4-1:0] node1497;
	wire [4-1:0] node1498;
	wire [4-1:0] node1501;
	wire [4-1:0] node1504;
	wire [4-1:0] node1505;
	wire [4-1:0] node1506;
	wire [4-1:0] node1510;
	wire [4-1:0] node1511;
	wire [4-1:0] node1514;
	wire [4-1:0] node1517;
	wire [4-1:0] node1518;
	wire [4-1:0] node1519;
	wire [4-1:0] node1521;
	wire [4-1:0] node1525;
	wire [4-1:0] node1527;
	wire [4-1:0] node1530;
	wire [4-1:0] node1531;
	wire [4-1:0] node1532;
	wire [4-1:0] node1533;
	wire [4-1:0] node1534;
	wire [4-1:0] node1535;
	wire [4-1:0] node1536;
	wire [4-1:0] node1537;
	wire [4-1:0] node1540;
	wire [4-1:0] node1542;
	wire [4-1:0] node1546;
	wire [4-1:0] node1547;
	wire [4-1:0] node1548;
	wire [4-1:0] node1549;
	wire [4-1:0] node1550;
	wire [4-1:0] node1556;
	wire [4-1:0] node1557;
	wire [4-1:0] node1561;
	wire [4-1:0] node1562;
	wire [4-1:0] node1563;
	wire [4-1:0] node1564;
	wire [4-1:0] node1566;
	wire [4-1:0] node1569;
	wire [4-1:0] node1571;
	wire [4-1:0] node1574;
	wire [4-1:0] node1575;
	wire [4-1:0] node1579;
	wire [4-1:0] node1580;
	wire [4-1:0] node1581;
	wire [4-1:0] node1583;
	wire [4-1:0] node1586;
	wire [4-1:0] node1588;
	wire [4-1:0] node1591;
	wire [4-1:0] node1593;
	wire [4-1:0] node1596;
	wire [4-1:0] node1597;
	wire [4-1:0] node1598;
	wire [4-1:0] node1599;
	wire [4-1:0] node1600;
	wire [4-1:0] node1601;
	wire [4-1:0] node1603;
	wire [4-1:0] node1608;
	wire [4-1:0] node1609;
	wire [4-1:0] node1610;
	wire [4-1:0] node1613;
	wire [4-1:0] node1614;
	wire [4-1:0] node1618;
	wire [4-1:0] node1619;
	wire [4-1:0] node1623;
	wire [4-1:0] node1624;
	wire [4-1:0] node1626;
	wire [4-1:0] node1628;
	wire [4-1:0] node1631;
	wire [4-1:0] node1632;
	wire [4-1:0] node1633;
	wire [4-1:0] node1635;
	wire [4-1:0] node1639;
	wire [4-1:0] node1640;
	wire [4-1:0] node1642;
	wire [4-1:0] node1645;
	wire [4-1:0] node1648;
	wire [4-1:0] node1649;
	wire [4-1:0] node1650;
	wire [4-1:0] node1651;
	wire [4-1:0] node1652;
	wire [4-1:0] node1653;
	wire [4-1:0] node1659;
	wire [4-1:0] node1661;
	wire [4-1:0] node1663;
	wire [4-1:0] node1666;
	wire [4-1:0] node1667;
	wire [4-1:0] node1668;
	wire [4-1:0] node1670;
	wire [4-1:0] node1673;
	wire [4-1:0] node1675;
	wire [4-1:0] node1678;
	wire [4-1:0] node1679;
	wire [4-1:0] node1680;
	wire [4-1:0] node1682;
	wire [4-1:0] node1685;
	wire [4-1:0] node1688;
	wire [4-1:0] node1690;
	wire [4-1:0] node1692;
	wire [4-1:0] node1695;
	wire [4-1:0] node1696;
	wire [4-1:0] node1697;
	wire [4-1:0] node1698;
	wire [4-1:0] node1699;
	wire [4-1:0] node1700;
	wire [4-1:0] node1704;
	wire [4-1:0] node1706;
	wire [4-1:0] node1707;
	wire [4-1:0] node1711;
	wire [4-1:0] node1712;
	wire [4-1:0] node1713;
	wire [4-1:0] node1714;
	wire [4-1:0] node1719;
	wire [4-1:0] node1720;
	wire [4-1:0] node1724;
	wire [4-1:0] node1725;
	wire [4-1:0] node1726;
	wire [4-1:0] node1728;
	wire [4-1:0] node1729;
	wire [4-1:0] node1731;
	wire [4-1:0] node1735;
	wire [4-1:0] node1736;
	wire [4-1:0] node1737;
	wire [4-1:0] node1741;
	wire [4-1:0] node1743;
	wire [4-1:0] node1746;
	wire [4-1:0] node1747;
	wire [4-1:0] node1748;
	wire [4-1:0] node1751;
	wire [4-1:0] node1753;
	wire [4-1:0] node1756;
	wire [4-1:0] node1757;
	wire [4-1:0] node1759;
	wire [4-1:0] node1762;
	wire [4-1:0] node1763;
	wire [4-1:0] node1767;
	wire [4-1:0] node1768;
	wire [4-1:0] node1769;
	wire [4-1:0] node1770;
	wire [4-1:0] node1771;
	wire [4-1:0] node1773;
	wire [4-1:0] node1776;
	wire [4-1:0] node1777;
	wire [4-1:0] node1782;
	wire [4-1:0] node1783;
	wire [4-1:0] node1784;
	wire [4-1:0] node1785;
	wire [4-1:0] node1789;
	wire [4-1:0] node1791;
	wire [4-1:0] node1794;
	wire [4-1:0] node1795;
	wire [4-1:0] node1799;
	wire [4-1:0] node1800;
	wire [4-1:0] node1801;
	wire [4-1:0] node1803;
	wire [4-1:0] node1806;
	wire [4-1:0] node1807;
	wire [4-1:0] node1808;
	wire [4-1:0] node1812;
	wire [4-1:0] node1813;
	wire [4-1:0] node1817;
	wire [4-1:0] node1818;
	wire [4-1:0] node1819;
	wire [4-1:0] node1820;
	wire [4-1:0] node1824;
	wire [4-1:0] node1826;
	wire [4-1:0] node1827;
	wire [4-1:0] node1831;
	wire [4-1:0] node1832;
	wire [4-1:0] node1835;
	wire [4-1:0] node1837;
	wire [4-1:0] node1841;
	wire [4-1:0] node1842;
	wire [4-1:0] node1843;
	wire [4-1:0] node1844;
	wire [4-1:0] node1845;
	wire [4-1:0] node1846;
	wire [4-1:0] node1847;
	wire [4-1:0] node1848;
	wire [4-1:0] node1849;
	wire [4-1:0] node1852;
	wire [4-1:0] node1853;
	wire [4-1:0] node1854;
	wire [4-1:0] node1858;
	wire [4-1:0] node1861;
	wire [4-1:0] node1862;
	wire [4-1:0] node1863;
	wire [4-1:0] node1865;
	wire [4-1:0] node1868;
	wire [4-1:0] node1871;
	wire [4-1:0] node1872;
	wire [4-1:0] node1875;
	wire [4-1:0] node1878;
	wire [4-1:0] node1879;
	wire [4-1:0] node1880;
	wire [4-1:0] node1883;
	wire [4-1:0] node1886;
	wire [4-1:0] node1887;
	wire [4-1:0] node1888;
	wire [4-1:0] node1891;
	wire [4-1:0] node1894;
	wire [4-1:0] node1895;
	wire [4-1:0] node1897;
	wire [4-1:0] node1900;
	wire [4-1:0] node1901;
	wire [4-1:0] node1904;
	wire [4-1:0] node1907;
	wire [4-1:0] node1908;
	wire [4-1:0] node1909;
	wire [4-1:0] node1910;
	wire [4-1:0] node1911;
	wire [4-1:0] node1912;
	wire [4-1:0] node1916;
	wire [4-1:0] node1918;
	wire [4-1:0] node1921;
	wire [4-1:0] node1922;
	wire [4-1:0] node1924;
	wire [4-1:0] node1928;
	wire [4-1:0] node1929;
	wire [4-1:0] node1930;
	wire [4-1:0] node1933;
	wire [4-1:0] node1934;
	wire [4-1:0] node1937;
	wire [4-1:0] node1940;
	wire [4-1:0] node1941;
	wire [4-1:0] node1942;
	wire [4-1:0] node1946;
	wire [4-1:0] node1949;
	wire [4-1:0] node1950;
	wire [4-1:0] node1952;
	wire [4-1:0] node1953;
	wire [4-1:0] node1956;
	wire [4-1:0] node1959;
	wire [4-1:0] node1960;
	wire [4-1:0] node1962;
	wire [4-1:0] node1965;
	wire [4-1:0] node1966;
	wire [4-1:0] node1970;
	wire [4-1:0] node1971;
	wire [4-1:0] node1972;
	wire [4-1:0] node1973;
	wire [4-1:0] node1974;
	wire [4-1:0] node1977;
	wire [4-1:0] node1978;
	wire [4-1:0] node1981;
	wire [4-1:0] node1984;
	wire [4-1:0] node1985;
	wire [4-1:0] node1988;
	wire [4-1:0] node1989;
	wire [4-1:0] node1993;
	wire [4-1:0] node1994;
	wire [4-1:0] node1995;
	wire [4-1:0] node1998;
	wire [4-1:0] node2000;
	wire [4-1:0] node2003;
	wire [4-1:0] node2004;
	wire [4-1:0] node2005;
	wire [4-1:0] node2008;
	wire [4-1:0] node2010;
	wire [4-1:0] node2013;
	wire [4-1:0] node2014;
	wire [4-1:0] node2017;
	wire [4-1:0] node2020;
	wire [4-1:0] node2021;
	wire [4-1:0] node2022;
	wire [4-1:0] node2023;
	wire [4-1:0] node2024;
	wire [4-1:0] node2028;
	wire [4-1:0] node2029;
	wire [4-1:0] node2032;
	wire [4-1:0] node2035;
	wire [4-1:0] node2036;
	wire [4-1:0] node2037;
	wire [4-1:0] node2041;
	wire [4-1:0] node2043;
	wire [4-1:0] node2047;
	wire [4-1:0] node2048;
	wire [4-1:0] node2049;
	wire [4-1:0] node2050;
	wire [4-1:0] node2051;
	wire [4-1:0] node2053;
	wire [4-1:0] node2056;
	wire [4-1:0] node2057;
	wire [4-1:0] node2058;
	wire [4-1:0] node2059;
	wire [4-1:0] node2063;
	wire [4-1:0] node2066;
	wire [4-1:0] node2068;
	wire [4-1:0] node2071;
	wire [4-1:0] node2072;
	wire [4-1:0] node2073;
	wire [4-1:0] node2074;
	wire [4-1:0] node2075;
	wire [4-1:0] node2078;
	wire [4-1:0] node2081;
	wire [4-1:0] node2084;
	wire [4-1:0] node2085;
	wire [4-1:0] node2086;
	wire [4-1:0] node2089;
	wire [4-1:0] node2092;
	wire [4-1:0] node2093;
	wire [4-1:0] node2096;
	wire [4-1:0] node2099;
	wire [4-1:0] node2100;
	wire [4-1:0] node2101;
	wire [4-1:0] node2103;
	wire [4-1:0] node2106;
	wire [4-1:0] node2107;
	wire [4-1:0] node2110;
	wire [4-1:0] node2113;
	wire [4-1:0] node2114;
	wire [4-1:0] node2117;
	wire [4-1:0] node2120;
	wire [4-1:0] node2121;
	wire [4-1:0] node2122;
	wire [4-1:0] node2123;
	wire [4-1:0] node2124;
	wire [4-1:0] node2125;
	wire [4-1:0] node2129;
	wire [4-1:0] node2132;
	wire [4-1:0] node2133;
	wire [4-1:0] node2134;
	wire [4-1:0] node2139;
	wire [4-1:0] node2140;
	wire [4-1:0] node2141;
	wire [4-1:0] node2142;
	wire [4-1:0] node2145;
	wire [4-1:0] node2148;
	wire [4-1:0] node2149;
	wire [4-1:0] node2152;
	wire [4-1:0] node2156;
	wire [4-1:0] node2157;
	wire [4-1:0] node2159;
	wire [4-1:0] node2162;
	wire [4-1:0] node2163;
	wire [4-1:0] node2164;
	wire [4-1:0] node2169;
	wire [4-1:0] node2170;
	wire [4-1:0] node2171;
	wire [4-1:0] node2172;
	wire [4-1:0] node2173;
	wire [4-1:0] node2174;
	wire [4-1:0] node2177;
	wire [4-1:0] node2180;
	wire [4-1:0] node2181;
	wire [4-1:0] node2185;
	wire [4-1:0] node2186;
	wire [4-1:0] node2187;
	wire [4-1:0] node2189;
	wire [4-1:0] node2193;
	wire [4-1:0] node2194;
	wire [4-1:0] node2196;
	wire [4-1:0] node2200;
	wire [4-1:0] node2201;
	wire [4-1:0] node2202;
	wire [4-1:0] node2203;
	wire [4-1:0] node2207;
	wire [4-1:0] node2210;
	wire [4-1:0] node2212;
	wire [4-1:0] node2213;
	wire [4-1:0] node2216;
	wire [4-1:0] node2219;
	wire [4-1:0] node2220;
	wire [4-1:0] node2221;
	wire [4-1:0] node2223;
	wire [4-1:0] node2224;
	wire [4-1:0] node2228;
	wire [4-1:0] node2229;
	wire [4-1:0] node2233;
	wire [4-1:0] node2234;
	wire [4-1:0] node2235;
	wire [4-1:0] node2237;
	wire [4-1:0] node2238;
	wire [4-1:0] node2242;
	wire [4-1:0] node2245;
	wire [4-1:0] node2246;
	wire [4-1:0] node2248;
	wire [4-1:0] node2251;
	wire [4-1:0] node2252;
	wire [4-1:0] node2256;
	wire [4-1:0] node2257;
	wire [4-1:0] node2258;
	wire [4-1:0] node2259;
	wire [4-1:0] node2260;
	wire [4-1:0] node2261;
	wire [4-1:0] node2262;
	wire [4-1:0] node2265;
	wire [4-1:0] node2268;
	wire [4-1:0] node2269;
	wire [4-1:0] node2270;
	wire [4-1:0] node2271;
	wire [4-1:0] node2276;
	wire [4-1:0] node2277;
	wire [4-1:0] node2278;
	wire [4-1:0] node2283;
	wire [4-1:0] node2284;
	wire [4-1:0] node2285;
	wire [4-1:0] node2286;
	wire [4-1:0] node2289;
	wire [4-1:0] node2290;
	wire [4-1:0] node2293;
	wire [4-1:0] node2296;
	wire [4-1:0] node2297;
	wire [4-1:0] node2298;
	wire [4-1:0] node2301;
	wire [4-1:0] node2304;
	wire [4-1:0] node2307;
	wire [4-1:0] node2308;
	wire [4-1:0] node2309;
	wire [4-1:0] node2312;
	wire [4-1:0] node2313;
	wire [4-1:0] node2317;
	wire [4-1:0] node2318;
	wire [4-1:0] node2322;
	wire [4-1:0] node2323;
	wire [4-1:0] node2324;
	wire [4-1:0] node2325;
	wire [4-1:0] node2327;
	wire [4-1:0] node2330;
	wire [4-1:0] node2331;
	wire [4-1:0] node2334;
	wire [4-1:0] node2337;
	wire [4-1:0] node2338;
	wire [4-1:0] node2340;
	wire [4-1:0] node2341;
	wire [4-1:0] node2346;
	wire [4-1:0] node2347;
	wire [4-1:0] node2348;
	wire [4-1:0] node2349;
	wire [4-1:0] node2353;
	wire [4-1:0] node2354;
	wire [4-1:0] node2355;
	wire [4-1:0] node2360;
	wire [4-1:0] node2361;
	wire [4-1:0] node2362;
	wire [4-1:0] node2365;
	wire [4-1:0] node2367;
	wire [4-1:0] node2370;
	wire [4-1:0] node2373;
	wire [4-1:0] node2374;
	wire [4-1:0] node2375;
	wire [4-1:0] node2376;
	wire [4-1:0] node2377;
	wire [4-1:0] node2378;
	wire [4-1:0] node2381;
	wire [4-1:0] node2385;
	wire [4-1:0] node2386;
	wire [4-1:0] node2388;
	wire [4-1:0] node2390;
	wire [4-1:0] node2393;
	wire [4-1:0] node2394;
	wire [4-1:0] node2397;
	wire [4-1:0] node2400;
	wire [4-1:0] node2401;
	wire [4-1:0] node2402;
	wire [4-1:0] node2403;
	wire [4-1:0] node2404;
	wire [4-1:0] node2408;
	wire [4-1:0] node2411;
	wire [4-1:0] node2412;
	wire [4-1:0] node2414;
	wire [4-1:0] node2418;
	wire [4-1:0] node2419;
	wire [4-1:0] node2420;
	wire [4-1:0] node2422;
	wire [4-1:0] node2425;
	wire [4-1:0] node2429;
	wire [4-1:0] node2430;
	wire [4-1:0] node2431;
	wire [4-1:0] node2432;
	wire [4-1:0] node2433;
	wire [4-1:0] node2434;
	wire [4-1:0] node2439;
	wire [4-1:0] node2442;
	wire [4-1:0] node2443;
	wire [4-1:0] node2445;
	wire [4-1:0] node2448;
	wire [4-1:0] node2449;
	wire [4-1:0] node2452;
	wire [4-1:0] node2455;
	wire [4-1:0] node2456;
	wire [4-1:0] node2457;
	wire [4-1:0] node2458;
	wire [4-1:0] node2459;
	wire [4-1:0] node2463;
	wire [4-1:0] node2465;
	wire [4-1:0] node2468;
	wire [4-1:0] node2469;
	wire [4-1:0] node2471;
	wire [4-1:0] node2474;
	wire [4-1:0] node2476;
	wire [4-1:0] node2479;
	wire [4-1:0] node2480;
	wire [4-1:0] node2481;
	wire [4-1:0] node2483;
	wire [4-1:0] node2487;
	wire [4-1:0] node2489;
	wire [4-1:0] node2492;
	wire [4-1:0] node2493;
	wire [4-1:0] node2494;
	wire [4-1:0] node2495;
	wire [4-1:0] node2496;
	wire [4-1:0] node2497;
	wire [4-1:0] node2498;
	wire [4-1:0] node2502;
	wire [4-1:0] node2503;
	wire [4-1:0] node2506;
	wire [4-1:0] node2509;
	wire [4-1:0] node2510;
	wire [4-1:0] node2511;
	wire [4-1:0] node2515;
	wire [4-1:0] node2518;
	wire [4-1:0] node2519;
	wire [4-1:0] node2520;
	wire [4-1:0] node2521;
	wire [4-1:0] node2524;
	wire [4-1:0] node2527;
	wire [4-1:0] node2528;
	wire [4-1:0] node2531;
	wire [4-1:0] node2534;
	wire [4-1:0] node2536;
	wire [4-1:0] node2539;
	wire [4-1:0] node2540;
	wire [4-1:0] node2541;
	wire [4-1:0] node2542;
	wire [4-1:0] node2543;
	wire [4-1:0] node2546;
	wire [4-1:0] node2549;
	wire [4-1:0] node2550;
	wire [4-1:0] node2553;
	wire [4-1:0] node2556;
	wire [4-1:0] node2557;
	wire [4-1:0] node2559;
	wire [4-1:0] node2562;
	wire [4-1:0] node2563;
	wire [4-1:0] node2567;
	wire [4-1:0] node2568;
	wire [4-1:0] node2569;
	wire [4-1:0] node2570;
	wire [4-1:0] node2574;
	wire [4-1:0] node2575;
	wire [4-1:0] node2579;
	wire [4-1:0] node2580;
	wire [4-1:0] node2583;
	wire [4-1:0] node2585;
	wire [4-1:0] node2588;
	wire [4-1:0] node2589;
	wire [4-1:0] node2590;
	wire [4-1:0] node2591;
	wire [4-1:0] node2593;
	wire [4-1:0] node2596;
	wire [4-1:0] node2598;
	wire [4-1:0] node2599;
	wire [4-1:0] node2600;
	wire [4-1:0] node2604;
	wire [4-1:0] node2605;
	wire [4-1:0] node2608;
	wire [4-1:0] node2611;
	wire [4-1:0] node2612;
	wire [4-1:0] node2614;
	wire [4-1:0] node2617;
	wire [4-1:0] node2618;
	wire [4-1:0] node2621;
	wire [4-1:0] node2624;
	wire [4-1:0] node2625;
	wire [4-1:0] node2626;
	wire [4-1:0] node2628;
	wire [4-1:0] node2631;
	wire [4-1:0] node2632;
	wire [4-1:0] node2633;
	wire [4-1:0] node2634;
	wire [4-1:0] node2637;
	wire [4-1:0] node2641;
	wire [4-1:0] node2642;
	wire [4-1:0] node2645;
	wire [4-1:0] node2649;
	wire [4-1:0] node2650;
	wire [4-1:0] node2651;
	wire [4-1:0] node2652;
	wire [4-1:0] node2653;
	wire [4-1:0] node2654;
	wire [4-1:0] node2655;
	wire [4-1:0] node2656;
	wire [4-1:0] node2657;
	wire [4-1:0] node2659;
	wire [4-1:0] node2662;
	wire [4-1:0] node2665;
	wire [4-1:0] node2666;
	wire [4-1:0] node2667;
	wire [4-1:0] node2670;
	wire [4-1:0] node2674;
	wire [4-1:0] node2675;
	wire [4-1:0] node2676;
	wire [4-1:0] node2680;
	wire [4-1:0] node2681;
	wire [4-1:0] node2683;
	wire [4-1:0] node2687;
	wire [4-1:0] node2688;
	wire [4-1:0] node2689;
	wire [4-1:0] node2690;
	wire [4-1:0] node2692;
	wire [4-1:0] node2695;
	wire [4-1:0] node2696;
	wire [4-1:0] node2700;
	wire [4-1:0] node2701;
	wire [4-1:0] node2705;
	wire [4-1:0] node2706;
	wire [4-1:0] node2708;
	wire [4-1:0] node2711;
	wire [4-1:0] node2712;
	wire [4-1:0] node2713;
	wire [4-1:0] node2717;
	wire [4-1:0] node2719;
	wire [4-1:0] node2722;
	wire [4-1:0] node2723;
	wire [4-1:0] node2724;
	wire [4-1:0] node2726;
	wire [4-1:0] node2727;
	wire [4-1:0] node2730;
	wire [4-1:0] node2733;
	wire [4-1:0] node2734;
	wire [4-1:0] node2735;
	wire [4-1:0] node2739;
	wire [4-1:0] node2740;
	wire [4-1:0] node2741;
	wire [4-1:0] node2746;
	wire [4-1:0] node2747;
	wire [4-1:0] node2748;
	wire [4-1:0] node2750;
	wire [4-1:0] node2752;
	wire [4-1:0] node2755;
	wire [4-1:0] node2756;
	wire [4-1:0] node2760;
	wire [4-1:0] node2763;
	wire [4-1:0] node2764;
	wire [4-1:0] node2765;
	wire [4-1:0] node2766;
	wire [4-1:0] node2767;
	wire [4-1:0] node2768;
	wire [4-1:0] node2772;
	wire [4-1:0] node2773;
	wire [4-1:0] node2776;
	wire [4-1:0] node2778;
	wire [4-1:0] node2781;
	wire [4-1:0] node2782;
	wire [4-1:0] node2783;
	wire [4-1:0] node2787;
	wire [4-1:0] node2788;
	wire [4-1:0] node2789;
	wire [4-1:0] node2794;
	wire [4-1:0] node2795;
	wire [4-1:0] node2797;
	wire [4-1:0] node2798;
	wire [4-1:0] node2800;
	wire [4-1:0] node2803;
	wire [4-1:0] node2804;
	wire [4-1:0] node2808;
	wire [4-1:0] node2809;
	wire [4-1:0] node2811;
	wire [4-1:0] node2814;
	wire [4-1:0] node2815;
	wire [4-1:0] node2818;
	wire [4-1:0] node2821;
	wire [4-1:0] node2822;
	wire [4-1:0] node2823;
	wire [4-1:0] node2824;
	wire [4-1:0] node2825;
	wire [4-1:0] node2828;
	wire [4-1:0] node2831;
	wire [4-1:0] node2832;
	wire [4-1:0] node2836;
	wire [4-1:0] node2837;
	wire [4-1:0] node2841;
	wire [4-1:0] node2842;
	wire [4-1:0] node2844;
	wire [4-1:0] node2845;
	wire [4-1:0] node2846;
	wire [4-1:0] node2849;
	wire [4-1:0] node2852;
	wire [4-1:0] node2855;
	wire [4-1:0] node2856;
	wire [4-1:0] node2857;
	wire [4-1:0] node2860;
	wire [4-1:0] node2862;
	wire [4-1:0] node2865;
	wire [4-1:0] node2867;
	wire [4-1:0] node2870;
	wire [4-1:0] node2871;
	wire [4-1:0] node2872;
	wire [4-1:0] node2873;
	wire [4-1:0] node2874;
	wire [4-1:0] node2875;
	wire [4-1:0] node2879;
	wire [4-1:0] node2880;
	wire [4-1:0] node2882;
	wire [4-1:0] node2885;
	wire [4-1:0] node2886;
	wire [4-1:0] node2889;
	wire [4-1:0] node2892;
	wire [4-1:0] node2893;
	wire [4-1:0] node2894;
	wire [4-1:0] node2897;
	wire [4-1:0] node2898;
	wire [4-1:0] node2902;
	wire [4-1:0] node2903;
	wire [4-1:0] node2904;
	wire [4-1:0] node2907;
	wire [4-1:0] node2910;
	wire [4-1:0] node2911;
	wire [4-1:0] node2914;
	wire [4-1:0] node2917;
	wire [4-1:0] node2918;
	wire [4-1:0] node2919;
	wire [4-1:0] node2920;
	wire [4-1:0] node2922;
	wire [4-1:0] node2926;
	wire [4-1:0] node2927;
	wire [4-1:0] node2929;
	wire [4-1:0] node2932;
	wire [4-1:0] node2935;
	wire [4-1:0] node2936;
	wire [4-1:0] node2937;
	wire [4-1:0] node2939;
	wire [4-1:0] node2942;
	wire [4-1:0] node2943;
	wire [4-1:0] node2947;
	wire [4-1:0] node2948;
	wire [4-1:0] node2949;
	wire [4-1:0] node2952;
	wire [4-1:0] node2955;
	wire [4-1:0] node2956;
	wire [4-1:0] node2959;
	wire [4-1:0] node2962;
	wire [4-1:0] node2963;
	wire [4-1:0] node2964;
	wire [4-1:0] node2965;
	wire [4-1:0] node2966;
	wire [4-1:0] node2967;
	wire [4-1:0] node2972;
	wire [4-1:0] node2973;
	wire [4-1:0] node2976;
	wire [4-1:0] node2978;
	wire [4-1:0] node2981;
	wire [4-1:0] node2982;
	wire [4-1:0] node2983;
	wire [4-1:0] node2985;
	wire [4-1:0] node2988;
	wire [4-1:0] node2989;
	wire [4-1:0] node2993;
	wire [4-1:0] node2995;
	wire [4-1:0] node2997;
	wire [4-1:0] node2999;
	wire [4-1:0] node3002;
	wire [4-1:0] node3003;
	wire [4-1:0] node3004;
	wire [4-1:0] node3005;
	wire [4-1:0] node3009;
	wire [4-1:0] node3010;
	wire [4-1:0] node3013;
	wire [4-1:0] node3017;
	wire [4-1:0] node3018;
	wire [4-1:0] node3019;
	wire [4-1:0] node3020;
	wire [4-1:0] node3021;
	wire [4-1:0] node3022;
	wire [4-1:0] node3023;
	wire [4-1:0] node3024;
	wire [4-1:0] node3025;
	wire [4-1:0] node3029;
	wire [4-1:0] node3032;
	wire [4-1:0] node3035;
	wire [4-1:0] node3036;
	wire [4-1:0] node3038;
	wire [4-1:0] node3041;
	wire [4-1:0] node3043;
	wire [4-1:0] node3046;
	wire [4-1:0] node3047;
	wire [4-1:0] node3048;
	wire [4-1:0] node3049;
	wire [4-1:0] node3050;
	wire [4-1:0] node3054;
	wire [4-1:0] node3055;
	wire [4-1:0] node3058;
	wire [4-1:0] node3061;
	wire [4-1:0] node3063;
	wire [4-1:0] node3064;
	wire [4-1:0] node3068;
	wire [4-1:0] node3069;
	wire [4-1:0] node3070;
	wire [4-1:0] node3073;
	wire [4-1:0] node3076;
	wire [4-1:0] node3077;
	wire [4-1:0] node3078;
	wire [4-1:0] node3081;
	wire [4-1:0] node3084;
	wire [4-1:0] node3085;
	wire [4-1:0] node3089;
	wire [4-1:0] node3090;
	wire [4-1:0] node3091;
	wire [4-1:0] node3092;
	wire [4-1:0] node3093;
	wire [4-1:0] node3096;
	wire [4-1:0] node3099;
	wire [4-1:0] node3100;
	wire [4-1:0] node3104;
	wire [4-1:0] node3105;
	wire [4-1:0] node3108;
	wire [4-1:0] node3109;
	wire [4-1:0] node3112;
	wire [4-1:0] node3115;
	wire [4-1:0] node3116;
	wire [4-1:0] node3117;
	wire [4-1:0] node3118;
	wire [4-1:0] node3122;
	wire [4-1:0] node3123;
	wire [4-1:0] node3127;
	wire [4-1:0] node3128;
	wire [4-1:0] node3129;
	wire [4-1:0] node3133;
	wire [4-1:0] node3134;
	wire [4-1:0] node3137;
	wire [4-1:0] node3140;
	wire [4-1:0] node3141;
	wire [4-1:0] node3142;
	wire [4-1:0] node3143;
	wire [4-1:0] node3144;
	wire [4-1:0] node3145;
	wire [4-1:0] node3148;
	wire [4-1:0] node3149;
	wire [4-1:0] node3153;
	wire [4-1:0] node3155;
	wire [4-1:0] node3158;
	wire [4-1:0] node3159;
	wire [4-1:0] node3160;
	wire [4-1:0] node3163;
	wire [4-1:0] node3166;
	wire [4-1:0] node3168;
	wire [4-1:0] node3171;
	wire [4-1:0] node3172;
	wire [4-1:0] node3173;
	wire [4-1:0] node3174;
	wire [4-1:0] node3178;
	wire [4-1:0] node3180;
	wire [4-1:0] node3183;
	wire [4-1:0] node3184;
	wire [4-1:0] node3185;
	wire [4-1:0] node3190;
	wire [4-1:0] node3191;
	wire [4-1:0] node3192;
	wire [4-1:0] node3193;
	wire [4-1:0] node3194;
	wire [4-1:0] node3198;
	wire [4-1:0] node3199;
	wire [4-1:0] node3200;
	wire [4-1:0] node3204;
	wire [4-1:0] node3206;
	wire [4-1:0] node3209;
	wire [4-1:0] node3210;
	wire [4-1:0] node3213;
	wire [4-1:0] node3215;
	wire [4-1:0] node3216;
	wire [4-1:0] node3219;
	wire [4-1:0] node3223;
	wire [4-1:0] node3224;
	wire [4-1:0] node3225;
	wire [4-1:0] node3226;
	wire [4-1:0] node3227;
	wire [4-1:0] node3228;
	wire [4-1:0] node3229;
	wire [4-1:0] node3230;
	wire [4-1:0] node3233;
	wire [4-1:0] node3237;
	wire [4-1:0] node3239;
	wire [4-1:0] node3242;
	wire [4-1:0] node3243;
	wire [4-1:0] node3244;
	wire [4-1:0] node3245;
	wire [4-1:0] node3249;
	wire [4-1:0] node3250;
	wire [4-1:0] node3254;
	wire [4-1:0] node3257;
	wire [4-1:0] node3258;
	wire [4-1:0] node3260;
	wire [4-1:0] node3262;
	wire [4-1:0] node3265;
	wire [4-1:0] node3266;
	wire [4-1:0] node3267;
	wire [4-1:0] node3270;
	wire [4-1:0] node3273;
	wire [4-1:0] node3274;
	wire [4-1:0] node3278;
	wire [4-1:0] node3279;
	wire [4-1:0] node3280;
	wire [4-1:0] node3281;
	wire [4-1:0] node3283;
	wire [4-1:0] node3286;
	wire [4-1:0] node3287;
	wire [4-1:0] node3291;
	wire [4-1:0] node3292;
	wire [4-1:0] node3294;
	wire [4-1:0] node3297;
	wire [4-1:0] node3298;
	wire [4-1:0] node3299;
	wire [4-1:0] node3305;
	wire [4-1:0] node3306;
	wire [4-1:0] node3307;
	wire [4-1:0] node3308;
	wire [4-1:0] node3309;
	wire [4-1:0] node3310;
	wire [4-1:0] node3311;
	wire [4-1:0] node3316;
	wire [4-1:0] node3317;
	wire [4-1:0] node3318;
	wire [4-1:0] node3322;
	wire [4-1:0] node3325;
	wire [4-1:0] node3326;
	wire [4-1:0] node3328;
	wire [4-1:0] node3329;
	wire [4-1:0] node3332;
	wire [4-1:0] node3335;
	wire [4-1:0] node3337;
	wire [4-1:0] node3338;
	wire [4-1:0] node3344;
	wire [4-1:0] node3345;
	wire [4-1:0] node3346;
	wire [4-1:0] node3347;
	wire [4-1:0] node3348;
	wire [4-1:0] node3350;
	wire [4-1:0] node3351;
	wire [4-1:0] node3352;
	wire [4-1:0] node3353;
	wire [4-1:0] node3354;
	wire [4-1:0] node3355;
	wire [4-1:0] node3356;
	wire [4-1:0] node3361;
	wire [4-1:0] node3362;
	wire [4-1:0] node3363;
	wire [4-1:0] node3364;
	wire [4-1:0] node3368;
	wire [4-1:0] node3371;
	wire [4-1:0] node3372;
	wire [4-1:0] node3376;
	wire [4-1:0] node3377;
	wire [4-1:0] node3379;
	wire [4-1:0] node3380;
	wire [4-1:0] node3384;
	wire [4-1:0] node3385;
	wire [4-1:0] node3389;
	wire [4-1:0] node3390;
	wire [4-1:0] node3391;
	wire [4-1:0] node3393;
	wire [4-1:0] node3394;
	wire [4-1:0] node3398;
	wire [4-1:0] node3399;
	wire [4-1:0] node3403;
	wire [4-1:0] node3404;
	wire [4-1:0] node3405;
	wire [4-1:0] node3407;
	wire [4-1:0] node3410;
	wire [4-1:0] node3411;
	wire [4-1:0] node3415;
	wire [4-1:0] node3416;
	wire [4-1:0] node3417;
	wire [4-1:0] node3419;
	wire [4-1:0] node3423;
	wire [4-1:0] node3424;
	wire [4-1:0] node3428;
	wire [4-1:0] node3430;
	wire [4-1:0] node3431;
	wire [4-1:0] node3432;
	wire [4-1:0] node3433;
	wire [4-1:0] node3434;
	wire [4-1:0] node3437;
	wire [4-1:0] node3441;
	wire [4-1:0] node3442;
	wire [4-1:0] node3443;
	wire [4-1:0] node3446;
	wire [4-1:0] node3450;
	wire [4-1:0] node3451;
	wire [4-1:0] node3452;
	wire [4-1:0] node3455;
	wire [4-1:0] node3456;
	wire [4-1:0] node3460;
	wire [4-1:0] node3461;
	wire [4-1:0] node3463;
	wire [4-1:0] node3464;
	wire [4-1:0] node3468;
	wire [4-1:0] node3469;
	wire [4-1:0] node3474;
	wire [4-1:0] node3475;
	wire [4-1:0] node3476;
	wire [4-1:0] node3477;
	wire [4-1:0] node3478;
	wire [4-1:0] node3479;
	wire [4-1:0] node3480;
	wire [4-1:0] node3481;
	wire [4-1:0] node3483;
	wire [4-1:0] node3486;
	wire [4-1:0] node3488;
	wire [4-1:0] node3491;
	wire [4-1:0] node3493;
	wire [4-1:0] node3494;
	wire [4-1:0] node3495;
	wire [4-1:0] node3498;
	wire [4-1:0] node3502;
	wire [4-1:0] node3503;
	wire [4-1:0] node3504;
	wire [4-1:0] node3506;
	wire [4-1:0] node3509;
	wire [4-1:0] node3511;
	wire [4-1:0] node3514;
	wire [4-1:0] node3515;
	wire [4-1:0] node3516;
	wire [4-1:0] node3518;
	wire [4-1:0] node3522;
	wire [4-1:0] node3523;
	wire [4-1:0] node3525;
	wire [4-1:0] node3529;
	wire [4-1:0] node3530;
	wire [4-1:0] node3531;
	wire [4-1:0] node3532;
	wire [4-1:0] node3533;
	wire [4-1:0] node3536;
	wire [4-1:0] node3539;
	wire [4-1:0] node3541;
	wire [4-1:0] node3542;
	wire [4-1:0] node3546;
	wire [4-1:0] node3547;
	wire [4-1:0] node3548;
	wire [4-1:0] node3552;
	wire [4-1:0] node3554;
	wire [4-1:0] node3557;
	wire [4-1:0] node3558;
	wire [4-1:0] node3559;
	wire [4-1:0] node3560;
	wire [4-1:0] node3564;
	wire [4-1:0] node3565;
	wire [4-1:0] node3567;
	wire [4-1:0] node3571;
	wire [4-1:0] node3572;
	wire [4-1:0] node3573;
	wire [4-1:0] node3575;
	wire [4-1:0] node3578;
	wire [4-1:0] node3582;
	wire [4-1:0] node3583;
	wire [4-1:0] node3584;
	wire [4-1:0] node3585;
	wire [4-1:0] node3586;
	wire [4-1:0] node3588;
	wire [4-1:0] node3592;
	wire [4-1:0] node3593;
	wire [4-1:0] node3594;
	wire [4-1:0] node3598;
	wire [4-1:0] node3599;
	wire [4-1:0] node3603;
	wire [4-1:0] node3604;
	wire [4-1:0] node3605;
	wire [4-1:0] node3609;
	wire [4-1:0] node3611;
	wire [4-1:0] node3614;
	wire [4-1:0] node3615;
	wire [4-1:0] node3616;
	wire [4-1:0] node3618;
	wire [4-1:0] node3619;
	wire [4-1:0] node3623;
	wire [4-1:0] node3624;
	wire [4-1:0] node3626;
	wire [4-1:0] node3629;
	wire [4-1:0] node3630;
	wire [4-1:0] node3634;
	wire [4-1:0] node3635;
	wire [4-1:0] node3636;
	wire [4-1:0] node3640;
	wire [4-1:0] node3641;
	wire [4-1:0] node3645;
	wire [4-1:0] node3646;
	wire [4-1:0] node3647;
	wire [4-1:0] node3648;
	wire [4-1:0] node3649;
	wire [4-1:0] node3650;
	wire [4-1:0] node3652;
	wire [4-1:0] node3656;
	wire [4-1:0] node3658;
	wire [4-1:0] node3659;
	wire [4-1:0] node3663;
	wire [4-1:0] node3664;
	wire [4-1:0] node3666;
	wire [4-1:0] node3669;
	wire [4-1:0] node3671;
	wire [4-1:0] node3674;
	wire [4-1:0] node3675;
	wire [4-1:0] node3676;
	wire [4-1:0] node3677;
	wire [4-1:0] node3678;
	wire [4-1:0] node3682;
	wire [4-1:0] node3684;
	wire [4-1:0] node3687;
	wire [4-1:0] node3688;
	wire [4-1:0] node3692;
	wire [4-1:0] node3693;
	wire [4-1:0] node3694;
	wire [4-1:0] node3698;
	wire [4-1:0] node3699;
	wire [4-1:0] node3700;
	wire [4-1:0] node3704;
	wire [4-1:0] node3705;
	wire [4-1:0] node3709;
	wire [4-1:0] node3710;
	wire [4-1:0] node3711;
	wire [4-1:0] node3712;
	wire [4-1:0] node3713;
	wire [4-1:0] node3714;
	wire [4-1:0] node3717;
	wire [4-1:0] node3718;
	wire [4-1:0] node3722;
	wire [4-1:0] node3723;
	wire [4-1:0] node3724;
	wire [4-1:0] node3728;
	wire [4-1:0] node3731;
	wire [4-1:0] node3732;
	wire [4-1:0] node3734;
	wire [4-1:0] node3737;
	wire [4-1:0] node3739;
	wire [4-1:0] node3742;
	wire [4-1:0] node3743;
	wire [4-1:0] node3744;
	wire [4-1:0] node3745;
	wire [4-1:0] node3748;
	wire [4-1:0] node3749;
	wire [4-1:0] node3753;
	wire [4-1:0] node3754;
	wire [4-1:0] node3755;
	wire [4-1:0] node3759;
	wire [4-1:0] node3760;
	wire [4-1:0] node3764;
	wire [4-1:0] node3765;
	wire [4-1:0] node3766;
	wire [4-1:0] node3770;
	wire [4-1:0] node3772;
	wire [4-1:0] node3775;
	wire [4-1:0] node3776;
	wire [4-1:0] node3777;
	wire [4-1:0] node3778;
	wire [4-1:0] node3779;
	wire [4-1:0] node3783;
	wire [4-1:0] node3784;
	wire [4-1:0] node3788;
	wire [4-1:0] node3789;
	wire [4-1:0] node3790;
	wire [4-1:0] node3792;
	wire [4-1:0] node3797;
	wire [4-1:0] node3798;
	wire [4-1:0] node3799;
	wire [4-1:0] node3800;
	wire [4-1:0] node3804;
	wire [4-1:0] node3805;
	wire [4-1:0] node3809;
	wire [4-1:0] node3810;
	wire [4-1:0] node3813;
	wire [4-1:0] node3814;
	wire [4-1:0] node3817;
	wire [4-1:0] node3818;
	wire [4-1:0] node3822;
	wire [4-1:0] node3824;
	wire [4-1:0] node3825;
	wire [4-1:0] node3826;
	wire [4-1:0] node3827;
	wire [4-1:0] node3828;
	wire [4-1:0] node3829;
	wire [4-1:0] node3830;
	wire [4-1:0] node3832;
	wire [4-1:0] node3836;
	wire [4-1:0] node3838;
	wire [4-1:0] node3841;
	wire [4-1:0] node3842;
	wire [4-1:0] node3843;
	wire [4-1:0] node3845;
	wire [4-1:0] node3849;
	wire [4-1:0] node3850;
	wire [4-1:0] node3852;
	wire [4-1:0] node3855;
	wire [4-1:0] node3858;
	wire [4-1:0] node3859;
	wire [4-1:0] node3860;
	wire [4-1:0] node3862;
	wire [4-1:0] node3866;
	wire [4-1:0] node3867;
	wire [4-1:0] node3871;
	wire [4-1:0] node3872;
	wire [4-1:0] node3873;
	wire [4-1:0] node3875;
	wire [4-1:0] node3876;
	wire [4-1:0] node3880;
	wire [4-1:0] node3881;
	wire [4-1:0] node3885;
	wire [4-1:0] node3886;
	wire [4-1:0] node3887;
	wire [4-1:0] node3888;
	wire [4-1:0] node3890;
	wire [4-1:0] node3894;
	wire [4-1:0] node3896;
	wire [4-1:0] node3899;
	wire [4-1:0] node3901;
	wire [4-1:0] node3903;
	wire [4-1:0] node3906;
	wire [4-1:0] node3908;
	wire [4-1:0] node3909;
	wire [4-1:0] node3910;
	wire [4-1:0] node3911;
	wire [4-1:0] node3912;
	wire [4-1:0] node3914;
	wire [4-1:0] node3917;
	wire [4-1:0] node3919;
	wire [4-1:0] node3923;
	wire [4-1:0] node3924;
	wire [4-1:0] node3925;
	wire [4-1:0] node3927;
	wire [4-1:0] node3931;
	wire [4-1:0] node3932;
	wire [4-1:0] node3936;
	wire [4-1:0] node3937;
	wire [4-1:0] node3938;
	wire [4-1:0] node3939;
	wire [4-1:0] node3943;
	wire [4-1:0] node3944;
	wire [4-1:0] node3948;
	wire [4-1:0] node3949;
	wire [4-1:0] node3951;
	wire [4-1:0] node3952;
	wire [4-1:0] node3955;
	wire [4-1:0] node3958;
	wire [4-1:0] node3959;
	wire [4-1:0] node3962;
	wire [4-1:0] node3966;
	wire [4-1:0] node3967;
	wire [4-1:0] node3968;
	wire [4-1:0] node3969;
	wire [4-1:0] node3970;
	wire [4-1:0] node3971;
	wire [4-1:0] node3972;
	wire [4-1:0] node3973;
	wire [4-1:0] node3974;
	wire [4-1:0] node3975;
	wire [4-1:0] node3976;
	wire [4-1:0] node3977;
	wire [4-1:0] node3981;
	wire [4-1:0] node3984;
	wire [4-1:0] node3985;
	wire [4-1:0] node3986;
	wire [4-1:0] node3990;
	wire [4-1:0] node3993;
	wire [4-1:0] node3994;
	wire [4-1:0] node3995;
	wire [4-1:0] node3996;
	wire [4-1:0] node4000;
	wire [4-1:0] node4001;
	wire [4-1:0] node4004;
	wire [4-1:0] node4007;
	wire [4-1:0] node4008;
	wire [4-1:0] node4009;
	wire [4-1:0] node4012;
	wire [4-1:0] node4015;
	wire [4-1:0] node4017;
	wire [4-1:0] node4020;
	wire [4-1:0] node4021;
	wire [4-1:0] node4022;
	wire [4-1:0] node4024;
	wire [4-1:0] node4028;
	wire [4-1:0] node4030;
	wire [4-1:0] node4033;
	wire [4-1:0] node4034;
	wire [4-1:0] node4035;
	wire [4-1:0] node4036;
	wire [4-1:0] node4037;
	wire [4-1:0] node4038;
	wire [4-1:0] node4042;
	wire [4-1:0] node4045;
	wire [4-1:0] node4046;
	wire [4-1:0] node4049;
	wire [4-1:0] node4052;
	wire [4-1:0] node4053;
	wire [4-1:0] node4054;
	wire [4-1:0] node4057;
	wire [4-1:0] node4060;
	wire [4-1:0] node4061;
	wire [4-1:0] node4063;
	wire [4-1:0] node4066;
	wire [4-1:0] node4068;
	wire [4-1:0] node4071;
	wire [4-1:0] node4072;
	wire [4-1:0] node4073;
	wire [4-1:0] node4075;
	wire [4-1:0] node4078;
	wire [4-1:0] node4079;
	wire [4-1:0] node4083;
	wire [4-1:0] node4084;
	wire [4-1:0] node4086;
	wire [4-1:0] node4089;
	wire [4-1:0] node4092;
	wire [4-1:0] node4093;
	wire [4-1:0] node4094;
	wire [4-1:0] node4095;
	wire [4-1:0] node4096;
	wire [4-1:0] node4098;
	wire [4-1:0] node4102;
	wire [4-1:0] node4103;
	wire [4-1:0] node4104;
	wire [4-1:0] node4108;
	wire [4-1:0] node4109;
	wire [4-1:0] node4113;
	wire [4-1:0] node4114;
	wire [4-1:0] node4115;
	wire [4-1:0] node4116;
	wire [4-1:0] node4117;
	wire [4-1:0] node4120;
	wire [4-1:0] node4123;
	wire [4-1:0] node4125;
	wire [4-1:0] node4128;
	wire [4-1:0] node4129;
	wire [4-1:0] node4132;
	wire [4-1:0] node4135;
	wire [4-1:0] node4136;
	wire [4-1:0] node4137;
	wire [4-1:0] node4141;
	wire [4-1:0] node4142;
	wire [4-1:0] node4146;
	wire [4-1:0] node4147;
	wire [4-1:0] node4148;
	wire [4-1:0] node4149;
	wire [4-1:0] node4151;
	wire [4-1:0] node4153;
	wire [4-1:0] node4157;
	wire [4-1:0] node4158;
	wire [4-1:0] node4159;
	wire [4-1:0] node4161;
	wire [4-1:0] node4164;
	wire [4-1:0] node4165;
	wire [4-1:0] node4170;
	wire [4-1:0] node4171;
	wire [4-1:0] node4172;
	wire [4-1:0] node4175;
	wire [4-1:0] node4178;
	wire [4-1:0] node4180;
	wire [4-1:0] node4182;
	wire [4-1:0] node4185;
	wire [4-1:0] node4186;
	wire [4-1:0] node4187;
	wire [4-1:0] node4188;
	wire [4-1:0] node4189;
	wire [4-1:0] node4190;
	wire [4-1:0] node4191;
	wire [4-1:0] node4192;
	wire [4-1:0] node4196;
	wire [4-1:0] node4197;
	wire [4-1:0] node4201;
	wire [4-1:0] node4202;
	wire [4-1:0] node4203;
	wire [4-1:0] node4206;
	wire [4-1:0] node4209;
	wire [4-1:0] node4210;
	wire [4-1:0] node4214;
	wire [4-1:0] node4215;
	wire [4-1:0] node4216;
	wire [4-1:0] node4219;
	wire [4-1:0] node4220;
	wire [4-1:0] node4224;
	wire [4-1:0] node4225;
	wire [4-1:0] node4226;
	wire [4-1:0] node4229;
	wire [4-1:0] node4232;
	wire [4-1:0] node4233;
	wire [4-1:0] node4236;
	wire [4-1:0] node4239;
	wire [4-1:0] node4240;
	wire [4-1:0] node4241;
	wire [4-1:0] node4243;
	wire [4-1:0] node4246;
	wire [4-1:0] node4247;
	wire [4-1:0] node4249;
	wire [4-1:0] node4252;
	wire [4-1:0] node4255;
	wire [4-1:0] node4256;
	wire [4-1:0] node4257;
	wire [4-1:0] node4258;
	wire [4-1:0] node4263;
	wire [4-1:0] node4265;
	wire [4-1:0] node4266;
	wire [4-1:0] node4270;
	wire [4-1:0] node4271;
	wire [4-1:0] node4272;
	wire [4-1:0] node4273;
	wire [4-1:0] node4274;
	wire [4-1:0] node4277;
	wire [4-1:0] node4280;
	wire [4-1:0] node4281;
	wire [4-1:0] node4284;
	wire [4-1:0] node4287;
	wire [4-1:0] node4288;
	wire [4-1:0] node4289;
	wire [4-1:0] node4290;
	wire [4-1:0] node4293;
	wire [4-1:0] node4297;
	wire [4-1:0] node4298;
	wire [4-1:0] node4300;
	wire [4-1:0] node4303;
	wire [4-1:0] node4306;
	wire [4-1:0] node4307;
	wire [4-1:0] node4308;
	wire [4-1:0] node4309;
	wire [4-1:0] node4312;
	wire [4-1:0] node4315;
	wire [4-1:0] node4316;
	wire [4-1:0] node4319;
	wire [4-1:0] node4322;
	wire [4-1:0] node4323;
	wire [4-1:0] node4324;
	wire [4-1:0] node4327;
	wire [4-1:0] node4330;
	wire [4-1:0] node4331;
	wire [4-1:0] node4334;
	wire [4-1:0] node4337;
	wire [4-1:0] node4338;
	wire [4-1:0] node4339;
	wire [4-1:0] node4340;
	wire [4-1:0] node4341;
	wire [4-1:0] node4342;
	wire [4-1:0] node4344;
	wire [4-1:0] node4347;
	wire [4-1:0] node4348;
	wire [4-1:0] node4351;
	wire [4-1:0] node4354;
	wire [4-1:0] node4355;
	wire [4-1:0] node4358;
	wire [4-1:0] node4361;
	wire [4-1:0] node4362;
	wire [4-1:0] node4363;
	wire [4-1:0] node4364;
	wire [4-1:0] node4368;
	wire [4-1:0] node4369;
	wire [4-1:0] node4372;
	wire [4-1:0] node4375;
	wire [4-1:0] node4376;
	wire [4-1:0] node4377;
	wire [4-1:0] node4380;
	wire [4-1:0] node4383;
	wire [4-1:0] node4384;
	wire [4-1:0] node4388;
	wire [4-1:0] node4389;
	wire [4-1:0] node4390;
	wire [4-1:0] node4392;
	wire [4-1:0] node4393;
	wire [4-1:0] node4397;
	wire [4-1:0] node4398;
	wire [4-1:0] node4399;
	wire [4-1:0] node4404;
	wire [4-1:0] node4405;
	wire [4-1:0] node4406;
	wire [4-1:0] node4410;
	wire [4-1:0] node4413;
	wire [4-1:0] node4414;
	wire [4-1:0] node4415;
	wire [4-1:0] node4417;
	wire [4-1:0] node4418;
	wire [4-1:0] node4419;
	wire [4-1:0] node4424;
	wire [4-1:0] node4425;
	wire [4-1:0] node4429;
	wire [4-1:0] node4430;
	wire [4-1:0] node4431;
	wire [4-1:0] node4432;
	wire [4-1:0] node4433;
	wire [4-1:0] node4437;
	wire [4-1:0] node4438;
	wire [4-1:0] node4441;
	wire [4-1:0] node4444;
	wire [4-1:0] node4445;
	wire [4-1:0] node4446;
	wire [4-1:0] node4449;
	wire [4-1:0] node4452;
	wire [4-1:0] node4455;
	wire [4-1:0] node4456;
	wire [4-1:0] node4457;
	wire [4-1:0] node4461;
	wire [4-1:0] node4464;
	wire [4-1:0] node4465;
	wire [4-1:0] node4466;
	wire [4-1:0] node4467;
	wire [4-1:0] node4468;
	wire [4-1:0] node4469;
	wire [4-1:0] node4470;
	wire [4-1:0] node4472;
	wire [4-1:0] node4475;
	wire [4-1:0] node4477;
	wire [4-1:0] node4480;
	wire [4-1:0] node4481;
	wire [4-1:0] node4483;
	wire [4-1:0] node4486;
	wire [4-1:0] node4489;
	wire [4-1:0] node4490;
	wire [4-1:0] node4492;
	wire [4-1:0] node4493;
	wire [4-1:0] node4497;
	wire [4-1:0] node4498;
	wire [4-1:0] node4502;
	wire [4-1:0] node4503;
	wire [4-1:0] node4504;
	wire [4-1:0] node4505;
	wire [4-1:0] node4509;
	wire [4-1:0] node4510;
	wire [4-1:0] node4514;
	wire [4-1:0] node4515;
	wire [4-1:0] node4516;
	wire [4-1:0] node4519;
	wire [4-1:0] node4520;
	wire [4-1:0] node4523;
	wire [4-1:0] node4526;
	wire [4-1:0] node4527;
	wire [4-1:0] node4528;
	wire [4-1:0] node4532;
	wire [4-1:0] node4535;
	wire [4-1:0] node4536;
	wire [4-1:0] node4537;
	wire [4-1:0] node4538;
	wire [4-1:0] node4539;
	wire [4-1:0] node4540;
	wire [4-1:0] node4544;
	wire [4-1:0] node4545;
	wire [4-1:0] node4549;
	wire [4-1:0] node4550;
	wire [4-1:0] node4553;
	wire [4-1:0] node4556;
	wire [4-1:0] node4557;
	wire [4-1:0] node4558;
	wire [4-1:0] node4559;
	wire [4-1:0] node4562;
	wire [4-1:0] node4565;
	wire [4-1:0] node4567;
	wire [4-1:0] node4570;
	wire [4-1:0] node4571;
	wire [4-1:0] node4572;
	wire [4-1:0] node4574;
	wire [4-1:0] node4577;
	wire [4-1:0] node4578;
	wire [4-1:0] node4581;
	wire [4-1:0] node4584;
	wire [4-1:0] node4585;
	wire [4-1:0] node4589;
	wire [4-1:0] node4590;
	wire [4-1:0] node4591;
	wire [4-1:0] node4592;
	wire [4-1:0] node4595;
	wire [4-1:0] node4596;
	wire [4-1:0] node4600;
	wire [4-1:0] node4601;
	wire [4-1:0] node4602;
	wire [4-1:0] node4606;
	wire [4-1:0] node4608;
	wire [4-1:0] node4611;
	wire [4-1:0] node4612;
	wire [4-1:0] node4614;
	wire [4-1:0] node4616;
	wire [4-1:0] node4619;
	wire [4-1:0] node4620;
	wire [4-1:0] node4623;
	wire [4-1:0] node4625;
	wire [4-1:0] node4628;
	wire [4-1:0] node4629;
	wire [4-1:0] node4630;
	wire [4-1:0] node4631;
	wire [4-1:0] node4632;
	wire [4-1:0] node4634;
	wire [4-1:0] node4635;
	wire [4-1:0] node4639;
	wire [4-1:0] node4642;
	wire [4-1:0] node4643;
	wire [4-1:0] node4644;
	wire [4-1:0] node4645;
	wire [4-1:0] node4649;
	wire [4-1:0] node4651;
	wire [4-1:0] node4654;
	wire [4-1:0] node4655;
	wire [4-1:0] node4657;
	wire [4-1:0] node4660;
	wire [4-1:0] node4661;
	wire [4-1:0] node4664;
	wire [4-1:0] node4667;
	wire [4-1:0] node4668;
	wire [4-1:0] node4669;
	wire [4-1:0] node4671;
	wire [4-1:0] node4673;
	wire [4-1:0] node4676;
	wire [4-1:0] node4677;
	wire [4-1:0] node4678;
	wire [4-1:0] node4680;
	wire [4-1:0] node4683;
	wire [4-1:0] node4684;
	wire [4-1:0] node4687;
	wire [4-1:0] node4690;
	wire [4-1:0] node4692;
	wire [4-1:0] node4695;
	wire [4-1:0] node4696;
	wire [4-1:0] node4697;
	wire [4-1:0] node4700;
	wire [4-1:0] node4701;
	wire [4-1:0] node4705;
	wire [4-1:0] node4706;
	wire [4-1:0] node4708;
	wire [4-1:0] node4710;
	wire [4-1:0] node4713;
	wire [4-1:0] node4714;
	wire [4-1:0] node4717;
	wire [4-1:0] node4720;
	wire [4-1:0] node4721;
	wire [4-1:0] node4722;
	wire [4-1:0] node4723;
	wire [4-1:0] node4724;
	wire [4-1:0] node4725;
	wire [4-1:0] node4729;
	wire [4-1:0] node4730;
	wire [4-1:0] node4733;
	wire [4-1:0] node4736;
	wire [4-1:0] node4737;
	wire [4-1:0] node4741;
	wire [4-1:0] node4742;
	wire [4-1:0] node4743;
	wire [4-1:0] node4746;
	wire [4-1:0] node4747;
	wire [4-1:0] node4751;
	wire [4-1:0] node4752;
	wire [4-1:0] node4755;
	wire [4-1:0] node4756;
	wire [4-1:0] node4757;
	wire [4-1:0] node4762;
	wire [4-1:0] node4763;
	wire [4-1:0] node4764;
	wire [4-1:0] node4766;
	wire [4-1:0] node4769;
	wire [4-1:0] node4772;
	wire [4-1:0] node4774;
	wire [4-1:0] node4777;
	wire [4-1:0] node4778;
	wire [4-1:0] node4779;
	wire [4-1:0] node4780;
	wire [4-1:0] node4781;
	wire [4-1:0] node4782;
	wire [4-1:0] node4783;
	wire [4-1:0] node4784;
	wire [4-1:0] node4785;
	wire [4-1:0] node4788;
	wire [4-1:0] node4789;
	wire [4-1:0] node4792;
	wire [4-1:0] node4795;
	wire [4-1:0] node4796;
	wire [4-1:0] node4797;
	wire [4-1:0] node4801;
	wire [4-1:0] node4803;
	wire [4-1:0] node4806;
	wire [4-1:0] node4807;
	wire [4-1:0] node4808;
	wire [4-1:0] node4809;
	wire [4-1:0] node4812;
	wire [4-1:0] node4815;
	wire [4-1:0] node4818;
	wire [4-1:0] node4820;
	wire [4-1:0] node4822;
	wire [4-1:0] node4825;
	wire [4-1:0] node4826;
	wire [4-1:0] node4827;
	wire [4-1:0] node4828;
	wire [4-1:0] node4831;
	wire [4-1:0] node4834;
	wire [4-1:0] node4835;
	wire [4-1:0] node4836;
	wire [4-1:0] node4840;
	wire [4-1:0] node4841;
	wire [4-1:0] node4845;
	wire [4-1:0] node4847;
	wire [4-1:0] node4848;
	wire [4-1:0] node4851;
	wire [4-1:0] node4852;
	wire [4-1:0] node4856;
	wire [4-1:0] node4857;
	wire [4-1:0] node4858;
	wire [4-1:0] node4859;
	wire [4-1:0] node4860;
	wire [4-1:0] node4864;
	wire [4-1:0] node4866;
	wire [4-1:0] node4869;
	wire [4-1:0] node4870;
	wire [4-1:0] node4874;
	wire [4-1:0] node4875;
	wire [4-1:0] node4876;
	wire [4-1:0] node4877;
	wire [4-1:0] node4880;
	wire [4-1:0] node4881;
	wire [4-1:0] node4885;
	wire [4-1:0] node4886;
	wire [4-1:0] node4887;
	wire [4-1:0] node4892;
	wire [4-1:0] node4893;
	wire [4-1:0] node4896;
	wire [4-1:0] node4899;
	wire [4-1:0] node4900;
	wire [4-1:0] node4901;
	wire [4-1:0] node4902;
	wire [4-1:0] node4903;
	wire [4-1:0] node4906;
	wire [4-1:0] node4908;
	wire [4-1:0] node4911;
	wire [4-1:0] node4912;
	wire [4-1:0] node4916;
	wire [4-1:0] node4917;
	wire [4-1:0] node4918;
	wire [4-1:0] node4920;
	wire [4-1:0] node4923;
	wire [4-1:0] node4924;
	wire [4-1:0] node4927;
	wire [4-1:0] node4930;
	wire [4-1:0] node4931;
	wire [4-1:0] node4932;
	wire [4-1:0] node4933;
	wire [4-1:0] node4936;
	wire [4-1:0] node4940;
	wire [4-1:0] node4941;
	wire [4-1:0] node4944;
	wire [4-1:0] node4947;
	wire [4-1:0] node4948;
	wire [4-1:0] node4949;
	wire [4-1:0] node4950;
	wire [4-1:0] node4951;
	wire [4-1:0] node4955;
	wire [4-1:0] node4958;
	wire [4-1:0] node4959;
	wire [4-1:0] node4960;
	wire [4-1:0] node4964;
	wire [4-1:0] node4967;
	wire [4-1:0] node4968;
	wire [4-1:0] node4970;
	wire [4-1:0] node4971;
	wire [4-1:0] node4975;
	wire [4-1:0] node4976;
	wire [4-1:0] node4977;
	wire [4-1:0] node4981;
	wire [4-1:0] node4984;
	wire [4-1:0] node4985;
	wire [4-1:0] node4986;
	wire [4-1:0] node4987;
	wire [4-1:0] node4988;
	wire [4-1:0] node4989;
	wire [4-1:0] node4992;
	wire [4-1:0] node4995;
	wire [4-1:0] node4996;
	wire [4-1:0] node4997;
	wire [4-1:0] node4999;
	wire [4-1:0] node5002;
	wire [4-1:0] node5005;
	wire [4-1:0] node5006;
	wire [4-1:0] node5010;
	wire [4-1:0] node5011;
	wire [4-1:0] node5012;
	wire [4-1:0] node5013;
	wire [4-1:0] node5017;
	wire [4-1:0] node5018;
	wire [4-1:0] node5022;
	wire [4-1:0] node5024;
	wire [4-1:0] node5025;
	wire [4-1:0] node5029;
	wire [4-1:0] node5030;
	wire [4-1:0] node5031;
	wire [4-1:0] node5032;
	wire [4-1:0] node5034;
	wire [4-1:0] node5037;
	wire [4-1:0] node5038;
	wire [4-1:0] node5040;
	wire [4-1:0] node5043;
	wire [4-1:0] node5045;
	wire [4-1:0] node5048;
	wire [4-1:0] node5049;
	wire [4-1:0] node5052;
	wire [4-1:0] node5054;
	wire [4-1:0] node5057;
	wire [4-1:0] node5058;
	wire [4-1:0] node5059;
	wire [4-1:0] node5060;
	wire [4-1:0] node5063;
	wire [4-1:0] node5065;
	wire [4-1:0] node5068;
	wire [4-1:0] node5069;
	wire [4-1:0] node5071;
	wire [4-1:0] node5075;
	wire [4-1:0] node5076;
	wire [4-1:0] node5077;
	wire [4-1:0] node5078;
	wire [4-1:0] node5081;
	wire [4-1:0] node5084;
	wire [4-1:0] node5085;
	wire [4-1:0] node5088;
	wire [4-1:0] node5092;
	wire [4-1:0] node5093;
	wire [4-1:0] node5094;
	wire [4-1:0] node5095;
	wire [4-1:0] node5096;
	wire [4-1:0] node5098;
	wire [4-1:0] node5101;
	wire [4-1:0] node5102;
	wire [4-1:0] node5105;
	wire [4-1:0] node5106;
	wire [4-1:0] node5110;
	wire [4-1:0] node5111;
	wire [4-1:0] node5112;
	wire [4-1:0] node5114;
	wire [4-1:0] node5119;
	wire [4-1:0] node5120;
	wire [4-1:0] node5121;
	wire [4-1:0] node5122;
	wire [4-1:0] node5124;
	wire [4-1:0] node5128;
	wire [4-1:0] node5129;
	wire [4-1:0] node5133;
	wire [4-1:0] node5134;
	wire [4-1:0] node5135;
	wire [4-1:0] node5139;
	wire [4-1:0] node5141;
	wire [4-1:0] node5143;
	wire [4-1:0] node5146;
	wire [4-1:0] node5147;
	wire [4-1:0] node5148;
	wire [4-1:0] node5149;
	wire [4-1:0] node5150;
	wire [4-1:0] node5153;
	wire [4-1:0] node5156;
	wire [4-1:0] node5158;
	wire [4-1:0] node5161;
	wire [4-1:0] node5162;
	wire [4-1:0] node5166;
	wire [4-1:0] node5167;
	wire [4-1:0] node5169;
	wire [4-1:0] node5170;
	wire [4-1:0] node5175;
	wire [4-1:0] node5176;
	wire [4-1:0] node5177;
	wire [4-1:0] node5178;
	wire [4-1:0] node5179;
	wire [4-1:0] node5180;
	wire [4-1:0] node5181;
	wire [4-1:0] node5182;
	wire [4-1:0] node5184;
	wire [4-1:0] node5187;
	wire [4-1:0] node5189;
	wire [4-1:0] node5192;
	wire [4-1:0] node5193;
	wire [4-1:0] node5194;
	wire [4-1:0] node5197;
	wire [4-1:0] node5200;
	wire [4-1:0] node5203;
	wire [4-1:0] node5204;
	wire [4-1:0] node5205;
	wire [4-1:0] node5207;
	wire [4-1:0] node5210;
	wire [4-1:0] node5214;
	wire [4-1:0] node5215;
	wire [4-1:0] node5216;
	wire [4-1:0] node5218;
	wire [4-1:0] node5219;
	wire [4-1:0] node5223;
	wire [4-1:0] node5224;
	wire [4-1:0] node5228;
	wire [4-1:0] node5229;
	wire [4-1:0] node5230;
	wire [4-1:0] node5233;
	wire [4-1:0] node5235;
	wire [4-1:0] node5238;
	wire [4-1:0] node5240;
	wire [4-1:0] node5243;
	wire [4-1:0] node5244;
	wire [4-1:0] node5245;
	wire [4-1:0] node5246;
	wire [4-1:0] node5248;
	wire [4-1:0] node5251;
	wire [4-1:0] node5252;
	wire [4-1:0] node5256;
	wire [4-1:0] node5257;
	wire [4-1:0] node5258;
	wire [4-1:0] node5261;
	wire [4-1:0] node5264;
	wire [4-1:0] node5265;
	wire [4-1:0] node5268;
	wire [4-1:0] node5271;
	wire [4-1:0] node5272;
	wire [4-1:0] node5273;
	wire [4-1:0] node5274;
	wire [4-1:0] node5276;
	wire [4-1:0] node5279;
	wire [4-1:0] node5282;
	wire [4-1:0] node5283;
	wire [4-1:0] node5286;
	wire [4-1:0] node5289;
	wire [4-1:0] node5290;
	wire [4-1:0] node5292;
	wire [4-1:0] node5295;
	wire [4-1:0] node5296;
	wire [4-1:0] node5298;
	wire [4-1:0] node5301;
	wire [4-1:0] node5302;
	wire [4-1:0] node5305;
	wire [4-1:0] node5308;
	wire [4-1:0] node5309;
	wire [4-1:0] node5310;
	wire [4-1:0] node5311;
	wire [4-1:0] node5312;
	wire [4-1:0] node5314;
	wire [4-1:0] node5316;
	wire [4-1:0] node5320;
	wire [4-1:0] node5321;
	wire [4-1:0] node5323;
	wire [4-1:0] node5326;
	wire [4-1:0] node5327;
	wire [4-1:0] node5329;
	wire [4-1:0] node5332;
	wire [4-1:0] node5335;
	wire [4-1:0] node5336;
	wire [4-1:0] node5337;
	wire [4-1:0] node5339;
	wire [4-1:0] node5341;
	wire [4-1:0] node5344;
	wire [4-1:0] node5345;
	wire [4-1:0] node5348;
	wire [4-1:0] node5351;
	wire [4-1:0] node5353;
	wire [4-1:0] node5354;
	wire [4-1:0] node5355;
	wire [4-1:0] node5359;
	wire [4-1:0] node5361;
	wire [4-1:0] node5364;
	wire [4-1:0] node5365;
	wire [4-1:0] node5366;
	wire [4-1:0] node5367;
	wire [4-1:0] node5369;
	wire [4-1:0] node5371;
	wire [4-1:0] node5374;
	wire [4-1:0] node5375;
	wire [4-1:0] node5376;
	wire [4-1:0] node5380;
	wire [4-1:0] node5381;
	wire [4-1:0] node5384;
	wire [4-1:0] node5387;
	wire [4-1:0] node5389;
	wire [4-1:0] node5392;
	wire [4-1:0] node5393;
	wire [4-1:0] node5394;
	wire [4-1:0] node5396;
	wire [4-1:0] node5399;
	wire [4-1:0] node5400;
	wire [4-1:0] node5403;
	wire [4-1:0] node5407;
	wire [4-1:0] node5408;
	wire [4-1:0] node5409;
	wire [4-1:0] node5410;
	wire [4-1:0] node5411;
	wire [4-1:0] node5413;
	wire [4-1:0] node5414;
	wire [4-1:0] node5418;
	wire [4-1:0] node5419;
	wire [4-1:0] node5420;
	wire [4-1:0] node5423;
	wire [4-1:0] node5424;
	wire [4-1:0] node5427;
	wire [4-1:0] node5430;
	wire [4-1:0] node5431;
	wire [4-1:0] node5432;
	wire [4-1:0] node5436;
	wire [4-1:0] node5439;
	wire [4-1:0] node5440;
	wire [4-1:0] node5441;
	wire [4-1:0] node5442;
	wire [4-1:0] node5444;
	wire [4-1:0] node5447;
	wire [4-1:0] node5448;
	wire [4-1:0] node5452;
	wire [4-1:0] node5453;
	wire [4-1:0] node5455;
	wire [4-1:0] node5458;
	wire [4-1:0] node5459;
	wire [4-1:0] node5463;
	wire [4-1:0] node5464;
	wire [4-1:0] node5466;
	wire [4-1:0] node5469;
	wire [4-1:0] node5471;
	wire [4-1:0] node5474;
	wire [4-1:0] node5475;
	wire [4-1:0] node5476;
	wire [4-1:0] node5477;
	wire [4-1:0] node5479;
	wire [4-1:0] node5480;
	wire [4-1:0] node5484;
	wire [4-1:0] node5485;
	wire [4-1:0] node5489;
	wire [4-1:0] node5490;
	wire [4-1:0] node5491;
	wire [4-1:0] node5493;
	wire [4-1:0] node5496;
	wire [4-1:0] node5499;
	wire [4-1:0] node5501;
	wire [4-1:0] node5504;
	wire [4-1:0] node5505;
	wire [4-1:0] node5506;
	wire [4-1:0] node5508;
	wire [4-1:0] node5511;
	wire [4-1:0] node5512;
	wire [4-1:0] node5513;
	wire [4-1:0] node5517;
	wire [4-1:0] node5519;
	wire [4-1:0] node5523;
	wire [4-1:0] node5524;
	wire [4-1:0] node5525;
	wire [4-1:0] node5526;
	wire [4-1:0] node5527;
	wire [4-1:0] node5528;
	wire [4-1:0] node5529;
	wire [4-1:0] node5533;
	wire [4-1:0] node5534;
	wire [4-1:0] node5538;
	wire [4-1:0] node5539;
	wire [4-1:0] node5540;
	wire [4-1:0] node5544;
	wire [4-1:0] node5547;
	wire [4-1:0] node5548;
	wire [4-1:0] node5549;
	wire [4-1:0] node5551;
	wire [4-1:0] node5555;
	wire [4-1:0] node5557;
	wire [4-1:0] node5558;
	wire [4-1:0] node5562;
	wire [4-1:0] node5563;
	wire [4-1:0] node5564;
	wire [4-1:0] node5565;
	wire [4-1:0] node5566;
	wire [4-1:0] node5571;
	wire [4-1:0] node5573;
	wire [4-1:0] node5577;
	wire [4-1:0] node5578;
	wire [4-1:0] node5579;
	wire [4-1:0] node5580;
	wire [4-1:0] node5581;
	wire [4-1:0] node5583;
	wire [4-1:0] node5587;
	wire [4-1:0] node5588;
	wire [4-1:0] node5589;
	wire [4-1:0] node5592;
	wire [4-1:0] node5598;
	wire [4-1:0] node5599;
	wire [4-1:0] node5600;
	wire [4-1:0] node5602;
	wire [4-1:0] node5603;
	wire [4-1:0] node5604;
	wire [4-1:0] node5605;
	wire [4-1:0] node5606;
	wire [4-1:0] node5608;
	wire [4-1:0] node5609;
	wire [4-1:0] node5613;
	wire [4-1:0] node5615;
	wire [4-1:0] node5618;
	wire [4-1:0] node5619;
	wire [4-1:0] node5620;
	wire [4-1:0] node5622;
	wire [4-1:0] node5625;
	wire [4-1:0] node5627;
	wire [4-1:0] node5630;
	wire [4-1:0] node5631;
	wire [4-1:0] node5633;
	wire [4-1:0] node5636;
	wire [4-1:0] node5637;
	wire [4-1:0] node5641;
	wire [4-1:0] node5642;
	wire [4-1:0] node5643;
	wire [4-1:0] node5645;
	wire [4-1:0] node5647;
	wire [4-1:0] node5648;
	wire [4-1:0] node5652;
	wire [4-1:0] node5654;
	wire [4-1:0] node5657;
	wire [4-1:0] node5658;
	wire [4-1:0] node5660;
	wire [4-1:0] node5661;
	wire [4-1:0] node5665;
	wire [4-1:0] node5667;
	wire [4-1:0] node5670;
	wire [4-1:0] node5672;
	wire [4-1:0] node5673;
	wire [4-1:0] node5674;
	wire [4-1:0] node5675;
	wire [4-1:0] node5676;
	wire [4-1:0] node5678;
	wire [4-1:0] node5681;
	wire [4-1:0] node5683;
	wire [4-1:0] node5687;
	wire [4-1:0] node5688;
	wire [4-1:0] node5689;
	wire [4-1:0] node5691;
	wire [4-1:0] node5696;
	wire [4-1:0] node5697;
	wire [4-1:0] node5698;
	wire [4-1:0] node5699;
	wire [4-1:0] node5701;
	wire [4-1:0] node5704;
	wire [4-1:0] node5705;
	wire [4-1:0] node5709;
	wire [4-1:0] node5711;
	wire [4-1:0] node5712;
	wire [4-1:0] node5716;
	wire [4-1:0] node5717;
	wire [4-1:0] node5719;
	wire [4-1:0] node5722;
	wire [4-1:0] node5726;
	wire [4-1:0] node5727;
	wire [4-1:0] node5728;
	wire [4-1:0] node5729;
	wire [4-1:0] node5730;
	wire [4-1:0] node5731;
	wire [4-1:0] node5732;
	wire [4-1:0] node5733;
	wire [4-1:0] node5734;
	wire [4-1:0] node5736;
	wire [4-1:0] node5739;
	wire [4-1:0] node5742;
	wire [4-1:0] node5744;
	wire [4-1:0] node5746;
	wire [4-1:0] node5749;
	wire [4-1:0] node5750;
	wire [4-1:0] node5751;
	wire [4-1:0] node5752;
	wire [4-1:0] node5756;
	wire [4-1:0] node5757;
	wire [4-1:0] node5760;
	wire [4-1:0] node5763;
	wire [4-1:0] node5764;
	wire [4-1:0] node5765;
	wire [4-1:0] node5769;
	wire [4-1:0] node5772;
	wire [4-1:0] node5773;
	wire [4-1:0] node5774;
	wire [4-1:0] node5775;
	wire [4-1:0] node5776;
	wire [4-1:0] node5781;
	wire [4-1:0] node5782;
	wire [4-1:0] node5783;
	wire [4-1:0] node5787;
	wire [4-1:0] node5790;
	wire [4-1:0] node5791;
	wire [4-1:0] node5793;
	wire [4-1:0] node5796;
	wire [4-1:0] node5797;
	wire [4-1:0] node5798;
	wire [4-1:0] node5801;
	wire [4-1:0] node5805;
	wire [4-1:0] node5806;
	wire [4-1:0] node5807;
	wire [4-1:0] node5808;
	wire [4-1:0] node5810;
	wire [4-1:0] node5811;
	wire [4-1:0] node5816;
	wire [4-1:0] node5817;
	wire [4-1:0] node5821;
	wire [4-1:0] node5822;
	wire [4-1:0] node5823;
	wire [4-1:0] node5825;
	wire [4-1:0] node5826;
	wire [4-1:0] node5830;
	wire [4-1:0] node5831;
	wire [4-1:0] node5834;
	wire [4-1:0] node5836;
	wire [4-1:0] node5839;
	wire [4-1:0] node5840;
	wire [4-1:0] node5842;
	wire [4-1:0] node5843;
	wire [4-1:0] node5847;
	wire [4-1:0] node5849;
	wire [4-1:0] node5852;
	wire [4-1:0] node5853;
	wire [4-1:0] node5854;
	wire [4-1:0] node5855;
	wire [4-1:0] node5856;
	wire [4-1:0] node5858;
	wire [4-1:0] node5861;
	wire [4-1:0] node5863;
	wire [4-1:0] node5866;
	wire [4-1:0] node5867;
	wire [4-1:0] node5870;
	wire [4-1:0] node5871;
	wire [4-1:0] node5875;
	wire [4-1:0] node5876;
	wire [4-1:0] node5877;
	wire [4-1:0] node5880;
	wire [4-1:0] node5883;
	wire [4-1:0] node5884;
	wire [4-1:0] node5886;
	wire [4-1:0] node5889;
	wire [4-1:0] node5890;
	wire [4-1:0] node5893;
	wire [4-1:0] node5896;
	wire [4-1:0] node5897;
	wire [4-1:0] node5898;
	wire [4-1:0] node5899;
	wire [4-1:0] node5900;
	wire [4-1:0] node5903;
	wire [4-1:0] node5906;
	wire [4-1:0] node5907;
	wire [4-1:0] node5910;
	wire [4-1:0] node5913;
	wire [4-1:0] node5914;
	wire [4-1:0] node5916;
	wire [4-1:0] node5920;
	wire [4-1:0] node5921;
	wire [4-1:0] node5922;
	wire [4-1:0] node5925;
	wire [4-1:0] node5928;
	wire [4-1:0] node5929;
	wire [4-1:0] node5933;
	wire [4-1:0] node5934;
	wire [4-1:0] node5935;
	wire [4-1:0] node5936;
	wire [4-1:0] node5937;
	wire [4-1:0] node5939;
	wire [4-1:0] node5942;
	wire [4-1:0] node5944;
	wire [4-1:0] node5946;
	wire [4-1:0] node5949;
	wire [4-1:0] node5950;
	wire [4-1:0] node5951;
	wire [4-1:0] node5953;
	wire [4-1:0] node5956;
	wire [4-1:0] node5957;
	wire [4-1:0] node5960;
	wire [4-1:0] node5963;
	wire [4-1:0] node5964;
	wire [4-1:0] node5965;
	wire [4-1:0] node5970;
	wire [4-1:0] node5971;
	wire [4-1:0] node5972;
	wire [4-1:0] node5973;
	wire [4-1:0] node5974;
	wire [4-1:0] node5978;
	wire [4-1:0] node5979;
	wire [4-1:0] node5981;
	wire [4-1:0] node5985;
	wire [4-1:0] node5986;
	wire [4-1:0] node5987;
	wire [4-1:0] node5988;
	wire [4-1:0] node5994;
	wire [4-1:0] node5995;
	wire [4-1:0] node5996;
	wire [4-1:0] node5997;
	wire [4-1:0] node6001;
	wire [4-1:0] node6002;
	wire [4-1:0] node6004;
	wire [4-1:0] node6007;
	wire [4-1:0] node6011;
	wire [4-1:0] node6012;
	wire [4-1:0] node6013;
	wire [4-1:0] node6014;
	wire [4-1:0] node6015;
	wire [4-1:0] node6017;
	wire [4-1:0] node6020;
	wire [4-1:0] node6023;
	wire [4-1:0] node6024;
	wire [4-1:0] node6025;
	wire [4-1:0] node6026;
	wire [4-1:0] node6029;
	wire [4-1:0] node6032;
	wire [4-1:0] node6033;
	wire [4-1:0] node6037;
	wire [4-1:0] node6040;
	wire [4-1:0] node6041;
	wire [4-1:0] node6042;
	wire [4-1:0] node6043;
	wire [4-1:0] node6044;
	wire [4-1:0] node6048;
	wire [4-1:0] node6051;
	wire [4-1:0] node6054;
	wire [4-1:0] node6055;
	wire [4-1:0] node6056;
	wire [4-1:0] node6061;
	wire [4-1:0] node6062;
	wire [4-1:0] node6063;
	wire [4-1:0] node6064;
	wire [4-1:0] node6065;
	wire [4-1:0] node6066;
	wire [4-1:0] node6069;
	wire [4-1:0] node6072;
	wire [4-1:0] node6074;
	wire [4-1:0] node6078;
	wire [4-1:0] node6079;
	wire [4-1:0] node6081;
	wire [4-1:0] node6082;
	wire [4-1:0] node6087;
	wire [4-1:0] node6088;
	wire [4-1:0] node6089;
	wire [4-1:0] node6090;
	wire [4-1:0] node6091;
	wire [4-1:0] node6098;
	wire [4-1:0] node6100;
	wire [4-1:0] node6101;
	wire [4-1:0] node6102;
	wire [4-1:0] node6103;
	wire [4-1:0] node6104;
	wire [4-1:0] node6105;
	wire [4-1:0] node6106;
	wire [4-1:0] node6110;
	wire [4-1:0] node6112;
	wire [4-1:0] node6115;
	wire [4-1:0] node6116;
	wire [4-1:0] node6118;
	wire [4-1:0] node6121;
	wire [4-1:0] node6122;
	wire [4-1:0] node6125;
	wire [4-1:0] node6128;
	wire [4-1:0] node6129;
	wire [4-1:0] node6130;
	wire [4-1:0] node6132;
	wire [4-1:0] node6135;
	wire [4-1:0] node6137;
	wire [4-1:0] node6138;
	wire [4-1:0] node6142;
	wire [4-1:0] node6143;
	wire [4-1:0] node6146;
	wire [4-1:0] node6147;
	wire [4-1:0] node6152;
	wire [4-1:0] node6153;
	wire [4-1:0] node6154;
	wire [4-1:0] node6155;
	wire [4-1:0] node6156;
	wire [4-1:0] node6159;
	wire [4-1:0] node6160;
	wire [4-1:0] node6161;
	wire [4-1:0] node6165;
	wire [4-1:0] node6168;
	wire [4-1:0] node6169;
	wire [4-1:0] node6170;
	wire [4-1:0] node6172;
	wire [4-1:0] node6175;
	wire [4-1:0] node6179;
	wire [4-1:0] node6180;
	wire [4-1:0] node6181;
	wire [4-1:0] node6183;
	wire [4-1:0] node6184;
	wire [4-1:0] node6187;
	wire [4-1:0] node6190;
	wire [4-1:0] node6191;
	wire [4-1:0] node6195;
	wire [4-1:0] node6196;
	wire [4-1:0] node6197;
	wire [4-1:0] node6200;
	wire [4-1:0] node6204;
	wire [4-1:0] node6205;
	wire [4-1:0] node6206;
	wire [4-1:0] node6207;
	wire [4-1:0] node6208;
	wire [4-1:0] node6210;
	wire [4-1:0] node6214;
	wire [4-1:0] node6215;
	wire [4-1:0] node6217;
	wire [4-1:0] node6221;
	wire [4-1:0] node6222;
	wire [4-1:0] node6223;
	wire [4-1:0] node6224;
	wire [4-1:0] node6227;
	wire [4-1:0] node6232;
	wire [4-1:0] node6233;
	wire [4-1:0] node6234;
	wire [4-1:0] node6236;
	wire [4-1:0] node6237;
	wire [4-1:0] node6240;
	wire [4-1:0] node6245;
	wire [4-1:0] node6246;
	wire [4-1:0] node6247;
	wire [4-1:0] node6248;
	wire [4-1:0] node6249;
	wire [4-1:0] node6250;
	wire [4-1:0] node6251;
	wire [4-1:0] node6252;
	wire [4-1:0] node6253;
	wire [4-1:0] node6254;
	wire [4-1:0] node6255;
	wire [4-1:0] node6257;
	wire [4-1:0] node6259;
	wire [4-1:0] node6262;
	wire [4-1:0] node6263;
	wire [4-1:0] node6265;
	wire [4-1:0] node6268;
	wire [4-1:0] node6270;
	wire [4-1:0] node6273;
	wire [4-1:0] node6274;
	wire [4-1:0] node6276;
	wire [4-1:0] node6280;
	wire [4-1:0] node6281;
	wire [4-1:0] node6282;
	wire [4-1:0] node6283;
	wire [4-1:0] node6285;
	wire [4-1:0] node6288;
	wire [4-1:0] node6290;
	wire [4-1:0] node6293;
	wire [4-1:0] node6294;
	wire [4-1:0] node6298;
	wire [4-1:0] node6299;
	wire [4-1:0] node6301;
	wire [4-1:0] node6304;
	wire [4-1:0] node6305;
	wire [4-1:0] node6306;
	wire [4-1:0] node6311;
	wire [4-1:0] node6312;
	wire [4-1:0] node6313;
	wire [4-1:0] node6314;
	wire [4-1:0] node6318;
	wire [4-1:0] node6319;
	wire [4-1:0] node6321;
	wire [4-1:0] node6324;
	wire [4-1:0] node6326;
	wire [4-1:0] node6329;
	wire [4-1:0] node6330;
	wire [4-1:0] node6331;
	wire [4-1:0] node6333;
	wire [4-1:0] node6337;
	wire [4-1:0] node6338;
	wire [4-1:0] node6340;
	wire [4-1:0] node6343;
	wire [4-1:0] node6345;
	wire [4-1:0] node6348;
	wire [4-1:0] node6349;
	wire [4-1:0] node6350;
	wire [4-1:0] node6351;
	wire [4-1:0] node6352;
	wire [4-1:0] node6353;
	wire [4-1:0] node6354;
	wire [4-1:0] node6358;
	wire [4-1:0] node6360;
	wire [4-1:0] node6362;
	wire [4-1:0] node6365;
	wire [4-1:0] node6367;
	wire [4-1:0] node6369;
	wire [4-1:0] node6372;
	wire [4-1:0] node6373;
	wire [4-1:0] node6374;
	wire [4-1:0] node6375;
	wire [4-1:0] node6379;
	wire [4-1:0] node6381;
	wire [4-1:0] node6382;
	wire [4-1:0] node6386;
	wire [4-1:0] node6387;
	wire [4-1:0] node6388;
	wire [4-1:0] node6390;
	wire [4-1:0] node6393;
	wire [4-1:0] node6395;
	wire [4-1:0] node6398;
	wire [4-1:0] node6399;
	wire [4-1:0] node6400;
	wire [4-1:0] node6404;
	wire [4-1:0] node6407;
	wire [4-1:0] node6408;
	wire [4-1:0] node6409;
	wire [4-1:0] node6410;
	wire [4-1:0] node6414;
	wire [4-1:0] node6415;
	wire [4-1:0] node6417;
	wire [4-1:0] node6420;
	wire [4-1:0] node6421;
	wire [4-1:0] node6425;
	wire [4-1:0] node6426;
	wire [4-1:0] node6427;
	wire [4-1:0] node6429;
	wire [4-1:0] node6433;
	wire [4-1:0] node6434;
	wire [4-1:0] node6436;
	wire [4-1:0] node6439;
	wire [4-1:0] node6440;
	wire [4-1:0] node6444;
	wire [4-1:0] node6445;
	wire [4-1:0] node6446;
	wire [4-1:0] node6447;
	wire [4-1:0] node6448;
	wire [4-1:0] node6450;
	wire [4-1:0] node6452;
	wire [4-1:0] node6455;
	wire [4-1:0] node6456;
	wire [4-1:0] node6459;
	wire [4-1:0] node6460;
	wire [4-1:0] node6464;
	wire [4-1:0] node6465;
	wire [4-1:0] node6467;
	wire [4-1:0] node6471;
	wire [4-1:0] node6472;
	wire [4-1:0] node6474;
	wire [4-1:0] node6475;
	wire [4-1:0] node6479;
	wire [4-1:0] node6480;
	wire [4-1:0] node6483;
	wire [4-1:0] node6484;
	wire [4-1:0] node6485;
	wire [4-1:0] node6490;
	wire [4-1:0] node6491;
	wire [4-1:0] node6492;
	wire [4-1:0] node6493;
	wire [4-1:0] node6496;
	wire [4-1:0] node6497;
	wire [4-1:0] node6501;
	wire [4-1:0] node6503;
	wire [4-1:0] node6506;
	wire [4-1:0] node6507;
	wire [4-1:0] node6508;
	wire [4-1:0] node6510;
	wire [4-1:0] node6514;
	wire [4-1:0] node6516;
	wire [4-1:0] node6517;
	wire [4-1:0] node6521;
	wire [4-1:0] node6522;
	wire [4-1:0] node6523;
	wire [4-1:0] node6524;
	wire [4-1:0] node6525;
	wire [4-1:0] node6526;
	wire [4-1:0] node6528;
	wire [4-1:0] node6531;
	wire [4-1:0] node6532;
	wire [4-1:0] node6533;
	wire [4-1:0] node6536;
	wire [4-1:0] node6537;
	wire [4-1:0] node6541;
	wire [4-1:0] node6543;
	wire [4-1:0] node6546;
	wire [4-1:0] node6547;
	wire [4-1:0] node6548;
	wire [4-1:0] node6550;
	wire [4-1:0] node6553;
	wire [4-1:0] node6555;
	wire [4-1:0] node6558;
	wire [4-1:0] node6559;
	wire [4-1:0] node6563;
	wire [4-1:0] node6564;
	wire [4-1:0] node6565;
	wire [4-1:0] node6567;
	wire [4-1:0] node6568;
	wire [4-1:0] node6572;
	wire [4-1:0] node6573;
	wire [4-1:0] node6575;
	wire [4-1:0] node6577;
	wire [4-1:0] node6580;
	wire [4-1:0] node6582;
	wire [4-1:0] node6585;
	wire [4-1:0] node6586;
	wire [4-1:0] node6587;
	wire [4-1:0] node6591;
	wire [4-1:0] node6593;
	wire [4-1:0] node6596;
	wire [4-1:0] node6597;
	wire [4-1:0] node6598;
	wire [4-1:0] node6599;
	wire [4-1:0] node6601;
	wire [4-1:0] node6602;
	wire [4-1:0] node6603;
	wire [4-1:0] node6608;
	wire [4-1:0] node6609;
	wire [4-1:0] node6610;
	wire [4-1:0] node6613;
	wire [4-1:0] node6615;
	wire [4-1:0] node6618;
	wire [4-1:0] node6620;
	wire [4-1:0] node6623;
	wire [4-1:0] node6624;
	wire [4-1:0] node6625;
	wire [4-1:0] node6628;
	wire [4-1:0] node6629;
	wire [4-1:0] node6633;
	wire [4-1:0] node6635;
	wire [4-1:0] node6638;
	wire [4-1:0] node6639;
	wire [4-1:0] node6640;
	wire [4-1:0] node6641;
	wire [4-1:0] node6642;
	wire [4-1:0] node6646;
	wire [4-1:0] node6647;
	wire [4-1:0] node6648;
	wire [4-1:0] node6652;
	wire [4-1:0] node6654;
	wire [4-1:0] node6657;
	wire [4-1:0] node6659;
	wire [4-1:0] node6660;
	wire [4-1:0] node6662;
	wire [4-1:0] node6665;
	wire [4-1:0] node6666;
	wire [4-1:0] node6670;
	wire [4-1:0] node6671;
	wire [4-1:0] node6672;
	wire [4-1:0] node6676;
	wire [4-1:0] node6677;
	wire [4-1:0] node6678;
	wire [4-1:0] node6682;
	wire [4-1:0] node6683;
	wire [4-1:0] node6687;
	wire [4-1:0] node6688;
	wire [4-1:0] node6689;
	wire [4-1:0] node6690;
	wire [4-1:0] node6691;
	wire [4-1:0] node6693;
	wire [4-1:0] node6697;
	wire [4-1:0] node6698;
	wire [4-1:0] node6699;
	wire [4-1:0] node6701;
	wire [4-1:0] node6704;
	wire [4-1:0] node6705;
	wire [4-1:0] node6707;
	wire [4-1:0] node6711;
	wire [4-1:0] node6712;
	wire [4-1:0] node6716;
	wire [4-1:0] node6717;
	wire [4-1:0] node6718;
	wire [4-1:0] node6720;
	wire [4-1:0] node6724;
	wire [4-1:0] node6725;
	wire [4-1:0] node6729;
	wire [4-1:0] node6730;
	wire [4-1:0] node6731;
	wire [4-1:0] node6732;
	wire [4-1:0] node6733;
	wire [4-1:0] node6735;
	wire [4-1:0] node6739;
	wire [4-1:0] node6740;
	wire [4-1:0] node6744;
	wire [4-1:0] node6745;
	wire [4-1:0] node6746;
	wire [4-1:0] node6748;
	wire [4-1:0] node6751;
	wire [4-1:0] node6754;
	wire [4-1:0] node6755;
	wire [4-1:0] node6759;
	wire [4-1:0] node6760;
	wire [4-1:0] node6761;
	wire [4-1:0] node6763;
	wire [4-1:0] node6767;
	wire [4-1:0] node6768;
	wire [4-1:0] node6772;
	wire [4-1:0] node6774;
	wire [4-1:0] node6775;
	wire [4-1:0] node6776;
	wire [4-1:0] node6778;
	wire [4-1:0] node6779;
	wire [4-1:0] node6780;
	wire [4-1:0] node6781;
	wire [4-1:0] node6783;
	wire [4-1:0] node6786;
	wire [4-1:0] node6788;
	wire [4-1:0] node6791;
	wire [4-1:0] node6793;
	wire [4-1:0] node6794;
	wire [4-1:0] node6797;
	wire [4-1:0] node6801;
	wire [4-1:0] node6802;
	wire [4-1:0] node6803;
	wire [4-1:0] node6804;
	wire [4-1:0] node6805;
	wire [4-1:0] node6806;
	wire [4-1:0] node6809;
	wire [4-1:0] node6811;
	wire [4-1:0] node6814;
	wire [4-1:0] node6816;
	wire [4-1:0] node6819;
	wire [4-1:0] node6820;
	wire [4-1:0] node6821;
	wire [4-1:0] node6822;
	wire [4-1:0] node6828;
	wire [4-1:0] node6829;
	wire [4-1:0] node6830;
	wire [4-1:0] node6832;
	wire [4-1:0] node6835;
	wire [4-1:0] node6837;
	wire [4-1:0] node6840;
	wire [4-1:0] node6841;
	wire [4-1:0] node6842;
	wire [4-1:0] node6844;
	wire [4-1:0] node6847;
	wire [4-1:0] node6849;
	wire [4-1:0] node6852;
	wire [4-1:0] node6853;
	wire [4-1:0] node6854;
	wire [4-1:0] node6857;
	wire [4-1:0] node6861;
	wire [4-1:0] node6863;
	wire [4-1:0] node6864;
	wire [4-1:0] node6865;
	wire [4-1:0] node6869;
	wire [4-1:0] node6870;
	wire [4-1:0] node6872;
	wire [4-1:0] node6875;
	wire [4-1:0] node6877;
	wire [4-1:0] node6880;
	wire [4-1:0] node6881;
	wire [4-1:0] node6882;
	wire [4-1:0] node6883;
	wire [4-1:0] node6884;
	wire [4-1:0] node6885;
	wire [4-1:0] node6889;
	wire [4-1:0] node6890;
	wire [4-1:0] node6893;
	wire [4-1:0] node6896;
	wire [4-1:0] node6897;
	wire [4-1:0] node6898;
	wire [4-1:0] node6899;
	wire [4-1:0] node6903;
	wire [4-1:0] node6904;
	wire [4-1:0] node6908;
	wire [4-1:0] node6909;
	wire [4-1:0] node6912;
	wire [4-1:0] node6913;
	wire [4-1:0] node6917;
	wire [4-1:0] node6918;
	wire [4-1:0] node6919;
	wire [4-1:0] node6920;
	wire [4-1:0] node6924;
	wire [4-1:0] node6925;
	wire [4-1:0] node6927;
	wire [4-1:0] node6930;
	wire [4-1:0] node6931;
	wire [4-1:0] node6935;
	wire [4-1:0] node6936;
	wire [4-1:0] node6937;
	wire [4-1:0] node6938;
	wire [4-1:0] node6942;
	wire [4-1:0] node6943;
	wire [4-1:0] node6947;
	wire [4-1:0] node6948;
	wire [4-1:0] node6949;
	wire [4-1:0] node6953;
	wire [4-1:0] node6954;
	wire [4-1:0] node6955;
	wire [4-1:0] node6959;
	wire [4-1:0] node6962;
	wire [4-1:0] node6963;
	wire [4-1:0] node6964;
	wire [4-1:0] node6965;
	wire [4-1:0] node6966;
	wire [4-1:0] node6967;
	wire [4-1:0] node6969;
	wire [4-1:0] node6973;
	wire [4-1:0] node6974;
	wire [4-1:0] node6976;
	wire [4-1:0] node6979;
	wire [4-1:0] node6980;
	wire [4-1:0] node6984;
	wire [4-1:0] node6985;
	wire [4-1:0] node6987;
	wire [4-1:0] node6990;
	wire [4-1:0] node6991;
	wire [4-1:0] node6995;
	wire [4-1:0] node6996;
	wire [4-1:0] node6997;
	wire [4-1:0] node6998;
	wire [4-1:0] node7001;
	wire [4-1:0] node7003;
	wire [4-1:0] node7007;
	wire [4-1:0] node7008;
	wire [4-1:0] node7010;
	wire [4-1:0] node7012;
	wire [4-1:0] node7015;
	wire [4-1:0] node7016;
	wire [4-1:0] node7020;
	wire [4-1:0] node7021;
	wire [4-1:0] node7022;
	wire [4-1:0] node7023;
	wire [4-1:0] node7024;
	wire [4-1:0] node7025;
	wire [4-1:0] node7029;
	wire [4-1:0] node7030;
	wire [4-1:0] node7035;
	wire [4-1:0] node7036;
	wire [4-1:0] node7038;
	wire [4-1:0] node7041;
	wire [4-1:0] node7042;
	wire [4-1:0] node7043;
	wire [4-1:0] node7047;
	wire [4-1:0] node7050;
	wire [4-1:0] node7051;
	wire [4-1:0] node7052;
	wire [4-1:0] node7054;
	wire [4-1:0] node7055;
	wire [4-1:0] node7059;
	wire [4-1:0] node7061;
	wire [4-1:0] node7064;
	wire [4-1:0] node7065;
	wire [4-1:0] node7066;
	wire [4-1:0] node7069;
	wire [4-1:0] node7072;
	wire [4-1:0] node7073;
	wire [4-1:0] node7076;
	wire [4-1:0] node7078;
	wire [4-1:0] node7082;
	wire [4-1:0] node7083;
	wire [4-1:0] node7084;
	wire [4-1:0] node7085;
	wire [4-1:0] node7086;
	wire [4-1:0] node7087;
	wire [4-1:0] node7088;
	wire [4-1:0] node7089;
	wire [4-1:0] node7090;
	wire [4-1:0] node7091;
	wire [4-1:0] node7092;
	wire [4-1:0] node7095;
	wire [4-1:0] node7098;
	wire [4-1:0] node7100;
	wire [4-1:0] node7103;
	wire [4-1:0] node7104;
	wire [4-1:0] node7105;
	wire [4-1:0] node7109;
	wire [4-1:0] node7110;
	wire [4-1:0] node7112;
	wire [4-1:0] node7115;
	wire [4-1:0] node7116;
	wire [4-1:0] node7119;
	wire [4-1:0] node7122;
	wire [4-1:0] node7123;
	wire [4-1:0] node7124;
	wire [4-1:0] node7126;
	wire [4-1:0] node7129;
	wire [4-1:0] node7130;
	wire [4-1:0] node7134;
	wire [4-1:0] node7135;
	wire [4-1:0] node7139;
	wire [4-1:0] node7140;
	wire [4-1:0] node7141;
	wire [4-1:0] node7143;
	wire [4-1:0] node7144;
	wire [4-1:0] node7146;
	wire [4-1:0] node7150;
	wire [4-1:0] node7151;
	wire [4-1:0] node7155;
	wire [4-1:0] node7156;
	wire [4-1:0] node7157;
	wire [4-1:0] node7158;
	wire [4-1:0] node7161;
	wire [4-1:0] node7163;
	wire [4-1:0] node7166;
	wire [4-1:0] node7167;
	wire [4-1:0] node7171;
	wire [4-1:0] node7172;
	wire [4-1:0] node7174;
	wire [4-1:0] node7177;
	wire [4-1:0] node7179;
	wire [4-1:0] node7182;
	wire [4-1:0] node7183;
	wire [4-1:0] node7184;
	wire [4-1:0] node7185;
	wire [4-1:0] node7186;
	wire [4-1:0] node7187;
	wire [4-1:0] node7190;
	wire [4-1:0] node7193;
	wire [4-1:0] node7195;
	wire [4-1:0] node7197;
	wire [4-1:0] node7200;
	wire [4-1:0] node7201;
	wire [4-1:0] node7202;
	wire [4-1:0] node7206;
	wire [4-1:0] node7207;
	wire [4-1:0] node7208;
	wire [4-1:0] node7211;
	wire [4-1:0] node7214;
	wire [4-1:0] node7215;
	wire [4-1:0] node7218;
	wire [4-1:0] node7221;
	wire [4-1:0] node7222;
	wire [4-1:0] node7223;
	wire [4-1:0] node7224;
	wire [4-1:0] node7225;
	wire [4-1:0] node7228;
	wire [4-1:0] node7232;
	wire [4-1:0] node7233;
	wire [4-1:0] node7237;
	wire [4-1:0] node7238;
	wire [4-1:0] node7240;
	wire [4-1:0] node7242;
	wire [4-1:0] node7245;
	wire [4-1:0] node7246;
	wire [4-1:0] node7249;
	wire [4-1:0] node7252;
	wire [4-1:0] node7253;
	wire [4-1:0] node7254;
	wire [4-1:0] node7255;
	wire [4-1:0] node7256;
	wire [4-1:0] node7259;
	wire [4-1:0] node7262;
	wire [4-1:0] node7263;
	wire [4-1:0] node7265;
	wire [4-1:0] node7268;
	wire [4-1:0] node7271;
	wire [4-1:0] node7272;
	wire [4-1:0] node7273;
	wire [4-1:0] node7274;
	wire [4-1:0] node7277;
	wire [4-1:0] node7280;
	wire [4-1:0] node7281;
	wire [4-1:0] node7284;
	wire [4-1:0] node7287;
	wire [4-1:0] node7288;
	wire [4-1:0] node7291;
	wire [4-1:0] node7294;
	wire [4-1:0] node7295;
	wire [4-1:0] node7296;
	wire [4-1:0] node7297;
	wire [4-1:0] node7298;
	wire [4-1:0] node7302;
	wire [4-1:0] node7305;
	wire [4-1:0] node7306;
	wire [4-1:0] node7309;
	wire [4-1:0] node7312;
	wire [4-1:0] node7313;
	wire [4-1:0] node7314;
	wire [4-1:0] node7316;
	wire [4-1:0] node7319;
	wire [4-1:0] node7321;
	wire [4-1:0] node7324;
	wire [4-1:0] node7325;
	wire [4-1:0] node7326;
	wire [4-1:0] node7330;
	wire [4-1:0] node7333;
	wire [4-1:0] node7334;
	wire [4-1:0] node7335;
	wire [4-1:0] node7336;
	wire [4-1:0] node7337;
	wire [4-1:0] node7338;
	wire [4-1:0] node7341;
	wire [4-1:0] node7342;
	wire [4-1:0] node7343;
	wire [4-1:0] node7347;
	wire [4-1:0] node7350;
	wire [4-1:0] node7352;
	wire [4-1:0] node7353;
	wire [4-1:0] node7355;
	wire [4-1:0] node7359;
	wire [4-1:0] node7360;
	wire [4-1:0] node7361;
	wire [4-1:0] node7363;
	wire [4-1:0] node7366;
	wire [4-1:0] node7367;
	wire [4-1:0] node7368;
	wire [4-1:0] node7373;
	wire [4-1:0] node7374;
	wire [4-1:0] node7375;
	wire [4-1:0] node7377;
	wire [4-1:0] node7380;
	wire [4-1:0] node7383;
	wire [4-1:0] node7384;
	wire [4-1:0] node7386;
	wire [4-1:0] node7389;
	wire [4-1:0] node7390;
	wire [4-1:0] node7394;
	wire [4-1:0] node7395;
	wire [4-1:0] node7396;
	wire [4-1:0] node7398;
	wire [4-1:0] node7401;
	wire [4-1:0] node7402;
	wire [4-1:0] node7403;
	wire [4-1:0] node7406;
	wire [4-1:0] node7407;
	wire [4-1:0] node7410;
	wire [4-1:0] node7413;
	wire [4-1:0] node7414;
	wire [4-1:0] node7417;
	wire [4-1:0] node7420;
	wire [4-1:0] node7421;
	wire [4-1:0] node7422;
	wire [4-1:0] node7423;
	wire [4-1:0] node7426;
	wire [4-1:0] node7429;
	wire [4-1:0] node7431;
	wire [4-1:0] node7434;
	wire [4-1:0] node7436;
	wire [4-1:0] node7439;
	wire [4-1:0] node7440;
	wire [4-1:0] node7441;
	wire [4-1:0] node7442;
	wire [4-1:0] node7443;
	wire [4-1:0] node7445;
	wire [4-1:0] node7448;
	wire [4-1:0] node7449;
	wire [4-1:0] node7452;
	wire [4-1:0] node7453;
	wire [4-1:0] node7456;
	wire [4-1:0] node7459;
	wire [4-1:0] node7460;
	wire [4-1:0] node7463;
	wire [4-1:0] node7465;
	wire [4-1:0] node7468;
	wire [4-1:0] node7469;
	wire [4-1:0] node7470;
	wire [4-1:0] node7472;
	wire [4-1:0] node7475;
	wire [4-1:0] node7476;
	wire [4-1:0] node7480;
	wire [4-1:0] node7481;
	wire [4-1:0] node7482;
	wire [4-1:0] node7485;
	wire [4-1:0] node7488;
	wire [4-1:0] node7489;
	wire [4-1:0] node7490;
	wire [4-1:0] node7493;
	wire [4-1:0] node7496;
	wire [4-1:0] node7497;
	wire [4-1:0] node7500;
	wire [4-1:0] node7503;
	wire [4-1:0] node7504;
	wire [4-1:0] node7505;
	wire [4-1:0] node7506;
	wire [4-1:0] node7508;
	wire [4-1:0] node7512;
	wire [4-1:0] node7513;
	wire [4-1:0] node7515;
	wire [4-1:0] node7519;
	wire [4-1:0] node7520;
	wire [4-1:0] node7521;
	wire [4-1:0] node7524;
	wire [4-1:0] node7525;
	wire [4-1:0] node7528;
	wire [4-1:0] node7530;
	wire [4-1:0] node7533;
	wire [4-1:0] node7535;
	wire [4-1:0] node7538;
	wire [4-1:0] node7539;
	wire [4-1:0] node7540;
	wire [4-1:0] node7541;
	wire [4-1:0] node7542;
	wire [4-1:0] node7543;
	wire [4-1:0] node7544;
	wire [4-1:0] node7546;
	wire [4-1:0] node7549;
	wire [4-1:0] node7552;
	wire [4-1:0] node7553;
	wire [4-1:0] node7554;
	wire [4-1:0] node7555;
	wire [4-1:0] node7559;
	wire [4-1:0] node7561;
	wire [4-1:0] node7564;
	wire [4-1:0] node7565;
	wire [4-1:0] node7568;
	wire [4-1:0] node7571;
	wire [4-1:0] node7572;
	wire [4-1:0] node7573;
	wire [4-1:0] node7574;
	wire [4-1:0] node7578;
	wire [4-1:0] node7580;
	wire [4-1:0] node7583;
	wire [4-1:0] node7584;
	wire [4-1:0] node7586;
	wire [4-1:0] node7589;
	wire [4-1:0] node7590;
	wire [4-1:0] node7594;
	wire [4-1:0] node7595;
	wire [4-1:0] node7596;
	wire [4-1:0] node7597;
	wire [4-1:0] node7600;
	wire [4-1:0] node7602;
	wire [4-1:0] node7605;
	wire [4-1:0] node7606;
	wire [4-1:0] node7608;
	wire [4-1:0] node7611;
	wire [4-1:0] node7613;
	wire [4-1:0] node7616;
	wire [4-1:0] node7617;
	wire [4-1:0] node7619;
	wire [4-1:0] node7622;
	wire [4-1:0] node7623;
	wire [4-1:0] node7626;
	wire [4-1:0] node7628;
	wire [4-1:0] node7631;
	wire [4-1:0] node7632;
	wire [4-1:0] node7633;
	wire [4-1:0] node7634;
	wire [4-1:0] node7635;
	wire [4-1:0] node7636;
	wire [4-1:0] node7639;
	wire [4-1:0] node7642;
	wire [4-1:0] node7643;
	wire [4-1:0] node7646;
	wire [4-1:0] node7649;
	wire [4-1:0] node7650;
	wire [4-1:0] node7652;
	wire [4-1:0] node7655;
	wire [4-1:0] node7656;
	wire [4-1:0] node7660;
	wire [4-1:0] node7661;
	wire [4-1:0] node7662;
	wire [4-1:0] node7664;
	wire [4-1:0] node7667;
	wire [4-1:0] node7668;
	wire [4-1:0] node7672;
	wire [4-1:0] node7673;
	wire [4-1:0] node7675;
	wire [4-1:0] node7678;
	wire [4-1:0] node7680;
	wire [4-1:0] node7683;
	wire [4-1:0] node7684;
	wire [4-1:0] node7685;
	wire [4-1:0] node7686;
	wire [4-1:0] node7688;
	wire [4-1:0] node7691;
	wire [4-1:0] node7692;
	wire [4-1:0] node7695;
	wire [4-1:0] node7698;
	wire [4-1:0] node7699;
	wire [4-1:0] node7700;
	wire [4-1:0] node7704;
	wire [4-1:0] node7705;
	wire [4-1:0] node7708;
	wire [4-1:0] node7711;
	wire [4-1:0] node7712;
	wire [4-1:0] node7713;
	wire [4-1:0] node7714;
	wire [4-1:0] node7717;
	wire [4-1:0] node7720;
	wire [4-1:0] node7722;
	wire [4-1:0] node7725;
	wire [4-1:0] node7726;
	wire [4-1:0] node7729;
	wire [4-1:0] node7730;
	wire [4-1:0] node7734;
	wire [4-1:0] node7735;
	wire [4-1:0] node7736;
	wire [4-1:0] node7737;
	wire [4-1:0] node7738;
	wire [4-1:0] node7739;
	wire [4-1:0] node7742;
	wire [4-1:0] node7744;
	wire [4-1:0] node7747;
	wire [4-1:0] node7748;
	wire [4-1:0] node7751;
	wire [4-1:0] node7754;
	wire [4-1:0] node7755;
	wire [4-1:0] node7757;
	wire [4-1:0] node7760;
	wire [4-1:0] node7761;
	wire [4-1:0] node7764;
	wire [4-1:0] node7766;
	wire [4-1:0] node7769;
	wire [4-1:0] node7770;
	wire [4-1:0] node7771;
	wire [4-1:0] node7773;
	wire [4-1:0] node7776;
	wire [4-1:0] node7777;
	wire [4-1:0] node7778;
	wire [4-1:0] node7781;
	wire [4-1:0] node7784;
	wire [4-1:0] node7785;
	wire [4-1:0] node7788;
	wire [4-1:0] node7791;
	wire [4-1:0] node7792;
	wire [4-1:0] node7793;
	wire [4-1:0] node7796;
	wire [4-1:0] node7797;
	wire [4-1:0] node7801;
	wire [4-1:0] node7802;
	wire [4-1:0] node7806;
	wire [4-1:0] node7807;
	wire [4-1:0] node7808;
	wire [4-1:0] node7809;
	wire [4-1:0] node7811;
	wire [4-1:0] node7814;
	wire [4-1:0] node7815;
	wire [4-1:0] node7819;
	wire [4-1:0] node7820;
	wire [4-1:0] node7822;
	wire [4-1:0] node7825;
	wire [4-1:0] node7826;
	wire [4-1:0] node7829;
	wire [4-1:0] node7832;
	wire [4-1:0] node7833;
	wire [4-1:0] node7835;
	wire [4-1:0] node7837;
	wire [4-1:0] node7840;
	wire [4-1:0] node7842;
	wire [4-1:0] node7845;
	wire [4-1:0] node7846;
	wire [4-1:0] node7847;
	wire [4-1:0] node7848;
	wire [4-1:0] node7850;
	wire [4-1:0] node7851;
	wire [4-1:0] node7852;
	wire [4-1:0] node7853;
	wire [4-1:0] node7855;
	wire [4-1:0] node7856;
	wire [4-1:0] node7860;
	wire [4-1:0] node7862;
	wire [4-1:0] node7865;
	wire [4-1:0] node7867;
	wire [4-1:0] node7868;
	wire [4-1:0] node7870;
	wire [4-1:0] node7875;
	wire [4-1:0] node7876;
	wire [4-1:0] node7877;
	wire [4-1:0] node7878;
	wire [4-1:0] node7879;
	wire [4-1:0] node7881;
	wire [4-1:0] node7884;
	wire [4-1:0] node7885;
	wire [4-1:0] node7889;
	wire [4-1:0] node7890;
	wire [4-1:0] node7891;
	wire [4-1:0] node7892;
	wire [4-1:0] node7896;
	wire [4-1:0] node7898;
	wire [4-1:0] node7901;
	wire [4-1:0] node7904;
	wire [4-1:0] node7905;
	wire [4-1:0] node7906;
	wire [4-1:0] node7907;
	wire [4-1:0] node7910;
	wire [4-1:0] node7912;
	wire [4-1:0] node7916;
	wire [4-1:0] node7917;
	wire [4-1:0] node7919;
	wire [4-1:0] node7922;
	wire [4-1:0] node7923;
	wire [4-1:0] node7925;
	wire [4-1:0] node7929;
	wire [4-1:0] node7931;
	wire [4-1:0] node7932;
	wire [4-1:0] node7933;
	wire [4-1:0] node7934;
	wire [4-1:0] node7935;
	wire [4-1:0] node7941;
	wire [4-1:0] node7942;
	wire [4-1:0] node7944;
	wire [4-1:0] node7945;
	wire [4-1:0] node7949;
	wire [4-1:0] node7951;
	wire [4-1:0] node7954;
	wire [4-1:0] node7955;
	wire [4-1:0] node7956;
	wire [4-1:0] node7957;
	wire [4-1:0] node7958;
	wire [4-1:0] node7960;
	wire [4-1:0] node7961;
	wire [4-1:0] node7963;
	wire [4-1:0] node7967;
	wire [4-1:0] node7968;
	wire [4-1:0] node7970;
	wire [4-1:0] node7973;
	wire [4-1:0] node7974;
	wire [4-1:0] node7977;
	wire [4-1:0] node7980;
	wire [4-1:0] node7981;
	wire [4-1:0] node7982;
	wire [4-1:0] node7984;
	wire [4-1:0] node7987;
	wire [4-1:0] node7989;
	wire [4-1:0] node7992;
	wire [4-1:0] node7993;
	wire [4-1:0] node7995;
	wire [4-1:0] node7997;
	wire [4-1:0] node8000;
	wire [4-1:0] node8001;
	wire [4-1:0] node8004;
	wire [4-1:0] node8007;
	wire [4-1:0] node8008;
	wire [4-1:0] node8009;
	wire [4-1:0] node8010;
	wire [4-1:0] node8014;
	wire [4-1:0] node8015;
	wire [4-1:0] node8016;
	wire [4-1:0] node8020;
	wire [4-1:0] node8022;
	wire [4-1:0] node8025;
	wire [4-1:0] node8026;
	wire [4-1:0] node8028;
	wire [4-1:0] node8031;
	wire [4-1:0] node8032;
	wire [4-1:0] node8033;
	wire [4-1:0] node8037;
	wire [4-1:0] node8039;
	wire [4-1:0] node8042;
	wire [4-1:0] node8043;
	wire [4-1:0] node8044;
	wire [4-1:0] node8045;
	wire [4-1:0] node8047;
	wire [4-1:0] node8050;
	wire [4-1:0] node8052;
	wire [4-1:0] node8055;
	wire [4-1:0] node8056;
	wire [4-1:0] node8057;
	wire [4-1:0] node8059;
	wire [4-1:0] node8060;
	wire [4-1:0] node8064;
	wire [4-1:0] node8065;
	wire [4-1:0] node8069;
	wire [4-1:0] node8070;
	wire [4-1:0] node8073;
	wire [4-1:0] node8074;
	wire [4-1:0] node8076;
	wire [4-1:0] node8080;
	wire [4-1:0] node8081;
	wire [4-1:0] node8082;
	wire [4-1:0] node8083;
	wire [4-1:0] node8085;
	wire [4-1:0] node8088;
	wire [4-1:0] node8091;
	wire [4-1:0] node8092;
	wire [4-1:0] node8093;
	wire [4-1:0] node8097;
	wire [4-1:0] node8098;
	wire [4-1:0] node8100;
	wire [4-1:0] node8104;
	wire [4-1:0] node8105;
	wire [4-1:0] node8107;
	wire [4-1:0] node8110;
	wire [4-1:0] node8111;
	wire [4-1:0] node8116;
	wire [4-1:0] node8117;
	wire [4-1:0] node8118;
	wire [4-1:0] node8119;
	wire [4-1:0] node8120;
	wire [4-1:0] node8121;
	wire [4-1:0] node8122;
	wire [4-1:0] node8123;
	wire [4-1:0] node8124;
	wire [4-1:0] node8125;
	wire [4-1:0] node8128;
	wire [4-1:0] node8130;
	wire [4-1:0] node8133;
	wire [4-1:0] node8134;
	wire [4-1:0] node8137;
	wire [4-1:0] node8140;
	wire [4-1:0] node8141;
	wire [4-1:0] node8142;
	wire [4-1:0] node8144;
	wire [4-1:0] node8148;
	wire [4-1:0] node8151;
	wire [4-1:0] node8152;
	wire [4-1:0] node8154;
	wire [4-1:0] node8157;
	wire [4-1:0] node8158;
	wire [4-1:0] node8161;
	wire [4-1:0] node8163;
	wire [4-1:0] node8166;
	wire [4-1:0] node8167;
	wire [4-1:0] node8168;
	wire [4-1:0] node8169;
	wire [4-1:0] node8172;
	wire [4-1:0] node8173;
	wire [4-1:0] node8174;
	wire [4-1:0] node8177;
	wire [4-1:0] node8180;
	wire [4-1:0] node8181;
	wire [4-1:0] node8185;
	wire [4-1:0] node8186;
	wire [4-1:0] node8187;
	wire [4-1:0] node8191;
	wire [4-1:0] node8192;
	wire [4-1:0] node8194;
	wire [4-1:0] node8198;
	wire [4-1:0] node8199;
	wire [4-1:0] node8200;
	wire [4-1:0] node8201;
	wire [4-1:0] node8204;
	wire [4-1:0] node8207;
	wire [4-1:0] node8208;
	wire [4-1:0] node8211;
	wire [4-1:0] node8214;
	wire [4-1:0] node8215;
	wire [4-1:0] node8216;
	wire [4-1:0] node8218;
	wire [4-1:0] node8222;
	wire [4-1:0] node8225;
	wire [4-1:0] node8226;
	wire [4-1:0] node8227;
	wire [4-1:0] node8228;
	wire [4-1:0] node8230;
	wire [4-1:0] node8233;
	wire [4-1:0] node8234;
	wire [4-1:0] node8236;
	wire [4-1:0] node8239;
	wire [4-1:0] node8240;
	wire [4-1:0] node8241;
	wire [4-1:0] node8245;
	wire [4-1:0] node8248;
	wire [4-1:0] node8249;
	wire [4-1:0] node8250;
	wire [4-1:0] node8253;
	wire [4-1:0] node8256;
	wire [4-1:0] node8257;
	wire [4-1:0] node8259;
	wire [4-1:0] node8261;
	wire [4-1:0] node8264;
	wire [4-1:0] node8266;
	wire [4-1:0] node8270;
	wire [4-1:0] node8271;
	wire [4-1:0] node8272;
	wire [4-1:0] node8273;
	wire [4-1:0] node8274;
	wire [4-1:0] node8275;
	wire [4-1:0] node8277;
	wire [4-1:0] node8280;
	wire [4-1:0] node8281;
	wire [4-1:0] node8285;
	wire [4-1:0] node8286;
	wire [4-1:0] node8290;
	wire [4-1:0] node8291;
	wire [4-1:0] node8292;
	wire [4-1:0] node8293;
	wire [4-1:0] node8298;
	wire [4-1:0] node8299;
	wire [4-1:0] node8301;
	wire [4-1:0] node8304;
	wire [4-1:0] node8305;
	wire [4-1:0] node8309;
	wire [4-1:0] node8310;
	wire [4-1:0] node8311;
	wire [4-1:0] node8312;
	wire [4-1:0] node8313;
	wire [4-1:0] node8316;
	wire [4-1:0] node8319;
	wire [4-1:0] node8320;
	wire [4-1:0] node8323;
	wire [4-1:0] node8326;
	wire [4-1:0] node8328;
	wire [4-1:0] node8329;
	wire [4-1:0] node8333;
	wire [4-1:0] node8334;
	wire [4-1:0] node8335;
	wire [4-1:0] node8336;
	wire [4-1:0] node8338;
	wire [4-1:0] node8341;
	wire [4-1:0] node8342;
	wire [4-1:0] node8346;
	wire [4-1:0] node8347;
	wire [4-1:0] node8350;
	wire [4-1:0] node8352;
	wire [4-1:0] node8356;
	wire [4-1:0] node8357;
	wire [4-1:0] node8358;
	wire [4-1:0] node8359;
	wire [4-1:0] node8360;
	wire [4-1:0] node8361;
	wire [4-1:0] node8362;
	wire [4-1:0] node8365;
	wire [4-1:0] node8368;
	wire [4-1:0] node8370;
	wire [4-1:0] node8373;
	wire [4-1:0] node8374;
	wire [4-1:0] node8376;
	wire [4-1:0] node8379;
	wire [4-1:0] node8382;
	wire [4-1:0] node8383;
	wire [4-1:0] node8384;
	wire [4-1:0] node8388;
	wire [4-1:0] node8389;
	wire [4-1:0] node8392;
	wire [4-1:0] node8395;
	wire [4-1:0] node8396;
	wire [4-1:0] node8397;
	wire [4-1:0] node8401;
	wire [4-1:0] node8402;
	wire [4-1:0] node8404;
	wire [4-1:0] node8408;
	wire [4-1:0] node8409;
	wire [4-1:0] node8410;
	wire [4-1:0] node8411;
	wire [4-1:0] node8414;
	wire [4-1:0] node8415;
	wire [4-1:0] node8419;
	wire [4-1:0] node8420;
	wire [4-1:0] node8422;
	wire [4-1:0] node8425;
	wire [4-1:0] node8426;
	wire [4-1:0] node8430;
	wire [4-1:0] node8431;
	wire [4-1:0] node8433;
	wire [4-1:0] node8436;
	wire [4-1:0] node8437;
	wire [4-1:0] node8440;
	wire [4-1:0] node8443;
	wire [4-1:0] node8444;
	wire [4-1:0] node8445;
	wire [4-1:0] node8446;
	wire [4-1:0] node8447;
	wire [4-1:0] node8448;
	wire [4-1:0] node8449;
	wire [4-1:0] node8450;
	wire [4-1:0] node8453;
	wire [4-1:0] node8457;
	wire [4-1:0] node8458;
	wire [4-1:0] node8460;
	wire [4-1:0] node8463;
	wire [4-1:0] node8465;
	wire [4-1:0] node8468;
	wire [4-1:0] node8469;
	wire [4-1:0] node8470;
	wire [4-1:0] node8471;
	wire [4-1:0] node8474;
	wire [4-1:0] node8475;
	wire [4-1:0] node8478;
	wire [4-1:0] node8481;
	wire [4-1:0] node8482;
	wire [4-1:0] node8483;
	wire [4-1:0] node8488;
	wire [4-1:0] node8489;
	wire [4-1:0] node8492;
	wire [4-1:0] node8495;
	wire [4-1:0] node8496;
	wire [4-1:0] node8497;
	wire [4-1:0] node8498;
	wire [4-1:0] node8499;
	wire [4-1:0] node8503;
	wire [4-1:0] node8505;
	wire [4-1:0] node8506;
	wire [4-1:0] node8510;
	wire [4-1:0] node8511;
	wire [4-1:0] node8513;
	wire [4-1:0] node8514;
	wire [4-1:0] node8517;
	wire [4-1:0] node8520;
	wire [4-1:0] node8521;
	wire [4-1:0] node8525;
	wire [4-1:0] node8526;
	wire [4-1:0] node8527;
	wire [4-1:0] node8528;
	wire [4-1:0] node8531;
	wire [4-1:0] node8532;
	wire [4-1:0] node8536;
	wire [4-1:0] node8537;
	wire [4-1:0] node8538;
	wire [4-1:0] node8542;
	wire [4-1:0] node8545;
	wire [4-1:0] node8546;
	wire [4-1:0] node8547;
	wire [4-1:0] node8549;
	wire [4-1:0] node8553;
	wire [4-1:0] node8555;
	wire [4-1:0] node8556;
	wire [4-1:0] node8560;
	wire [4-1:0] node8561;
	wire [4-1:0] node8562;
	wire [4-1:0] node8563;
	wire [4-1:0] node8564;
	wire [4-1:0] node8565;
	wire [4-1:0] node8568;
	wire [4-1:0] node8571;
	wire [4-1:0] node8572;
	wire [4-1:0] node8573;
	wire [4-1:0] node8578;
	wire [4-1:0] node8579;
	wire [4-1:0] node8582;
	wire [4-1:0] node8583;
	wire [4-1:0] node8587;
	wire [4-1:0] node8588;
	wire [4-1:0] node8589;
	wire [4-1:0] node8591;
	wire [4-1:0] node8594;
	wire [4-1:0] node8596;
	wire [4-1:0] node8599;
	wire [4-1:0] node8600;
	wire [4-1:0] node8601;
	wire [4-1:0] node8602;
	wire [4-1:0] node8605;
	wire [4-1:0] node8608;
	wire [4-1:0] node8609;
	wire [4-1:0] node8612;
	wire [4-1:0] node8615;
	wire [4-1:0] node8616;
	wire [4-1:0] node8619;
	wire [4-1:0] node8622;
	wire [4-1:0] node8623;
	wire [4-1:0] node8624;
	wire [4-1:0] node8625;
	wire [4-1:0] node8626;
	wire [4-1:0] node8630;
	wire [4-1:0] node8631;
	wire [4-1:0] node8634;
	wire [4-1:0] node8637;
	wire [4-1:0] node8638;
	wire [4-1:0] node8642;
	wire [4-1:0] node8644;
	wire [4-1:0] node8645;
	wire [4-1:0] node8646;
	wire [4-1:0] node8651;
	wire [4-1:0] node8652;
	wire [4-1:0] node8653;
	wire [4-1:0] node8654;
	wire [4-1:0] node8655;
	wire [4-1:0] node8656;
	wire [4-1:0] node8659;
	wire [4-1:0] node8662;
	wire [4-1:0] node8664;
	wire [4-1:0] node8665;
	wire [4-1:0] node8666;
	wire [4-1:0] node8671;
	wire [4-1:0] node8672;
	wire [4-1:0] node8673;
	wire [4-1:0] node8674;
	wire [4-1:0] node8675;
	wire [4-1:0] node8678;
	wire [4-1:0] node8681;
	wire [4-1:0] node8682;
	wire [4-1:0] node8686;
	wire [4-1:0] node8687;
	wire [4-1:0] node8688;
	wire [4-1:0] node8691;
	wire [4-1:0] node8694;
	wire [4-1:0] node8697;
	wire [4-1:0] node8698;
	wire [4-1:0] node8701;
	wire [4-1:0] node8703;
	wire [4-1:0] node8704;
	wire [4-1:0] node8707;
	wire [4-1:0] node8710;
	wire [4-1:0] node8711;
	wire [4-1:0] node8712;
	wire [4-1:0] node8713;
	wire [4-1:0] node8714;
	wire [4-1:0] node8717;
	wire [4-1:0] node8718;
	wire [4-1:0] node8722;
	wire [4-1:0] node8723;
	wire [4-1:0] node8724;
	wire [4-1:0] node8729;
	wire [4-1:0] node8730;
	wire [4-1:0] node8733;
	wire [4-1:0] node8736;
	wire [4-1:0] node8737;
	wire [4-1:0] node8738;
	wire [4-1:0] node8739;
	wire [4-1:0] node8742;
	wire [4-1:0] node8745;
	wire [4-1:0] node8747;
	wire [4-1:0] node8750;
	wire [4-1:0] node8751;
	wire [4-1:0] node8752;
	wire [4-1:0] node8753;
	wire [4-1:0] node8756;
	wire [4-1:0] node8759;
	wire [4-1:0] node8761;
	wire [4-1:0] node8764;
	wire [4-1:0] node8767;
	wire [4-1:0] node8768;
	wire [4-1:0] node8769;
	wire [4-1:0] node8771;
	wire [4-1:0] node8772;
	wire [4-1:0] node8775;
	wire [4-1:0] node8777;
	wire [4-1:0] node8780;
	wire [4-1:0] node8781;
	wire [4-1:0] node8782;
	wire [4-1:0] node8785;
	wire [4-1:0] node8786;
	wire [4-1:0] node8789;
	wire [4-1:0] node8792;
	wire [4-1:0] node8793;
	wire [4-1:0] node8794;
	wire [4-1:0] node8797;
	wire [4-1:0] node8800;
	wire [4-1:0] node8801;
	wire [4-1:0] node8805;
	wire [4-1:0] node8806;
	wire [4-1:0] node8807;
	wire [4-1:0] node8809;
	wire [4-1:0] node8812;
	wire [4-1:0] node8813;
	wire [4-1:0] node8816;
	wire [4-1:0] node8820;
	wire [4-1:0] node8821;
	wire [4-1:0] node8822;
	wire [4-1:0] node8823;
	wire [4-1:0] node8824;
	wire [4-1:0] node8825;
	wire [4-1:0] node8826;
	wire [4-1:0] node8827;
	wire [4-1:0] node8828;
	wire [4-1:0] node8832;
	wire [4-1:0] node8833;
	wire [4-1:0] node8837;
	wire [4-1:0] node8838;
	wire [4-1:0] node8840;
	wire [4-1:0] node8843;
	wire [4-1:0] node8844;
	wire [4-1:0] node8845;
	wire [4-1:0] node8850;
	wire [4-1:0] node8851;
	wire [4-1:0] node8852;
	wire [4-1:0] node8853;
	wire [4-1:0] node8856;
	wire [4-1:0] node8859;
	wire [4-1:0] node8861;
	wire [4-1:0] node8862;
	wire [4-1:0] node8865;
	wire [4-1:0] node8868;
	wire [4-1:0] node8869;
	wire [4-1:0] node8871;
	wire [4-1:0] node8874;
	wire [4-1:0] node8875;
	wire [4-1:0] node8878;
	wire [4-1:0] node8881;
	wire [4-1:0] node8882;
	wire [4-1:0] node8883;
	wire [4-1:0] node8884;
	wire [4-1:0] node8886;
	wire [4-1:0] node8889;
	wire [4-1:0] node8891;
	wire [4-1:0] node8894;
	wire [4-1:0] node8895;
	wire [4-1:0] node8897;
	wire [4-1:0] node8900;
	wire [4-1:0] node8901;
	wire [4-1:0] node8905;
	wire [4-1:0] node8906;
	wire [4-1:0] node8907;
	wire [4-1:0] node8909;
	wire [4-1:0] node8911;
	wire [4-1:0] node8914;
	wire [4-1:0] node8917;
	wire [4-1:0] node8918;
	wire [4-1:0] node8921;
	wire [4-1:0] node8922;
	wire [4-1:0] node8926;
	wire [4-1:0] node8927;
	wire [4-1:0] node8928;
	wire [4-1:0] node8929;
	wire [4-1:0] node8930;
	wire [4-1:0] node8931;
	wire [4-1:0] node8932;
	wire [4-1:0] node8937;
	wire [4-1:0] node8938;
	wire [4-1:0] node8941;
	wire [4-1:0] node8943;
	wire [4-1:0] node8946;
	wire [4-1:0] node8947;
	wire [4-1:0] node8949;
	wire [4-1:0] node8951;
	wire [4-1:0] node8954;
	wire [4-1:0] node8955;
	wire [4-1:0] node8956;
	wire [4-1:0] node8960;
	wire [4-1:0] node8963;
	wire [4-1:0] node8964;
	wire [4-1:0] node8965;
	wire [4-1:0] node8966;
	wire [4-1:0] node8967;
	wire [4-1:0] node8970;
	wire [4-1:0] node8973;
	wire [4-1:0] node8975;
	wire [4-1:0] node8978;
	wire [4-1:0] node8979;
	wire [4-1:0] node8980;
	wire [4-1:0] node8984;
	wire [4-1:0] node8985;
	wire [4-1:0] node8989;
	wire [4-1:0] node8990;
	wire [4-1:0] node8991;
	wire [4-1:0] node8994;
	wire [4-1:0] node8996;
	wire [4-1:0] node8999;
	wire [4-1:0] node9001;
	wire [4-1:0] node9003;
	wire [4-1:0] node9006;
	wire [4-1:0] node9007;
	wire [4-1:0] node9008;
	wire [4-1:0] node9010;
	wire [4-1:0] node9013;
	wire [4-1:0] node9014;
	wire [4-1:0] node9017;
	wire [4-1:0] node9018;
	wire [4-1:0] node9022;
	wire [4-1:0] node9023;
	wire [4-1:0] node9024;
	wire [4-1:0] node9025;
	wire [4-1:0] node9028;
	wire [4-1:0] node9031;
	wire [4-1:0] node9032;
	wire [4-1:0] node9035;
	wire [4-1:0] node9038;
	wire [4-1:0] node9039;
	wire [4-1:0] node9040;
	wire [4-1:0] node9043;
	wire [4-1:0] node9046;
	wire [4-1:0] node9047;
	wire [4-1:0] node9050;
	wire [4-1:0] node9053;
	wire [4-1:0] node9054;
	wire [4-1:0] node9055;
	wire [4-1:0] node9056;
	wire [4-1:0] node9057;
	wire [4-1:0] node9058;
	wire [4-1:0] node9059;
	wire [4-1:0] node9061;
	wire [4-1:0] node9065;
	wire [4-1:0] node9067;
	wire [4-1:0] node9068;
	wire [4-1:0] node9071;
	wire [4-1:0] node9074;
	wire [4-1:0] node9075;
	wire [4-1:0] node9076;
	wire [4-1:0] node9077;
	wire [4-1:0] node9081;
	wire [4-1:0] node9083;
	wire [4-1:0] node9086;
	wire [4-1:0] node9087;
	wire [4-1:0] node9090;
	wire [4-1:0] node9093;
	wire [4-1:0] node9094;
	wire [4-1:0] node9095;
	wire [4-1:0] node9096;
	wire [4-1:0] node9098;
	wire [4-1:0] node9101;
	wire [4-1:0] node9104;
	wire [4-1:0] node9106;
	wire [4-1:0] node9108;
	wire [4-1:0] node9111;
	wire [4-1:0] node9112;
	wire [4-1:0] node9113;
	wire [4-1:0] node9114;
	wire [4-1:0] node9117;
	wire [4-1:0] node9120;
	wire [4-1:0] node9123;
	wire [4-1:0] node9126;
	wire [4-1:0] node9127;
	wire [4-1:0] node9128;
	wire [4-1:0] node9130;
	wire [4-1:0] node9133;
	wire [4-1:0] node9134;
	wire [4-1:0] node9135;
	wire [4-1:0] node9138;
	wire [4-1:0] node9139;
	wire [4-1:0] node9143;
	wire [4-1:0] node9146;
	wire [4-1:0] node9147;
	wire [4-1:0] node9148;
	wire [4-1:0] node9149;
	wire [4-1:0] node9153;
	wire [4-1:0] node9154;
	wire [4-1:0] node9155;
	wire [4-1:0] node9159;
	wire [4-1:0] node9162;
	wire [4-1:0] node9163;
	wire [4-1:0] node9165;
	wire [4-1:0] node9167;
	wire [4-1:0] node9170;
	wire [4-1:0] node9171;
	wire [4-1:0] node9175;
	wire [4-1:0] node9176;
	wire [4-1:0] node9177;
	wire [4-1:0] node9179;
	wire [4-1:0] node9180;
	wire [4-1:0] node9183;
	wire [4-1:0] node9184;
	wire [4-1:0] node9188;
	wire [4-1:0] node9189;
	wire [4-1:0] node9191;
	wire [4-1:0] node9192;
	wire [4-1:0] node9194;
	wire [4-1:0] node9197;
	wire [4-1:0] node9199;
	wire [4-1:0] node9202;
	wire [4-1:0] node9203;
	wire [4-1:0] node9204;
	wire [4-1:0] node9208;
	wire [4-1:0] node9209;
	wire [4-1:0] node9212;
	wire [4-1:0] node9215;
	wire [4-1:0] node9216;
	wire [4-1:0] node9217;
	wire [4-1:0] node9218;
	wire [4-1:0] node9219;
	wire [4-1:0] node9224;
	wire [4-1:0] node9225;
	wire [4-1:0] node9226;
	wire [4-1:0] node9230;
	wire [4-1:0] node9231;
	wire [4-1:0] node9236;
	wire [4-1:0] node9237;
	wire [4-1:0] node9238;
	wire [4-1:0] node9239;
	wire [4-1:0] node9240;
	wire [4-1:0] node9241;
	wire [4-1:0] node9242;
	wire [4-1:0] node9243;
	wire [4-1:0] node9245;
	wire [4-1:0] node9248;
	wire [4-1:0] node9249;
	wire [4-1:0] node9253;
	wire [4-1:0] node9254;
	wire [4-1:0] node9257;
	wire [4-1:0] node9260;
	wire [4-1:0] node9261;
	wire [4-1:0] node9262;
	wire [4-1:0] node9264;
	wire [4-1:0] node9269;
	wire [4-1:0] node9270;
	wire [4-1:0] node9271;
	wire [4-1:0] node9272;
	wire [4-1:0] node9276;
	wire [4-1:0] node9278;
	wire [4-1:0] node9279;
	wire [4-1:0] node9283;
	wire [4-1:0] node9284;
	wire [4-1:0] node9285;
	wire [4-1:0] node9289;
	wire [4-1:0] node9290;
	wire [4-1:0] node9294;
	wire [4-1:0] node9295;
	wire [4-1:0] node9296;
	wire [4-1:0] node9297;
	wire [4-1:0] node9298;
	wire [4-1:0] node9301;
	wire [4-1:0] node9304;
	wire [4-1:0] node9305;
	wire [4-1:0] node9306;
	wire [4-1:0] node9311;
	wire [4-1:0] node9312;
	wire [4-1:0] node9314;
	wire [4-1:0] node9315;
	wire [4-1:0] node9319;
	wire [4-1:0] node9320;
	wire [4-1:0] node9323;
	wire [4-1:0] node9324;
	wire [4-1:0] node9328;
	wire [4-1:0] node9329;
	wire [4-1:0] node9330;
	wire [4-1:0] node9331;
	wire [4-1:0] node9332;
	wire [4-1:0] node9337;
	wire [4-1:0] node9338;
	wire [4-1:0] node9341;
	wire [4-1:0] node9344;
	wire [4-1:0] node9345;
	wire [4-1:0] node9346;
	wire [4-1:0] node9349;
	wire [4-1:0] node9352;
	wire [4-1:0] node9353;
	wire [4-1:0] node9355;
	wire [4-1:0] node9359;
	wire [4-1:0] node9360;
	wire [4-1:0] node9361;
	wire [4-1:0] node9362;
	wire [4-1:0] node9363;
	wire [4-1:0] node9365;
	wire [4-1:0] node9368;
	wire [4-1:0] node9369;
	wire [4-1:0] node9372;
	wire [4-1:0] node9373;
	wire [4-1:0] node9377;
	wire [4-1:0] node9378;
	wire [4-1:0] node9381;
	wire [4-1:0] node9382;
	wire [4-1:0] node9383;
	wire [4-1:0] node9387;
	wire [4-1:0] node9390;
	wire [4-1:0] node9391;
	wire [4-1:0] node9392;
	wire [4-1:0] node9393;
	wire [4-1:0] node9394;
	wire [4-1:0] node9398;
	wire [4-1:0] node9401;
	wire [4-1:0] node9403;
	wire [4-1:0] node9406;
	wire [4-1:0] node9407;
	wire [4-1:0] node9408;
	wire [4-1:0] node9412;
	wire [4-1:0] node9413;
	wire [4-1:0] node9416;
	wire [4-1:0] node9418;
	wire [4-1:0] node9421;
	wire [4-1:0] node9422;
	wire [4-1:0] node9423;
	wire [4-1:0] node9424;
	wire [4-1:0] node9425;
	wire [4-1:0] node9429;
	wire [4-1:0] node9430;
	wire [4-1:0] node9434;
	wire [4-1:0] node9436;
	wire [4-1:0] node9438;
	wire [4-1:0] node9442;
	wire [4-1:0] node9443;
	wire [4-1:0] node9444;
	wire [4-1:0] node9445;
	wire [4-1:0] node9446;
	wire [4-1:0] node9447;
	wire [4-1:0] node9450;
	wire [4-1:0] node9451;
	wire [4-1:0] node9455;
	wire [4-1:0] node9456;
	wire [4-1:0] node9458;
	wire [4-1:0] node9459;
	wire [4-1:0] node9462;
	wire [4-1:0] node9466;
	wire [4-1:0] node9467;
	wire [4-1:0] node9468;
	wire [4-1:0] node9470;
	wire [4-1:0] node9471;
	wire [4-1:0] node9474;
	wire [4-1:0] node9477;
	wire [4-1:0] node9478;
	wire [4-1:0] node9479;
	wire [4-1:0] node9483;
	wire [4-1:0] node9484;
	wire [4-1:0] node9488;
	wire [4-1:0] node9489;
	wire [4-1:0] node9490;
	wire [4-1:0] node9494;
	wire [4-1:0] node9495;
	wire [4-1:0] node9497;
	wire [4-1:0] node9500;
	wire [4-1:0] node9503;
	wire [4-1:0] node9504;
	wire [4-1:0] node9505;
	wire [4-1:0] node9506;
	wire [4-1:0] node9507;
	wire [4-1:0] node9510;
	wire [4-1:0] node9511;
	wire [4-1:0] node9515;
	wire [4-1:0] node9516;
	wire [4-1:0] node9520;
	wire [4-1:0] node9521;
	wire [4-1:0] node9522;
	wire [4-1:0] node9523;
	wire [4-1:0] node9528;
	wire [4-1:0] node9530;
	wire [4-1:0] node9531;
	wire [4-1:0] node9536;
	wire [4-1:0] node9537;
	wire [4-1:0] node9538;
	wire [4-1:0] node9539;
	wire [4-1:0] node9541;
	wire [4-1:0] node9542;
	wire [4-1:0] node9544;
	wire [4-1:0] node9547;
	wire [4-1:0] node9550;
	wire [4-1:0] node9551;
	wire [4-1:0] node9552;
	wire [4-1:0] node9554;
	wire [4-1:0] node9558;
	wire [4-1:0] node9559;
	wire [4-1:0] node9560;
	wire [4-1:0] node9567;
	wire [4-1:0] node9568;
	wire [4-1:0] node9569;
	wire [4-1:0] node9570;
	wire [4-1:0] node9571;
	wire [4-1:0] node9573;
	wire [4-1:0] node9574;
	wire [4-1:0] node9575;
	wire [4-1:0] node9577;
	wire [4-1:0] node9578;
	wire [4-1:0] node9579;
	wire [4-1:0] node9581;
	wire [4-1:0] node9582;
	wire [4-1:0] node9586;
	wire [4-1:0] node9587;
	wire [4-1:0] node9591;
	wire [4-1:0] node9593;
	wire [4-1:0] node9594;
	wire [4-1:0] node9596;
	wire [4-1:0] node9599;
	wire [4-1:0] node9602;
	wire [4-1:0] node9603;
	wire [4-1:0] node9604;
	wire [4-1:0] node9605;
	wire [4-1:0] node9606;
	wire [4-1:0] node9608;
	wire [4-1:0] node9611;
	wire [4-1:0] node9614;
	wire [4-1:0] node9616;
	wire [4-1:0] node9618;
	wire [4-1:0] node9621;
	wire [4-1:0] node9622;
	wire [4-1:0] node9623;
	wire [4-1:0] node9628;
	wire [4-1:0] node9629;
	wire [4-1:0] node9630;
	wire [4-1:0] node9631;
	wire [4-1:0] node9635;
	wire [4-1:0] node9638;
	wire [4-1:0] node9639;
	wire [4-1:0] node9641;
	wire [4-1:0] node9644;
	wire [4-1:0] node9647;
	wire [4-1:0] node9649;
	wire [4-1:0] node9651;
	wire [4-1:0] node9652;
	wire [4-1:0] node9653;
	wire [4-1:0] node9655;
	wire [4-1:0] node9656;
	wire [4-1:0] node9660;
	wire [4-1:0] node9662;
	wire [4-1:0] node9665;
	wire [4-1:0] node9667;
	wire [4-1:0] node9669;
	wire [4-1:0] node9671;
	wire [4-1:0] node9674;
	wire [4-1:0] node9675;
	wire [4-1:0] node9676;
	wire [4-1:0] node9677;
	wire [4-1:0] node9678;
	wire [4-1:0] node9679;
	wire [4-1:0] node9680;
	wire [4-1:0] node9681;
	wire [4-1:0] node9685;
	wire [4-1:0] node9687;
	wire [4-1:0] node9690;
	wire [4-1:0] node9691;
	wire [4-1:0] node9692;
	wire [4-1:0] node9694;
	wire [4-1:0] node9698;
	wire [4-1:0] node9700;
	wire [4-1:0] node9703;
	wire [4-1:0] node9704;
	wire [4-1:0] node9705;
	wire [4-1:0] node9706;
	wire [4-1:0] node9708;
	wire [4-1:0] node9711;
	wire [4-1:0] node9714;
	wire [4-1:0] node9715;
	wire [4-1:0] node9716;
	wire [4-1:0] node9721;
	wire [4-1:0] node9722;
	wire [4-1:0] node9723;
	wire [4-1:0] node9727;
	wire [4-1:0] node9729;
	wire [4-1:0] node9732;
	wire [4-1:0] node9733;
	wire [4-1:0] node9734;
	wire [4-1:0] node9735;
	wire [4-1:0] node9736;
	wire [4-1:0] node9740;
	wire [4-1:0] node9741;
	wire [4-1:0] node9743;
	wire [4-1:0] node9746;
	wire [4-1:0] node9747;
	wire [4-1:0] node9751;
	wire [4-1:0] node9752;
	wire [4-1:0] node9753;
	wire [4-1:0] node9757;
	wire [4-1:0] node9758;
	wire [4-1:0] node9760;
	wire [4-1:0] node9764;
	wire [4-1:0] node9765;
	wire [4-1:0] node9766;
	wire [4-1:0] node9767;
	wire [4-1:0] node9770;
	wire [4-1:0] node9772;
	wire [4-1:0] node9775;
	wire [4-1:0] node9777;
	wire [4-1:0] node9779;
	wire [4-1:0] node9782;
	wire [4-1:0] node9783;
	wire [4-1:0] node9785;
	wire [4-1:0] node9788;
	wire [4-1:0] node9789;
	wire [4-1:0] node9793;
	wire [4-1:0] node9794;
	wire [4-1:0] node9795;
	wire [4-1:0] node9796;
	wire [4-1:0] node9798;
	wire [4-1:0] node9799;
	wire [4-1:0] node9803;
	wire [4-1:0] node9804;
	wire [4-1:0] node9808;
	wire [4-1:0] node9809;
	wire [4-1:0] node9810;
	wire [4-1:0] node9814;
	wire [4-1:0] node9817;
	wire [4-1:0] node9818;
	wire [4-1:0] node9819;
	wire [4-1:0] node9820;
	wire [4-1:0] node9821;
	wire [4-1:0] node9825;
	wire [4-1:0] node9827;
	wire [4-1:0] node9830;
	wire [4-1:0] node9831;
	wire [4-1:0] node9832;
	wire [4-1:0] node9836;
	wire [4-1:0] node9838;
	wire [4-1:0] node9841;
	wire [4-1:0] node9842;
	wire [4-1:0] node9844;
	wire [4-1:0] node9847;
	wire [4-1:0] node9849;
	wire [4-1:0] node9852;
	wire [4-1:0] node9853;
	wire [4-1:0] node9854;
	wire [4-1:0] node9855;
	wire [4-1:0] node9856;
	wire [4-1:0] node9857;
	wire [4-1:0] node9860;
	wire [4-1:0] node9861;
	wire [4-1:0] node9864;
	wire [4-1:0] node9865;
	wire [4-1:0] node9869;
	wire [4-1:0] node9870;
	wire [4-1:0] node9871;
	wire [4-1:0] node9875;
	wire [4-1:0] node9877;
	wire [4-1:0] node9880;
	wire [4-1:0] node9881;
	wire [4-1:0] node9882;
	wire [4-1:0] node9883;
	wire [4-1:0] node9887;
	wire [4-1:0] node9890;
	wire [4-1:0] node9891;
	wire [4-1:0] node9892;
	wire [4-1:0] node9893;
	wire [4-1:0] node9898;
	wire [4-1:0] node9899;
	wire [4-1:0] node9900;
	wire [4-1:0] node9905;
	wire [4-1:0] node9906;
	wire [4-1:0] node9907;
	wire [4-1:0] node9908;
	wire [4-1:0] node9910;
	wire [4-1:0] node9913;
	wire [4-1:0] node9916;
	wire [4-1:0] node9917;
	wire [4-1:0] node9918;
	wire [4-1:0] node9921;
	wire [4-1:0] node9922;
	wire [4-1:0] node9926;
	wire [4-1:0] node9928;
	wire [4-1:0] node9931;
	wire [4-1:0] node9932;
	wire [4-1:0] node9933;
	wire [4-1:0] node9934;
	wire [4-1:0] node9937;
	wire [4-1:0] node9940;
	wire [4-1:0] node9942;
	wire [4-1:0] node9943;
	wire [4-1:0] node9946;
	wire [4-1:0] node9949;
	wire [4-1:0] node9950;
	wire [4-1:0] node9952;
	wire [4-1:0] node9955;
	wire [4-1:0] node9957;
	wire [4-1:0] node9960;
	wire [4-1:0] node9961;
	wire [4-1:0] node9962;
	wire [4-1:0] node9963;
	wire [4-1:0] node9964;
	wire [4-1:0] node9967;
	wire [4-1:0] node9969;
	wire [4-1:0] node9972;
	wire [4-1:0] node9974;
	wire [4-1:0] node9977;
	wire [4-1:0] node9978;
	wire [4-1:0] node9979;
	wire [4-1:0] node9983;
	wire [4-1:0] node9984;
	wire [4-1:0] node9985;
	wire [4-1:0] node9989;
	wire [4-1:0] node9990;
	wire [4-1:0] node9994;
	wire [4-1:0] node9995;
	wire [4-1:0] node9996;
	wire [4-1:0] node9997;
	wire [4-1:0] node9998;
	wire [4-1:0] node10002;
	wire [4-1:0] node10003;
	wire [4-1:0] node10007;
	wire [4-1:0] node10008;
	wire [4-1:0] node10009;
	wire [4-1:0] node10013;
	wire [4-1:0] node10014;
	wire [4-1:0] node10018;
	wire [4-1:0] node10019;
	wire [4-1:0] node10021;
	wire [4-1:0] node10024;
	wire [4-1:0] node10026;
	wire [4-1:0] node10029;
	wire [4-1:0] node10031;
	wire [4-1:0] node10033;
	wire [4-1:0] node10034;
	wire [4-1:0] node10036;
	wire [4-1:0] node10037;
	wire [4-1:0] node10038;
	wire [4-1:0] node10039;
	wire [4-1:0] node10040;
	wire [4-1:0] node10045;
	wire [4-1:0] node10047;
	wire [4-1:0] node10048;
	wire [4-1:0] node10049;
	wire [4-1:0] node10052;
	wire [4-1:0] node10055;
	wire [4-1:0] node10057;
	wire [4-1:0] node10061;
	wire [4-1:0] node10062;
	wire [4-1:0] node10063;
	wire [4-1:0] node10064;
	wire [4-1:0] node10065;
	wire [4-1:0] node10066;
	wire [4-1:0] node10070;
	wire [4-1:0] node10072;
	wire [4-1:0] node10074;
	wire [4-1:0] node10077;
	wire [4-1:0] node10078;
	wire [4-1:0] node10080;
	wire [4-1:0] node10083;
	wire [4-1:0] node10085;
	wire [4-1:0] node10088;
	wire [4-1:0] node10089;
	wire [4-1:0] node10090;
	wire [4-1:0] node10092;
	wire [4-1:0] node10095;
	wire [4-1:0] node10096;
	wire [4-1:0] node10100;
	wire [4-1:0] node10101;
	wire [4-1:0] node10103;
	wire [4-1:0] node10106;
	wire [4-1:0] node10107;
	wire [4-1:0] node10108;
	wire [4-1:0] node10112;
	wire [4-1:0] node10114;
	wire [4-1:0] node10117;
	wire [4-1:0] node10119;
	wire [4-1:0] node10120;
	wire [4-1:0] node10121;
	wire [4-1:0] node10123;
	wire [4-1:0] node10124;
	wire [4-1:0] node10128;
	wire [4-1:0] node10129;
	wire [4-1:0] node10133;
	wire [4-1:0] node10135;
	wire [4-1:0] node10136;
	wire [4-1:0] node10139;
	wire [4-1:0] node10140;
	wire [4-1:0] node10144;
	wire [4-1:0] node10145;
	wire [4-1:0] node10146;
	wire [4-1:0] node10147;
	wire [4-1:0] node10148;
	wire [4-1:0] node10149;
	wire [4-1:0] node10150;
	wire [4-1:0] node10151;
	wire [4-1:0] node10152;
	wire [4-1:0] node10156;
	wire [4-1:0] node10157;
	wire [4-1:0] node10158;
	wire [4-1:0] node10160;
	wire [4-1:0] node10163;
	wire [4-1:0] node10166;
	wire [4-1:0] node10167;
	wire [4-1:0] node10171;
	wire [4-1:0] node10173;
	wire [4-1:0] node10176;
	wire [4-1:0] node10177;
	wire [4-1:0] node10178;
	wire [4-1:0] node10179;
	wire [4-1:0] node10182;
	wire [4-1:0] node10184;
	wire [4-1:0] node10186;
	wire [4-1:0] node10189;
	wire [4-1:0] node10190;
	wire [4-1:0] node10191;
	wire [4-1:0] node10193;
	wire [4-1:0] node10196;
	wire [4-1:0] node10199;
	wire [4-1:0] node10200;
	wire [4-1:0] node10204;
	wire [4-1:0] node10205;
	wire [4-1:0] node10206;
	wire [4-1:0] node10208;
	wire [4-1:0] node10211;
	wire [4-1:0] node10213;
	wire [4-1:0] node10214;
	wire [4-1:0] node10217;
	wire [4-1:0] node10220;
	wire [4-1:0] node10221;
	wire [4-1:0] node10222;
	wire [4-1:0] node10224;
	wire [4-1:0] node10227;
	wire [4-1:0] node10228;
	wire [4-1:0] node10231;
	wire [4-1:0] node10234;
	wire [4-1:0] node10236;
	wire [4-1:0] node10239;
	wire [4-1:0] node10240;
	wire [4-1:0] node10241;
	wire [4-1:0] node10242;
	wire [4-1:0] node10243;
	wire [4-1:0] node10244;
	wire [4-1:0] node10246;
	wire [4-1:0] node10249;
	wire [4-1:0] node10252;
	wire [4-1:0] node10253;
	wire [4-1:0] node10255;
	wire [4-1:0] node10259;
	wire [4-1:0] node10260;
	wire [4-1:0] node10264;
	wire [4-1:0] node10265;
	wire [4-1:0] node10266;
	wire [4-1:0] node10267;
	wire [4-1:0] node10270;
	wire [4-1:0] node10273;
	wire [4-1:0] node10275;
	wire [4-1:0] node10278;
	wire [4-1:0] node10279;
	wire [4-1:0] node10280;
	wire [4-1:0] node10281;
	wire [4-1:0] node10284;
	wire [4-1:0] node10287;
	wire [4-1:0] node10288;
	wire [4-1:0] node10292;
	wire [4-1:0] node10293;
	wire [4-1:0] node10294;
	wire [4-1:0] node10298;
	wire [4-1:0] node10301;
	wire [4-1:0] node10302;
	wire [4-1:0] node10303;
	wire [4-1:0] node10305;
	wire [4-1:0] node10308;
	wire [4-1:0] node10309;
	wire [4-1:0] node10310;
	wire [4-1:0] node10313;
	wire [4-1:0] node10314;
	wire [4-1:0] node10319;
	wire [4-1:0] node10320;
	wire [4-1:0] node10321;
	wire [4-1:0] node10323;
	wire [4-1:0] node10326;
	wire [4-1:0] node10329;
	wire [4-1:0] node10330;
	wire [4-1:0] node10331;
	wire [4-1:0] node10332;
	wire [4-1:0] node10335;
	wire [4-1:0] node10338;
	wire [4-1:0] node10339;
	wire [4-1:0] node10342;
	wire [4-1:0] node10345;
	wire [4-1:0] node10346;
	wire [4-1:0] node10348;
	wire [4-1:0] node10351;
	wire [4-1:0] node10354;
	wire [4-1:0] node10355;
	wire [4-1:0] node10356;
	wire [4-1:0] node10357;
	wire [4-1:0] node10358;
	wire [4-1:0] node10360;
	wire [4-1:0] node10363;
	wire [4-1:0] node10364;
	wire [4-1:0] node10365;
	wire [4-1:0] node10369;
	wire [4-1:0] node10372;
	wire [4-1:0] node10373;
	wire [4-1:0] node10374;
	wire [4-1:0] node10376;
	wire [4-1:0] node10377;
	wire [4-1:0] node10381;
	wire [4-1:0] node10382;
	wire [4-1:0] node10386;
	wire [4-1:0] node10387;
	wire [4-1:0] node10389;
	wire [4-1:0] node10391;
	wire [4-1:0] node10394;
	wire [4-1:0] node10396;
	wire [4-1:0] node10399;
	wire [4-1:0] node10400;
	wire [4-1:0] node10401;
	wire [4-1:0] node10402;
	wire [4-1:0] node10403;
	wire [4-1:0] node10404;
	wire [4-1:0] node10408;
	wire [4-1:0] node10409;
	wire [4-1:0] node10413;
	wire [4-1:0] node10414;
	wire [4-1:0] node10417;
	wire [4-1:0] node10420;
	wire [4-1:0] node10421;
	wire [4-1:0] node10422;
	wire [4-1:0] node10423;
	wire [4-1:0] node10428;
	wire [4-1:0] node10429;
	wire [4-1:0] node10432;
	wire [4-1:0] node10435;
	wire [4-1:0] node10436;
	wire [4-1:0] node10437;
	wire [4-1:0] node10439;
	wire [4-1:0] node10440;
	wire [4-1:0] node10444;
	wire [4-1:0] node10445;
	wire [4-1:0] node10449;
	wire [4-1:0] node10450;
	wire [4-1:0] node10452;
	wire [4-1:0] node10455;
	wire [4-1:0] node10456;
	wire [4-1:0] node10458;
	wire [4-1:0] node10462;
	wire [4-1:0] node10463;
	wire [4-1:0] node10464;
	wire [4-1:0] node10465;
	wire [4-1:0] node10466;
	wire [4-1:0] node10467;
	wire [4-1:0] node10469;
	wire [4-1:0] node10472;
	wire [4-1:0] node10474;
	wire [4-1:0] node10477;
	wire [4-1:0] node10480;
	wire [4-1:0] node10481;
	wire [4-1:0] node10484;
	wire [4-1:0] node10485;
	wire [4-1:0] node10487;
	wire [4-1:0] node10490;
	wire [4-1:0] node10493;
	wire [4-1:0] node10494;
	wire [4-1:0] node10495;
	wire [4-1:0] node10496;
	wire [4-1:0] node10499;
	wire [4-1:0] node10500;
	wire [4-1:0] node10504;
	wire [4-1:0] node10505;
	wire [4-1:0] node10507;
	wire [4-1:0] node10510;
	wire [4-1:0] node10511;
	wire [4-1:0] node10514;
	wire [4-1:0] node10517;
	wire [4-1:0] node10518;
	wire [4-1:0] node10519;
	wire [4-1:0] node10523;
	wire [4-1:0] node10525;
	wire [4-1:0] node10527;
	wire [4-1:0] node10530;
	wire [4-1:0] node10531;
	wire [4-1:0] node10532;
	wire [4-1:0] node10533;
	wire [4-1:0] node10535;
	wire [4-1:0] node10538;
	wire [4-1:0] node10541;
	wire [4-1:0] node10543;
	wire [4-1:0] node10544;
	wire [4-1:0] node10547;
	wire [4-1:0] node10550;
	wire [4-1:0] node10551;
	wire [4-1:0] node10552;
	wire [4-1:0] node10554;
	wire [4-1:0] node10557;
	wire [4-1:0] node10558;
	wire [4-1:0] node10559;
	wire [4-1:0] node10563;
	wire [4-1:0] node10565;
	wire [4-1:0] node10568;
	wire [4-1:0] node10569;
	wire [4-1:0] node10571;
	wire [4-1:0] node10573;
	wire [4-1:0] node10576;
	wire [4-1:0] node10579;
	wire [4-1:0] node10580;
	wire [4-1:0] node10581;
	wire [4-1:0] node10582;
	wire [4-1:0] node10583;
	wire [4-1:0] node10584;
	wire [4-1:0] node10585;
	wire [4-1:0] node10587;
	wire [4-1:0] node10590;
	wire [4-1:0] node10593;
	wire [4-1:0] node10594;
	wire [4-1:0] node10595;
	wire [4-1:0] node10598;
	wire [4-1:0] node10600;
	wire [4-1:0] node10603;
	wire [4-1:0] node10604;
	wire [4-1:0] node10608;
	wire [4-1:0] node10609;
	wire [4-1:0] node10610;
	wire [4-1:0] node10611;
	wire [4-1:0] node10616;
	wire [4-1:0] node10617;
	wire [4-1:0] node10618;
	wire [4-1:0] node10622;
	wire [4-1:0] node10624;
	wire [4-1:0] node10627;
	wire [4-1:0] node10628;
	wire [4-1:0] node10629;
	wire [4-1:0] node10630;
	wire [4-1:0] node10632;
	wire [4-1:0] node10635;
	wire [4-1:0] node10636;
	wire [4-1:0] node10638;
	wire [4-1:0] node10642;
	wire [4-1:0] node10643;
	wire [4-1:0] node10644;
	wire [4-1:0] node10648;
	wire [4-1:0] node10649;
	wire [4-1:0] node10650;
	wire [4-1:0] node10655;
	wire [4-1:0] node10656;
	wire [4-1:0] node10657;
	wire [4-1:0] node10658;
	wire [4-1:0] node10661;
	wire [4-1:0] node10662;
	wire [4-1:0] node10666;
	wire [4-1:0] node10667;
	wire [4-1:0] node10668;
	wire [4-1:0] node10673;
	wire [4-1:0] node10674;
	wire [4-1:0] node10675;
	wire [4-1:0] node10679;
	wire [4-1:0] node10680;
	wire [4-1:0] node10684;
	wire [4-1:0] node10685;
	wire [4-1:0] node10686;
	wire [4-1:0] node10687;
	wire [4-1:0] node10688;
	wire [4-1:0] node10691;
	wire [4-1:0] node10694;
	wire [4-1:0] node10695;
	wire [4-1:0] node10696;
	wire [4-1:0] node10699;
	wire [4-1:0] node10700;
	wire [4-1:0] node10703;
	wire [4-1:0] node10706;
	wire [4-1:0] node10707;
	wire [4-1:0] node10710;
	wire [4-1:0] node10713;
	wire [4-1:0] node10714;
	wire [4-1:0] node10715;
	wire [4-1:0] node10716;
	wire [4-1:0] node10720;
	wire [4-1:0] node10722;
	wire [4-1:0] node10725;
	wire [4-1:0] node10726;
	wire [4-1:0] node10727;
	wire [4-1:0] node10730;
	wire [4-1:0] node10733;
	wire [4-1:0] node10734;
	wire [4-1:0] node10736;
	wire [4-1:0] node10739;
	wire [4-1:0] node10740;
	wire [4-1:0] node10743;
	wire [4-1:0] node10746;
	wire [4-1:0] node10747;
	wire [4-1:0] node10748;
	wire [4-1:0] node10750;
	wire [4-1:0] node10753;
	wire [4-1:0] node10754;
	wire [4-1:0] node10755;
	wire [4-1:0] node10758;
	wire [4-1:0] node10761;
	wire [4-1:0] node10763;
	wire [4-1:0] node10766;
	wire [4-1:0] node10767;
	wire [4-1:0] node10768;
	wire [4-1:0] node10771;
	wire [4-1:0] node10772;
	wire [4-1:0] node10776;
	wire [4-1:0] node10777;
	wire [4-1:0] node10779;
	wire [4-1:0] node10780;
	wire [4-1:0] node10783;
	wire [4-1:0] node10786;
	wire [4-1:0] node10789;
	wire [4-1:0] node10790;
	wire [4-1:0] node10791;
	wire [4-1:0] node10792;
	wire [4-1:0] node10793;
	wire [4-1:0] node10794;
	wire [4-1:0] node10797;
	wire [4-1:0] node10800;
	wire [4-1:0] node10801;
	wire [4-1:0] node10802;
	wire [4-1:0] node10806;
	wire [4-1:0] node10807;
	wire [4-1:0] node10810;
	wire [4-1:0] node10813;
	wire [4-1:0] node10814;
	wire [4-1:0] node10815;
	wire [4-1:0] node10816;
	wire [4-1:0] node10819;
	wire [4-1:0] node10822;
	wire [4-1:0] node10823;
	wire [4-1:0] node10826;
	wire [4-1:0] node10829;
	wire [4-1:0] node10830;
	wire [4-1:0] node10833;
	wire [4-1:0] node10836;
	wire [4-1:0] node10837;
	wire [4-1:0] node10838;
	wire [4-1:0] node10840;
	wire [4-1:0] node10843;
	wire [4-1:0] node10844;
	wire [4-1:0] node10848;
	wire [4-1:0] node10849;
	wire [4-1:0] node10850;
	wire [4-1:0] node10851;
	wire [4-1:0] node10854;
	wire [4-1:0] node10855;
	wire [4-1:0] node10859;
	wire [4-1:0] node10860;
	wire [4-1:0] node10864;
	wire [4-1:0] node10865;
	wire [4-1:0] node10867;
	wire [4-1:0] node10870;
	wire [4-1:0] node10873;
	wire [4-1:0] node10874;
	wire [4-1:0] node10875;
	wire [4-1:0] node10876;
	wire [4-1:0] node10877;
	wire [4-1:0] node10880;
	wire [4-1:0] node10884;
	wire [4-1:0] node10885;
	wire [4-1:0] node10886;
	wire [4-1:0] node10887;
	wire [4-1:0] node10888;
	wire [4-1:0] node10891;
	wire [4-1:0] node10894;
	wire [4-1:0] node10895;
	wire [4-1:0] node10898;
	wire [4-1:0] node10901;
	wire [4-1:0] node10902;
	wire [4-1:0] node10906;
	wire [4-1:0] node10908;
	wire [4-1:0] node10911;
	wire [4-1:0] node10912;
	wire [4-1:0] node10913;
	wire [4-1:0] node10916;
	wire [4-1:0] node10917;
	wire [4-1:0] node10921;
	wire [4-1:0] node10923;
	wire [4-1:0] node10926;
	wire [4-1:0] node10927;
	wire [4-1:0] node10928;
	wire [4-1:0] node10929;
	wire [4-1:0] node10930;
	wire [4-1:0] node10931;
	wire [4-1:0] node10932;
	wire [4-1:0] node10933;
	wire [4-1:0] node10934;
	wire [4-1:0] node10937;
	wire [4-1:0] node10938;
	wire [4-1:0] node10942;
	wire [4-1:0] node10943;
	wire [4-1:0] node10946;
	wire [4-1:0] node10949;
	wire [4-1:0] node10950;
	wire [4-1:0] node10951;
	wire [4-1:0] node10952;
	wire [4-1:0] node10955;
	wire [4-1:0] node10958;
	wire [4-1:0] node10959;
	wire [4-1:0] node10963;
	wire [4-1:0] node10964;
	wire [4-1:0] node10967;
	wire [4-1:0] node10970;
	wire [4-1:0] node10971;
	wire [4-1:0] node10972;
	wire [4-1:0] node10973;
	wire [4-1:0] node10976;
	wire [4-1:0] node10979;
	wire [4-1:0] node10980;
	wire [4-1:0] node10982;
	wire [4-1:0] node10985;
	wire [4-1:0] node10988;
	wire [4-1:0] node10989;
	wire [4-1:0] node10990;
	wire [4-1:0] node10993;
	wire [4-1:0] node10996;
	wire [4-1:0] node10997;
	wire [4-1:0] node11000;
	wire [4-1:0] node11002;
	wire [4-1:0] node11005;
	wire [4-1:0] node11006;
	wire [4-1:0] node11007;
	wire [4-1:0] node11009;
	wire [4-1:0] node11012;
	wire [4-1:0] node11013;
	wire [4-1:0] node11014;
	wire [4-1:0] node11018;
	wire [4-1:0] node11019;
	wire [4-1:0] node11023;
	wire [4-1:0] node11024;
	wire [4-1:0] node11025;
	wire [4-1:0] node11026;
	wire [4-1:0] node11030;
	wire [4-1:0] node11031;
	wire [4-1:0] node11032;
	wire [4-1:0] node11036;
	wire [4-1:0] node11037;
	wire [4-1:0] node11041;
	wire [4-1:0] node11042;
	wire [4-1:0] node11043;
	wire [4-1:0] node11047;
	wire [4-1:0] node11048;
	wire [4-1:0] node11051;
	wire [4-1:0] node11054;
	wire [4-1:0] node11055;
	wire [4-1:0] node11056;
	wire [4-1:0] node11057;
	wire [4-1:0] node11058;
	wire [4-1:0] node11060;
	wire [4-1:0] node11061;
	wire [4-1:0] node11065;
	wire [4-1:0] node11066;
	wire [4-1:0] node11069;
	wire [4-1:0] node11072;
	wire [4-1:0] node11073;
	wire [4-1:0] node11075;
	wire [4-1:0] node11076;
	wire [4-1:0] node11079;
	wire [4-1:0] node11082;
	wire [4-1:0] node11083;
	wire [4-1:0] node11084;
	wire [4-1:0] node11089;
	wire [4-1:0] node11090;
	wire [4-1:0] node11091;
	wire [4-1:0] node11092;
	wire [4-1:0] node11096;
	wire [4-1:0] node11098;
	wire [4-1:0] node11100;
	wire [4-1:0] node11103;
	wire [4-1:0] node11104;
	wire [4-1:0] node11106;
	wire [4-1:0] node11107;
	wire [4-1:0] node11110;
	wire [4-1:0] node11113;
	wire [4-1:0] node11114;
	wire [4-1:0] node11115;
	wire [4-1:0] node11119;
	wire [4-1:0] node11121;
	wire [4-1:0] node11124;
	wire [4-1:0] node11125;
	wire [4-1:0] node11126;
	wire [4-1:0] node11127;
	wire [4-1:0] node11128;
	wire [4-1:0] node11130;
	wire [4-1:0] node11133;
	wire [4-1:0] node11136;
	wire [4-1:0] node11137;
	wire [4-1:0] node11140;
	wire [4-1:0] node11143;
	wire [4-1:0] node11144;
	wire [4-1:0] node11145;
	wire [4-1:0] node11149;
	wire [4-1:0] node11150;
	wire [4-1:0] node11152;
	wire [4-1:0] node11156;
	wire [4-1:0] node11157;
	wire [4-1:0] node11158;
	wire [4-1:0] node11160;
	wire [4-1:0] node11161;
	wire [4-1:0] node11165;
	wire [4-1:0] node11166;
	wire [4-1:0] node11168;
	wire [4-1:0] node11172;
	wire [4-1:0] node11173;
	wire [4-1:0] node11174;
	wire [4-1:0] node11177;
	wire [4-1:0] node11178;
	wire [4-1:0] node11181;
	wire [4-1:0] node11184;
	wire [4-1:0] node11185;
	wire [4-1:0] node11187;
	wire [4-1:0] node11190;
	wire [4-1:0] node11193;
	wire [4-1:0] node11194;
	wire [4-1:0] node11195;
	wire [4-1:0] node11196;
	wire [4-1:0] node11197;
	wire [4-1:0] node11199;
	wire [4-1:0] node11200;
	wire [4-1:0] node11204;
	wire [4-1:0] node11205;
	wire [4-1:0] node11209;
	wire [4-1:0] node11210;
	wire [4-1:0] node11211;
	wire [4-1:0] node11212;
	wire [4-1:0] node11215;
	wire [4-1:0] node11218;
	wire [4-1:0] node11219;
	wire [4-1:0] node11222;
	wire [4-1:0] node11225;
	wire [4-1:0] node11226;
	wire [4-1:0] node11228;
	wire [4-1:0] node11231;
	wire [4-1:0] node11234;
	wire [4-1:0] node11235;
	wire [4-1:0] node11236;
	wire [4-1:0] node11237;
	wire [4-1:0] node11240;
	wire [4-1:0] node11241;
	wire [4-1:0] node11245;
	wire [4-1:0] node11246;
	wire [4-1:0] node11248;
	wire [4-1:0] node11251;
	wire [4-1:0] node11252;
	wire [4-1:0] node11256;
	wire [4-1:0] node11257;
	wire [4-1:0] node11258;
	wire [4-1:0] node11260;
	wire [4-1:0] node11263;
	wire [4-1:0] node11265;
	wire [4-1:0] node11268;
	wire [4-1:0] node11269;
	wire [4-1:0] node11270;
	wire [4-1:0] node11273;
	wire [4-1:0] node11276;
	wire [4-1:0] node11277;
	wire [4-1:0] node11280;
	wire [4-1:0] node11283;
	wire [4-1:0] node11284;
	wire [4-1:0] node11285;
	wire [4-1:0] node11286;
	wire [4-1:0] node11287;
	wire [4-1:0] node11290;
	wire [4-1:0] node11293;
	wire [4-1:0] node11294;
	wire [4-1:0] node11295;
	wire [4-1:0] node11298;
	wire [4-1:0] node11302;
	wire [4-1:0] node11303;
	wire [4-1:0] node11305;
	wire [4-1:0] node11306;
	wire [4-1:0] node11310;
	wire [4-1:0] node11311;
	wire [4-1:0] node11313;
	wire [4-1:0] node11316;
	wire [4-1:0] node11317;
	wire [4-1:0] node11321;
	wire [4-1:0] node11322;
	wire [4-1:0] node11323;
	wire [4-1:0] node11324;
	wire [4-1:0] node11327;
	wire [4-1:0] node11330;
	wire [4-1:0] node11331;
	wire [4-1:0] node11332;
	wire [4-1:0] node11336;
	wire [4-1:0] node11337;
	wire [4-1:0] node11341;
	wire [4-1:0] node11342;
	wire [4-1:0] node11344;
	wire [4-1:0] node11348;
	wire [4-1:0] node11349;
	wire [4-1:0] node11350;
	wire [4-1:0] node11351;
	wire [4-1:0] node11352;
	wire [4-1:0] node11353;
	wire [4-1:0] node11354;
	wire [4-1:0] node11355;
	wire [4-1:0] node11359;
	wire [4-1:0] node11361;
	wire [4-1:0] node11364;
	wire [4-1:0] node11365;
	wire [4-1:0] node11366;
	wire [4-1:0] node11369;
	wire [4-1:0] node11371;
	wire [4-1:0] node11374;
	wire [4-1:0] node11375;
	wire [4-1:0] node11379;
	wire [4-1:0] node11380;
	wire [4-1:0] node11381;
	wire [4-1:0] node11383;
	wire [4-1:0] node11385;
	wire [4-1:0] node11388;
	wire [4-1:0] node11389;
	wire [4-1:0] node11392;
	wire [4-1:0] node11395;
	wire [4-1:0] node11396;
	wire [4-1:0] node11397;
	wire [4-1:0] node11399;
	wire [4-1:0] node11402;
	wire [4-1:0] node11403;
	wire [4-1:0] node11407;
	wire [4-1:0] node11408;
	wire [4-1:0] node11411;
	wire [4-1:0] node11414;
	wire [4-1:0] node11415;
	wire [4-1:0] node11416;
	wire [4-1:0] node11417;
	wire [4-1:0] node11418;
	wire [4-1:0] node11421;
	wire [4-1:0] node11425;
	wire [4-1:0] node11426;
	wire [4-1:0] node11427;
	wire [4-1:0] node11431;
	wire [4-1:0] node11433;
	wire [4-1:0] node11436;
	wire [4-1:0] node11437;
	wire [4-1:0] node11438;
	wire [4-1:0] node11439;
	wire [4-1:0] node11443;
	wire [4-1:0] node11444;
	wire [4-1:0] node11447;
	wire [4-1:0] node11450;
	wire [4-1:0] node11451;
	wire [4-1:0] node11453;
	wire [4-1:0] node11456;
	wire [4-1:0] node11458;
	wire [4-1:0] node11461;
	wire [4-1:0] node11462;
	wire [4-1:0] node11463;
	wire [4-1:0] node11464;
	wire [4-1:0] node11465;
	wire [4-1:0] node11466;
	wire [4-1:0] node11468;
	wire [4-1:0] node11471;
	wire [4-1:0] node11474;
	wire [4-1:0] node11476;
	wire [4-1:0] node11477;
	wire [4-1:0] node11481;
	wire [4-1:0] node11482;
	wire [4-1:0] node11483;
	wire [4-1:0] node11485;
	wire [4-1:0] node11488;
	wire [4-1:0] node11491;
	wire [4-1:0] node11492;
	wire [4-1:0] node11493;
	wire [4-1:0] node11498;
	wire [4-1:0] node11499;
	wire [4-1:0] node11501;
	wire [4-1:0] node11502;
	wire [4-1:0] node11503;
	wire [4-1:0] node11506;
	wire [4-1:0] node11509;
	wire [4-1:0] node11510;
	wire [4-1:0] node11513;
	wire [4-1:0] node11516;
	wire [4-1:0] node11517;
	wire [4-1:0] node11519;
	wire [4-1:0] node11520;
	wire [4-1:0] node11524;
	wire [4-1:0] node11525;
	wire [4-1:0] node11527;
	wire [4-1:0] node11530;
	wire [4-1:0] node11531;
	wire [4-1:0] node11535;
	wire [4-1:0] node11536;
	wire [4-1:0] node11537;
	wire [4-1:0] node11538;
	wire [4-1:0] node11539;
	wire [4-1:0] node11542;
	wire [4-1:0] node11545;
	wire [4-1:0] node11546;
	wire [4-1:0] node11550;
	wire [4-1:0] node11551;
	wire [4-1:0] node11552;
	wire [4-1:0] node11556;
	wire [4-1:0] node11557;
	wire [4-1:0] node11561;
	wire [4-1:0] node11563;
	wire [4-1:0] node11565;
	wire [4-1:0] node11568;
	wire [4-1:0] node11569;
	wire [4-1:0] node11570;
	wire [4-1:0] node11571;
	wire [4-1:0] node11572;
	wire [4-1:0] node11573;
	wire [4-1:0] node11574;
	wire [4-1:0] node11579;
	wire [4-1:0] node11580;
	wire [4-1:0] node11581;
	wire [4-1:0] node11582;
	wire [4-1:0] node11585;
	wire [4-1:0] node11588;
	wire [4-1:0] node11589;
	wire [4-1:0] node11592;
	wire [4-1:0] node11595;
	wire [4-1:0] node11596;
	wire [4-1:0] node11599;
	wire [4-1:0] node11600;
	wire [4-1:0] node11604;
	wire [4-1:0] node11605;
	wire [4-1:0] node11606;
	wire [4-1:0] node11607;
	wire [4-1:0] node11609;
	wire [4-1:0] node11612;
	wire [4-1:0] node11613;
	wire [4-1:0] node11617;
	wire [4-1:0] node11618;
	wire [4-1:0] node11621;
	wire [4-1:0] node11623;
	wire [4-1:0] node11626;
	wire [4-1:0] node11627;
	wire [4-1:0] node11628;
	wire [4-1:0] node11629;
	wire [4-1:0] node11632;
	wire [4-1:0] node11636;
	wire [4-1:0] node11639;
	wire [4-1:0] node11640;
	wire [4-1:0] node11641;
	wire [4-1:0] node11642;
	wire [4-1:0] node11643;
	wire [4-1:0] node11644;
	wire [4-1:0] node11647;
	wire [4-1:0] node11650;
	wire [4-1:0] node11652;
	wire [4-1:0] node11656;
	wire [4-1:0] node11657;
	wire [4-1:0] node11658;
	wire [4-1:0] node11661;
	wire [4-1:0] node11662;
	wire [4-1:0] node11666;
	wire [4-1:0] node11667;
	wire [4-1:0] node11669;
	wire [4-1:0] node11673;
	wire [4-1:0] node11674;
	wire [4-1:0] node11675;
	wire [4-1:0] node11676;
	wire [4-1:0] node11680;
	wire [4-1:0] node11682;
	wire [4-1:0] node11686;
	wire [4-1:0] node11687;
	wire [4-1:0] node11688;
	wire [4-1:0] node11689;
	wire [4-1:0] node11690;
	wire [4-1:0] node11691;
	wire [4-1:0] node11693;
	wire [4-1:0] node11697;
	wire [4-1:0] node11699;
	wire [4-1:0] node11700;
	wire [4-1:0] node11705;
	wire [4-1:0] node11706;
	wire [4-1:0] node11708;
	wire [4-1:0] node11709;
	wire [4-1:0] node11711;
	wire [4-1:0] node11714;
	wire [4-1:0] node11716;
	wire [4-1:0] node11720;
	wire [4-1:0] node11721;
	wire [4-1:0] node11722;
	wire [4-1:0] node11723;
	wire [4-1:0] node11724;
	wire [4-1:0] node11725;
	wire [4-1:0] node11729;
	wire [4-1:0] node11731;
	wire [4-1:0] node11734;
	wire [4-1:0] node11735;
	wire [4-1:0] node11738;
	wire [4-1:0] node11740;
	wire [4-1:0] node11745;
	wire [4-1:0] node11747;
	wire [4-1:0] node11748;
	wire [4-1:0] node11749;
	wire [4-1:0] node11751;
	wire [4-1:0] node11752;
	wire [4-1:0] node11753;
	wire [4-1:0] node11755;
	wire [4-1:0] node11756;
	wire [4-1:0] node11759;
	wire [4-1:0] node11761;
	wire [4-1:0] node11762;
	wire [4-1:0] node11766;
	wire [4-1:0] node11767;
	wire [4-1:0] node11768;
	wire [4-1:0] node11769;
	wire [4-1:0] node11770;
	wire [4-1:0] node11773;
	wire [4-1:0] node11776;
	wire [4-1:0] node11777;
	wire [4-1:0] node11779;
	wire [4-1:0] node11782;
	wire [4-1:0] node11784;
	wire [4-1:0] node11787;
	wire [4-1:0] node11788;
	wire [4-1:0] node11790;
	wire [4-1:0] node11793;
	wire [4-1:0] node11796;
	wire [4-1:0] node11797;
	wire [4-1:0] node11798;
	wire [4-1:0] node11800;
	wire [4-1:0] node11801;
	wire [4-1:0] node11804;
	wire [4-1:0] node11807;
	wire [4-1:0] node11809;
	wire [4-1:0] node11811;
	wire [4-1:0] node11814;
	wire [4-1:0] node11815;
	wire [4-1:0] node11817;
	wire [4-1:0] node11820;
	wire [4-1:0] node11822;
	wire [4-1:0] node11825;
	wire [4-1:0] node11827;
	wire [4-1:0] node11829;
	wire [4-1:0] node11830;
	wire [4-1:0] node11831;
	wire [4-1:0] node11833;
	wire [4-1:0] node11836;
	wire [4-1:0] node11838;
	wire [4-1:0] node11841;
	wire [4-1:0] node11843;
	wire [4-1:0] node11844;
	wire [4-1:0] node11845;
	wire [4-1:0] node11850;
	wire [4-1:0] node11851;
	wire [4-1:0] node11852;
	wire [4-1:0] node11853;
	wire [4-1:0] node11854;
	wire [4-1:0] node11855;
	wire [4-1:0] node11856;
	wire [4-1:0] node11857;
	wire [4-1:0] node11860;
	wire [4-1:0] node11863;
	wire [4-1:0] node11864;
	wire [4-1:0] node11868;
	wire [4-1:0] node11869;
	wire [4-1:0] node11872;
	wire [4-1:0] node11873;
	wire [4-1:0] node11877;
	wire [4-1:0] node11878;
	wire [4-1:0] node11879;
	wire [4-1:0] node11880;
	wire [4-1:0] node11884;
	wire [4-1:0] node11885;
	wire [4-1:0] node11889;
	wire [4-1:0] node11890;
	wire [4-1:0] node11891;
	wire [4-1:0] node11894;
	wire [4-1:0] node11895;
	wire [4-1:0] node11898;
	wire [4-1:0] node11901;
	wire [4-1:0] node11902;
	wire [4-1:0] node11903;
	wire [4-1:0] node11908;
	wire [4-1:0] node11909;
	wire [4-1:0] node11910;
	wire [4-1:0] node11911;
	wire [4-1:0] node11912;
	wire [4-1:0] node11915;
	wire [4-1:0] node11918;
	wire [4-1:0] node11919;
	wire [4-1:0] node11922;
	wire [4-1:0] node11925;
	wire [4-1:0] node11926;
	wire [4-1:0] node11928;
	wire [4-1:0] node11931;
	wire [4-1:0] node11933;
	wire [4-1:0] node11934;
	wire [4-1:0] node11937;
	wire [4-1:0] node11940;
	wire [4-1:0] node11941;
	wire [4-1:0] node11942;
	wire [4-1:0] node11944;
	wire [4-1:0] node11945;
	wire [4-1:0] node11949;
	wire [4-1:0] node11950;
	wire [4-1:0] node11954;
	wire [4-1:0] node11955;
	wire [4-1:0] node11956;
	wire [4-1:0] node11959;
	wire [4-1:0] node11960;
	wire [4-1:0] node11963;
	wire [4-1:0] node11966;
	wire [4-1:0] node11967;
	wire [4-1:0] node11969;
	wire [4-1:0] node11972;
	wire [4-1:0] node11975;
	wire [4-1:0] node11976;
	wire [4-1:0] node11977;
	wire [4-1:0] node11978;
	wire [4-1:0] node11980;
	wire [4-1:0] node11982;
	wire [4-1:0] node11985;
	wire [4-1:0] node11986;
	wire [4-1:0] node11988;
	wire [4-1:0] node11991;
	wire [4-1:0] node11993;
	wire [4-1:0] node11996;
	wire [4-1:0] node11997;
	wire [4-1:0] node11998;
	wire [4-1:0] node12001;
	wire [4-1:0] node12002;
	wire [4-1:0] node12005;
	wire [4-1:0] node12008;
	wire [4-1:0] node12009;
	wire [4-1:0] node12011;
	wire [4-1:0] node12014;
	wire [4-1:0] node12016;
	wire [4-1:0] node12019;
	wire [4-1:0] node12020;
	wire [4-1:0] node12021;
	wire [4-1:0] node12022;
	wire [4-1:0] node12024;
	wire [4-1:0] node12027;
	wire [4-1:0] node12028;
	wire [4-1:0] node12032;
	wire [4-1:0] node12033;
	wire [4-1:0] node12035;
	wire [4-1:0] node12039;
	wire [4-1:0] node12040;
	wire [4-1:0] node12041;
	wire [4-1:0] node12042;
	wire [4-1:0] node12045;
	wire [4-1:0] node12048;
	wire [4-1:0] node12049;
	wire [4-1:0] node12051;
	wire [4-1:0] node12055;
	wire [4-1:0] node12056;
	wire [4-1:0] node12057;
	wire [4-1:0] node12060;
	wire [4-1:0] node12061;
	wire [4-1:0] node12066;
	wire [4-1:0] node12067;
	wire [4-1:0] node12068;
	wire [4-1:0] node12069;
	wire [4-1:0] node12070;
	wire [4-1:0] node12071;
	wire [4-1:0] node12073;
	wire [4-1:0] node12076;
	wire [4-1:0] node12077;
	wire [4-1:0] node12078;
	wire [4-1:0] node12082;
	wire [4-1:0] node12084;
	wire [4-1:0] node12087;
	wire [4-1:0] node12088;
	wire [4-1:0] node12089;
	wire [4-1:0] node12090;
	wire [4-1:0] node12093;
	wire [4-1:0] node12096;
	wire [4-1:0] node12098;
	wire [4-1:0] node12101;
	wire [4-1:0] node12102;
	wire [4-1:0] node12105;
	wire [4-1:0] node12108;
	wire [4-1:0] node12109;
	wire [4-1:0] node12110;
	wire [4-1:0] node12112;
	wire [4-1:0] node12115;
	wire [4-1:0] node12116;
	wire [4-1:0] node12120;
	wire [4-1:0] node12121;
	wire [4-1:0] node12122;
	wire [4-1:0] node12127;
	wire [4-1:0] node12128;
	wire [4-1:0] node12129;
	wire [4-1:0] node12130;
	wire [4-1:0] node12132;
	wire [4-1:0] node12135;
	wire [4-1:0] node12137;
	wire [4-1:0] node12140;
	wire [4-1:0] node12141;
	wire [4-1:0] node12142;
	wire [4-1:0] node12146;
	wire [4-1:0] node12148;
	wire [4-1:0] node12151;
	wire [4-1:0] node12152;
	wire [4-1:0] node12153;
	wire [4-1:0] node12155;
	wire [4-1:0] node12156;
	wire [4-1:0] node12160;
	wire [4-1:0] node12161;
	wire [4-1:0] node12162;
	wire [4-1:0] node12165;
	wire [4-1:0] node12168;
	wire [4-1:0] node12171;
	wire [4-1:0] node12172;
	wire [4-1:0] node12173;
	wire [4-1:0] node12178;
	wire [4-1:0] node12179;
	wire [4-1:0] node12180;
	wire [4-1:0] node12181;
	wire [4-1:0] node12182;
	wire [4-1:0] node12183;
	wire [4-1:0] node12188;
	wire [4-1:0] node12189;
	wire [4-1:0] node12190;
	wire [4-1:0] node12191;
	wire [4-1:0] node12196;
	wire [4-1:0] node12198;
	wire [4-1:0] node12201;
	wire [4-1:0] node12202;
	wire [4-1:0] node12203;
	wire [4-1:0] node12204;
	wire [4-1:0] node12208;
	wire [4-1:0] node12209;
	wire [4-1:0] node12213;
	wire [4-1:0] node12214;
	wire [4-1:0] node12215;
	wire [4-1:0] node12216;
	wire [4-1:0] node12220;
	wire [4-1:0] node12221;
	wire [4-1:0] node12226;
	wire [4-1:0] node12227;
	wire [4-1:0] node12228;
	wire [4-1:0] node12229;
	wire [4-1:0] node12233;
	wire [4-1:0] node12235;
	wire [4-1:0] node12236;
	wire [4-1:0] node12237;
	wire [4-1:0] node12241;
	wire [4-1:0] node12242;
	wire [4-1:0] node12246;
	wire [4-1:0] node12247;
	wire [4-1:0] node12248;
	wire [4-1:0] node12249;
	wire [4-1:0] node12250;
	wire [4-1:0] node12253;
	wire [4-1:0] node12259;
	wire [4-1:0] node12261;
	wire [4-1:0] node12263;
	wire [4-1:0] node12264;
	wire [4-1:0] node12266;
	wire [4-1:0] node12267;
	wire [4-1:0] node12268;
	wire [4-1:0] node12269;
	wire [4-1:0] node12270;
	wire [4-1:0] node12274;
	wire [4-1:0] node12276;
	wire [4-1:0] node12279;
	wire [4-1:0] node12280;
	wire [4-1:0] node12282;
	wire [4-1:0] node12287;
	wire [4-1:0] node12288;
	wire [4-1:0] node12289;
	wire [4-1:0] node12290;
	wire [4-1:0] node12291;
	wire [4-1:0] node12292;
	wire [4-1:0] node12293;
	wire [4-1:0] node12297;
	wire [4-1:0] node12300;
	wire [4-1:0] node12301;
	wire [4-1:0] node12304;
	wire [4-1:0] node12307;
	wire [4-1:0] node12308;
	wire [4-1:0] node12309;
	wire [4-1:0] node12314;
	wire [4-1:0] node12315;
	wire [4-1:0] node12316;
	wire [4-1:0] node12317;
	wire [4-1:0] node12320;
	wire [4-1:0] node12324;
	wire [4-1:0] node12325;
	wire [4-1:0] node12326;
	wire [4-1:0] node12330;
	wire [4-1:0] node12331;
	wire [4-1:0] node12333;
	wire [4-1:0] node12337;
	wire [4-1:0] node12339;
	wire [4-1:0] node12340;
	wire [4-1:0] node12341;
	wire [4-1:0] node12343;
	wire [4-1:0] node12347;
	wire [4-1:0] node12349;
	wire [4-1:0] node12351;
	wire [4-1:0] node12354;
	wire [4-1:0] node12355;
	wire [4-1:0] node12356;
	wire [4-1:0] node12357;
	wire [4-1:0] node12358;
	wire [4-1:0] node12359;
	wire [4-1:0] node12360;
	wire [4-1:0] node12361;
	wire [4-1:0] node12362;
	wire [4-1:0] node12363;
	wire [4-1:0] node12364;
	wire [4-1:0] node12365;
	wire [4-1:0] node12367;
	wire [4-1:0] node12369;
	wire [4-1:0] node12373;
	wire [4-1:0] node12374;
	wire [4-1:0] node12375;
	wire [4-1:0] node12379;
	wire [4-1:0] node12380;
	wire [4-1:0] node12381;
	wire [4-1:0] node12385;
	wire [4-1:0] node12387;
	wire [4-1:0] node12390;
	wire [4-1:0] node12391;
	wire [4-1:0] node12393;
	wire [4-1:0] node12396;
	wire [4-1:0] node12397;
	wire [4-1:0] node12398;
	wire [4-1:0] node12402;
	wire [4-1:0] node12403;
	wire [4-1:0] node12407;
	wire [4-1:0] node12408;
	wire [4-1:0] node12409;
	wire [4-1:0] node12410;
	wire [4-1:0] node12412;
	wire [4-1:0] node12415;
	wire [4-1:0] node12416;
	wire [4-1:0] node12420;
	wire [4-1:0] node12421;
	wire [4-1:0] node12423;
	wire [4-1:0] node12425;
	wire [4-1:0] node12428;
	wire [4-1:0] node12429;
	wire [4-1:0] node12432;
	wire [4-1:0] node12433;
	wire [4-1:0] node12437;
	wire [4-1:0] node12438;
	wire [4-1:0] node12439;
	wire [4-1:0] node12441;
	wire [4-1:0] node12442;
	wire [4-1:0] node12446;
	wire [4-1:0] node12448;
	wire [4-1:0] node12449;
	wire [4-1:0] node12451;
	wire [4-1:0] node12454;
	wire [4-1:0] node12457;
	wire [4-1:0] node12458;
	wire [4-1:0] node12461;
	wire [4-1:0] node12463;
	wire [4-1:0] node12466;
	wire [4-1:0] node12467;
	wire [4-1:0] node12468;
	wire [4-1:0] node12469;
	wire [4-1:0] node12470;
	wire [4-1:0] node12471;
	wire [4-1:0] node12475;
	wire [4-1:0] node12476;
	wire [4-1:0] node12478;
	wire [4-1:0] node12481;
	wire [4-1:0] node12482;
	wire [4-1:0] node12486;
	wire [4-1:0] node12488;
	wire [4-1:0] node12489;
	wire [4-1:0] node12491;
	wire [4-1:0] node12493;
	wire [4-1:0] node12496;
	wire [4-1:0] node12497;
	wire [4-1:0] node12501;
	wire [4-1:0] node12502;
	wire [4-1:0] node12503;
	wire [4-1:0] node12507;
	wire [4-1:0] node12508;
	wire [4-1:0] node12510;
	wire [4-1:0] node12513;
	wire [4-1:0] node12515;
	wire [4-1:0] node12518;
	wire [4-1:0] node12519;
	wire [4-1:0] node12520;
	wire [4-1:0] node12521;
	wire [4-1:0] node12522;
	wire [4-1:0] node12526;
	wire [4-1:0] node12527;
	wire [4-1:0] node12529;
	wire [4-1:0] node12532;
	wire [4-1:0] node12533;
	wire [4-1:0] node12537;
	wire [4-1:0] node12538;
	wire [4-1:0] node12539;
	wire [4-1:0] node12543;
	wire [4-1:0] node12544;
	wire [4-1:0] node12545;
	wire [4-1:0] node12549;
	wire [4-1:0] node12550;
	wire [4-1:0] node12554;
	wire [4-1:0] node12555;
	wire [4-1:0] node12556;
	wire [4-1:0] node12558;
	wire [4-1:0] node12561;
	wire [4-1:0] node12562;
	wire [4-1:0] node12566;
	wire [4-1:0] node12568;
	wire [4-1:0] node12571;
	wire [4-1:0] node12572;
	wire [4-1:0] node12573;
	wire [4-1:0] node12574;
	wire [4-1:0] node12575;
	wire [4-1:0] node12577;
	wire [4-1:0] node12578;
	wire [4-1:0] node12582;
	wire [4-1:0] node12584;
	wire [4-1:0] node12587;
	wire [4-1:0] node12588;
	wire [4-1:0] node12589;
	wire [4-1:0] node12590;
	wire [4-1:0] node12591;
	wire [4-1:0] node12595;
	wire [4-1:0] node12598;
	wire [4-1:0] node12599;
	wire [4-1:0] node12603;
	wire [4-1:0] node12604;
	wire [4-1:0] node12606;
	wire [4-1:0] node12607;
	wire [4-1:0] node12611;
	wire [4-1:0] node12613;
	wire [4-1:0] node12616;
	wire [4-1:0] node12617;
	wire [4-1:0] node12618;
	wire [4-1:0] node12619;
	wire [4-1:0] node12621;
	wire [4-1:0] node12624;
	wire [4-1:0] node12626;
	wire [4-1:0] node12629;
	wire [4-1:0] node12630;
	wire [4-1:0] node12632;
	wire [4-1:0] node12633;
	wire [4-1:0] node12637;
	wire [4-1:0] node12638;
	wire [4-1:0] node12642;
	wire [4-1:0] node12643;
	wire [4-1:0] node12645;
	wire [4-1:0] node12646;
	wire [4-1:0] node12650;
	wire [4-1:0] node12652;
	wire [4-1:0] node12655;
	wire [4-1:0] node12656;
	wire [4-1:0] node12657;
	wire [4-1:0] node12658;
	wire [4-1:0] node12659;
	wire [4-1:0] node12661;
	wire [4-1:0] node12664;
	wire [4-1:0] node12665;
	wire [4-1:0] node12668;
	wire [4-1:0] node12670;
	wire [4-1:0] node12673;
	wire [4-1:0] node12674;
	wire [4-1:0] node12675;
	wire [4-1:0] node12676;
	wire [4-1:0] node12680;
	wire [4-1:0] node12682;
	wire [4-1:0] node12685;
	wire [4-1:0] node12686;
	wire [4-1:0] node12690;
	wire [4-1:0] node12691;
	wire [4-1:0] node12692;
	wire [4-1:0] node12693;
	wire [4-1:0] node12695;
	wire [4-1:0] node12698;
	wire [4-1:0] node12701;
	wire [4-1:0] node12702;
	wire [4-1:0] node12704;
	wire [4-1:0] node12707;
	wire [4-1:0] node12709;
	wire [4-1:0] node12712;
	wire [4-1:0] node12713;
	wire [4-1:0] node12715;
	wire [4-1:0] node12717;
	wire [4-1:0] node12720;
	wire [4-1:0] node12722;
	wire [4-1:0] node12725;
	wire [4-1:0] node12726;
	wire [4-1:0] node12727;
	wire [4-1:0] node12728;
	wire [4-1:0] node12730;
	wire [4-1:0] node12731;
	wire [4-1:0] node12732;
	wire [4-1:0] node12737;
	wire [4-1:0] node12739;
	wire [4-1:0] node12742;
	wire [4-1:0] node12743;
	wire [4-1:0] node12745;
	wire [4-1:0] node12747;
	wire [4-1:0] node12748;
	wire [4-1:0] node12751;
	wire [4-1:0] node12754;
	wire [4-1:0] node12755;
	wire [4-1:0] node12757;
	wire [4-1:0] node12758;
	wire [4-1:0] node12762;
	wire [4-1:0] node12765;
	wire [4-1:0] node12766;
	wire [4-1:0] node12767;
	wire [4-1:0] node12768;
	wire [4-1:0] node12770;
	wire [4-1:0] node12773;
	wire [4-1:0] node12776;
	wire [4-1:0] node12777;
	wire [4-1:0] node12778;
	wire [4-1:0] node12782;
	wire [4-1:0] node12783;
	wire [4-1:0] node12787;
	wire [4-1:0] node12788;
	wire [4-1:0] node12789;
	wire [4-1:0] node12791;
	wire [4-1:0] node12792;
	wire [4-1:0] node12797;
	wire [4-1:0] node12798;
	wire [4-1:0] node12802;
	wire [4-1:0] node12804;
	wire [4-1:0] node12805;
	wire [4-1:0] node12806;
	wire [4-1:0] node12807;
	wire [4-1:0] node12808;
	wire [4-1:0] node12809;
	wire [4-1:0] node12810;
	wire [4-1:0] node12812;
	wire [4-1:0] node12813;
	wire [4-1:0] node12817;
	wire [4-1:0] node12820;
	wire [4-1:0] node12822;
	wire [4-1:0] node12825;
	wire [4-1:0] node12826;
	wire [4-1:0] node12827;
	wire [4-1:0] node12828;
	wire [4-1:0] node12830;
	wire [4-1:0] node12834;
	wire [4-1:0] node12835;
	wire [4-1:0] node12837;
	wire [4-1:0] node12841;
	wire [4-1:0] node12842;
	wire [4-1:0] node12845;
	wire [4-1:0] node12846;
	wire [4-1:0] node12849;
	wire [4-1:0] node12853;
	wire [4-1:0] node12854;
	wire [4-1:0] node12855;
	wire [4-1:0] node12856;
	wire [4-1:0] node12857;
	wire [4-1:0] node12858;
	wire [4-1:0] node12862;
	wire [4-1:0] node12863;
	wire [4-1:0] node12865;
	wire [4-1:0] node12869;
	wire [4-1:0] node12870;
	wire [4-1:0] node12871;
	wire [4-1:0] node12874;
	wire [4-1:0] node12875;
	wire [4-1:0] node12879;
	wire [4-1:0] node12881;
	wire [4-1:0] node12884;
	wire [4-1:0] node12885;
	wire [4-1:0] node12886;
	wire [4-1:0] node12889;
	wire [4-1:0] node12890;
	wire [4-1:0] node12891;
	wire [4-1:0] node12895;
	wire [4-1:0] node12896;
	wire [4-1:0] node12900;
	wire [4-1:0] node12902;
	wire [4-1:0] node12904;
	wire [4-1:0] node12906;
	wire [4-1:0] node12909;
	wire [4-1:0] node12910;
	wire [4-1:0] node12911;
	wire [4-1:0] node12913;
	wire [4-1:0] node12916;
	wire [4-1:0] node12917;
	wire [4-1:0] node12919;
	wire [4-1:0] node12922;
	wire [4-1:0] node12924;
	wire [4-1:0] node12927;
	wire [4-1:0] node12928;
	wire [4-1:0] node12929;
	wire [4-1:0] node12931;
	wire [4-1:0] node12934;
	wire [4-1:0] node12936;
	wire [4-1:0] node12939;
	wire [4-1:0] node12941;
	wire [4-1:0] node12944;
	wire [4-1:0] node12945;
	wire [4-1:0] node12946;
	wire [4-1:0] node12947;
	wire [4-1:0] node12948;
	wire [4-1:0] node12949;
	wire [4-1:0] node12950;
	wire [4-1:0] node12954;
	wire [4-1:0] node12957;
	wire [4-1:0] node12958;
	wire [4-1:0] node12959;
	wire [4-1:0] node12963;
	wire [4-1:0] node12964;
	wire [4-1:0] node12965;
	wire [4-1:0] node12969;
	wire [4-1:0] node12971;
	wire [4-1:0] node12974;
	wire [4-1:0] node12975;
	wire [4-1:0] node12977;
	wire [4-1:0] node12979;
	wire [4-1:0] node12982;
	wire [4-1:0] node12983;
	wire [4-1:0] node12987;
	wire [4-1:0] node12988;
	wire [4-1:0] node12989;
	wire [4-1:0] node12990;
	wire [4-1:0] node12992;
	wire [4-1:0] node12995;
	wire [4-1:0] node12997;
	wire [4-1:0] node13000;
	wire [4-1:0] node13001;
	wire [4-1:0] node13005;
	wire [4-1:0] node13006;
	wire [4-1:0] node13007;
	wire [4-1:0] node13009;
	wire [4-1:0] node13012;
	wire [4-1:0] node13015;
	wire [4-1:0] node13016;
	wire [4-1:0] node13017;
	wire [4-1:0] node13021;
	wire [4-1:0] node13023;
	wire [4-1:0] node13026;
	wire [4-1:0] node13027;
	wire [4-1:0] node13028;
	wire [4-1:0] node13029;
	wire [4-1:0] node13030;
	wire [4-1:0] node13033;
	wire [4-1:0] node13035;
	wire [4-1:0] node13038;
	wire [4-1:0] node13039;
	wire [4-1:0] node13040;
	wire [4-1:0] node13044;
	wire [4-1:0] node13046;
	wire [4-1:0] node13049;
	wire [4-1:0] node13050;
	wire [4-1:0] node13051;
	wire [4-1:0] node13052;
	wire [4-1:0] node13056;
	wire [4-1:0] node13057;
	wire [4-1:0] node13061;
	wire [4-1:0] node13062;
	wire [4-1:0] node13066;
	wire [4-1:0] node13067;
	wire [4-1:0] node13068;
	wire [4-1:0] node13070;
	wire [4-1:0] node13071;
	wire [4-1:0] node13075;
	wire [4-1:0] node13076;
	wire [4-1:0] node13080;
	wire [4-1:0] node13081;
	wire [4-1:0] node13082;
	wire [4-1:0] node13083;
	wire [4-1:0] node13084;
	wire [4-1:0] node13090;
	wire [4-1:0] node13091;
	wire [4-1:0] node13093;
	wire [4-1:0] node13094;
	wire [4-1:0] node13098;
	wire [4-1:0] node13100;
	wire [4-1:0] node13104;
	wire [4-1:0] node13105;
	wire [4-1:0] node13106;
	wire [4-1:0] node13107;
	wire [4-1:0] node13108;
	wire [4-1:0] node13109;
	wire [4-1:0] node13110;
	wire [4-1:0] node13111;
	wire [4-1:0] node13112;
	wire [4-1:0] node13113;
	wire [4-1:0] node13116;
	wire [4-1:0] node13117;
	wire [4-1:0] node13118;
	wire [4-1:0] node13122;
	wire [4-1:0] node13123;
	wire [4-1:0] node13127;
	wire [4-1:0] node13128;
	wire [4-1:0] node13130;
	wire [4-1:0] node13133;
	wire [4-1:0] node13134;
	wire [4-1:0] node13137;
	wire [4-1:0] node13140;
	wire [4-1:0] node13141;
	wire [4-1:0] node13143;
	wire [4-1:0] node13145;
	wire [4-1:0] node13148;
	wire [4-1:0] node13149;
	wire [4-1:0] node13150;
	wire [4-1:0] node13153;
	wire [4-1:0] node13154;
	wire [4-1:0] node13158;
	wire [4-1:0] node13159;
	wire [4-1:0] node13162;
	wire [4-1:0] node13165;
	wire [4-1:0] node13166;
	wire [4-1:0] node13167;
	wire [4-1:0] node13168;
	wire [4-1:0] node13170;
	wire [4-1:0] node13173;
	wire [4-1:0] node13174;
	wire [4-1:0] node13178;
	wire [4-1:0] node13179;
	wire [4-1:0] node13182;
	wire [4-1:0] node13185;
	wire [4-1:0] node13186;
	wire [4-1:0] node13187;
	wire [4-1:0] node13188;
	wire [4-1:0] node13190;
	wire [4-1:0] node13193;
	wire [4-1:0] node13194;
	wire [4-1:0] node13199;
	wire [4-1:0] node13200;
	wire [4-1:0] node13202;
	wire [4-1:0] node13203;
	wire [4-1:0] node13207;
	wire [4-1:0] node13208;
	wire [4-1:0] node13212;
	wire [4-1:0] node13213;
	wire [4-1:0] node13214;
	wire [4-1:0] node13215;
	wire [4-1:0] node13216;
	wire [4-1:0] node13217;
	wire [4-1:0] node13221;
	wire [4-1:0] node13222;
	wire [4-1:0] node13225;
	wire [4-1:0] node13226;
	wire [4-1:0] node13229;
	wire [4-1:0] node13232;
	wire [4-1:0] node13233;
	wire [4-1:0] node13234;
	wire [4-1:0] node13238;
	wire [4-1:0] node13239;
	wire [4-1:0] node13243;
	wire [4-1:0] node13244;
	wire [4-1:0] node13245;
	wire [4-1:0] node13248;
	wire [4-1:0] node13249;
	wire [4-1:0] node13253;
	wire [4-1:0] node13254;
	wire [4-1:0] node13255;
	wire [4-1:0] node13258;
	wire [4-1:0] node13261;
	wire [4-1:0] node13262;
	wire [4-1:0] node13265;
	wire [4-1:0] node13266;
	wire [4-1:0] node13270;
	wire [4-1:0] node13271;
	wire [4-1:0] node13272;
	wire [4-1:0] node13274;
	wire [4-1:0] node13276;
	wire [4-1:0] node13279;
	wire [4-1:0] node13281;
	wire [4-1:0] node13283;
	wire [4-1:0] node13285;
	wire [4-1:0] node13288;
	wire [4-1:0] node13289;
	wire [4-1:0] node13290;
	wire [4-1:0] node13291;
	wire [4-1:0] node13292;
	wire [4-1:0] node13296;
	wire [4-1:0] node13299;
	wire [4-1:0] node13301;
	wire [4-1:0] node13304;
	wire [4-1:0] node13305;
	wire [4-1:0] node13306;
	wire [4-1:0] node13307;
	wire [4-1:0] node13311;
	wire [4-1:0] node13314;
	wire [4-1:0] node13315;
	wire [4-1:0] node13319;
	wire [4-1:0] node13320;
	wire [4-1:0] node13321;
	wire [4-1:0] node13322;
	wire [4-1:0] node13324;
	wire [4-1:0] node13325;
	wire [4-1:0] node13326;
	wire [4-1:0] node13329;
	wire [4-1:0] node13333;
	wire [4-1:0] node13334;
	wire [4-1:0] node13335;
	wire [4-1:0] node13336;
	wire [4-1:0] node13339;
	wire [4-1:0] node13342;
	wire [4-1:0] node13343;
	wire [4-1:0] node13344;
	wire [4-1:0] node13348;
	wire [4-1:0] node13351;
	wire [4-1:0] node13352;
	wire [4-1:0] node13355;
	wire [4-1:0] node13356;
	wire [4-1:0] node13357;
	wire [4-1:0] node13360;
	wire [4-1:0] node13364;
	wire [4-1:0] node13365;
	wire [4-1:0] node13366;
	wire [4-1:0] node13367;
	wire [4-1:0] node13369;
	wire [4-1:0] node13372;
	wire [4-1:0] node13373;
	wire [4-1:0] node13377;
	wire [4-1:0] node13378;
	wire [4-1:0] node13380;
	wire [4-1:0] node13381;
	wire [4-1:0] node13385;
	wire [4-1:0] node13386;
	wire [4-1:0] node13388;
	wire [4-1:0] node13392;
	wire [4-1:0] node13393;
	wire [4-1:0] node13395;
	wire [4-1:0] node13396;
	wire [4-1:0] node13399;
	wire [4-1:0] node13402;
	wire [4-1:0] node13403;
	wire [4-1:0] node13406;
	wire [4-1:0] node13407;
	wire [4-1:0] node13409;
	wire [4-1:0] node13413;
	wire [4-1:0] node13414;
	wire [4-1:0] node13415;
	wire [4-1:0] node13416;
	wire [4-1:0] node13417;
	wire [4-1:0] node13419;
	wire [4-1:0] node13420;
	wire [4-1:0] node13424;
	wire [4-1:0] node13425;
	wire [4-1:0] node13428;
	wire [4-1:0] node13429;
	wire [4-1:0] node13433;
	wire [4-1:0] node13434;
	wire [4-1:0] node13435;
	wire [4-1:0] node13438;
	wire [4-1:0] node13440;
	wire [4-1:0] node13443;
	wire [4-1:0] node13444;
	wire [4-1:0] node13447;
	wire [4-1:0] node13448;
	wire [4-1:0] node13452;
	wire [4-1:0] node13453;
	wire [4-1:0] node13454;
	wire [4-1:0] node13456;
	wire [4-1:0] node13457;
	wire [4-1:0] node13461;
	wire [4-1:0] node13462;
	wire [4-1:0] node13463;
	wire [4-1:0] node13468;
	wire [4-1:0] node13469;
	wire [4-1:0] node13471;
	wire [4-1:0] node13474;
	wire [4-1:0] node13475;
	wire [4-1:0] node13479;
	wire [4-1:0] node13480;
	wire [4-1:0] node13481;
	wire [4-1:0] node13482;
	wire [4-1:0] node13483;
	wire [4-1:0] node13487;
	wire [4-1:0] node13488;
	wire [4-1:0] node13492;
	wire [4-1:0] node13493;
	wire [4-1:0] node13494;
	wire [4-1:0] node13497;
	wire [4-1:0] node13498;
	wire [4-1:0] node13502;
	wire [4-1:0] node13503;
	wire [4-1:0] node13505;
	wire [4-1:0] node13508;
	wire [4-1:0] node13511;
	wire [4-1:0] node13512;
	wire [4-1:0] node13513;
	wire [4-1:0] node13514;
	wire [4-1:0] node13517;
	wire [4-1:0] node13520;
	wire [4-1:0] node13522;
	wire [4-1:0] node13523;
	wire [4-1:0] node13527;
	wire [4-1:0] node13528;
	wire [4-1:0] node13529;
	wire [4-1:0] node13532;
	wire [4-1:0] node13535;
	wire [4-1:0] node13537;
	wire [4-1:0] node13540;
	wire [4-1:0] node13541;
	wire [4-1:0] node13542;
	wire [4-1:0] node13543;
	wire [4-1:0] node13544;
	wire [4-1:0] node13545;
	wire [4-1:0] node13546;
	wire [4-1:0] node13548;
	wire [4-1:0] node13551;
	wire [4-1:0] node13553;
	wire [4-1:0] node13556;
	wire [4-1:0] node13557;
	wire [4-1:0] node13560;
	wire [4-1:0] node13561;
	wire [4-1:0] node13565;
	wire [4-1:0] node13566;
	wire [4-1:0] node13567;
	wire [4-1:0] node13568;
	wire [4-1:0] node13571;
	wire [4-1:0] node13572;
	wire [4-1:0] node13576;
	wire [4-1:0] node13577;
	wire [4-1:0] node13580;
	wire [4-1:0] node13581;
	wire [4-1:0] node13585;
	wire [4-1:0] node13586;
	wire [4-1:0] node13587;
	wire [4-1:0] node13591;
	wire [4-1:0] node13593;
	wire [4-1:0] node13596;
	wire [4-1:0] node13597;
	wire [4-1:0] node13598;
	wire [4-1:0] node13599;
	wire [4-1:0] node13602;
	wire [4-1:0] node13603;
	wire [4-1:0] node13607;
	wire [4-1:0] node13608;
	wire [4-1:0] node13610;
	wire [4-1:0] node13614;
	wire [4-1:0] node13615;
	wire [4-1:0] node13617;
	wire [4-1:0] node13620;
	wire [4-1:0] node13621;
	wire [4-1:0] node13623;
	wire [4-1:0] node13626;
	wire [4-1:0] node13627;
	wire [4-1:0] node13631;
	wire [4-1:0] node13632;
	wire [4-1:0] node13633;
	wire [4-1:0] node13634;
	wire [4-1:0] node13635;
	wire [4-1:0] node13637;
	wire [4-1:0] node13640;
	wire [4-1:0] node13641;
	wire [4-1:0] node13645;
	wire [4-1:0] node13646;
	wire [4-1:0] node13647;
	wire [4-1:0] node13648;
	wire [4-1:0] node13652;
	wire [4-1:0] node13653;
	wire [4-1:0] node13656;
	wire [4-1:0] node13659;
	wire [4-1:0] node13660;
	wire [4-1:0] node13663;
	wire [4-1:0] node13666;
	wire [4-1:0] node13667;
	wire [4-1:0] node13668;
	wire [4-1:0] node13671;
	wire [4-1:0] node13673;
	wire [4-1:0] node13676;
	wire [4-1:0] node13677;
	wire [4-1:0] node13678;
	wire [4-1:0] node13681;
	wire [4-1:0] node13685;
	wire [4-1:0] node13686;
	wire [4-1:0] node13687;
	wire [4-1:0] node13688;
	wire [4-1:0] node13690;
	wire [4-1:0] node13693;
	wire [4-1:0] node13694;
	wire [4-1:0] node13696;
	wire [4-1:0] node13699;
	wire [4-1:0] node13700;
	wire [4-1:0] node13704;
	wire [4-1:0] node13705;
	wire [4-1:0] node13706;
	wire [4-1:0] node13710;
	wire [4-1:0] node13711;
	wire [4-1:0] node13715;
	wire [4-1:0] node13716;
	wire [4-1:0] node13717;
	wire [4-1:0] node13718;
	wire [4-1:0] node13721;
	wire [4-1:0] node13724;
	wire [4-1:0] node13725;
	wire [4-1:0] node13727;
	wire [4-1:0] node13730;
	wire [4-1:0] node13731;
	wire [4-1:0] node13735;
	wire [4-1:0] node13736;
	wire [4-1:0] node13738;
	wire [4-1:0] node13741;
	wire [4-1:0] node13744;
	wire [4-1:0] node13745;
	wire [4-1:0] node13746;
	wire [4-1:0] node13747;
	wire [4-1:0] node13749;
	wire [4-1:0] node13750;
	wire [4-1:0] node13751;
	wire [4-1:0] node13756;
	wire [4-1:0] node13757;
	wire [4-1:0] node13758;
	wire [4-1:0] node13759;
	wire [4-1:0] node13763;
	wire [4-1:0] node13764;
	wire [4-1:0] node13767;
	wire [4-1:0] node13770;
	wire [4-1:0] node13771;
	wire [4-1:0] node13774;
	wire [4-1:0] node13777;
	wire [4-1:0] node13778;
	wire [4-1:0] node13779;
	wire [4-1:0] node13780;
	wire [4-1:0] node13782;
	wire [4-1:0] node13785;
	wire [4-1:0] node13786;
	wire [4-1:0] node13790;
	wire [4-1:0] node13791;
	wire [4-1:0] node13793;
	wire [4-1:0] node13796;
	wire [4-1:0] node13797;
	wire [4-1:0] node13801;
	wire [4-1:0] node13802;
	wire [4-1:0] node13804;
	wire [4-1:0] node13807;
	wire [4-1:0] node13808;
	wire [4-1:0] node13812;
	wire [4-1:0] node13813;
	wire [4-1:0] node13814;
	wire [4-1:0] node13815;
	wire [4-1:0] node13817;
	wire [4-1:0] node13820;
	wire [4-1:0] node13821;
	wire [4-1:0] node13824;
	wire [4-1:0] node13827;
	wire [4-1:0] node13828;
	wire [4-1:0] node13829;
	wire [4-1:0] node13833;
	wire [4-1:0] node13834;
	wire [4-1:0] node13837;
	wire [4-1:0] node13840;
	wire [4-1:0] node13841;
	wire [4-1:0] node13842;
	wire [4-1:0] node13844;
	wire [4-1:0] node13848;
	wire [4-1:0] node13849;
	wire [4-1:0] node13853;
	wire [4-1:0] node13854;
	wire [4-1:0] node13855;
	wire [4-1:0] node13856;
	wire [4-1:0] node13857;
	wire [4-1:0] node13858;
	wire [4-1:0] node13859;
	wire [4-1:0] node13860;
	wire [4-1:0] node13861;
	wire [4-1:0] node13863;
	wire [4-1:0] node13866;
	wire [4-1:0] node13869;
	wire [4-1:0] node13870;
	wire [4-1:0] node13875;
	wire [4-1:0] node13876;
	wire [4-1:0] node13877;
	wire [4-1:0] node13879;
	wire [4-1:0] node13880;
	wire [4-1:0] node13883;
	wire [4-1:0] node13886;
	wire [4-1:0] node13887;
	wire [4-1:0] node13890;
	wire [4-1:0] node13891;
	wire [4-1:0] node13895;
	wire [4-1:0] node13896;
	wire [4-1:0] node13898;
	wire [4-1:0] node13901;
	wire [4-1:0] node13902;
	wire [4-1:0] node13906;
	wire [4-1:0] node13907;
	wire [4-1:0] node13908;
	wire [4-1:0] node13909;
	wire [4-1:0] node13911;
	wire [4-1:0] node13914;
	wire [4-1:0] node13916;
	wire [4-1:0] node13919;
	wire [4-1:0] node13920;
	wire [4-1:0] node13921;
	wire [4-1:0] node13922;
	wire [4-1:0] node13926;
	wire [4-1:0] node13928;
	wire [4-1:0] node13931;
	wire [4-1:0] node13934;
	wire [4-1:0] node13935;
	wire [4-1:0] node13936;
	wire [4-1:0] node13938;
	wire [4-1:0] node13941;
	wire [4-1:0] node13942;
	wire [4-1:0] node13946;
	wire [4-1:0] node13947;
	wire [4-1:0] node13948;
	wire [4-1:0] node13950;
	wire [4-1:0] node13953;
	wire [4-1:0] node13956;
	wire [4-1:0] node13959;
	wire [4-1:0] node13960;
	wire [4-1:0] node13961;
	wire [4-1:0] node13962;
	wire [4-1:0] node13963;
	wire [4-1:0] node13964;
	wire [4-1:0] node13968;
	wire [4-1:0] node13969;
	wire [4-1:0] node13974;
	wire [4-1:0] node13975;
	wire [4-1:0] node13976;
	wire [4-1:0] node13978;
	wire [4-1:0] node13981;
	wire [4-1:0] node13983;
	wire [4-1:0] node13986;
	wire [4-1:0] node13987;
	wire [4-1:0] node13991;
	wire [4-1:0] node13992;
	wire [4-1:0] node13993;
	wire [4-1:0] node13994;
	wire [4-1:0] node13996;
	wire [4-1:0] node13999;
	wire [4-1:0] node14001;
	wire [4-1:0] node14004;
	wire [4-1:0] node14005;
	wire [4-1:0] node14009;
	wire [4-1:0] node14010;
	wire [4-1:0] node14011;
	wire [4-1:0] node14013;
	wire [4-1:0] node14016;
	wire [4-1:0] node14017;
	wire [4-1:0] node14021;
	wire [4-1:0] node14022;
	wire [4-1:0] node14026;
	wire [4-1:0] node14027;
	wire [4-1:0] node14028;
	wire [4-1:0] node14029;
	wire [4-1:0] node14030;
	wire [4-1:0] node14031;
	wire [4-1:0] node14032;
	wire [4-1:0] node14036;
	wire [4-1:0] node14038;
	wire [4-1:0] node14042;
	wire [4-1:0] node14043;
	wire [4-1:0] node14045;
	wire [4-1:0] node14046;
	wire [4-1:0] node14050;
	wire [4-1:0] node14052;
	wire [4-1:0] node14055;
	wire [4-1:0] node14056;
	wire [4-1:0] node14057;
	wire [4-1:0] node14058;
	wire [4-1:0] node14059;
	wire [4-1:0] node14063;
	wire [4-1:0] node14064;
	wire [4-1:0] node14068;
	wire [4-1:0] node14069;
	wire [4-1:0] node14070;
	wire [4-1:0] node14074;
	wire [4-1:0] node14076;
	wire [4-1:0] node14079;
	wire [4-1:0] node14080;
	wire [4-1:0] node14082;
	wire [4-1:0] node14083;
	wire [4-1:0] node14087;
	wire [4-1:0] node14089;
	wire [4-1:0] node14092;
	wire [4-1:0] node14093;
	wire [4-1:0] node14094;
	wire [4-1:0] node14095;
	wire [4-1:0] node14096;
	wire [4-1:0] node14097;
	wire [4-1:0] node14099;
	wire [4-1:0] node14103;
	wire [4-1:0] node14105;
	wire [4-1:0] node14108;
	wire [4-1:0] node14109;
	wire [4-1:0] node14111;
	wire [4-1:0] node14112;
	wire [4-1:0] node14116;
	wire [4-1:0] node14119;
	wire [4-1:0] node14120;
	wire [4-1:0] node14121;
	wire [4-1:0] node14123;
	wire [4-1:0] node14126;
	wire [4-1:0] node14129;
	wire [4-1:0] node14130;
	wire [4-1:0] node14131;
	wire [4-1:0] node14133;
	wire [4-1:0] node14136;
	wire [4-1:0] node14137;
	wire [4-1:0] node14141;
	wire [4-1:0] node14142;
	wire [4-1:0] node14146;
	wire [4-1:0] node14147;
	wire [4-1:0] node14148;
	wire [4-1:0] node14149;
	wire [4-1:0] node14151;
	wire [4-1:0] node14155;
	wire [4-1:0] node14156;
	wire [4-1:0] node14157;
	wire [4-1:0] node14158;
	wire [4-1:0] node14162;
	wire [4-1:0] node14164;
	wire [4-1:0] node14167;
	wire [4-1:0] node14169;
	wire [4-1:0] node14170;
	wire [4-1:0] node14173;
	wire [4-1:0] node14176;
	wire [4-1:0] node14177;
	wire [4-1:0] node14178;
	wire [4-1:0] node14181;
	wire [4-1:0] node14183;
	wire [4-1:0] node14186;
	wire [4-1:0] node14187;
	wire [4-1:0] node14189;
	wire [4-1:0] node14192;
	wire [4-1:0] node14193;
	wire [4-1:0] node14194;
	wire [4-1:0] node14198;
	wire [4-1:0] node14200;
	wire [4-1:0] node14204;
	wire [4-1:0] node14205;
	wire [4-1:0] node14206;
	wire [4-1:0] node14207;
	wire [4-1:0] node14208;
	wire [4-1:0] node14209;
	wire [4-1:0] node14210;
	wire [4-1:0] node14211;
	wire [4-1:0] node14212;
	wire [4-1:0] node14214;
	wire [4-1:0] node14218;
	wire [4-1:0] node14219;
	wire [4-1:0] node14221;
	wire [4-1:0] node14224;
	wire [4-1:0] node14225;
	wire [4-1:0] node14229;
	wire [4-1:0] node14230;
	wire [4-1:0] node14231;
	wire [4-1:0] node14232;
	wire [4-1:0] node14237;
	wire [4-1:0] node14238;
	wire [4-1:0] node14240;
	wire [4-1:0] node14243;
	wire [4-1:0] node14246;
	wire [4-1:0] node14247;
	wire [4-1:0] node14248;
	wire [4-1:0] node14249;
	wire [4-1:0] node14250;
	wire [4-1:0] node14251;
	wire [4-1:0] node14255;
	wire [4-1:0] node14258;
	wire [4-1:0] node14259;
	wire [4-1:0] node14260;
	wire [4-1:0] node14265;
	wire [4-1:0] node14267;
	wire [4-1:0] node14268;
	wire [4-1:0] node14272;
	wire [4-1:0] node14273;
	wire [4-1:0] node14274;
	wire [4-1:0] node14275;
	wire [4-1:0] node14277;
	wire [4-1:0] node14280;
	wire [4-1:0] node14281;
	wire [4-1:0] node14285;
	wire [4-1:0] node14286;
	wire [4-1:0] node14289;
	wire [4-1:0] node14290;
	wire [4-1:0] node14294;
	wire [4-1:0] node14295;
	wire [4-1:0] node14296;
	wire [4-1:0] node14299;
	wire [4-1:0] node14302;
	wire [4-1:0] node14303;
	wire [4-1:0] node14307;
	wire [4-1:0] node14308;
	wire [4-1:0] node14309;
	wire [4-1:0] node14310;
	wire [4-1:0] node14311;
	wire [4-1:0] node14312;
	wire [4-1:0] node14316;
	wire [4-1:0] node14317;
	wire [4-1:0] node14320;
	wire [4-1:0] node14322;
	wire [4-1:0] node14325;
	wire [4-1:0] node14326;
	wire [4-1:0] node14327;
	wire [4-1:0] node14330;
	wire [4-1:0] node14333;
	wire [4-1:0] node14334;
	wire [4-1:0] node14337;
	wire [4-1:0] node14339;
	wire [4-1:0] node14342;
	wire [4-1:0] node14343;
	wire [4-1:0] node14344;
	wire [4-1:0] node14346;
	wire [4-1:0] node14347;
	wire [4-1:0] node14351;
	wire [4-1:0] node14354;
	wire [4-1:0] node14355;
	wire [4-1:0] node14357;
	wire [4-1:0] node14360;
	wire [4-1:0] node14361;
	wire [4-1:0] node14364;
	wire [4-1:0] node14366;
	wire [4-1:0] node14369;
	wire [4-1:0] node14370;
	wire [4-1:0] node14371;
	wire [4-1:0] node14373;
	wire [4-1:0] node14376;
	wire [4-1:0] node14377;
	wire [4-1:0] node14378;
	wire [4-1:0] node14381;
	wire [4-1:0] node14384;
	wire [4-1:0] node14386;
	wire [4-1:0] node14389;
	wire [4-1:0] node14390;
	wire [4-1:0] node14392;
	wire [4-1:0] node14393;
	wire [4-1:0] node14397;
	wire [4-1:0] node14398;
	wire [4-1:0] node14402;
	wire [4-1:0] node14403;
	wire [4-1:0] node14404;
	wire [4-1:0] node14405;
	wire [4-1:0] node14406;
	wire [4-1:0] node14407;
	wire [4-1:0] node14408;
	wire [4-1:0] node14412;
	wire [4-1:0] node14413;
	wire [4-1:0] node14416;
	wire [4-1:0] node14419;
	wire [4-1:0] node14420;
	wire [4-1:0] node14423;
	wire [4-1:0] node14424;
	wire [4-1:0] node14428;
	wire [4-1:0] node14429;
	wire [4-1:0] node14430;
	wire [4-1:0] node14431;
	wire [4-1:0] node14432;
	wire [4-1:0] node14437;
	wire [4-1:0] node14439;
	wire [4-1:0] node14440;
	wire [4-1:0] node14444;
	wire [4-1:0] node14445;
	wire [4-1:0] node14448;
	wire [4-1:0] node14449;
	wire [4-1:0] node14453;
	wire [4-1:0] node14454;
	wire [4-1:0] node14455;
	wire [4-1:0] node14456;
	wire [4-1:0] node14459;
	wire [4-1:0] node14461;
	wire [4-1:0] node14464;
	wire [4-1:0] node14465;
	wire [4-1:0] node14466;
	wire [4-1:0] node14470;
	wire [4-1:0] node14472;
	wire [4-1:0] node14475;
	wire [4-1:0] node14476;
	wire [4-1:0] node14477;
	wire [4-1:0] node14478;
	wire [4-1:0] node14479;
	wire [4-1:0] node14483;
	wire [4-1:0] node14486;
	wire [4-1:0] node14487;
	wire [4-1:0] node14489;
	wire [4-1:0] node14492;
	wire [4-1:0] node14495;
	wire [4-1:0] node14496;
	wire [4-1:0] node14498;
	wire [4-1:0] node14501;
	wire [4-1:0] node14502;
	wire [4-1:0] node14504;
	wire [4-1:0] node14507;
	wire [4-1:0] node14510;
	wire [4-1:0] node14511;
	wire [4-1:0] node14512;
	wire [4-1:0] node14513;
	wire [4-1:0] node14514;
	wire [4-1:0] node14516;
	wire [4-1:0] node14519;
	wire [4-1:0] node14520;
	wire [4-1:0] node14523;
	wire [4-1:0] node14526;
	wire [4-1:0] node14527;
	wire [4-1:0] node14528;
	wire [4-1:0] node14531;
	wire [4-1:0] node14532;
	wire [4-1:0] node14536;
	wire [4-1:0] node14537;
	wire [4-1:0] node14538;
	wire [4-1:0] node14542;
	wire [4-1:0] node14545;
	wire [4-1:0] node14546;
	wire [4-1:0] node14547;
	wire [4-1:0] node14548;
	wire [4-1:0] node14549;
	wire [4-1:0] node14553;
	wire [4-1:0] node14554;
	wire [4-1:0] node14557;
	wire [4-1:0] node14560;
	wire [4-1:0] node14561;
	wire [4-1:0] node14565;
	wire [4-1:0] node14566;
	wire [4-1:0] node14567;
	wire [4-1:0] node14571;
	wire [4-1:0] node14573;
	wire [4-1:0] node14577;
	wire [4-1:0] node14578;
	wire [4-1:0] node14579;
	wire [4-1:0] node14580;
	wire [4-1:0] node14581;
	wire [4-1:0] node14582;
	wire [4-1:0] node14583;
	wire [4-1:0] node14585;
	wire [4-1:0] node14588;
	wire [4-1:0] node14589;
	wire [4-1:0] node14593;
	wire [4-1:0] node14594;
	wire [4-1:0] node14595;
	wire [4-1:0] node14599;
	wire [4-1:0] node14600;
	wire [4-1:0] node14603;
	wire [4-1:0] node14604;
	wire [4-1:0] node14608;
	wire [4-1:0] node14609;
	wire [4-1:0] node14610;
	wire [4-1:0] node14611;
	wire [4-1:0] node14612;
	wire [4-1:0] node14615;
	wire [4-1:0] node14619;
	wire [4-1:0] node14620;
	wire [4-1:0] node14623;
	wire [4-1:0] node14626;
	wire [4-1:0] node14627;
	wire [4-1:0] node14630;
	wire [4-1:0] node14631;
	wire [4-1:0] node14632;
	wire [4-1:0] node14637;
	wire [4-1:0] node14638;
	wire [4-1:0] node14639;
	wire [4-1:0] node14641;
	wire [4-1:0] node14642;
	wire [4-1:0] node14644;
	wire [4-1:0] node14647;
	wire [4-1:0] node14650;
	wire [4-1:0] node14652;
	wire [4-1:0] node14653;
	wire [4-1:0] node14654;
	wire [4-1:0] node14658;
	wire [4-1:0] node14661;
	wire [4-1:0] node14662;
	wire [4-1:0] node14663;
	wire [4-1:0] node14664;
	wire [4-1:0] node14667;
	wire [4-1:0] node14670;
	wire [4-1:0] node14672;
	wire [4-1:0] node14675;
	wire [4-1:0] node14676;
	wire [4-1:0] node14677;
	wire [4-1:0] node14678;
	wire [4-1:0] node14682;
	wire [4-1:0] node14685;
	wire [4-1:0] node14686;
	wire [4-1:0] node14689;
	wire [4-1:0] node14691;
	wire [4-1:0] node14694;
	wire [4-1:0] node14695;
	wire [4-1:0] node14696;
	wire [4-1:0] node14697;
	wire [4-1:0] node14698;
	wire [4-1:0] node14699;
	wire [4-1:0] node14701;
	wire [4-1:0] node14704;
	wire [4-1:0] node14706;
	wire [4-1:0] node14709;
	wire [4-1:0] node14710;
	wire [4-1:0] node14712;
	wire [4-1:0] node14715;
	wire [4-1:0] node14718;
	wire [4-1:0] node14719;
	wire [4-1:0] node14720;
	wire [4-1:0] node14721;
	wire [4-1:0] node14726;
	wire [4-1:0] node14727;
	wire [4-1:0] node14729;
	wire [4-1:0] node14733;
	wire [4-1:0] node14734;
	wire [4-1:0] node14735;
	wire [4-1:0] node14737;
	wire [4-1:0] node14738;
	wire [4-1:0] node14742;
	wire [4-1:0] node14743;
	wire [4-1:0] node14744;
	wire [4-1:0] node14748;
	wire [4-1:0] node14749;
	wire [4-1:0] node14753;
	wire [4-1:0] node14754;
	wire [4-1:0] node14755;
	wire [4-1:0] node14758;
	wire [4-1:0] node14759;
	wire [4-1:0] node14763;
	wire [4-1:0] node14766;
	wire [4-1:0] node14767;
	wire [4-1:0] node14768;
	wire [4-1:0] node14769;
	wire [4-1:0] node14770;
	wire [4-1:0] node14771;
	wire [4-1:0] node14775;
	wire [4-1:0] node14776;
	wire [4-1:0] node14780;
	wire [4-1:0] node14781;
	wire [4-1:0] node14785;
	wire [4-1:0] node14786;
	wire [4-1:0] node14787;
	wire [4-1:0] node14788;
	wire [4-1:0] node14793;
	wire [4-1:0] node14794;
	wire [4-1:0] node14795;
	wire [4-1:0] node14798;
	wire [4-1:0] node14801;
	wire [4-1:0] node14804;
	wire [4-1:0] node14805;
	wire [4-1:0] node14806;
	wire [4-1:0] node14808;
	wire [4-1:0] node14809;
	wire [4-1:0] node14813;
	wire [4-1:0] node14814;
	wire [4-1:0] node14817;
	wire [4-1:0] node14818;
	wire [4-1:0] node14822;
	wire [4-1:0] node14823;
	wire [4-1:0] node14824;
	wire [4-1:0] node14827;
	wire [4-1:0] node14830;
	wire [4-1:0] node14831;
	wire [4-1:0] node14834;
	wire [4-1:0] node14837;
	wire [4-1:0] node14838;
	wire [4-1:0] node14839;
	wire [4-1:0] node14840;
	wire [4-1:0] node14841;
	wire [4-1:0] node14843;
	wire [4-1:0] node14845;
	wire [4-1:0] node14848;
	wire [4-1:0] node14850;
	wire [4-1:0] node14851;
	wire [4-1:0] node14855;
	wire [4-1:0] node14856;
	wire [4-1:0] node14857;
	wire [4-1:0] node14860;
	wire [4-1:0] node14863;
	wire [4-1:0] node14864;
	wire [4-1:0] node14865;
	wire [4-1:0] node14869;
	wire [4-1:0] node14870;
	wire [4-1:0] node14873;
	wire [4-1:0] node14876;
	wire [4-1:0] node14877;
	wire [4-1:0] node14878;
	wire [4-1:0] node14879;
	wire [4-1:0] node14880;
	wire [4-1:0] node14884;
	wire [4-1:0] node14885;
	wire [4-1:0] node14888;
	wire [4-1:0] node14891;
	wire [4-1:0] node14892;
	wire [4-1:0] node14894;
	wire [4-1:0] node14897;
	wire [4-1:0] node14899;
	wire [4-1:0] node14902;
	wire [4-1:0] node14903;
	wire [4-1:0] node14904;
	wire [4-1:0] node14906;
	wire [4-1:0] node14910;
	wire [4-1:0] node14912;
	wire [4-1:0] node14915;
	wire [4-1:0] node14916;
	wire [4-1:0] node14917;
	wire [4-1:0] node14918;
	wire [4-1:0] node14919;
	wire [4-1:0] node14923;
	wire [4-1:0] node14924;
	wire [4-1:0] node14926;
	wire [4-1:0] node14929;
	wire [4-1:0] node14930;
	wire [4-1:0] node14931;
	wire [4-1:0] node14934;
	wire [4-1:0] node14938;
	wire [4-1:0] node14939;
	wire [4-1:0] node14940;
	wire [4-1:0] node14941;
	wire [4-1:0] node14945;
	wire [4-1:0] node14948;
	wire [4-1:0] node14949;
	wire [4-1:0] node14950;
	wire [4-1:0] node14953;
	wire [4-1:0] node14956;
	wire [4-1:0] node14958;
	wire [4-1:0] node14961;
	wire [4-1:0] node14962;
	wire [4-1:0] node14963;
	wire [4-1:0] node14965;
	wire [4-1:0] node14968;
	wire [4-1:0] node14970;
	wire [4-1:0] node14974;
	wire [4-1:0] node14975;
	wire [4-1:0] node14976;
	wire [4-1:0] node14977;
	wire [4-1:0] node14978;
	wire [4-1:0] node14979;
	wire [4-1:0] node14980;
	wire [4-1:0] node14981;
	wire [4-1:0] node14983;
	wire [4-1:0] node14986;
	wire [4-1:0] node14987;
	wire [4-1:0] node14990;
	wire [4-1:0] node14991;
	wire [4-1:0] node14995;
	wire [4-1:0] node14996;
	wire [4-1:0] node14997;
	wire [4-1:0] node14998;
	wire [4-1:0] node15002;
	wire [4-1:0] node15004;
	wire [4-1:0] node15007;
	wire [4-1:0] node15008;
	wire [4-1:0] node15011;
	wire [4-1:0] node15014;
	wire [4-1:0] node15015;
	wire [4-1:0] node15016;
	wire [4-1:0] node15018;
	wire [4-1:0] node15021;
	wire [4-1:0] node15022;
	wire [4-1:0] node15025;
	wire [4-1:0] node15028;
	wire [4-1:0] node15030;
	wire [4-1:0] node15031;
	wire [4-1:0] node15033;
	wire [4-1:0] node15037;
	wire [4-1:0] node15038;
	wire [4-1:0] node15039;
	wire [4-1:0] node15040;
	wire [4-1:0] node15041;
	wire [4-1:0] node15042;
	wire [4-1:0] node15045;
	wire [4-1:0] node15049;
	wire [4-1:0] node15051;
	wire [4-1:0] node15054;
	wire [4-1:0] node15055;
	wire [4-1:0] node15056;
	wire [4-1:0] node15059;
	wire [4-1:0] node15060;
	wire [4-1:0] node15064;
	wire [4-1:0] node15065;
	wire [4-1:0] node15066;
	wire [4-1:0] node15069;
	wire [4-1:0] node15072;
	wire [4-1:0] node15073;
	wire [4-1:0] node15076;
	wire [4-1:0] node15079;
	wire [4-1:0] node15080;
	wire [4-1:0] node15081;
	wire [4-1:0] node15082;
	wire [4-1:0] node15085;
	wire [4-1:0] node15088;
	wire [4-1:0] node15089;
	wire [4-1:0] node15092;
	wire [4-1:0] node15095;
	wire [4-1:0] node15096;
	wire [4-1:0] node15098;
	wire [4-1:0] node15101;
	wire [4-1:0] node15102;
	wire [4-1:0] node15106;
	wire [4-1:0] node15107;
	wire [4-1:0] node15108;
	wire [4-1:0] node15109;
	wire [4-1:0] node15110;
	wire [4-1:0] node15111;
	wire [4-1:0] node15114;
	wire [4-1:0] node15115;
	wire [4-1:0] node15119;
	wire [4-1:0] node15120;
	wire [4-1:0] node15121;
	wire [4-1:0] node15125;
	wire [4-1:0] node15126;
	wire [4-1:0] node15130;
	wire [4-1:0] node15131;
	wire [4-1:0] node15133;
	wire [4-1:0] node15134;
	wire [4-1:0] node15138;
	wire [4-1:0] node15140;
	wire [4-1:0] node15143;
	wire [4-1:0] node15144;
	wire [4-1:0] node15145;
	wire [4-1:0] node15146;
	wire [4-1:0] node15149;
	wire [4-1:0] node15151;
	wire [4-1:0] node15154;
	wire [4-1:0] node15155;
	wire [4-1:0] node15156;
	wire [4-1:0] node15159;
	wire [4-1:0] node15163;
	wire [4-1:0] node15164;
	wire [4-1:0] node15165;
	wire [4-1:0] node15166;
	wire [4-1:0] node15169;
	wire [4-1:0] node15172;
	wire [4-1:0] node15173;
	wire [4-1:0] node15177;
	wire [4-1:0] node15178;
	wire [4-1:0] node15180;
	wire [4-1:0] node15183;
	wire [4-1:0] node15186;
	wire [4-1:0] node15187;
	wire [4-1:0] node15188;
	wire [4-1:0] node15189;
	wire [4-1:0] node15191;
	wire [4-1:0] node15193;
	wire [4-1:0] node15197;
	wire [4-1:0] node15198;
	wire [4-1:0] node15201;
	wire [4-1:0] node15203;
	wire [4-1:0] node15204;
	wire [4-1:0] node15208;
	wire [4-1:0] node15209;
	wire [4-1:0] node15210;
	wire [4-1:0] node15211;
	wire [4-1:0] node15215;
	wire [4-1:0] node15216;
	wire [4-1:0] node15219;
	wire [4-1:0] node15220;
	wire [4-1:0] node15223;
	wire [4-1:0] node15226;
	wire [4-1:0] node15227;
	wire [4-1:0] node15228;
	wire [4-1:0] node15231;
	wire [4-1:0] node15234;
	wire [4-1:0] node15236;
	wire [4-1:0] node15239;
	wire [4-1:0] node15240;
	wire [4-1:0] node15241;
	wire [4-1:0] node15242;
	wire [4-1:0] node15243;
	wire [4-1:0] node15244;
	wire [4-1:0] node15247;
	wire [4-1:0] node15248;
	wire [4-1:0] node15250;
	wire [4-1:0] node15253;
	wire [4-1:0] node15254;
	wire [4-1:0] node15258;
	wire [4-1:0] node15259;
	wire [4-1:0] node15260;
	wire [4-1:0] node15264;
	wire [4-1:0] node15265;
	wire [4-1:0] node15268;
	wire [4-1:0] node15271;
	wire [4-1:0] node15272;
	wire [4-1:0] node15274;
	wire [4-1:0] node15275;
	wire [4-1:0] node15278;
	wire [4-1:0] node15281;
	wire [4-1:0] node15282;
	wire [4-1:0] node15283;
	wire [4-1:0] node15286;
	wire [4-1:0] node15289;
	wire [4-1:0] node15290;
	wire [4-1:0] node15293;
	wire [4-1:0] node15296;
	wire [4-1:0] node15297;
	wire [4-1:0] node15298;
	wire [4-1:0] node15299;
	wire [4-1:0] node15300;
	wire [4-1:0] node15304;
	wire [4-1:0] node15307;
	wire [4-1:0] node15308;
	wire [4-1:0] node15309;
	wire [4-1:0] node15312;
	wire [4-1:0] node15315;
	wire [4-1:0] node15317;
	wire [4-1:0] node15320;
	wire [4-1:0] node15321;
	wire [4-1:0] node15322;
	wire [4-1:0] node15324;
	wire [4-1:0] node15327;
	wire [4-1:0] node15328;
	wire [4-1:0] node15331;
	wire [4-1:0] node15334;
	wire [4-1:0] node15335;
	wire [4-1:0] node15337;
	wire [4-1:0] node15340;
	wire [4-1:0] node15341;
	wire [4-1:0] node15344;
	wire [4-1:0] node15347;
	wire [4-1:0] node15348;
	wire [4-1:0] node15349;
	wire [4-1:0] node15350;
	wire [4-1:0] node15351;
	wire [4-1:0] node15352;
	wire [4-1:0] node15353;
	wire [4-1:0] node15358;
	wire [4-1:0] node15359;
	wire [4-1:0] node15362;
	wire [4-1:0] node15365;
	wire [4-1:0] node15366;
	wire [4-1:0] node15369;
	wire [4-1:0] node15372;
	wire [4-1:0] node15374;
	wire [4-1:0] node15376;
	wire [4-1:0] node15377;
	wire [4-1:0] node15379;
	wire [4-1:0] node15382;
	wire [4-1:0] node15385;
	wire [4-1:0] node15386;
	wire [4-1:0] node15387;
	wire [4-1:0] node15388;
	wire [4-1:0] node15390;
	wire [4-1:0] node15393;
	wire [4-1:0] node15394;
	wire [4-1:0] node15398;
	wire [4-1:0] node15399;
	wire [4-1:0] node15401;
	wire [4-1:0] node15402;
	wire [4-1:0] node15408;
	wire [4-1:0] node15409;
	wire [4-1:0] node15410;
	wire [4-1:0] node15411;
	wire [4-1:0] node15412;
	wire [4-1:0] node15413;
	wire [4-1:0] node15414;
	wire [4-1:0] node15416;
	wire [4-1:0] node15419;
	wire [4-1:0] node15421;
	wire [4-1:0] node15424;
	wire [4-1:0] node15425;
	wire [4-1:0] node15426;
	wire [4-1:0] node15428;
	wire [4-1:0] node15431;
	wire [4-1:0] node15434;
	wire [4-1:0] node15436;
	wire [4-1:0] node15439;
	wire [4-1:0] node15440;
	wire [4-1:0] node15441;
	wire [4-1:0] node15443;
	wire [4-1:0] node15445;
	wire [4-1:0] node15448;
	wire [4-1:0] node15449;
	wire [4-1:0] node15450;
	wire [4-1:0] node15453;
	wire [4-1:0] node15457;
	wire [4-1:0] node15458;
	wire [4-1:0] node15461;
	wire [4-1:0] node15462;
	wire [4-1:0] node15464;
	wire [4-1:0] node15467;
	wire [4-1:0] node15468;
	wire [4-1:0] node15472;
	wire [4-1:0] node15473;
	wire [4-1:0] node15474;
	wire [4-1:0] node15475;
	wire [4-1:0] node15476;
	wire [4-1:0] node15480;
	wire [4-1:0] node15481;
	wire [4-1:0] node15485;
	wire [4-1:0] node15486;
	wire [4-1:0] node15487;
	wire [4-1:0] node15490;
	wire [4-1:0] node15493;
	wire [4-1:0] node15495;
	wire [4-1:0] node15498;
	wire [4-1:0] node15499;
	wire [4-1:0] node15500;
	wire [4-1:0] node15502;
	wire [4-1:0] node15503;
	wire [4-1:0] node15507;
	wire [4-1:0] node15508;
	wire [4-1:0] node15510;
	wire [4-1:0] node15513;
	wire [4-1:0] node15514;
	wire [4-1:0] node15518;
	wire [4-1:0] node15519;
	wire [4-1:0] node15521;
	wire [4-1:0] node15524;
	wire [4-1:0] node15525;
	wire [4-1:0] node15527;
	wire [4-1:0] node15531;
	wire [4-1:0] node15532;
	wire [4-1:0] node15533;
	wire [4-1:0] node15534;
	wire [4-1:0] node15535;
	wire [4-1:0] node15536;
	wire [4-1:0] node15539;
	wire [4-1:0] node15542;
	wire [4-1:0] node15543;
	wire [4-1:0] node15546;
	wire [4-1:0] node15549;
	wire [4-1:0] node15550;
	wire [4-1:0] node15553;
	wire [4-1:0] node15554;
	wire [4-1:0] node15558;
	wire [4-1:0] node15559;
	wire [4-1:0] node15560;
	wire [4-1:0] node15563;
	wire [4-1:0] node15565;
	wire [4-1:0] node15568;
	wire [4-1:0] node15569;
	wire [4-1:0] node15570;
	wire [4-1:0] node15574;
	wire [4-1:0] node15576;
	wire [4-1:0] node15577;
	wire [4-1:0] node15581;
	wire [4-1:0] node15582;
	wire [4-1:0] node15583;
	wire [4-1:0] node15584;
	wire [4-1:0] node15585;
	wire [4-1:0] node15589;
	wire [4-1:0] node15590;
	wire [4-1:0] node15591;
	wire [4-1:0] node15594;
	wire [4-1:0] node15597;
	wire [4-1:0] node15598;
	wire [4-1:0] node15602;
	wire [4-1:0] node15603;
	wire [4-1:0] node15604;
	wire [4-1:0] node15607;
	wire [4-1:0] node15610;
	wire [4-1:0] node15612;
	wire [4-1:0] node15616;
	wire [4-1:0] node15617;
	wire [4-1:0] node15618;
	wire [4-1:0] node15619;
	wire [4-1:0] node15620;
	wire [4-1:0] node15621;
	wire [4-1:0] node15625;
	wire [4-1:0] node15626;
	wire [4-1:0] node15627;
	wire [4-1:0] node15631;
	wire [4-1:0] node15632;
	wire [4-1:0] node15634;
	wire [4-1:0] node15638;
	wire [4-1:0] node15639;
	wire [4-1:0] node15640;
	wire [4-1:0] node15641;
	wire [4-1:0] node15642;
	wire [4-1:0] node15645;
	wire [4-1:0] node15649;
	wire [4-1:0] node15650;
	wire [4-1:0] node15651;
	wire [4-1:0] node15655;
	wire [4-1:0] node15658;
	wire [4-1:0] node15660;
	wire [4-1:0] node15661;
	wire [4-1:0] node15662;
	wire [4-1:0] node15665;
	wire [4-1:0] node15669;
	wire [4-1:0] node15670;
	wire [4-1:0] node15671;
	wire [4-1:0] node15672;
	wire [4-1:0] node15673;
	wire [4-1:0] node15674;
	wire [4-1:0] node15678;
	wire [4-1:0] node15681;
	wire [4-1:0] node15683;
	wire [4-1:0] node15685;
	wire [4-1:0] node15688;
	wire [4-1:0] node15689;
	wire [4-1:0] node15691;
	wire [4-1:0] node15694;
	wire [4-1:0] node15695;
	wire [4-1:0] node15700;
	wire [4-1:0] node15701;
	wire [4-1:0] node15702;
	wire [4-1:0] node15703;
	wire [4-1:0] node15704;
	wire [4-1:0] node15705;
	wire [4-1:0] node15707;
	wire [4-1:0] node15711;
	wire [4-1:0] node15712;
	wire [4-1:0] node15714;
	wire [4-1:0] node15717;
	wire [4-1:0] node15719;
	wire [4-1:0] node15722;
	wire [4-1:0] node15723;
	wire [4-1:0] node15724;
	wire [4-1:0] node15726;
	wire [4-1:0] node15730;
	wire [4-1:0] node15731;
	wire [4-1:0] node15732;
	wire [4-1:0] node15736;
	wire [4-1:0] node15737;
	wire [4-1:0] node15743;
	wire [4-1:0] node15744;
	wire [4-1:0] node15745;
	wire [4-1:0] node15746;
	wire [4-1:0] node15748;
	wire [4-1:0] node15749;
	wire [4-1:0] node15750;
	wire [4-1:0] node15751;
	wire [4-1:0] node15752;
	wire [4-1:0] node15753;
	wire [4-1:0] node15754;
	wire [4-1:0] node15757;
	wire [4-1:0] node15758;
	wire [4-1:0] node15761;
	wire [4-1:0] node15762;
	wire [4-1:0] node15766;
	wire [4-1:0] node15768;
	wire [4-1:0] node15770;
	wire [4-1:0] node15771;
	wire [4-1:0] node15775;
	wire [4-1:0] node15776;
	wire [4-1:0] node15777;
	wire [4-1:0] node15780;
	wire [4-1:0] node15783;
	wire [4-1:0] node15784;
	wire [4-1:0] node15785;
	wire [4-1:0] node15786;
	wire [4-1:0] node15790;
	wire [4-1:0] node15791;
	wire [4-1:0] node15795;
	wire [4-1:0] node15796;
	wire [4-1:0] node15801;
	wire [4-1:0] node15802;
	wire [4-1:0] node15803;
	wire [4-1:0] node15804;
	wire [4-1:0] node15805;
	wire [4-1:0] node15807;
	wire [4-1:0] node15810;
	wire [4-1:0] node15812;
	wire [4-1:0] node15815;
	wire [4-1:0] node15817;
	wire [4-1:0] node15820;
	wire [4-1:0] node15821;
	wire [4-1:0] node15823;
	wire [4-1:0] node15825;
	wire [4-1:0] node15828;
	wire [4-1:0] node15829;
	wire [4-1:0] node15833;
	wire [4-1:0] node15834;
	wire [4-1:0] node15835;
	wire [4-1:0] node15836;
	wire [4-1:0] node15837;
	wire [4-1:0] node15838;
	wire [4-1:0] node15841;
	wire [4-1:0] node15844;
	wire [4-1:0] node15846;
	wire [4-1:0] node15849;
	wire [4-1:0] node15852;
	wire [4-1:0] node15853;
	wire [4-1:0] node15854;
	wire [4-1:0] node15857;
	wire [4-1:0] node15858;
	wire [4-1:0] node15862;
	wire [4-1:0] node15864;
	wire [4-1:0] node15867;
	wire [4-1:0] node15868;
	wire [4-1:0] node15870;
	wire [4-1:0] node15871;
	wire [4-1:0] node15875;
	wire [4-1:0] node15877;
	wire [4-1:0] node15881;
	wire [4-1:0] node15882;
	wire [4-1:0] node15883;
	wire [4-1:0] node15884;
	wire [4-1:0] node15885;
	wire [4-1:0] node15886;
	wire [4-1:0] node15887;
	wire [4-1:0] node15888;
	wire [4-1:0] node15890;
	wire [4-1:0] node15893;
	wire [4-1:0] node15895;
	wire [4-1:0] node15898;
	wire [4-1:0] node15899;
	wire [4-1:0] node15901;
	wire [4-1:0] node15904;
	wire [4-1:0] node15905;
	wire [4-1:0] node15909;
	wire [4-1:0] node15910;
	wire [4-1:0] node15912;
	wire [4-1:0] node15915;
	wire [4-1:0] node15916;
	wire [4-1:0] node15920;
	wire [4-1:0] node15921;
	wire [4-1:0] node15922;
	wire [4-1:0] node15923;
	wire [4-1:0] node15924;
	wire [4-1:0] node15929;
	wire [4-1:0] node15930;
	wire [4-1:0] node15932;
	wire [4-1:0] node15935;
	wire [4-1:0] node15936;
	wire [4-1:0] node15940;
	wire [4-1:0] node15941;
	wire [4-1:0] node15943;
	wire [4-1:0] node15946;
	wire [4-1:0] node15948;
	wire [4-1:0] node15951;
	wire [4-1:0] node15952;
	wire [4-1:0] node15953;
	wire [4-1:0] node15954;
	wire [4-1:0] node15955;
	wire [4-1:0] node15956;
	wire [4-1:0] node15957;
	wire [4-1:0] node15960;
	wire [4-1:0] node15964;
	wire [4-1:0] node15965;
	wire [4-1:0] node15967;
	wire [4-1:0] node15971;
	wire [4-1:0] node15973;
	wire [4-1:0] node15974;
	wire [4-1:0] node15978;
	wire [4-1:0] node15979;
	wire [4-1:0] node15980;
	wire [4-1:0] node15981;
	wire [4-1:0] node15985;
	wire [4-1:0] node15987;
	wire [4-1:0] node15990;
	wire [4-1:0] node15991;
	wire [4-1:0] node15992;
	wire [4-1:0] node15994;
	wire [4-1:0] node15997;
	wire [4-1:0] node16000;
	wire [4-1:0] node16001;
	wire [4-1:0] node16004;
	wire [4-1:0] node16007;
	wire [4-1:0] node16008;
	wire [4-1:0] node16009;
	wire [4-1:0] node16010;
	wire [4-1:0] node16012;
	wire [4-1:0] node16015;
	wire [4-1:0] node16016;
	wire [4-1:0] node16019;
	wire [4-1:0] node16020;
	wire [4-1:0] node16024;
	wire [4-1:0] node16025;
	wire [4-1:0] node16028;
	wire [4-1:0] node16029;
	wire [4-1:0] node16032;
	wire [4-1:0] node16035;
	wire [4-1:0] node16036;
	wire [4-1:0] node16037;
	wire [4-1:0] node16038;
	wire [4-1:0] node16042;
	wire [4-1:0] node16043;
	wire [4-1:0] node16047;
	wire [4-1:0] node16048;
	wire [4-1:0] node16049;
	wire [4-1:0] node16051;
	wire [4-1:0] node16054;
	wire [4-1:0] node16056;
	wire [4-1:0] node16059;
	wire [4-1:0] node16061;
	wire [4-1:0] node16064;
	wire [4-1:0] node16065;
	wire [4-1:0] node16066;
	wire [4-1:0] node16067;
	wire [4-1:0] node16068;
	wire [4-1:0] node16069;
	wire [4-1:0] node16071;
	wire [4-1:0] node16075;
	wire [4-1:0] node16076;
	wire [4-1:0] node16077;
	wire [4-1:0] node16081;
	wire [4-1:0] node16083;
	wire [4-1:0] node16086;
	wire [4-1:0] node16087;
	wire [4-1:0] node16089;
	wire [4-1:0] node16092;
	wire [4-1:0] node16094;
	wire [4-1:0] node16097;
	wire [4-1:0] node16098;
	wire [4-1:0] node16099;
	wire [4-1:0] node16101;
	wire [4-1:0] node16104;
	wire [4-1:0] node16105;
	wire [4-1:0] node16109;
	wire [4-1:0] node16110;
	wire [4-1:0] node16111;
	wire [4-1:0] node16113;
	wire [4-1:0] node16116;
	wire [4-1:0] node16117;
	wire [4-1:0] node16121;
	wire [4-1:0] node16123;
	wire [4-1:0] node16126;
	wire [4-1:0] node16127;
	wire [4-1:0] node16128;
	wire [4-1:0] node16129;
	wire [4-1:0] node16130;
	wire [4-1:0] node16131;
	wire [4-1:0] node16135;
	wire [4-1:0] node16137;
	wire [4-1:0] node16140;
	wire [4-1:0] node16141;
	wire [4-1:0] node16142;
	wire [4-1:0] node16143;
	wire [4-1:0] node16147;
	wire [4-1:0] node16149;
	wire [4-1:0] node16152;
	wire [4-1:0] node16154;
	wire [4-1:0] node16155;
	wire [4-1:0] node16159;
	wire [4-1:0] node16160;
	wire [4-1:0] node16161;
	wire [4-1:0] node16163;
	wire [4-1:0] node16166;
	wire [4-1:0] node16167;
	wire [4-1:0] node16171;
	wire [4-1:0] node16172;
	wire [4-1:0] node16174;
	wire [4-1:0] node16177;
	wire [4-1:0] node16179;
	wire [4-1:0] node16182;
	wire [4-1:0] node16183;
	wire [4-1:0] node16184;
	wire [4-1:0] node16185;
	wire [4-1:0] node16186;
	wire [4-1:0] node16190;
	wire [4-1:0] node16191;
	wire [4-1:0] node16195;
	wire [4-1:0] node16196;
	wire [4-1:0] node16198;
	wire [4-1:0] node16199;
	wire [4-1:0] node16202;
	wire [4-1:0] node16205;
	wire [4-1:0] node16206;
	wire [4-1:0] node16210;
	wire [4-1:0] node16211;
	wire [4-1:0] node16212;
	wire [4-1:0] node16213;
	wire [4-1:0] node16217;
	wire [4-1:0] node16218;
	wire [4-1:0] node16222;
	wire [4-1:0] node16223;
	wire [4-1:0] node16225;
	wire [4-1:0] node16228;
	wire [4-1:0] node16229;
	wire [4-1:0] node16233;
	wire [4-1:0] node16235;
	wire [4-1:0] node16236;
	wire [4-1:0] node16237;
	wire [4-1:0] node16238;
	wire [4-1:0] node16239;
	wire [4-1:0] node16241;
	wire [4-1:0] node16242;
	wire [4-1:0] node16244;
	wire [4-1:0] node16248;
	wire [4-1:0] node16249;
	wire [4-1:0] node16252;
	wire [4-1:0] node16254;
	wire [4-1:0] node16257;
	wire [4-1:0] node16258;
	wire [4-1:0] node16260;
	wire [4-1:0] node16262;
	wire [4-1:0] node16265;
	wire [4-1:0] node16266;
	wire [4-1:0] node16270;
	wire [4-1:0] node16271;
	wire [4-1:0] node16272;
	wire [4-1:0] node16273;
	wire [4-1:0] node16274;
	wire [4-1:0] node16278;
	wire [4-1:0] node16280;
	wire [4-1:0] node16283;
	wire [4-1:0] node16284;
	wire [4-1:0] node16287;
	wire [4-1:0] node16289;
	wire [4-1:0] node16292;
	wire [4-1:0] node16293;
	wire [4-1:0] node16294;
	wire [4-1:0] node16296;
	wire [4-1:0] node16300;
	wire [4-1:0] node16302;
	wire [4-1:0] node16305;
	wire [4-1:0] node16307;
	wire [4-1:0] node16308;
	wire [4-1:0] node16309;
	wire [4-1:0] node16310;
	wire [4-1:0] node16312;
	wire [4-1:0] node16315;
	wire [4-1:0] node16318;
	wire [4-1:0] node16320;
	wire [4-1:0] node16322;
	wire [4-1:0] node16324;
	wire [4-1:0] node16327;
	wire [4-1:0] node16328;
	wire [4-1:0] node16329;
	wire [4-1:0] node16330;
	wire [4-1:0] node16332;
	wire [4-1:0] node16335;
	wire [4-1:0] node16339;
	wire [4-1:0] node16340;
	wire [4-1:0] node16341;
	wire [4-1:0] node16345;
	wire [4-1:0] node16346;
	wire [4-1:0] node16347;
	wire [4-1:0] node16352;
	wire [4-1:0] node16353;
	wire [4-1:0] node16354;
	wire [4-1:0] node16355;
	wire [4-1:0] node16356;
	wire [4-1:0] node16357;
	wire [4-1:0] node16358;
	wire [4-1:0] node16359;
	wire [4-1:0] node16363;
	wire [4-1:0] node16364;
	wire [4-1:0] node16366;
	wire [4-1:0] node16369;
	wire [4-1:0] node16370;
	wire [4-1:0] node16372;
	wire [4-1:0] node16373;
	wire [4-1:0] node16378;
	wire [4-1:0] node16379;
	wire [4-1:0] node16380;
	wire [4-1:0] node16382;
	wire [4-1:0] node16385;
	wire [4-1:0] node16387;
	wire [4-1:0] node16390;
	wire [4-1:0] node16391;
	wire [4-1:0] node16392;
	wire [4-1:0] node16393;
	wire [4-1:0] node16396;
	wire [4-1:0] node16399;
	wire [4-1:0] node16402;
	wire [4-1:0] node16404;
	wire [4-1:0] node16405;
	wire [4-1:0] node16409;
	wire [4-1:0] node16410;
	wire [4-1:0] node16411;
	wire [4-1:0] node16412;
	wire [4-1:0] node16413;
	wire [4-1:0] node16414;
	wire [4-1:0] node16417;
	wire [4-1:0] node16418;
	wire [4-1:0] node16422;
	wire [4-1:0] node16423;
	wire [4-1:0] node16424;
	wire [4-1:0] node16429;
	wire [4-1:0] node16430;
	wire [4-1:0] node16432;
	wire [4-1:0] node16433;
	wire [4-1:0] node16437;
	wire [4-1:0] node16438;
	wire [4-1:0] node16440;
	wire [4-1:0] node16443;
	wire [4-1:0] node16445;
	wire [4-1:0] node16448;
	wire [4-1:0] node16449;
	wire [4-1:0] node16450;
	wire [4-1:0] node16451;
	wire [4-1:0] node16454;
	wire [4-1:0] node16457;
	wire [4-1:0] node16458;
	wire [4-1:0] node16461;
	wire [4-1:0] node16464;
	wire [4-1:0] node16466;
	wire [4-1:0] node16468;
	wire [4-1:0] node16471;
	wire [4-1:0] node16472;
	wire [4-1:0] node16473;
	wire [4-1:0] node16475;
	wire [4-1:0] node16476;
	wire [4-1:0] node16477;
	wire [4-1:0] node16481;
	wire [4-1:0] node16484;
	wire [4-1:0] node16485;
	wire [4-1:0] node16487;
	wire [4-1:0] node16489;
	wire [4-1:0] node16492;
	wire [4-1:0] node16495;
	wire [4-1:0] node16496;
	wire [4-1:0] node16497;
	wire [4-1:0] node16498;
	wire [4-1:0] node16499;
	wire [4-1:0] node16502;
	wire [4-1:0] node16506;
	wire [4-1:0] node16507;
	wire [4-1:0] node16510;
	wire [4-1:0] node16513;
	wire [4-1:0] node16514;
	wire [4-1:0] node16516;
	wire [4-1:0] node16519;
	wire [4-1:0] node16520;
	wire [4-1:0] node16524;
	wire [4-1:0] node16525;
	wire [4-1:0] node16526;
	wire [4-1:0] node16527;
	wire [4-1:0] node16528;
	wire [4-1:0] node16529;
	wire [4-1:0] node16530;
	wire [4-1:0] node16532;
	wire [4-1:0] node16535;
	wire [4-1:0] node16538;
	wire [4-1:0] node16539;
	wire [4-1:0] node16540;
	wire [4-1:0] node16543;
	wire [4-1:0] node16546;
	wire [4-1:0] node16547;
	wire [4-1:0] node16550;
	wire [4-1:0] node16553;
	wire [4-1:0] node16554;
	wire [4-1:0] node16556;
	wire [4-1:0] node16559;
	wire [4-1:0] node16560;
	wire [4-1:0] node16562;
	wire [4-1:0] node16566;
	wire [4-1:0] node16567;
	wire [4-1:0] node16568;
	wire [4-1:0] node16569;
	wire [4-1:0] node16571;
	wire [4-1:0] node16574;
	wire [4-1:0] node16577;
	wire [4-1:0] node16578;
	wire [4-1:0] node16579;
	wire [4-1:0] node16584;
	wire [4-1:0] node16585;
	wire [4-1:0] node16587;
	wire [4-1:0] node16590;
	wire [4-1:0] node16591;
	wire [4-1:0] node16595;
	wire [4-1:0] node16596;
	wire [4-1:0] node16597;
	wire [4-1:0] node16598;
	wire [4-1:0] node16601;
	wire [4-1:0] node16602;
	wire [4-1:0] node16605;
	wire [4-1:0] node16608;
	wire [4-1:0] node16609;
	wire [4-1:0] node16610;
	wire [4-1:0] node16613;
	wire [4-1:0] node16615;
	wire [4-1:0] node16618;
	wire [4-1:0] node16619;
	wire [4-1:0] node16622;
	wire [4-1:0] node16624;
	wire [4-1:0] node16627;
	wire [4-1:0] node16628;
	wire [4-1:0] node16629;
	wire [4-1:0] node16632;
	wire [4-1:0] node16633;
	wire [4-1:0] node16637;
	wire [4-1:0] node16638;
	wire [4-1:0] node16640;
	wire [4-1:0] node16643;
	wire [4-1:0] node16646;
	wire [4-1:0] node16647;
	wire [4-1:0] node16648;
	wire [4-1:0] node16649;
	wire [4-1:0] node16650;
	wire [4-1:0] node16652;
	wire [4-1:0] node16655;
	wire [4-1:0] node16658;
	wire [4-1:0] node16659;
	wire [4-1:0] node16660;
	wire [4-1:0] node16661;
	wire [4-1:0] node16664;
	wire [4-1:0] node16668;
	wire [4-1:0] node16669;
	wire [4-1:0] node16672;
	wire [4-1:0] node16675;
	wire [4-1:0] node16676;
	wire [4-1:0] node16677;
	wire [4-1:0] node16678;
	wire [4-1:0] node16681;
	wire [4-1:0] node16684;
	wire [4-1:0] node16685;
	wire [4-1:0] node16688;
	wire [4-1:0] node16691;
	wire [4-1:0] node16692;
	wire [4-1:0] node16693;
	wire [4-1:0] node16694;
	wire [4-1:0] node16699;
	wire [4-1:0] node16700;
	wire [4-1:0] node16703;
	wire [4-1:0] node16705;
	wire [4-1:0] node16708;
	wire [4-1:0] node16709;
	wire [4-1:0] node16710;
	wire [4-1:0] node16711;
	wire [4-1:0] node16712;
	wire [4-1:0] node16716;
	wire [4-1:0] node16718;
	wire [4-1:0] node16721;
	wire [4-1:0] node16722;
	wire [4-1:0] node16725;
	wire [4-1:0] node16727;
	wire [4-1:0] node16730;
	wire [4-1:0] node16731;
	wire [4-1:0] node16732;
	wire [4-1:0] node16735;
	wire [4-1:0] node16736;
	wire [4-1:0] node16740;
	wire [4-1:0] node16741;
	wire [4-1:0] node16742;
	wire [4-1:0] node16743;
	wire [4-1:0] node16747;
	wire [4-1:0] node16748;
	wire [4-1:0] node16751;
	wire [4-1:0] node16754;
	wire [4-1:0] node16755;
	wire [4-1:0] node16756;
	wire [4-1:0] node16760;
	wire [4-1:0] node16763;
	wire [4-1:0] node16764;
	wire [4-1:0] node16765;
	wire [4-1:0] node16766;
	wire [4-1:0] node16767;
	wire [4-1:0] node16768;
	wire [4-1:0] node16769;
	wire [4-1:0] node16770;
	wire [4-1:0] node16772;
	wire [4-1:0] node16776;
	wire [4-1:0] node16777;
	wire [4-1:0] node16780;
	wire [4-1:0] node16781;
	wire [4-1:0] node16785;
	wire [4-1:0] node16786;
	wire [4-1:0] node16788;
	wire [4-1:0] node16791;
	wire [4-1:0] node16792;
	wire [4-1:0] node16796;
	wire [4-1:0] node16797;
	wire [4-1:0] node16798;
	wire [4-1:0] node16800;
	wire [4-1:0] node16803;
	wire [4-1:0] node16804;
	wire [4-1:0] node16808;
	wire [4-1:0] node16809;
	wire [4-1:0] node16811;
	wire [4-1:0] node16814;
	wire [4-1:0] node16815;
	wire [4-1:0] node16818;
	wire [4-1:0] node16821;
	wire [4-1:0] node16822;
	wire [4-1:0] node16823;
	wire [4-1:0] node16824;
	wire [4-1:0] node16825;
	wire [4-1:0] node16826;
	wire [4-1:0] node16829;
	wire [4-1:0] node16833;
	wire [4-1:0] node16835;
	wire [4-1:0] node16838;
	wire [4-1:0] node16839;
	wire [4-1:0] node16841;
	wire [4-1:0] node16843;
	wire [4-1:0] node16846;
	wire [4-1:0] node16847;
	wire [4-1:0] node16851;
	wire [4-1:0] node16852;
	wire [4-1:0] node16853;
	wire [4-1:0] node16854;
	wire [4-1:0] node16855;
	wire [4-1:0] node16860;
	wire [4-1:0] node16861;
	wire [4-1:0] node16863;
	wire [4-1:0] node16867;
	wire [4-1:0] node16868;
	wire [4-1:0] node16869;
	wire [4-1:0] node16870;
	wire [4-1:0] node16874;
	wire [4-1:0] node16877;
	wire [4-1:0] node16879;
	wire [4-1:0] node16880;
	wire [4-1:0] node16884;
	wire [4-1:0] node16885;
	wire [4-1:0] node16886;
	wire [4-1:0] node16887;
	wire [4-1:0] node16888;
	wire [4-1:0] node16892;
	wire [4-1:0] node16893;
	wire [4-1:0] node16894;
	wire [4-1:0] node16896;
	wire [4-1:0] node16899;
	wire [4-1:0] node16902;
	wire [4-1:0] node16903;
	wire [4-1:0] node16907;
	wire [4-1:0] node16908;
	wire [4-1:0] node16909;
	wire [4-1:0] node16911;
	wire [4-1:0] node16912;
	wire [4-1:0] node16916;
	wire [4-1:0] node16918;
	wire [4-1:0] node16920;
	wire [4-1:0] node16923;
	wire [4-1:0] node16925;
	wire [4-1:0] node16926;
	wire [4-1:0] node16927;
	wire [4-1:0] node16932;
	wire [4-1:0] node16933;
	wire [4-1:0] node16934;
	wire [4-1:0] node16935;
	wire [4-1:0] node16938;
	wire [4-1:0] node16940;
	wire [4-1:0] node16942;
	wire [4-1:0] node16945;
	wire [4-1:0] node16946;
	wire [4-1:0] node16947;
	wire [4-1:0] node16949;
	wire [4-1:0] node16953;
	wire [4-1:0] node16955;
	wire [4-1:0] node16957;
	wire [4-1:0] node16960;
	wire [4-1:0] node16961;
	wire [4-1:0] node16962;
	wire [4-1:0] node16963;
	wire [4-1:0] node16966;
	wire [4-1:0] node16969;
	wire [4-1:0] node16971;
	wire [4-1:0] node16974;
	wire [4-1:0] node16975;
	wire [4-1:0] node16976;
	wire [4-1:0] node16978;
	wire [4-1:0] node16981;
	wire [4-1:0] node16984;
	wire [4-1:0] node16985;
	wire [4-1:0] node16987;
	wire [4-1:0] node16990;
	wire [4-1:0] node16993;
	wire [4-1:0] node16994;
	wire [4-1:0] node16995;
	wire [4-1:0] node16996;
	wire [4-1:0] node16997;
	wire [4-1:0] node16998;
	wire [4-1:0] node16999;
	wire [4-1:0] node17002;
	wire [4-1:0] node17006;
	wire [4-1:0] node17007;
	wire [4-1:0] node17008;
	wire [4-1:0] node17011;
	wire [4-1:0] node17014;
	wire [4-1:0] node17017;
	wire [4-1:0] node17018;
	wire [4-1:0] node17020;
	wire [4-1:0] node17023;
	wire [4-1:0] node17024;
	wire [4-1:0] node17026;
	wire [4-1:0] node17030;
	wire [4-1:0] node17031;
	wire [4-1:0] node17032;
	wire [4-1:0] node17033;
	wire [4-1:0] node17034;
	wire [4-1:0] node17037;
	wire [4-1:0] node17040;
	wire [4-1:0] node17042;
	wire [4-1:0] node17045;
	wire [4-1:0] node17046;
	wire [4-1:0] node17047;
	wire [4-1:0] node17048;
	wire [4-1:0] node17051;
	wire [4-1:0] node17054;
	wire [4-1:0] node17055;
	wire [4-1:0] node17058;
	wire [4-1:0] node17061;
	wire [4-1:0] node17062;
	wire [4-1:0] node17065;
	wire [4-1:0] node17068;
	wire [4-1:0] node17069;
	wire [4-1:0] node17070;
	wire [4-1:0] node17071;
	wire [4-1:0] node17074;
	wire [4-1:0] node17077;
	wire [4-1:0] node17078;
	wire [4-1:0] node17081;
	wire [4-1:0] node17084;
	wire [4-1:0] node17086;
	wire [4-1:0] node17087;
	wire [4-1:0] node17091;
	wire [4-1:0] node17092;
	wire [4-1:0] node17093;
	wire [4-1:0] node17094;
	wire [4-1:0] node17096;
	wire [4-1:0] node17099;
	wire [4-1:0] node17102;
	wire [4-1:0] node17103;
	wire [4-1:0] node17104;
	wire [4-1:0] node17107;
	wire [4-1:0] node17110;
	wire [4-1:0] node17111;
	wire [4-1:0] node17114;
	wire [4-1:0] node17117;
	wire [4-1:0] node17118;
	wire [4-1:0] node17119;
	wire [4-1:0] node17121;
	wire [4-1:0] node17124;
	wire [4-1:0] node17127;
	wire [4-1:0] node17128;
	wire [4-1:0] node17132;
	wire [4-1:0] node17133;
	wire [4-1:0] node17134;
	wire [4-1:0] node17135;
	wire [4-1:0] node17136;
	wire [4-1:0] node17137;
	wire [4-1:0] node17138;
	wire [4-1:0] node17139;
	wire [4-1:0] node17140;
	wire [4-1:0] node17143;
	wire [4-1:0] node17145;
	wire [4-1:0] node17148;
	wire [4-1:0] node17150;
	wire [4-1:0] node17152;
	wire [4-1:0] node17155;
	wire [4-1:0] node17156;
	wire [4-1:0] node17157;
	wire [4-1:0] node17160;
	wire [4-1:0] node17162;
	wire [4-1:0] node17165;
	wire [4-1:0] node17167;
	wire [4-1:0] node17170;
	wire [4-1:0] node17171;
	wire [4-1:0] node17172;
	wire [4-1:0] node17173;
	wire [4-1:0] node17176;
	wire [4-1:0] node17177;
	wire [4-1:0] node17181;
	wire [4-1:0] node17182;
	wire [4-1:0] node17184;
	wire [4-1:0] node17187;
	wire [4-1:0] node17190;
	wire [4-1:0] node17191;
	wire [4-1:0] node17192;
	wire [4-1:0] node17195;
	wire [4-1:0] node17198;
	wire [4-1:0] node17199;
	wire [4-1:0] node17202;
	wire [4-1:0] node17205;
	wire [4-1:0] node17206;
	wire [4-1:0] node17207;
	wire [4-1:0] node17209;
	wire [4-1:0] node17211;
	wire [4-1:0] node17214;
	wire [4-1:0] node17216;
	wire [4-1:0] node17219;
	wire [4-1:0] node17220;
	wire [4-1:0] node17221;
	wire [4-1:0] node17222;
	wire [4-1:0] node17223;
	wire [4-1:0] node17226;
	wire [4-1:0] node17230;
	wire [4-1:0] node17232;
	wire [4-1:0] node17233;
	wire [4-1:0] node17236;
	wire [4-1:0] node17239;
	wire [4-1:0] node17240;
	wire [4-1:0] node17242;
	wire [4-1:0] node17243;
	wire [4-1:0] node17246;
	wire [4-1:0] node17249;
	wire [4-1:0] node17252;
	wire [4-1:0] node17253;
	wire [4-1:0] node17254;
	wire [4-1:0] node17255;
	wire [4-1:0] node17256;
	wire [4-1:0] node17257;
	wire [4-1:0] node17261;
	wire [4-1:0] node17264;
	wire [4-1:0] node17266;
	wire [4-1:0] node17267;
	wire [4-1:0] node17271;
	wire [4-1:0] node17272;
	wire [4-1:0] node17273;
	wire [4-1:0] node17275;
	wire [4-1:0] node17278;
	wire [4-1:0] node17279;
	wire [4-1:0] node17283;
	wire [4-1:0] node17284;
	wire [4-1:0] node17287;
	wire [4-1:0] node17290;
	wire [4-1:0] node17291;
	wire [4-1:0] node17292;
	wire [4-1:0] node17293;
	wire [4-1:0] node17294;
	wire [4-1:0] node17297;
	wire [4-1:0] node17300;
	wire [4-1:0] node17302;
	wire [4-1:0] node17305;
	wire [4-1:0] node17306;
	wire [4-1:0] node17308;
	wire [4-1:0] node17311;
	wire [4-1:0] node17314;
	wire [4-1:0] node17315;
	wire [4-1:0] node17317;
	wire [4-1:0] node17320;
	wire [4-1:0] node17322;
	wire [4-1:0] node17325;
	wire [4-1:0] node17326;
	wire [4-1:0] node17327;
	wire [4-1:0] node17328;
	wire [4-1:0] node17329;
	wire [4-1:0] node17330;
	wire [4-1:0] node17331;
	wire [4-1:0] node17334;
	wire [4-1:0] node17337;
	wire [4-1:0] node17338;
	wire [4-1:0] node17340;
	wire [4-1:0] node17343;
	wire [4-1:0] node17346;
	wire [4-1:0] node17347;
	wire [4-1:0] node17348;
	wire [4-1:0] node17349;
	wire [4-1:0] node17353;
	wire [4-1:0] node17356;
	wire [4-1:0] node17359;
	wire [4-1:0] node17360;
	wire [4-1:0] node17361;
	wire [4-1:0] node17362;
	wire [4-1:0] node17365;
	wire [4-1:0] node17368;
	wire [4-1:0] node17369;
	wire [4-1:0] node17373;
	wire [4-1:0] node17374;
	wire [4-1:0] node17376;
	wire [4-1:0] node17377;
	wire [4-1:0] node17381;
	wire [4-1:0] node17382;
	wire [4-1:0] node17383;
	wire [4-1:0] node17386;
	wire [4-1:0] node17389;
	wire [4-1:0] node17391;
	wire [4-1:0] node17394;
	wire [4-1:0] node17395;
	wire [4-1:0] node17396;
	wire [4-1:0] node17397;
	wire [4-1:0] node17400;
	wire [4-1:0] node17401;
	wire [4-1:0] node17405;
	wire [4-1:0] node17406;
	wire [4-1:0] node17408;
	wire [4-1:0] node17412;
	wire [4-1:0] node17413;
	wire [4-1:0] node17415;
	wire [4-1:0] node17417;
	wire [4-1:0] node17420;
	wire [4-1:0] node17421;
	wire [4-1:0] node17423;
	wire [4-1:0] node17427;
	wire [4-1:0] node17428;
	wire [4-1:0] node17429;
	wire [4-1:0] node17430;
	wire [4-1:0] node17431;
	wire [4-1:0] node17432;
	wire [4-1:0] node17436;
	wire [4-1:0] node17437;
	wire [4-1:0] node17439;
	wire [4-1:0] node17442;
	wire [4-1:0] node17445;
	wire [4-1:0] node17446;
	wire [4-1:0] node17448;
	wire [4-1:0] node17451;
	wire [4-1:0] node17453;
	wire [4-1:0] node17454;
	wire [4-1:0] node17458;
	wire [4-1:0] node17459;
	wire [4-1:0] node17460;
	wire [4-1:0] node17461;
	wire [4-1:0] node17464;
	wire [4-1:0] node17468;
	wire [4-1:0] node17469;
	wire [4-1:0] node17470;
	wire [4-1:0] node17471;
	wire [4-1:0] node17476;
	wire [4-1:0] node17477;
	wire [4-1:0] node17479;
	wire [4-1:0] node17483;
	wire [4-1:0] node17484;
	wire [4-1:0] node17485;
	wire [4-1:0] node17486;
	wire [4-1:0] node17487;
	wire [4-1:0] node17491;
	wire [4-1:0] node17492;
	wire [4-1:0] node17496;
	wire [4-1:0] node17497;
	wire [4-1:0] node17501;
	wire [4-1:0] node17502;
	wire [4-1:0] node17503;
	wire [4-1:0] node17505;
	wire [4-1:0] node17510;
	wire [4-1:0] node17511;
	wire [4-1:0] node17512;
	wire [4-1:0] node17513;
	wire [4-1:0] node17514;
	wire [4-1:0] node17515;
	wire [4-1:0] node17516;
	wire [4-1:0] node17517;
	wire [4-1:0] node17520;
	wire [4-1:0] node17521;
	wire [4-1:0] node17525;
	wire [4-1:0] node17526;
	wire [4-1:0] node17529;
	wire [4-1:0] node17530;
	wire [4-1:0] node17534;
	wire [4-1:0] node17535;
	wire [4-1:0] node17536;
	wire [4-1:0] node17540;
	wire [4-1:0] node17542;
	wire [4-1:0] node17545;
	wire [4-1:0] node17546;
	wire [4-1:0] node17547;
	wire [4-1:0] node17548;
	wire [4-1:0] node17549;
	wire [4-1:0] node17553;
	wire [4-1:0] node17556;
	wire [4-1:0] node17558;
	wire [4-1:0] node17561;
	wire [4-1:0] node17562;
	wire [4-1:0] node17565;
	wire [4-1:0] node17566;
	wire [4-1:0] node17569;
	wire [4-1:0] node17572;
	wire [4-1:0] node17573;
	wire [4-1:0] node17574;
	wire [4-1:0] node17575;
	wire [4-1:0] node17576;
	wire [4-1:0] node17577;
	wire [4-1:0] node17580;
	wire [4-1:0] node17583;
	wire [4-1:0] node17584;
	wire [4-1:0] node17587;
	wire [4-1:0] node17590;
	wire [4-1:0] node17591;
	wire [4-1:0] node17594;
	wire [4-1:0] node17597;
	wire [4-1:0] node17598;
	wire [4-1:0] node17599;
	wire [4-1:0] node17603;
	wire [4-1:0] node17605;
	wire [4-1:0] node17608;
	wire [4-1:0] node17609;
	wire [4-1:0] node17610;
	wire [4-1:0] node17612;
	wire [4-1:0] node17615;
	wire [4-1:0] node17617;
	wire [4-1:0] node17620;
	wire [4-1:0] node17621;
	wire [4-1:0] node17622;
	wire [4-1:0] node17625;
	wire [4-1:0] node17628;
	wire [4-1:0] node17629;
	wire [4-1:0] node17632;
	wire [4-1:0] node17633;
	wire [4-1:0] node17637;
	wire [4-1:0] node17638;
	wire [4-1:0] node17639;
	wire [4-1:0] node17640;
	wire [4-1:0] node17641;
	wire [4-1:0] node17642;
	wire [4-1:0] node17646;
	wire [4-1:0] node17647;
	wire [4-1:0] node17650;
	wire [4-1:0] node17653;
	wire [4-1:0] node17654;
	wire [4-1:0] node17655;
	wire [4-1:0] node17656;
	wire [4-1:0] node17661;
	wire [4-1:0] node17662;
	wire [4-1:0] node17665;
	wire [4-1:0] node17668;
	wire [4-1:0] node17669;
	wire [4-1:0] node17670;
	wire [4-1:0] node17672;
	wire [4-1:0] node17675;
	wire [4-1:0] node17677;
	wire [4-1:0] node17680;
	wire [4-1:0] node17681;
	wire [4-1:0] node17682;
	wire [4-1:0] node17686;
	wire [4-1:0] node17687;
	wire [4-1:0] node17688;
	wire [4-1:0] node17691;
	wire [4-1:0] node17694;
	wire [4-1:0] node17695;
	wire [4-1:0] node17698;
	wire [4-1:0] node17701;
	wire [4-1:0] node17702;
	wire [4-1:0] node17703;
	wire [4-1:0] node17704;
	wire [4-1:0] node17706;
	wire [4-1:0] node17707;
	wire [4-1:0] node17710;
	wire [4-1:0] node17713;
	wire [4-1:0] node17714;
	wire [4-1:0] node17717;
	wire [4-1:0] node17720;
	wire [4-1:0] node17721;
	wire [4-1:0] node17722;
	wire [4-1:0] node17726;
	wire [4-1:0] node17727;
	wire [4-1:0] node17729;
	wire [4-1:0] node17732;
	wire [4-1:0] node17735;
	wire [4-1:0] node17736;
	wire [4-1:0] node17737;
	wire [4-1:0] node17739;
	wire [4-1:0] node17741;
	wire [4-1:0] node17744;
	wire [4-1:0] node17745;
	wire [4-1:0] node17748;
	wire [4-1:0] node17750;
	wire [4-1:0] node17754;
	wire [4-1:0] node17755;
	wire [4-1:0] node17756;
	wire [4-1:0] node17757;
	wire [4-1:0] node17758;
	wire [4-1:0] node17759;
	wire [4-1:0] node17760;
	wire [4-1:0] node17761;
	wire [4-1:0] node17766;
	wire [4-1:0] node17767;
	wire [4-1:0] node17768;
	wire [4-1:0] node17772;
	wire [4-1:0] node17775;
	wire [4-1:0] node17776;
	wire [4-1:0] node17777;
	wire [4-1:0] node17779;
	wire [4-1:0] node17782;
	wire [4-1:0] node17783;
	wire [4-1:0] node17787;
	wire [4-1:0] node17788;
	wire [4-1:0] node17791;
	wire [4-1:0] node17792;
	wire [4-1:0] node17796;
	wire [4-1:0] node17797;
	wire [4-1:0] node17799;
	wire [4-1:0] node17801;
	wire [4-1:0] node17803;
	wire [4-1:0] node17806;
	wire [4-1:0] node17807;
	wire [4-1:0] node17810;
	wire [4-1:0] node17811;
	wire [4-1:0] node17815;
	wire [4-1:0] node17816;
	wire [4-1:0] node17817;
	wire [4-1:0] node17818;
	wire [4-1:0] node17819;
	wire [4-1:0] node17822;
	wire [4-1:0] node17825;
	wire [4-1:0] node17826;
	wire [4-1:0] node17827;
	wire [4-1:0] node17831;
	wire [4-1:0] node17832;
	wire [4-1:0] node17836;
	wire [4-1:0] node17838;
	wire [4-1:0] node17839;
	wire [4-1:0] node17843;
	wire [4-1:0] node17844;
	wire [4-1:0] node17845;
	wire [4-1:0] node17848;
	wire [4-1:0] node17852;
	wire [4-1:0] node17853;
	wire [4-1:0] node17854;
	wire [4-1:0] node17855;
	wire [4-1:0] node17857;
	wire [4-1:0] node17858;
	wire [4-1:0] node17859;
	wire [4-1:0] node17863;
	wire [4-1:0] node17864;
	wire [4-1:0] node17868;
	wire [4-1:0] node17869;
	wire [4-1:0] node17870;
	wire [4-1:0] node17874;
	wire [4-1:0] node17876;
	wire [4-1:0] node17877;
	wire [4-1:0] node17881;
	wire [4-1:0] node17882;
	wire [4-1:0] node17883;
	wire [4-1:0] node17884;
	wire [4-1:0] node17888;
	wire [4-1:0] node17890;
	wire [4-1:0] node17892;
	wire [4-1:0] node17896;
	wire [4-1:0] node17897;
	wire [4-1:0] node17898;
	wire [4-1:0] node17899;
	wire [4-1:0] node17901;
	wire [4-1:0] node17904;
	wire [4-1:0] node17905;
	wire [4-1:0] node17908;
	wire [4-1:0] node17910;
	wire [4-1:0] node17915;
	wire [4-1:0] node17917;
	wire [4-1:0] node17918;
	wire [4-1:0] node17919;
	wire [4-1:0] node17921;
	wire [4-1:0] node17922;
	wire [4-1:0] node17923;
	wire [4-1:0] node17924;
	wire [4-1:0] node17925;
	wire [4-1:0] node17927;
	wire [4-1:0] node17930;
	wire [4-1:0] node17931;
	wire [4-1:0] node17932;
	wire [4-1:0] node17936;
	wire [4-1:0] node17937;
	wire [4-1:0] node17941;
	wire [4-1:0] node17942;
	wire [4-1:0] node17944;
	wire [4-1:0] node17947;
	wire [4-1:0] node17948;
	wire [4-1:0] node17950;
	wire [4-1:0] node17954;
	wire [4-1:0] node17955;
	wire [4-1:0] node17956;
	wire [4-1:0] node17957;
	wire [4-1:0] node17958;
	wire [4-1:0] node17963;
	wire [4-1:0] node17964;
	wire [4-1:0] node17965;
	wire [4-1:0] node17968;
	wire [4-1:0] node17971;
	wire [4-1:0] node17972;
	wire [4-1:0] node17976;
	wire [4-1:0] node17977;
	wire [4-1:0] node17979;
	wire [4-1:0] node17982;
	wire [4-1:0] node17984;
	wire [4-1:0] node17987;
	wire [4-1:0] node17989;
	wire [4-1:0] node17990;
	wire [4-1:0] node17991;
	wire [4-1:0] node17993;
	wire [4-1:0] node17994;
	wire [4-1:0] node17995;
	wire [4-1:0] node18000;
	wire [4-1:0] node18001;
	wire [4-1:0] node18003;
	wire [4-1:0] node18004;
	wire [4-1:0] node18008;
	wire [4-1:0] node18011;
	wire [4-1:0] node18012;
	wire [4-1:0] node18013;
	wire [4-1:0] node18015;
	wire [4-1:0] node18018;
	wire [4-1:0] node18019;
	wire [4-1:0] node18020;
	wire [4-1:0] node18025;
	wire [4-1:0] node18026;
	wire [4-1:0] node18027;
	wire [4-1:0] node18031;
	wire [4-1:0] node18035;
	wire [4-1:0] node18036;
	wire [4-1:0] node18037;
	wire [4-1:0] node18038;
	wire [4-1:0] node18039;
	wire [4-1:0] node18040;
	wire [4-1:0] node18041;
	wire [4-1:0] node18042;
	wire [4-1:0] node18043;
	wire [4-1:0] node18047;
	wire [4-1:0] node18049;
	wire [4-1:0] node18052;
	wire [4-1:0] node18054;
	wire [4-1:0] node18057;
	wire [4-1:0] node18058;
	wire [4-1:0] node18059;
	wire [4-1:0] node18060;
	wire [4-1:0] node18063;
	wire [4-1:0] node18064;
	wire [4-1:0] node18068;
	wire [4-1:0] node18069;
	wire [4-1:0] node18070;
	wire [4-1:0] node18073;
	wire [4-1:0] node18076;
	wire [4-1:0] node18077;
	wire [4-1:0] node18080;
	wire [4-1:0] node18083;
	wire [4-1:0] node18085;
	wire [4-1:0] node18086;
	wire [4-1:0] node18089;
	wire [4-1:0] node18092;
	wire [4-1:0] node18093;
	wire [4-1:0] node18094;
	wire [4-1:0] node18095;
	wire [4-1:0] node18096;
	wire [4-1:0] node18098;
	wire [4-1:0] node18101;
	wire [4-1:0] node18102;
	wire [4-1:0] node18106;
	wire [4-1:0] node18107;
	wire [4-1:0] node18111;
	wire [4-1:0] node18112;
	wire [4-1:0] node18115;
	wire [4-1:0] node18116;
	wire [4-1:0] node18120;
	wire [4-1:0] node18121;
	wire [4-1:0] node18122;
	wire [4-1:0] node18125;
	wire [4-1:0] node18126;
	wire [4-1:0] node18130;
	wire [4-1:0] node18131;
	wire [4-1:0] node18132;
	wire [4-1:0] node18135;
	wire [4-1:0] node18138;
	wire [4-1:0] node18139;
	wire [4-1:0] node18142;
	wire [4-1:0] node18145;
	wire [4-1:0] node18146;
	wire [4-1:0] node18147;
	wire [4-1:0] node18148;
	wire [4-1:0] node18149;
	wire [4-1:0] node18150;
	wire [4-1:0] node18152;
	wire [4-1:0] node18155;
	wire [4-1:0] node18158;
	wire [4-1:0] node18159;
	wire [4-1:0] node18161;
	wire [4-1:0] node18165;
	wire [4-1:0] node18166;
	wire [4-1:0] node18167;
	wire [4-1:0] node18169;
	wire [4-1:0] node18172;
	wire [4-1:0] node18175;
	wire [4-1:0] node18178;
	wire [4-1:0] node18179;
	wire [4-1:0] node18180;
	wire [4-1:0] node18182;
	wire [4-1:0] node18185;
	wire [4-1:0] node18186;
	wire [4-1:0] node18190;
	wire [4-1:0] node18191;
	wire [4-1:0] node18192;
	wire [4-1:0] node18194;
	wire [4-1:0] node18197;
	wire [4-1:0] node18200;
	wire [4-1:0] node18201;
	wire [4-1:0] node18202;
	wire [4-1:0] node18205;
	wire [4-1:0] node18208;
	wire [4-1:0] node18210;
	wire [4-1:0] node18213;
	wire [4-1:0] node18214;
	wire [4-1:0] node18215;
	wire [4-1:0] node18216;
	wire [4-1:0] node18217;
	wire [4-1:0] node18220;
	wire [4-1:0] node18223;
	wire [4-1:0] node18224;
	wire [4-1:0] node18227;
	wire [4-1:0] node18230;
	wire [4-1:0] node18231;
	wire [4-1:0] node18233;
	wire [4-1:0] node18237;
	wire [4-1:0] node18238;
	wire [4-1:0] node18239;
	wire [4-1:0] node18242;
	wire [4-1:0] node18245;
	wire [4-1:0] node18246;
	wire [4-1:0] node18250;
	wire [4-1:0] node18251;
	wire [4-1:0] node18252;
	wire [4-1:0] node18253;
	wire [4-1:0] node18254;
	wire [4-1:0] node18255;
	wire [4-1:0] node18256;
	wire [4-1:0] node18257;
	wire [4-1:0] node18262;
	wire [4-1:0] node18263;
	wire [4-1:0] node18266;
	wire [4-1:0] node18268;
	wire [4-1:0] node18271;
	wire [4-1:0] node18272;
	wire [4-1:0] node18274;
	wire [4-1:0] node18277;
	wire [4-1:0] node18279;
	wire [4-1:0] node18282;
	wire [4-1:0] node18283;
	wire [4-1:0] node18284;
	wire [4-1:0] node18285;
	wire [4-1:0] node18288;
	wire [4-1:0] node18291;
	wire [4-1:0] node18292;
	wire [4-1:0] node18293;
	wire [4-1:0] node18297;
	wire [4-1:0] node18299;
	wire [4-1:0] node18302;
	wire [4-1:0] node18303;
	wire [4-1:0] node18304;
	wire [4-1:0] node18308;
	wire [4-1:0] node18309;
	wire [4-1:0] node18310;
	wire [4-1:0] node18313;
	wire [4-1:0] node18316;
	wire [4-1:0] node18318;
	wire [4-1:0] node18321;
	wire [4-1:0] node18322;
	wire [4-1:0] node18323;
	wire [4-1:0] node18324;
	wire [4-1:0] node18325;
	wire [4-1:0] node18328;
	wire [4-1:0] node18331;
	wire [4-1:0] node18332;
	wire [4-1:0] node18335;
	wire [4-1:0] node18338;
	wire [4-1:0] node18339;
	wire [4-1:0] node18341;
	wire [4-1:0] node18344;
	wire [4-1:0] node18345;
	wire [4-1:0] node18349;
	wire [4-1:0] node18350;
	wire [4-1:0] node18351;
	wire [4-1:0] node18352;
	wire [4-1:0] node18357;
	wire [4-1:0] node18358;
	wire [4-1:0] node18359;
	wire [4-1:0] node18364;
	wire [4-1:0] node18365;
	wire [4-1:0] node18366;
	wire [4-1:0] node18367;
	wire [4-1:0] node18368;
	wire [4-1:0] node18370;
	wire [4-1:0] node18371;
	wire [4-1:0] node18375;
	wire [4-1:0] node18376;
	wire [4-1:0] node18377;
	wire [4-1:0] node18381;
	wire [4-1:0] node18384;
	wire [4-1:0] node18385;
	wire [4-1:0] node18387;
	wire [4-1:0] node18390;
	wire [4-1:0] node18392;
	wire [4-1:0] node18395;
	wire [4-1:0] node18396;
	wire [4-1:0] node18397;
	wire [4-1:0] node18398;
	wire [4-1:0] node18399;
	wire [4-1:0] node18403;
	wire [4-1:0] node18407;
	wire [4-1:0] node18408;
	wire [4-1:0] node18409;
	wire [4-1:0] node18414;
	wire [4-1:0] node18415;
	wire [4-1:0] node18416;
	wire [4-1:0] node18417;
	wire [4-1:0] node18418;
	wire [4-1:0] node18419;
	wire [4-1:0] node18424;
	wire [4-1:0] node18425;
	wire [4-1:0] node18426;
	wire [4-1:0] node18431;
	wire [4-1:0] node18432;
	wire [4-1:0] node18433;
	wire [4-1:0] node18435;
	wire [4-1:0] node18440;
	wire [4-1:0] node18441;
	wire [4-1:0] node18442;
	wire [4-1:0] node18447;
	wire [4-1:0] node18449;
	wire [4-1:0] node18450;
	wire [4-1:0] node18451;
	wire [4-1:0] node18452;
	wire [4-1:0] node18453;
	wire [4-1:0] node18454;
	wire [4-1:0] node18458;
	wire [4-1:0] node18459;
	wire [4-1:0] node18460;
	wire [4-1:0] node18462;
	wire [4-1:0] node18465;
	wire [4-1:0] node18467;
	wire [4-1:0] node18470;
	wire [4-1:0] node18472;
	wire [4-1:0] node18475;
	wire [4-1:0] node18476;
	wire [4-1:0] node18477;
	wire [4-1:0] node18478;
	wire [4-1:0] node18482;
	wire [4-1:0] node18483;
	wire [4-1:0] node18484;
	wire [4-1:0] node18489;
	wire [4-1:0] node18490;
	wire [4-1:0] node18491;
	wire [4-1:0] node18495;
	wire [4-1:0] node18496;
	wire [4-1:0] node18497;
	wire [4-1:0] node18501;
	wire [4-1:0] node18502;
	wire [4-1:0] node18507;
	wire [4-1:0] node18508;
	wire [4-1:0] node18509;
	wire [4-1:0] node18510;
	wire [4-1:0] node18511;
	wire [4-1:0] node18512;
	wire [4-1:0] node18515;
	wire [4-1:0] node18516;
	wire [4-1:0] node18521;
	wire [4-1:0] node18522;
	wire [4-1:0] node18523;
	wire [4-1:0] node18527;
	wire [4-1:0] node18528;
	wire [4-1:0] node18532;
	wire [4-1:0] node18533;
	wire [4-1:0] node18534;
	wire [4-1:0] node18536;
	wire [4-1:0] node18537;
	wire [4-1:0] node18541;
	wire [4-1:0] node18542;
	wire [4-1:0] node18543;
	wire [4-1:0] node18546;
	wire [4-1:0] node18549;
	wire [4-1:0] node18550;
	wire [4-1:0] node18554;
	wire [4-1:0] node18555;
	wire [4-1:0] node18556;
	wire [4-1:0] node18561;
	wire [4-1:0] node18562;
	wire [4-1:0] node18563;
	wire [4-1:0] node18564;
	wire [4-1:0] node18565;
	wire [4-1:0] node18566;
	wire [4-1:0] node18572;
	wire [4-1:0] node18573;
	wire [4-1:0] node18574;
	wire [4-1:0] node18575;
	wire [4-1:0] node18578;
	wire [4-1:0] node18582;
	wire [4-1:0] node18584;
	wire [4-1:0] node18585;
	wire [4-1:0] node18589;
	wire [4-1:0] node18591;
	wire [4-1:0] node18592;
	wire [4-1:0] node18593;
	wire [4-1:0] node18598;
	wire [4-1:0] node18599;
	wire [4-1:0] node18600;
	wire [4-1:0] node18601;
	wire [4-1:0] node18602;
	wire [4-1:0] node18603;
	wire [4-1:0] node18604;
	wire [4-1:0] node18605;
	wire [4-1:0] node18606;
	wire [4-1:0] node18608;
	wire [4-1:0] node18609;
	wire [4-1:0] node18610;
	wire [4-1:0] node18612;
	wire [4-1:0] node18614;
	wire [4-1:0] node18617;
	wire [4-1:0] node18618;
	wire [4-1:0] node18619;
	wire [4-1:0] node18624;
	wire [4-1:0] node18626;
	wire [4-1:0] node18628;
	wire [4-1:0] node18632;
	wire [4-1:0] node18633;
	wire [4-1:0] node18634;
	wire [4-1:0] node18635;
	wire [4-1:0] node18636;
	wire [4-1:0] node18638;
	wire [4-1:0] node18641;
	wire [4-1:0] node18642;
	wire [4-1:0] node18646;
	wire [4-1:0] node18647;
	wire [4-1:0] node18648;
	wire [4-1:0] node18651;
	wire [4-1:0] node18653;
	wire [4-1:0] node18656;
	wire [4-1:0] node18657;
	wire [4-1:0] node18661;
	wire [4-1:0] node18662;
	wire [4-1:0] node18663;
	wire [4-1:0] node18664;
	wire [4-1:0] node18666;
	wire [4-1:0] node18670;
	wire [4-1:0] node18671;
	wire [4-1:0] node18672;
	wire [4-1:0] node18676;
	wire [4-1:0] node18679;
	wire [4-1:0] node18680;
	wire [4-1:0] node18682;
	wire [4-1:0] node18685;
	wire [4-1:0] node18688;
	wire [4-1:0] node18690;
	wire [4-1:0] node18691;
	wire [4-1:0] node18692;
	wire [4-1:0] node18695;
	wire [4-1:0] node18696;
	wire [4-1:0] node18698;
	wire [4-1:0] node18702;
	wire [4-1:0] node18703;
	wire [4-1:0] node18705;
	wire [4-1:0] node18709;
	wire [4-1:0] node18710;
	wire [4-1:0] node18711;
	wire [4-1:0] node18712;
	wire [4-1:0] node18713;
	wire [4-1:0] node18714;
	wire [4-1:0] node18716;
	wire [4-1:0] node18719;
	wire [4-1:0] node18720;
	wire [4-1:0] node18724;
	wire [4-1:0] node18725;
	wire [4-1:0] node18727;
	wire [4-1:0] node18730;
	wire [4-1:0] node18731;
	wire [4-1:0] node18735;
	wire [4-1:0] node18736;
	wire [4-1:0] node18738;
	wire [4-1:0] node18741;
	wire [4-1:0] node18742;
	wire [4-1:0] node18744;
	wire [4-1:0] node18748;
	wire [4-1:0] node18749;
	wire [4-1:0] node18750;
	wire [4-1:0] node18751;
	wire [4-1:0] node18752;
	wire [4-1:0] node18756;
	wire [4-1:0] node18757;
	wire [4-1:0] node18761;
	wire [4-1:0] node18762;
	wire [4-1:0] node18763;
	wire [4-1:0] node18766;
	wire [4-1:0] node18767;
	wire [4-1:0] node18772;
	wire [4-1:0] node18773;
	wire [4-1:0] node18774;
	wire [4-1:0] node18777;
	wire [4-1:0] node18779;
	wire [4-1:0] node18780;
	wire [4-1:0] node18784;
	wire [4-1:0] node18785;
	wire [4-1:0] node18787;
	wire [4-1:0] node18788;
	wire [4-1:0] node18791;
	wire [4-1:0] node18794;
	wire [4-1:0] node18795;
	wire [4-1:0] node18799;
	wire [4-1:0] node18800;
	wire [4-1:0] node18801;
	wire [4-1:0] node18802;
	wire [4-1:0] node18803;
	wire [4-1:0] node18804;
	wire [4-1:0] node18805;
	wire [4-1:0] node18811;
	wire [4-1:0] node18812;
	wire [4-1:0] node18813;
	wire [4-1:0] node18817;
	wire [4-1:0] node18819;
	wire [4-1:0] node18821;
	wire [4-1:0] node18824;
	wire [4-1:0] node18825;
	wire [4-1:0] node18826;
	wire [4-1:0] node18828;
	wire [4-1:0] node18831;
	wire [4-1:0] node18832;
	wire [4-1:0] node18836;
	wire [4-1:0] node18837;
	wire [4-1:0] node18839;
	wire [4-1:0] node18840;
	wire [4-1:0] node18843;
	wire [4-1:0] node18846;
	wire [4-1:0] node18848;
	wire [4-1:0] node18849;
	wire [4-1:0] node18853;
	wire [4-1:0] node18854;
	wire [4-1:0] node18855;
	wire [4-1:0] node18856;
	wire [4-1:0] node18857;
	wire [4-1:0] node18861;
	wire [4-1:0] node18864;
	wire [4-1:0] node18865;
	wire [4-1:0] node18866;
	wire [4-1:0] node18870;
	wire [4-1:0] node18872;
	wire [4-1:0] node18873;
	wire [4-1:0] node18877;
	wire [4-1:0] node18878;
	wire [4-1:0] node18880;
	wire [4-1:0] node18883;
	wire [4-1:0] node18884;
	wire [4-1:0] node18885;
	wire [4-1:0] node18889;
	wire [4-1:0] node18891;
	wire [4-1:0] node18894;
	wire [4-1:0] node18895;
	wire [4-1:0] node18896;
	wire [4-1:0] node18897;
	wire [4-1:0] node18898;
	wire [4-1:0] node18899;
	wire [4-1:0] node18900;
	wire [4-1:0] node18904;
	wire [4-1:0] node18905;
	wire [4-1:0] node18907;
	wire [4-1:0] node18911;
	wire [4-1:0] node18912;
	wire [4-1:0] node18913;
	wire [4-1:0] node18917;
	wire [4-1:0] node18919;
	wire [4-1:0] node18920;
	wire [4-1:0] node18924;
	wire [4-1:0] node18925;
	wire [4-1:0] node18926;
	wire [4-1:0] node18930;
	wire [4-1:0] node18931;
	wire [4-1:0] node18933;
	wire [4-1:0] node18937;
	wire [4-1:0] node18938;
	wire [4-1:0] node18939;
	wire [4-1:0] node18941;
	wire [4-1:0] node18944;
	wire [4-1:0] node18945;
	wire [4-1:0] node18947;
	wire [4-1:0] node18950;
	wire [4-1:0] node18952;
	wire [4-1:0] node18955;
	wire [4-1:0] node18956;
	wire [4-1:0] node18957;
	wire [4-1:0] node18958;
	wire [4-1:0] node18962;
	wire [4-1:0] node18964;
	wire [4-1:0] node18966;
	wire [4-1:0] node18969;
	wire [4-1:0] node18970;
	wire [4-1:0] node18972;
	wire [4-1:0] node18975;
	wire [4-1:0] node18976;
	wire [4-1:0] node18977;
	wire [4-1:0] node18981;
	wire [4-1:0] node18982;
	wire [4-1:0] node18986;
	wire [4-1:0] node18987;
	wire [4-1:0] node18988;
	wire [4-1:0] node18989;
	wire [4-1:0] node18990;
	wire [4-1:0] node18991;
	wire [4-1:0] node18995;
	wire [4-1:0] node18997;
	wire [4-1:0] node19000;
	wire [4-1:0] node19001;
	wire [4-1:0] node19002;
	wire [4-1:0] node19004;
	wire [4-1:0] node19007;
	wire [4-1:0] node19008;
	wire [4-1:0] node19012;
	wire [4-1:0] node19013;
	wire [4-1:0] node19014;
	wire [4-1:0] node19018;
	wire [4-1:0] node19021;
	wire [4-1:0] node19022;
	wire [4-1:0] node19023;
	wire [4-1:0] node19024;
	wire [4-1:0] node19028;
	wire [4-1:0] node19029;
	wire [4-1:0] node19031;
	wire [4-1:0] node19034;
	wire [4-1:0] node19036;
	wire [4-1:0] node19039;
	wire [4-1:0] node19040;
	wire [4-1:0] node19042;
	wire [4-1:0] node19045;
	wire [4-1:0] node19047;
	wire [4-1:0] node19050;
	wire [4-1:0] node19051;
	wire [4-1:0] node19052;
	wire [4-1:0] node19053;
	wire [4-1:0] node19054;
	wire [4-1:0] node19058;
	wire [4-1:0] node19059;
	wire [4-1:0] node19063;
	wire [4-1:0] node19064;
	wire [4-1:0] node19066;
	wire [4-1:0] node19069;
	wire [4-1:0] node19070;
	wire [4-1:0] node19072;
	wire [4-1:0] node19075;
	wire [4-1:0] node19077;
	wire [4-1:0] node19080;
	wire [4-1:0] node19081;
	wire [4-1:0] node19082;
	wire [4-1:0] node19083;
	wire [4-1:0] node19085;
	wire [4-1:0] node19089;
	wire [4-1:0] node19090;
	wire [4-1:0] node19093;
	wire [4-1:0] node19096;
	wire [4-1:0] node19097;
	wire [4-1:0] node19099;
	wire [4-1:0] node19102;
	wire [4-1:0] node19103;
	wire [4-1:0] node19104;
	wire [4-1:0] node19109;
	wire [4-1:0] node19111;
	wire [4-1:0] node19112;
	wire [4-1:0] node19113;
	wire [4-1:0] node19114;
	wire [4-1:0] node19116;
	wire [4-1:0] node19117;
	wire [4-1:0] node19119;
	wire [4-1:0] node19122;
	wire [4-1:0] node19124;
	wire [4-1:0] node19125;
	wire [4-1:0] node19129;
	wire [4-1:0] node19130;
	wire [4-1:0] node19131;
	wire [4-1:0] node19132;
	wire [4-1:0] node19133;
	wire [4-1:0] node19137;
	wire [4-1:0] node19138;
	wire [4-1:0] node19142;
	wire [4-1:0] node19143;
	wire [4-1:0] node19144;
	wire [4-1:0] node19145;
	wire [4-1:0] node19151;
	wire [4-1:0] node19152;
	wire [4-1:0] node19153;
	wire [4-1:0] node19155;
	wire [4-1:0] node19158;
	wire [4-1:0] node19159;
	wire [4-1:0] node19161;
	wire [4-1:0] node19165;
	wire [4-1:0] node19166;
	wire [4-1:0] node19167;
	wire [4-1:0] node19169;
	wire [4-1:0] node19173;
	wire [4-1:0] node19174;
	wire [4-1:0] node19177;
	wire [4-1:0] node19180;
	wire [4-1:0] node19182;
	wire [4-1:0] node19184;
	wire [4-1:0] node19185;
	wire [4-1:0] node19187;
	wire [4-1:0] node19190;
	wire [4-1:0] node19191;
	wire [4-1:0] node19192;
	wire [4-1:0] node19194;
	wire [4-1:0] node19199;
	wire [4-1:0] node19200;
	wire [4-1:0] node19201;
	wire [4-1:0] node19202;
	wire [4-1:0] node19203;
	wire [4-1:0] node19204;
	wire [4-1:0] node19205;
	wire [4-1:0] node19209;
	wire [4-1:0] node19210;
	wire [4-1:0] node19214;
	wire [4-1:0] node19215;
	wire [4-1:0] node19216;
	wire [4-1:0] node19219;
	wire [4-1:0] node19222;
	wire [4-1:0] node19224;
	wire [4-1:0] node19225;
	wire [4-1:0] node19228;
	wire [4-1:0] node19231;
	wire [4-1:0] node19232;
	wire [4-1:0] node19233;
	wire [4-1:0] node19235;
	wire [4-1:0] node19239;
	wire [4-1:0] node19240;
	wire [4-1:0] node19242;
	wire [4-1:0] node19246;
	wire [4-1:0] node19247;
	wire [4-1:0] node19248;
	wire [4-1:0] node19249;
	wire [4-1:0] node19252;
	wire [4-1:0] node19254;
	wire [4-1:0] node19257;
	wire [4-1:0] node19258;
	wire [4-1:0] node19262;
	wire [4-1:0] node19263;
	wire [4-1:0] node19264;
	wire [4-1:0] node19265;
	wire [4-1:0] node19269;
	wire [4-1:0] node19271;
	wire [4-1:0] node19274;
	wire [4-1:0] node19275;
	wire [4-1:0] node19277;
	wire [4-1:0] node19281;
	wire [4-1:0] node19282;
	wire [4-1:0] node19283;
	wire [4-1:0] node19284;
	wire [4-1:0] node19285;
	wire [4-1:0] node19286;
	wire [4-1:0] node19290;
	wire [4-1:0] node19291;
	wire [4-1:0] node19295;
	wire [4-1:0] node19296;
	wire [4-1:0] node19299;
	wire [4-1:0] node19300;
	wire [4-1:0] node19303;
	wire [4-1:0] node19304;
	wire [4-1:0] node19307;
	wire [4-1:0] node19310;
	wire [4-1:0] node19311;
	wire [4-1:0] node19312;
	wire [4-1:0] node19316;
	wire [4-1:0] node19317;
	wire [4-1:0] node19319;
	wire [4-1:0] node19323;
	wire [4-1:0] node19324;
	wire [4-1:0] node19325;
	wire [4-1:0] node19326;
	wire [4-1:0] node19327;
	wire [4-1:0] node19331;
	wire [4-1:0] node19332;
	wire [4-1:0] node19336;
	wire [4-1:0] node19337;
	wire [4-1:0] node19339;
	wire [4-1:0] node19340;
	wire [4-1:0] node19344;
	wire [4-1:0] node19346;
	wire [4-1:0] node19348;
	wire [4-1:0] node19351;
	wire [4-1:0] node19352;
	wire [4-1:0] node19354;
	wire [4-1:0] node19355;
	wire [4-1:0] node19356;
	wire [4-1:0] node19361;
	wire [4-1:0] node19362;
	wire [4-1:0] node19364;
	wire [4-1:0] node19367;
	wire [4-1:0] node19368;
	wire [4-1:0] node19369;
	wire [4-1:0] node19375;
	wire [4-1:0] node19376;
	wire [4-1:0] node19377;
	wire [4-1:0] node19378;
	wire [4-1:0] node19379;
	wire [4-1:0] node19380;
	wire [4-1:0] node19381;
	wire [4-1:0] node19382;
	wire [4-1:0] node19383;
	wire [4-1:0] node19384;
	wire [4-1:0] node19387;
	wire [4-1:0] node19390;
	wire [4-1:0] node19391;
	wire [4-1:0] node19392;
	wire [4-1:0] node19395;
	wire [4-1:0] node19398;
	wire [4-1:0] node19399;
	wire [4-1:0] node19403;
	wire [4-1:0] node19404;
	wire [4-1:0] node19406;
	wire [4-1:0] node19409;
	wire [4-1:0] node19412;
	wire [4-1:0] node19413;
	wire [4-1:0] node19414;
	wire [4-1:0] node19415;
	wire [4-1:0] node19416;
	wire [4-1:0] node19419;
	wire [4-1:0] node19420;
	wire [4-1:0] node19424;
	wire [4-1:0] node19425;
	wire [4-1:0] node19427;
	wire [4-1:0] node19431;
	wire [4-1:0] node19432;
	wire [4-1:0] node19434;
	wire [4-1:0] node19437;
	wire [4-1:0] node19438;
	wire [4-1:0] node19441;
	wire [4-1:0] node19444;
	wire [4-1:0] node19445;
	wire [4-1:0] node19446;
	wire [4-1:0] node19449;
	wire [4-1:0] node19450;
	wire [4-1:0] node19454;
	wire [4-1:0] node19455;
	wire [4-1:0] node19456;
	wire [4-1:0] node19458;
	wire [4-1:0] node19462;
	wire [4-1:0] node19463;
	wire [4-1:0] node19466;
	wire [4-1:0] node19467;
	wire [4-1:0] node19471;
	wire [4-1:0] node19472;
	wire [4-1:0] node19473;
	wire [4-1:0] node19474;
	wire [4-1:0] node19475;
	wire [4-1:0] node19476;
	wire [4-1:0] node19480;
	wire [4-1:0] node19482;
	wire [4-1:0] node19485;
	wire [4-1:0] node19486;
	wire [4-1:0] node19488;
	wire [4-1:0] node19492;
	wire [4-1:0] node19493;
	wire [4-1:0] node19495;
	wire [4-1:0] node19498;
	wire [4-1:0] node19499;
	wire [4-1:0] node19501;
	wire [4-1:0] node19505;
	wire [4-1:0] node19506;
	wire [4-1:0] node19507;
	wire [4-1:0] node19508;
	wire [4-1:0] node19511;
	wire [4-1:0] node19513;
	wire [4-1:0] node19516;
	wire [4-1:0] node19517;
	wire [4-1:0] node19518;
	wire [4-1:0] node19523;
	wire [4-1:0] node19524;
	wire [4-1:0] node19525;
	wire [4-1:0] node19527;
	wire [4-1:0] node19531;
	wire [4-1:0] node19532;
	wire [4-1:0] node19533;
	wire [4-1:0] node19535;
	wire [4-1:0] node19538;
	wire [4-1:0] node19541;
	wire [4-1:0] node19542;
	wire [4-1:0] node19545;
	wire [4-1:0] node19547;
	wire [4-1:0] node19550;
	wire [4-1:0] node19551;
	wire [4-1:0] node19552;
	wire [4-1:0] node19553;
	wire [4-1:0] node19554;
	wire [4-1:0] node19555;
	wire [4-1:0] node19557;
	wire [4-1:0] node19558;
	wire [4-1:0] node19562;
	wire [4-1:0] node19563;
	wire [4-1:0] node19567;
	wire [4-1:0] node19569;
	wire [4-1:0] node19570;
	wire [4-1:0] node19574;
	wire [4-1:0] node19575;
	wire [4-1:0] node19577;
	wire [4-1:0] node19578;
	wire [4-1:0] node19580;
	wire [4-1:0] node19584;
	wire [4-1:0] node19585;
	wire [4-1:0] node19586;
	wire [4-1:0] node19588;
	wire [4-1:0] node19591;
	wire [4-1:0] node19592;
	wire [4-1:0] node19596;
	wire [4-1:0] node19598;
	wire [4-1:0] node19599;
	wire [4-1:0] node19603;
	wire [4-1:0] node19604;
	wire [4-1:0] node19605;
	wire [4-1:0] node19606;
	wire [4-1:0] node19608;
	wire [4-1:0] node19612;
	wire [4-1:0] node19613;
	wire [4-1:0] node19615;
	wire [4-1:0] node19618;
	wire [4-1:0] node19619;
	wire [4-1:0] node19622;
	wire [4-1:0] node19625;
	wire [4-1:0] node19626;
	wire [4-1:0] node19627;
	wire [4-1:0] node19628;
	wire [4-1:0] node19629;
	wire [4-1:0] node19633;
	wire [4-1:0] node19634;
	wire [4-1:0] node19638;
	wire [4-1:0] node19639;
	wire [4-1:0] node19640;
	wire [4-1:0] node19643;
	wire [4-1:0] node19646;
	wire [4-1:0] node19649;
	wire [4-1:0] node19651;
	wire [4-1:0] node19652;
	wire [4-1:0] node19656;
	wire [4-1:0] node19657;
	wire [4-1:0] node19658;
	wire [4-1:0] node19659;
	wire [4-1:0] node19661;
	wire [4-1:0] node19663;
	wire [4-1:0] node19666;
	wire [4-1:0] node19667;
	wire [4-1:0] node19668;
	wire [4-1:0] node19669;
	wire [4-1:0] node19673;
	wire [4-1:0] node19677;
	wire [4-1:0] node19678;
	wire [4-1:0] node19679;
	wire [4-1:0] node19680;
	wire [4-1:0] node19681;
	wire [4-1:0] node19685;
	wire [4-1:0] node19686;
	wire [4-1:0] node19689;
	wire [4-1:0] node19692;
	wire [4-1:0] node19693;
	wire [4-1:0] node19694;
	wire [4-1:0] node19698;
	wire [4-1:0] node19700;
	wire [4-1:0] node19703;
	wire [4-1:0] node19704;
	wire [4-1:0] node19706;
	wire [4-1:0] node19709;
	wire [4-1:0] node19711;
	wire [4-1:0] node19714;
	wire [4-1:0] node19715;
	wire [4-1:0] node19716;
	wire [4-1:0] node19717;
	wire [4-1:0] node19719;
	wire [4-1:0] node19723;
	wire [4-1:0] node19724;
	wire [4-1:0] node19725;
	wire [4-1:0] node19726;
	wire [4-1:0] node19730;
	wire [4-1:0] node19733;
	wire [4-1:0] node19734;
	wire [4-1:0] node19737;
	wire [4-1:0] node19740;
	wire [4-1:0] node19741;
	wire [4-1:0] node19742;
	wire [4-1:0] node19743;
	wire [4-1:0] node19746;
	wire [4-1:0] node19747;
	wire [4-1:0] node19751;
	wire [4-1:0] node19752;
	wire [4-1:0] node19755;
	wire [4-1:0] node19758;
	wire [4-1:0] node19759;
	wire [4-1:0] node19761;
	wire [4-1:0] node19764;
	wire [4-1:0] node19765;
	wire [4-1:0] node19769;
	wire [4-1:0] node19770;
	wire [4-1:0] node19771;
	wire [4-1:0] node19772;
	wire [4-1:0] node19773;
	wire [4-1:0] node19774;
	wire [4-1:0] node19776;
	wire [4-1:0] node19777;
	wire [4-1:0] node19781;
	wire [4-1:0] node19782;
	wire [4-1:0] node19783;
	wire [4-1:0] node19787;
	wire [4-1:0] node19789;
	wire [4-1:0] node19792;
	wire [4-1:0] node19793;
	wire [4-1:0] node19794;
	wire [4-1:0] node19795;
	wire [4-1:0] node19798;
	wire [4-1:0] node19801;
	wire [4-1:0] node19802;
	wire [4-1:0] node19803;
	wire [4-1:0] node19807;
	wire [4-1:0] node19809;
	wire [4-1:0] node19812;
	wire [4-1:0] node19813;
	wire [4-1:0] node19814;
	wire [4-1:0] node19817;
	wire [4-1:0] node19820;
	wire [4-1:0] node19821;
	wire [4-1:0] node19824;
	wire [4-1:0] node19827;
	wire [4-1:0] node19828;
	wire [4-1:0] node19829;
	wire [4-1:0] node19831;
	wire [4-1:0] node19834;
	wire [4-1:0] node19836;
	wire [4-1:0] node19837;
	wire [4-1:0] node19841;
	wire [4-1:0] node19842;
	wire [4-1:0] node19843;
	wire [4-1:0] node19844;
	wire [4-1:0] node19848;
	wire [4-1:0] node19850;
	wire [4-1:0] node19853;
	wire [4-1:0] node19855;
	wire [4-1:0] node19856;
	wire [4-1:0] node19860;
	wire [4-1:0] node19861;
	wire [4-1:0] node19862;
	wire [4-1:0] node19863;
	wire [4-1:0] node19864;
	wire [4-1:0] node19866;
	wire [4-1:0] node19869;
	wire [4-1:0] node19872;
	wire [4-1:0] node19873;
	wire [4-1:0] node19874;
	wire [4-1:0] node19877;
	wire [4-1:0] node19880;
	wire [4-1:0] node19881;
	wire [4-1:0] node19884;
	wire [4-1:0] node19887;
	wire [4-1:0] node19888;
	wire [4-1:0] node19889;
	wire [4-1:0] node19890;
	wire [4-1:0] node19893;
	wire [4-1:0] node19897;
	wire [4-1:0] node19898;
	wire [4-1:0] node19900;
	wire [4-1:0] node19903;
	wire [4-1:0] node19904;
	wire [4-1:0] node19908;
	wire [4-1:0] node19909;
	wire [4-1:0] node19910;
	wire [4-1:0] node19912;
	wire [4-1:0] node19913;
	wire [4-1:0] node19917;
	wire [4-1:0] node19918;
	wire [4-1:0] node19919;
	wire [4-1:0] node19920;
	wire [4-1:0] node19924;
	wire [4-1:0] node19927;
	wire [4-1:0] node19930;
	wire [4-1:0] node19931;
	wire [4-1:0] node19932;
	wire [4-1:0] node19933;
	wire [4-1:0] node19936;
	wire [4-1:0] node19939;
	wire [4-1:0] node19940;
	wire [4-1:0] node19944;
	wire [4-1:0] node19945;
	wire [4-1:0] node19947;
	wire [4-1:0] node19950;
	wire [4-1:0] node19953;
	wire [4-1:0] node19954;
	wire [4-1:0] node19955;
	wire [4-1:0] node19956;
	wire [4-1:0] node19957;
	wire [4-1:0] node19960;
	wire [4-1:0] node19961;
	wire [4-1:0] node19962;
	wire [4-1:0] node19966;
	wire [4-1:0] node19967;
	wire [4-1:0] node19971;
	wire [4-1:0] node19972;
	wire [4-1:0] node19973;
	wire [4-1:0] node19977;
	wire [4-1:0] node19978;
	wire [4-1:0] node19980;
	wire [4-1:0] node19983;
	wire [4-1:0] node19984;
	wire [4-1:0] node19986;
	wire [4-1:0] node19989;
	wire [4-1:0] node19990;
	wire [4-1:0] node19994;
	wire [4-1:0] node19995;
	wire [4-1:0] node19996;
	wire [4-1:0] node19998;
	wire [4-1:0] node20001;
	wire [4-1:0] node20002;
	wire [4-1:0] node20003;
	wire [4-1:0] node20006;
	wire [4-1:0] node20010;
	wire [4-1:0] node20011;
	wire [4-1:0] node20012;
	wire [4-1:0] node20014;
	wire [4-1:0] node20017;
	wire [4-1:0] node20018;
	wire [4-1:0] node20022;
	wire [4-1:0] node20023;
	wire [4-1:0] node20024;
	wire [4-1:0] node20027;
	wire [4-1:0] node20030;
	wire [4-1:0] node20032;
	wire [4-1:0] node20033;
	wire [4-1:0] node20037;
	wire [4-1:0] node20038;
	wire [4-1:0] node20039;
	wire [4-1:0] node20040;
	wire [4-1:0] node20042;
	wire [4-1:0] node20045;
	wire [4-1:0] node20046;
	wire [4-1:0] node20047;
	wire [4-1:0] node20050;
	wire [4-1:0] node20053;
	wire [4-1:0] node20054;
	wire [4-1:0] node20055;
	wire [4-1:0] node20058;
	wire [4-1:0] node20062;
	wire [4-1:0] node20063;
	wire [4-1:0] node20065;
	wire [4-1:0] node20068;
	wire [4-1:0] node20069;
	wire [4-1:0] node20072;
	wire [4-1:0] node20075;
	wire [4-1:0] node20076;
	wire [4-1:0] node20078;
	wire [4-1:0] node20079;
	wire [4-1:0] node20083;
	wire [4-1:0] node20084;
	wire [4-1:0] node20088;
	wire [4-1:0] node20089;
	wire [4-1:0] node20090;
	wire [4-1:0] node20091;
	wire [4-1:0] node20093;
	wire [4-1:0] node20094;
	wire [4-1:0] node20095;
	wire [4-1:0] node20097;
	wire [4-1:0] node20099;
	wire [4-1:0] node20102;
	wire [4-1:0] node20103;
	wire [4-1:0] node20104;
	wire [4-1:0] node20105;
	wire [4-1:0] node20109;
	wire [4-1:0] node20110;
	wire [4-1:0] node20114;
	wire [4-1:0] node20118;
	wire [4-1:0] node20119;
	wire [4-1:0] node20120;
	wire [4-1:0] node20121;
	wire [4-1:0] node20122;
	wire [4-1:0] node20124;
	wire [4-1:0] node20127;
	wire [4-1:0] node20128;
	wire [4-1:0] node20131;
	wire [4-1:0] node20134;
	wire [4-1:0] node20135;
	wire [4-1:0] node20136;
	wire [4-1:0] node20140;
	wire [4-1:0] node20142;
	wire [4-1:0] node20145;
	wire [4-1:0] node20146;
	wire [4-1:0] node20147;
	wire [4-1:0] node20148;
	wire [4-1:0] node20149;
	wire [4-1:0] node20152;
	wire [4-1:0] node20156;
	wire [4-1:0] node20157;
	wire [4-1:0] node20159;
	wire [4-1:0] node20162;
	wire [4-1:0] node20165;
	wire [4-1:0] node20166;
	wire [4-1:0] node20168;
	wire [4-1:0] node20171;
	wire [4-1:0] node20173;
	wire [4-1:0] node20176;
	wire [4-1:0] node20178;
	wire [4-1:0] node20179;
	wire [4-1:0] node20180;
	wire [4-1:0] node20182;
	wire [4-1:0] node20183;
	wire [4-1:0] node20187;
	wire [4-1:0] node20188;
	wire [4-1:0] node20191;
	wire [4-1:0] node20193;
	wire [4-1:0] node20196;
	wire [4-1:0] node20198;
	wire [4-1:0] node20200;
	wire [4-1:0] node20203;
	wire [4-1:0] node20204;
	wire [4-1:0] node20205;
	wire [4-1:0] node20206;
	wire [4-1:0] node20207;
	wire [4-1:0] node20208;
	wire [4-1:0] node20210;
	wire [4-1:0] node20213;
	wire [4-1:0] node20214;
	wire [4-1:0] node20218;
	wire [4-1:0] node20219;
	wire [4-1:0] node20220;
	wire [4-1:0] node20224;
	wire [4-1:0] node20225;
	wire [4-1:0] node20227;
	wire [4-1:0] node20230;
	wire [4-1:0] node20231;
	wire [4-1:0] node20235;
	wire [4-1:0] node20236;
	wire [4-1:0] node20237;
	wire [4-1:0] node20239;
	wire [4-1:0] node20242;
	wire [4-1:0] node20243;
	wire [4-1:0] node20244;
	wire [4-1:0] node20249;
	wire [4-1:0] node20250;
	wire [4-1:0] node20251;
	wire [4-1:0] node20254;
	wire [4-1:0] node20255;
	wire [4-1:0] node20259;
	wire [4-1:0] node20260;
	wire [4-1:0] node20264;
	wire [4-1:0] node20265;
	wire [4-1:0] node20266;
	wire [4-1:0] node20268;
	wire [4-1:0] node20271;
	wire [4-1:0] node20273;
	wire [4-1:0] node20274;
	wire [4-1:0] node20278;
	wire [4-1:0] node20279;
	wire [4-1:0] node20280;
	wire [4-1:0] node20282;
	wire [4-1:0] node20285;
	wire [4-1:0] node20287;
	wire [4-1:0] node20290;
	wire [4-1:0] node20291;
	wire [4-1:0] node20293;
	wire [4-1:0] node20296;
	wire [4-1:0] node20297;
	wire [4-1:0] node20301;
	wire [4-1:0] node20302;
	wire [4-1:0] node20303;
	wire [4-1:0] node20304;
	wire [4-1:0] node20305;
	wire [4-1:0] node20309;
	wire [4-1:0] node20310;
	wire [4-1:0] node20312;
	wire [4-1:0] node20315;
	wire [4-1:0] node20318;
	wire [4-1:0] node20319;
	wire [4-1:0] node20321;
	wire [4-1:0] node20322;
	wire [4-1:0] node20326;
	wire [4-1:0] node20327;
	wire [4-1:0] node20329;
	wire [4-1:0] node20332;
	wire [4-1:0] node20333;
	wire [4-1:0] node20337;
	wire [4-1:0] node20338;
	wire [4-1:0] node20339;
	wire [4-1:0] node20340;
	wire [4-1:0] node20342;
	wire [4-1:0] node20345;
	wire [4-1:0] node20346;
	wire [4-1:0] node20350;
	wire [4-1:0] node20351;
	wire [4-1:0] node20352;
	wire [4-1:0] node20353;
	wire [4-1:0] node20357;
	wire [4-1:0] node20360;
	wire [4-1:0] node20361;
	wire [4-1:0] node20362;
	wire [4-1:0] node20366;
	wire [4-1:0] node20369;
	wire [4-1:0] node20370;
	wire [4-1:0] node20371;
	wire [4-1:0] node20372;
	wire [4-1:0] node20376;
	wire [4-1:0] node20378;
	wire [4-1:0] node20381;
	wire [4-1:0] node20383;
	wire [4-1:0] node20384;
	wire [4-1:0] node20386;
	wire [4-1:0] node20389;
	wire [4-1:0] node20391;
	wire [4-1:0] node20395;
	wire [4-1:0] node20396;
	wire [4-1:0] node20397;
	wire [4-1:0] node20398;
	wire [4-1:0] node20399;
	wire [4-1:0] node20400;
	wire [4-1:0] node20401;
	wire [4-1:0] node20402;
	wire [4-1:0] node20403;
	wire [4-1:0] node20404;
	wire [4-1:0] node20408;
	wire [4-1:0] node20409;
	wire [4-1:0] node20410;
	wire [4-1:0] node20415;
	wire [4-1:0] node20417;
	wire [4-1:0] node20420;
	wire [4-1:0] node20421;
	wire [4-1:0] node20422;
	wire [4-1:0] node20425;
	wire [4-1:0] node20427;
	wire [4-1:0] node20430;
	wire [4-1:0] node20432;
	wire [4-1:0] node20435;
	wire [4-1:0] node20436;
	wire [4-1:0] node20437;
	wire [4-1:0] node20438;
	wire [4-1:0] node20440;
	wire [4-1:0] node20443;
	wire [4-1:0] node20445;
	wire [4-1:0] node20448;
	wire [4-1:0] node20449;
	wire [4-1:0] node20450;
	wire [4-1:0] node20453;
	wire [4-1:0] node20455;
	wire [4-1:0] node20458;
	wire [4-1:0] node20459;
	wire [4-1:0] node20460;
	wire [4-1:0] node20464;
	wire [4-1:0] node20467;
	wire [4-1:0] node20468;
	wire [4-1:0] node20469;
	wire [4-1:0] node20470;
	wire [4-1:0] node20474;
	wire [4-1:0] node20475;
	wire [4-1:0] node20479;
	wire [4-1:0] node20481;
	wire [4-1:0] node20483;
	wire [4-1:0] node20486;
	wire [4-1:0] node20487;
	wire [4-1:0] node20488;
	wire [4-1:0] node20489;
	wire [4-1:0] node20490;
	wire [4-1:0] node20494;
	wire [4-1:0] node20495;
	wire [4-1:0] node20496;
	wire [4-1:0] node20500;
	wire [4-1:0] node20502;
	wire [4-1:0] node20505;
	wire [4-1:0] node20506;
	wire [4-1:0] node20507;
	wire [4-1:0] node20508;
	wire [4-1:0] node20509;
	wire [4-1:0] node20512;
	wire [4-1:0] node20515;
	wire [4-1:0] node20517;
	wire [4-1:0] node20521;
	wire [4-1:0] node20522;
	wire [4-1:0] node20524;
	wire [4-1:0] node20527;
	wire [4-1:0] node20528;
	wire [4-1:0] node20531;
	wire [4-1:0] node20534;
	wire [4-1:0] node20535;
	wire [4-1:0] node20536;
	wire [4-1:0] node20537;
	wire [4-1:0] node20538;
	wire [4-1:0] node20540;
	wire [4-1:0] node20543;
	wire [4-1:0] node20544;
	wire [4-1:0] node20548;
	wire [4-1:0] node20549;
	wire [4-1:0] node20550;
	wire [4-1:0] node20554;
	wire [4-1:0] node20557;
	wire [4-1:0] node20558;
	wire [4-1:0] node20560;
	wire [4-1:0] node20564;
	wire [4-1:0] node20565;
	wire [4-1:0] node20566;
	wire [4-1:0] node20568;
	wire [4-1:0] node20569;
	wire [4-1:0] node20573;
	wire [4-1:0] node20574;
	wire [4-1:0] node20577;
	wire [4-1:0] node20580;
	wire [4-1:0] node20581;
	wire [4-1:0] node20583;
	wire [4-1:0] node20586;
	wire [4-1:0] node20587;
	wire [4-1:0] node20591;
	wire [4-1:0] node20592;
	wire [4-1:0] node20593;
	wire [4-1:0] node20594;
	wire [4-1:0] node20595;
	wire [4-1:0] node20597;
	wire [4-1:0] node20598;
	wire [4-1:0] node20600;
	wire [4-1:0] node20604;
	wire [4-1:0] node20605;
	wire [4-1:0] node20606;
	wire [4-1:0] node20610;
	wire [4-1:0] node20612;
	wire [4-1:0] node20614;
	wire [4-1:0] node20617;
	wire [4-1:0] node20618;
	wire [4-1:0] node20619;
	wire [4-1:0] node20620;
	wire [4-1:0] node20623;
	wire [4-1:0] node20626;
	wire [4-1:0] node20627;
	wire [4-1:0] node20631;
	wire [4-1:0] node20632;
	wire [4-1:0] node20633;
	wire [4-1:0] node20637;
	wire [4-1:0] node20638;
	wire [4-1:0] node20642;
	wire [4-1:0] node20643;
	wire [4-1:0] node20644;
	wire [4-1:0] node20645;
	wire [4-1:0] node20646;
	wire [4-1:0] node20648;
	wire [4-1:0] node20651;
	wire [4-1:0] node20653;
	wire [4-1:0] node20656;
	wire [4-1:0] node20657;
	wire [4-1:0] node20659;
	wire [4-1:0] node20663;
	wire [4-1:0] node20664;
	wire [4-1:0] node20665;
	wire [4-1:0] node20668;
	wire [4-1:0] node20669;
	wire [4-1:0] node20673;
	wire [4-1:0] node20674;
	wire [4-1:0] node20677;
	wire [4-1:0] node20678;
	wire [4-1:0] node20682;
	wire [4-1:0] node20683;
	wire [4-1:0] node20684;
	wire [4-1:0] node20685;
	wire [4-1:0] node20689;
	wire [4-1:0] node20691;
	wire [4-1:0] node20694;
	wire [4-1:0] node20696;
	wire [4-1:0] node20699;
	wire [4-1:0] node20700;
	wire [4-1:0] node20702;
	wire [4-1:0] node20703;
	wire [4-1:0] node20704;
	wire [4-1:0] node20707;
	wire [4-1:0] node20710;
	wire [4-1:0] node20712;
	wire [4-1:0] node20716;
	wire [4-1:0] node20717;
	wire [4-1:0] node20718;
	wire [4-1:0] node20719;
	wire [4-1:0] node20720;
	wire [4-1:0] node20721;
	wire [4-1:0] node20722;
	wire [4-1:0] node20723;
	wire [4-1:0] node20726;
	wire [4-1:0] node20728;
	wire [4-1:0] node20731;
	wire [4-1:0] node20732;
	wire [4-1:0] node20735;
	wire [4-1:0] node20736;
	wire [4-1:0] node20739;
	wire [4-1:0] node20742;
	wire [4-1:0] node20743;
	wire [4-1:0] node20744;
	wire [4-1:0] node20747;
	wire [4-1:0] node20748;
	wire [4-1:0] node20751;
	wire [4-1:0] node20755;
	wire [4-1:0] node20756;
	wire [4-1:0] node20758;
	wire [4-1:0] node20760;
	wire [4-1:0] node20763;
	wire [4-1:0] node20764;
	wire [4-1:0] node20765;
	wire [4-1:0] node20768;
	wire [4-1:0] node20772;
	wire [4-1:0] node20773;
	wire [4-1:0] node20774;
	wire [4-1:0] node20775;
	wire [4-1:0] node20776;
	wire [4-1:0] node20779;
	wire [4-1:0] node20780;
	wire [4-1:0] node20784;
	wire [4-1:0] node20786;
	wire [4-1:0] node20789;
	wire [4-1:0] node20790;
	wire [4-1:0] node20791;
	wire [4-1:0] node20792;
	wire [4-1:0] node20797;
	wire [4-1:0] node20799;
	wire [4-1:0] node20801;
	wire [4-1:0] node20804;
	wire [4-1:0] node20805;
	wire [4-1:0] node20806;
	wire [4-1:0] node20807;
	wire [4-1:0] node20809;
	wire [4-1:0] node20812;
	wire [4-1:0] node20815;
	wire [4-1:0] node20816;
	wire [4-1:0] node20820;
	wire [4-1:0] node20821;
	wire [4-1:0] node20822;
	wire [4-1:0] node20824;
	wire [4-1:0] node20827;
	wire [4-1:0] node20831;
	wire [4-1:0] node20832;
	wire [4-1:0] node20833;
	wire [4-1:0] node20834;
	wire [4-1:0] node20835;
	wire [4-1:0] node20838;
	wire [4-1:0] node20841;
	wire [4-1:0] node20842;
	wire [4-1:0] node20844;
	wire [4-1:0] node20847;
	wire [4-1:0] node20848;
	wire [4-1:0] node20851;
	wire [4-1:0] node20854;
	wire [4-1:0] node20856;
	wire [4-1:0] node20857;
	wire [4-1:0] node20859;
	wire [4-1:0] node20860;
	wire [4-1:0] node20863;
	wire [4-1:0] node20867;
	wire [4-1:0] node20868;
	wire [4-1:0] node20869;
	wire [4-1:0] node20870;
	wire [4-1:0] node20871;
	wire [4-1:0] node20874;
	wire [4-1:0] node20877;
	wire [4-1:0] node20878;
	wire [4-1:0] node20881;
	wire [4-1:0] node20884;
	wire [4-1:0] node20885;
	wire [4-1:0] node20886;
	wire [4-1:0] node20889;
	wire [4-1:0] node20892;
	wire [4-1:0] node20893;
	wire [4-1:0] node20897;
	wire [4-1:0] node20898;
	wire [4-1:0] node20899;
	wire [4-1:0] node20903;
	wire [4-1:0] node20904;
	wire [4-1:0] node20905;
	wire [4-1:0] node20910;
	wire [4-1:0] node20911;
	wire [4-1:0] node20912;
	wire [4-1:0] node20913;
	wire [4-1:0] node20914;
	wire [4-1:0] node20915;
	wire [4-1:0] node20916;
	wire [4-1:0] node20917;
	wire [4-1:0] node20921;
	wire [4-1:0] node20922;
	wire [4-1:0] node20926;
	wire [4-1:0] node20927;
	wire [4-1:0] node20930;
	wire [4-1:0] node20933;
	wire [4-1:0] node20934;
	wire [4-1:0] node20935;
	wire [4-1:0] node20939;
	wire [4-1:0] node20940;
	wire [4-1:0] node20944;
	wire [4-1:0] node20945;
	wire [4-1:0] node20946;
	wire [4-1:0] node20947;
	wire [4-1:0] node20951;
	wire [4-1:0] node20953;
	wire [4-1:0] node20956;
	wire [4-1:0] node20957;
	wire [4-1:0] node20958;
	wire [4-1:0] node20962;
	wire [4-1:0] node20964;
	wire [4-1:0] node20967;
	wire [4-1:0] node20968;
	wire [4-1:0] node20969;
	wire [4-1:0] node20970;
	wire [4-1:0] node20971;
	wire [4-1:0] node20973;
	wire [4-1:0] node20976;
	wire [4-1:0] node20977;
	wire [4-1:0] node20981;
	wire [4-1:0] node20982;
	wire [4-1:0] node20983;
	wire [4-1:0] node20987;
	wire [4-1:0] node20990;
	wire [4-1:0] node20991;
	wire [4-1:0] node20992;
	wire [4-1:0] node20993;
	wire [4-1:0] node20996;
	wire [4-1:0] node20999;
	wire [4-1:0] node21000;
	wire [4-1:0] node21004;
	wire [4-1:0] node21005;
	wire [4-1:0] node21006;
	wire [4-1:0] node21010;
	wire [4-1:0] node21013;
	wire [4-1:0] node21014;
	wire [4-1:0] node21016;
	wire [4-1:0] node21017;
	wire [4-1:0] node21021;
	wire [4-1:0] node21022;
	wire [4-1:0] node21025;
	wire [4-1:0] node21027;
	wire [4-1:0] node21030;
	wire [4-1:0] node21031;
	wire [4-1:0] node21032;
	wire [4-1:0] node21033;
	wire [4-1:0] node21034;
	wire [4-1:0] node21035;
	wire [4-1:0] node21036;
	wire [4-1:0] node21039;
	wire [4-1:0] node21042;
	wire [4-1:0] node21043;
	wire [4-1:0] node21047;
	wire [4-1:0] node21048;
	wire [4-1:0] node21051;
	wire [4-1:0] node21053;
	wire [4-1:0] node21056;
	wire [4-1:0] node21057;
	wire [4-1:0] node21059;
	wire [4-1:0] node21062;
	wire [4-1:0] node21064;
	wire [4-1:0] node21065;
	wire [4-1:0] node21069;
	wire [4-1:0] node21070;
	wire [4-1:0] node21072;
	wire [4-1:0] node21075;
	wire [4-1:0] node21076;
	wire [4-1:0] node21080;
	wire [4-1:0] node21082;
	wire [4-1:0] node21083;
	wire [4-1:0] node21085;
	wire [4-1:0] node21086;
	wire [4-1:0] node21090;
	wire [4-1:0] node21091;
	wire [4-1:0] node21093;
	wire [4-1:0] node21095;
	wire [4-1:0] node21098;
	wire [4-1:0] node21100;
	wire [4-1:0] node21102;
	wire [4-1:0] node21105;
	wire [4-1:0] node21106;
	wire [4-1:0] node21107;
	wire [4-1:0] node21108;
	wire [4-1:0] node21109;
	wire [4-1:0] node21110;
	wire [4-1:0] node21111;
	wire [4-1:0] node21113;
	wire [4-1:0] node21116;
	wire [4-1:0] node21117;
	wire [4-1:0] node21118;
	wire [4-1:0] node21122;
	wire [4-1:0] node21123;
	wire [4-1:0] node21126;
	wire [4-1:0] node21127;
	wire [4-1:0] node21131;
	wire [4-1:0] node21132;
	wire [4-1:0] node21134;
	wire [4-1:0] node21135;
	wire [4-1:0] node21138;
	wire [4-1:0] node21140;
	wire [4-1:0] node21143;
	wire [4-1:0] node21144;
	wire [4-1:0] node21146;
	wire [4-1:0] node21149;
	wire [4-1:0] node21150;
	wire [4-1:0] node21154;
	wire [4-1:0] node21155;
	wire [4-1:0] node21156;
	wire [4-1:0] node21157;
	wire [4-1:0] node21159;
	wire [4-1:0] node21162;
	wire [4-1:0] node21163;
	wire [4-1:0] node21166;
	wire [4-1:0] node21168;
	wire [4-1:0] node21171;
	wire [4-1:0] node21172;
	wire [4-1:0] node21173;
	wire [4-1:0] node21174;
	wire [4-1:0] node21177;
	wire [4-1:0] node21182;
	wire [4-1:0] node21183;
	wire [4-1:0] node21184;
	wire [4-1:0] node21185;
	wire [4-1:0] node21188;
	wire [4-1:0] node21191;
	wire [4-1:0] node21192;
	wire [4-1:0] node21196;
	wire [4-1:0] node21197;
	wire [4-1:0] node21198;
	wire [4-1:0] node21201;
	wire [4-1:0] node21202;
	wire [4-1:0] node21206;
	wire [4-1:0] node21207;
	wire [4-1:0] node21211;
	wire [4-1:0] node21212;
	wire [4-1:0] node21213;
	wire [4-1:0] node21214;
	wire [4-1:0] node21215;
	wire [4-1:0] node21216;
	wire [4-1:0] node21217;
	wire [4-1:0] node21222;
	wire [4-1:0] node21224;
	wire [4-1:0] node21226;
	wire [4-1:0] node21229;
	wire [4-1:0] node21230;
	wire [4-1:0] node21231;
	wire [4-1:0] node21233;
	wire [4-1:0] node21236;
	wire [4-1:0] node21239;
	wire [4-1:0] node21240;
	wire [4-1:0] node21243;
	wire [4-1:0] node21246;
	wire [4-1:0] node21247;
	wire [4-1:0] node21248;
	wire [4-1:0] node21250;
	wire [4-1:0] node21251;
	wire [4-1:0] node21256;
	wire [4-1:0] node21257;
	wire [4-1:0] node21258;
	wire [4-1:0] node21259;
	wire [4-1:0] node21263;
	wire [4-1:0] node21264;
	wire [4-1:0] node21267;
	wire [4-1:0] node21270;
	wire [4-1:0] node21272;
	wire [4-1:0] node21275;
	wire [4-1:0] node21276;
	wire [4-1:0] node21277;
	wire [4-1:0] node21278;
	wire [4-1:0] node21279;
	wire [4-1:0] node21280;
	wire [4-1:0] node21284;
	wire [4-1:0] node21285;
	wire [4-1:0] node21288;
	wire [4-1:0] node21291;
	wire [4-1:0] node21292;
	wire [4-1:0] node21294;
	wire [4-1:0] node21297;
	wire [4-1:0] node21300;
	wire [4-1:0] node21301;
	wire [4-1:0] node21302;
	wire [4-1:0] node21305;
	wire [4-1:0] node21308;
	wire [4-1:0] node21309;
	wire [4-1:0] node21311;
	wire [4-1:0] node21314;
	wire [4-1:0] node21316;
	wire [4-1:0] node21319;
	wire [4-1:0] node21320;
	wire [4-1:0] node21321;
	wire [4-1:0] node21322;
	wire [4-1:0] node21326;
	wire [4-1:0] node21328;
	wire [4-1:0] node21330;
	wire [4-1:0] node21333;
	wire [4-1:0] node21334;
	wire [4-1:0] node21335;
	wire [4-1:0] node21337;
	wire [4-1:0] node21340;
	wire [4-1:0] node21342;
	wire [4-1:0] node21345;
	wire [4-1:0] node21346;
	wire [4-1:0] node21347;
	wire [4-1:0] node21351;
	wire [4-1:0] node21352;
	wire [4-1:0] node21356;
	wire [4-1:0] node21357;
	wire [4-1:0] node21358;
	wire [4-1:0] node21359;
	wire [4-1:0] node21360;
	wire [4-1:0] node21361;
	wire [4-1:0] node21362;
	wire [4-1:0] node21367;
	wire [4-1:0] node21368;
	wire [4-1:0] node21369;
	wire [4-1:0] node21373;
	wire [4-1:0] node21375;
	wire [4-1:0] node21378;
	wire [4-1:0] node21379;
	wire [4-1:0] node21380;
	wire [4-1:0] node21383;
	wire [4-1:0] node21384;
	wire [4-1:0] node21387;
	wire [4-1:0] node21390;
	wire [4-1:0] node21391;
	wire [4-1:0] node21393;
	wire [4-1:0] node21396;
	wire [4-1:0] node21398;
	wire [4-1:0] node21401;
	wire [4-1:0] node21402;
	wire [4-1:0] node21403;
	wire [4-1:0] node21404;
	wire [4-1:0] node21405;
	wire [4-1:0] node21409;
	wire [4-1:0] node21410;
	wire [4-1:0] node21414;
	wire [4-1:0] node21415;
	wire [4-1:0] node21417;
	wire [4-1:0] node21420;
	wire [4-1:0] node21422;
	wire [4-1:0] node21425;
	wire [4-1:0] node21426;
	wire [4-1:0] node21427;
	wire [4-1:0] node21428;
	wire [4-1:0] node21432;
	wire [4-1:0] node21434;
	wire [4-1:0] node21437;
	wire [4-1:0] node21438;
	wire [4-1:0] node21439;
	wire [4-1:0] node21443;
	wire [4-1:0] node21444;
	wire [4-1:0] node21447;
	wire [4-1:0] node21450;
	wire [4-1:0] node21451;
	wire [4-1:0] node21452;
	wire [4-1:0] node21453;
	wire [4-1:0] node21455;
	wire [4-1:0] node21457;
	wire [4-1:0] node21461;
	wire [4-1:0] node21462;
	wire [4-1:0] node21463;
	wire [4-1:0] node21466;
	wire [4-1:0] node21469;
	wire [4-1:0] node21470;
	wire [4-1:0] node21471;
	wire [4-1:0] node21476;
	wire [4-1:0] node21477;
	wire [4-1:0] node21478;
	wire [4-1:0] node21480;
	wire [4-1:0] node21481;
	wire [4-1:0] node21482;
	wire [4-1:0] node21485;
	wire [4-1:0] node21488;
	wire [4-1:0] node21490;
	wire [4-1:0] node21493;
	wire [4-1:0] node21494;
	wire [4-1:0] node21497;
	wire [4-1:0] node21499;
	wire [4-1:0] node21502;
	wire [4-1:0] node21504;
	wire [4-1:0] node21505;
	wire [4-1:0] node21506;
	wire [4-1:0] node21511;
	wire [4-1:0] node21512;
	wire [4-1:0] node21513;
	wire [4-1:0] node21514;
	wire [4-1:0] node21515;
	wire [4-1:0] node21516;
	wire [4-1:0] node21517;
	wire [4-1:0] node21518;
	wire [4-1:0] node21521;
	wire [4-1:0] node21523;
	wire [4-1:0] node21526;
	wire [4-1:0] node21529;
	wire [4-1:0] node21530;
	wire [4-1:0] node21532;
	wire [4-1:0] node21535;
	wire [4-1:0] node21536;
	wire [4-1:0] node21537;
	wire [4-1:0] node21541;
	wire [4-1:0] node21544;
	wire [4-1:0] node21545;
	wire [4-1:0] node21546;
	wire [4-1:0] node21548;
	wire [4-1:0] node21551;
	wire [4-1:0] node21552;
	wire [4-1:0] node21553;
	wire [4-1:0] node21557;
	wire [4-1:0] node21560;
	wire [4-1:0] node21561;
	wire [4-1:0] node21562;
	wire [4-1:0] node21565;
	wire [4-1:0] node21568;
	wire [4-1:0] node21570;
	wire [4-1:0] node21572;
	wire [4-1:0] node21575;
	wire [4-1:0] node21576;
	wire [4-1:0] node21577;
	wire [4-1:0] node21578;
	wire [4-1:0] node21580;
	wire [4-1:0] node21583;
	wire [4-1:0] node21585;
	wire [4-1:0] node21588;
	wire [4-1:0] node21589;
	wire [4-1:0] node21590;
	wire [4-1:0] node21592;
	wire [4-1:0] node21595;
	wire [4-1:0] node21598;
	wire [4-1:0] node21599;
	wire [4-1:0] node21602;
	wire [4-1:0] node21604;
	wire [4-1:0] node21607;
	wire [4-1:0] node21608;
	wire [4-1:0] node21609;
	wire [4-1:0] node21610;
	wire [4-1:0] node21611;
	wire [4-1:0] node21615;
	wire [4-1:0] node21616;
	wire [4-1:0] node21620;
	wire [4-1:0] node21622;
	wire [4-1:0] node21625;
	wire [4-1:0] node21626;
	wire [4-1:0] node21627;
	wire [4-1:0] node21629;
	wire [4-1:0] node21632;
	wire [4-1:0] node21634;
	wire [4-1:0] node21637;
	wire [4-1:0] node21638;
	wire [4-1:0] node21642;
	wire [4-1:0] node21643;
	wire [4-1:0] node21644;
	wire [4-1:0] node21645;
	wire [4-1:0] node21646;
	wire [4-1:0] node21649;
	wire [4-1:0] node21651;
	wire [4-1:0] node21654;
	wire [4-1:0] node21655;
	wire [4-1:0] node21657;
	wire [4-1:0] node21660;
	wire [4-1:0] node21663;
	wire [4-1:0] node21664;
	wire [4-1:0] node21665;
	wire [4-1:0] node21667;
	wire [4-1:0] node21670;
	wire [4-1:0] node21673;
	wire [4-1:0] node21674;
	wire [4-1:0] node21675;
	wire [4-1:0] node21678;
	wire [4-1:0] node21682;
	wire [4-1:0] node21683;
	wire [4-1:0] node21684;
	wire [4-1:0] node21685;
	wire [4-1:0] node21686;
	wire [4-1:0] node21687;
	wire [4-1:0] node21691;
	wire [4-1:0] node21693;
	wire [4-1:0] node21697;
	wire [4-1:0] node21698;
	wire [4-1:0] node21700;
	wire [4-1:0] node21703;
	wire [4-1:0] node21705;
	wire [4-1:0] node21709;
	wire [4-1:0] node21710;
	wire [4-1:0] node21711;
	wire [4-1:0] node21712;
	wire [4-1:0] node21713;
	wire [4-1:0] node21714;
	wire [4-1:0] node21715;
	wire [4-1:0] node21716;
	wire [4-1:0] node21721;
	wire [4-1:0] node21722;
	wire [4-1:0] node21724;
	wire [4-1:0] node21728;
	wire [4-1:0] node21729;
	wire [4-1:0] node21730;
	wire [4-1:0] node21732;
	wire [4-1:0] node21736;
	wire [4-1:0] node21737;
	wire [4-1:0] node21740;
	wire [4-1:0] node21743;
	wire [4-1:0] node21744;
	wire [4-1:0] node21745;
	wire [4-1:0] node21747;
	wire [4-1:0] node21750;
	wire [4-1:0] node21751;
	wire [4-1:0] node21752;
	wire [4-1:0] node21756;
	wire [4-1:0] node21757;
	wire [4-1:0] node21761;
	wire [4-1:0] node21762;
	wire [4-1:0] node21764;
	wire [4-1:0] node21766;
	wire [4-1:0] node21769;
	wire [4-1:0] node21770;
	wire [4-1:0] node21771;
	wire [4-1:0] node21775;
	wire [4-1:0] node21776;
	wire [4-1:0] node21780;
	wire [4-1:0] node21781;
	wire [4-1:0] node21782;
	wire [4-1:0] node21783;
	wire [4-1:0] node21784;
	wire [4-1:0] node21786;
	wire [4-1:0] node21789;
	wire [4-1:0] node21791;
	wire [4-1:0] node21794;
	wire [4-1:0] node21796;
	wire [4-1:0] node21799;
	wire [4-1:0] node21800;
	wire [4-1:0] node21801;
	wire [4-1:0] node21805;
	wire [4-1:0] node21806;
	wire [4-1:0] node21808;
	wire [4-1:0] node21811;
	wire [4-1:0] node21812;
	wire [4-1:0] node21815;
	wire [4-1:0] node21819;
	wire [4-1:0] node21820;
	wire [4-1:0] node21821;
	wire [4-1:0] node21822;
	wire [4-1:0] node21823;
	wire [4-1:0] node21825;
	wire [4-1:0] node21828;
	wire [4-1:0] node21829;
	wire [4-1:0] node21830;
	wire [4-1:0] node21833;
	wire [4-1:0] node21836;
	wire [4-1:0] node21837;
	wire [4-1:0] node21840;
	wire [4-1:0] node21843;
	wire [4-1:0] node21845;
	wire [4-1:0] node21846;
	wire [4-1:0] node21847;
	wire [4-1:0] node21851;
	wire [4-1:0] node21853;
	wire [4-1:0] node21858;
	wire [4-1:0] node21859;
	wire [4-1:0] node21860;
	wire [4-1:0] node21861;
	wire [4-1:0] node21863;
	wire [4-1:0] node21864;
	wire [4-1:0] node21865;
	wire [4-1:0] node21866;
	wire [4-1:0] node21868;
	wire [4-1:0] node21869;
	wire [4-1:0] node21870;
	wire [4-1:0] node21873;
	wire [4-1:0] node21874;
	wire [4-1:0] node21876;
	wire [4-1:0] node21879;
	wire [4-1:0] node21882;
	wire [4-1:0] node21884;
	wire [4-1:0] node21886;
	wire [4-1:0] node21888;
	wire [4-1:0] node21892;
	wire [4-1:0] node21893;
	wire [4-1:0] node21894;
	wire [4-1:0] node21895;
	wire [4-1:0] node21896;
	wire [4-1:0] node21897;
	wire [4-1:0] node21901;
	wire [4-1:0] node21903;
	wire [4-1:0] node21906;
	wire [4-1:0] node21907;
	wire [4-1:0] node21908;
	wire [4-1:0] node21910;
	wire [4-1:0] node21913;
	wire [4-1:0] node21915;
	wire [4-1:0] node21918;
	wire [4-1:0] node21920;
	wire [4-1:0] node21923;
	wire [4-1:0] node21924;
	wire [4-1:0] node21925;
	wire [4-1:0] node21927;
	wire [4-1:0] node21930;
	wire [4-1:0] node21931;
	wire [4-1:0] node21935;
	wire [4-1:0] node21936;
	wire [4-1:0] node21937;
	wire [4-1:0] node21939;
	wire [4-1:0] node21942;
	wire [4-1:0] node21944;
	wire [4-1:0] node21947;
	wire [4-1:0] node21948;
	wire [4-1:0] node21950;
	wire [4-1:0] node21954;
	wire [4-1:0] node21956;
	wire [4-1:0] node21957;
	wire [4-1:0] node21959;
	wire [4-1:0] node21960;
	wire [4-1:0] node21964;
	wire [4-1:0] node21965;
	wire [4-1:0] node21966;
	wire [4-1:0] node21968;
	wire [4-1:0] node21971;
	wire [4-1:0] node21974;
	wire [4-1:0] node21976;
	wire [4-1:0] node21977;
	wire [4-1:0] node21982;
	wire [4-1:0] node21983;
	wire [4-1:0] node21984;
	wire [4-1:0] node21985;
	wire [4-1:0] node21986;
	wire [4-1:0] node21987;
	wire [4-1:0] node21988;
	wire [4-1:0] node21989;
	wire [4-1:0] node21992;
	wire [4-1:0] node21994;
	wire [4-1:0] node21997;
	wire [4-1:0] node21998;
	wire [4-1:0] node21999;
	wire [4-1:0] node22002;
	wire [4-1:0] node22004;
	wire [4-1:0] node22007;
	wire [4-1:0] node22009;
	wire [4-1:0] node22012;
	wire [4-1:0] node22013;
	wire [4-1:0] node22014;
	wire [4-1:0] node22016;
	wire [4-1:0] node22019;
	wire [4-1:0] node22021;
	wire [4-1:0] node22024;
	wire [4-1:0] node22026;
	wire [4-1:0] node22029;
	wire [4-1:0] node22030;
	wire [4-1:0] node22031;
	wire [4-1:0] node22032;
	wire [4-1:0] node22034;
	wire [4-1:0] node22037;
	wire [4-1:0] node22039;
	wire [4-1:0] node22042;
	wire [4-1:0] node22044;
	wire [4-1:0] node22047;
	wire [4-1:0] node22048;
	wire [4-1:0] node22050;
	wire [4-1:0] node22051;
	wire [4-1:0] node22054;
	wire [4-1:0] node22056;
	wire [4-1:0] node22059;
	wire [4-1:0] node22060;
	wire [4-1:0] node22063;
	wire [4-1:0] node22065;
	wire [4-1:0] node22068;
	wire [4-1:0] node22069;
	wire [4-1:0] node22070;
	wire [4-1:0] node22071;
	wire [4-1:0] node22072;
	wire [4-1:0] node22073;
	wire [4-1:0] node22074;
	wire [4-1:0] node22079;
	wire [4-1:0] node22080;
	wire [4-1:0] node22083;
	wire [4-1:0] node22084;
	wire [4-1:0] node22088;
	wire [4-1:0] node22089;
	wire [4-1:0] node22091;
	wire [4-1:0] node22095;
	wire [4-1:0] node22096;
	wire [4-1:0] node22098;
	wire [4-1:0] node22101;
	wire [4-1:0] node22102;
	wire [4-1:0] node22106;
	wire [4-1:0] node22107;
	wire [4-1:0] node22108;
	wire [4-1:0] node22109;
	wire [4-1:0] node22111;
	wire [4-1:0] node22114;
	wire [4-1:0] node22116;
	wire [4-1:0] node22119;
	wire [4-1:0] node22120;
	wire [4-1:0] node22123;
	wire [4-1:0] node22124;
	wire [4-1:0] node22126;
	wire [4-1:0] node22130;
	wire [4-1:0] node22131;
	wire [4-1:0] node22132;
	wire [4-1:0] node22133;
	wire [4-1:0] node22134;
	wire [4-1:0] node22139;
	wire [4-1:0] node22142;
	wire [4-1:0] node22143;
	wire [4-1:0] node22145;
	wire [4-1:0] node22148;
	wire [4-1:0] node22150;
	wire [4-1:0] node22153;
	wire [4-1:0] node22154;
	wire [4-1:0] node22155;
	wire [4-1:0] node22156;
	wire [4-1:0] node22157;
	wire [4-1:0] node22158;
	wire [4-1:0] node22159;
	wire [4-1:0] node22163;
	wire [4-1:0] node22164;
	wire [4-1:0] node22168;
	wire [4-1:0] node22170;
	wire [4-1:0] node22173;
	wire [4-1:0] node22174;
	wire [4-1:0] node22175;
	wire [4-1:0] node22177;
	wire [4-1:0] node22179;
	wire [4-1:0] node22183;
	wire [4-1:0] node22184;
	wire [4-1:0] node22188;
	wire [4-1:0] node22189;
	wire [4-1:0] node22190;
	wire [4-1:0] node22191;
	wire [4-1:0] node22193;
	wire [4-1:0] node22196;
	wire [4-1:0] node22198;
	wire [4-1:0] node22201;
	wire [4-1:0] node22202;
	wire [4-1:0] node22206;
	wire [4-1:0] node22207;
	wire [4-1:0] node22209;
	wire [4-1:0] node22212;
	wire [4-1:0] node22214;
	wire [4-1:0] node22217;
	wire [4-1:0] node22218;
	wire [4-1:0] node22219;
	wire [4-1:0] node22220;
	wire [4-1:0] node22221;
	wire [4-1:0] node22223;
	wire [4-1:0] node22226;
	wire [4-1:0] node22229;
	wire [4-1:0] node22230;
	wire [4-1:0] node22231;
	wire [4-1:0] node22234;
	wire [4-1:0] node22236;
	wire [4-1:0] node22239;
	wire [4-1:0] node22240;
	wire [4-1:0] node22244;
	wire [4-1:0] node22245;
	wire [4-1:0] node22246;
	wire [4-1:0] node22247;
	wire [4-1:0] node22250;
	wire [4-1:0] node22252;
	wire [4-1:0] node22255;
	wire [4-1:0] node22257;
	wire [4-1:0] node22259;
	wire [4-1:0] node22262;
	wire [4-1:0] node22263;
	wire [4-1:0] node22264;
	wire [4-1:0] node22268;
	wire [4-1:0] node22269;
	wire [4-1:0] node22273;
	wire [4-1:0] node22274;
	wire [4-1:0] node22275;
	wire [4-1:0] node22276;
	wire [4-1:0] node22277;
	wire [4-1:0] node22281;
	wire [4-1:0] node22284;
	wire [4-1:0] node22285;
	wire [4-1:0] node22286;
	wire [4-1:0] node22288;
	wire [4-1:0] node22292;
	wire [4-1:0] node22295;
	wire [4-1:0] node22296;
	wire [4-1:0] node22297;
	wire [4-1:0] node22298;
	wire [4-1:0] node22301;
	wire [4-1:0] node22305;
	wire [4-1:0] node22306;
	wire [4-1:0] node22308;
	wire [4-1:0] node22311;
	wire [4-1:0] node22313;
	wire [4-1:0] node22316;
	wire [4-1:0] node22318;
	wire [4-1:0] node22319;
	wire [4-1:0] node22320;
	wire [4-1:0] node22322;
	wire [4-1:0] node22323;
	wire [4-1:0] node22324;
	wire [4-1:0] node22328;
	wire [4-1:0] node22330;
	wire [4-1:0] node22332;
	wire [4-1:0] node22333;
	wire [4-1:0] node22338;
	wire [4-1:0] node22339;
	wire [4-1:0] node22340;
	wire [4-1:0] node22341;
	wire [4-1:0] node22342;
	wire [4-1:0] node22343;
	wire [4-1:0] node22346;
	wire [4-1:0] node22349;
	wire [4-1:0] node22351;
	wire [4-1:0] node22352;
	wire [4-1:0] node22355;
	wire [4-1:0] node22358;
	wire [4-1:0] node22359;
	wire [4-1:0] node22361;
	wire [4-1:0] node22364;
	wire [4-1:0] node22366;
	wire [4-1:0] node22369;
	wire [4-1:0] node22370;
	wire [4-1:0] node22371;
	wire [4-1:0] node22372;
	wire [4-1:0] node22374;
	wire [4-1:0] node22377;
	wire [4-1:0] node22380;
	wire [4-1:0] node22381;
	wire [4-1:0] node22383;
	wire [4-1:0] node22386;
	wire [4-1:0] node22388;
	wire [4-1:0] node22391;
	wire [4-1:0] node22392;
	wire [4-1:0] node22393;
	wire [4-1:0] node22397;
	wire [4-1:0] node22399;
	wire [4-1:0] node22402;
	wire [4-1:0] node22404;
	wire [4-1:0] node22405;
	wire [4-1:0] node22406;
	wire [4-1:0] node22407;
	wire [4-1:0] node22408;
	wire [4-1:0] node22413;
	wire [4-1:0] node22416;
	wire [4-1:0] node22418;
	wire [4-1:0] node22421;
	wire [4-1:0] node22422;
	wire [4-1:0] node22423;
	wire [4-1:0] node22424;
	wire [4-1:0] node22425;
	wire [4-1:0] node22426;
	wire [4-1:0] node22427;
	wire [4-1:0] node22428;
	wire [4-1:0] node22431;
	wire [4-1:0] node22432;
	wire [4-1:0] node22436;
	wire [4-1:0] node22437;
	wire [4-1:0] node22438;
	wire [4-1:0] node22441;
	wire [4-1:0] node22444;
	wire [4-1:0] node22445;
	wire [4-1:0] node22448;
	wire [4-1:0] node22451;
	wire [4-1:0] node22452;
	wire [4-1:0] node22453;
	wire [4-1:0] node22454;
	wire [4-1:0] node22457;
	wire [4-1:0] node22458;
	wire [4-1:0] node22462;
	wire [4-1:0] node22463;
	wire [4-1:0] node22464;
	wire [4-1:0] node22465;
	wire [4-1:0] node22469;
	wire [4-1:0] node22470;
	wire [4-1:0] node22473;
	wire [4-1:0] node22476;
	wire [4-1:0] node22477;
	wire [4-1:0] node22480;
	wire [4-1:0] node22483;
	wire [4-1:0] node22484;
	wire [4-1:0] node22487;
	wire [4-1:0] node22488;
	wire [4-1:0] node22492;
	wire [4-1:0] node22493;
	wire [4-1:0] node22494;
	wire [4-1:0] node22495;
	wire [4-1:0] node22496;
	wire [4-1:0] node22497;
	wire [4-1:0] node22500;
	wire [4-1:0] node22503;
	wire [4-1:0] node22504;
	wire [4-1:0] node22507;
	wire [4-1:0] node22508;
	wire [4-1:0] node22512;
	wire [4-1:0] node22513;
	wire [4-1:0] node22515;
	wire [4-1:0] node22518;
	wire [4-1:0] node22521;
	wire [4-1:0] node22522;
	wire [4-1:0] node22523;
	wire [4-1:0] node22525;
	wire [4-1:0] node22528;
	wire [4-1:0] node22529;
	wire [4-1:0] node22533;
	wire [4-1:0] node22534;
	wire [4-1:0] node22535;
	wire [4-1:0] node22536;
	wire [4-1:0] node22540;
	wire [4-1:0] node22543;
	wire [4-1:0] node22544;
	wire [4-1:0] node22545;
	wire [4-1:0] node22548;
	wire [4-1:0] node22551;
	wire [4-1:0] node22553;
	wire [4-1:0] node22556;
	wire [4-1:0] node22557;
	wire [4-1:0] node22558;
	wire [4-1:0] node22559;
	wire [4-1:0] node22560;
	wire [4-1:0] node22563;
	wire [4-1:0] node22566;
	wire [4-1:0] node22567;
	wire [4-1:0] node22571;
	wire [4-1:0] node22572;
	wire [4-1:0] node22573;
	wire [4-1:0] node22576;
	wire [4-1:0] node22579;
	wire [4-1:0] node22580;
	wire [4-1:0] node22581;
	wire [4-1:0] node22584;
	wire [4-1:0] node22587;
	wire [4-1:0] node22589;
	wire [4-1:0] node22592;
	wire [4-1:0] node22593;
	wire [4-1:0] node22594;
	wire [4-1:0] node22596;
	wire [4-1:0] node22599;
	wire [4-1:0] node22602;
	wire [4-1:0] node22603;
	wire [4-1:0] node22604;
	wire [4-1:0] node22605;
	wire [4-1:0] node22609;
	wire [4-1:0] node22610;
	wire [4-1:0] node22614;
	wire [4-1:0] node22615;
	wire [4-1:0] node22616;
	wire [4-1:0] node22619;
	wire [4-1:0] node22623;
	wire [4-1:0] node22624;
	wire [4-1:0] node22625;
	wire [4-1:0] node22626;
	wire [4-1:0] node22627;
	wire [4-1:0] node22628;
	wire [4-1:0] node22632;
	wire [4-1:0] node22633;
	wire [4-1:0] node22635;
	wire [4-1:0] node22638;
	wire [4-1:0] node22639;
	wire [4-1:0] node22643;
	wire [4-1:0] node22644;
	wire [4-1:0] node22646;
	wire [4-1:0] node22647;
	wire [4-1:0] node22648;
	wire [4-1:0] node22651;
	wire [4-1:0] node22655;
	wire [4-1:0] node22656;
	wire [4-1:0] node22660;
	wire [4-1:0] node22661;
	wire [4-1:0] node22662;
	wire [4-1:0] node22663;
	wire [4-1:0] node22667;
	wire [4-1:0] node22669;
	wire [4-1:0] node22670;
	wire [4-1:0] node22672;
	wire [4-1:0] node22676;
	wire [4-1:0] node22677;
	wire [4-1:0] node22678;
	wire [4-1:0] node22680;
	wire [4-1:0] node22683;
	wire [4-1:0] node22684;
	wire [4-1:0] node22687;
	wire [4-1:0] node22690;
	wire [4-1:0] node22691;
	wire [4-1:0] node22692;
	wire [4-1:0] node22697;
	wire [4-1:0] node22698;
	wire [4-1:0] node22699;
	wire [4-1:0] node22700;
	wire [4-1:0] node22701;
	wire [4-1:0] node22702;
	wire [4-1:0] node22704;
	wire [4-1:0] node22707;
	wire [4-1:0] node22710;
	wire [4-1:0] node22711;
	wire [4-1:0] node22714;
	wire [4-1:0] node22715;
	wire [4-1:0] node22719;
	wire [4-1:0] node22720;
	wire [4-1:0] node22721;
	wire [4-1:0] node22724;
	wire [4-1:0] node22725;
	wire [4-1:0] node22728;
	wire [4-1:0] node22731;
	wire [4-1:0] node22732;
	wire [4-1:0] node22733;
	wire [4-1:0] node22736;
	wire [4-1:0] node22739;
	wire [4-1:0] node22741;
	wire [4-1:0] node22744;
	wire [4-1:0] node22745;
	wire [4-1:0] node22746;
	wire [4-1:0] node22747;
	wire [4-1:0] node22750;
	wire [4-1:0] node22753;
	wire [4-1:0] node22754;
	wire [4-1:0] node22756;
	wire [4-1:0] node22760;
	wire [4-1:0] node22761;
	wire [4-1:0] node22762;
	wire [4-1:0] node22766;
	wire [4-1:0] node22767;
	wire [4-1:0] node22771;
	wire [4-1:0] node22772;
	wire [4-1:0] node22773;
	wire [4-1:0] node22774;
	wire [4-1:0] node22775;
	wire [4-1:0] node22777;
	wire [4-1:0] node22780;
	wire [4-1:0] node22781;
	wire [4-1:0] node22785;
	wire [4-1:0] node22786;
	wire [4-1:0] node22789;
	wire [4-1:0] node22792;
	wire [4-1:0] node22793;
	wire [4-1:0] node22795;
	wire [4-1:0] node22798;
	wire [4-1:0] node22799;
	wire [4-1:0] node22802;
	wire [4-1:0] node22805;
	wire [4-1:0] node22806;
	wire [4-1:0] node22807;
	wire [4-1:0] node22808;
	wire [4-1:0] node22810;
	wire [4-1:0] node22813;
	wire [4-1:0] node22816;
	wire [4-1:0] node22817;
	wire [4-1:0] node22818;
	wire [4-1:0] node22822;
	wire [4-1:0] node22825;
	wire [4-1:0] node22826;
	wire [4-1:0] node22828;
	wire [4-1:0] node22831;
	wire [4-1:0] node22834;
	wire [4-1:0] node22835;
	wire [4-1:0] node22836;
	wire [4-1:0] node22837;
	wire [4-1:0] node22838;
	wire [4-1:0] node22839;
	wire [4-1:0] node22840;
	wire [4-1:0] node22844;
	wire [4-1:0] node22846;
	wire [4-1:0] node22847;
	wire [4-1:0] node22850;
	wire [4-1:0] node22853;
	wire [4-1:0] node22855;
	wire [4-1:0] node22858;
	wire [4-1:0] node22859;
	wire [4-1:0] node22860;
	wire [4-1:0] node22861;
	wire [4-1:0] node22863;
	wire [4-1:0] node22866;
	wire [4-1:0] node22870;
	wire [4-1:0] node22871;
	wire [4-1:0] node22872;
	wire [4-1:0] node22873;
	wire [4-1:0] node22877;
	wire [4-1:0] node22879;
	wire [4-1:0] node22882;
	wire [4-1:0] node22884;
	wire [4-1:0] node22885;
	wire [4-1:0] node22889;
	wire [4-1:0] node22890;
	wire [4-1:0] node22891;
	wire [4-1:0] node22892;
	wire [4-1:0] node22893;
	wire [4-1:0] node22896;
	wire [4-1:0] node22897;
	wire [4-1:0] node22900;
	wire [4-1:0] node22903;
	wire [4-1:0] node22904;
	wire [4-1:0] node22907;
	wire [4-1:0] node22908;
	wire [4-1:0] node22912;
	wire [4-1:0] node22913;
	wire [4-1:0] node22914;
	wire [4-1:0] node22915;
	wire [4-1:0] node22918;
	wire [4-1:0] node22921;
	wire [4-1:0] node22922;
	wire [4-1:0] node22926;
	wire [4-1:0] node22927;
	wire [4-1:0] node22930;
	wire [4-1:0] node22931;
	wire [4-1:0] node22935;
	wire [4-1:0] node22936;
	wire [4-1:0] node22937;
	wire [4-1:0] node22939;
	wire [4-1:0] node22942;
	wire [4-1:0] node22944;
	wire [4-1:0] node22945;
	wire [4-1:0] node22949;
	wire [4-1:0] node22950;
	wire [4-1:0] node22951;
	wire [4-1:0] node22952;
	wire [4-1:0] node22956;
	wire [4-1:0] node22957;
	wire [4-1:0] node22960;
	wire [4-1:0] node22963;
	wire [4-1:0] node22964;
	wire [4-1:0] node22966;
	wire [4-1:0] node22969;
	wire [4-1:0] node22970;
	wire [4-1:0] node22974;
	wire [4-1:0] node22975;
	wire [4-1:0] node22976;
	wire [4-1:0] node22977;
	wire [4-1:0] node22978;
	wire [4-1:0] node22980;
	wire [4-1:0] node22982;
	wire [4-1:0] node22986;
	wire [4-1:0] node22987;
	wire [4-1:0] node22989;
	wire [4-1:0] node22992;
	wire [4-1:0] node22994;
	wire [4-1:0] node22995;
	wire [4-1:0] node22998;
	wire [4-1:0] node23001;
	wire [4-1:0] node23002;
	wire [4-1:0] node23003;
	wire [4-1:0] node23004;
	wire [4-1:0] node23007;
	wire [4-1:0] node23008;
	wire [4-1:0] node23012;
	wire [4-1:0] node23013;
	wire [4-1:0] node23015;
	wire [4-1:0] node23019;
	wire [4-1:0] node23020;
	wire [4-1:0] node23021;
	wire [4-1:0] node23024;
	wire [4-1:0] node23027;
	wire [4-1:0] node23029;
	wire [4-1:0] node23032;
	wire [4-1:0] node23033;
	wire [4-1:0] node23034;
	wire [4-1:0] node23035;
	wire [4-1:0] node23036;
	wire [4-1:0] node23038;
	wire [4-1:0] node23042;
	wire [4-1:0] node23043;
	wire [4-1:0] node23044;
	wire [4-1:0] node23047;
	wire [4-1:0] node23050;
	wire [4-1:0] node23051;
	wire [4-1:0] node23055;
	wire [4-1:0] node23056;
	wire [4-1:0] node23058;
	wire [4-1:0] node23059;
	wire [4-1:0] node23063;
	wire [4-1:0] node23064;
	wire [4-1:0] node23065;
	wire [4-1:0] node23068;
	wire [4-1:0] node23071;
	wire [4-1:0] node23073;
	wire [4-1:0] node23076;
	wire [4-1:0] node23077;
	wire [4-1:0] node23078;
	wire [4-1:0] node23079;
	wire [4-1:0] node23083;
	wire [4-1:0] node23084;
	wire [4-1:0] node23086;
	wire [4-1:0] node23089;
	wire [4-1:0] node23090;
	wire [4-1:0] node23093;
	wire [4-1:0] node23096;
	wire [4-1:0] node23097;
	wire [4-1:0] node23101;
	wire [4-1:0] node23102;
	wire [4-1:0] node23103;
	wire [4-1:0] node23104;
	wire [4-1:0] node23105;
	wire [4-1:0] node23106;
	wire [4-1:0] node23107;
	wire [4-1:0] node23108;
	wire [4-1:0] node23111;
	wire [4-1:0] node23114;
	wire [4-1:0] node23115;
	wire [4-1:0] node23116;
	wire [4-1:0] node23118;
	wire [4-1:0] node23121;
	wire [4-1:0] node23122;
	wire [4-1:0] node23126;
	wire [4-1:0] node23127;
	wire [4-1:0] node23128;
	wire [4-1:0] node23132;
	wire [4-1:0] node23133;
	wire [4-1:0] node23137;
	wire [4-1:0] node23138;
	wire [4-1:0] node23139;
	wire [4-1:0] node23140;
	wire [4-1:0] node23141;
	wire [4-1:0] node23145;
	wire [4-1:0] node23147;
	wire [4-1:0] node23150;
	wire [4-1:0] node23151;
	wire [4-1:0] node23154;
	wire [4-1:0] node23157;
	wire [4-1:0] node23158;
	wire [4-1:0] node23159;
	wire [4-1:0] node23161;
	wire [4-1:0] node23164;
	wire [4-1:0] node23166;
	wire [4-1:0] node23169;
	wire [4-1:0] node23170;
	wire [4-1:0] node23173;
	wire [4-1:0] node23174;
	wire [4-1:0] node23177;
	wire [4-1:0] node23180;
	wire [4-1:0] node23181;
	wire [4-1:0] node23182;
	wire [4-1:0] node23183;
	wire [4-1:0] node23187;
	wire [4-1:0] node23189;
	wire [4-1:0] node23190;
	wire [4-1:0] node23194;
	wire [4-1:0] node23195;
	wire [4-1:0] node23196;
	wire [4-1:0] node23197;
	wire [4-1:0] node23201;
	wire [4-1:0] node23203;
	wire [4-1:0] node23204;
	wire [4-1:0] node23208;
	wire [4-1:0] node23210;
	wire [4-1:0] node23211;
	wire [4-1:0] node23215;
	wire [4-1:0] node23216;
	wire [4-1:0] node23217;
	wire [4-1:0] node23218;
	wire [4-1:0] node23219;
	wire [4-1:0] node23221;
	wire [4-1:0] node23224;
	wire [4-1:0] node23227;
	wire [4-1:0] node23228;
	wire [4-1:0] node23229;
	wire [4-1:0] node23232;
	wire [4-1:0] node23233;
	wire [4-1:0] node23237;
	wire [4-1:0] node23238;
	wire [4-1:0] node23241;
	wire [4-1:0] node23244;
	wire [4-1:0] node23245;
	wire [4-1:0] node23246;
	wire [4-1:0] node23247;
	wire [4-1:0] node23250;
	wire [4-1:0] node23253;
	wire [4-1:0] node23255;
	wire [4-1:0] node23256;
	wire [4-1:0] node23260;
	wire [4-1:0] node23261;
	wire [4-1:0] node23264;
	wire [4-1:0] node23267;
	wire [4-1:0] node23268;
	wire [4-1:0] node23269;
	wire [4-1:0] node23270;
	wire [4-1:0] node23271;
	wire [4-1:0] node23272;
	wire [4-1:0] node23276;
	wire [4-1:0] node23279;
	wire [4-1:0] node23281;
	wire [4-1:0] node23284;
	wire [4-1:0] node23285;
	wire [4-1:0] node23286;
	wire [4-1:0] node23287;
	wire [4-1:0] node23292;
	wire [4-1:0] node23293;
	wire [4-1:0] node23294;
	wire [4-1:0] node23298;
	wire [4-1:0] node23301;
	wire [4-1:0] node23302;
	wire [4-1:0] node23303;
	wire [4-1:0] node23304;
	wire [4-1:0] node23307;
	wire [4-1:0] node23310;
	wire [4-1:0] node23311;
	wire [4-1:0] node23314;
	wire [4-1:0] node23317;
	wire [4-1:0] node23318;
	wire [4-1:0] node23319;
	wire [4-1:0] node23322;
	wire [4-1:0] node23325;
	wire [4-1:0] node23326;
	wire [4-1:0] node23329;
	wire [4-1:0] node23332;
	wire [4-1:0] node23333;
	wire [4-1:0] node23334;
	wire [4-1:0] node23335;
	wire [4-1:0] node23336;
	wire [4-1:0] node23337;
	wire [4-1:0] node23340;
	wire [4-1:0] node23343;
	wire [4-1:0] node23344;
	wire [4-1:0] node23346;
	wire [4-1:0] node23349;
	wire [4-1:0] node23352;
	wire [4-1:0] node23353;
	wire [4-1:0] node23354;
	wire [4-1:0] node23357;
	wire [4-1:0] node23360;
	wire [4-1:0] node23361;
	wire [4-1:0] node23363;
	wire [4-1:0] node23366;
	wire [4-1:0] node23367;
	wire [4-1:0] node23370;
	wire [4-1:0] node23373;
	wire [4-1:0] node23374;
	wire [4-1:0] node23375;
	wire [4-1:0] node23376;
	wire [4-1:0] node23377;
	wire [4-1:0] node23380;
	wire [4-1:0] node23384;
	wire [4-1:0] node23385;
	wire [4-1:0] node23387;
	wire [4-1:0] node23391;
	wire [4-1:0] node23392;
	wire [4-1:0] node23393;
	wire [4-1:0] node23394;
	wire [4-1:0] node23398;
	wire [4-1:0] node23401;
	wire [4-1:0] node23402;
	wire [4-1:0] node23404;
	wire [4-1:0] node23407;
	wire [4-1:0] node23409;
	wire [4-1:0] node23412;
	wire [4-1:0] node23413;
	wire [4-1:0] node23414;
	wire [4-1:0] node23415;
	wire [4-1:0] node23416;
	wire [4-1:0] node23418;
	wire [4-1:0] node23422;
	wire [4-1:0] node23423;
	wire [4-1:0] node23426;
	wire [4-1:0] node23429;
	wire [4-1:0] node23430;
	wire [4-1:0] node23431;
	wire [4-1:0] node23435;
	wire [4-1:0] node23436;
	wire [4-1:0] node23438;
	wire [4-1:0] node23441;
	wire [4-1:0] node23444;
	wire [4-1:0] node23445;
	wire [4-1:0] node23446;
	wire [4-1:0] node23447;
	wire [4-1:0] node23449;
	wire [4-1:0] node23452;
	wire [4-1:0] node23455;
	wire [4-1:0] node23456;
	wire [4-1:0] node23457;
	wire [4-1:0] node23461;
	wire [4-1:0] node23462;
	wire [4-1:0] node23465;
	wire [4-1:0] node23468;
	wire [4-1:0] node23469;
	wire [4-1:0] node23471;
	wire [4-1:0] node23475;
	wire [4-1:0] node23476;
	wire [4-1:0] node23477;
	wire [4-1:0] node23478;
	wire [4-1:0] node23479;
	wire [4-1:0] node23480;
	wire [4-1:0] node23481;
	wire [4-1:0] node23482;
	wire [4-1:0] node23485;
	wire [4-1:0] node23486;
	wire [4-1:0] node23490;
	wire [4-1:0] node23491;
	wire [4-1:0] node23494;
	wire [4-1:0] node23495;
	wire [4-1:0] node23499;
	wire [4-1:0] node23500;
	wire [4-1:0] node23502;
	wire [4-1:0] node23503;
	wire [4-1:0] node23508;
	wire [4-1:0] node23509;
	wire [4-1:0] node23510;
	wire [4-1:0] node23511;
	wire [4-1:0] node23515;
	wire [4-1:0] node23516;
	wire [4-1:0] node23517;
	wire [4-1:0] node23521;
	wire [4-1:0] node23522;
	wire [4-1:0] node23525;
	wire [4-1:0] node23528;
	wire [4-1:0] node23529;
	wire [4-1:0] node23531;
	wire [4-1:0] node23534;
	wire [4-1:0] node23535;
	wire [4-1:0] node23538;
	wire [4-1:0] node23541;
	wire [4-1:0] node23542;
	wire [4-1:0] node23543;
	wire [4-1:0] node23544;
	wire [4-1:0] node23548;
	wire [4-1:0] node23549;
	wire [4-1:0] node23551;
	wire [4-1:0] node23553;
	wire [4-1:0] node23556;
	wire [4-1:0] node23558;
	wire [4-1:0] node23561;
	wire [4-1:0] node23562;
	wire [4-1:0] node23563;
	wire [4-1:0] node23564;
	wire [4-1:0] node23568;
	wire [4-1:0] node23569;
	wire [4-1:0] node23573;
	wire [4-1:0] node23574;
	wire [4-1:0] node23575;
	wire [4-1:0] node23578;
	wire [4-1:0] node23579;
	wire [4-1:0] node23583;
	wire [4-1:0] node23584;
	wire [4-1:0] node23587;
	wire [4-1:0] node23588;
	wire [4-1:0] node23592;
	wire [4-1:0] node23593;
	wire [4-1:0] node23594;
	wire [4-1:0] node23595;
	wire [4-1:0] node23596;
	wire [4-1:0] node23597;
	wire [4-1:0] node23598;
	wire [4-1:0] node23602;
	wire [4-1:0] node23603;
	wire [4-1:0] node23607;
	wire [4-1:0] node23608;
	wire [4-1:0] node23612;
	wire [4-1:0] node23615;
	wire [4-1:0] node23616;
	wire [4-1:0] node23617;
	wire [4-1:0] node23618;
	wire [4-1:0] node23620;
	wire [4-1:0] node23624;
	wire [4-1:0] node23625;
	wire [4-1:0] node23626;
	wire [4-1:0] node23629;
	wire [4-1:0] node23633;
	wire [4-1:0] node23634;
	wire [4-1:0] node23635;
	wire [4-1:0] node23638;
	wire [4-1:0] node23641;
	wire [4-1:0] node23644;
	wire [4-1:0] node23645;
	wire [4-1:0] node23646;
	wire [4-1:0] node23647;
	wire [4-1:0] node23649;
	wire [4-1:0] node23651;
	wire [4-1:0] node23654;
	wire [4-1:0] node23655;
	wire [4-1:0] node23656;
	wire [4-1:0] node23660;
	wire [4-1:0] node23663;
	wire [4-1:0] node23664;
	wire [4-1:0] node23665;
	wire [4-1:0] node23669;
	wire [4-1:0] node23672;
	wire [4-1:0] node23673;
	wire [4-1:0] node23674;
	wire [4-1:0] node23676;
	wire [4-1:0] node23678;
	wire [4-1:0] node23681;
	wire [4-1:0] node23682;
	wire [4-1:0] node23685;
	wire [4-1:0] node23689;
	wire [4-1:0] node23690;
	wire [4-1:0] node23691;
	wire [4-1:0] node23692;
	wire [4-1:0] node23693;
	wire [4-1:0] node23694;
	wire [4-1:0] node23695;
	wire [4-1:0] node23696;
	wire [4-1:0] node23699;
	wire [4-1:0] node23703;
	wire [4-1:0] node23705;
	wire [4-1:0] node23706;
	wire [4-1:0] node23710;
	wire [4-1:0] node23711;
	wire [4-1:0] node23712;
	wire [4-1:0] node23713;
	wire [4-1:0] node23718;
	wire [4-1:0] node23719;
	wire [4-1:0] node23723;
	wire [4-1:0] node23724;
	wire [4-1:0] node23726;
	wire [4-1:0] node23728;
	wire [4-1:0] node23729;
	wire [4-1:0] node23732;
	wire [4-1:0] node23735;
	wire [4-1:0] node23736;
	wire [4-1:0] node23737;
	wire [4-1:0] node23740;
	wire [4-1:0] node23741;
	wire [4-1:0] node23745;
	wire [4-1:0] node23746;
	wire [4-1:0] node23749;
	wire [4-1:0] node23750;
	wire [4-1:0] node23754;
	wire [4-1:0] node23755;
	wire [4-1:0] node23756;
	wire [4-1:0] node23757;
	wire [4-1:0] node23758;
	wire [4-1:0] node23762;
	wire [4-1:0] node23763;
	wire [4-1:0] node23766;
	wire [4-1:0] node23767;
	wire [4-1:0] node23771;
	wire [4-1:0] node23772;
	wire [4-1:0] node23773;
	wire [4-1:0] node23777;
	wire [4-1:0] node23779;
	wire [4-1:0] node23782;
	wire [4-1:0] node23783;
	wire [4-1:0] node23784;
	wire [4-1:0] node23785;
	wire [4-1:0] node23789;
	wire [4-1:0] node23790;
	wire [4-1:0] node23795;
	wire [4-1:0] node23796;
	wire [4-1:0] node23797;
	wire [4-1:0] node23798;
	wire [4-1:0] node23799;
	wire [4-1:0] node23802;
	wire [4-1:0] node23803;
	wire [4-1:0] node23807;
	wire [4-1:0] node23808;
	wire [4-1:0] node23810;
	wire [4-1:0] node23813;
	wire [4-1:0] node23814;
	wire [4-1:0] node23818;
	wire [4-1:0] node23819;
	wire [4-1:0] node23820;
	wire [4-1:0] node23821;
	wire [4-1:0] node23825;
	wire [4-1:0] node23827;
	wire [4-1:0] node23831;
	wire [4-1:0] node23833;
	wire [4-1:0] node23835;
	wire [4-1:0] node23836;
	wire [4-1:0] node23838;
	wire [4-1:0] node23842;
	wire [4-1:0] node23844;
	wire [4-1:0] node23845;
	wire [4-1:0] node23846;
	wire [4-1:0] node23848;
	wire [4-1:0] node23849;
	wire [4-1:0] node23850;
	wire [4-1:0] node23851;
	wire [4-1:0] node23852;
	wire [4-1:0] node23854;
	wire [4-1:0] node23860;
	wire [4-1:0] node23861;
	wire [4-1:0] node23862;
	wire [4-1:0] node23863;
	wire [4-1:0] node23864;
	wire [4-1:0] node23866;
	wire [4-1:0] node23869;
	wire [4-1:0] node23871;
	wire [4-1:0] node23874;
	wire [4-1:0] node23875;
	wire [4-1:0] node23876;
	wire [4-1:0] node23877;
	wire [4-1:0] node23881;
	wire [4-1:0] node23884;
	wire [4-1:0] node23885;
	wire [4-1:0] node23887;
	wire [4-1:0] node23890;
	wire [4-1:0] node23893;
	wire [4-1:0] node23894;
	wire [4-1:0] node23895;
	wire [4-1:0] node23896;
	wire [4-1:0] node23900;
	wire [4-1:0] node23901;
	wire [4-1:0] node23905;
	wire [4-1:0] node23906;
	wire [4-1:0] node23907;
	wire [4-1:0] node23908;
	wire [4-1:0] node23911;
	wire [4-1:0] node23915;
	wire [4-1:0] node23916;
	wire [4-1:0] node23920;
	wire [4-1:0] node23922;
	wire [4-1:0] node23923;
	wire [4-1:0] node23925;
	wire [4-1:0] node23926;
	wire [4-1:0] node23927;
	wire [4-1:0] node23930;
	wire [4-1:0] node23935;
	wire [4-1:0] node23936;
	wire [4-1:0] node23937;
	wire [4-1:0] node23938;
	wire [4-1:0] node23939;
	wire [4-1:0] node23940;
	wire [4-1:0] node23941;
	wire [4-1:0] node23944;
	wire [4-1:0] node23945;
	wire [4-1:0] node23949;
	wire [4-1:0] node23950;
	wire [4-1:0] node23951;
	wire [4-1:0] node23952;
	wire [4-1:0] node23956;
	wire [4-1:0] node23959;
	wire [4-1:0] node23961;
	wire [4-1:0] node23964;
	wire [4-1:0] node23965;
	wire [4-1:0] node23966;
	wire [4-1:0] node23969;
	wire [4-1:0] node23971;
	wire [4-1:0] node23974;
	wire [4-1:0] node23976;
	wire [4-1:0] node23979;
	wire [4-1:0] node23980;
	wire [4-1:0] node23981;
	wire [4-1:0] node23982;
	wire [4-1:0] node23983;
	wire [4-1:0] node23986;
	wire [4-1:0] node23989;
	wire [4-1:0] node23990;
	wire [4-1:0] node23994;
	wire [4-1:0] node23995;
	wire [4-1:0] node23996;
	wire [4-1:0] node23998;
	wire [4-1:0] node24001;
	wire [4-1:0] node24003;
	wire [4-1:0] node24006;
	wire [4-1:0] node24007;
	wire [4-1:0] node24009;
	wire [4-1:0] node24013;
	wire [4-1:0] node24014;
	wire [4-1:0] node24016;
	wire [4-1:0] node24017;
	wire [4-1:0] node24021;
	wire [4-1:0] node24022;
	wire [4-1:0] node24025;
	wire [4-1:0] node24026;
	wire [4-1:0] node24027;
	wire [4-1:0] node24030;
	wire [4-1:0] node24033;
	wire [4-1:0] node24036;
	wire [4-1:0] node24037;
	wire [4-1:0] node24038;
	wire [4-1:0] node24039;
	wire [4-1:0] node24041;
	wire [4-1:0] node24042;
	wire [4-1:0] node24044;
	wire [4-1:0] node24047;
	wire [4-1:0] node24050;
	wire [4-1:0] node24051;
	wire [4-1:0] node24054;
	wire [4-1:0] node24055;
	wire [4-1:0] node24058;
	wire [4-1:0] node24061;
	wire [4-1:0] node24062;
	wire [4-1:0] node24063;
	wire [4-1:0] node24064;
	wire [4-1:0] node24067;
	wire [4-1:0] node24070;
	wire [4-1:0] node24073;
	wire [4-1:0] node24074;
	wire [4-1:0] node24075;
	wire [4-1:0] node24078;
	wire [4-1:0] node24081;
	wire [4-1:0] node24083;
	wire [4-1:0] node24086;
	wire [4-1:0] node24087;
	wire [4-1:0] node24088;
	wire [4-1:0] node24089;
	wire [4-1:0] node24090;
	wire [4-1:0] node24091;
	wire [4-1:0] node24096;
	wire [4-1:0] node24098;
	wire [4-1:0] node24101;
	wire [4-1:0] node24102;
	wire [4-1:0] node24103;
	wire [4-1:0] node24104;
	wire [4-1:0] node24108;
	wire [4-1:0] node24110;
	wire [4-1:0] node24113;
	wire [4-1:0] node24115;
	wire [4-1:0] node24118;
	wire [4-1:0] node24119;
	wire [4-1:0] node24120;
	wire [4-1:0] node24121;
	wire [4-1:0] node24124;
	wire [4-1:0] node24126;
	wire [4-1:0] node24129;
	wire [4-1:0] node24130;
	wire [4-1:0] node24133;
	wire [4-1:0] node24136;
	wire [4-1:0] node24137;
	wire [4-1:0] node24139;
	wire [4-1:0] node24141;
	wire [4-1:0] node24145;
	wire [4-1:0] node24146;
	wire [4-1:0] node24147;
	wire [4-1:0] node24148;
	wire [4-1:0] node24149;
	wire [4-1:0] node24150;
	wire [4-1:0] node24151;
	wire [4-1:0] node24155;
	wire [4-1:0] node24156;
	wire [4-1:0] node24157;
	wire [4-1:0] node24162;
	wire [4-1:0] node24163;
	wire [4-1:0] node24164;
	wire [4-1:0] node24165;
	wire [4-1:0] node24168;
	wire [4-1:0] node24172;
	wire [4-1:0] node24173;
	wire [4-1:0] node24175;
	wire [4-1:0] node24178;
	wire [4-1:0] node24180;
	wire [4-1:0] node24183;
	wire [4-1:0] node24184;
	wire [4-1:0] node24185;
	wire [4-1:0] node24187;
	wire [4-1:0] node24190;
	wire [4-1:0] node24191;
	wire [4-1:0] node24193;
	wire [4-1:0] node24196;
	wire [4-1:0] node24199;
	wire [4-1:0] node24201;
	wire [4-1:0] node24202;
	wire [4-1:0] node24203;
	wire [4-1:0] node24208;
	wire [4-1:0] node24209;
	wire [4-1:0] node24210;
	wire [4-1:0] node24211;
	wire [4-1:0] node24213;
	wire [4-1:0] node24216;
	wire [4-1:0] node24217;
	wire [4-1:0] node24220;
	wire [4-1:0] node24223;
	wire [4-1:0] node24224;
	wire [4-1:0] node24226;
	wire [4-1:0] node24229;
	wire [4-1:0] node24230;
	wire [4-1:0] node24231;
	wire [4-1:0] node24235;
	wire [4-1:0] node24236;
	wire [4-1:0] node24240;
	wire [4-1:0] node24241;
	wire [4-1:0] node24242;
	wire [4-1:0] node24244;
	wire [4-1:0] node24247;
	wire [4-1:0] node24248;
	wire [4-1:0] node24253;
	wire [4-1:0] node24254;
	wire [4-1:0] node24255;
	wire [4-1:0] node24256;
	wire [4-1:0] node24257;
	wire [4-1:0] node24259;
	wire [4-1:0] node24263;
	wire [4-1:0] node24264;
	wire [4-1:0] node24267;
	wire [4-1:0] node24269;
	wire [4-1:0] node24272;
	wire [4-1:0] node24273;
	wire [4-1:0] node24274;
	wire [4-1:0] node24277;
	wire [4-1:0] node24279;
	wire [4-1:0] node24282;
	wire [4-1:0] node24283;
	wire [4-1:0] node24287;
	wire [4-1:0] node24288;
	wire [4-1:0] node24289;
	wire [4-1:0] node24290;
	wire [4-1:0] node24291;
	wire [4-1:0] node24296;
	wire [4-1:0] node24298;
	wire [4-1:0] node24299;
	wire [4-1:0] node24303;
	wire [4-1:0] node24304;
	wire [4-1:0] node24305;
	wire [4-1:0] node24310;
	wire [4-1:0] node24312;
	wire [4-1:0] node24314;
	wire [4-1:0] node24315;
	wire [4-1:0] node24316;
	wire [4-1:0] node24318;
	wire [4-1:0] node24320;
	wire [4-1:0] node24321;
	wire [4-1:0] node24325;
	wire [4-1:0] node24326;
	wire [4-1:0] node24327;
	wire [4-1:0] node24328;
	wire [4-1:0] node24329;
	wire [4-1:0] node24331;
	wire [4-1:0] node24334;
	wire [4-1:0] node24337;
	wire [4-1:0] node24338;
	wire [4-1:0] node24341;
	wire [4-1:0] node24342;
	wire [4-1:0] node24346;
	wire [4-1:0] node24347;
	wire [4-1:0] node24348;
	wire [4-1:0] node24351;
	wire [4-1:0] node24353;
	wire [4-1:0] node24356;
	wire [4-1:0] node24357;
	wire [4-1:0] node24361;
	wire [4-1:0] node24362;
	wire [4-1:0] node24363;
	wire [4-1:0] node24365;
	wire [4-1:0] node24368;
	wire [4-1:0] node24369;
	wire [4-1:0] node24373;
	wire [4-1:0] node24374;
	wire [4-1:0] node24375;
	wire [4-1:0] node24380;
	wire [4-1:0] node24382;
	wire [4-1:0] node24383;
	wire [4-1:0] node24384;
	wire [4-1:0] node24386;
	wire [4-1:0] node24388;
	wire [4-1:0] node24389;

	assign outp = (inp[8]) ? node12354 : node1;
		assign node1 = (inp[9]) ? node6245 : node2;
			assign node2 = (inp[15]) ? node3344 : node3;
				assign node3 = (inp[6]) ? node775 : node4;
					assign node4 = (inp[0]) ? 4'b1101 : node5;
						assign node5 = (inp[2]) ? node475 : node6;
							assign node6 = (inp[1]) ? node242 : node7;
								assign node7 = (inp[14]) ? node91 : node8;
									assign node8 = (inp[13]) ? node54 : node9;
										assign node9 = (inp[12]) ? node23 : node10;
											assign node10 = (inp[3]) ? node18 : node11;
												assign node11 = (inp[7]) ? node13 : 4'b0000;
													assign node13 = (inp[4]) ? 4'b0000 : node14;
														assign node14 = (inp[5]) ? 4'b0100 : 4'b1111;
												assign node18 = (inp[7]) ? node20 : 4'b0100;
													assign node20 = (inp[4]) ? 4'b0100 : 4'b0000;
											assign node23 = (inp[10]) ? node41 : node24;
												assign node24 = (inp[3]) ? node36 : node25;
													assign node25 = (inp[5]) ? node31 : node26;
														assign node26 = (inp[4]) ? node28 : 4'b1111;
															assign node28 = (inp[7]) ? 4'b1111 : 4'b1000;
														assign node31 = (inp[4]) ? node33 : 4'b1100;
															assign node33 = (inp[7]) ? 4'b1100 : 4'b1000;
													assign node36 = (inp[4]) ? node38 : 4'b1000;
														assign node38 = (inp[7]) ? 4'b1000 : 4'b1100;
												assign node41 = (inp[3]) ? node49 : node42;
													assign node42 = (inp[7]) ? node44 : 4'b0000;
														assign node44 = (inp[4]) ? 4'b0000 : node45;
															assign node45 = (inp[5]) ? 4'b0100 : 4'b1111;
													assign node49 = (inp[7]) ? node51 : 4'b0100;
														assign node51 = (inp[4]) ? 4'b0100 : 4'b0000;
										assign node54 = (inp[3]) ? node74 : node55;
											assign node55 = (inp[4]) ? node69 : node56;
												assign node56 = (inp[7]) ? node62 : node57;
													assign node57 = (inp[10]) ? 4'b1000 : node58;
														assign node58 = (inp[12]) ? 4'b0000 : 4'b1000;
													assign node62 = (inp[5]) ? node64 : 4'b1111;
														assign node64 = (inp[10]) ? 4'b1100 : node65;
															assign node65 = (inp[12]) ? 4'b0100 : 4'b1100;
												assign node69 = (inp[12]) ? node71 : 4'b1000;
													assign node71 = (inp[10]) ? 4'b1000 : 4'b0000;
											assign node74 = (inp[7]) ? node80 : node75;
												assign node75 = (inp[10]) ? 4'b1100 : node76;
													assign node76 = (inp[12]) ? 4'b0100 : 4'b1100;
												assign node80 = (inp[4]) ? node86 : node81;
													assign node81 = (inp[12]) ? node83 : 4'b1000;
														assign node83 = (inp[10]) ? 4'b1000 : 4'b0000;
													assign node86 = (inp[10]) ? 4'b1100 : node87;
														assign node87 = (inp[12]) ? 4'b0100 : 4'b1100;
									assign node91 = (inp[11]) ? node161 : node92;
										assign node92 = (inp[13]) ? node130 : node93;
											assign node93 = (inp[12]) ? node117 : node94;
												assign node94 = (inp[10]) ? node104 : node95;
													assign node95 = (inp[3]) ? 4'b1001 : node96;
														assign node96 = (inp[4]) ? node100 : node97;
															assign node97 = (inp[5]) ? 4'b1101 : 4'b1111;
															assign node100 = (inp[7]) ? 4'b1111 : 4'b1001;
													assign node104 = (inp[3]) ? node112 : node105;
														assign node105 = (inp[7]) ? node107 : 4'b0001;
															assign node107 = (inp[4]) ? 4'b0001 : node108;
																assign node108 = (inp[5]) ? 4'b0101 : 4'b1111;
														assign node112 = (inp[4]) ? 4'b0101 : node113;
															assign node113 = (inp[7]) ? 4'b0001 : 4'b0101;
												assign node117 = (inp[3]) ? node125 : node118;
													assign node118 = (inp[5]) ? node120 : 4'b1111;
														assign node120 = (inp[4]) ? node122 : 4'b1101;
															assign node122 = (inp[7]) ? 4'b1101 : 4'b1001;
													assign node125 = (inp[4]) ? node127 : 4'b1001;
														assign node127 = (inp[7]) ? 4'b1001 : 4'b1101;
											assign node130 = (inp[3]) ? node144 : node131;
												assign node131 = (inp[7]) ? node137 : node132;
													assign node132 = (inp[10]) ? node134 : 4'b0001;
														assign node134 = (inp[12]) ? 4'b0001 : 4'b1001;
													assign node137 = (inp[4]) ? node141 : node138;
														assign node138 = (inp[5]) ? 4'b0101 : 4'b1111;
														assign node141 = (inp[10]) ? 4'b1001 : 4'b0001;
												assign node144 = (inp[12]) ? node156 : node145;
													assign node145 = (inp[10]) ? node151 : node146;
														assign node146 = (inp[4]) ? 4'b0101 : node147;
															assign node147 = (inp[7]) ? 4'b0001 : 4'b0101;
														assign node151 = (inp[7]) ? node153 : 4'b1101;
															assign node153 = (inp[4]) ? 4'b1101 : 4'b1001;
													assign node156 = (inp[4]) ? 4'b0101 : node157;
														assign node157 = (inp[7]) ? 4'b0001 : 4'b0101;
										assign node161 = (inp[13]) ? node203 : node162;
											assign node162 = (inp[12]) ? node176 : node163;
												assign node163 = (inp[3]) ? node171 : node164;
													assign node164 = (inp[4]) ? 4'b0000 : node165;
														assign node165 = (inp[7]) ? node167 : 4'b0000;
															assign node167 = (inp[5]) ? 4'b0100 : 4'b1111;
													assign node171 = (inp[4]) ? 4'b0100 : node172;
														assign node172 = (inp[7]) ? 4'b0000 : 4'b0100;
												assign node176 = (inp[10]) ? node190 : node177;
													assign node177 = (inp[3]) ? node185 : node178;
														assign node178 = (inp[5]) ? node180 : 4'b1111;
															assign node180 = (inp[7]) ? 4'b1100 : node181;
																assign node181 = (inp[4]) ? 4'b1000 : 4'b1100;
														assign node185 = (inp[7]) ? 4'b1000 : node186;
															assign node186 = (inp[4]) ? 4'b1100 : 4'b1000;
													assign node190 = (inp[7]) ? node194 : node191;
														assign node191 = (inp[3]) ? 4'b0100 : 4'b0000;
														assign node194 = (inp[3]) ? node200 : node195;
															assign node195 = (inp[4]) ? 4'b0000 : node196;
																assign node196 = (inp[5]) ? 4'b0100 : 4'b1111;
															assign node200 = (inp[4]) ? 4'b0100 : 4'b0000;
											assign node203 = (inp[10]) ? node229 : node204;
												assign node204 = (inp[12]) ? node216 : node205;
													assign node205 = (inp[3]) ? node213 : node206;
														assign node206 = (inp[7]) ? node208 : 4'b1000;
															assign node208 = (inp[4]) ? 4'b1000 : node209;
																assign node209 = (inp[5]) ? 4'b1100 : 4'b1111;
														assign node213 = (inp[7]) ? 4'b1000 : 4'b1100;
													assign node216 = (inp[3]) ? node224 : node217;
														assign node217 = (inp[4]) ? 4'b0000 : node218;
															assign node218 = (inp[7]) ? node220 : 4'b0000;
																assign node220 = (inp[5]) ? 4'b0100 : 4'b1111;
														assign node224 = (inp[7]) ? node226 : 4'b0100;
															assign node226 = (inp[4]) ? 4'b0100 : 4'b0000;
												assign node229 = (inp[3]) ? node237 : node230;
													assign node230 = (inp[7]) ? node232 : 4'b1000;
														assign node232 = (inp[4]) ? 4'b1000 : node233;
															assign node233 = (inp[5]) ? 4'b1100 : 4'b1111;
													assign node237 = (inp[4]) ? 4'b1100 : node238;
														assign node238 = (inp[7]) ? 4'b1000 : 4'b1100;
								assign node242 = (inp[14]) ? node324 : node243;
									assign node243 = (inp[13]) ? node287 : node244;
										assign node244 = (inp[10]) ? node274 : node245;
											assign node245 = (inp[12]) ? node257 : node246;
												assign node246 = (inp[3]) ? node252 : node247;
													assign node247 = (inp[4]) ? 4'b0001 : node248;
														assign node248 = (inp[5]) ? 4'b0101 : 4'b0001;
													assign node252 = (inp[4]) ? 4'b0101 : node253;
														assign node253 = (inp[7]) ? 4'b0001 : 4'b0101;
												assign node257 = (inp[3]) ? node269 : node258;
													assign node258 = (inp[5]) ? node264 : node259;
														assign node259 = (inp[4]) ? node261 : 4'b1111;
															assign node261 = (inp[7]) ? 4'b1111 : 4'b1001;
														assign node264 = (inp[7]) ? 4'b1101 : node265;
															assign node265 = (inp[4]) ? 4'b1001 : 4'b1101;
													assign node269 = (inp[7]) ? 4'b1001 : node270;
														assign node270 = (inp[4]) ? 4'b1101 : 4'b1001;
											assign node274 = (inp[3]) ? node282 : node275;
												assign node275 = (inp[7]) ? node277 : 4'b0001;
													assign node277 = (inp[4]) ? 4'b0001 : node278;
														assign node278 = (inp[5]) ? 4'b0101 : 4'b1111;
												assign node282 = (inp[4]) ? 4'b0101 : node283;
													assign node283 = (inp[7]) ? 4'b0001 : 4'b0101;
										assign node287 = (inp[3]) ? node307 : node288;
											assign node288 = (inp[4]) ? node302 : node289;
												assign node289 = (inp[7]) ? node295 : node290;
													assign node290 = (inp[12]) ? node292 : 4'b1001;
														assign node292 = (inp[10]) ? 4'b1001 : 4'b0001;
													assign node295 = (inp[5]) ? node297 : 4'b1111;
														assign node297 = (inp[10]) ? 4'b1101 : node298;
															assign node298 = (inp[11]) ? 4'b0101 : 4'b1101;
												assign node302 = (inp[12]) ? node304 : 4'b1001;
													assign node304 = (inp[10]) ? 4'b1001 : 4'b0001;
											assign node307 = (inp[10]) ? node319 : node308;
												assign node308 = (inp[12]) ? node314 : node309;
													assign node309 = (inp[7]) ? node311 : 4'b1101;
														assign node311 = (inp[4]) ? 4'b1101 : 4'b1001;
													assign node314 = (inp[4]) ? 4'b0101 : node315;
														assign node315 = (inp[7]) ? 4'b0001 : 4'b0101;
												assign node319 = (inp[4]) ? 4'b1101 : node320;
													assign node320 = (inp[7]) ? 4'b1001 : 4'b1101;
									assign node324 = (inp[11]) ? node400 : node325;
										assign node325 = (inp[13]) ? node367 : node326;
											assign node326 = (inp[10]) ? node354 : node327;
												assign node327 = (inp[12]) ? node337 : node328;
													assign node328 = (inp[5]) ? node330 : 4'b0100;
														assign node330 = (inp[7]) ? node332 : 4'b0000;
															assign node332 = (inp[4]) ? 4'b0100 : node333;
																assign node333 = (inp[3]) ? 4'b0000 : 4'b0100;
													assign node337 = (inp[3]) ? node349 : node338;
														assign node338 = (inp[5]) ? node344 : node339;
															assign node339 = (inp[7]) ? 4'b1111 : node340;
																assign node340 = (inp[4]) ? 4'b1000 : 4'b1111;
															assign node344 = (inp[7]) ? 4'b1100 : node345;
																assign node345 = (inp[4]) ? 4'b1000 : 4'b1100;
														assign node349 = (inp[4]) ? node351 : 4'b1000;
															assign node351 = (inp[7]) ? 4'b1000 : 4'b1100;
												assign node354 = (inp[3]) ? node362 : node355;
													assign node355 = (inp[7]) ? node357 : 4'b0000;
														assign node357 = (inp[4]) ? 4'b0000 : node358;
															assign node358 = (inp[5]) ? 4'b0100 : 4'b1111;
													assign node362 = (inp[4]) ? 4'b0100 : node363;
														assign node363 = (inp[7]) ? 4'b0000 : 4'b0100;
											assign node367 = (inp[3]) ? node383 : node368;
												assign node368 = (inp[4]) ? node378 : node369;
													assign node369 = (inp[7]) ? node375 : node370;
														assign node370 = (inp[12]) ? node372 : 4'b1000;
															assign node372 = (inp[10]) ? 4'b1000 : 4'b0000;
														assign node375 = (inp[5]) ? 4'b1100 : 4'b1111;
													assign node378 = (inp[12]) ? node380 : 4'b1000;
														assign node380 = (inp[10]) ? 4'b1000 : 4'b0000;
												assign node383 = (inp[7]) ? node389 : node384;
													assign node384 = (inp[10]) ? 4'b1100 : node385;
														assign node385 = (inp[12]) ? 4'b0100 : 4'b1100;
													assign node389 = (inp[4]) ? node395 : node390;
														assign node390 = (inp[10]) ? 4'b1000 : node391;
															assign node391 = (inp[12]) ? 4'b0000 : 4'b1000;
														assign node395 = (inp[10]) ? 4'b1100 : node396;
															assign node396 = (inp[12]) ? 4'b0100 : 4'b1100;
										assign node400 = (inp[3]) ? node442 : node401;
											assign node401 = (inp[4]) ? node427 : node402;
												assign node402 = (inp[7]) ? node416 : node403;
													assign node403 = (inp[13]) ? node411 : node404;
														assign node404 = (inp[12]) ? node406 : 4'b0001;
															assign node406 = (inp[10]) ? 4'b0001 : node407;
																assign node407 = (inp[5]) ? 4'b1101 : 4'b1111;
														assign node411 = (inp[12]) ? node413 : 4'b1001;
															assign node413 = (inp[10]) ? 4'b1001 : 4'b0001;
													assign node416 = (inp[5]) ? node418 : 4'b1111;
														assign node418 = (inp[10]) ? node424 : node419;
															assign node419 = (inp[12]) ? node421 : 4'b1101;
																assign node421 = (inp[13]) ? 4'b0101 : 4'b1101;
															assign node424 = (inp[13]) ? 4'b1101 : 4'b0101;
												assign node427 = (inp[13]) ? node437 : node428;
													assign node428 = (inp[10]) ? 4'b0001 : node429;
														assign node429 = (inp[12]) ? node431 : 4'b0001;
															assign node431 = (inp[7]) ? node433 : 4'b1001;
																assign node433 = (inp[5]) ? 4'b1101 : 4'b1111;
													assign node437 = (inp[10]) ? 4'b1001 : node438;
														assign node438 = (inp[12]) ? 4'b0001 : 4'b1001;
											assign node442 = (inp[7]) ? node456 : node443;
												assign node443 = (inp[13]) ? node451 : node444;
													assign node444 = (inp[12]) ? node446 : 4'b0101;
														assign node446 = (inp[10]) ? 4'b0101 : node447;
															assign node447 = (inp[4]) ? 4'b1101 : 4'b1001;
													assign node451 = (inp[10]) ? 4'b1101 : node452;
														assign node452 = (inp[12]) ? 4'b0101 : 4'b1101;
												assign node456 = (inp[4]) ? node466 : node457;
													assign node457 = (inp[12]) ? node459 : 4'b0001;
														assign node459 = (inp[10]) ? node463 : node460;
															assign node460 = (inp[13]) ? 4'b0001 : 4'b1001;
															assign node463 = (inp[13]) ? 4'b1001 : 4'b0001;
													assign node466 = (inp[10]) ? node472 : node467;
														assign node467 = (inp[13]) ? node469 : 4'b1001;
															assign node469 = (inp[12]) ? 4'b0101 : 4'b1101;
														assign node472 = (inp[13]) ? 4'b1101 : 4'b0101;
							assign node475 = (inp[5]) ? node477 : 4'b1111;
								assign node477 = (inp[3]) ? node595 : node478;
									assign node478 = (inp[4]) ? node526 : node479;
										assign node479 = (inp[7]) ? 4'b1111 : node480;
											assign node480 = (inp[13]) ? node502 : node481;
												assign node481 = (inp[10]) ? node491 : node482;
													assign node482 = (inp[12]) ? 4'b1111 : node483;
														assign node483 = (inp[14]) ? node487 : node484;
															assign node484 = (inp[1]) ? 4'b0001 : 4'b0000;
															assign node487 = (inp[11]) ? 4'b0000 : 4'b1111;
													assign node491 = (inp[1]) ? node497 : node492;
														assign node492 = (inp[12]) ? 4'b0000 : node493;
															assign node493 = (inp[11]) ? 4'b0000 : 4'b0001;
														assign node497 = (inp[11]) ? 4'b0001 : node498;
															assign node498 = (inp[14]) ? 4'b0000 : 4'b0001;
												assign node502 = (inp[10]) ? node516 : node503;
													assign node503 = (inp[12]) ? node509 : node504;
														assign node504 = (inp[1]) ? node506 : 4'b1000;
															assign node506 = (inp[14]) ? 4'b1000 : 4'b1001;
														assign node509 = (inp[14]) ? node511 : 4'b0000;
															assign node511 = (inp[1]) ? node513 : 4'b0001;
																assign node513 = (inp[11]) ? 4'b0001 : 4'b0000;
													assign node516 = (inp[1]) ? node520 : node517;
														assign node517 = (inp[11]) ? 4'b1000 : 4'b1001;
														assign node520 = (inp[11]) ? 4'b1001 : node521;
															assign node521 = (inp[14]) ? 4'b1000 : 4'b1001;
										assign node526 = (inp[1]) ? node568 : node527;
											assign node527 = (inp[11]) ? node555 : node528;
												assign node528 = (inp[14]) ? node542 : node529;
													assign node529 = (inp[12]) ? node533 : node530;
														assign node530 = (inp[13]) ? 4'b1000 : 4'b0000;
														assign node533 = (inp[7]) ? node539 : node534;
															assign node534 = (inp[13]) ? 4'b0000 : node535;
																assign node535 = (inp[10]) ? 4'b0000 : 4'b1000;
															assign node539 = (inp[13]) ? 4'b0000 : 4'b1111;
													assign node542 = (inp[13]) ? node550 : node543;
														assign node543 = (inp[10]) ? node547 : node544;
															assign node544 = (inp[7]) ? 4'b1111 : 4'b1001;
															assign node547 = (inp[12]) ? 4'b1001 : 4'b0001;
														assign node550 = (inp[10]) ? node552 : 4'b0001;
															assign node552 = (inp[12]) ? 4'b0001 : 4'b1001;
												assign node555 = (inp[13]) ? node563 : node556;
													assign node556 = (inp[12]) ? node558 : 4'b0000;
														assign node558 = (inp[10]) ? 4'b0000 : node559;
															assign node559 = (inp[7]) ? 4'b1111 : 4'b1000;
													assign node563 = (inp[10]) ? 4'b1000 : node564;
														assign node564 = (inp[12]) ? 4'b0000 : 4'b1000;
											assign node568 = (inp[13]) ? node582 : node569;
												assign node569 = (inp[10]) ? node577 : node570;
													assign node570 = (inp[12]) ? node574 : node571;
														assign node571 = (inp[11]) ? 4'b0001 : 4'b0000;
														assign node574 = (inp[7]) ? 4'b1111 : 4'b1001;
													assign node577 = (inp[14]) ? node579 : 4'b0001;
														assign node579 = (inp[11]) ? 4'b0001 : 4'b0000;
												assign node582 = (inp[10]) ? node590 : node583;
													assign node583 = (inp[12]) ? node585 : 4'b1001;
														assign node585 = (inp[14]) ? node587 : 4'b0001;
															assign node587 = (inp[11]) ? 4'b0001 : 4'b0000;
													assign node590 = (inp[11]) ? 4'b1001 : node591;
														assign node591 = (inp[14]) ? 4'b1000 : 4'b1001;
									assign node595 = (inp[4]) ? node705 : node596;
										assign node596 = (inp[7]) ? node650 : node597;
											assign node597 = (inp[1]) ? node625 : node598;
												assign node598 = (inp[11]) ? node616 : node599;
													assign node599 = (inp[14]) ? node609 : node600;
														assign node600 = (inp[10]) ? 4'b0100 : node601;
															assign node601 = (inp[13]) ? node605 : node602;
																assign node602 = (inp[12]) ? 4'b1000 : 4'b0100;
																assign node605 = (inp[12]) ? 4'b0100 : 4'b1100;
														assign node609 = (inp[13]) ? 4'b0101 : node610;
															assign node610 = (inp[10]) ? node612 : 4'b1001;
																assign node612 = (inp[12]) ? 4'b1001 : 4'b0101;
													assign node616 = (inp[12]) ? node620 : node617;
														assign node617 = (inp[13]) ? 4'b1100 : 4'b0100;
														assign node620 = (inp[10]) ? 4'b0100 : node621;
															assign node621 = (inp[13]) ? 4'b0100 : 4'b1000;
												assign node625 = (inp[11]) ? node639 : node626;
													assign node626 = (inp[14]) ? node632 : node627;
														assign node627 = (inp[13]) ? node629 : 4'b0101;
															assign node629 = (inp[10]) ? 4'b1101 : 4'b0101;
														assign node632 = (inp[12]) ? node636 : node633;
															assign node633 = (inp[13]) ? 4'b1100 : 4'b0100;
															assign node636 = (inp[13]) ? 4'b0100 : 4'b1000;
													assign node639 = (inp[13]) ? node645 : node640;
														assign node640 = (inp[10]) ? 4'b0101 : node641;
															assign node641 = (inp[12]) ? 4'b1001 : 4'b0101;
														assign node645 = (inp[12]) ? node647 : 4'b1101;
															assign node647 = (inp[10]) ? 4'b1101 : 4'b0101;
											assign node650 = (inp[1]) ? node676 : node651;
												assign node651 = (inp[11]) ? node667 : node652;
													assign node652 = (inp[14]) ? node660 : node653;
														assign node653 = (inp[12]) ? node655 : 4'b0000;
															assign node655 = (inp[10]) ? 4'b0000 : node656;
																assign node656 = (inp[13]) ? 4'b0000 : 4'b1000;
														assign node660 = (inp[13]) ? 4'b0001 : node661;
															assign node661 = (inp[12]) ? 4'b1001 : node662;
																assign node662 = (inp[10]) ? 4'b0001 : 4'b1001;
													assign node667 = (inp[13]) ? node673 : node668;
														assign node668 = (inp[12]) ? node670 : 4'b0000;
															assign node670 = (inp[10]) ? 4'b0000 : 4'b1000;
														assign node673 = (inp[12]) ? 4'b0000 : 4'b1000;
												assign node676 = (inp[14]) ? node688 : node677;
													assign node677 = (inp[13]) ? node683 : node678;
														assign node678 = (inp[10]) ? 4'b0001 : node679;
															assign node679 = (inp[12]) ? 4'b1001 : 4'b0001;
														assign node683 = (inp[10]) ? 4'b1001 : node684;
															assign node684 = (inp[12]) ? 4'b0001 : 4'b1001;
													assign node688 = (inp[11]) ? node700 : node689;
														assign node689 = (inp[13]) ? node695 : node690;
															assign node690 = (inp[12]) ? node692 : 4'b0000;
																assign node692 = (inp[10]) ? 4'b0000 : 4'b1000;
															assign node695 = (inp[10]) ? 4'b1000 : node696;
																assign node696 = (inp[12]) ? 4'b0000 : 4'b1000;
														assign node700 = (inp[13]) ? 4'b1001 : node701;
															assign node701 = (inp[12]) ? 4'b1001 : 4'b0001;
										assign node705 = (inp[1]) ? node747 : node706;
											assign node706 = (inp[11]) ? node734 : node707;
												assign node707 = (inp[14]) ? node721 : node708;
													assign node708 = (inp[13]) ? node716 : node709;
														assign node709 = (inp[10]) ? 4'b0100 : node710;
															assign node710 = (inp[7]) ? 4'b1000 : node711;
																assign node711 = (inp[12]) ? 4'b1100 : 4'b0100;
														assign node716 = (inp[10]) ? 4'b1100 : node717;
															assign node717 = (inp[12]) ? 4'b0100 : 4'b1100;
													assign node721 = (inp[13]) ? node729 : node722;
														assign node722 = (inp[12]) ? node726 : node723;
															assign node723 = (inp[10]) ? 4'b0101 : 4'b1101;
															assign node726 = (inp[7]) ? 4'b1001 : 4'b1101;
														assign node729 = (inp[10]) ? node731 : 4'b0101;
															assign node731 = (inp[12]) ? 4'b0101 : 4'b1101;
												assign node734 = (inp[13]) ? node742 : node735;
													assign node735 = (inp[10]) ? 4'b0100 : node736;
														assign node736 = (inp[12]) ? node738 : 4'b0100;
															assign node738 = (inp[7]) ? 4'b1000 : 4'b1100;
													assign node742 = (inp[10]) ? 4'b1100 : node743;
														assign node743 = (inp[12]) ? 4'b0100 : 4'b1100;
											assign node747 = (inp[13]) ? node763 : node748;
												assign node748 = (inp[10]) ? 4'b0101 : node749;
													assign node749 = (inp[12]) ? node755 : node750;
														assign node750 = (inp[11]) ? 4'b0101 : node751;
															assign node751 = (inp[14]) ? 4'b0100 : 4'b0101;
														assign node755 = (inp[7]) ? node757 : 4'b1101;
															assign node757 = (inp[14]) ? node759 : 4'b1001;
																assign node759 = (inp[11]) ? 4'b1001 : 4'b1000;
												assign node763 = (inp[10]) ? node769 : node764;
													assign node764 = (inp[12]) ? 4'b0101 : node765;
														assign node765 = (inp[14]) ? 4'b1100 : 4'b1101;
													assign node769 = (inp[14]) ? node771 : 4'b1101;
														assign node771 = (inp[11]) ? 4'b1101 : 4'b1100;
					assign node775 = (inp[5]) ? node1841 : node776;
						assign node776 = (inp[0]) ? node1530 : node777;
							assign node777 = (inp[11]) ? node1207 : node778;
								assign node778 = (inp[10]) ? node1004 : node779;
									assign node779 = (inp[12]) ? node885 : node780;
										assign node780 = (inp[4]) ? node826 : node781;
											assign node781 = (inp[7]) ? node797 : node782;
												assign node782 = (inp[3]) ? 4'b0000 : node783;
													assign node783 = (inp[2]) ? node785 : 4'b0000;
														assign node785 = (inp[13]) ? node789 : node786;
															assign node786 = (inp[1]) ? 4'b0001 : 4'b0000;
															assign node789 = (inp[1]) ? node793 : node790;
																assign node790 = (inp[14]) ? 4'b0001 : 4'b1000;
																assign node793 = (inp[14]) ? 4'b1000 : 4'b1001;
												assign node797 = (inp[13]) ? node817 : node798;
													assign node798 = (inp[2]) ? node804 : node799;
														assign node799 = (inp[1]) ? node801 : 4'b0100;
															assign node801 = (inp[14]) ? 4'b0100 : 4'b0101;
														assign node804 = (inp[3]) ? node810 : node805;
															assign node805 = (inp[14]) ? 4'b0100 : node806;
																assign node806 = (inp[1]) ? 4'b0101 : 4'b0100;
															assign node810 = (inp[1]) ? node814 : node811;
																assign node811 = (inp[14]) ? 4'b1001 : 4'b0000;
																assign node814 = (inp[14]) ? 4'b0000 : 4'b0001;
													assign node817 = (inp[2]) ? node819 : 4'b0000;
														assign node819 = (inp[3]) ? 4'b0000 : node820;
															assign node820 = (inp[1]) ? 4'b1100 : node821;
																assign node821 = (inp[14]) ? 4'b0101 : 4'b1100;
											assign node826 = (inp[13]) ? node858 : node827;
												assign node827 = (inp[7]) ? node841 : node828;
													assign node828 = (inp[3]) ? node834 : node829;
														assign node829 = (inp[2]) ? node831 : 4'b0100;
															assign node831 = (inp[14]) ? 4'b1001 : 4'b0001;
														assign node834 = (inp[2]) ? 4'b0100 : node835;
															assign node835 = (inp[1]) ? 4'b1000 : node836;
																assign node836 = (inp[14]) ? 4'b0000 : 4'b0001;
													assign node841 = (inp[1]) ? node849 : node842;
														assign node842 = (inp[2]) ? node846 : node843;
															assign node843 = (inp[14]) ? 4'b0000 : 4'b0001;
															assign node846 = (inp[3]) ? 4'b0000 : 4'b1101;
														assign node849 = (inp[2]) ? node853 : node850;
															assign node850 = (inp[3]) ? 4'b1000 : 4'b0000;
															assign node853 = (inp[14]) ? 4'b0000 : node854;
																assign node854 = (inp[3]) ? 4'b0000 : 4'b0001;
												assign node858 = (inp[2]) ? node876 : node859;
													assign node859 = (inp[3]) ? node861 : 4'b0100;
														assign node861 = (inp[7]) ? node869 : node862;
															assign node862 = (inp[1]) ? node866 : node863;
																assign node863 = (inp[14]) ? 4'b1100 : 4'b1101;
																assign node866 = (inp[14]) ? 4'b1101 : 4'b0100;
															assign node869 = (inp[1]) ? node873 : node870;
																assign node870 = (inp[14]) ? 4'b1000 : 4'b1001;
																assign node873 = (inp[14]) ? 4'b1001 : 4'b0100;
													assign node876 = (inp[3]) ? 4'b0100 : node877;
														assign node877 = (inp[1]) ? node881 : node878;
															assign node878 = (inp[14]) ? 4'b0001 : 4'b1000;
															assign node881 = (inp[14]) ? 4'b1000 : 4'b1001;
										assign node885 = (inp[1]) ? node949 : node886;
											assign node886 = (inp[14]) ? node916 : node887;
												assign node887 = (inp[13]) ? node893 : node888;
													assign node888 = (inp[4]) ? 4'b1000 : node889;
														assign node889 = (inp[2]) ? 4'b1000 : 4'b1100;
													assign node893 = (inp[2]) ? node905 : node894;
														assign node894 = (inp[4]) ? node900 : node895;
															assign node895 = (inp[7]) ? node897 : 4'b1000;
																assign node897 = (inp[3]) ? 4'b1100 : 4'b0100;
															assign node900 = (inp[3]) ? 4'b0101 : node901;
																assign node901 = (inp[7]) ? 4'b1000 : 4'b1100;
														assign node905 = (inp[3]) ? node911 : node906;
															assign node906 = (inp[4]) ? 4'b0000 : node907;
																assign node907 = (inp[7]) ? 4'b0100 : 4'b0000;
															assign node911 = (inp[4]) ? 4'b1100 : node912;
																assign node912 = (inp[7]) ? 4'b0000 : 4'b1000;
												assign node916 = (inp[3]) ? node940 : node917;
													assign node917 = (inp[2]) ? node931 : node918;
														assign node918 = (inp[4]) ? node926 : node919;
															assign node919 = (inp[7]) ? node923 : node920;
																assign node920 = (inp[13]) ? 4'b1000 : 4'b1101;
																assign node923 = (inp[13]) ? 4'b0101 : 4'b1101;
															assign node926 = (inp[7]) ? 4'b1000 : node927;
																assign node927 = (inp[13]) ? 4'b1100 : 4'b1000;
														assign node931 = (inp[13]) ? node935 : node932;
															assign node932 = (inp[4]) ? 4'b1001 : 4'b1101;
															assign node935 = (inp[7]) ? node937 : 4'b0001;
																assign node937 = (inp[4]) ? 4'b0001 : 4'b0101;
													assign node940 = (inp[13]) ? node944 : node941;
														assign node941 = (inp[4]) ? 4'b1000 : 4'b1001;
														assign node944 = (inp[4]) ? node946 : 4'b1000;
															assign node946 = (inp[7]) ? 4'b1000 : 4'b1100;
											assign node949 = (inp[3]) ? node977 : node950;
												assign node950 = (inp[13]) ? node968 : node951;
													assign node951 = (inp[2]) ? node961 : node952;
														assign node952 = (inp[7]) ? node956 : node953;
															assign node953 = (inp[4]) ? 4'b0100 : 4'b0000;
															assign node956 = (inp[4]) ? 4'b0000 : node957;
																assign node957 = (inp[14]) ? 4'b1100 : 4'b1101;
														assign node961 = (inp[14]) ? 4'b1100 : node962;
															assign node962 = (inp[7]) ? 4'b1101 : node963;
																assign node963 = (inp[4]) ? 4'b1001 : 4'b1101;
													assign node968 = (inp[4]) ? node974 : node969;
														assign node969 = (inp[2]) ? node971 : 4'b0000;
															assign node971 = (inp[7]) ? 4'b0100 : 4'b0000;
														assign node974 = (inp[2]) ? 4'b0001 : 4'b0100;
												assign node977 = (inp[4]) ? node989 : node978;
													assign node978 = (inp[13]) ? 4'b0000 : node979;
														assign node979 = (inp[2]) ? node983 : node980;
															assign node980 = (inp[7]) ? 4'b0100 : 4'b0000;
															assign node983 = (inp[14]) ? node985 : 4'b1001;
																assign node985 = (inp[7]) ? 4'b1000 : 4'b0000;
													assign node989 = (inp[13]) ? node999 : node990;
														assign node990 = (inp[14]) ? node996 : node991;
															assign node991 = (inp[7]) ? 4'b0000 : node992;
																assign node992 = (inp[2]) ? 4'b0100 : 4'b0000;
															assign node996 = (inp[7]) ? 4'b0000 : 4'b0001;
														assign node999 = (inp[2]) ? 4'b0100 : node1000;
															assign node1000 = (inp[14]) ? 4'b1101 : 4'b1000;
									assign node1004 = (inp[4]) ? node1096 : node1005;
										assign node1005 = (inp[7]) ? node1051 : node1006;
											assign node1006 = (inp[1]) ? node1032 : node1007;
												assign node1007 = (inp[12]) ? node1019 : node1008;
													assign node1008 = (inp[3]) ? node1014 : node1009;
														assign node1009 = (inp[13]) ? 4'b1000 : node1010;
															assign node1010 = (inp[14]) ? 4'b0001 : 4'b0000;
														assign node1014 = (inp[13]) ? node1016 : 4'b1000;
															assign node1016 = (inp[2]) ? 4'b1000 : 4'b0001;
													assign node1019 = (inp[2]) ? node1025 : node1020;
														assign node1020 = (inp[3]) ? node1022 : 4'b0000;
															assign node1022 = (inp[14]) ? 4'b0000 : 4'b0001;
														assign node1025 = (inp[3]) ? 4'b0000 : node1026;
															assign node1026 = (inp[14]) ? 4'b1101 : node1027;
																assign node1027 = (inp[13]) ? 4'b1000 : 4'b0000;
												assign node1032 = (inp[3]) ? node1042 : node1033;
													assign node1033 = (inp[2]) ? node1035 : 4'b1000;
														assign node1035 = (inp[14]) ? node1039 : node1036;
															assign node1036 = (inp[13]) ? 4'b1001 : 4'b0001;
															assign node1039 = (inp[13]) ? 4'b1000 : 4'b0000;
													assign node1042 = (inp[2]) ? 4'b1000 : node1043;
														assign node1043 = (inp[14]) ? node1045 : 4'b1000;
															assign node1045 = (inp[12]) ? 4'b0001 : node1046;
																assign node1046 = (inp[13]) ? 4'b1001 : 4'b1000;
											assign node1051 = (inp[13]) ? node1077 : node1052;
												assign node1052 = (inp[3]) ? node1062 : node1053;
													assign node1053 = (inp[1]) ? node1059 : node1054;
														assign node1054 = (inp[14]) ? node1056 : 4'b0100;
															assign node1056 = (inp[12]) ? 4'b1101 : 4'b0101;
														assign node1059 = (inp[14]) ? 4'b0100 : 4'b0101;
													assign node1062 = (inp[2]) ? node1068 : node1063;
														assign node1063 = (inp[1]) ? 4'b1100 : node1064;
															assign node1064 = (inp[14]) ? 4'b0100 : 4'b1100;
														assign node1068 = (inp[1]) ? node1074 : node1069;
															assign node1069 = (inp[14]) ? node1071 : 4'b0000;
																assign node1071 = (inp[12]) ? 4'b1001 : 4'b0001;
															assign node1074 = (inp[14]) ? 4'b0000 : 4'b0001;
												assign node1077 = (inp[1]) ? node1089 : node1078;
													assign node1078 = (inp[12]) ? node1084 : node1079;
														assign node1079 = (inp[3]) ? 4'b1000 : node1080;
															assign node1080 = (inp[14]) ? 4'b1101 : 4'b1100;
														assign node1084 = (inp[3]) ? 4'b0000 : node1085;
															assign node1085 = (inp[2]) ? 4'b0101 : 4'b0000;
													assign node1089 = (inp[2]) ? node1091 : 4'b1000;
														assign node1091 = (inp[3]) ? 4'b1000 : node1092;
															assign node1092 = (inp[14]) ? 4'b1100 : 4'b1101;
										assign node1096 = (inp[13]) ? node1158 : node1097;
											assign node1097 = (inp[7]) ? node1127 : node1098;
												assign node1098 = (inp[3]) ? node1114 : node1099;
													assign node1099 = (inp[2]) ? node1105 : node1100;
														assign node1100 = (inp[12]) ? node1102 : 4'b1100;
															assign node1102 = (inp[1]) ? 4'b1100 : 4'b0100;
														assign node1105 = (inp[14]) ? node1109 : node1106;
															assign node1106 = (inp[1]) ? 4'b0001 : 4'b0000;
															assign node1109 = (inp[1]) ? 4'b0000 : node1110;
																assign node1110 = (inp[12]) ? 4'b1001 : 4'b0001;
													assign node1114 = (inp[2]) ? node1122 : node1115;
														assign node1115 = (inp[1]) ? node1119 : node1116;
															assign node1116 = (inp[14]) ? 4'b1000 : 4'b1001;
															assign node1119 = (inp[14]) ? 4'b1001 : 4'b0100;
														assign node1122 = (inp[1]) ? 4'b1100 : node1123;
															assign node1123 = (inp[12]) ? 4'b0100 : 4'b1100;
												assign node1127 = (inp[3]) ? node1145 : node1128;
													assign node1128 = (inp[2]) ? node1134 : node1129;
														assign node1129 = (inp[1]) ? 4'b1000 : node1130;
															assign node1130 = (inp[12]) ? 4'b0000 : 4'b1000;
														assign node1134 = (inp[12]) ? node1142 : node1135;
															assign node1135 = (inp[1]) ? node1139 : node1136;
																assign node1136 = (inp[14]) ? 4'b0001 : 4'b0000;
																assign node1139 = (inp[14]) ? 4'b0000 : 4'b0001;
															assign node1142 = (inp[14]) ? 4'b1101 : 4'b0000;
													assign node1145 = (inp[2]) ? node1153 : node1146;
														assign node1146 = (inp[1]) ? node1150 : node1147;
															assign node1147 = (inp[14]) ? 4'b1000 : 4'b1001;
															assign node1150 = (inp[14]) ? 4'b0001 : 4'b0000;
														assign node1153 = (inp[12]) ? node1155 : 4'b1000;
															assign node1155 = (inp[1]) ? 4'b1000 : 4'b0000;
											assign node1158 = (inp[3]) ? node1188 : node1159;
												assign node1159 = (inp[2]) ? node1165 : node1160;
													assign node1160 = (inp[1]) ? 4'b1100 : node1161;
														assign node1161 = (inp[12]) ? 4'b0100 : 4'b1100;
													assign node1165 = (inp[7]) ? node1175 : node1166;
														assign node1166 = (inp[14]) ? node1170 : node1167;
															assign node1167 = (inp[1]) ? 4'b1001 : 4'b1000;
															assign node1170 = (inp[1]) ? 4'b1000 : node1171;
																assign node1171 = (inp[12]) ? 4'b0001 : 4'b1001;
														assign node1175 = (inp[12]) ? node1183 : node1176;
															assign node1176 = (inp[14]) ? node1180 : node1177;
																assign node1177 = (inp[1]) ? 4'b1001 : 4'b1000;
																assign node1180 = (inp[1]) ? 4'b1000 : 4'b1001;
															assign node1183 = (inp[14]) ? 4'b1000 : node1184;
																assign node1184 = (inp[1]) ? 4'b1001 : 4'b1000;
												assign node1188 = (inp[12]) ? node1196 : node1189;
													assign node1189 = (inp[2]) ? 4'b1100 : node1190;
														assign node1190 = (inp[1]) ? node1192 : 4'b0100;
															assign node1192 = (inp[14]) ? 4'b1101 : 4'b1100;
													assign node1196 = (inp[1]) ? node1202 : node1197;
														assign node1197 = (inp[2]) ? 4'b0100 : node1198;
															assign node1198 = (inp[7]) ? 4'b0101 : 4'b0100;
														assign node1202 = (inp[2]) ? 4'b1100 : node1203;
															assign node1203 = (inp[14]) ? 4'b0101 : 4'b1100;
								assign node1207 = (inp[1]) ? node1407 : node1208;
									assign node1208 = (inp[2]) ? node1308 : node1209;
										assign node1209 = (inp[3]) ? node1261 : node1210;
											assign node1210 = (inp[4]) ? node1234 : node1211;
												assign node1211 = (inp[7]) ? node1221 : node1212;
													assign node1212 = (inp[12]) ? node1216 : node1213;
														assign node1213 = (inp[10]) ? 4'b1001 : 4'b0001;
														assign node1216 = (inp[10]) ? 4'b0001 : node1217;
															assign node1217 = (inp[14]) ? 4'b1001 : 4'b1100;
													assign node1221 = (inp[13]) ? node1227 : node1222;
														assign node1222 = (inp[10]) ? 4'b0100 : node1223;
															assign node1223 = (inp[12]) ? 4'b1100 : 4'b0100;
														assign node1227 = (inp[10]) ? node1231 : node1228;
															assign node1228 = (inp[12]) ? 4'b0100 : 4'b0001;
															assign node1231 = (inp[12]) ? 4'b0001 : 4'b1001;
												assign node1234 = (inp[7]) ? node1248 : node1235;
													assign node1235 = (inp[13]) ? node1241 : node1236;
														assign node1236 = (inp[12]) ? 4'b1001 : node1237;
															assign node1237 = (inp[10]) ? 4'b1101 : 4'b0101;
														assign node1241 = (inp[10]) ? node1245 : node1242;
															assign node1242 = (inp[12]) ? 4'b1101 : 4'b0101;
															assign node1245 = (inp[12]) ? 4'b0101 : 4'b1101;
													assign node1248 = (inp[13]) ? node1254 : node1249;
														assign node1249 = (inp[10]) ? 4'b1001 : node1250;
															assign node1250 = (inp[12]) ? 4'b1001 : 4'b0001;
														assign node1254 = (inp[12]) ? node1258 : node1255;
															assign node1255 = (inp[10]) ? 4'b1101 : 4'b0101;
															assign node1258 = (inp[10]) ? 4'b0101 : 4'b1001;
											assign node1261 = (inp[4]) ? node1291 : node1262;
												assign node1262 = (inp[13]) ? node1278 : node1263;
													assign node1263 = (inp[7]) ? node1271 : node1264;
														assign node1264 = (inp[10]) ? node1268 : node1265;
															assign node1265 = (inp[12]) ? 4'b1101 : 4'b0001;
															assign node1268 = (inp[12]) ? 4'b0001 : 4'b1001;
														assign node1271 = (inp[12]) ? node1275 : node1272;
															assign node1272 = (inp[10]) ? 4'b1101 : 4'b0101;
															assign node1275 = (inp[10]) ? 4'b0101 : 4'b1101;
													assign node1278 = (inp[10]) ? node1284 : node1279;
														assign node1279 = (inp[12]) ? node1281 : 4'b0001;
															assign node1281 = (inp[7]) ? 4'b1101 : 4'b1001;
														assign node1284 = (inp[12]) ? node1288 : node1285;
															assign node1285 = (inp[7]) ? 4'b1001 : 4'b1000;
															assign node1288 = (inp[7]) ? 4'b0001 : 4'b0000;
												assign node1291 = (inp[13]) ? node1301 : node1292;
													assign node1292 = (inp[12]) ? node1298 : node1293;
														assign node1293 = (inp[7]) ? 4'b0000 : node1294;
															assign node1294 = (inp[10]) ? 4'b0100 : 4'b0000;
														assign node1298 = (inp[10]) ? 4'b1000 : 4'b0000;
													assign node1301 = (inp[10]) ? node1305 : node1302;
														assign node1302 = (inp[7]) ? 4'b1000 : 4'b1100;
														assign node1305 = (inp[12]) ? 4'b0100 : 4'b1100;
										assign node1308 = (inp[3]) ? node1342 : node1309;
											assign node1309 = (inp[7]) ? node1321 : node1310;
												assign node1310 = (inp[13]) ? node1316 : node1311;
													assign node1311 = (inp[10]) ? 4'b0000 : node1312;
														assign node1312 = (inp[12]) ? 4'b1000 : 4'b0000;
													assign node1316 = (inp[10]) ? 4'b1000 : node1317;
														assign node1317 = (inp[12]) ? 4'b0000 : 4'b1000;
												assign node1321 = (inp[4]) ? node1333 : node1322;
													assign node1322 = (inp[12]) ? node1324 : 4'b1100;
														assign node1324 = (inp[14]) ? 4'b0100 : node1325;
															assign node1325 = (inp[13]) ? node1329 : node1326;
																assign node1326 = (inp[10]) ? 4'b0100 : 4'b1100;
																assign node1329 = (inp[10]) ? 4'b1100 : 4'b0100;
													assign node1333 = (inp[10]) ? node1339 : node1334;
														assign node1334 = (inp[13]) ? 4'b0000 : node1335;
															assign node1335 = (inp[12]) ? 4'b1100 : 4'b0000;
														assign node1339 = (inp[13]) ? 4'b1000 : 4'b0000;
											assign node1342 = (inp[4]) ? node1374 : node1343;
												assign node1343 = (inp[7]) ? node1361 : node1344;
													assign node1344 = (inp[13]) ? node1354 : node1345;
														assign node1345 = (inp[14]) ? 4'b0001 : node1346;
															assign node1346 = (inp[10]) ? node1350 : node1347;
																assign node1347 = (inp[12]) ? 4'b1000 : 4'b0001;
																assign node1350 = (inp[12]) ? 4'b0001 : 4'b1001;
														assign node1354 = (inp[10]) ? node1358 : node1355;
															assign node1355 = (inp[12]) ? 4'b1001 : 4'b0001;
															assign node1358 = (inp[12]) ? 4'b0001 : 4'b1001;
													assign node1361 = (inp[13]) ? node1367 : node1362;
														assign node1362 = (inp[10]) ? 4'b0000 : node1363;
															assign node1363 = (inp[12]) ? 4'b1000 : 4'b0000;
														assign node1367 = (inp[12]) ? node1371 : node1368;
															assign node1368 = (inp[10]) ? 4'b1001 : 4'b0001;
															assign node1371 = (inp[10]) ? 4'b0001 : 4'b0000;
												assign node1374 = (inp[7]) ? node1392 : node1375;
													assign node1375 = (inp[13]) ? node1383 : node1376;
														assign node1376 = (inp[10]) ? node1380 : node1377;
															assign node1377 = (inp[12]) ? 4'b1001 : 4'b0101;
															assign node1380 = (inp[12]) ? 4'b0101 : 4'b1101;
														assign node1383 = (inp[14]) ? 4'b0101 : node1384;
															assign node1384 = (inp[12]) ? node1388 : node1385;
																assign node1385 = (inp[10]) ? 4'b1101 : 4'b0101;
																assign node1388 = (inp[10]) ? 4'b0101 : 4'b1101;
													assign node1392 = (inp[13]) ? node1400 : node1393;
														assign node1393 = (inp[12]) ? node1397 : node1394;
															assign node1394 = (inp[10]) ? 4'b1001 : 4'b0001;
															assign node1397 = (inp[10]) ? 4'b0001 : 4'b1001;
														assign node1400 = (inp[12]) ? node1404 : node1401;
															assign node1401 = (inp[10]) ? 4'b1101 : 4'b0101;
															assign node1404 = (inp[10]) ? 4'b0101 : 4'b1001;
									assign node1407 = (inp[10]) ? node1473 : node1408;
										assign node1408 = (inp[4]) ? node1438 : node1409;
											assign node1409 = (inp[7]) ? node1419 : node1410;
												assign node1410 = (inp[3]) ? 4'b0001 : node1411;
													assign node1411 = (inp[2]) ? node1413 : 4'b0001;
														assign node1413 = (inp[13]) ? node1415 : 4'b0001;
															assign node1415 = (inp[14]) ? 4'b0001 : 4'b1001;
												assign node1419 = (inp[3]) ? node1429 : node1420;
													assign node1420 = (inp[13]) ? node1424 : node1421;
														assign node1421 = (inp[12]) ? 4'b1101 : 4'b0101;
														assign node1424 = (inp[2]) ? node1426 : 4'b0001;
															assign node1426 = (inp[12]) ? 4'b0101 : 4'b1101;
													assign node1429 = (inp[2]) ? node1433 : node1430;
														assign node1430 = (inp[13]) ? 4'b0001 : 4'b0101;
														assign node1433 = (inp[13]) ? 4'b0001 : node1434;
															assign node1434 = (inp[12]) ? 4'b1001 : 4'b0001;
											assign node1438 = (inp[13]) ? node1460 : node1439;
												assign node1439 = (inp[7]) ? node1449 : node1440;
													assign node1440 = (inp[3]) ? node1444 : node1441;
														assign node1441 = (inp[2]) ? 4'b1001 : 4'b0101;
														assign node1444 = (inp[2]) ? 4'b0101 : node1445;
															assign node1445 = (inp[12]) ? 4'b0001 : 4'b1001;
													assign node1449 = (inp[2]) ? node1455 : node1450;
														assign node1450 = (inp[12]) ? 4'b0001 : node1451;
															assign node1451 = (inp[14]) ? 4'b1001 : 4'b0001;
														assign node1455 = (inp[3]) ? 4'b0001 : node1456;
															assign node1456 = (inp[12]) ? 4'b1101 : 4'b0001;
												assign node1460 = (inp[2]) ? node1468 : node1461;
													assign node1461 = (inp[12]) ? node1463 : 4'b0101;
														assign node1463 = (inp[3]) ? node1465 : 4'b0101;
															assign node1465 = (inp[7]) ? 4'b1001 : 4'b1101;
													assign node1468 = (inp[3]) ? 4'b0101 : node1469;
														assign node1469 = (inp[12]) ? 4'b0001 : 4'b1001;
										assign node1473 = (inp[13]) ? node1517 : node1474;
											assign node1474 = (inp[2]) ? node1504 : node1475;
												assign node1475 = (inp[14]) ? node1489 : node1476;
													assign node1476 = (inp[4]) ? node1482 : node1477;
														assign node1477 = (inp[7]) ? node1479 : 4'b1001;
															assign node1479 = (inp[3]) ? 4'b1101 : 4'b0101;
														assign node1482 = (inp[7]) ? node1486 : node1483;
															assign node1483 = (inp[12]) ? 4'b1101 : 4'b0101;
															assign node1486 = (inp[3]) ? 4'b0001 : 4'b1001;
													assign node1489 = (inp[3]) ? node1497 : node1490;
														assign node1490 = (inp[4]) ? node1494 : node1491;
															assign node1491 = (inp[7]) ? 4'b0101 : 4'b1001;
															assign node1494 = (inp[7]) ? 4'b1001 : 4'b1101;
														assign node1497 = (inp[4]) ? node1501 : node1498;
															assign node1498 = (inp[7]) ? 4'b1101 : 4'b1001;
															assign node1501 = (inp[7]) ? 4'b0001 : 4'b0101;
												assign node1504 = (inp[3]) ? node1510 : node1505;
													assign node1505 = (inp[4]) ? 4'b0001 : node1506;
														assign node1506 = (inp[7]) ? 4'b0101 : 4'b0001;
													assign node1510 = (inp[4]) ? node1514 : node1511;
														assign node1511 = (inp[7]) ? 4'b0001 : 4'b1001;
														assign node1514 = (inp[7]) ? 4'b1001 : 4'b1101;
											assign node1517 = (inp[4]) ? node1525 : node1518;
												assign node1518 = (inp[3]) ? 4'b1001 : node1519;
													assign node1519 = (inp[7]) ? node1521 : 4'b1001;
														assign node1521 = (inp[2]) ? 4'b1101 : 4'b1001;
												assign node1525 = (inp[2]) ? node1527 : 4'b1101;
													assign node1527 = (inp[3]) ? 4'b1101 : 4'b1001;
							assign node1530 = (inp[2]) ? 4'b1101 : node1531;
								assign node1531 = (inp[1]) ? node1695 : node1532;
									assign node1532 = (inp[14]) ? node1596 : node1533;
										assign node1533 = (inp[3]) ? node1561 : node1534;
											assign node1534 = (inp[4]) ? node1546 : node1535;
												assign node1535 = (inp[7]) ? 4'b1101 : node1536;
													assign node1536 = (inp[13]) ? node1540 : node1537;
														assign node1537 = (inp[10]) ? 4'b0000 : 4'b1101;
														assign node1540 = (inp[12]) ? node1542 : 4'b1000;
															assign node1542 = (inp[10]) ? 4'b1000 : 4'b0000;
												assign node1546 = (inp[13]) ? node1556 : node1547;
													assign node1547 = (inp[11]) ? 4'b0000 : node1548;
														assign node1548 = (inp[10]) ? 4'b0000 : node1549;
															assign node1549 = (inp[7]) ? 4'b1101 : node1550;
																assign node1550 = (inp[12]) ? 4'b1000 : 4'b0000;
													assign node1556 = (inp[10]) ? 4'b1000 : node1557;
														assign node1557 = (inp[12]) ? 4'b0000 : 4'b1000;
											assign node1561 = (inp[13]) ? node1579 : node1562;
												assign node1562 = (inp[4]) ? node1574 : node1563;
													assign node1563 = (inp[7]) ? node1569 : node1564;
														assign node1564 = (inp[12]) ? node1566 : 4'b0100;
															assign node1566 = (inp[10]) ? 4'b0100 : 4'b1000;
														assign node1569 = (inp[12]) ? node1571 : 4'b0000;
															assign node1571 = (inp[10]) ? 4'b0000 : 4'b1000;
													assign node1574 = (inp[10]) ? 4'b0100 : node1575;
														assign node1575 = (inp[12]) ? 4'b1100 : 4'b0100;
												assign node1579 = (inp[10]) ? node1591 : node1580;
													assign node1580 = (inp[12]) ? node1586 : node1581;
														assign node1581 = (inp[7]) ? node1583 : 4'b1100;
															assign node1583 = (inp[4]) ? 4'b1100 : 4'b1000;
														assign node1586 = (inp[7]) ? node1588 : 4'b0100;
															assign node1588 = (inp[4]) ? 4'b0100 : 4'b0000;
													assign node1591 = (inp[7]) ? node1593 : 4'b1100;
														assign node1593 = (inp[4]) ? 4'b1100 : 4'b1000;
										assign node1596 = (inp[11]) ? node1648 : node1597;
											assign node1597 = (inp[13]) ? node1623 : node1598;
												assign node1598 = (inp[3]) ? node1608 : node1599;
													assign node1599 = (inp[7]) ? 4'b1101 : node1600;
														assign node1600 = (inp[4]) ? 4'b1001 : node1601;
															assign node1601 = (inp[10]) ? node1603 : 4'b1101;
																assign node1603 = (inp[12]) ? 4'b1101 : 4'b0001;
													assign node1608 = (inp[12]) ? node1618 : node1609;
														assign node1609 = (inp[10]) ? node1613 : node1610;
															assign node1610 = (inp[7]) ? 4'b1001 : 4'b1101;
															assign node1613 = (inp[4]) ? 4'b0101 : node1614;
																assign node1614 = (inp[7]) ? 4'b0001 : 4'b0101;
														assign node1618 = (inp[7]) ? 4'b1001 : node1619;
															assign node1619 = (inp[4]) ? 4'b1101 : 4'b1001;
												assign node1623 = (inp[10]) ? node1631 : node1624;
													assign node1624 = (inp[3]) ? node1626 : 4'b0001;
														assign node1626 = (inp[7]) ? node1628 : 4'b0101;
															assign node1628 = (inp[4]) ? 4'b0101 : 4'b0001;
													assign node1631 = (inp[12]) ? node1639 : node1632;
														assign node1632 = (inp[3]) ? 4'b1101 : node1633;
															assign node1633 = (inp[7]) ? node1635 : 4'b1001;
																assign node1635 = (inp[4]) ? 4'b1001 : 4'b1101;
														assign node1639 = (inp[3]) ? node1645 : node1640;
															assign node1640 = (inp[7]) ? node1642 : 4'b0001;
																assign node1642 = (inp[4]) ? 4'b0001 : 4'b1101;
															assign node1645 = (inp[7]) ? 4'b0001 : 4'b0101;
											assign node1648 = (inp[3]) ? node1666 : node1649;
												assign node1649 = (inp[4]) ? node1659 : node1650;
													assign node1650 = (inp[7]) ? 4'b1101 : node1651;
														assign node1651 = (inp[13]) ? 4'b1000 : node1652;
															assign node1652 = (inp[10]) ? 4'b0000 : node1653;
																assign node1653 = (inp[12]) ? 4'b1101 : 4'b0000;
													assign node1659 = (inp[13]) ? node1661 : 4'b0000;
														assign node1661 = (inp[12]) ? node1663 : 4'b1000;
															assign node1663 = (inp[10]) ? 4'b1000 : 4'b0000;
												assign node1666 = (inp[7]) ? node1678 : node1667;
													assign node1667 = (inp[13]) ? node1673 : node1668;
														assign node1668 = (inp[12]) ? node1670 : 4'b0100;
															assign node1670 = (inp[10]) ? 4'b0100 : 4'b1100;
														assign node1673 = (inp[12]) ? node1675 : 4'b1100;
															assign node1675 = (inp[10]) ? 4'b1100 : 4'b0100;
													assign node1678 = (inp[4]) ? node1688 : node1679;
														assign node1679 = (inp[10]) ? node1685 : node1680;
															assign node1680 = (inp[12]) ? node1682 : 4'b1000;
																assign node1682 = (inp[13]) ? 4'b0000 : 4'b1000;
															assign node1685 = (inp[13]) ? 4'b1000 : 4'b0000;
														assign node1688 = (inp[12]) ? node1690 : 4'b1100;
															assign node1690 = (inp[10]) ? node1692 : 4'b0100;
																assign node1692 = (inp[13]) ? 4'b1100 : 4'b0100;
									assign node1695 = (inp[13]) ? node1767 : node1696;
										assign node1696 = (inp[12]) ? node1724 : node1697;
											assign node1697 = (inp[3]) ? node1711 : node1698;
												assign node1698 = (inp[7]) ? node1704 : node1699;
													assign node1699 = (inp[11]) ? 4'b0001 : node1700;
														assign node1700 = (inp[14]) ? 4'b0000 : 4'b0001;
													assign node1704 = (inp[4]) ? node1706 : 4'b1101;
														assign node1706 = (inp[11]) ? 4'b0001 : node1707;
															assign node1707 = (inp[14]) ? 4'b0000 : 4'b0001;
												assign node1711 = (inp[11]) ? node1719 : node1712;
													assign node1712 = (inp[14]) ? 4'b0100 : node1713;
														assign node1713 = (inp[4]) ? 4'b0101 : node1714;
															assign node1714 = (inp[7]) ? 4'b0001 : 4'b0101;
													assign node1719 = (inp[4]) ? 4'b0101 : node1720;
														assign node1720 = (inp[7]) ? 4'b0001 : 4'b0101;
											assign node1724 = (inp[10]) ? node1746 : node1725;
												assign node1725 = (inp[3]) ? node1735 : node1726;
													assign node1726 = (inp[4]) ? node1728 : 4'b1101;
														assign node1728 = (inp[7]) ? 4'b1101 : node1729;
															assign node1729 = (inp[14]) ? node1731 : 4'b1001;
																assign node1731 = (inp[11]) ? 4'b1001 : 4'b1000;
													assign node1735 = (inp[4]) ? node1741 : node1736;
														assign node1736 = (inp[11]) ? 4'b1001 : node1737;
															assign node1737 = (inp[14]) ? 4'b1000 : 4'b1001;
														assign node1741 = (inp[7]) ? node1743 : 4'b1101;
															assign node1743 = (inp[11]) ? 4'b1001 : 4'b1000;
												assign node1746 = (inp[3]) ? node1756 : node1747;
													assign node1747 = (inp[4]) ? node1751 : node1748;
														assign node1748 = (inp[7]) ? 4'b1101 : 4'b0001;
														assign node1751 = (inp[14]) ? node1753 : 4'b0001;
															assign node1753 = (inp[11]) ? 4'b0001 : 4'b0000;
													assign node1756 = (inp[4]) ? node1762 : node1757;
														assign node1757 = (inp[7]) ? node1759 : 4'b0101;
															assign node1759 = (inp[14]) ? 4'b0000 : 4'b0001;
														assign node1762 = (inp[11]) ? 4'b0101 : node1763;
															assign node1763 = (inp[14]) ? 4'b0100 : 4'b0101;
										assign node1767 = (inp[3]) ? node1799 : node1768;
											assign node1768 = (inp[4]) ? node1782 : node1769;
												assign node1769 = (inp[7]) ? 4'b1101 : node1770;
													assign node1770 = (inp[10]) ? node1776 : node1771;
														assign node1771 = (inp[14]) ? node1773 : 4'b0001;
															assign node1773 = (inp[11]) ? 4'b0001 : 4'b0000;
														assign node1776 = (inp[11]) ? 4'b1001 : node1777;
															assign node1777 = (inp[14]) ? 4'b1000 : 4'b1001;
												assign node1782 = (inp[10]) ? node1794 : node1783;
													assign node1783 = (inp[12]) ? node1789 : node1784;
														assign node1784 = (inp[11]) ? 4'b1001 : node1785;
															assign node1785 = (inp[14]) ? 4'b1000 : 4'b1001;
														assign node1789 = (inp[14]) ? node1791 : 4'b0001;
															assign node1791 = (inp[11]) ? 4'b0001 : 4'b0000;
													assign node1794 = (inp[11]) ? 4'b1001 : node1795;
														assign node1795 = (inp[14]) ? 4'b1000 : 4'b1001;
											assign node1799 = (inp[14]) ? node1817 : node1800;
												assign node1800 = (inp[12]) ? node1806 : node1801;
													assign node1801 = (inp[7]) ? node1803 : 4'b1101;
														assign node1803 = (inp[4]) ? 4'b1101 : 4'b1001;
													assign node1806 = (inp[10]) ? node1812 : node1807;
														assign node1807 = (inp[4]) ? 4'b0101 : node1808;
															assign node1808 = (inp[7]) ? 4'b0001 : 4'b0101;
														assign node1812 = (inp[4]) ? 4'b1101 : node1813;
															assign node1813 = (inp[7]) ? 4'b1001 : 4'b1101;
												assign node1817 = (inp[11]) ? node1831 : node1818;
													assign node1818 = (inp[7]) ? node1824 : node1819;
														assign node1819 = (inp[10]) ? 4'b1100 : node1820;
															assign node1820 = (inp[12]) ? 4'b0100 : 4'b1100;
														assign node1824 = (inp[4]) ? node1826 : 4'b1000;
															assign node1826 = (inp[10]) ? 4'b1100 : node1827;
																assign node1827 = (inp[12]) ? 4'b0100 : 4'b1100;
													assign node1831 = (inp[4]) ? node1835 : node1832;
														assign node1832 = (inp[7]) ? 4'b1001 : 4'b1101;
														assign node1835 = (inp[12]) ? node1837 : 4'b1101;
															assign node1837 = (inp[10]) ? 4'b1101 : 4'b0101;
						assign node1841 = (inp[3]) ? node2649 : node1842;
							assign node1842 = (inp[1]) ? node2256 : node1843;
								assign node1843 = (inp[4]) ? node2047 : node1844;
									assign node1844 = (inp[7]) ? node1970 : node1845;
										assign node1845 = (inp[2]) ? node1907 : node1846;
											assign node1846 = (inp[11]) ? node1878 : node1847;
												assign node1847 = (inp[0]) ? node1861 : node1848;
													assign node1848 = (inp[12]) ? node1852 : node1849;
														assign node1849 = (inp[13]) ? 4'b0101 : 4'b0001;
														assign node1852 = (inp[10]) ? node1858 : node1853;
															assign node1853 = (inp[13]) ? 4'b1001 : node1854;
																assign node1854 = (inp[14]) ? 4'b1100 : 4'b1101;
															assign node1858 = (inp[13]) ? 4'b1101 : 4'b1001;
													assign node1861 = (inp[13]) ? node1871 : node1862;
														assign node1862 = (inp[14]) ? node1868 : node1863;
															assign node1863 = (inp[12]) ? node1865 : 4'b0000;
																assign node1865 = (inp[10]) ? 4'b0000 : 4'b1100;
															assign node1868 = (inp[10]) ? 4'b1000 : 4'b1101;
														assign node1871 = (inp[10]) ? node1875 : node1872;
															assign node1872 = (inp[12]) ? 4'b1000 : 4'b0000;
															assign node1875 = (inp[12]) ? 4'b0000 : 4'b1000;
												assign node1878 = (inp[0]) ? node1886 : node1879;
													assign node1879 = (inp[10]) ? node1883 : node1880;
														assign node1880 = (inp[13]) ? 4'b0101 : 4'b0001;
														assign node1883 = (inp[13]) ? 4'b0000 : 4'b0001;
													assign node1886 = (inp[13]) ? node1894 : node1887;
														assign node1887 = (inp[12]) ? node1891 : node1888;
															assign node1888 = (inp[10]) ? 4'b1001 : 4'b0001;
															assign node1891 = (inp[10]) ? 4'b0001 : 4'b1100;
														assign node1894 = (inp[14]) ? node1900 : node1895;
															assign node1895 = (inp[12]) ? node1897 : 4'b0001;
																assign node1897 = (inp[10]) ? 4'b0001 : 4'b1001;
															assign node1900 = (inp[12]) ? node1904 : node1901;
																assign node1901 = (inp[10]) ? 4'b1001 : 4'b0001;
																assign node1904 = (inp[10]) ? 4'b0001 : 4'b1001;
											assign node1907 = (inp[11]) ? node1949 : node1908;
												assign node1908 = (inp[12]) ? node1928 : node1909;
													assign node1909 = (inp[13]) ? node1921 : node1910;
														assign node1910 = (inp[10]) ? node1916 : node1911;
															assign node1911 = (inp[14]) ? 4'b0000 : node1912;
																assign node1912 = (inp[0]) ? 4'b0000 : 4'b0001;
															assign node1916 = (inp[0]) ? node1918 : 4'b1001;
																assign node1918 = (inp[14]) ? 4'b0001 : 4'b0000;
														assign node1921 = (inp[0]) ? 4'b1001 : node1922;
															assign node1922 = (inp[10]) ? node1924 : 4'b1000;
																assign node1924 = (inp[14]) ? 4'b0100 : 4'b0101;
													assign node1928 = (inp[13]) ? node1940 : node1929;
														assign node1929 = (inp[10]) ? node1933 : node1930;
															assign node1930 = (inp[0]) ? 4'b1101 : 4'b1100;
															assign node1933 = (inp[14]) ? node1937 : node1934;
																assign node1934 = (inp[0]) ? 4'b0000 : 4'b1001;
																assign node1937 = (inp[0]) ? 4'b1101 : 4'b1000;
														assign node1940 = (inp[10]) ? node1946 : node1941;
															assign node1941 = (inp[14]) ? 4'b0000 : node1942;
																assign node1942 = (inp[0]) ? 4'b0000 : 4'b0001;
															assign node1946 = (inp[14]) ? 4'b0001 : 4'b1000;
												assign node1949 = (inp[13]) ? node1959 : node1950;
													assign node1950 = (inp[12]) ? node1952 : 4'b0000;
														assign node1952 = (inp[0]) ? node1956 : node1953;
															assign node1953 = (inp[10]) ? 4'b1000 : 4'b0000;
															assign node1956 = (inp[10]) ? 4'b0000 : 4'b1101;
													assign node1959 = (inp[10]) ? node1965 : node1960;
														assign node1960 = (inp[0]) ? node1962 : 4'b1000;
															assign node1962 = (inp[14]) ? 4'b1000 : 4'b0000;
														assign node1965 = (inp[0]) ? 4'b1000 : node1966;
															assign node1966 = (inp[12]) ? 4'b0100 : 4'b1100;
										assign node1970 = (inp[2]) ? node2020 : node1971;
											assign node1971 = (inp[13]) ? node1993 : node1972;
												assign node1972 = (inp[11]) ? node1984 : node1973;
													assign node1973 = (inp[12]) ? node1977 : node1974;
														assign node1974 = (inp[14]) ? 4'b0101 : 4'b0100;
														assign node1977 = (inp[0]) ? node1981 : node1978;
															assign node1978 = (inp[14]) ? 4'b1100 : 4'b1101;
															assign node1981 = (inp[14]) ? 4'b1101 : 4'b0100;
													assign node1984 = (inp[0]) ? node1988 : node1985;
														assign node1985 = (inp[10]) ? 4'b0001 : 4'b0100;
														assign node1988 = (inp[10]) ? 4'b0100 : node1989;
															assign node1989 = (inp[12]) ? 4'b1100 : 4'b0100;
												assign node1993 = (inp[0]) ? node2003 : node1994;
													assign node1994 = (inp[10]) ? node1998 : node1995;
														assign node1995 = (inp[14]) ? 4'b1001 : 4'b0001;
														assign node1998 = (inp[12]) ? node2000 : 4'b0101;
															assign node2000 = (inp[11]) ? 4'b0101 : 4'b1001;
													assign node2003 = (inp[10]) ? node2013 : node2004;
														assign node2004 = (inp[12]) ? node2008 : node2005;
															assign node2005 = (inp[11]) ? 4'b0001 : 4'b0000;
															assign node2008 = (inp[14]) ? node2010 : 4'b0100;
																assign node2010 = (inp[11]) ? 4'b0100 : 4'b0101;
														assign node2013 = (inp[11]) ? node2017 : node2014;
															assign node2014 = (inp[14]) ? 4'b1000 : 4'b0000;
															assign node2017 = (inp[12]) ? 4'b0001 : 4'b1001;
											assign node2020 = (inp[0]) ? 4'b1101 : node2021;
												assign node2021 = (inp[13]) ? node2035 : node2022;
													assign node2022 = (inp[11]) ? node2028 : node2023;
														assign node2023 = (inp[12]) ? 4'b1100 : node2024;
															assign node2024 = (inp[10]) ? 4'b1100 : 4'b0100;
														assign node2028 = (inp[12]) ? node2032 : node2029;
															assign node2029 = (inp[10]) ? 4'b0000 : 4'b0101;
															assign node2032 = (inp[10]) ? 4'b0101 : 4'b1101;
													assign node2035 = (inp[11]) ? node2041 : node2036;
														assign node2036 = (inp[14]) ? 4'b0000 : node2037;
															assign node2037 = (inp[10]) ? 4'b0001 : 4'b1001;
														assign node2041 = (inp[10]) ? node2043 : 4'b1000;
															assign node2043 = (inp[12]) ? 4'b0000 : 4'b1000;
									assign node2047 = (inp[0]) ? node2169 : node2048;
										assign node2048 = (inp[2]) ? node2120 : node2049;
											assign node2049 = (inp[10]) ? node2071 : node2050;
												assign node2050 = (inp[14]) ? node2056 : node2051;
													assign node2051 = (inp[11]) ? node2053 : 4'b0000;
														assign node2053 = (inp[13]) ? 4'b0001 : 4'b0000;
													assign node2056 = (inp[13]) ? node2066 : node2057;
														assign node2057 = (inp[11]) ? node2063 : node2058;
															assign node2058 = (inp[7]) ? 4'b1101 : node2059;
																assign node2059 = (inp[12]) ? 4'b1001 : 4'b0001;
															assign node2063 = (inp[12]) ? 4'b0000 : 4'b1000;
														assign node2066 = (inp[11]) ? node2068 : 4'b0000;
															assign node2068 = (inp[12]) ? 4'b0001 : 4'b1001;
												assign node2071 = (inp[7]) ? node2099 : node2072;
													assign node2072 = (inp[13]) ? node2084 : node2073;
														assign node2073 = (inp[14]) ? node2081 : node2074;
															assign node2074 = (inp[11]) ? node2078 : node2075;
																assign node2075 = (inp[12]) ? 4'b0100 : 4'b1100;
																assign node2078 = (inp[12]) ? 4'b1100 : 4'b0001;
															assign node2081 = (inp[11]) ? 4'b0001 : 4'b0101;
														assign node2084 = (inp[14]) ? node2092 : node2085;
															assign node2085 = (inp[11]) ? node2089 : node2086;
																assign node2086 = (inp[12]) ? 4'b0001 : 4'b1001;
																assign node2089 = (inp[12]) ? 4'b1000 : 4'b0000;
															assign node2092 = (inp[11]) ? node2096 : node2093;
																assign node2093 = (inp[12]) ? 4'b0000 : 4'b1000;
																assign node2096 = (inp[12]) ? 4'b1000 : 4'b0000;
													assign node2099 = (inp[12]) ? node2113 : node2100;
														assign node2100 = (inp[14]) ? node2106 : node2101;
															assign node2101 = (inp[11]) ? node2103 : 4'b1000;
																assign node2103 = (inp[13]) ? 4'b0000 : 4'b1000;
															assign node2106 = (inp[13]) ? node2110 : node2107;
																assign node2107 = (inp[11]) ? 4'b1000 : 4'b0001;
																assign node2110 = (inp[11]) ? 4'b0000 : 4'b1000;
														assign node2113 = (inp[11]) ? node2117 : node2114;
															assign node2114 = (inp[13]) ? 4'b1000 : 4'b0001;
															assign node2117 = (inp[13]) ? 4'b1001 : 4'b1000;
											assign node2120 = (inp[11]) ? node2156 : node2121;
												assign node2121 = (inp[12]) ? node2139 : node2122;
													assign node2122 = (inp[14]) ? node2132 : node2123;
														assign node2123 = (inp[10]) ? node2129 : node2124;
															assign node2124 = (inp[7]) ? 4'b0001 : node2125;
																assign node2125 = (inp[13]) ? 4'b0101 : 4'b0001;
															assign node2129 = (inp[13]) ? 4'b0000 : 4'b0001;
														assign node2132 = (inp[13]) ? 4'b0101 : node2133;
															assign node2133 = (inp[10]) ? 4'b0001 : node2134;
																assign node2134 = (inp[7]) ? 4'b0100 : 4'b0001;
													assign node2139 = (inp[13]) ? 4'b1001 : node2140;
														assign node2140 = (inp[14]) ? node2148 : node2141;
															assign node2141 = (inp[10]) ? node2145 : node2142;
																assign node2142 = (inp[7]) ? 4'b1001 : 4'b1101;
																assign node2145 = (inp[7]) ? 4'b1101 : 4'b1001;
															assign node2148 = (inp[7]) ? node2152 : node2149;
																assign node2149 = (inp[10]) ? 4'b1001 : 4'b1100;
																assign node2152 = (inp[10]) ? 4'b1100 : 4'b1000;
												assign node2156 = (inp[13]) ? node2162 : node2157;
													assign node2157 = (inp[7]) ? node2159 : 4'b0001;
														assign node2159 = (inp[10]) ? 4'b0001 : 4'b0100;
													assign node2162 = (inp[10]) ? 4'b0000 : node2163;
														assign node2163 = (inp[7]) ? 4'b0001 : node2164;
															assign node2164 = (inp[12]) ? 4'b0101 : 4'b0000;
										assign node2169 = (inp[2]) ? node2219 : node2170;
											assign node2170 = (inp[11]) ? node2200 : node2171;
												assign node2171 = (inp[13]) ? node2185 : node2172;
													assign node2172 = (inp[7]) ? node2180 : node2173;
														assign node2173 = (inp[12]) ? node2177 : node2174;
															assign node2174 = (inp[10]) ? 4'b1100 : 4'b0100;
															assign node2177 = (inp[10]) ? 4'b0100 : 4'b1000;
														assign node2180 = (inp[10]) ? 4'b0000 : node2181;
															assign node2181 = (inp[12]) ? 4'b1000 : 4'b0000;
													assign node2185 = (inp[14]) ? node2193 : node2186;
														assign node2186 = (inp[10]) ? 4'b0001 : node2187;
															assign node2187 = (inp[12]) ? node2189 : 4'b0100;
																assign node2189 = (inp[7]) ? 4'b1000 : 4'b0001;
														assign node2193 = (inp[10]) ? 4'b0000 : node2194;
															assign node2194 = (inp[12]) ? node2196 : 4'b0100;
																assign node2196 = (inp[7]) ? 4'b1000 : 4'b0000;
												assign node2200 = (inp[13]) ? node2210 : node2201;
													assign node2201 = (inp[12]) ? node2207 : node2202;
														assign node2202 = (inp[10]) ? 4'b0000 : node2203;
															assign node2203 = (inp[7]) ? 4'b0001 : 4'b0101;
														assign node2207 = (inp[10]) ? 4'b0001 : 4'b1001;
													assign node2210 = (inp[7]) ? node2212 : 4'b1000;
														assign node2212 = (inp[10]) ? node2216 : node2213;
															assign node2213 = (inp[12]) ? 4'b1001 : 4'b0101;
															assign node2216 = (inp[12]) ? 4'b0000 : 4'b1000;
											assign node2219 = (inp[14]) ? node2233 : node2220;
												assign node2220 = (inp[13]) ? node2228 : node2221;
													assign node2221 = (inp[12]) ? node2223 : 4'b0000;
														assign node2223 = (inp[10]) ? 4'b0000 : node2224;
															assign node2224 = (inp[7]) ? 4'b1101 : 4'b1000;
													assign node2228 = (inp[10]) ? 4'b1000 : node2229;
														assign node2229 = (inp[12]) ? 4'b0000 : 4'b1000;
												assign node2233 = (inp[11]) ? node2245 : node2234;
													assign node2234 = (inp[13]) ? node2242 : node2235;
														assign node2235 = (inp[7]) ? node2237 : 4'b1001;
															assign node2237 = (inp[12]) ? 4'b1101 : node2238;
																assign node2238 = (inp[10]) ? 4'b0001 : 4'b1101;
														assign node2242 = (inp[12]) ? 4'b0001 : 4'b1001;
													assign node2245 = (inp[13]) ? node2251 : node2246;
														assign node2246 = (inp[12]) ? node2248 : 4'b0000;
															assign node2248 = (inp[7]) ? 4'b0000 : 4'b1000;
														assign node2251 = (inp[10]) ? 4'b1000 : node2252;
															assign node2252 = (inp[12]) ? 4'b0000 : 4'b1000;
								assign node2256 = (inp[11]) ? node2492 : node2257;
									assign node2257 = (inp[4]) ? node2373 : node2258;
										assign node2258 = (inp[7]) ? node2322 : node2259;
											assign node2259 = (inp[13]) ? node2283 : node2260;
												assign node2260 = (inp[2]) ? node2268 : node2261;
													assign node2261 = (inp[0]) ? node2265 : node2262;
														assign node2262 = (inp[12]) ? 4'b0001 : 4'b1001;
														assign node2265 = (inp[10]) ? 4'b1000 : 4'b0000;
													assign node2268 = (inp[0]) ? node2276 : node2269;
														assign node2269 = (inp[14]) ? 4'b0001 : node2270;
															assign node2270 = (inp[10]) ? 4'b0000 : node2271;
																assign node2271 = (inp[12]) ? 4'b0000 : 4'b1000;
														assign node2276 = (inp[14]) ? 4'b0000 : node2277;
															assign node2277 = (inp[10]) ? 4'b0001 : node2278;
																assign node2278 = (inp[12]) ? 4'b1101 : 4'b0001;
												assign node2283 = (inp[0]) ? node2307 : node2284;
													assign node2284 = (inp[2]) ? node2296 : node2285;
														assign node2285 = (inp[10]) ? node2289 : node2286;
															assign node2286 = (inp[12]) ? 4'b0101 : 4'b1101;
															assign node2289 = (inp[12]) ? node2293 : node2290;
																assign node2290 = (inp[14]) ? 4'b1000 : 4'b1001;
																assign node2293 = (inp[14]) ? 4'b0000 : 4'b0001;
														assign node2296 = (inp[14]) ? node2304 : node2297;
															assign node2297 = (inp[12]) ? node2301 : node2298;
																assign node2298 = (inp[10]) ? 4'b1100 : 4'b0100;
																assign node2301 = (inp[10]) ? 4'b1100 : 4'b1000;
															assign node2304 = (inp[10]) ? 4'b1101 : 4'b1001;
													assign node2307 = (inp[14]) ? node2317 : node2308;
														assign node2308 = (inp[2]) ? node2312 : node2309;
															assign node2309 = (inp[10]) ? 4'b1000 : 4'b0000;
															assign node2312 = (inp[10]) ? 4'b1001 : node2313;
																assign node2313 = (inp[12]) ? 4'b0001 : 4'b1001;
														assign node2317 = (inp[10]) ? 4'b1000 : node2318;
															assign node2318 = (inp[12]) ? 4'b0000 : 4'b1000;
											assign node2322 = (inp[13]) ? node2346 : node2323;
												assign node2323 = (inp[0]) ? node2337 : node2324;
													assign node2324 = (inp[10]) ? node2330 : node2325;
														assign node2325 = (inp[14]) ? node2327 : 4'b0100;
															assign node2327 = (inp[2]) ? 4'b0100 : 4'b0101;
														assign node2330 = (inp[2]) ? node2334 : node2331;
															assign node2331 = (inp[12]) ? 4'b0001 : 4'b1001;
															assign node2334 = (inp[14]) ? 4'b0001 : 4'b0000;
													assign node2337 = (inp[2]) ? 4'b1101 : node2338;
														assign node2338 = (inp[14]) ? node2340 : 4'b0101;
															assign node2340 = (inp[10]) ? 4'b0100 : node2341;
																assign node2341 = (inp[12]) ? 4'b1100 : 4'b0100;
												assign node2346 = (inp[10]) ? node2360 : node2347;
													assign node2347 = (inp[2]) ? node2353 : node2348;
														assign node2348 = (inp[0]) ? 4'b0000 : node2349;
															assign node2349 = (inp[12]) ? 4'b0001 : 4'b1001;
														assign node2353 = (inp[0]) ? 4'b1101 : node2354;
															assign node2354 = (inp[14]) ? 4'b1001 : node2355;
																assign node2355 = (inp[12]) ? 4'b1000 : 4'b0000;
													assign node2360 = (inp[0]) ? node2370 : node2361;
														assign node2361 = (inp[2]) ? node2365 : node2362;
															assign node2362 = (inp[12]) ? 4'b0101 : 4'b1101;
															assign node2365 = (inp[14]) ? node2367 : 4'b1000;
																assign node2367 = (inp[12]) ? 4'b0001 : 4'b1001;
														assign node2370 = (inp[2]) ? 4'b1101 : 4'b1000;
										assign node2373 = (inp[2]) ? node2429 : node2374;
											assign node2374 = (inp[10]) ? node2400 : node2375;
												assign node2375 = (inp[0]) ? node2385 : node2376;
													assign node2376 = (inp[12]) ? 4'b1000 : node2377;
														assign node2377 = (inp[13]) ? node2381 : node2378;
															assign node2378 = (inp[14]) ? 4'b1000 : 4'b1001;
															assign node2381 = (inp[7]) ? 4'b0000 : 4'b0100;
													assign node2385 = (inp[14]) ? node2393 : node2386;
														assign node2386 = (inp[12]) ? node2388 : 4'b0000;
															assign node2388 = (inp[7]) ? node2390 : 4'b0100;
																assign node2390 = (inp[13]) ? 4'b0100 : 4'b0000;
														assign node2393 = (inp[13]) ? node2397 : node2394;
															assign node2394 = (inp[12]) ? 4'b0000 : 4'b0100;
															assign node2397 = (inp[7]) ? 4'b0100 : 4'b1001;
												assign node2400 = (inp[14]) ? node2418 : node2401;
													assign node2401 = (inp[7]) ? node2411 : node2402;
														assign node2402 = (inp[13]) ? node2408 : node2403;
															assign node2403 = (inp[0]) ? 4'b0000 : node2404;
																assign node2404 = (inp[12]) ? 4'b0000 : 4'b1000;
															assign node2408 = (inp[0]) ? 4'b1000 : 4'b0000;
														assign node2411 = (inp[13]) ? 4'b1000 : node2412;
															assign node2412 = (inp[12]) ? node2414 : 4'b0101;
																assign node2414 = (inp[0]) ? 4'b1000 : 4'b1001;
													assign node2418 = (inp[13]) ? 4'b0001 : node2419;
														assign node2419 = (inp[12]) ? node2425 : node2420;
															assign node2420 = (inp[0]) ? node2422 : 4'b1000;
																assign node2422 = (inp[7]) ? 4'b1000 : 4'b0001;
															assign node2425 = (inp[7]) ? 4'b1000 : 4'b1100;
											assign node2429 = (inp[14]) ? node2455 : node2430;
												assign node2430 = (inp[12]) ? node2442 : node2431;
													assign node2431 = (inp[0]) ? node2439 : node2432;
														assign node2432 = (inp[10]) ? 4'b1001 : node2433;
															assign node2433 = (inp[13]) ? 4'b1001 : node2434;
																assign node2434 = (inp[7]) ? 4'b1100 : 4'b1001;
														assign node2439 = (inp[13]) ? 4'b1001 : 4'b0001;
													assign node2442 = (inp[0]) ? node2448 : node2443;
														assign node2443 = (inp[7]) ? node2445 : 4'b0001;
															assign node2445 = (inp[13]) ? 4'b0001 : 4'b0100;
														assign node2448 = (inp[10]) ? node2452 : node2449;
															assign node2449 = (inp[13]) ? 4'b0001 : 4'b1101;
															assign node2452 = (inp[13]) ? 4'b1001 : 4'b0001;
												assign node2455 = (inp[0]) ? node2479 : node2456;
													assign node2456 = (inp[13]) ? node2468 : node2457;
														assign node2457 = (inp[12]) ? node2463 : node2458;
															assign node2458 = (inp[10]) ? 4'b1001 : node2459;
																assign node2459 = (inp[7]) ? 4'b0101 : 4'b1001;
															assign node2463 = (inp[7]) ? node2465 : 4'b0001;
																assign node2465 = (inp[10]) ? 4'b0001 : 4'b0101;
														assign node2468 = (inp[7]) ? node2474 : node2469;
															assign node2469 = (inp[10]) ? node2471 : 4'b0000;
																assign node2471 = (inp[12]) ? 4'b0000 : 4'b1000;
															assign node2474 = (inp[12]) ? node2476 : 4'b1001;
																assign node2476 = (inp[10]) ? 4'b0000 : 4'b0001;
													assign node2479 = (inp[13]) ? node2487 : node2480;
														assign node2480 = (inp[10]) ? 4'b0000 : node2481;
															assign node2481 = (inp[12]) ? node2483 : 4'b0000;
																assign node2483 = (inp[7]) ? 4'b1101 : 4'b1000;
														assign node2487 = (inp[12]) ? node2489 : 4'b1000;
															assign node2489 = (inp[10]) ? 4'b1000 : 4'b0000;
									assign node2492 = (inp[10]) ? node2588 : node2493;
										assign node2493 = (inp[2]) ? node2539 : node2494;
											assign node2494 = (inp[0]) ? node2518 : node2495;
												assign node2495 = (inp[4]) ? node2509 : node2496;
													assign node2496 = (inp[12]) ? node2502 : node2497;
														assign node2497 = (inp[14]) ? 4'b1001 : node2498;
															assign node2498 = (inp[7]) ? 4'b1101 : 4'b1001;
														assign node2502 = (inp[7]) ? node2506 : node2503;
															assign node2503 = (inp[13]) ? 4'b1101 : 4'b1001;
															assign node2506 = (inp[13]) ? 4'b1001 : 4'b0101;
													assign node2509 = (inp[12]) ? node2515 : node2510;
														assign node2510 = (inp[13]) ? 4'b0001 : node2511;
															assign node2511 = (inp[7]) ? 4'b0001 : 4'b0101;
														assign node2515 = (inp[13]) ? 4'b0101 : 4'b1001;
												assign node2518 = (inp[13]) ? node2534 : node2519;
													assign node2519 = (inp[12]) ? node2527 : node2520;
														assign node2520 = (inp[7]) ? node2524 : node2521;
															assign node2521 = (inp[4]) ? 4'b0101 : 4'b0001;
															assign node2524 = (inp[4]) ? 4'b0001 : 4'b0101;
														assign node2527 = (inp[7]) ? node2531 : node2528;
															assign node2528 = (inp[4]) ? 4'b0101 : 4'b0001;
															assign node2531 = (inp[4]) ? 4'b0001 : 4'b1101;
													assign node2534 = (inp[4]) ? node2536 : 4'b0001;
														assign node2536 = (inp[12]) ? 4'b0101 : 4'b0001;
											assign node2539 = (inp[7]) ? node2567 : node2540;
												assign node2540 = (inp[4]) ? node2556 : node2541;
													assign node2541 = (inp[13]) ? node2549 : node2542;
														assign node2542 = (inp[0]) ? node2546 : node2543;
															assign node2543 = (inp[12]) ? 4'b0001 : 4'b1001;
															assign node2546 = (inp[12]) ? 4'b1101 : 4'b0001;
														assign node2549 = (inp[12]) ? node2553 : node2550;
															assign node2550 = (inp[0]) ? 4'b1001 : 4'b0101;
															assign node2553 = (inp[0]) ? 4'b0001 : 4'b1001;
													assign node2556 = (inp[0]) ? node2562 : node2557;
														assign node2557 = (inp[12]) ? node2559 : 4'b1001;
															assign node2559 = (inp[13]) ? 4'b0001 : 4'b1001;
														assign node2562 = (inp[13]) ? 4'b0001 : node2563;
															assign node2563 = (inp[12]) ? 4'b1001 : 4'b0001;
												assign node2567 = (inp[13]) ? node2579 : node2568;
													assign node2568 = (inp[0]) ? node2574 : node2569;
														assign node2569 = (inp[12]) ? 4'b0101 : node2570;
															assign node2570 = (inp[4]) ? 4'b1101 : 4'b0101;
														assign node2574 = (inp[12]) ? 4'b1101 : node2575;
															assign node2575 = (inp[4]) ? 4'b0001 : 4'b1101;
													assign node2579 = (inp[4]) ? node2583 : node2580;
														assign node2580 = (inp[0]) ? 4'b1101 : 4'b0001;
														assign node2583 = (inp[12]) ? node2585 : 4'b1001;
															assign node2585 = (inp[0]) ? 4'b0001 : 4'b1001;
										assign node2588 = (inp[13]) ? node2624 : node2589;
											assign node2589 = (inp[2]) ? node2611 : node2590;
												assign node2590 = (inp[7]) ? node2596 : node2591;
													assign node2591 = (inp[4]) ? node2593 : 4'b1001;
														assign node2593 = (inp[0]) ? 4'b0001 : 4'b1001;
													assign node2596 = (inp[14]) ? node2598 : 4'b1001;
														assign node2598 = (inp[12]) ? node2604 : node2599;
															assign node2599 = (inp[4]) ? 4'b0101 : node2600;
																assign node2600 = (inp[0]) ? 4'b0101 : 4'b1001;
															assign node2604 = (inp[4]) ? node2608 : node2605;
																assign node2605 = (inp[0]) ? 4'b0101 : 4'b1001;
																assign node2608 = (inp[0]) ? 4'b1001 : 4'b0101;
												assign node2611 = (inp[7]) ? node2617 : node2612;
													assign node2612 = (inp[4]) ? node2614 : 4'b0001;
														assign node2614 = (inp[0]) ? 4'b0001 : 4'b1001;
													assign node2617 = (inp[4]) ? node2621 : node2618;
														assign node2618 = (inp[0]) ? 4'b1101 : 4'b0001;
														assign node2621 = (inp[0]) ? 4'b0001 : 4'b1001;
											assign node2624 = (inp[4]) ? 4'b1001 : node2625;
												assign node2625 = (inp[7]) ? node2631 : node2626;
													assign node2626 = (inp[2]) ? node2628 : 4'b1001;
														assign node2628 = (inp[0]) ? 4'b1001 : 4'b1101;
													assign node2631 = (inp[12]) ? node2641 : node2632;
														assign node2632 = (inp[14]) ? 4'b1001 : node2633;
															assign node2633 = (inp[2]) ? node2637 : node2634;
																assign node2634 = (inp[0]) ? 4'b1001 : 4'b1101;
																assign node2637 = (inp[0]) ? 4'b1101 : 4'b1001;
														assign node2641 = (inp[2]) ? node2645 : node2642;
															assign node2642 = (inp[0]) ? 4'b1001 : 4'b1101;
															assign node2645 = (inp[0]) ? 4'b1101 : 4'b1001;
							assign node2649 = (inp[4]) ? node3017 : node2650;
								assign node2650 = (inp[11]) ? node2870 : node2651;
									assign node2651 = (inp[10]) ? node2763 : node2652;
										assign node2652 = (inp[1]) ? node2722 : node2653;
											assign node2653 = (inp[0]) ? node2687 : node2654;
												assign node2654 = (inp[7]) ? node2674 : node2655;
													assign node2655 = (inp[14]) ? node2665 : node2656;
														assign node2656 = (inp[2]) ? node2662 : node2657;
															assign node2657 = (inp[12]) ? node2659 : 4'b0001;
																assign node2659 = (inp[13]) ? 4'b0000 : 4'b0001;
															assign node2662 = (inp[13]) ? 4'b0001 : 4'b0000;
														assign node2665 = (inp[12]) ? 4'b0001 : node2666;
															assign node2666 = (inp[2]) ? node2670 : node2667;
																assign node2667 = (inp[13]) ? 4'b0000 : 4'b0001;
																assign node2670 = (inp[13]) ? 4'b0001 : 4'b0000;
													assign node2674 = (inp[2]) ? node2680 : node2675;
														assign node2675 = (inp[12]) ? 4'b0000 : node2676;
															assign node2676 = (inp[13]) ? 4'b1000 : 4'b0000;
														assign node2680 = (inp[13]) ? 4'b1001 : node2681;
															assign node2681 = (inp[14]) ? node2683 : 4'b0000;
																assign node2683 = (inp[12]) ? 4'b1001 : 4'b0001;
												assign node2687 = (inp[12]) ? node2705 : node2688;
													assign node2688 = (inp[2]) ? node2700 : node2689;
														assign node2689 = (inp[7]) ? node2695 : node2690;
															assign node2690 = (inp[13]) ? node2692 : 4'b0001;
																assign node2692 = (inp[14]) ? 4'b1001 : 4'b1000;
															assign node2695 = (inp[13]) ? 4'b0001 : node2696;
																assign node2696 = (inp[14]) ? 4'b0000 : 4'b0001;
														assign node2700 = (inp[13]) ? 4'b0000 : node2701;
															assign node2701 = (inp[7]) ? 4'b1001 : 4'b0000;
													assign node2705 = (inp[7]) ? node2711 : node2706;
														assign node2706 = (inp[14]) ? node2708 : 4'b1000;
															assign node2708 = (inp[13]) ? 4'b1000 : 4'b1001;
														assign node2711 = (inp[13]) ? node2717 : node2712;
															assign node2712 = (inp[2]) ? 4'b1001 : node2713;
																assign node2713 = (inp[14]) ? 4'b1000 : 4'b1001;
															assign node2717 = (inp[2]) ? node2719 : 4'b1001;
																assign node2719 = (inp[14]) ? 4'b0001 : 4'b0000;
											assign node2722 = (inp[2]) ? node2746 : node2723;
												assign node2723 = (inp[13]) ? node2733 : node2724;
													assign node2724 = (inp[0]) ? node2726 : 4'b0001;
														assign node2726 = (inp[12]) ? node2730 : node2727;
															assign node2727 = (inp[7]) ? 4'b0001 : 4'b1001;
															assign node2730 = (inp[7]) ? 4'b0000 : 4'b0001;
													assign node2733 = (inp[0]) ? node2739 : node2734;
														assign node2734 = (inp[14]) ? 4'b0001 : node2735;
															assign node2735 = (inp[12]) ? 4'b0000 : 4'b0001;
														assign node2739 = (inp[14]) ? 4'b0000 : node2740;
															assign node2740 = (inp[7]) ? 4'b0001 : node2741;
																assign node2741 = (inp[12]) ? 4'b0001 : 4'b0000;
												assign node2746 = (inp[13]) ? node2760 : node2747;
													assign node2747 = (inp[12]) ? node2755 : node2748;
														assign node2748 = (inp[0]) ? node2750 : 4'b0000;
															assign node2750 = (inp[7]) ? node2752 : 4'b0000;
																assign node2752 = (inp[14]) ? 4'b0000 : 4'b0001;
														assign node2755 = (inp[7]) ? 4'b1001 : node2756;
															assign node2756 = (inp[0]) ? 4'b0000 : 4'b1000;
													assign node2760 = (inp[0]) ? 4'b0000 : 4'b0001;
										assign node2763 = (inp[2]) ? node2821 : node2764;
											assign node2764 = (inp[1]) ? node2794 : node2765;
												assign node2765 = (inp[13]) ? node2781 : node2766;
													assign node2766 = (inp[12]) ? node2772 : node2767;
														assign node2767 = (inp[7]) ? 4'b0001 : node2768;
															assign node2768 = (inp[0]) ? 4'b0001 : 4'b1001;
														assign node2772 = (inp[0]) ? node2776 : node2773;
															assign node2773 = (inp[7]) ? 4'b0001 : 4'b1000;
															assign node2776 = (inp[14]) ? node2778 : 4'b1001;
																assign node2778 = (inp[7]) ? 4'b1000 : 4'b1001;
													assign node2781 = (inp[7]) ? node2787 : node2782;
														assign node2782 = (inp[0]) ? 4'b1000 : node2783;
															assign node2783 = (inp[14]) ? 4'b0001 : 4'b1000;
														assign node2787 = (inp[14]) ? 4'b1001 : node2788;
															assign node2788 = (inp[0]) ? 4'b0000 : node2789;
																assign node2789 = (inp[12]) ? 4'b0001 : 4'b1001;
												assign node2794 = (inp[0]) ? node2808 : node2795;
													assign node2795 = (inp[7]) ? node2797 : 4'b0000;
														assign node2797 = (inp[14]) ? node2803 : node2798;
															assign node2798 = (inp[13]) ? node2800 : 4'b1001;
																assign node2800 = (inp[12]) ? 4'b1001 : 4'b0000;
															assign node2803 = (inp[12]) ? 4'b1000 : node2804;
																assign node2804 = (inp[13]) ? 4'b0000 : 4'b1000;
													assign node2808 = (inp[13]) ? node2814 : node2809;
														assign node2809 = (inp[7]) ? node2811 : 4'b0001;
															assign node2811 = (inp[12]) ? 4'b0001 : 4'b1001;
														assign node2814 = (inp[14]) ? node2818 : node2815;
															assign node2815 = (inp[12]) ? 4'b0000 : 4'b1000;
															assign node2818 = (inp[7]) ? 4'b0000 : 4'b0001;
											assign node2821 = (inp[13]) ? node2841 : node2822;
												assign node2822 = (inp[7]) ? node2836 : node2823;
													assign node2823 = (inp[1]) ? node2831 : node2824;
														assign node2824 = (inp[0]) ? node2828 : node2825;
															assign node2825 = (inp[14]) ? 4'b0000 : 4'b1000;
															assign node2828 = (inp[12]) ? 4'b0000 : 4'b1000;
														assign node2831 = (inp[0]) ? 4'b1000 : node2832;
															assign node2832 = (inp[14]) ? 4'b1001 : 4'b1000;
													assign node2836 = (inp[0]) ? 4'b0000 : node2837;
														assign node2837 = (inp[1]) ? 4'b0000 : 4'b1000;
												assign node2841 = (inp[0]) ? node2855 : node2842;
													assign node2842 = (inp[14]) ? node2844 : 4'b0000;
														assign node2844 = (inp[1]) ? node2852 : node2845;
															assign node2845 = (inp[12]) ? node2849 : node2846;
																assign node2846 = (inp[7]) ? 4'b0001 : 4'b0000;
																assign node2849 = (inp[7]) ? 4'b0001 : 4'b1001;
															assign node2852 = (inp[7]) ? 4'b0000 : 4'b0001;
													assign node2855 = (inp[7]) ? node2865 : node2856;
														assign node2856 = (inp[1]) ? node2860 : node2857;
															assign node2857 = (inp[14]) ? 4'b0000 : 4'b0001;
															assign node2860 = (inp[14]) ? node2862 : 4'b1000;
																assign node2862 = (inp[12]) ? 4'b0001 : 4'b1001;
														assign node2865 = (inp[12]) ? node2867 : 4'b1000;
															assign node2867 = (inp[1]) ? 4'b1000 : 4'b0000;
									assign node2870 = (inp[1]) ? node2962 : node2871;
										assign node2871 = (inp[7]) ? node2917 : node2872;
											assign node2872 = (inp[2]) ? node2892 : node2873;
												assign node2873 = (inp[13]) ? node2879 : node2874;
													assign node2874 = (inp[0]) ? 4'b0001 : node2875;
														assign node2875 = (inp[10]) ? 4'b0000 : 4'b1001;
													assign node2879 = (inp[10]) ? node2885 : node2880;
														assign node2880 = (inp[0]) ? node2882 : 4'b1000;
															assign node2882 = (inp[12]) ? 4'b1000 : 4'b0000;
														assign node2885 = (inp[12]) ? node2889 : node2886;
															assign node2886 = (inp[0]) ? 4'b0000 : 4'b0001;
															assign node2889 = (inp[0]) ? 4'b1001 : 4'b0000;
												assign node2892 = (inp[10]) ? node2902 : node2893;
													assign node2893 = (inp[12]) ? node2897 : node2894;
														assign node2894 = (inp[0]) ? 4'b0001 : 4'b1001;
														assign node2897 = (inp[13]) ? 4'b1001 : node2898;
															assign node2898 = (inp[0]) ? 4'b1000 : 4'b0001;
													assign node2902 = (inp[12]) ? node2910 : node2903;
														assign node2903 = (inp[13]) ? node2907 : node2904;
															assign node2904 = (inp[0]) ? 4'b1001 : 4'b1000;
															assign node2907 = (inp[0]) ? 4'b1000 : 4'b1001;
														assign node2910 = (inp[13]) ? node2914 : node2911;
															assign node2911 = (inp[0]) ? 4'b0001 : 4'b0000;
															assign node2914 = (inp[0]) ? 4'b0000 : 4'b0001;
											assign node2917 = (inp[0]) ? node2935 : node2918;
												assign node2918 = (inp[2]) ? node2926 : node2919;
													assign node2919 = (inp[10]) ? 4'b0000 : node2920;
														assign node2920 = (inp[13]) ? node2922 : 4'b1000;
															assign node2922 = (inp[14]) ? 4'b1001 : 4'b0001;
													assign node2926 = (inp[13]) ? node2932 : node2927;
														assign node2927 = (inp[10]) ? node2929 : 4'b1000;
															assign node2929 = (inp[12]) ? 4'b1001 : 4'b0001;
														assign node2932 = (inp[10]) ? 4'b1000 : 4'b0000;
												assign node2935 = (inp[13]) ? node2947 : node2936;
													assign node2936 = (inp[12]) ? node2942 : node2937;
														assign node2937 = (inp[10]) ? node2939 : 4'b0000;
															assign node2939 = (inp[2]) ? 4'b0000 : 4'b0001;
														assign node2942 = (inp[10]) ? 4'b0000 : node2943;
															assign node2943 = (inp[2]) ? 4'b1000 : 4'b0000;
													assign node2947 = (inp[10]) ? node2955 : node2948;
														assign node2948 = (inp[12]) ? node2952 : node2949;
															assign node2949 = (inp[2]) ? 4'b0001 : 4'b0000;
															assign node2952 = (inp[2]) ? 4'b0000 : 4'b0001;
														assign node2955 = (inp[2]) ? node2959 : node2956;
															assign node2956 = (inp[12]) ? 4'b0000 : 4'b0001;
															assign node2959 = (inp[12]) ? 4'b0001 : 4'b1001;
										assign node2962 = (inp[10]) ? node3002 : node2963;
											assign node2963 = (inp[0]) ? node2981 : node2964;
												assign node2964 = (inp[13]) ? node2972 : node2965;
													assign node2965 = (inp[2]) ? 4'b0001 : node2966;
														assign node2966 = (inp[7]) ? 4'b1001 : node2967;
															assign node2967 = (inp[12]) ? 4'b1001 : 4'b0001;
													assign node2972 = (inp[2]) ? node2976 : node2973;
														assign node2973 = (inp[7]) ? 4'b0001 : 4'b1001;
														assign node2976 = (inp[12]) ? node2978 : 4'b1001;
															assign node2978 = (inp[7]) ? 4'b1001 : 4'b0001;
												assign node2981 = (inp[2]) ? node2993 : node2982;
													assign node2982 = (inp[12]) ? node2988 : node2983;
														assign node2983 = (inp[13]) ? node2985 : 4'b1001;
															assign node2985 = (inp[7]) ? 4'b1001 : 4'b0001;
														assign node2988 = (inp[13]) ? 4'b0001 : node2989;
															assign node2989 = (inp[14]) ? 4'b1001 : 4'b0001;
													assign node2993 = (inp[12]) ? node2995 : 4'b0001;
														assign node2995 = (inp[14]) ? node2997 : 4'b0001;
															assign node2997 = (inp[7]) ? node2999 : 4'b0001;
																assign node2999 = (inp[13]) ? 4'b0001 : 4'b1001;
											assign node3002 = (inp[13]) ? 4'b1001 : node3003;
												assign node3003 = (inp[0]) ? node3009 : node3004;
													assign node3004 = (inp[7]) ? 4'b0001 : node3005;
														assign node3005 = (inp[2]) ? 4'b0001 : 4'b1001;
													assign node3009 = (inp[2]) ? node3013 : node3010;
														assign node3010 = (inp[7]) ? 4'b1001 : 4'b0001;
														assign node3013 = (inp[7]) ? 4'b0001 : 4'b1001;
								assign node3017 = (inp[13]) ? node3223 : node3018;
									assign node3018 = (inp[1]) ? node3140 : node3019;
										assign node3019 = (inp[11]) ? node3089 : node3020;
											assign node3020 = (inp[10]) ? node3046 : node3021;
												assign node3021 = (inp[0]) ? node3035 : node3022;
													assign node3022 = (inp[12]) ? node3032 : node3023;
														assign node3023 = (inp[7]) ? node3029 : node3024;
															assign node3024 = (inp[14]) ? 4'b1001 : node3025;
																assign node3025 = (inp[2]) ? 4'b1001 : 4'b0000;
															assign node3029 = (inp[14]) ? 4'b1000 : 4'b1001;
														assign node3032 = (inp[2]) ? 4'b0001 : 4'b1001;
													assign node3035 = (inp[14]) ? node3041 : node3036;
														assign node3036 = (inp[2]) ? node3038 : 4'b0001;
															assign node3038 = (inp[12]) ? 4'b1001 : 4'b0001;
														assign node3041 = (inp[7]) ? node3043 : 4'b0001;
															assign node3043 = (inp[12]) ? 4'b1000 : 4'b0000;
												assign node3046 = (inp[2]) ? node3068 : node3047;
													assign node3047 = (inp[14]) ? node3061 : node3048;
														assign node3048 = (inp[7]) ? node3054 : node3049;
															assign node3049 = (inp[0]) ? 4'b0001 : node3050;
																assign node3050 = (inp[12]) ? 4'b1000 : 4'b0001;
															assign node3054 = (inp[12]) ? node3058 : node3055;
																assign node3055 = (inp[0]) ? 4'b0000 : 4'b1000;
																assign node3058 = (inp[0]) ? 4'b1000 : 4'b0000;
														assign node3061 = (inp[7]) ? node3063 : 4'b0000;
															assign node3063 = (inp[12]) ? 4'b0001 : node3064;
																assign node3064 = (inp[0]) ? 4'b0000 : 4'b0001;
													assign node3068 = (inp[7]) ? node3076 : node3069;
														assign node3069 = (inp[14]) ? node3073 : node3070;
															assign node3070 = (inp[0]) ? 4'b1000 : 4'b0000;
															assign node3073 = (inp[12]) ? 4'b1001 : 4'b0001;
														assign node3076 = (inp[14]) ? node3084 : node3077;
															assign node3077 = (inp[12]) ? node3081 : node3078;
																assign node3078 = (inp[0]) ? 4'b0001 : 4'b1001;
																assign node3081 = (inp[0]) ? 4'b1001 : 4'b0001;
															assign node3084 = (inp[0]) ? 4'b1000 : node3085;
																assign node3085 = (inp[12]) ? 4'b0000 : 4'b1000;
											assign node3089 = (inp[2]) ? node3115 : node3090;
												assign node3090 = (inp[7]) ? node3104 : node3091;
													assign node3091 = (inp[12]) ? node3099 : node3092;
														assign node3092 = (inp[0]) ? node3096 : node3093;
															assign node3093 = (inp[10]) ? 4'b0000 : 4'b0001;
															assign node3096 = (inp[10]) ? 4'b0001 : 4'b0000;
														assign node3099 = (inp[10]) ? 4'b0001 : node3100;
															assign node3100 = (inp[0]) ? 4'b1001 : 4'b1000;
													assign node3104 = (inp[10]) ? node3108 : node3105;
														assign node3105 = (inp[0]) ? 4'b1000 : 4'b0000;
														assign node3108 = (inp[12]) ? node3112 : node3109;
															assign node3109 = (inp[0]) ? 4'b0000 : 4'b1000;
															assign node3112 = (inp[0]) ? 4'b0001 : 4'b0000;
												assign node3115 = (inp[0]) ? node3127 : node3116;
													assign node3116 = (inp[10]) ? node3122 : node3117;
														assign node3117 = (inp[7]) ? 4'b0001 : node3118;
															assign node3118 = (inp[12]) ? 4'b0000 : 4'b1000;
														assign node3122 = (inp[7]) ? 4'b0000 : node3123;
															assign node3123 = (inp[12]) ? 4'b0001 : 4'b0000;
													assign node3127 = (inp[12]) ? node3133 : node3128;
														assign node3128 = (inp[10]) ? 4'b0001 : node3129;
															assign node3129 = (inp[7]) ? 4'b0000 : 4'b0001;
														assign node3133 = (inp[7]) ? node3137 : node3134;
															assign node3134 = (inp[10]) ? 4'b1000 : 4'b0001;
															assign node3137 = (inp[10]) ? 4'b0001 : 4'b0000;
										assign node3140 = (inp[11]) ? node3190 : node3141;
											assign node3141 = (inp[0]) ? node3171 : node3142;
												assign node3142 = (inp[12]) ? node3158 : node3143;
													assign node3143 = (inp[14]) ? node3153 : node3144;
														assign node3144 = (inp[7]) ? node3148 : node3145;
															assign node3145 = (inp[10]) ? 4'b0001 : 4'b1000;
															assign node3148 = (inp[10]) ? 4'b0000 : node3149;
																assign node3149 = (inp[2]) ? 4'b0001 : 4'b0000;
														assign node3153 = (inp[2]) ? node3155 : 4'b0001;
															assign node3155 = (inp[7]) ? 4'b0001 : 4'b0000;
													assign node3158 = (inp[7]) ? node3166 : node3159;
														assign node3159 = (inp[14]) ? node3163 : node3160;
															assign node3160 = (inp[10]) ? 4'b1000 : 4'b0000;
															assign node3163 = (inp[2]) ? 4'b0000 : 4'b0001;
														assign node3166 = (inp[2]) ? node3168 : 4'b0000;
															assign node3168 = (inp[14]) ? 4'b1000 : 4'b0000;
												assign node3171 = (inp[7]) ? node3183 : node3172;
													assign node3172 = (inp[10]) ? node3178 : node3173;
														assign node3173 = (inp[12]) ? 4'b0001 : node3174;
															assign node3174 = (inp[14]) ? 4'b1000 : 4'b1001;
														assign node3178 = (inp[14]) ? node3180 : 4'b0000;
															assign node3180 = (inp[2]) ? 4'b1000 : 4'b0000;
													assign node3183 = (inp[14]) ? 4'b0001 : node3184;
														assign node3184 = (inp[10]) ? 4'b0001 : node3185;
															assign node3185 = (inp[2]) ? 4'b1000 : 4'b0001;
											assign node3190 = (inp[10]) ? 4'b0001 : node3191;
												assign node3191 = (inp[2]) ? node3209 : node3192;
													assign node3192 = (inp[12]) ? node3198 : node3193;
														assign node3193 = (inp[0]) ? 4'b0001 : node3194;
															assign node3194 = (inp[7]) ? 4'b1001 : 4'b0001;
														assign node3198 = (inp[14]) ? node3204 : node3199;
															assign node3199 = (inp[7]) ? 4'b0001 : node3200;
																assign node3200 = (inp[0]) ? 4'b0001 : 4'b1001;
															assign node3204 = (inp[7]) ? node3206 : 4'b1001;
																assign node3206 = (inp[0]) ? 4'b1001 : 4'b0001;
													assign node3209 = (inp[0]) ? node3213 : node3210;
														assign node3210 = (inp[12]) ? 4'b0001 : 4'b1001;
														assign node3213 = (inp[14]) ? node3215 : 4'b1001;
															assign node3215 = (inp[7]) ? node3219 : node3216;
																assign node3216 = (inp[12]) ? 4'b1001 : 4'b0001;
																assign node3219 = (inp[12]) ? 4'b0001 : 4'b1001;
									assign node3223 = (inp[10]) ? node3305 : node3224;
										assign node3224 = (inp[1]) ? node3278 : node3225;
											assign node3225 = (inp[11]) ? node3257 : node3226;
												assign node3226 = (inp[14]) ? node3242 : node3227;
													assign node3227 = (inp[12]) ? node3237 : node3228;
														assign node3228 = (inp[2]) ? 4'b0000 : node3229;
															assign node3229 = (inp[0]) ? node3233 : node3230;
																assign node3230 = (inp[7]) ? 4'b0000 : 4'b0001;
																assign node3233 = (inp[7]) ? 4'b0001 : 4'b0000;
														assign node3237 = (inp[7]) ? node3239 : 4'b0000;
															assign node3239 = (inp[2]) ? 4'b0001 : 4'b0000;
													assign node3242 = (inp[7]) ? node3254 : node3243;
														assign node3243 = (inp[0]) ? node3249 : node3244;
															assign node3244 = (inp[12]) ? 4'b0000 : node3245;
																assign node3245 = (inp[2]) ? 4'b0000 : 4'b0001;
															assign node3249 = (inp[12]) ? 4'b0001 : node3250;
																assign node3250 = (inp[2]) ? 4'b0001 : 4'b0000;
														assign node3254 = (inp[0]) ? 4'b0000 : 4'b0001;
												assign node3257 = (inp[0]) ? node3265 : node3258;
													assign node3258 = (inp[7]) ? node3260 : 4'b0000;
														assign node3260 = (inp[12]) ? node3262 : 4'b0000;
															assign node3262 = (inp[2]) ? 4'b0001 : 4'b0000;
													assign node3265 = (inp[12]) ? node3273 : node3266;
														assign node3266 = (inp[2]) ? node3270 : node3267;
															assign node3267 = (inp[7]) ? 4'b0001 : 4'b0000;
															assign node3270 = (inp[7]) ? 4'b0000 : 4'b0001;
														assign node3273 = (inp[2]) ? 4'b0000 : node3274;
															assign node3274 = (inp[14]) ? 4'b0000 : 4'b0001;
											assign node3278 = (inp[11]) ? 4'b0001 : node3279;
												assign node3279 = (inp[0]) ? node3291 : node3280;
													assign node3280 = (inp[2]) ? node3286 : node3281;
														assign node3281 = (inp[14]) ? node3283 : 4'b0000;
															assign node3283 = (inp[7]) ? 4'b0001 : 4'b0000;
														assign node3286 = (inp[7]) ? 4'b0000 : node3287;
															assign node3287 = (inp[14]) ? 4'b0000 : 4'b0001;
													assign node3291 = (inp[14]) ? node3297 : node3292;
														assign node3292 = (inp[2]) ? node3294 : 4'b0001;
															assign node3294 = (inp[12]) ? 4'b0000 : 4'b0001;
														assign node3297 = (inp[2]) ? 4'b0001 : node3298;
															assign node3298 = (inp[7]) ? 4'b0000 : node3299;
																assign node3299 = (inp[12]) ? 4'b0001 : 4'b0000;
										assign node3305 = (inp[11]) ? 4'b0000 : node3306;
											assign node3306 = (inp[1]) ? 4'b0000 : node3307;
												assign node3307 = (inp[0]) ? node3325 : node3308;
													assign node3308 = (inp[7]) ? node3316 : node3309;
														assign node3309 = (inp[12]) ? 4'b0000 : node3310;
															assign node3310 = (inp[2]) ? 4'b0000 : node3311;
																assign node3311 = (inp[14]) ? 4'b0001 : 4'b0000;
														assign node3316 = (inp[2]) ? node3322 : node3317;
															assign node3317 = (inp[14]) ? 4'b0000 : node3318;
																assign node3318 = (inp[12]) ? 4'b0000 : 4'b0001;
															assign node3322 = (inp[12]) ? 4'b0001 : 4'b0000;
													assign node3325 = (inp[14]) ? node3335 : node3326;
														assign node3326 = (inp[2]) ? node3328 : 4'b0000;
															assign node3328 = (inp[12]) ? node3332 : node3329;
																assign node3329 = (inp[7]) ? 4'b0001 : 4'b0000;
																assign node3332 = (inp[7]) ? 4'b0000 : 4'b0001;
														assign node3335 = (inp[7]) ? node3337 : 4'b0001;
															assign node3337 = (inp[12]) ? 4'b0000 : node3338;
																assign node3338 = (inp[2]) ? 4'b0000 : 4'b0001;
				assign node3344 = (inp[6]) ? node3966 : node3345;
					assign node3345 = (inp[0]) ? 4'b1001 : node3346;
						assign node3346 = (inp[5]) ? node3474 : node3347;
							assign node3347 = (inp[2]) ? 4'b1011 : node3348;
								assign node3348 = (inp[3]) ? node3350 : 4'b1011;
									assign node3350 = (inp[7]) ? node3428 : node3351;
										assign node3351 = (inp[1]) ? node3389 : node3352;
											assign node3352 = (inp[11]) ? node3376 : node3353;
												assign node3353 = (inp[14]) ? node3361 : node3354;
													assign node3354 = (inp[4]) ? 4'b0000 : node3355;
														assign node3355 = (inp[13]) ? 4'b1000 : node3356;
															assign node3356 = (inp[10]) ? 4'b0000 : 4'b1011;
													assign node3361 = (inp[13]) ? node3371 : node3362;
														assign node3362 = (inp[4]) ? node3368 : node3363;
															assign node3363 = (inp[12]) ? 4'b1011 : node3364;
																assign node3364 = (inp[10]) ? 4'b0001 : 4'b1011;
															assign node3368 = (inp[12]) ? 4'b1001 : 4'b0001;
														assign node3371 = (inp[12]) ? 4'b0001 : node3372;
															assign node3372 = (inp[10]) ? 4'b1001 : 4'b0001;
												assign node3376 = (inp[13]) ? node3384 : node3377;
													assign node3377 = (inp[12]) ? node3379 : 4'b0000;
														assign node3379 = (inp[10]) ? 4'b0000 : node3380;
															assign node3380 = (inp[14]) ? 4'b1000 : 4'b1011;
													assign node3384 = (inp[10]) ? 4'b1000 : node3385;
														assign node3385 = (inp[12]) ? 4'b0000 : 4'b1000;
											assign node3389 = (inp[14]) ? node3403 : node3390;
												assign node3390 = (inp[13]) ? node3398 : node3391;
													assign node3391 = (inp[12]) ? node3393 : 4'b0001;
														assign node3393 = (inp[10]) ? 4'b0001 : node3394;
															assign node3394 = (inp[4]) ? 4'b1001 : 4'b1011;
													assign node3398 = (inp[10]) ? 4'b1001 : node3399;
														assign node3399 = (inp[12]) ? 4'b0001 : 4'b1001;
												assign node3403 = (inp[11]) ? node3415 : node3404;
													assign node3404 = (inp[13]) ? node3410 : node3405;
														assign node3405 = (inp[12]) ? node3407 : 4'b0000;
															assign node3407 = (inp[4]) ? 4'b1000 : 4'b1011;
														assign node3410 = (inp[10]) ? 4'b1000 : node3411;
															assign node3411 = (inp[12]) ? 4'b0000 : 4'b1000;
													assign node3415 = (inp[13]) ? node3423 : node3416;
														assign node3416 = (inp[10]) ? 4'b0001 : node3417;
															assign node3417 = (inp[4]) ? node3419 : 4'b1011;
																assign node3419 = (inp[12]) ? 4'b1001 : 4'b0001;
														assign node3423 = (inp[10]) ? 4'b1001 : node3424;
															assign node3424 = (inp[12]) ? 4'b0001 : 4'b1001;
										assign node3428 = (inp[4]) ? node3430 : 4'b1011;
											assign node3430 = (inp[13]) ? node3450 : node3431;
												assign node3431 = (inp[10]) ? node3441 : node3432;
													assign node3432 = (inp[12]) ? 4'b1011 : node3433;
														assign node3433 = (inp[14]) ? node3437 : node3434;
															assign node3434 = (inp[1]) ? 4'b0001 : 4'b0000;
															assign node3437 = (inp[1]) ? 4'b0000 : 4'b1011;
													assign node3441 = (inp[11]) ? 4'b0000 : node3442;
														assign node3442 = (inp[14]) ? node3446 : node3443;
															assign node3443 = (inp[1]) ? 4'b0001 : 4'b0000;
															assign node3446 = (inp[1]) ? 4'b0000 : 4'b1011;
												assign node3450 = (inp[1]) ? node3460 : node3451;
													assign node3451 = (inp[10]) ? node3455 : node3452;
														assign node3452 = (inp[12]) ? 4'b0000 : 4'b1000;
														assign node3455 = (inp[11]) ? 4'b1000 : node3456;
															assign node3456 = (inp[12]) ? 4'b1000 : 4'b1001;
													assign node3460 = (inp[10]) ? node3468 : node3461;
														assign node3461 = (inp[12]) ? node3463 : 4'b1001;
															assign node3463 = (inp[11]) ? 4'b0001 : node3464;
																assign node3464 = (inp[14]) ? 4'b0000 : 4'b0001;
														assign node3468 = (inp[11]) ? 4'b1001 : node3469;
															assign node3469 = (inp[14]) ? 4'b1000 : 4'b1001;
							assign node3474 = (inp[2]) ? node3822 : node3475;
								assign node3475 = (inp[1]) ? node3645 : node3476;
									assign node3476 = (inp[11]) ? node3582 : node3477;
										assign node3477 = (inp[14]) ? node3529 : node3478;
											assign node3478 = (inp[13]) ? node3502 : node3479;
												assign node3479 = (inp[12]) ? node3491 : node3480;
													assign node3480 = (inp[3]) ? node3486 : node3481;
														assign node3481 = (inp[7]) ? node3483 : 4'b0100;
															assign node3483 = (inp[10]) ? 4'b0100 : 4'b0000;
														assign node3486 = (inp[7]) ? node3488 : 4'b0000;
															assign node3488 = (inp[4]) ? 4'b0000 : 4'b0100;
													assign node3491 = (inp[10]) ? node3493 : 4'b1000;
														assign node3493 = (inp[4]) ? 4'b0000 : node3494;
															assign node3494 = (inp[7]) ? node3498 : node3495;
																assign node3495 = (inp[3]) ? 4'b0000 : 4'b0100;
																assign node3498 = (inp[3]) ? 4'b0100 : 4'b0000;
												assign node3502 = (inp[12]) ? node3514 : node3503;
													assign node3503 = (inp[3]) ? node3509 : node3504;
														assign node3504 = (inp[7]) ? node3506 : 4'b1100;
															assign node3506 = (inp[4]) ? 4'b1100 : 4'b1000;
														assign node3509 = (inp[7]) ? node3511 : 4'b1000;
															assign node3511 = (inp[4]) ? 4'b1000 : 4'b1100;
													assign node3514 = (inp[10]) ? node3522 : node3515;
														assign node3515 = (inp[4]) ? 4'b0000 : node3516;
															assign node3516 = (inp[7]) ? node3518 : 4'b0100;
																assign node3518 = (inp[3]) ? 4'b0100 : 4'b0000;
														assign node3522 = (inp[3]) ? 4'b1000 : node3523;
															assign node3523 = (inp[7]) ? node3525 : 4'b1100;
																assign node3525 = (inp[4]) ? 4'b1100 : 4'b1000;
											assign node3529 = (inp[13]) ? node3557 : node3530;
												assign node3530 = (inp[12]) ? node3546 : node3531;
													assign node3531 = (inp[10]) ? node3539 : node3532;
														assign node3532 = (inp[3]) ? node3536 : node3533;
															assign node3533 = (inp[4]) ? 4'b1101 : 4'b1001;
															assign node3536 = (inp[7]) ? 4'b1101 : 4'b1001;
														assign node3539 = (inp[3]) ? node3541 : 4'b0101;
															assign node3541 = (inp[4]) ? 4'b0001 : node3542;
																assign node3542 = (inp[7]) ? 4'b0101 : 4'b0001;
													assign node3546 = (inp[3]) ? node3552 : node3547;
														assign node3547 = (inp[7]) ? 4'b1001 : node3548;
															assign node3548 = (inp[4]) ? 4'b1101 : 4'b1001;
														assign node3552 = (inp[4]) ? node3554 : 4'b1101;
															assign node3554 = (inp[7]) ? 4'b1101 : 4'b1001;
												assign node3557 = (inp[3]) ? node3571 : node3558;
													assign node3558 = (inp[10]) ? node3564 : node3559;
														assign node3559 = (inp[4]) ? 4'b0101 : node3560;
															assign node3560 = (inp[7]) ? 4'b0001 : 4'b0101;
														assign node3564 = (inp[12]) ? 4'b0101 : node3565;
															assign node3565 = (inp[7]) ? node3567 : 4'b1101;
																assign node3567 = (inp[4]) ? 4'b1101 : 4'b1001;
													assign node3571 = (inp[12]) ? 4'b0001 : node3572;
														assign node3572 = (inp[10]) ? node3578 : node3573;
															assign node3573 = (inp[7]) ? node3575 : 4'b0001;
																assign node3575 = (inp[4]) ? 4'b0001 : 4'b0101;
															assign node3578 = (inp[7]) ? 4'b1101 : 4'b1001;
										assign node3582 = (inp[13]) ? node3614 : node3583;
											assign node3583 = (inp[10]) ? node3603 : node3584;
												assign node3584 = (inp[12]) ? node3592 : node3585;
													assign node3585 = (inp[3]) ? 4'b0000 : node3586;
														assign node3586 = (inp[7]) ? node3588 : 4'b0100;
															assign node3588 = (inp[4]) ? 4'b0100 : 4'b0000;
													assign node3592 = (inp[3]) ? node3598 : node3593;
														assign node3593 = (inp[7]) ? 4'b1000 : node3594;
															assign node3594 = (inp[4]) ? 4'b1100 : 4'b1000;
														assign node3598 = (inp[7]) ? 4'b1100 : node3599;
															assign node3599 = (inp[4]) ? 4'b1000 : 4'b1100;
												assign node3603 = (inp[3]) ? node3609 : node3604;
													assign node3604 = (inp[4]) ? 4'b0100 : node3605;
														assign node3605 = (inp[7]) ? 4'b0000 : 4'b0100;
													assign node3609 = (inp[7]) ? node3611 : 4'b0000;
														assign node3611 = (inp[4]) ? 4'b0000 : 4'b0100;
											assign node3614 = (inp[10]) ? node3634 : node3615;
												assign node3615 = (inp[12]) ? node3623 : node3616;
													assign node3616 = (inp[3]) ? node3618 : 4'b1100;
														assign node3618 = (inp[4]) ? 4'b1000 : node3619;
															assign node3619 = (inp[7]) ? 4'b1100 : 4'b1000;
													assign node3623 = (inp[3]) ? node3629 : node3624;
														assign node3624 = (inp[7]) ? node3626 : 4'b0100;
															assign node3626 = (inp[4]) ? 4'b0100 : 4'b0000;
														assign node3629 = (inp[4]) ? 4'b0000 : node3630;
															assign node3630 = (inp[7]) ? 4'b0100 : 4'b0000;
												assign node3634 = (inp[3]) ? node3640 : node3635;
													assign node3635 = (inp[4]) ? 4'b1100 : node3636;
														assign node3636 = (inp[7]) ? 4'b1000 : 4'b1100;
													assign node3640 = (inp[4]) ? 4'b1000 : node3641;
														assign node3641 = (inp[7]) ? 4'b1100 : 4'b1000;
									assign node3645 = (inp[14]) ? node3709 : node3646;
										assign node3646 = (inp[13]) ? node3674 : node3647;
											assign node3647 = (inp[10]) ? node3663 : node3648;
												assign node3648 = (inp[12]) ? node3656 : node3649;
													assign node3649 = (inp[3]) ? 4'b0001 : node3650;
														assign node3650 = (inp[7]) ? node3652 : 4'b0101;
															assign node3652 = (inp[4]) ? 4'b0101 : 4'b0001;
													assign node3656 = (inp[3]) ? node3658 : 4'b1001;
														assign node3658 = (inp[7]) ? 4'b1101 : node3659;
															assign node3659 = (inp[4]) ? 4'b1001 : 4'b1101;
												assign node3663 = (inp[3]) ? node3669 : node3664;
													assign node3664 = (inp[7]) ? node3666 : 4'b0101;
														assign node3666 = (inp[4]) ? 4'b0101 : 4'b0001;
													assign node3669 = (inp[7]) ? node3671 : 4'b0001;
														assign node3671 = (inp[4]) ? 4'b0001 : 4'b0101;
											assign node3674 = (inp[3]) ? node3692 : node3675;
												assign node3675 = (inp[4]) ? node3687 : node3676;
													assign node3676 = (inp[7]) ? node3682 : node3677;
														assign node3677 = (inp[10]) ? 4'b1101 : node3678;
															assign node3678 = (inp[12]) ? 4'b0101 : 4'b1101;
														assign node3682 = (inp[12]) ? node3684 : 4'b1001;
															assign node3684 = (inp[10]) ? 4'b1001 : 4'b0001;
													assign node3687 = (inp[10]) ? 4'b1101 : node3688;
														assign node3688 = (inp[12]) ? 4'b0101 : 4'b1101;
												assign node3692 = (inp[12]) ? node3698 : node3693;
													assign node3693 = (inp[4]) ? 4'b1001 : node3694;
														assign node3694 = (inp[7]) ? 4'b1101 : 4'b1001;
													assign node3698 = (inp[10]) ? node3704 : node3699;
														assign node3699 = (inp[4]) ? 4'b0001 : node3700;
															assign node3700 = (inp[7]) ? 4'b0101 : 4'b0001;
														assign node3704 = (inp[4]) ? 4'b1001 : node3705;
															assign node3705 = (inp[7]) ? 4'b1101 : 4'b1001;
										assign node3709 = (inp[11]) ? node3775 : node3710;
											assign node3710 = (inp[13]) ? node3742 : node3711;
												assign node3711 = (inp[10]) ? node3731 : node3712;
													assign node3712 = (inp[12]) ? node3722 : node3713;
														assign node3713 = (inp[3]) ? node3717 : node3714;
															assign node3714 = (inp[4]) ? 4'b0100 : 4'b0000;
															assign node3717 = (inp[4]) ? 4'b0000 : node3718;
																assign node3718 = (inp[7]) ? 4'b0100 : 4'b0000;
														assign node3722 = (inp[7]) ? node3728 : node3723;
															assign node3723 = (inp[3]) ? 4'b1000 : node3724;
																assign node3724 = (inp[4]) ? 4'b1100 : 4'b1000;
															assign node3728 = (inp[3]) ? 4'b1100 : 4'b1000;
													assign node3731 = (inp[3]) ? node3737 : node3732;
														assign node3732 = (inp[7]) ? node3734 : 4'b0100;
															assign node3734 = (inp[4]) ? 4'b0100 : 4'b0000;
														assign node3737 = (inp[7]) ? node3739 : 4'b0000;
															assign node3739 = (inp[4]) ? 4'b0000 : 4'b0100;
												assign node3742 = (inp[10]) ? node3764 : node3743;
													assign node3743 = (inp[12]) ? node3753 : node3744;
														assign node3744 = (inp[7]) ? node3748 : node3745;
															assign node3745 = (inp[3]) ? 4'b1000 : 4'b1100;
															assign node3748 = (inp[4]) ? 4'b1000 : node3749;
																assign node3749 = (inp[3]) ? 4'b1100 : 4'b1000;
														assign node3753 = (inp[3]) ? node3759 : node3754;
															assign node3754 = (inp[4]) ? 4'b0100 : node3755;
																assign node3755 = (inp[7]) ? 4'b0000 : 4'b0100;
															assign node3759 = (inp[4]) ? 4'b0000 : node3760;
																assign node3760 = (inp[7]) ? 4'b0100 : 4'b0000;
													assign node3764 = (inp[3]) ? node3770 : node3765;
														assign node3765 = (inp[4]) ? 4'b1100 : node3766;
															assign node3766 = (inp[7]) ? 4'b1000 : 4'b1100;
														assign node3770 = (inp[7]) ? node3772 : 4'b1000;
															assign node3772 = (inp[4]) ? 4'b1000 : 4'b1100;
											assign node3775 = (inp[13]) ? node3797 : node3776;
												assign node3776 = (inp[3]) ? node3788 : node3777;
													assign node3777 = (inp[4]) ? node3783 : node3778;
														assign node3778 = (inp[7]) ? 4'b0001 : node3779;
															assign node3779 = (inp[12]) ? 4'b1001 : 4'b0101;
														assign node3783 = (inp[10]) ? 4'b0101 : node3784;
															assign node3784 = (inp[12]) ? 4'b1101 : 4'b0101;
													assign node3788 = (inp[4]) ? 4'b0001 : node3789;
														assign node3789 = (inp[7]) ? 4'b0101 : node3790;
															assign node3790 = (inp[12]) ? node3792 : 4'b0001;
																assign node3792 = (inp[10]) ? 4'b0001 : 4'b1101;
												assign node3797 = (inp[12]) ? node3809 : node3798;
													assign node3798 = (inp[3]) ? node3804 : node3799;
														assign node3799 = (inp[4]) ? 4'b1101 : node3800;
															assign node3800 = (inp[7]) ? 4'b1001 : 4'b1101;
														assign node3804 = (inp[4]) ? 4'b1001 : node3805;
															assign node3805 = (inp[7]) ? 4'b1101 : 4'b1001;
													assign node3809 = (inp[10]) ? node3813 : node3810;
														assign node3810 = (inp[3]) ? 4'b0001 : 4'b0101;
														assign node3813 = (inp[7]) ? node3817 : node3814;
															assign node3814 = (inp[4]) ? 4'b1101 : 4'b1001;
															assign node3817 = (inp[4]) ? 4'b1001 : node3818;
																assign node3818 = (inp[3]) ? 4'b1101 : 4'b1001;
								assign node3822 = (inp[3]) ? node3824 : 4'b1011;
									assign node3824 = (inp[7]) ? node3906 : node3825;
										assign node3825 = (inp[1]) ? node3871 : node3826;
											assign node3826 = (inp[11]) ? node3858 : node3827;
												assign node3827 = (inp[14]) ? node3841 : node3828;
													assign node3828 = (inp[13]) ? node3836 : node3829;
														assign node3829 = (inp[10]) ? 4'b0000 : node3830;
															assign node3830 = (inp[4]) ? node3832 : 4'b1011;
																assign node3832 = (inp[12]) ? 4'b1000 : 4'b0000;
														assign node3836 = (inp[4]) ? node3838 : 4'b1000;
															assign node3838 = (inp[10]) ? 4'b1000 : 4'b0000;
													assign node3841 = (inp[4]) ? node3849 : node3842;
														assign node3842 = (inp[12]) ? 4'b1011 : node3843;
															assign node3843 = (inp[10]) ? node3845 : 4'b1011;
																assign node3845 = (inp[13]) ? 4'b1001 : 4'b0001;
														assign node3849 = (inp[13]) ? node3855 : node3850;
															assign node3850 = (inp[10]) ? node3852 : 4'b1001;
																assign node3852 = (inp[12]) ? 4'b1001 : 4'b0001;
															assign node3855 = (inp[10]) ? 4'b1001 : 4'b0001;
												assign node3858 = (inp[13]) ? node3866 : node3859;
													assign node3859 = (inp[10]) ? 4'b0000 : node3860;
														assign node3860 = (inp[12]) ? node3862 : 4'b0000;
															assign node3862 = (inp[4]) ? 4'b1000 : 4'b1011;
													assign node3866 = (inp[10]) ? 4'b1000 : node3867;
														assign node3867 = (inp[12]) ? 4'b0000 : 4'b1000;
											assign node3871 = (inp[14]) ? node3885 : node3872;
												assign node3872 = (inp[13]) ? node3880 : node3873;
													assign node3873 = (inp[12]) ? node3875 : 4'b0001;
														assign node3875 = (inp[10]) ? 4'b0001 : node3876;
															assign node3876 = (inp[4]) ? 4'b1001 : 4'b1011;
													assign node3880 = (inp[10]) ? 4'b1001 : node3881;
														assign node3881 = (inp[12]) ? 4'b0001 : 4'b1001;
												assign node3885 = (inp[11]) ? node3899 : node3886;
													assign node3886 = (inp[13]) ? node3894 : node3887;
														assign node3887 = (inp[10]) ? 4'b0000 : node3888;
															assign node3888 = (inp[12]) ? node3890 : 4'b0000;
																assign node3890 = (inp[4]) ? 4'b1000 : 4'b1011;
														assign node3894 = (inp[12]) ? node3896 : 4'b1000;
															assign node3896 = (inp[10]) ? 4'b1000 : 4'b0000;
													assign node3899 = (inp[13]) ? node3901 : 4'b0001;
														assign node3901 = (inp[12]) ? node3903 : 4'b1001;
															assign node3903 = (inp[10]) ? 4'b1001 : 4'b0001;
										assign node3906 = (inp[4]) ? node3908 : 4'b1011;
											assign node3908 = (inp[13]) ? node3936 : node3909;
												assign node3909 = (inp[10]) ? node3923 : node3910;
													assign node3910 = (inp[12]) ? 4'b1011 : node3911;
														assign node3911 = (inp[1]) ? node3917 : node3912;
															assign node3912 = (inp[14]) ? node3914 : 4'b0000;
																assign node3914 = (inp[11]) ? 4'b0000 : 4'b1011;
															assign node3917 = (inp[14]) ? node3919 : 4'b0001;
																assign node3919 = (inp[11]) ? 4'b0001 : 4'b0000;
													assign node3923 = (inp[1]) ? node3931 : node3924;
														assign node3924 = (inp[11]) ? 4'b0000 : node3925;
															assign node3925 = (inp[14]) ? node3927 : 4'b0000;
																assign node3927 = (inp[12]) ? 4'b1011 : 4'b0001;
														assign node3931 = (inp[11]) ? 4'b0001 : node3932;
															assign node3932 = (inp[14]) ? 4'b0000 : 4'b0001;
												assign node3936 = (inp[12]) ? node3948 : node3937;
													assign node3937 = (inp[1]) ? node3943 : node3938;
														assign node3938 = (inp[11]) ? 4'b1000 : node3939;
															assign node3939 = (inp[10]) ? 4'b1000 : 4'b0001;
														assign node3943 = (inp[11]) ? 4'b1001 : node3944;
															assign node3944 = (inp[14]) ? 4'b1000 : 4'b1001;
													assign node3948 = (inp[10]) ? node3958 : node3949;
														assign node3949 = (inp[14]) ? node3951 : 4'b0001;
															assign node3951 = (inp[11]) ? node3955 : node3952;
																assign node3952 = (inp[1]) ? 4'b0000 : 4'b0001;
																assign node3955 = (inp[1]) ? 4'b0001 : 4'b0000;
														assign node3958 = (inp[14]) ? node3962 : node3959;
															assign node3959 = (inp[1]) ? 4'b1001 : 4'b1000;
															assign node3962 = (inp[1]) ? 4'b1001 : 4'b0001;
					assign node3966 = (inp[0]) ? node5598 : node3967;
						assign node3967 = (inp[5]) ? node4777 : node3968;
							assign node3968 = (inp[11]) ? node4464 : node3969;
								assign node3969 = (inp[2]) ? node4185 : node3970;
									assign node3970 = (inp[4]) ? node4092 : node3971;
										assign node3971 = (inp[7]) ? node4033 : node3972;
											assign node3972 = (inp[3]) ? node4020 : node3973;
												assign node3973 = (inp[13]) ? node3993 : node3974;
													assign node3974 = (inp[10]) ? node3984 : node3975;
														assign node3975 = (inp[1]) ? node3981 : node3976;
															assign node3976 = (inp[14]) ? 4'b1001 : node3977;
																assign node3977 = (inp[12]) ? 4'b1000 : 4'b0100;
															assign node3981 = (inp[14]) ? 4'b0100 : 4'b0101;
														assign node3984 = (inp[12]) ? node3990 : node3985;
															assign node3985 = (inp[1]) ? 4'b0100 : node3986;
																assign node3986 = (inp[14]) ? 4'b0101 : 4'b0100;
															assign node3990 = (inp[1]) ? 4'b0101 : 4'b0100;
													assign node3993 = (inp[10]) ? node4007 : node3994;
														assign node3994 = (inp[12]) ? node4000 : node3995;
															assign node3995 = (inp[14]) ? 4'b0101 : node3996;
																assign node3996 = (inp[1]) ? 4'b1101 : 4'b1100;
															assign node4000 = (inp[14]) ? node4004 : node4001;
																assign node4001 = (inp[1]) ? 4'b0101 : 4'b0100;
																assign node4004 = (inp[1]) ? 4'b0100 : 4'b0101;
														assign node4007 = (inp[12]) ? node4015 : node4008;
															assign node4008 = (inp[1]) ? node4012 : node4009;
																assign node4009 = (inp[14]) ? 4'b1101 : 4'b1100;
																assign node4012 = (inp[14]) ? 4'b1100 : 4'b1101;
															assign node4015 = (inp[1]) ? node4017 : 4'b1100;
																assign node4017 = (inp[14]) ? 4'b1100 : 4'b1101;
												assign node4020 = (inp[10]) ? node4028 : node4021;
													assign node4021 = (inp[1]) ? 4'b0100 : node4022;
														assign node4022 = (inp[12]) ? node4024 : 4'b0100;
															assign node4024 = (inp[13]) ? 4'b1100 : 4'b1000;
													assign node4028 = (inp[12]) ? node4030 : 4'b1100;
														assign node4030 = (inp[1]) ? 4'b1100 : 4'b0100;
											assign node4033 = (inp[3]) ? node4071 : node4034;
												assign node4034 = (inp[13]) ? node4052 : node4035;
													assign node4035 = (inp[10]) ? node4045 : node4036;
														assign node4036 = (inp[14]) ? node4042 : node4037;
															assign node4037 = (inp[12]) ? 4'b1001 : node4038;
																assign node4038 = (inp[1]) ? 4'b0001 : 4'b0000;
															assign node4042 = (inp[1]) ? 4'b1000 : 4'b1001;
														assign node4045 = (inp[1]) ? node4049 : node4046;
															assign node4046 = (inp[14]) ? 4'b0001 : 4'b0000;
															assign node4049 = (inp[14]) ? 4'b0000 : 4'b0001;
													assign node4052 = (inp[10]) ? node4060 : node4053;
														assign node4053 = (inp[1]) ? node4057 : node4054;
															assign node4054 = (inp[14]) ? 4'b0001 : 4'b0000;
															assign node4057 = (inp[14]) ? 4'b1000 : 4'b1001;
														assign node4060 = (inp[12]) ? node4066 : node4061;
															assign node4061 = (inp[1]) ? node4063 : 4'b1001;
																assign node4063 = (inp[14]) ? 4'b1000 : 4'b1001;
															assign node4066 = (inp[1]) ? node4068 : 4'b1000;
																assign node4068 = (inp[14]) ? 4'b1000 : 4'b1001;
												assign node4071 = (inp[13]) ? node4083 : node4072;
													assign node4072 = (inp[10]) ? node4078 : node4073;
														assign node4073 = (inp[12]) ? node4075 : 4'b0000;
															assign node4075 = (inp[1]) ? 4'b0000 : 4'b1000;
														assign node4078 = (inp[1]) ? 4'b1000 : node4079;
															assign node4079 = (inp[12]) ? 4'b0000 : 4'b1000;
													assign node4083 = (inp[1]) ? node4089 : node4084;
														assign node4084 = (inp[10]) ? node4086 : 4'b1000;
															assign node4086 = (inp[12]) ? 4'b0100 : 4'b1100;
														assign node4089 = (inp[10]) ? 4'b1100 : 4'b0100;
										assign node4092 = (inp[13]) ? node4146 : node4093;
											assign node4093 = (inp[7]) ? node4113 : node4094;
												assign node4094 = (inp[10]) ? node4102 : node4095;
													assign node4095 = (inp[1]) ? 4'b0000 : node4096;
														assign node4096 = (inp[12]) ? node4098 : 4'b0000;
															assign node4098 = (inp[3]) ? 4'b1100 : 4'b1101;
													assign node4102 = (inp[3]) ? node4108 : node4103;
														assign node4103 = (inp[1]) ? 4'b1000 : node4104;
															assign node4104 = (inp[12]) ? 4'b0000 : 4'b1000;
														assign node4108 = (inp[1]) ? 4'b0001 : node4109;
															assign node4109 = (inp[12]) ? 4'b0000 : 4'b1000;
												assign node4113 = (inp[3]) ? node4135 : node4114;
													assign node4114 = (inp[10]) ? node4128 : node4115;
														assign node4115 = (inp[12]) ? node4123 : node4116;
															assign node4116 = (inp[14]) ? node4120 : node4117;
																assign node4117 = (inp[1]) ? 4'b0101 : 4'b0100;
																assign node4120 = (inp[1]) ? 4'b0100 : 4'b1001;
															assign node4123 = (inp[14]) ? node4125 : 4'b1000;
																assign node4125 = (inp[1]) ? 4'b1000 : 4'b1001;
														assign node4128 = (inp[1]) ? node4132 : node4129;
															assign node4129 = (inp[14]) ? 4'b0101 : 4'b0100;
															assign node4132 = (inp[14]) ? 4'b0100 : 4'b0101;
													assign node4135 = (inp[10]) ? node4141 : node4136;
														assign node4136 = (inp[1]) ? 4'b0100 : node4137;
															assign node4137 = (inp[12]) ? 4'b1100 : 4'b0100;
														assign node4141 = (inp[1]) ? 4'b1100 : node4142;
															assign node4142 = (inp[12]) ? 4'b0100 : 4'b1100;
											assign node4146 = (inp[10]) ? node4170 : node4147;
												assign node4147 = (inp[12]) ? node4157 : node4148;
													assign node4148 = (inp[7]) ? 4'b0000 : node4149;
														assign node4149 = (inp[3]) ? node4151 : 4'b0000;
															assign node4151 = (inp[14]) ? node4153 : 4'b0000;
																assign node4153 = (inp[1]) ? 4'b1001 : 4'b1000;
													assign node4157 = (inp[1]) ? 4'b0000 : node4158;
														assign node4158 = (inp[7]) ? node4164 : node4159;
															assign node4159 = (inp[3]) ? node4161 : 4'b1000;
																assign node4161 = (inp[14]) ? 4'b0000 : 4'b0001;
															assign node4164 = (inp[3]) ? 4'b1100 : node4165;
																assign node4165 = (inp[14]) ? 4'b0101 : 4'b0100;
												assign node4170 = (inp[1]) ? node4178 : node4171;
													assign node4171 = (inp[3]) ? node4175 : node4172;
														assign node4172 = (inp[12]) ? 4'b0000 : 4'b1000;
														assign node4175 = (inp[14]) ? 4'b0000 : 4'b0001;
													assign node4178 = (inp[14]) ? node4180 : 4'b1000;
														assign node4180 = (inp[3]) ? node4182 : 4'b1000;
															assign node4182 = (inp[12]) ? 4'b0001 : 4'b1001;
									assign node4185 = (inp[3]) ? node4337 : node4186;
										assign node4186 = (inp[4]) ? node4270 : node4187;
											assign node4187 = (inp[7]) ? node4239 : node4188;
												assign node4188 = (inp[13]) ? node4214 : node4189;
													assign node4189 = (inp[10]) ? node4201 : node4190;
														assign node4190 = (inp[12]) ? node4196 : node4191;
															assign node4191 = (inp[14]) ? 4'b1001 : node4192;
																assign node4192 = (inp[1]) ? 4'b0101 : 4'b0100;
															assign node4196 = (inp[14]) ? 4'b1001 : node4197;
																assign node4197 = (inp[1]) ? 4'b1001 : 4'b1000;
														assign node4201 = (inp[12]) ? node4209 : node4202;
															assign node4202 = (inp[14]) ? node4206 : node4203;
																assign node4203 = (inp[1]) ? 4'b0101 : 4'b0100;
																assign node4206 = (inp[1]) ? 4'b0100 : 4'b0101;
															assign node4209 = (inp[1]) ? 4'b0100 : node4210;
																assign node4210 = (inp[14]) ? 4'b1001 : 4'b0100;
													assign node4214 = (inp[12]) ? node4224 : node4215;
														assign node4215 = (inp[10]) ? node4219 : node4216;
															assign node4216 = (inp[14]) ? 4'b1100 : 4'b1101;
															assign node4219 = (inp[1]) ? 4'b1101 : node4220;
																assign node4220 = (inp[14]) ? 4'b1101 : 4'b1100;
														assign node4224 = (inp[10]) ? node4232 : node4225;
															assign node4225 = (inp[1]) ? node4229 : node4226;
																assign node4226 = (inp[14]) ? 4'b0101 : 4'b0100;
																assign node4229 = (inp[14]) ? 4'b0100 : 4'b0101;
															assign node4232 = (inp[1]) ? node4236 : node4233;
																assign node4233 = (inp[14]) ? 4'b0101 : 4'b1100;
																assign node4236 = (inp[14]) ? 4'b1100 : 4'b1101;
												assign node4239 = (inp[13]) ? node4255 : node4240;
													assign node4240 = (inp[12]) ? node4246 : node4241;
														assign node4241 = (inp[1]) ? node4243 : 4'b0000;
															assign node4243 = (inp[14]) ? 4'b0000 : 4'b0001;
														assign node4246 = (inp[10]) ? node4252 : node4247;
															assign node4247 = (inp[1]) ? node4249 : 4'b1001;
																assign node4249 = (inp[14]) ? 4'b1000 : 4'b1001;
															assign node4252 = (inp[14]) ? 4'b0000 : 4'b0001;
													assign node4255 = (inp[1]) ? node4263 : node4256;
														assign node4256 = (inp[14]) ? 4'b0001 : node4257;
															assign node4257 = (inp[10]) ? 4'b1000 : node4258;
																assign node4258 = (inp[12]) ? 4'b0000 : 4'b1000;
														assign node4263 = (inp[14]) ? node4265 : 4'b1001;
															assign node4265 = (inp[10]) ? 4'b1000 : node4266;
																assign node4266 = (inp[12]) ? 4'b0000 : 4'b1000;
											assign node4270 = (inp[13]) ? node4306 : node4271;
												assign node4271 = (inp[12]) ? node4287 : node4272;
													assign node4272 = (inp[7]) ? node4280 : node4273;
														assign node4273 = (inp[14]) ? node4277 : node4274;
															assign node4274 = (inp[1]) ? 4'b0101 : 4'b0100;
															assign node4277 = (inp[1]) ? 4'b0100 : 4'b0101;
														assign node4280 = (inp[1]) ? node4284 : node4281;
															assign node4281 = (inp[14]) ? 4'b1001 : 4'b0100;
															assign node4284 = (inp[14]) ? 4'b0100 : 4'b0101;
													assign node4287 = (inp[10]) ? node4297 : node4288;
														assign node4288 = (inp[7]) ? 4'b1000 : node4289;
															assign node4289 = (inp[1]) ? node4293 : node4290;
																assign node4290 = (inp[14]) ? 4'b1101 : 4'b1100;
																assign node4293 = (inp[14]) ? 4'b1100 : 4'b1101;
														assign node4297 = (inp[1]) ? node4303 : node4298;
															assign node4298 = (inp[14]) ? node4300 : 4'b0100;
																assign node4300 = (inp[7]) ? 4'b1001 : 4'b1101;
															assign node4303 = (inp[14]) ? 4'b0100 : 4'b0101;
												assign node4306 = (inp[12]) ? node4322 : node4307;
													assign node4307 = (inp[7]) ? node4315 : node4308;
														assign node4308 = (inp[14]) ? node4312 : node4309;
															assign node4309 = (inp[1]) ? 4'b1101 : 4'b1100;
															assign node4312 = (inp[1]) ? 4'b1100 : 4'b0101;
														assign node4315 = (inp[14]) ? node4319 : node4316;
															assign node4316 = (inp[1]) ? 4'b1101 : 4'b1100;
															assign node4319 = (inp[1]) ? 4'b1100 : 4'b1101;
													assign node4322 = (inp[10]) ? node4330 : node4323;
														assign node4323 = (inp[1]) ? node4327 : node4324;
															assign node4324 = (inp[14]) ? 4'b0101 : 4'b0100;
															assign node4327 = (inp[14]) ? 4'b0100 : 4'b0101;
														assign node4330 = (inp[1]) ? node4334 : node4331;
															assign node4331 = (inp[14]) ? 4'b0101 : 4'b1100;
															assign node4334 = (inp[14]) ? 4'b1100 : 4'b1101;
										assign node4337 = (inp[4]) ? node4413 : node4338;
											assign node4338 = (inp[7]) ? node4388 : node4339;
												assign node4339 = (inp[13]) ? node4361 : node4340;
													assign node4340 = (inp[10]) ? node4354 : node4341;
														assign node4341 = (inp[12]) ? node4347 : node4342;
															assign node4342 = (inp[1]) ? node4344 : 4'b1101;
																assign node4344 = (inp[14]) ? 4'b0000 : 4'b0001;
															assign node4347 = (inp[14]) ? node4351 : node4348;
																assign node4348 = (inp[1]) ? 4'b1101 : 4'b1100;
																assign node4351 = (inp[1]) ? 4'b1100 : 4'b1101;
														assign node4354 = (inp[14]) ? node4358 : node4355;
															assign node4355 = (inp[1]) ? 4'b0001 : 4'b0000;
															assign node4358 = (inp[1]) ? 4'b0000 : 4'b1101;
													assign node4361 = (inp[12]) ? node4375 : node4362;
														assign node4362 = (inp[10]) ? node4368 : node4363;
															assign node4363 = (inp[14]) ? 4'b1000 : node4364;
																assign node4364 = (inp[1]) ? 4'b1001 : 4'b1000;
															assign node4368 = (inp[14]) ? node4372 : node4369;
																assign node4369 = (inp[1]) ? 4'b1001 : 4'b1000;
																assign node4372 = (inp[1]) ? 4'b1000 : 4'b1001;
														assign node4375 = (inp[10]) ? node4383 : node4376;
															assign node4376 = (inp[1]) ? node4380 : node4377;
																assign node4377 = (inp[14]) ? 4'b0001 : 4'b0000;
																assign node4380 = (inp[14]) ? 4'b0000 : 4'b0001;
															assign node4383 = (inp[1]) ? 4'b1000 : node4384;
																assign node4384 = (inp[14]) ? 4'b0001 : 4'b1000;
												assign node4388 = (inp[13]) ? node4404 : node4389;
													assign node4389 = (inp[1]) ? node4397 : node4390;
														assign node4390 = (inp[14]) ? node4392 : 4'b1100;
															assign node4392 = (inp[12]) ? 4'b1101 : node4393;
																assign node4393 = (inp[10]) ? 4'b0101 : 4'b1101;
														assign node4397 = (inp[14]) ? 4'b0100 : node4398;
															assign node4398 = (inp[10]) ? 4'b0101 : node4399;
																assign node4399 = (inp[12]) ? 4'b1101 : 4'b0101;
													assign node4404 = (inp[1]) ? node4410 : node4405;
														assign node4405 = (inp[10]) ? 4'b1101 : node4406;
															assign node4406 = (inp[14]) ? 4'b0101 : 4'b0100;
														assign node4410 = (inp[14]) ? 4'b1100 : 4'b1101;
											assign node4413 = (inp[7]) ? node4429 : node4414;
												assign node4414 = (inp[10]) ? node4424 : node4415;
													assign node4415 = (inp[12]) ? node4417 : 4'b0000;
														assign node4417 = (inp[1]) ? 4'b0000 : node4418;
															assign node4418 = (inp[13]) ? 4'b1000 : node4419;
																assign node4419 = (inp[14]) ? 4'b1001 : 4'b1000;
													assign node4424 = (inp[1]) ? 4'b1000 : node4425;
														assign node4425 = (inp[12]) ? 4'b0000 : 4'b1000;
												assign node4429 = (inp[13]) ? node4455 : node4430;
													assign node4430 = (inp[12]) ? node4444 : node4431;
														assign node4431 = (inp[10]) ? node4437 : node4432;
															assign node4432 = (inp[1]) ? 4'b0000 : node4433;
																assign node4433 = (inp[14]) ? 4'b1101 : 4'b0000;
															assign node4437 = (inp[14]) ? node4441 : node4438;
																assign node4438 = (inp[1]) ? 4'b0001 : 4'b0000;
																assign node4441 = (inp[1]) ? 4'b0000 : 4'b0001;
														assign node4444 = (inp[10]) ? node4452 : node4445;
															assign node4445 = (inp[14]) ? node4449 : node4446;
																assign node4446 = (inp[1]) ? 4'b1101 : 4'b1100;
																assign node4449 = (inp[1]) ? 4'b1100 : 4'b1101;
															assign node4452 = (inp[1]) ? 4'b0000 : 4'b1101;
													assign node4455 = (inp[10]) ? node4461 : node4456;
														assign node4456 = (inp[1]) ? 4'b0000 : node4457;
															assign node4457 = (inp[12]) ? 4'b0001 : 4'b0000;
														assign node4461 = (inp[12]) ? 4'b0000 : 4'b1000;
								assign node4464 = (inp[1]) ? node4628 : node4465;
									assign node4465 = (inp[3]) ? node4535 : node4466;
										assign node4466 = (inp[7]) ? node4502 : node4467;
											assign node4467 = (inp[2]) ? node4489 : node4468;
												assign node4468 = (inp[4]) ? node4480 : node4469;
													assign node4469 = (inp[13]) ? node4475 : node4470;
														assign node4470 = (inp[12]) ? node4472 : 4'b0100;
															assign node4472 = (inp[10]) ? 4'b0100 : 4'b1000;
														assign node4475 = (inp[12]) ? node4477 : 4'b1100;
															assign node4477 = (inp[10]) ? 4'b1100 : 4'b0100;
													assign node4480 = (inp[10]) ? node4486 : node4481;
														assign node4481 = (inp[12]) ? node4483 : 4'b0001;
															assign node4483 = (inp[13]) ? 4'b1001 : 4'b1100;
														assign node4486 = (inp[12]) ? 4'b0001 : 4'b1001;
												assign node4489 = (inp[13]) ? node4497 : node4490;
													assign node4490 = (inp[12]) ? node4492 : 4'b0100;
														assign node4492 = (inp[10]) ? 4'b0100 : node4493;
															assign node4493 = (inp[4]) ? 4'b1100 : 4'b1000;
													assign node4497 = (inp[10]) ? 4'b1100 : node4498;
														assign node4498 = (inp[12]) ? 4'b0100 : 4'b1100;
											assign node4502 = (inp[4]) ? node4514 : node4503;
												assign node4503 = (inp[13]) ? node4509 : node4504;
													assign node4504 = (inp[10]) ? 4'b0000 : node4505;
														assign node4505 = (inp[12]) ? 4'b1000 : 4'b0000;
													assign node4509 = (inp[10]) ? 4'b1000 : node4510;
														assign node4510 = (inp[12]) ? 4'b0000 : 4'b1000;
												assign node4514 = (inp[2]) ? node4526 : node4515;
													assign node4515 = (inp[13]) ? node4519 : node4516;
														assign node4516 = (inp[12]) ? 4'b1000 : 4'b0100;
														assign node4519 = (inp[12]) ? node4523 : node4520;
															assign node4520 = (inp[10]) ? 4'b1001 : 4'b0001;
															assign node4523 = (inp[10]) ? 4'b0001 : 4'b0100;
													assign node4526 = (inp[13]) ? node4532 : node4527;
														assign node4527 = (inp[10]) ? 4'b0100 : node4528;
															assign node4528 = (inp[12]) ? 4'b1000 : 4'b0100;
														assign node4532 = (inp[10]) ? 4'b1100 : 4'b0100;
										assign node4535 = (inp[2]) ? node4589 : node4536;
											assign node4536 = (inp[4]) ? node4556 : node4537;
												assign node4537 = (inp[13]) ? node4549 : node4538;
													assign node4538 = (inp[7]) ? node4544 : node4539;
														assign node4539 = (inp[12]) ? 4'b1001 : node4540;
															assign node4540 = (inp[10]) ? 4'b1101 : 4'b0101;
														assign node4544 = (inp[12]) ? 4'b1001 : node4545;
															assign node4545 = (inp[10]) ? 4'b1001 : 4'b0001;
													assign node4549 = (inp[10]) ? node4553 : node4550;
														assign node4550 = (inp[12]) ? 4'b1101 : 4'b0101;
														assign node4553 = (inp[12]) ? 4'b0101 : 4'b1101;
												assign node4556 = (inp[7]) ? node4570 : node4557;
													assign node4557 = (inp[13]) ? node4565 : node4558;
														assign node4558 = (inp[10]) ? node4562 : node4559;
															assign node4559 = (inp[12]) ? 4'b1101 : 4'b0001;
															assign node4562 = (inp[12]) ? 4'b0001 : 4'b0000;
														assign node4565 = (inp[12]) ? node4567 : 4'b1000;
															assign node4567 = (inp[10]) ? 4'b0000 : 4'b1000;
													assign node4570 = (inp[13]) ? node4584 : node4571;
														assign node4571 = (inp[14]) ? node4577 : node4572;
															assign node4572 = (inp[10]) ? node4574 : 4'b1101;
																assign node4574 = (inp[12]) ? 4'b0101 : 4'b1101;
															assign node4577 = (inp[10]) ? node4581 : node4578;
																assign node4578 = (inp[12]) ? 4'b1101 : 4'b0101;
																assign node4581 = (inp[12]) ? 4'b0101 : 4'b1101;
														assign node4584 = (inp[12]) ? 4'b1101 : node4585;
															assign node4585 = (inp[10]) ? 4'b1000 : 4'b0001;
											assign node4589 = (inp[4]) ? node4611 : node4590;
												assign node4590 = (inp[7]) ? node4600 : node4591;
													assign node4591 = (inp[12]) ? node4595 : node4592;
														assign node4592 = (inp[13]) ? 4'b1000 : 4'b0000;
														assign node4595 = (inp[13]) ? 4'b0000 : node4596;
															assign node4596 = (inp[10]) ? 4'b0000 : 4'b1100;
													assign node4600 = (inp[13]) ? node4606 : node4601;
														assign node4601 = (inp[10]) ? 4'b0100 : node4602;
															assign node4602 = (inp[12]) ? 4'b1100 : 4'b0100;
														assign node4606 = (inp[12]) ? node4608 : 4'b1100;
															assign node4608 = (inp[10]) ? 4'b1100 : 4'b0100;
												assign node4611 = (inp[12]) ? node4619 : node4612;
													assign node4612 = (inp[10]) ? node4614 : 4'b0001;
														assign node4614 = (inp[7]) ? node4616 : 4'b1001;
															assign node4616 = (inp[13]) ? 4'b1001 : 4'b0000;
													assign node4619 = (inp[10]) ? node4623 : node4620;
														assign node4620 = (inp[7]) ? 4'b0000 : 4'b1000;
														assign node4623 = (inp[7]) ? node4625 : 4'b0001;
															assign node4625 = (inp[13]) ? 4'b0001 : 4'b0000;
									assign node4628 = (inp[13]) ? node4720 : node4629;
										assign node4629 = (inp[12]) ? node4667 : node4630;
											assign node4630 = (inp[3]) ? node4642 : node4631;
												assign node4631 = (inp[7]) ? node4639 : node4632;
													assign node4632 = (inp[4]) ? node4634 : 4'b0101;
														assign node4634 = (inp[2]) ? 4'b0101 : node4635;
															assign node4635 = (inp[10]) ? 4'b1001 : 4'b0001;
													assign node4639 = (inp[4]) ? 4'b0101 : 4'b0001;
												assign node4642 = (inp[10]) ? node4654 : node4643;
													assign node4643 = (inp[7]) ? node4649 : node4644;
														assign node4644 = (inp[4]) ? 4'b0001 : node4645;
															assign node4645 = (inp[2]) ? 4'b0001 : 4'b0101;
														assign node4649 = (inp[14]) ? node4651 : 4'b0101;
															assign node4651 = (inp[4]) ? 4'b0101 : 4'b0001;
													assign node4654 = (inp[2]) ? node4660 : node4655;
														assign node4655 = (inp[7]) ? node4657 : 4'b0001;
															assign node4657 = (inp[4]) ? 4'b1101 : 4'b1001;
														assign node4660 = (inp[7]) ? node4664 : node4661;
															assign node4661 = (inp[4]) ? 4'b1001 : 4'b0001;
															assign node4664 = (inp[4]) ? 4'b0001 : 4'b0101;
											assign node4667 = (inp[10]) ? node4695 : node4668;
												assign node4668 = (inp[3]) ? node4676 : node4669;
													assign node4669 = (inp[4]) ? node4671 : 4'b1001;
														assign node4671 = (inp[2]) ? node4673 : 4'b0001;
															assign node4673 = (inp[7]) ? 4'b1001 : 4'b1101;
													assign node4676 = (inp[2]) ? node4690 : node4677;
														assign node4677 = (inp[14]) ? node4683 : node4678;
															assign node4678 = (inp[4]) ? node4680 : 4'b0101;
																assign node4680 = (inp[7]) ? 4'b0101 : 4'b0001;
															assign node4683 = (inp[4]) ? node4687 : node4684;
																assign node4684 = (inp[7]) ? 4'b0001 : 4'b0101;
																assign node4687 = (inp[7]) ? 4'b0101 : 4'b0001;
														assign node4690 = (inp[4]) ? node4692 : 4'b1101;
															assign node4692 = (inp[7]) ? 4'b1101 : 4'b0001;
												assign node4695 = (inp[3]) ? node4705 : node4696;
													assign node4696 = (inp[4]) ? node4700 : node4697;
														assign node4697 = (inp[7]) ? 4'b0001 : 4'b0101;
														assign node4700 = (inp[7]) ? 4'b0101 : node4701;
															assign node4701 = (inp[2]) ? 4'b0101 : 4'b1001;
													assign node4705 = (inp[2]) ? node4713 : node4706;
														assign node4706 = (inp[14]) ? node4708 : 4'b1101;
															assign node4708 = (inp[7]) ? node4710 : 4'b0001;
																assign node4710 = (inp[4]) ? 4'b1101 : 4'b1001;
														assign node4713 = (inp[4]) ? node4717 : node4714;
															assign node4714 = (inp[7]) ? 4'b0101 : 4'b0001;
															assign node4717 = (inp[7]) ? 4'b0001 : 4'b1001;
										assign node4720 = (inp[10]) ? node4762 : node4721;
											assign node4721 = (inp[12]) ? node4741 : node4722;
												assign node4722 = (inp[4]) ? node4736 : node4723;
													assign node4723 = (inp[2]) ? node4729 : node4724;
														assign node4724 = (inp[3]) ? 4'b0101 : node4725;
															assign node4725 = (inp[7]) ? 4'b1001 : 4'b1101;
														assign node4729 = (inp[7]) ? node4733 : node4730;
															assign node4730 = (inp[3]) ? 4'b1001 : 4'b1101;
															assign node4733 = (inp[3]) ? 4'b1101 : 4'b1001;
													assign node4736 = (inp[3]) ? 4'b0001 : node4737;
														assign node4737 = (inp[2]) ? 4'b1101 : 4'b0001;
												assign node4741 = (inp[4]) ? node4751 : node4742;
													assign node4742 = (inp[3]) ? node4746 : node4743;
														assign node4743 = (inp[7]) ? 4'b0001 : 4'b0101;
														assign node4746 = (inp[7]) ? 4'b0101 : node4747;
															assign node4747 = (inp[2]) ? 4'b0001 : 4'b0101;
													assign node4751 = (inp[3]) ? node4755 : node4752;
														assign node4752 = (inp[2]) ? 4'b0101 : 4'b0001;
														assign node4755 = (inp[14]) ? 4'b0001 : node4756;
															assign node4756 = (inp[2]) ? 4'b0001 : node4757;
																assign node4757 = (inp[7]) ? 4'b0001 : 4'b1001;
											assign node4762 = (inp[4]) ? node4772 : node4763;
												assign node4763 = (inp[7]) ? node4769 : node4764;
													assign node4764 = (inp[3]) ? node4766 : 4'b1101;
														assign node4766 = (inp[2]) ? 4'b1001 : 4'b1101;
													assign node4769 = (inp[3]) ? 4'b1101 : 4'b1001;
												assign node4772 = (inp[2]) ? node4774 : 4'b1001;
													assign node4774 = (inp[3]) ? 4'b1001 : 4'b1101;
							assign node4777 = (inp[3]) ? node5175 : node4778;
								assign node4778 = (inp[4]) ? node4984 : node4779;
									assign node4779 = (inp[11]) ? node4899 : node4780;
										assign node4780 = (inp[2]) ? node4856 : node4781;
											assign node4781 = (inp[13]) ? node4825 : node4782;
												assign node4782 = (inp[7]) ? node4806 : node4783;
													assign node4783 = (inp[1]) ? node4795 : node4784;
														assign node4784 = (inp[14]) ? node4788 : node4785;
															assign node4785 = (inp[10]) ? 4'b1101 : 4'b1001;
															assign node4788 = (inp[12]) ? node4792 : node4789;
																assign node4789 = (inp[10]) ? 4'b1100 : 4'b0100;
																assign node4792 = (inp[10]) ? 4'b1100 : 4'b1000;
														assign node4795 = (inp[14]) ? node4801 : node4796;
															assign node4796 = (inp[10]) ? 4'b0100 : node4797;
																assign node4797 = (inp[12]) ? 4'b0100 : 4'b1100;
															assign node4801 = (inp[12]) ? node4803 : 4'b0101;
																assign node4803 = (inp[10]) ? 4'b1101 : 4'b0101;
													assign node4806 = (inp[10]) ? node4818 : node4807;
														assign node4807 = (inp[14]) ? node4815 : node4808;
															assign node4808 = (inp[1]) ? node4812 : node4809;
																assign node4809 = (inp[12]) ? 4'b1001 : 4'b0001;
																assign node4812 = (inp[12]) ? 4'b0000 : 4'b1000;
															assign node4815 = (inp[1]) ? 4'b0001 : 4'b0000;
														assign node4818 = (inp[14]) ? node4820 : 4'b0100;
															assign node4820 = (inp[1]) ? node4822 : 4'b1000;
																assign node4822 = (inp[12]) ? 4'b1001 : 4'b0101;
												assign node4825 = (inp[10]) ? node4845 : node4826;
													assign node4826 = (inp[7]) ? node4834 : node4827;
														assign node4827 = (inp[14]) ? node4831 : node4828;
															assign node4828 = (inp[12]) ? 4'b0101 : 4'b0001;
															assign node4831 = (inp[12]) ? 4'b0001 : 4'b1001;
														assign node4834 = (inp[1]) ? node4840 : node4835;
															assign node4835 = (inp[14]) ? 4'b0100 : node4836;
																assign node4836 = (inp[12]) ? 4'b0101 : 4'b1101;
															assign node4840 = (inp[14]) ? 4'b1101 : node4841;
																assign node4841 = (inp[12]) ? 4'b1100 : 4'b0100;
													assign node4845 = (inp[14]) ? node4847 : 4'b0001;
														assign node4847 = (inp[12]) ? node4851 : node4848;
															assign node4848 = (inp[1]) ? 4'b1001 : 4'b0001;
															assign node4851 = (inp[7]) ? 4'b0100 : node4852;
																assign node4852 = (inp[1]) ? 4'b0001 : 4'b1001;
											assign node4856 = (inp[10]) ? node4874 : node4857;
												assign node4857 = (inp[1]) ? node4869 : node4858;
													assign node4858 = (inp[12]) ? node4864 : node4859;
														assign node4859 = (inp[13]) ? 4'b0100 : node4860;
															assign node4860 = (inp[7]) ? 4'b0000 : 4'b0100;
														assign node4864 = (inp[13]) ? node4866 : 4'b1000;
															assign node4866 = (inp[7]) ? 4'b1000 : 4'b1100;
													assign node4869 = (inp[13]) ? 4'b0100 : node4870;
														assign node4870 = (inp[7]) ? 4'b0000 : 4'b0100;
												assign node4874 = (inp[1]) ? node4892 : node4875;
													assign node4875 = (inp[12]) ? node4885 : node4876;
														assign node4876 = (inp[13]) ? node4880 : node4877;
															assign node4877 = (inp[7]) ? 4'b1000 : 4'b1100;
															assign node4880 = (inp[7]) ? 4'b1100 : node4881;
																assign node4881 = (inp[14]) ? 4'b0000 : 4'b0001;
														assign node4885 = (inp[14]) ? 4'b0100 : node4886;
															assign node4886 = (inp[13]) ? 4'b0001 : node4887;
																assign node4887 = (inp[7]) ? 4'b0000 : 4'b0100;
													assign node4892 = (inp[7]) ? node4896 : node4893;
														assign node4893 = (inp[13]) ? 4'b1000 : 4'b1100;
														assign node4896 = (inp[13]) ? 4'b1100 : 4'b1000;
										assign node4899 = (inp[1]) ? node4947 : node4900;
											assign node4900 = (inp[2]) ? node4916 : node4901;
												assign node4901 = (inp[13]) ? node4911 : node4902;
													assign node4902 = (inp[7]) ? node4906 : node4903;
														assign node4903 = (inp[10]) ? 4'b1100 : 4'b0100;
														assign node4906 = (inp[10]) ? node4908 : 4'b0000;
															assign node4908 = (inp[12]) ? 4'b1000 : 4'b0100;
													assign node4911 = (inp[10]) ? 4'b0001 : node4912;
														assign node4912 = (inp[7]) ? 4'b1100 : 4'b0001;
												assign node4916 = (inp[7]) ? node4930 : node4917;
													assign node4917 = (inp[13]) ? node4923 : node4918;
														assign node4918 = (inp[10]) ? node4920 : 4'b1001;
															assign node4920 = (inp[12]) ? 4'b0101 : 4'b1101;
														assign node4923 = (inp[10]) ? node4927 : node4924;
															assign node4924 = (inp[12]) ? 4'b1101 : 4'b0101;
															assign node4927 = (inp[12]) ? 4'b0000 : 4'b1000;
													assign node4930 = (inp[13]) ? node4940 : node4931;
														assign node4931 = (inp[14]) ? 4'b1001 : node4932;
															assign node4932 = (inp[12]) ? node4936 : node4933;
																assign node4933 = (inp[10]) ? 4'b1001 : 4'b0001;
																assign node4936 = (inp[10]) ? 4'b0001 : 4'b1001;
														assign node4940 = (inp[12]) ? node4944 : node4941;
															assign node4941 = (inp[10]) ? 4'b1101 : 4'b0101;
															assign node4944 = (inp[10]) ? 4'b0101 : 4'b1001;
											assign node4947 = (inp[13]) ? node4967 : node4948;
												assign node4948 = (inp[7]) ? node4958 : node4949;
													assign node4949 = (inp[10]) ? node4955 : node4950;
														assign node4950 = (inp[12]) ? 4'b0101 : node4951;
															assign node4951 = (inp[2]) ? 4'b0101 : 4'b1101;
														assign node4955 = (inp[2]) ? 4'b1101 : 4'b0101;
													assign node4958 = (inp[10]) ? node4964 : node4959;
														assign node4959 = (inp[12]) ? 4'b0001 : node4960;
															assign node4960 = (inp[2]) ? 4'b0001 : 4'b1001;
														assign node4964 = (inp[2]) ? 4'b1001 : 4'b0101;
												assign node4967 = (inp[7]) ? node4975 : node4968;
													assign node4968 = (inp[2]) ? node4970 : 4'b1001;
														assign node4970 = (inp[10]) ? 4'b1001 : node4971;
															assign node4971 = (inp[12]) ? 4'b0101 : 4'b0001;
													assign node4975 = (inp[10]) ? node4981 : node4976;
														assign node4976 = (inp[2]) ? 4'b0101 : node4977;
															assign node4977 = (inp[12]) ? 4'b1101 : 4'b0101;
														assign node4981 = (inp[2]) ? 4'b1101 : 4'b1001;
									assign node4984 = (inp[1]) ? node5092 : node4985;
										assign node4985 = (inp[12]) ? node5029 : node4986;
											assign node4986 = (inp[2]) ? node5010 : node4987;
												assign node4987 = (inp[13]) ? node4995 : node4988;
													assign node4988 = (inp[10]) ? node4992 : node4989;
														assign node4989 = (inp[7]) ? 4'b0001 : 4'b0101;
														assign node4992 = (inp[7]) ? 4'b0101 : 4'b1000;
													assign node4995 = (inp[11]) ? node5005 : node4996;
														assign node4996 = (inp[14]) ? node5002 : node4997;
															assign node4997 = (inp[10]) ? node4999 : 4'b1000;
																assign node4999 = (inp[7]) ? 4'b0100 : 4'b1000;
															assign node5002 = (inp[10]) ? 4'b1000 : 4'b1001;
														assign node5005 = (inp[10]) ? 4'b0001 : node5006;
															assign node5006 = (inp[7]) ? 4'b0000 : 4'b0100;
												assign node5010 = (inp[13]) ? node5022 : node5011;
													assign node5011 = (inp[10]) ? node5017 : node5012;
														assign node5012 = (inp[14]) ? 4'b0000 : node5013;
															assign node5013 = (inp[11]) ? 4'b0000 : 4'b0001;
														assign node5017 = (inp[11]) ? 4'b0000 : node5018;
															assign node5018 = (inp[14]) ? 4'b1000 : 4'b1001;
													assign node5022 = (inp[7]) ? node5024 : 4'b0001;
														assign node5024 = (inp[10]) ? 4'b0001 : node5025;
															assign node5025 = (inp[11]) ? 4'b1000 : 4'b1001;
											assign node5029 = (inp[13]) ? node5057 : node5030;
												assign node5030 = (inp[11]) ? node5048 : node5031;
													assign node5031 = (inp[2]) ? node5037 : node5032;
														assign node5032 = (inp[10]) ? node5034 : 4'b1001;
															assign node5034 = (inp[7]) ? 4'b1001 : 4'b0001;
														assign node5037 = (inp[14]) ? node5043 : node5038;
															assign node5038 = (inp[7]) ? node5040 : 4'b1001;
																assign node5040 = (inp[10]) ? 4'b1001 : 4'b1100;
															assign node5043 = (inp[7]) ? node5045 : 4'b1000;
																assign node5045 = (inp[10]) ? 4'b1000 : 4'b1100;
													assign node5048 = (inp[14]) ? node5052 : node5049;
														assign node5049 = (inp[10]) ? 4'b1000 : 4'b0000;
														assign node5052 = (inp[10]) ? node5054 : 4'b0101;
															assign node5054 = (inp[7]) ? 4'b0101 : 4'b1000;
												assign node5057 = (inp[2]) ? node5075 : node5058;
													assign node5058 = (inp[14]) ? node5068 : node5059;
														assign node5059 = (inp[7]) ? node5063 : node5060;
															assign node5060 = (inp[11]) ? 4'b1001 : 4'b1000;
															assign node5063 = (inp[10]) ? node5065 : 4'b1000;
																assign node5065 = (inp[11]) ? 4'b0100 : 4'b1000;
														assign node5068 = (inp[11]) ? 4'b1000 : node5069;
															assign node5069 = (inp[10]) ? node5071 : 4'b0001;
																assign node5071 = (inp[7]) ? 4'b1001 : 4'b1000;
													assign node5075 = (inp[11]) ? 4'b0001 : node5076;
														assign node5076 = (inp[14]) ? node5084 : node5077;
															assign node5077 = (inp[7]) ? node5081 : node5078;
																assign node5078 = (inp[10]) ? 4'b1001 : 4'b0101;
																assign node5081 = (inp[10]) ? 4'b0101 : 4'b0001;
															assign node5084 = (inp[7]) ? node5088 : node5085;
																assign node5085 = (inp[10]) ? 4'b1001 : 4'b0100;
																assign node5088 = (inp[10]) ? 4'b0100 : 4'b0000;
										assign node5092 = (inp[11]) ? node5146 : node5093;
											assign node5093 = (inp[12]) ? node5119 : node5094;
												assign node5094 = (inp[13]) ? node5110 : node5095;
													assign node5095 = (inp[10]) ? node5101 : node5096;
														assign node5096 = (inp[2]) ? node5098 : 4'b1101;
															assign node5098 = (inp[14]) ? 4'b0001 : 4'b1000;
														assign node5101 = (inp[2]) ? node5105 : node5102;
															assign node5102 = (inp[14]) ? 4'b0000 : 4'b0001;
															assign node5105 = (inp[14]) ? 4'b0101 : node5106;
																assign node5106 = (inp[7]) ? 4'b0000 : 4'b0100;
													assign node5110 = (inp[2]) ? 4'b1001 : node5111;
														assign node5111 = (inp[10]) ? 4'b1000 : node5112;
															assign node5112 = (inp[7]) ? node5114 : 4'b0000;
																assign node5114 = (inp[14]) ? 4'b0000 : 4'b0001;
												assign node5119 = (inp[13]) ? node5133 : node5120;
													assign node5120 = (inp[2]) ? node5128 : node5121;
														assign node5121 = (inp[14]) ? 4'b0101 : node5122;
															assign node5122 = (inp[7]) ? node5124 : 4'b1001;
																assign node5124 = (inp[10]) ? 4'b0101 : 4'b0001;
														assign node5128 = (inp[14]) ? 4'b0001 : node5129;
															assign node5129 = (inp[7]) ? 4'b0000 : 4'b0100;
													assign node5133 = (inp[2]) ? node5139 : node5134;
														assign node5134 = (inp[10]) ? 4'b0000 : node5135;
															assign node5135 = (inp[7]) ? 4'b0001 : 4'b0101;
														assign node5139 = (inp[7]) ? node5141 : 4'b0001;
															assign node5141 = (inp[14]) ? node5143 : 4'b1000;
																assign node5143 = (inp[10]) ? 4'b0001 : 4'b1001;
											assign node5146 = (inp[13]) ? node5166 : node5147;
												assign node5147 = (inp[10]) ? node5161 : node5148;
													assign node5148 = (inp[7]) ? node5156 : node5149;
														assign node5149 = (inp[12]) ? node5153 : node5150;
															assign node5150 = (inp[2]) ? 4'b1001 : 4'b0001;
															assign node5153 = (inp[2]) ? 4'b0001 : 4'b1101;
														assign node5156 = (inp[2]) ? node5158 : 4'b1001;
															assign node5158 = (inp[14]) ? 4'b1001 : 4'b0001;
													assign node5161 = (inp[7]) ? 4'b0001 : node5162;
														assign node5162 = (inp[2]) ? 4'b0101 : 4'b0001;
												assign node5166 = (inp[10]) ? 4'b1001 : node5167;
													assign node5167 = (inp[2]) ? node5169 : 4'b0001;
														assign node5169 = (inp[12]) ? 4'b1001 : node5170;
															assign node5170 = (inp[7]) ? 4'b0101 : 4'b1001;
								assign node5175 = (inp[4]) ? node5407 : node5176;
									assign node5176 = (inp[1]) ? node5308 : node5177;
										assign node5177 = (inp[10]) ? node5243 : node5178;
											assign node5178 = (inp[7]) ? node5214 : node5179;
												assign node5179 = (inp[2]) ? node5203 : node5180;
													assign node5180 = (inp[12]) ? node5192 : node5181;
														assign node5181 = (inp[14]) ? node5187 : node5182;
															assign node5182 = (inp[13]) ? node5184 : 4'b0001;
																assign node5184 = (inp[11]) ? 4'b0001 : 4'b0000;
															assign node5187 = (inp[13]) ? node5189 : 4'b1000;
																assign node5189 = (inp[11]) ? 4'b0001 : 4'b1001;
														assign node5192 = (inp[11]) ? node5200 : node5193;
															assign node5193 = (inp[13]) ? node5197 : node5194;
																assign node5194 = (inp[14]) ? 4'b0000 : 4'b0001;
																assign node5197 = (inp[14]) ? 4'b1001 : 4'b1000;
															assign node5200 = (inp[13]) ? 4'b0000 : 4'b1000;
													assign node5203 = (inp[13]) ? 4'b0000 : node5204;
														assign node5204 = (inp[11]) ? node5210 : node5205;
															assign node5205 = (inp[14]) ? node5207 : 4'b0000;
																assign node5207 = (inp[12]) ? 4'b1001 : 4'b0001;
															assign node5210 = (inp[12]) ? 4'b0000 : 4'b1000;
												assign node5214 = (inp[11]) ? node5228 : node5215;
													assign node5215 = (inp[2]) ? node5223 : node5216;
														assign node5216 = (inp[13]) ? node5218 : 4'b0000;
															assign node5218 = (inp[12]) ? 4'b0001 : node5219;
																assign node5219 = (inp[14]) ? 4'b0001 : 4'b0000;
														assign node5223 = (inp[13]) ? 4'b0000 : node5224;
															assign node5224 = (inp[12]) ? 4'b1001 : 4'b0001;
													assign node5228 = (inp[12]) ? node5238 : node5229;
														assign node5229 = (inp[14]) ? node5233 : node5230;
															assign node5230 = (inp[2]) ? 4'b0001 : 4'b1001;
															assign node5233 = (inp[13]) ? node5235 : 4'b1001;
																assign node5235 = (inp[2]) ? 4'b1001 : 4'b1000;
														assign node5238 = (inp[13]) ? node5240 : 4'b0001;
															assign node5240 = (inp[2]) ? 4'b0001 : 4'b0000;
											assign node5243 = (inp[7]) ? node5271 : node5244;
												assign node5244 = (inp[11]) ? node5256 : node5245;
													assign node5245 = (inp[2]) ? node5251 : node5246;
														assign node5246 = (inp[13]) ? node5248 : 4'b0001;
															assign node5248 = (inp[14]) ? 4'b1000 : 4'b1001;
														assign node5251 = (inp[13]) ? 4'b0001 : node5252;
															assign node5252 = (inp[14]) ? 4'b0001 : 4'b1000;
													assign node5256 = (inp[12]) ? node5264 : node5257;
														assign node5257 = (inp[13]) ? node5261 : node5258;
															assign node5258 = (inp[2]) ? 4'b0001 : 4'b1001;
															assign node5261 = (inp[2]) ? 4'b1001 : 4'b0001;
														assign node5264 = (inp[13]) ? node5268 : node5265;
															assign node5265 = (inp[2]) ? 4'b1000 : 4'b1001;
															assign node5268 = (inp[2]) ? 4'b1001 : 4'b0001;
												assign node5271 = (inp[11]) ? node5289 : node5272;
													assign node5272 = (inp[13]) ? node5282 : node5273;
														assign node5273 = (inp[14]) ? node5279 : node5274;
															assign node5274 = (inp[2]) ? node5276 : 4'b0001;
																assign node5276 = (inp[12]) ? 4'b0000 : 4'b1000;
															assign node5279 = (inp[2]) ? 4'b0001 : 4'b0000;
														assign node5282 = (inp[2]) ? node5286 : node5283;
															assign node5283 = (inp[12]) ? 4'b1000 : 4'b0000;
															assign node5286 = (inp[14]) ? 4'b1000 : 4'b1001;
													assign node5289 = (inp[13]) ? node5295 : node5290;
														assign node5290 = (inp[12]) ? node5292 : 4'b1000;
															assign node5292 = (inp[2]) ? 4'b1000 : 4'b0000;
														assign node5295 = (inp[14]) ? node5301 : node5296;
															assign node5296 = (inp[2]) ? node5298 : 4'b0000;
																assign node5298 = (inp[12]) ? 4'b1000 : 4'b0000;
															assign node5301 = (inp[12]) ? node5305 : node5302;
																assign node5302 = (inp[2]) ? 4'b0000 : 4'b1000;
																assign node5305 = (inp[2]) ? 4'b1000 : 4'b0000;
										assign node5308 = (inp[11]) ? node5364 : node5309;
											assign node5309 = (inp[10]) ? node5335 : node5310;
												assign node5310 = (inp[13]) ? node5320 : node5311;
													assign node5311 = (inp[2]) ? 4'b1001 : node5312;
														assign node5312 = (inp[14]) ? node5314 : 4'b0000;
															assign node5314 = (inp[12]) ? node5316 : 4'b0001;
																assign node5316 = (inp[7]) ? 4'b1000 : 4'b1001;
													assign node5320 = (inp[12]) ? node5326 : node5321;
														assign node5321 = (inp[7]) ? node5323 : 4'b1000;
															assign node5323 = (inp[2]) ? 4'b0000 : 4'b0001;
														assign node5326 = (inp[2]) ? node5332 : node5327;
															assign node5327 = (inp[7]) ? node5329 : 4'b1000;
																assign node5329 = (inp[14]) ? 4'b1000 : 4'b1001;
															assign node5332 = (inp[7]) ? 4'b1000 : 4'b0001;
												assign node5335 = (inp[7]) ? node5351 : node5336;
													assign node5336 = (inp[2]) ? node5344 : node5337;
														assign node5337 = (inp[14]) ? node5339 : 4'b0001;
															assign node5339 = (inp[12]) ? node5341 : 4'b0000;
																assign node5341 = (inp[13]) ? 4'b1001 : 4'b0001;
														assign node5344 = (inp[13]) ? node5348 : node5345;
															assign node5345 = (inp[12]) ? 4'b0000 : 4'b1000;
															assign node5348 = (inp[14]) ? 4'b0000 : 4'b0001;
													assign node5351 = (inp[12]) ? node5353 : 4'b0001;
														assign node5353 = (inp[14]) ? node5359 : node5354;
															assign node5354 = (inp[13]) ? 4'b0000 : node5355;
																assign node5355 = (inp[2]) ? 4'b1001 : 4'b0001;
															assign node5359 = (inp[13]) ? node5361 : 4'b0001;
																assign node5361 = (inp[2]) ? 4'b0001 : 4'b1001;
											assign node5364 = (inp[10]) ? node5392 : node5365;
												assign node5365 = (inp[13]) ? node5387 : node5366;
													assign node5366 = (inp[14]) ? node5374 : node5367;
														assign node5367 = (inp[7]) ? node5369 : 4'b0001;
															assign node5369 = (inp[12]) ? node5371 : 4'b0001;
																assign node5371 = (inp[2]) ? 4'b1001 : 4'b0001;
														assign node5374 = (inp[7]) ? node5380 : node5375;
															assign node5375 = (inp[12]) ? 4'b1001 : node5376;
																assign node5376 = (inp[2]) ? 4'b0001 : 4'b1001;
															assign node5380 = (inp[2]) ? node5384 : node5381;
																assign node5381 = (inp[12]) ? 4'b0001 : 4'b1001;
																assign node5384 = (inp[12]) ? 4'b1001 : 4'b0001;
													assign node5387 = (inp[2]) ? node5389 : 4'b0001;
														assign node5389 = (inp[12]) ? 4'b1001 : 4'b0001;
												assign node5392 = (inp[13]) ? 4'b1001 : node5393;
													assign node5393 = (inp[14]) ? node5399 : node5394;
														assign node5394 = (inp[7]) ? node5396 : 4'b1001;
															assign node5396 = (inp[2]) ? 4'b0001 : 4'b1001;
														assign node5399 = (inp[2]) ? node5403 : node5400;
															assign node5400 = (inp[7]) ? 4'b1001 : 4'b0001;
															assign node5403 = (inp[7]) ? 4'b0001 : 4'b1001;
									assign node5407 = (inp[13]) ? node5523 : node5408;
										assign node5408 = (inp[10]) ? node5474 : node5409;
											assign node5409 = (inp[1]) ? node5439 : node5410;
												assign node5410 = (inp[7]) ? node5418 : node5411;
													assign node5411 = (inp[2]) ? node5413 : 4'b1000;
														assign node5413 = (inp[11]) ? 4'b0000 : node5414;
															assign node5414 = (inp[12]) ? 4'b0000 : 4'b1000;
													assign node5418 = (inp[14]) ? node5430 : node5419;
														assign node5419 = (inp[11]) ? node5423 : node5420;
															assign node5420 = (inp[2]) ? 4'b0000 : 4'b1000;
															assign node5423 = (inp[12]) ? node5427 : node5424;
																assign node5424 = (inp[2]) ? 4'b0001 : 4'b1001;
																assign node5427 = (inp[2]) ? 4'b1000 : 4'b0001;
														assign node5430 = (inp[11]) ? node5436 : node5431;
															assign node5431 = (inp[12]) ? 4'b0001 : node5432;
																assign node5432 = (inp[2]) ? 4'b0001 : 4'b1001;
															assign node5436 = (inp[2]) ? 4'b1000 : 4'b0001;
												assign node5439 = (inp[11]) ? node5463 : node5440;
													assign node5440 = (inp[7]) ? node5452 : node5441;
														assign node5441 = (inp[12]) ? node5447 : node5442;
															assign node5442 = (inp[14]) ? node5444 : 4'b0001;
																assign node5444 = (inp[2]) ? 4'b0001 : 4'b0000;
															assign node5447 = (inp[14]) ? 4'b1001 : node5448;
																assign node5448 = (inp[2]) ? 4'b1000 : 4'b1001;
														assign node5452 = (inp[2]) ? node5458 : node5453;
															assign node5453 = (inp[14]) ? node5455 : 4'b1000;
																assign node5455 = (inp[12]) ? 4'b0001 : 4'b1001;
															assign node5458 = (inp[12]) ? 4'b1000 : node5459;
																assign node5459 = (inp[14]) ? 4'b1000 : 4'b0000;
													assign node5463 = (inp[12]) ? node5469 : node5464;
														assign node5464 = (inp[7]) ? node5466 : 4'b0001;
															assign node5466 = (inp[2]) ? 4'b1001 : 4'b0001;
														assign node5469 = (inp[7]) ? node5471 : 4'b1001;
															assign node5471 = (inp[2]) ? 4'b0001 : 4'b1001;
											assign node5474 = (inp[1]) ? node5504 : node5475;
												assign node5475 = (inp[7]) ? node5489 : node5476;
													assign node5476 = (inp[2]) ? node5484 : node5477;
														assign node5477 = (inp[12]) ? node5479 : 4'b0001;
															assign node5479 = (inp[11]) ? 4'b1000 : node5480;
																assign node5480 = (inp[14]) ? 4'b1000 : 4'b1001;
														assign node5484 = (inp[12]) ? 4'b0000 : node5485;
															assign node5485 = (inp[11]) ? 4'b1000 : 4'b0000;
													assign node5489 = (inp[11]) ? node5499 : node5490;
														assign node5490 = (inp[12]) ? node5496 : node5491;
															assign node5491 = (inp[2]) ? node5493 : 4'b1000;
																assign node5493 = (inp[14]) ? 4'b1001 : 4'b0000;
															assign node5496 = (inp[2]) ? 4'b0001 : 4'b0000;
														assign node5499 = (inp[12]) ? node5501 : 4'b0001;
															assign node5501 = (inp[2]) ? 4'b1000 : 4'b0001;
												assign node5504 = (inp[11]) ? 4'b0001 : node5505;
													assign node5505 = (inp[7]) ? node5511 : node5506;
														assign node5506 = (inp[2]) ? node5508 : 4'b0001;
															assign node5508 = (inp[14]) ? 4'b0000 : 4'b0001;
														assign node5511 = (inp[12]) ? node5517 : node5512;
															assign node5512 = (inp[14]) ? 4'b1000 : node5513;
																assign node5513 = (inp[2]) ? 4'b1000 : 4'b0000;
															assign node5517 = (inp[14]) ? node5519 : 4'b0000;
																assign node5519 = (inp[2]) ? 4'b0001 : 4'b0000;
										assign node5523 = (inp[10]) ? node5577 : node5524;
											assign node5524 = (inp[1]) ? node5562 : node5525;
												assign node5525 = (inp[2]) ? node5547 : node5526;
													assign node5526 = (inp[7]) ? node5538 : node5527;
														assign node5527 = (inp[12]) ? node5533 : node5528;
															assign node5528 = (inp[14]) ? 4'b0000 : node5529;
																assign node5529 = (inp[11]) ? 4'b0000 : 4'b0001;
															assign node5533 = (inp[11]) ? 4'b0001 : node5534;
																assign node5534 = (inp[14]) ? 4'b0000 : 4'b0001;
														assign node5538 = (inp[12]) ? node5544 : node5539;
															assign node5539 = (inp[14]) ? 4'b0001 : node5540;
																assign node5540 = (inp[11]) ? 4'b0001 : 4'b0000;
															assign node5544 = (inp[11]) ? 4'b0000 : 4'b0001;
													assign node5547 = (inp[12]) ? node5555 : node5548;
														assign node5548 = (inp[14]) ? 4'b0001 : node5549;
															assign node5549 = (inp[7]) ? node5551 : 4'b0000;
																assign node5551 = (inp[11]) ? 4'b0000 : 4'b0001;
														assign node5555 = (inp[7]) ? node5557 : 4'b0000;
															assign node5557 = (inp[11]) ? 4'b0000 : node5558;
																assign node5558 = (inp[14]) ? 4'b0000 : 4'b0001;
												assign node5562 = (inp[11]) ? 4'b0001 : node5563;
													assign node5563 = (inp[14]) ? node5571 : node5564;
														assign node5564 = (inp[2]) ? 4'b0000 : node5565;
															assign node5565 = (inp[7]) ? 4'b0001 : node5566;
																assign node5566 = (inp[12]) ? 4'b0000 : 4'b0001;
														assign node5571 = (inp[7]) ? node5573 : 4'b0001;
															assign node5573 = (inp[2]) ? 4'b0001 : 4'b0000;
											assign node5577 = (inp[11]) ? 4'b0000 : node5578;
												assign node5578 = (inp[1]) ? 4'b0000 : node5579;
													assign node5579 = (inp[12]) ? node5587 : node5580;
														assign node5580 = (inp[2]) ? 4'b0001 : node5581;
															assign node5581 = (inp[7]) ? node5583 : 4'b0000;
																assign node5583 = (inp[14]) ? 4'b0001 : 4'b0000;
														assign node5587 = (inp[2]) ? 4'b0000 : node5588;
															assign node5588 = (inp[7]) ? node5592 : node5589;
																assign node5589 = (inp[14]) ? 4'b0001 : 4'b0000;
																assign node5592 = (inp[14]) ? 4'b0000 : 4'b0001;
						assign node5598 = (inp[5]) ? node5726 : node5599;
							assign node5599 = (inp[2]) ? 4'b1001 : node5600;
								assign node5600 = (inp[3]) ? node5602 : 4'b1001;
									assign node5602 = (inp[7]) ? node5670 : node5603;
										assign node5603 = (inp[1]) ? node5641 : node5604;
											assign node5604 = (inp[14]) ? node5618 : node5605;
												assign node5605 = (inp[13]) ? node5613 : node5606;
													assign node5606 = (inp[12]) ? node5608 : 4'b0000;
														assign node5608 = (inp[10]) ? 4'b0000 : node5609;
															assign node5609 = (inp[4]) ? 4'b1000 : 4'b1001;
													assign node5613 = (inp[12]) ? node5615 : 4'b1000;
														assign node5615 = (inp[10]) ? 4'b1000 : 4'b0000;
												assign node5618 = (inp[11]) ? node5630 : node5619;
													assign node5619 = (inp[13]) ? node5625 : node5620;
														assign node5620 = (inp[10]) ? node5622 : 4'b1001;
															assign node5622 = (inp[12]) ? 4'b1001 : 4'b0001;
														assign node5625 = (inp[10]) ? node5627 : 4'b0001;
															assign node5627 = (inp[12]) ? 4'b0001 : 4'b1001;
													assign node5630 = (inp[13]) ? node5636 : node5631;
														assign node5631 = (inp[12]) ? node5633 : 4'b0000;
															assign node5633 = (inp[10]) ? 4'b0000 : 4'b1000;
														assign node5636 = (inp[10]) ? 4'b1000 : node5637;
															assign node5637 = (inp[12]) ? 4'b0000 : 4'b1000;
											assign node5641 = (inp[13]) ? node5657 : node5642;
												assign node5642 = (inp[10]) ? node5652 : node5643;
													assign node5643 = (inp[12]) ? node5645 : 4'b0001;
														assign node5645 = (inp[14]) ? node5647 : 4'b1001;
															assign node5647 = (inp[11]) ? 4'b1001 : node5648;
																assign node5648 = (inp[4]) ? 4'b1000 : 4'b1001;
													assign node5652 = (inp[14]) ? node5654 : 4'b0001;
														assign node5654 = (inp[11]) ? 4'b0001 : 4'b0000;
												assign node5657 = (inp[11]) ? node5665 : node5658;
													assign node5658 = (inp[14]) ? node5660 : 4'b1001;
														assign node5660 = (inp[10]) ? 4'b1000 : node5661;
															assign node5661 = (inp[12]) ? 4'b0000 : 4'b1000;
													assign node5665 = (inp[12]) ? node5667 : 4'b1001;
														assign node5667 = (inp[10]) ? 4'b1001 : 4'b0001;
										assign node5670 = (inp[4]) ? node5672 : 4'b1001;
											assign node5672 = (inp[13]) ? node5696 : node5673;
												assign node5673 = (inp[10]) ? node5687 : node5674;
													assign node5674 = (inp[12]) ? 4'b1001 : node5675;
														assign node5675 = (inp[1]) ? node5681 : node5676;
															assign node5676 = (inp[14]) ? node5678 : 4'b0000;
																assign node5678 = (inp[11]) ? 4'b0000 : 4'b1001;
															assign node5681 = (inp[14]) ? node5683 : 4'b0001;
																assign node5683 = (inp[11]) ? 4'b0001 : 4'b0000;
													assign node5687 = (inp[1]) ? 4'b0001 : node5688;
														assign node5688 = (inp[11]) ? 4'b0000 : node5689;
															assign node5689 = (inp[14]) ? node5691 : 4'b0000;
																assign node5691 = (inp[12]) ? 4'b1001 : 4'b0001;
												assign node5696 = (inp[10]) ? node5716 : node5697;
													assign node5697 = (inp[12]) ? node5709 : node5698;
														assign node5698 = (inp[1]) ? node5704 : node5699;
															assign node5699 = (inp[14]) ? node5701 : 4'b1000;
																assign node5701 = (inp[11]) ? 4'b1000 : 4'b0001;
															assign node5704 = (inp[11]) ? 4'b1001 : node5705;
																assign node5705 = (inp[14]) ? 4'b1000 : 4'b1001;
														assign node5709 = (inp[14]) ? node5711 : 4'b0001;
															assign node5711 = (inp[11]) ? 4'b0000 : node5712;
																assign node5712 = (inp[1]) ? 4'b0000 : 4'b0001;
													assign node5716 = (inp[1]) ? node5722 : node5717;
														assign node5717 = (inp[14]) ? node5719 : 4'b1000;
															assign node5719 = (inp[11]) ? 4'b1000 : 4'b1001;
														assign node5722 = (inp[11]) ? 4'b1001 : 4'b1000;
							assign node5726 = (inp[2]) ? node6098 : node5727;
								assign node5727 = (inp[3]) ? node5933 : node5728;
									assign node5728 = (inp[11]) ? node5852 : node5729;
										assign node5729 = (inp[4]) ? node5805 : node5730;
											assign node5730 = (inp[7]) ? node5772 : node5731;
												assign node5731 = (inp[13]) ? node5749 : node5732;
													assign node5732 = (inp[12]) ? node5742 : node5733;
														assign node5733 = (inp[1]) ? node5739 : node5734;
															assign node5734 = (inp[14]) ? node5736 : 4'b0100;
																assign node5736 = (inp[10]) ? 4'b0101 : 4'b1001;
															assign node5739 = (inp[14]) ? 4'b0100 : 4'b0101;
														assign node5742 = (inp[10]) ? node5744 : 4'b1001;
															assign node5744 = (inp[14]) ? node5746 : 4'b0100;
																assign node5746 = (inp[1]) ? 4'b0100 : 4'b1001;
													assign node5749 = (inp[12]) ? node5763 : node5750;
														assign node5750 = (inp[10]) ? node5756 : node5751;
															assign node5751 = (inp[14]) ? 4'b1100 : node5752;
																assign node5752 = (inp[1]) ? 4'b1101 : 4'b1100;
															assign node5756 = (inp[14]) ? node5760 : node5757;
																assign node5757 = (inp[1]) ? 4'b1101 : 4'b1100;
																assign node5760 = (inp[1]) ? 4'b1100 : 4'b1101;
														assign node5763 = (inp[10]) ? node5769 : node5764;
															assign node5764 = (inp[1]) ? 4'b0101 : node5765;
																assign node5765 = (inp[14]) ? 4'b0101 : 4'b0100;
															assign node5769 = (inp[1]) ? 4'b1101 : 4'b0101;
												assign node5772 = (inp[14]) ? node5790 : node5773;
													assign node5773 = (inp[1]) ? node5781 : node5774;
														assign node5774 = (inp[13]) ? 4'b1000 : node5775;
															assign node5775 = (inp[10]) ? 4'b0000 : node5776;
																assign node5776 = (inp[12]) ? 4'b1000 : 4'b0000;
														assign node5781 = (inp[13]) ? node5787 : node5782;
															assign node5782 = (inp[10]) ? 4'b0001 : node5783;
																assign node5783 = (inp[12]) ? 4'b1001 : 4'b0001;
															assign node5787 = (inp[10]) ? 4'b1001 : 4'b0001;
													assign node5790 = (inp[1]) ? node5796 : node5791;
														assign node5791 = (inp[13]) ? node5793 : 4'b1001;
															assign node5793 = (inp[10]) ? 4'b1001 : 4'b0001;
														assign node5796 = (inp[10]) ? 4'b1000 : node5797;
															assign node5797 = (inp[13]) ? node5801 : node5798;
																assign node5798 = (inp[12]) ? 4'b1000 : 4'b0000;
																assign node5801 = (inp[12]) ? 4'b0000 : 4'b1000;
											assign node5805 = (inp[7]) ? node5821 : node5806;
												assign node5806 = (inp[10]) ? node5816 : node5807;
													assign node5807 = (inp[1]) ? 4'b0000 : node5808;
														assign node5808 = (inp[12]) ? node5810 : 4'b0000;
															assign node5810 = (inp[13]) ? 4'b1000 : node5811;
																assign node5811 = (inp[14]) ? 4'b1101 : 4'b1100;
													assign node5816 = (inp[1]) ? 4'b1000 : node5817;
														assign node5817 = (inp[12]) ? 4'b0000 : 4'b1000;
												assign node5821 = (inp[13]) ? node5839 : node5822;
													assign node5822 = (inp[12]) ? node5830 : node5823;
														assign node5823 = (inp[14]) ? node5825 : 4'b0100;
															assign node5825 = (inp[1]) ? 4'b0100 : node5826;
																assign node5826 = (inp[10]) ? 4'b0101 : 4'b1001;
														assign node5830 = (inp[10]) ? node5834 : node5831;
															assign node5831 = (inp[14]) ? 4'b1000 : 4'b1001;
															assign node5834 = (inp[14]) ? node5836 : 4'b0100;
																assign node5836 = (inp[1]) ? 4'b0100 : 4'b1001;
													assign node5839 = (inp[10]) ? node5847 : node5840;
														assign node5840 = (inp[12]) ? node5842 : 4'b0000;
															assign node5842 = (inp[1]) ? 4'b0000 : node5843;
																assign node5843 = (inp[14]) ? 4'b0101 : 4'b0100;
														assign node5847 = (inp[12]) ? node5849 : 4'b1000;
															assign node5849 = (inp[1]) ? 4'b1000 : 4'b0000;
										assign node5852 = (inp[1]) ? node5896 : node5853;
											assign node5853 = (inp[4]) ? node5875 : node5854;
												assign node5854 = (inp[7]) ? node5866 : node5855;
													assign node5855 = (inp[13]) ? node5861 : node5856;
														assign node5856 = (inp[12]) ? node5858 : 4'b0100;
															assign node5858 = (inp[10]) ? 4'b0100 : 4'b1000;
														assign node5861 = (inp[12]) ? node5863 : 4'b1100;
															assign node5863 = (inp[10]) ? 4'b1100 : 4'b0100;
													assign node5866 = (inp[13]) ? node5870 : node5867;
														assign node5867 = (inp[10]) ? 4'b0000 : 4'b1000;
														assign node5870 = (inp[10]) ? 4'b1000 : node5871;
															assign node5871 = (inp[12]) ? 4'b0000 : 4'b1000;
												assign node5875 = (inp[7]) ? node5883 : node5876;
													assign node5876 = (inp[10]) ? node5880 : node5877;
														assign node5877 = (inp[12]) ? 4'b1100 : 4'b0001;
														assign node5880 = (inp[12]) ? 4'b0001 : 4'b1001;
													assign node5883 = (inp[13]) ? node5889 : node5884;
														assign node5884 = (inp[12]) ? node5886 : 4'b0100;
															assign node5886 = (inp[10]) ? 4'b0100 : 4'b1000;
														assign node5889 = (inp[12]) ? node5893 : node5890;
															assign node5890 = (inp[10]) ? 4'b1001 : 4'b0001;
															assign node5893 = (inp[10]) ? 4'b0001 : 4'b0100;
											assign node5896 = (inp[10]) ? node5920 : node5897;
												assign node5897 = (inp[4]) ? node5913 : node5898;
													assign node5898 = (inp[7]) ? node5906 : node5899;
														assign node5899 = (inp[13]) ? node5903 : node5900;
															assign node5900 = (inp[12]) ? 4'b1001 : 4'b0101;
															assign node5903 = (inp[12]) ? 4'b0101 : 4'b1101;
														assign node5906 = (inp[13]) ? node5910 : node5907;
															assign node5907 = (inp[12]) ? 4'b1001 : 4'b0001;
															assign node5910 = (inp[12]) ? 4'b0001 : 4'b1001;
													assign node5913 = (inp[13]) ? 4'b0001 : node5914;
														assign node5914 = (inp[7]) ? node5916 : 4'b0001;
															assign node5916 = (inp[14]) ? 4'b0101 : 4'b1001;
												assign node5920 = (inp[13]) ? node5928 : node5921;
													assign node5921 = (inp[4]) ? node5925 : node5922;
														assign node5922 = (inp[7]) ? 4'b0001 : 4'b0101;
														assign node5925 = (inp[7]) ? 4'b0101 : 4'b1001;
													assign node5928 = (inp[4]) ? 4'b1001 : node5929;
														assign node5929 = (inp[7]) ? 4'b1001 : 4'b1101;
									assign node5933 = (inp[4]) ? node6011 : node5934;
										assign node5934 = (inp[13]) ? node5970 : node5935;
											assign node5935 = (inp[11]) ? node5949 : node5936;
												assign node5936 = (inp[1]) ? node5942 : node5937;
													assign node5937 = (inp[14]) ? node5939 : 4'b1000;
														assign node5939 = (inp[7]) ? 4'b0000 : 4'b1000;
													assign node5942 = (inp[14]) ? node5944 : 4'b0000;
														assign node5944 = (inp[12]) ? node5946 : 4'b0001;
															assign node5946 = (inp[10]) ? 4'b1000 : 4'b0000;
												assign node5949 = (inp[1]) ? node5963 : node5950;
													assign node5950 = (inp[7]) ? node5956 : node5951;
														assign node5951 = (inp[10]) ? node5953 : 4'b0000;
															assign node5953 = (inp[12]) ? 4'b1000 : 4'b0000;
														assign node5956 = (inp[12]) ? node5960 : node5957;
															assign node5957 = (inp[10]) ? 4'b0000 : 4'b0001;
															assign node5960 = (inp[10]) ? 4'b0001 : 4'b1001;
													assign node5963 = (inp[12]) ? 4'b0001 : node5964;
														assign node5964 = (inp[7]) ? 4'b0001 : node5965;
															assign node5965 = (inp[10]) ? 4'b0001 : 4'b1001;
											assign node5970 = (inp[1]) ? node5994 : node5971;
												assign node5971 = (inp[10]) ? node5985 : node5972;
													assign node5972 = (inp[7]) ? node5978 : node5973;
														assign node5973 = (inp[11]) ? 4'b0001 : node5974;
															assign node5974 = (inp[12]) ? 4'b0000 : 4'b0001;
														assign node5978 = (inp[11]) ? 4'b1000 : node5979;
															assign node5979 = (inp[12]) ? node5981 : 4'b1001;
																assign node5981 = (inp[14]) ? 4'b0000 : 4'b0001;
													assign node5985 = (inp[7]) ? 4'b0001 : node5986;
														assign node5986 = (inp[11]) ? 4'b0000 : node5987;
															assign node5987 = (inp[12]) ? 4'b1001 : node5988;
																assign node5988 = (inp[14]) ? 4'b0001 : 4'b0000;
												assign node5994 = (inp[11]) ? 4'b1001 : node5995;
													assign node5995 = (inp[12]) ? node6001 : node5996;
														assign node5996 = (inp[7]) ? 4'b1001 : node5997;
															assign node5997 = (inp[14]) ? 4'b1000 : 4'b1001;
														assign node6001 = (inp[10]) ? node6007 : node6002;
															assign node6002 = (inp[7]) ? node6004 : 4'b0001;
																assign node6004 = (inp[14]) ? 4'b1001 : 4'b1000;
															assign node6007 = (inp[14]) ? 4'b0000 : 4'b0001;
										assign node6011 = (inp[13]) ? node6061 : node6012;
											assign node6012 = (inp[1]) ? node6040 : node6013;
												assign node6013 = (inp[7]) ? node6023 : node6014;
													assign node6014 = (inp[10]) ? node6020 : node6015;
														assign node6015 = (inp[11]) ? node6017 : 4'b0000;
															assign node6017 = (inp[12]) ? 4'b0001 : 4'b1001;
														assign node6020 = (inp[11]) ? 4'b0000 : 4'b0001;
													assign node6023 = (inp[11]) ? node6037 : node6024;
														assign node6024 = (inp[12]) ? node6032 : node6025;
															assign node6025 = (inp[10]) ? node6029 : node6026;
																assign node6026 = (inp[14]) ? 4'b0001 : 4'b0000;
																assign node6029 = (inp[14]) ? 4'b0000 : 4'b0001;
															assign node6032 = (inp[10]) ? 4'b1000 : node6033;
																assign node6033 = (inp[14]) ? 4'b1001 : 4'b0000;
														assign node6037 = (inp[12]) ? 4'b0000 : 4'b1000;
												assign node6040 = (inp[11]) ? node6054 : node6041;
													assign node6041 = (inp[10]) ? node6051 : node6042;
														assign node6042 = (inp[12]) ? node6048 : node6043;
															assign node6043 = (inp[7]) ? 4'b0000 : node6044;
																assign node6044 = (inp[14]) ? 4'b0001 : 4'b0000;
															assign node6048 = (inp[14]) ? 4'b1000 : 4'b1001;
														assign node6051 = (inp[7]) ? 4'b0001 : 4'b0000;
													assign node6054 = (inp[7]) ? 4'b0001 : node6055;
														assign node6055 = (inp[10]) ? 4'b0001 : node6056;
															assign node6056 = (inp[12]) ? 4'b0001 : 4'b1001;
											assign node6061 = (inp[10]) ? node6087 : node6062;
												assign node6062 = (inp[1]) ? node6078 : node6063;
													assign node6063 = (inp[11]) ? 4'b0000 : node6064;
														assign node6064 = (inp[12]) ? node6072 : node6065;
															assign node6065 = (inp[7]) ? node6069 : node6066;
																assign node6066 = (inp[14]) ? 4'b0001 : 4'b0000;
																assign node6069 = (inp[14]) ? 4'b0000 : 4'b0001;
															assign node6072 = (inp[14]) ? node6074 : 4'b0000;
																assign node6074 = (inp[7]) ? 4'b0000 : 4'b0001;
													assign node6078 = (inp[11]) ? 4'b0001 : node6079;
														assign node6079 = (inp[14]) ? node6081 : 4'b0000;
															assign node6081 = (inp[12]) ? 4'b0000 : node6082;
																assign node6082 = (inp[7]) ? 4'b0001 : 4'b0000;
												assign node6087 = (inp[1]) ? 4'b0000 : node6088;
													assign node6088 = (inp[11]) ? 4'b0000 : node6089;
														assign node6089 = (inp[12]) ? 4'b0000 : node6090;
															assign node6090 = (inp[14]) ? 4'b0000 : node6091;
																assign node6091 = (inp[7]) ? 4'b0000 : 4'b0001;
								assign node6098 = (inp[3]) ? node6100 : 4'b1001;
									assign node6100 = (inp[4]) ? node6152 : node6101;
										assign node6101 = (inp[7]) ? 4'b1001 : node6102;
											assign node6102 = (inp[1]) ? node6128 : node6103;
												assign node6103 = (inp[14]) ? node6115 : node6104;
													assign node6104 = (inp[13]) ? node6110 : node6105;
														assign node6105 = (inp[10]) ? 4'b0000 : node6106;
															assign node6106 = (inp[12]) ? 4'b1001 : 4'b0000;
														assign node6110 = (inp[12]) ? node6112 : 4'b1000;
															assign node6112 = (inp[10]) ? 4'b1000 : 4'b0000;
													assign node6115 = (inp[11]) ? node6121 : node6116;
														assign node6116 = (inp[12]) ? node6118 : 4'b1001;
															assign node6118 = (inp[13]) ? 4'b0001 : 4'b1001;
														assign node6121 = (inp[10]) ? node6125 : node6122;
															assign node6122 = (inp[13]) ? 4'b0000 : 4'b1001;
															assign node6125 = (inp[13]) ? 4'b1000 : 4'b0000;
												assign node6128 = (inp[13]) ? node6142 : node6129;
													assign node6129 = (inp[12]) ? node6135 : node6130;
														assign node6130 = (inp[14]) ? node6132 : 4'b0001;
															assign node6132 = (inp[11]) ? 4'b0001 : 4'b0000;
														assign node6135 = (inp[10]) ? node6137 : 4'b1001;
															assign node6137 = (inp[11]) ? 4'b0001 : node6138;
																assign node6138 = (inp[14]) ? 4'b0000 : 4'b0001;
													assign node6142 = (inp[11]) ? node6146 : node6143;
														assign node6143 = (inp[14]) ? 4'b1000 : 4'b1001;
														assign node6146 = (inp[10]) ? 4'b1001 : node6147;
															assign node6147 = (inp[12]) ? 4'b0001 : 4'b1001;
										assign node6152 = (inp[10]) ? node6204 : node6153;
											assign node6153 = (inp[13]) ? node6179 : node6154;
												assign node6154 = (inp[12]) ? node6168 : node6155;
													assign node6155 = (inp[7]) ? node6159 : node6156;
														assign node6156 = (inp[11]) ? 4'b0001 : 4'b0000;
														assign node6159 = (inp[1]) ? node6165 : node6160;
															assign node6160 = (inp[11]) ? 4'b0000 : node6161;
																assign node6161 = (inp[14]) ? 4'b1001 : 4'b0000;
															assign node6165 = (inp[14]) ? 4'b0000 : 4'b0001;
													assign node6168 = (inp[7]) ? 4'b1001 : node6169;
														assign node6169 = (inp[1]) ? node6175 : node6170;
															assign node6170 = (inp[14]) ? node6172 : 4'b1000;
																assign node6172 = (inp[11]) ? 4'b1000 : 4'b1001;
															assign node6175 = (inp[11]) ? 4'b0001 : 4'b0000;
												assign node6179 = (inp[11]) ? node6195 : node6180;
													assign node6180 = (inp[1]) ? node6190 : node6181;
														assign node6181 = (inp[14]) ? node6183 : 4'b0001;
															assign node6183 = (inp[7]) ? node6187 : node6184;
																assign node6184 = (inp[12]) ? 4'b0000 : 4'b0001;
																assign node6187 = (inp[12]) ? 4'b0001 : 4'b0000;
														assign node6190 = (inp[14]) ? 4'b0000 : node6191;
															assign node6191 = (inp[12]) ? 4'b0001 : 4'b0000;
													assign node6195 = (inp[1]) ? 4'b0001 : node6196;
														assign node6196 = (inp[12]) ? node6200 : node6197;
															assign node6197 = (inp[7]) ? 4'b0001 : 4'b0000;
															assign node6200 = (inp[7]) ? 4'b0000 : 4'b0001;
											assign node6204 = (inp[13]) ? node6232 : node6205;
												assign node6205 = (inp[1]) ? node6221 : node6206;
													assign node6206 = (inp[14]) ? node6214 : node6207;
														assign node6207 = (inp[7]) ? 4'b0000 : node6208;
															assign node6208 = (inp[11]) ? node6210 : 4'b0000;
																assign node6210 = (inp[12]) ? 4'b0001 : 4'b0000;
														assign node6214 = (inp[11]) ? 4'b0000 : node6215;
															assign node6215 = (inp[7]) ? node6217 : 4'b0000;
																assign node6217 = (inp[12]) ? 4'b1001 : 4'b0001;
													assign node6221 = (inp[11]) ? 4'b0001 : node6222;
														assign node6222 = (inp[7]) ? 4'b0001 : node6223;
															assign node6223 = (inp[12]) ? node6227 : node6224;
																assign node6224 = (inp[14]) ? 4'b0001 : 4'b0000;
																assign node6227 = (inp[14]) ? 4'b1000 : 4'b0000;
												assign node6232 = (inp[11]) ? 4'b0000 : node6233;
													assign node6233 = (inp[1]) ? 4'b0000 : node6234;
														assign node6234 = (inp[12]) ? node6236 : 4'b0000;
															assign node6236 = (inp[14]) ? node6240 : node6237;
																assign node6237 = (inp[7]) ? 4'b0001 : 4'b0000;
																assign node6240 = (inp[7]) ? 4'b0000 : 4'b0001;
			assign node6245 = (inp[15]) ? node9567 : node6246;
				assign node6246 = (inp[6]) ? node7082 : node6247;
					assign node6247 = (inp[0]) ? 4'b0101 : node6248;
						assign node6248 = (inp[2]) ? node6772 : node6249;
							assign node6249 = (inp[1]) ? node6521 : node6250;
								assign node6250 = (inp[14]) ? node6348 : node6251;
									assign node6251 = (inp[3]) ? node6311 : node6252;
										assign node6252 = (inp[5]) ? node6280 : node6253;
											assign node6253 = (inp[7]) ? node6273 : node6254;
												assign node6254 = (inp[4]) ? node6262 : node6255;
													assign node6255 = (inp[13]) ? node6257 : 4'b0111;
														assign node6257 = (inp[12]) ? node6259 : 4'b0000;
															assign node6259 = (inp[10]) ? 4'b0000 : 4'b0111;
													assign node6262 = (inp[13]) ? node6268 : node6263;
														assign node6263 = (inp[12]) ? node6265 : 4'b1000;
															assign node6265 = (inp[10]) ? 4'b1000 : 4'b0000;
														assign node6268 = (inp[12]) ? node6270 : 4'b0000;
															assign node6270 = (inp[10]) ? 4'b0000 : 4'b1000;
												assign node6273 = (inp[12]) ? 4'b0111 : node6274;
													assign node6274 = (inp[13]) ? node6276 : 4'b0111;
														assign node6276 = (inp[4]) ? 4'b0000 : 4'b0111;
											assign node6280 = (inp[13]) ? node6298 : node6281;
												assign node6281 = (inp[10]) ? node6293 : node6282;
													assign node6282 = (inp[12]) ? node6288 : node6283;
														assign node6283 = (inp[4]) ? node6285 : 4'b1100;
															assign node6285 = (inp[7]) ? 4'b1100 : 4'b1000;
														assign node6288 = (inp[4]) ? node6290 : 4'b0100;
															assign node6290 = (inp[7]) ? 4'b0100 : 4'b0000;
													assign node6293 = (inp[7]) ? 4'b1100 : node6294;
														assign node6294 = (inp[4]) ? 4'b1000 : 4'b1100;
												assign node6298 = (inp[12]) ? node6304 : node6299;
													assign node6299 = (inp[7]) ? node6301 : 4'b0000;
														assign node6301 = (inp[4]) ? 4'b0000 : 4'b0100;
													assign node6304 = (inp[10]) ? 4'b0000 : node6305;
														assign node6305 = (inp[7]) ? 4'b1100 : node6306;
															assign node6306 = (inp[4]) ? 4'b1000 : 4'b1100;
										assign node6311 = (inp[13]) ? node6329 : node6312;
											assign node6312 = (inp[4]) ? node6318 : node6313;
												assign node6313 = (inp[10]) ? 4'b1000 : node6314;
													assign node6314 = (inp[12]) ? 4'b0000 : 4'b1000;
												assign node6318 = (inp[7]) ? node6324 : node6319;
													assign node6319 = (inp[12]) ? node6321 : 4'b1100;
														assign node6321 = (inp[10]) ? 4'b1100 : 4'b0100;
													assign node6324 = (inp[12]) ? node6326 : 4'b1000;
														assign node6326 = (inp[10]) ? 4'b1000 : 4'b0000;
											assign node6329 = (inp[7]) ? node6337 : node6330;
												assign node6330 = (inp[10]) ? 4'b0100 : node6331;
													assign node6331 = (inp[12]) ? node6333 : 4'b0100;
														assign node6333 = (inp[4]) ? 4'b1100 : 4'b1000;
												assign node6337 = (inp[4]) ? node6343 : node6338;
													assign node6338 = (inp[12]) ? node6340 : 4'b0000;
														assign node6340 = (inp[10]) ? 4'b0000 : 4'b1000;
													assign node6343 = (inp[12]) ? node6345 : 4'b0100;
														assign node6345 = (inp[10]) ? 4'b0100 : 4'b1000;
									assign node6348 = (inp[11]) ? node6444 : node6349;
										assign node6349 = (inp[3]) ? node6407 : node6350;
											assign node6350 = (inp[5]) ? node6372 : node6351;
												assign node6351 = (inp[7]) ? node6365 : node6352;
													assign node6352 = (inp[4]) ? node6358 : node6353;
														assign node6353 = (inp[12]) ? 4'b0111 : node6354;
															assign node6354 = (inp[10]) ? 4'b0001 : 4'b0111;
														assign node6358 = (inp[13]) ? node6360 : 4'b0001;
															assign node6360 = (inp[10]) ? node6362 : 4'b1001;
																assign node6362 = (inp[12]) ? 4'b1001 : 4'b0001;
													assign node6365 = (inp[10]) ? node6367 : 4'b0111;
														assign node6367 = (inp[4]) ? node6369 : 4'b0111;
															assign node6369 = (inp[13]) ? 4'b0001 : 4'b0111;
												assign node6372 = (inp[4]) ? node6386 : node6373;
													assign node6373 = (inp[13]) ? node6379 : node6374;
														assign node6374 = (inp[12]) ? 4'b0101 : node6375;
															assign node6375 = (inp[10]) ? 4'b1101 : 4'b0101;
														assign node6379 = (inp[10]) ? node6381 : 4'b1101;
															assign node6381 = (inp[12]) ? 4'b1101 : node6382;
																assign node6382 = (inp[7]) ? 4'b0101 : 4'b0001;
													assign node6386 = (inp[7]) ? node6398 : node6387;
														assign node6387 = (inp[13]) ? node6393 : node6388;
															assign node6388 = (inp[10]) ? node6390 : 4'b0001;
																assign node6390 = (inp[12]) ? 4'b0001 : 4'b1001;
															assign node6393 = (inp[10]) ? node6395 : 4'b1001;
																assign node6395 = (inp[12]) ? 4'b1001 : 4'b0001;
														assign node6398 = (inp[13]) ? node6404 : node6399;
															assign node6399 = (inp[12]) ? 4'b0101 : node6400;
																assign node6400 = (inp[10]) ? 4'b1101 : 4'b0101;
															assign node6404 = (inp[10]) ? 4'b0001 : 4'b1101;
											assign node6407 = (inp[13]) ? node6425 : node6408;
												assign node6408 = (inp[10]) ? node6414 : node6409;
													assign node6409 = (inp[7]) ? 4'b0001 : node6410;
														assign node6410 = (inp[4]) ? 4'b0101 : 4'b0001;
													assign node6414 = (inp[12]) ? node6420 : node6415;
														assign node6415 = (inp[4]) ? node6417 : 4'b1001;
															assign node6417 = (inp[7]) ? 4'b1001 : 4'b1101;
														assign node6420 = (inp[7]) ? 4'b0001 : node6421;
															assign node6421 = (inp[4]) ? 4'b0101 : 4'b0001;
												assign node6425 = (inp[4]) ? node6433 : node6426;
													assign node6426 = (inp[12]) ? 4'b1001 : node6427;
														assign node6427 = (inp[10]) ? node6429 : 4'b1001;
															assign node6429 = (inp[7]) ? 4'b0001 : 4'b0101;
													assign node6433 = (inp[7]) ? node6439 : node6434;
														assign node6434 = (inp[10]) ? node6436 : 4'b1101;
															assign node6436 = (inp[12]) ? 4'b1101 : 4'b0101;
														assign node6439 = (inp[12]) ? 4'b1001 : node6440;
															assign node6440 = (inp[10]) ? 4'b0101 : 4'b1001;
										assign node6444 = (inp[3]) ? node6490 : node6445;
											assign node6445 = (inp[5]) ? node6471 : node6446;
												assign node6446 = (inp[7]) ? node6464 : node6447;
													assign node6447 = (inp[4]) ? node6455 : node6448;
														assign node6448 = (inp[13]) ? node6450 : 4'b0111;
															assign node6450 = (inp[12]) ? node6452 : 4'b0000;
																assign node6452 = (inp[10]) ? 4'b0000 : 4'b0111;
														assign node6455 = (inp[13]) ? node6459 : node6456;
															assign node6456 = (inp[12]) ? 4'b0000 : 4'b1000;
															assign node6459 = (inp[10]) ? 4'b0000 : node6460;
																assign node6460 = (inp[12]) ? 4'b1000 : 4'b0000;
													assign node6464 = (inp[12]) ? 4'b0111 : node6465;
														assign node6465 = (inp[4]) ? node6467 : 4'b0111;
															assign node6467 = (inp[13]) ? 4'b0000 : 4'b0111;
												assign node6471 = (inp[13]) ? node6479 : node6472;
													assign node6472 = (inp[12]) ? node6474 : 4'b1100;
														assign node6474 = (inp[10]) ? 4'b1100 : node6475;
															assign node6475 = (inp[4]) ? 4'b0000 : 4'b0100;
													assign node6479 = (inp[12]) ? node6483 : node6480;
														assign node6480 = (inp[4]) ? 4'b0000 : 4'b0100;
														assign node6483 = (inp[10]) ? 4'b0000 : node6484;
															assign node6484 = (inp[7]) ? 4'b1100 : node6485;
																assign node6485 = (inp[4]) ? 4'b1000 : 4'b1100;
											assign node6490 = (inp[13]) ? node6506 : node6491;
												assign node6491 = (inp[10]) ? node6501 : node6492;
													assign node6492 = (inp[12]) ? node6496 : node6493;
														assign node6493 = (inp[7]) ? 4'b1000 : 4'b1100;
														assign node6496 = (inp[7]) ? 4'b0000 : node6497;
															assign node6497 = (inp[4]) ? 4'b0100 : 4'b0000;
													assign node6501 = (inp[4]) ? node6503 : 4'b1000;
														assign node6503 = (inp[7]) ? 4'b1000 : 4'b1100;
												assign node6506 = (inp[7]) ? node6514 : node6507;
													assign node6507 = (inp[5]) ? 4'b0100 : node6508;
														assign node6508 = (inp[4]) ? node6510 : 4'b0100;
															assign node6510 = (inp[10]) ? 4'b0100 : 4'b1100;
													assign node6514 = (inp[4]) ? node6516 : 4'b0000;
														assign node6516 = (inp[10]) ? 4'b0100 : node6517;
															assign node6517 = (inp[12]) ? 4'b1000 : 4'b0100;
								assign node6521 = (inp[11]) ? node6687 : node6522;
									assign node6522 = (inp[14]) ? node6596 : node6523;
										assign node6523 = (inp[13]) ? node6563 : node6524;
											assign node6524 = (inp[3]) ? node6546 : node6525;
												assign node6525 = (inp[5]) ? node6531 : node6526;
													assign node6526 = (inp[4]) ? node6528 : 4'b0111;
														assign node6528 = (inp[7]) ? 4'b0111 : 4'b1001;
													assign node6531 = (inp[10]) ? node6541 : node6532;
														assign node6532 = (inp[12]) ? node6536 : node6533;
															assign node6533 = (inp[7]) ? 4'b1101 : 4'b1001;
															assign node6536 = (inp[7]) ? 4'b0101 : node6537;
																assign node6537 = (inp[4]) ? 4'b0001 : 4'b0101;
														assign node6541 = (inp[4]) ? node6543 : 4'b1101;
															assign node6543 = (inp[7]) ? 4'b1101 : 4'b1001;
												assign node6546 = (inp[7]) ? node6558 : node6547;
													assign node6547 = (inp[4]) ? node6553 : node6548;
														assign node6548 = (inp[12]) ? node6550 : 4'b1001;
															assign node6550 = (inp[10]) ? 4'b1001 : 4'b0001;
														assign node6553 = (inp[12]) ? node6555 : 4'b1101;
															assign node6555 = (inp[10]) ? 4'b1101 : 4'b0101;
													assign node6558 = (inp[10]) ? 4'b1001 : node6559;
														assign node6559 = (inp[12]) ? 4'b0001 : 4'b1001;
											assign node6563 = (inp[10]) ? node6585 : node6564;
												assign node6564 = (inp[12]) ? node6572 : node6565;
													assign node6565 = (inp[3]) ? node6567 : 4'b0001;
														assign node6567 = (inp[4]) ? 4'b0101 : node6568;
															assign node6568 = (inp[7]) ? 4'b0001 : 4'b0101;
													assign node6572 = (inp[3]) ? node6580 : node6573;
														assign node6573 = (inp[5]) ? node6575 : 4'b0111;
															assign node6575 = (inp[4]) ? node6577 : 4'b1101;
																assign node6577 = (inp[7]) ? 4'b1101 : 4'b1001;
														assign node6580 = (inp[4]) ? node6582 : 4'b1001;
															assign node6582 = (inp[7]) ? 4'b1001 : 4'b1101;
												assign node6585 = (inp[3]) ? node6591 : node6586;
													assign node6586 = (inp[4]) ? 4'b0001 : node6587;
														assign node6587 = (inp[7]) ? 4'b0101 : 4'b0001;
													assign node6591 = (inp[7]) ? node6593 : 4'b0101;
														assign node6593 = (inp[4]) ? 4'b0101 : 4'b0001;
										assign node6596 = (inp[13]) ? node6638 : node6597;
											assign node6597 = (inp[3]) ? node6623 : node6598;
												assign node6598 = (inp[5]) ? node6608 : node6599;
													assign node6599 = (inp[4]) ? node6601 : 4'b0111;
														assign node6601 = (inp[7]) ? 4'b0111 : node6602;
															assign node6602 = (inp[10]) ? 4'b1000 : node6603;
																assign node6603 = (inp[12]) ? 4'b0000 : 4'b1000;
													assign node6608 = (inp[7]) ? node6618 : node6609;
														assign node6609 = (inp[4]) ? node6613 : node6610;
															assign node6610 = (inp[12]) ? 4'b0100 : 4'b1100;
															assign node6613 = (inp[12]) ? node6615 : 4'b1000;
																assign node6615 = (inp[10]) ? 4'b1000 : 4'b0000;
														assign node6618 = (inp[12]) ? node6620 : 4'b1100;
															assign node6620 = (inp[10]) ? 4'b1100 : 4'b0100;
												assign node6623 = (inp[7]) ? node6633 : node6624;
													assign node6624 = (inp[4]) ? node6628 : node6625;
														assign node6625 = (inp[10]) ? 4'b1000 : 4'b0000;
														assign node6628 = (inp[10]) ? 4'b1100 : node6629;
															assign node6629 = (inp[12]) ? 4'b0100 : 4'b1100;
													assign node6633 = (inp[12]) ? node6635 : 4'b1000;
														assign node6635 = (inp[10]) ? 4'b1000 : 4'b0000;
											assign node6638 = (inp[3]) ? node6670 : node6639;
												assign node6639 = (inp[5]) ? node6657 : node6640;
													assign node6640 = (inp[4]) ? node6646 : node6641;
														assign node6641 = (inp[7]) ? 4'b0111 : node6642;
															assign node6642 = (inp[12]) ? 4'b0111 : 4'b0000;
														assign node6646 = (inp[7]) ? node6652 : node6647;
															assign node6647 = (inp[10]) ? 4'b0000 : node6648;
																assign node6648 = (inp[12]) ? 4'b1000 : 4'b0000;
															assign node6652 = (inp[12]) ? node6654 : 4'b0000;
																assign node6654 = (inp[10]) ? 4'b0000 : 4'b0111;
													assign node6657 = (inp[12]) ? node6659 : 4'b0000;
														assign node6659 = (inp[10]) ? node6665 : node6660;
															assign node6660 = (inp[4]) ? node6662 : 4'b1100;
																assign node6662 = (inp[7]) ? 4'b1100 : 4'b1000;
															assign node6665 = (inp[4]) ? 4'b0000 : node6666;
																assign node6666 = (inp[7]) ? 4'b0100 : 4'b0000;
												assign node6670 = (inp[12]) ? node6676 : node6671;
													assign node6671 = (inp[4]) ? 4'b0100 : node6672;
														assign node6672 = (inp[7]) ? 4'b0000 : 4'b0100;
													assign node6676 = (inp[10]) ? node6682 : node6677;
														assign node6677 = (inp[7]) ? 4'b1000 : node6678;
															assign node6678 = (inp[4]) ? 4'b1100 : 4'b1000;
														assign node6682 = (inp[4]) ? 4'b0100 : node6683;
															assign node6683 = (inp[7]) ? 4'b0000 : 4'b0100;
									assign node6687 = (inp[13]) ? node6729 : node6688;
										assign node6688 = (inp[3]) ? node6716 : node6689;
											assign node6689 = (inp[5]) ? node6697 : node6690;
												assign node6690 = (inp[7]) ? 4'b0111 : node6691;
													assign node6691 = (inp[4]) ? node6693 : 4'b0111;
														assign node6693 = (inp[10]) ? 4'b1001 : 4'b0001;
												assign node6697 = (inp[7]) ? node6711 : node6698;
													assign node6698 = (inp[4]) ? node6704 : node6699;
														assign node6699 = (inp[12]) ? node6701 : 4'b1101;
															assign node6701 = (inp[10]) ? 4'b1101 : 4'b0101;
														assign node6704 = (inp[14]) ? 4'b1001 : node6705;
															assign node6705 = (inp[12]) ? node6707 : 4'b1001;
																assign node6707 = (inp[10]) ? 4'b1001 : 4'b0001;
													assign node6711 = (inp[10]) ? 4'b1101 : node6712;
														assign node6712 = (inp[12]) ? 4'b0101 : 4'b1101;
											assign node6716 = (inp[10]) ? node6724 : node6717;
												assign node6717 = (inp[12]) ? 4'b0001 : node6718;
													assign node6718 = (inp[4]) ? node6720 : 4'b1001;
														assign node6720 = (inp[7]) ? 4'b1001 : 4'b1101;
												assign node6724 = (inp[7]) ? 4'b1001 : node6725;
													assign node6725 = (inp[4]) ? 4'b1101 : 4'b1001;
										assign node6729 = (inp[10]) ? node6759 : node6730;
											assign node6730 = (inp[12]) ? node6744 : node6731;
												assign node6731 = (inp[3]) ? node6739 : node6732;
													assign node6732 = (inp[4]) ? 4'b0001 : node6733;
														assign node6733 = (inp[7]) ? node6735 : 4'b0001;
															assign node6735 = (inp[5]) ? 4'b0101 : 4'b0111;
													assign node6739 = (inp[4]) ? 4'b0101 : node6740;
														assign node6740 = (inp[7]) ? 4'b0001 : 4'b0101;
												assign node6744 = (inp[3]) ? node6754 : node6745;
													assign node6745 = (inp[5]) ? node6751 : node6746;
														assign node6746 = (inp[4]) ? node6748 : 4'b0111;
															assign node6748 = (inp[7]) ? 4'b0111 : 4'b1001;
														assign node6751 = (inp[7]) ? 4'b1101 : 4'b1001;
													assign node6754 = (inp[7]) ? 4'b1001 : node6755;
														assign node6755 = (inp[4]) ? 4'b1101 : 4'b1001;
											assign node6759 = (inp[3]) ? node6767 : node6760;
												assign node6760 = (inp[4]) ? 4'b0001 : node6761;
													assign node6761 = (inp[7]) ? node6763 : 4'b0001;
														assign node6763 = (inp[5]) ? 4'b0101 : 4'b0111;
												assign node6767 = (inp[4]) ? 4'b0101 : node6768;
													assign node6768 = (inp[7]) ? 4'b0001 : 4'b0101;
							assign node6772 = (inp[5]) ? node6774 : 4'b0111;
								assign node6774 = (inp[3]) ? node6880 : node6775;
									assign node6775 = (inp[4]) ? node6801 : node6776;
										assign node6776 = (inp[13]) ? node6778 : 4'b0111;
											assign node6778 = (inp[7]) ? 4'b0111 : node6779;
												assign node6779 = (inp[12]) ? node6791 : node6780;
													assign node6780 = (inp[1]) ? node6786 : node6781;
														assign node6781 = (inp[14]) ? node6783 : 4'b0000;
															assign node6783 = (inp[11]) ? 4'b0000 : 4'b0111;
														assign node6786 = (inp[14]) ? node6788 : 4'b0001;
															assign node6788 = (inp[11]) ? 4'b0001 : 4'b0000;
													assign node6791 = (inp[10]) ? node6793 : 4'b0111;
														assign node6793 = (inp[14]) ? node6797 : node6794;
															assign node6794 = (inp[1]) ? 4'b0001 : 4'b0000;
															assign node6797 = (inp[1]) ? 4'b0001 : 4'b0111;
										assign node6801 = (inp[7]) ? node6861 : node6802;
											assign node6802 = (inp[1]) ? node6828 : node6803;
												assign node6803 = (inp[13]) ? node6819 : node6804;
													assign node6804 = (inp[11]) ? node6814 : node6805;
														assign node6805 = (inp[14]) ? node6809 : node6806;
															assign node6806 = (inp[10]) ? 4'b1000 : 4'b0000;
															assign node6809 = (inp[10]) ? node6811 : 4'b0001;
																assign node6811 = (inp[12]) ? 4'b0001 : 4'b1001;
														assign node6814 = (inp[12]) ? node6816 : 4'b1000;
															assign node6816 = (inp[10]) ? 4'b1000 : 4'b0000;
													assign node6819 = (inp[11]) ? 4'b0000 : node6820;
														assign node6820 = (inp[14]) ? 4'b0001 : node6821;
															assign node6821 = (inp[10]) ? 4'b0000 : node6822;
																assign node6822 = (inp[12]) ? 4'b1000 : 4'b0000;
												assign node6828 = (inp[14]) ? node6840 : node6829;
													assign node6829 = (inp[13]) ? node6835 : node6830;
														assign node6830 = (inp[12]) ? node6832 : 4'b1001;
															assign node6832 = (inp[10]) ? 4'b1001 : 4'b0001;
														assign node6835 = (inp[12]) ? node6837 : 4'b0001;
															assign node6837 = (inp[10]) ? 4'b0001 : 4'b1001;
													assign node6840 = (inp[11]) ? node6852 : node6841;
														assign node6841 = (inp[13]) ? node6847 : node6842;
															assign node6842 = (inp[12]) ? node6844 : 4'b1000;
																assign node6844 = (inp[10]) ? 4'b1000 : 4'b0000;
															assign node6847 = (inp[12]) ? node6849 : 4'b0000;
																assign node6849 = (inp[10]) ? 4'b0000 : 4'b1000;
														assign node6852 = (inp[10]) ? 4'b1001 : node6853;
															assign node6853 = (inp[13]) ? node6857 : node6854;
																assign node6854 = (inp[12]) ? 4'b0001 : 4'b1001;
																assign node6857 = (inp[12]) ? 4'b1001 : 4'b0001;
											assign node6861 = (inp[13]) ? node6863 : 4'b0111;
												assign node6863 = (inp[10]) ? node6869 : node6864;
													assign node6864 = (inp[12]) ? 4'b0111 : node6865;
														assign node6865 = (inp[1]) ? 4'b0001 : 4'b0000;
													assign node6869 = (inp[1]) ? node6875 : node6870;
														assign node6870 = (inp[14]) ? node6872 : 4'b0000;
															assign node6872 = (inp[11]) ? 4'b0000 : 4'b0111;
														assign node6875 = (inp[14]) ? node6877 : 4'b0001;
															assign node6877 = (inp[11]) ? 4'b0001 : 4'b0000;
									assign node6880 = (inp[4]) ? node6962 : node6881;
										assign node6881 = (inp[1]) ? node6917 : node6882;
											assign node6882 = (inp[14]) ? node6896 : node6883;
												assign node6883 = (inp[13]) ? node6889 : node6884;
													assign node6884 = (inp[10]) ? 4'b1000 : node6885;
														assign node6885 = (inp[12]) ? 4'b0000 : 4'b1000;
													assign node6889 = (inp[12]) ? node6893 : node6890;
														assign node6890 = (inp[7]) ? 4'b0000 : 4'b0100;
														assign node6893 = (inp[10]) ? 4'b0000 : 4'b1000;
												assign node6896 = (inp[11]) ? node6908 : node6897;
													assign node6897 = (inp[13]) ? node6903 : node6898;
														assign node6898 = (inp[7]) ? 4'b0001 : node6899;
															assign node6899 = (inp[12]) ? 4'b0001 : 4'b1001;
														assign node6903 = (inp[12]) ? 4'b1001 : node6904;
															assign node6904 = (inp[10]) ? 4'b0001 : 4'b1001;
													assign node6908 = (inp[12]) ? node6912 : node6909;
														assign node6909 = (inp[13]) ? 4'b0000 : 4'b1000;
														assign node6912 = (inp[13]) ? 4'b1000 : node6913;
															assign node6913 = (inp[10]) ? 4'b1000 : 4'b0000;
											assign node6917 = (inp[13]) ? node6935 : node6918;
												assign node6918 = (inp[12]) ? node6924 : node6919;
													assign node6919 = (inp[11]) ? 4'b1001 : node6920;
														assign node6920 = (inp[14]) ? 4'b1000 : 4'b1001;
													assign node6924 = (inp[10]) ? node6930 : node6925;
														assign node6925 = (inp[14]) ? node6927 : 4'b0001;
															assign node6927 = (inp[11]) ? 4'b0001 : 4'b0000;
														assign node6930 = (inp[11]) ? 4'b1001 : node6931;
															assign node6931 = (inp[14]) ? 4'b1000 : 4'b1001;
												assign node6935 = (inp[7]) ? node6947 : node6936;
													assign node6936 = (inp[12]) ? node6942 : node6937;
														assign node6937 = (inp[11]) ? 4'b0101 : node6938;
															assign node6938 = (inp[14]) ? 4'b0100 : 4'b0101;
														assign node6942 = (inp[10]) ? 4'b0101 : node6943;
															assign node6943 = (inp[11]) ? 4'b1001 : 4'b1000;
													assign node6947 = (inp[12]) ? node6953 : node6948;
														assign node6948 = (inp[11]) ? 4'b0001 : node6949;
															assign node6949 = (inp[14]) ? 4'b0000 : 4'b0001;
														assign node6953 = (inp[10]) ? node6959 : node6954;
															assign node6954 = (inp[11]) ? 4'b1001 : node6955;
																assign node6955 = (inp[14]) ? 4'b1000 : 4'b1001;
															assign node6959 = (inp[14]) ? 4'b0000 : 4'b0001;
										assign node6962 = (inp[7]) ? node7020 : node6963;
											assign node6963 = (inp[1]) ? node6995 : node6964;
												assign node6964 = (inp[11]) ? node6984 : node6965;
													assign node6965 = (inp[14]) ? node6973 : node6966;
														assign node6966 = (inp[10]) ? 4'b1100 : node6967;
															assign node6967 = (inp[13]) ? node6969 : 4'b0100;
																assign node6969 = (inp[12]) ? 4'b1100 : 4'b0100;
														assign node6973 = (inp[13]) ? node6979 : node6974;
															assign node6974 = (inp[10]) ? node6976 : 4'b0101;
																assign node6976 = (inp[12]) ? 4'b0101 : 4'b1101;
															assign node6979 = (inp[12]) ? 4'b1101 : node6980;
																assign node6980 = (inp[10]) ? 4'b0101 : 4'b1101;
													assign node6984 = (inp[13]) ? node6990 : node6985;
														assign node6985 = (inp[12]) ? node6987 : 4'b1100;
															assign node6987 = (inp[10]) ? 4'b1100 : 4'b0100;
														assign node6990 = (inp[10]) ? 4'b0100 : node6991;
															assign node6991 = (inp[12]) ? 4'b1100 : 4'b0100;
												assign node6995 = (inp[13]) ? node7007 : node6996;
													assign node6996 = (inp[11]) ? 4'b1101 : node6997;
														assign node6997 = (inp[14]) ? node7001 : node6998;
															assign node6998 = (inp[12]) ? 4'b0101 : 4'b1101;
															assign node7001 = (inp[12]) ? node7003 : 4'b1100;
																assign node7003 = (inp[10]) ? 4'b1100 : 4'b0100;
													assign node7007 = (inp[11]) ? node7015 : node7008;
														assign node7008 = (inp[14]) ? node7010 : 4'b0101;
															assign node7010 = (inp[12]) ? node7012 : 4'b0100;
																assign node7012 = (inp[10]) ? 4'b0100 : 4'b1100;
														assign node7015 = (inp[10]) ? 4'b0101 : node7016;
															assign node7016 = (inp[12]) ? 4'b1101 : 4'b0101;
											assign node7020 = (inp[13]) ? node7050 : node7021;
												assign node7021 = (inp[1]) ? node7035 : node7022;
													assign node7022 = (inp[10]) ? 4'b1000 : node7023;
														assign node7023 = (inp[12]) ? node7029 : node7024;
															assign node7024 = (inp[11]) ? 4'b1000 : node7025;
																assign node7025 = (inp[14]) ? 4'b0001 : 4'b1000;
															assign node7029 = (inp[11]) ? 4'b0000 : node7030;
																assign node7030 = (inp[14]) ? 4'b0001 : 4'b0000;
													assign node7035 = (inp[12]) ? node7041 : node7036;
														assign node7036 = (inp[14]) ? node7038 : 4'b1001;
															assign node7038 = (inp[11]) ? 4'b1001 : 4'b1000;
														assign node7041 = (inp[10]) ? node7047 : node7042;
															assign node7042 = (inp[11]) ? 4'b0001 : node7043;
																assign node7043 = (inp[14]) ? 4'b0000 : 4'b0001;
															assign node7047 = (inp[11]) ? 4'b1001 : 4'b1000;
												assign node7050 = (inp[12]) ? node7064 : node7051;
													assign node7051 = (inp[1]) ? node7059 : node7052;
														assign node7052 = (inp[14]) ? node7054 : 4'b0100;
															assign node7054 = (inp[11]) ? 4'b0100 : node7055;
																assign node7055 = (inp[10]) ? 4'b0101 : 4'b1001;
														assign node7059 = (inp[14]) ? node7061 : 4'b0101;
															assign node7061 = (inp[11]) ? 4'b0101 : 4'b0100;
													assign node7064 = (inp[10]) ? node7072 : node7065;
														assign node7065 = (inp[1]) ? node7069 : node7066;
															assign node7066 = (inp[11]) ? 4'b1000 : 4'b1001;
															assign node7069 = (inp[11]) ? 4'b1001 : 4'b1000;
														assign node7072 = (inp[1]) ? node7076 : node7073;
															assign node7073 = (inp[11]) ? 4'b0100 : 4'b1001;
															assign node7076 = (inp[14]) ? node7078 : 4'b0101;
																assign node7078 = (inp[11]) ? 4'b0101 : 4'b0100;
					assign node7082 = (inp[5]) ? node8116 : node7083;
						assign node7083 = (inp[0]) ? node7845 : node7084;
							assign node7084 = (inp[11]) ? node7538 : node7085;
								assign node7085 = (inp[3]) ? node7333 : node7086;
									assign node7086 = (inp[2]) ? node7182 : node7087;
										assign node7087 = (inp[10]) ? node7139 : node7088;
											assign node7088 = (inp[4]) ? node7122 : node7089;
												assign node7089 = (inp[13]) ? node7103 : node7090;
													assign node7090 = (inp[12]) ? node7098 : node7091;
														assign node7091 = (inp[14]) ? node7095 : node7092;
															assign node7092 = (inp[1]) ? 4'b1101 : 4'b1100;
															assign node7095 = (inp[1]) ? 4'b1100 : 4'b0101;
														assign node7098 = (inp[14]) ? node7100 : 4'b0101;
															assign node7100 = (inp[1]) ? 4'b0100 : 4'b0101;
													assign node7103 = (inp[7]) ? node7109 : node7104;
														assign node7104 = (inp[1]) ? 4'b1000 : node7105;
															assign node7105 = (inp[12]) ? 4'b0000 : 4'b1000;
														assign node7109 = (inp[12]) ? node7115 : node7110;
															assign node7110 = (inp[1]) ? node7112 : 4'b1101;
																assign node7112 = (inp[14]) ? 4'b0100 : 4'b0101;
															assign node7115 = (inp[1]) ? node7119 : node7116;
																assign node7116 = (inp[14]) ? 4'b1101 : 4'b1100;
																assign node7119 = (inp[14]) ? 4'b1100 : 4'b1101;
												assign node7122 = (inp[7]) ? node7134 : node7123;
													assign node7123 = (inp[13]) ? node7129 : node7124;
														assign node7124 = (inp[12]) ? node7126 : 4'b1000;
															assign node7126 = (inp[1]) ? 4'b1000 : 4'b0000;
														assign node7129 = (inp[1]) ? 4'b1100 : node7130;
															assign node7130 = (inp[12]) ? 4'b0100 : 4'b1100;
													assign node7134 = (inp[1]) ? 4'b1000 : node7135;
														assign node7135 = (inp[12]) ? 4'b0000 : 4'b1000;
											assign node7139 = (inp[12]) ? node7155 : node7140;
												assign node7140 = (inp[4]) ? node7150 : node7141;
													assign node7141 = (inp[7]) ? node7143 : 4'b0000;
														assign node7143 = (inp[13]) ? 4'b0000 : node7144;
															assign node7144 = (inp[1]) ? node7146 : 4'b1100;
																assign node7146 = (inp[14]) ? 4'b1100 : 4'b1101;
													assign node7150 = (inp[13]) ? 4'b0100 : node7151;
														assign node7151 = (inp[7]) ? 4'b0000 : 4'b0100;
												assign node7155 = (inp[1]) ? node7171 : node7156;
													assign node7156 = (inp[4]) ? node7166 : node7157;
														assign node7157 = (inp[14]) ? node7161 : node7158;
															assign node7158 = (inp[13]) ? 4'b0100 : 4'b1100;
															assign node7161 = (inp[13]) ? node7163 : 4'b0101;
																assign node7163 = (inp[7]) ? 4'b1101 : 4'b1000;
														assign node7166 = (inp[7]) ? 4'b1000 : node7167;
															assign node7167 = (inp[13]) ? 4'b1100 : 4'b1000;
													assign node7171 = (inp[4]) ? node7177 : node7172;
														assign node7172 = (inp[7]) ? node7174 : 4'b0000;
															assign node7174 = (inp[14]) ? 4'b0000 : 4'b1101;
														assign node7177 = (inp[7]) ? node7179 : 4'b0100;
															assign node7179 = (inp[13]) ? 4'b0100 : 4'b0000;
										assign node7182 = (inp[7]) ? node7252 : node7183;
											assign node7183 = (inp[4]) ? node7221 : node7184;
												assign node7184 = (inp[13]) ? node7200 : node7185;
													assign node7185 = (inp[12]) ? node7193 : node7186;
														assign node7186 = (inp[14]) ? node7190 : node7187;
															assign node7187 = (inp[1]) ? 4'b1101 : 4'b1100;
															assign node7190 = (inp[1]) ? 4'b1100 : 4'b1101;
														assign node7193 = (inp[10]) ? node7195 : 4'b0100;
															assign node7195 = (inp[1]) ? node7197 : 4'b0101;
																assign node7197 = (inp[14]) ? 4'b1100 : 4'b1101;
													assign node7200 = (inp[10]) ? node7206 : node7201;
														assign node7201 = (inp[14]) ? 4'b1101 : node7202;
															assign node7202 = (inp[1]) ? 4'b1101 : 4'b1100;
														assign node7206 = (inp[12]) ? node7214 : node7207;
															assign node7207 = (inp[14]) ? node7211 : node7208;
																assign node7208 = (inp[1]) ? 4'b0001 : 4'b0000;
																assign node7211 = (inp[1]) ? 4'b0000 : 4'b0001;
															assign node7214 = (inp[14]) ? node7218 : node7215;
																assign node7215 = (inp[1]) ? 4'b0001 : 4'b0000;
																assign node7218 = (inp[1]) ? 4'b0000 : 4'b1101;
												assign node7221 = (inp[10]) ? node7237 : node7222;
													assign node7222 = (inp[14]) ? node7232 : node7223;
														assign node7223 = (inp[1]) ? 4'b0001 : node7224;
															assign node7224 = (inp[13]) ? node7228 : node7225;
																assign node7225 = (inp[12]) ? 4'b0000 : 4'b1000;
																assign node7228 = (inp[12]) ? 4'b1000 : 4'b0000;
														assign node7232 = (inp[1]) ? 4'b0000 : node7233;
															assign node7233 = (inp[13]) ? 4'b1001 : 4'b0001;
													assign node7237 = (inp[13]) ? node7245 : node7238;
														assign node7238 = (inp[12]) ? node7240 : 4'b1001;
															assign node7240 = (inp[1]) ? node7242 : 4'b1000;
																assign node7242 = (inp[14]) ? 4'b1000 : 4'b1001;
														assign node7245 = (inp[1]) ? node7249 : node7246;
															assign node7246 = (inp[14]) ? 4'b1001 : 4'b0000;
															assign node7249 = (inp[14]) ? 4'b0000 : 4'b0001;
											assign node7252 = (inp[13]) ? node7294 : node7253;
												assign node7253 = (inp[12]) ? node7271 : node7254;
													assign node7254 = (inp[4]) ? node7262 : node7255;
														assign node7255 = (inp[1]) ? node7259 : node7256;
															assign node7256 = (inp[14]) ? 4'b1101 : 4'b1100;
															assign node7259 = (inp[14]) ? 4'b1100 : 4'b1101;
														assign node7262 = (inp[1]) ? node7268 : node7263;
															assign node7263 = (inp[14]) ? node7265 : 4'b1100;
																assign node7265 = (inp[10]) ? 4'b1101 : 4'b0101;
															assign node7268 = (inp[14]) ? 4'b1100 : 4'b1101;
													assign node7271 = (inp[10]) ? node7287 : node7272;
														assign node7272 = (inp[4]) ? node7280 : node7273;
															assign node7273 = (inp[14]) ? node7277 : node7274;
																assign node7274 = (inp[1]) ? 4'b0101 : 4'b0100;
																assign node7277 = (inp[1]) ? 4'b0100 : 4'b0101;
															assign node7280 = (inp[14]) ? node7284 : node7281;
																assign node7281 = (inp[1]) ? 4'b0101 : 4'b0100;
																assign node7284 = (inp[1]) ? 4'b0100 : 4'b0101;
														assign node7287 = (inp[14]) ? node7291 : node7288;
															assign node7288 = (inp[1]) ? 4'b1101 : 4'b1100;
															assign node7291 = (inp[1]) ? 4'b1100 : 4'b0101;
												assign node7294 = (inp[10]) ? node7312 : node7295;
													assign node7295 = (inp[12]) ? node7305 : node7296;
														assign node7296 = (inp[14]) ? node7302 : node7297;
															assign node7297 = (inp[4]) ? 4'b0001 : node7298;
																assign node7298 = (inp[1]) ? 4'b0101 : 4'b0100;
															assign node7302 = (inp[1]) ? 4'b0100 : 4'b1101;
														assign node7305 = (inp[14]) ? node7309 : node7306;
															assign node7306 = (inp[1]) ? 4'b1101 : 4'b1100;
															assign node7309 = (inp[1]) ? 4'b1100 : 4'b1101;
													assign node7312 = (inp[4]) ? node7324 : node7313;
														assign node7313 = (inp[12]) ? node7319 : node7314;
															assign node7314 = (inp[14]) ? node7316 : 4'b0100;
																assign node7316 = (inp[1]) ? 4'b0100 : 4'b0101;
															assign node7319 = (inp[1]) ? node7321 : 4'b0100;
																assign node7321 = (inp[14]) ? 4'b0100 : 4'b0101;
														assign node7324 = (inp[12]) ? node7330 : node7325;
															assign node7325 = (inp[1]) ? 4'b0001 : node7326;
																assign node7326 = (inp[14]) ? 4'b0001 : 4'b0000;
															assign node7330 = (inp[14]) ? 4'b0000 : 4'b0001;
									assign node7333 = (inp[10]) ? node7439 : node7334;
										assign node7334 = (inp[1]) ? node7394 : node7335;
											assign node7335 = (inp[12]) ? node7359 : node7336;
												assign node7336 = (inp[2]) ? node7350 : node7337;
													assign node7337 = (inp[4]) ? node7341 : node7338;
														assign node7338 = (inp[7]) ? 4'b1100 : 4'b1000;
														assign node7341 = (inp[14]) ? node7347 : node7342;
															assign node7342 = (inp[13]) ? 4'b0001 : node7343;
																assign node7343 = (inp[7]) ? 4'b1000 : 4'b1001;
															assign node7347 = (inp[7]) ? 4'b0000 : 4'b0100;
													assign node7350 = (inp[14]) ? node7352 : 4'b1000;
														assign node7352 = (inp[4]) ? 4'b1000 : node7353;
															assign node7353 = (inp[13]) ? node7355 : 4'b0001;
																assign node7355 = (inp[7]) ? 4'b1001 : 4'b1000;
												assign node7359 = (inp[13]) ? node7373 : node7360;
													assign node7360 = (inp[4]) ? node7366 : node7361;
														assign node7361 = (inp[2]) ? node7363 : 4'b0100;
															assign node7363 = (inp[14]) ? 4'b0001 : 4'b0000;
														assign node7366 = (inp[2]) ? 4'b0000 : node7367;
															assign node7367 = (inp[14]) ? 4'b0000 : node7368;
																assign node7368 = (inp[7]) ? 4'b0000 : 4'b0001;
													assign node7373 = (inp[7]) ? node7383 : node7374;
														assign node7374 = (inp[2]) ? node7380 : node7375;
															assign node7375 = (inp[4]) ? node7377 : 4'b0000;
																assign node7377 = (inp[14]) ? 4'b1000 : 4'b1001;
															assign node7380 = (inp[4]) ? 4'b0100 : 4'b0000;
														assign node7383 = (inp[2]) ? node7389 : node7384;
															assign node7384 = (inp[4]) ? node7386 : 4'b0100;
																assign node7386 = (inp[14]) ? 4'b1000 : 4'b1001;
															assign node7389 = (inp[4]) ? 4'b0000 : node7390;
																assign node7390 = (inp[14]) ? 4'b1001 : 4'b1000;
											assign node7394 = (inp[2]) ? node7420 : node7395;
												assign node7395 = (inp[4]) ? node7401 : node7396;
													assign node7396 = (inp[13]) ? node7398 : 4'b1100;
														assign node7398 = (inp[7]) ? 4'b1100 : 4'b1000;
													assign node7401 = (inp[14]) ? node7413 : node7402;
														assign node7402 = (inp[7]) ? node7406 : node7403;
															assign node7403 = (inp[13]) ? 4'b1100 : 4'b0000;
															assign node7406 = (inp[12]) ? node7410 : node7407;
																assign node7407 = (inp[13]) ? 4'b1000 : 4'b0000;
																assign node7410 = (inp[13]) ? 4'b0000 : 4'b1000;
														assign node7413 = (inp[13]) ? node7417 : node7414;
															assign node7414 = (inp[7]) ? 4'b1000 : 4'b1001;
															assign node7417 = (inp[7]) ? 4'b0001 : 4'b0101;
												assign node7420 = (inp[4]) ? node7434 : node7421;
													assign node7421 = (inp[14]) ? node7429 : node7422;
														assign node7422 = (inp[13]) ? node7426 : node7423;
															assign node7423 = (inp[12]) ? 4'b0001 : 4'b1001;
															assign node7426 = (inp[7]) ? 4'b1001 : 4'b1000;
														assign node7429 = (inp[12]) ? node7431 : 4'b1000;
															assign node7431 = (inp[13]) ? 4'b1000 : 4'b0000;
													assign node7434 = (inp[13]) ? node7436 : 4'b1000;
														assign node7436 = (inp[7]) ? 4'b1000 : 4'b1100;
										assign node7439 = (inp[1]) ? node7503 : node7440;
											assign node7440 = (inp[12]) ? node7468 : node7441;
												assign node7441 = (inp[2]) ? node7459 : node7442;
													assign node7442 = (inp[4]) ? node7448 : node7443;
														assign node7443 = (inp[7]) ? node7445 : 4'b0000;
															assign node7445 = (inp[13]) ? 4'b0000 : 4'b0100;
														assign node7448 = (inp[13]) ? node7452 : node7449;
															assign node7449 = (inp[14]) ? 4'b0000 : 4'b0001;
															assign node7452 = (inp[7]) ? node7456 : node7453;
																assign node7453 = (inp[14]) ? 4'b1100 : 4'b1101;
																assign node7456 = (inp[14]) ? 4'b1000 : 4'b1001;
													assign node7459 = (inp[4]) ? node7463 : node7460;
														assign node7460 = (inp[7]) ? 4'b1000 : 4'b0000;
														assign node7463 = (inp[7]) ? node7465 : 4'b0100;
															assign node7465 = (inp[13]) ? 4'b0100 : 4'b0000;
												assign node7468 = (inp[13]) ? node7480 : node7469;
													assign node7469 = (inp[4]) ? node7475 : node7470;
														assign node7470 = (inp[2]) ? node7472 : 4'b1100;
															assign node7472 = (inp[14]) ? 4'b0001 : 4'b1000;
														assign node7475 = (inp[2]) ? 4'b1000 : node7476;
															assign node7476 = (inp[14]) ? 4'b0000 : 4'b0001;
													assign node7480 = (inp[14]) ? node7488 : node7481;
														assign node7481 = (inp[2]) ? node7485 : node7482;
															assign node7482 = (inp[7]) ? 4'b1100 : 4'b1101;
															assign node7485 = (inp[7]) ? 4'b1000 : 4'b1100;
														assign node7488 = (inp[2]) ? node7496 : node7489;
															assign node7489 = (inp[4]) ? node7493 : node7490;
																assign node7490 = (inp[7]) ? 4'b1100 : 4'b1000;
																assign node7493 = (inp[7]) ? 4'b1000 : 4'b1100;
															assign node7496 = (inp[7]) ? node7500 : node7497;
																assign node7497 = (inp[4]) ? 4'b1100 : 4'b1000;
																assign node7500 = (inp[4]) ? 4'b1000 : 4'b1001;
											assign node7503 = (inp[4]) ? node7519 : node7504;
												assign node7504 = (inp[7]) ? node7512 : node7505;
													assign node7505 = (inp[2]) ? 4'b0000 : node7506;
														assign node7506 = (inp[13]) ? node7508 : 4'b0000;
															assign node7508 = (inp[12]) ? 4'b0000 : 4'b0001;
													assign node7512 = (inp[13]) ? 4'b0000 : node7513;
														assign node7513 = (inp[2]) ? node7515 : 4'b0100;
															assign node7515 = (inp[14]) ? 4'b1000 : 4'b1001;
												assign node7519 = (inp[2]) ? node7533 : node7520;
													assign node7520 = (inp[14]) ? node7524 : node7521;
														assign node7521 = (inp[13]) ? 4'b0100 : 4'b1000;
														assign node7524 = (inp[13]) ? node7528 : node7525;
															assign node7525 = (inp[12]) ? 4'b0001 : 4'b1001;
															assign node7528 = (inp[12]) ? node7530 : 4'b0101;
																assign node7530 = (inp[7]) ? 4'b1001 : 4'b1101;
													assign node7533 = (inp[7]) ? node7535 : 4'b0100;
														assign node7535 = (inp[13]) ? 4'b0100 : 4'b0000;
								assign node7538 = (inp[1]) ? node7734 : node7539;
									assign node7539 = (inp[3]) ? node7631 : node7540;
										assign node7540 = (inp[2]) ? node7594 : node7541;
											assign node7541 = (inp[4]) ? node7571 : node7542;
												assign node7542 = (inp[13]) ? node7552 : node7543;
													assign node7543 = (inp[12]) ? node7549 : node7544;
														assign node7544 = (inp[10]) ? node7546 : 4'b1100;
															assign node7546 = (inp[7]) ? 4'b1100 : 4'b0001;
														assign node7549 = (inp[10]) ? 4'b1100 : 4'b0100;
													assign node7552 = (inp[7]) ? node7564 : node7553;
														assign node7553 = (inp[14]) ? node7559 : node7554;
															assign node7554 = (inp[10]) ? 4'b0001 : node7555;
																assign node7555 = (inp[12]) ? 4'b0001 : 4'b1001;
															assign node7559 = (inp[10]) ? node7561 : 4'b1001;
																assign node7561 = (inp[12]) ? 4'b1001 : 4'b0001;
														assign node7564 = (inp[12]) ? node7568 : node7565;
															assign node7565 = (inp[10]) ? 4'b0001 : 4'b0100;
															assign node7568 = (inp[10]) ? 4'b0100 : 4'b1100;
												assign node7571 = (inp[10]) ? node7583 : node7572;
													assign node7572 = (inp[12]) ? node7578 : node7573;
														assign node7573 = (inp[7]) ? 4'b1001 : node7574;
															assign node7574 = (inp[13]) ? 4'b1101 : 4'b1001;
														assign node7578 = (inp[13]) ? node7580 : 4'b0001;
															assign node7580 = (inp[7]) ? 4'b0001 : 4'b0101;
													assign node7583 = (inp[12]) ? node7589 : node7584;
														assign node7584 = (inp[7]) ? node7586 : 4'b0101;
															assign node7586 = (inp[13]) ? 4'b0101 : 4'b0001;
														assign node7589 = (inp[7]) ? 4'b1001 : node7590;
															assign node7590 = (inp[13]) ? 4'b1101 : 4'b1001;
											assign node7594 = (inp[7]) ? node7616 : node7595;
												assign node7595 = (inp[4]) ? node7605 : node7596;
													assign node7596 = (inp[13]) ? node7600 : node7597;
														assign node7597 = (inp[10]) ? 4'b1100 : 4'b0100;
														assign node7600 = (inp[12]) ? node7602 : 4'b0000;
															assign node7602 = (inp[10]) ? 4'b0000 : 4'b1100;
													assign node7605 = (inp[13]) ? node7611 : node7606;
														assign node7606 = (inp[12]) ? node7608 : 4'b1000;
															assign node7608 = (inp[10]) ? 4'b1000 : 4'b0000;
														assign node7611 = (inp[12]) ? node7613 : 4'b0000;
															assign node7613 = (inp[10]) ? 4'b0000 : 4'b1000;
												assign node7616 = (inp[13]) ? node7622 : node7617;
													assign node7617 = (inp[12]) ? node7619 : 4'b1100;
														assign node7619 = (inp[10]) ? 4'b1100 : 4'b0100;
													assign node7622 = (inp[12]) ? node7626 : node7623;
														assign node7623 = (inp[4]) ? 4'b0000 : 4'b0100;
														assign node7626 = (inp[10]) ? node7628 : 4'b1100;
															assign node7628 = (inp[4]) ? 4'b0000 : 4'b0100;
										assign node7631 = (inp[2]) ? node7683 : node7632;
											assign node7632 = (inp[4]) ? node7660 : node7633;
												assign node7633 = (inp[13]) ? node7649 : node7634;
													assign node7634 = (inp[7]) ? node7642 : node7635;
														assign node7635 = (inp[10]) ? node7639 : node7636;
															assign node7636 = (inp[12]) ? 4'b0101 : 4'b1101;
															assign node7639 = (inp[12]) ? 4'b1101 : 4'b0001;
														assign node7642 = (inp[12]) ? node7646 : node7643;
															assign node7643 = (inp[10]) ? 4'b0101 : 4'b1101;
															assign node7646 = (inp[10]) ? 4'b1101 : 4'b0101;
													assign node7649 = (inp[7]) ? node7655 : node7650;
														assign node7650 = (inp[12]) ? node7652 : 4'b0000;
															assign node7652 = (inp[10]) ? 4'b1001 : 4'b0001;
														assign node7655 = (inp[12]) ? 4'b1101 : node7656;
															assign node7656 = (inp[10]) ? 4'b0001 : 4'b1101;
												assign node7660 = (inp[13]) ? node7672 : node7661;
													assign node7661 = (inp[12]) ? node7667 : node7662;
														assign node7662 = (inp[7]) ? node7664 : 4'b1000;
															assign node7664 = (inp[14]) ? 4'b1001 : 4'b1000;
														assign node7667 = (inp[10]) ? 4'b0000 : node7668;
															assign node7668 = (inp[7]) ? 4'b0001 : 4'b1000;
													assign node7672 = (inp[7]) ? node7678 : node7673;
														assign node7673 = (inp[12]) ? node7675 : 4'b0100;
															assign node7675 = (inp[10]) ? 4'b1100 : 4'b0100;
														assign node7678 = (inp[10]) ? node7680 : 4'b0000;
															assign node7680 = (inp[12]) ? 4'b1000 : 4'b0100;
											assign node7683 = (inp[4]) ? node7711 : node7684;
												assign node7684 = (inp[7]) ? node7698 : node7685;
													assign node7685 = (inp[13]) ? node7691 : node7686;
														assign node7686 = (inp[12]) ? node7688 : 4'b0001;
															assign node7688 = (inp[10]) ? 4'b1000 : 4'b0000;
														assign node7691 = (inp[10]) ? node7695 : node7692;
															assign node7692 = (inp[12]) ? 4'b0001 : 4'b1001;
															assign node7695 = (inp[12]) ? 4'b1001 : 4'b0001;
													assign node7698 = (inp[13]) ? node7704 : node7699;
														assign node7699 = (inp[10]) ? 4'b1000 : node7700;
															assign node7700 = (inp[12]) ? 4'b0000 : 4'b1000;
														assign node7704 = (inp[12]) ? node7708 : node7705;
															assign node7705 = (inp[10]) ? 4'b0001 : 4'b0000;
															assign node7708 = (inp[10]) ? 4'b0000 : 4'b1000;
												assign node7711 = (inp[7]) ? node7725 : node7712;
													assign node7712 = (inp[13]) ? node7720 : node7713;
														assign node7713 = (inp[12]) ? node7717 : node7714;
															assign node7714 = (inp[10]) ? 4'b0101 : 4'b1001;
															assign node7717 = (inp[10]) ? 4'b1001 : 4'b0001;
														assign node7720 = (inp[10]) ? node7722 : 4'b0101;
															assign node7722 = (inp[12]) ? 4'b1101 : 4'b0101;
													assign node7725 = (inp[10]) ? node7729 : node7726;
														assign node7726 = (inp[12]) ? 4'b0001 : 4'b1001;
														assign node7729 = (inp[12]) ? 4'b1001 : node7730;
															assign node7730 = (inp[13]) ? 4'b0101 : 4'b0001;
									assign node7734 = (inp[10]) ? node7806 : node7735;
										assign node7735 = (inp[3]) ? node7769 : node7736;
											assign node7736 = (inp[4]) ? node7754 : node7737;
												assign node7737 = (inp[7]) ? node7747 : node7738;
													assign node7738 = (inp[13]) ? node7742 : node7739;
														assign node7739 = (inp[12]) ? 4'b0101 : 4'b1101;
														assign node7742 = (inp[2]) ? node7744 : 4'b1001;
															assign node7744 = (inp[12]) ? 4'b1101 : 4'b0001;
													assign node7747 = (inp[12]) ? node7751 : node7748;
														assign node7748 = (inp[13]) ? 4'b0101 : 4'b1101;
														assign node7751 = (inp[13]) ? 4'b1101 : 4'b0101;
												assign node7754 = (inp[2]) ? node7760 : node7755;
													assign node7755 = (inp[13]) ? node7757 : 4'b1001;
														assign node7757 = (inp[7]) ? 4'b1001 : 4'b1101;
													assign node7760 = (inp[13]) ? node7764 : node7761;
														assign node7761 = (inp[12]) ? 4'b0101 : 4'b1101;
														assign node7764 = (inp[12]) ? node7766 : 4'b0001;
															assign node7766 = (inp[7]) ? 4'b1101 : 4'b1001;
											assign node7769 = (inp[2]) ? node7791 : node7770;
												assign node7770 = (inp[4]) ? node7776 : node7771;
													assign node7771 = (inp[13]) ? node7773 : 4'b1101;
														assign node7773 = (inp[7]) ? 4'b1101 : 4'b1001;
													assign node7776 = (inp[7]) ? node7784 : node7777;
														assign node7777 = (inp[13]) ? node7781 : node7778;
															assign node7778 = (inp[12]) ? 4'b1001 : 4'b0001;
															assign node7781 = (inp[12]) ? 4'b0101 : 4'b1101;
														assign node7784 = (inp[13]) ? node7788 : node7785;
															assign node7785 = (inp[12]) ? 4'b1001 : 4'b0001;
															assign node7788 = (inp[12]) ? 4'b0001 : 4'b1001;
												assign node7791 = (inp[4]) ? node7801 : node7792;
													assign node7792 = (inp[13]) ? node7796 : node7793;
														assign node7793 = (inp[12]) ? 4'b0001 : 4'b1001;
														assign node7796 = (inp[12]) ? 4'b1001 : node7797;
															assign node7797 = (inp[14]) ? 4'b0001 : 4'b1001;
													assign node7801 = (inp[7]) ? 4'b1001 : node7802;
														assign node7802 = (inp[13]) ? 4'b1101 : 4'b1001;
										assign node7806 = (inp[13]) ? node7832 : node7807;
											assign node7807 = (inp[2]) ? node7819 : node7808;
												assign node7808 = (inp[4]) ? node7814 : node7809;
													assign node7809 = (inp[7]) ? node7811 : 4'b0001;
														assign node7811 = (inp[3]) ? 4'b0101 : 4'b1101;
													assign node7814 = (inp[3]) ? 4'b1001 : node7815;
														assign node7815 = (inp[7]) ? 4'b0001 : 4'b0101;
												assign node7819 = (inp[3]) ? node7825 : node7820;
													assign node7820 = (inp[4]) ? node7822 : 4'b1101;
														assign node7822 = (inp[7]) ? 4'b1101 : 4'b1001;
													assign node7825 = (inp[4]) ? node7829 : node7826;
														assign node7826 = (inp[7]) ? 4'b1001 : 4'b0001;
														assign node7829 = (inp[7]) ? 4'b0001 : 4'b0101;
											assign node7832 = (inp[4]) ? node7840 : node7833;
												assign node7833 = (inp[2]) ? node7835 : 4'b0001;
													assign node7835 = (inp[7]) ? node7837 : 4'b0001;
														assign node7837 = (inp[3]) ? 4'b0001 : 4'b0101;
												assign node7840 = (inp[2]) ? node7842 : 4'b0101;
													assign node7842 = (inp[3]) ? 4'b0101 : 4'b0001;
							assign node7845 = (inp[2]) ? 4'b0101 : node7846;
								assign node7846 = (inp[3]) ? node7954 : node7847;
									assign node7847 = (inp[4]) ? node7875 : node7848;
										assign node7848 = (inp[13]) ? node7850 : 4'b0101;
											assign node7850 = (inp[7]) ? 4'b0101 : node7851;
												assign node7851 = (inp[12]) ? node7865 : node7852;
													assign node7852 = (inp[1]) ? node7860 : node7853;
														assign node7853 = (inp[14]) ? node7855 : 4'b0000;
															assign node7855 = (inp[11]) ? 4'b0000 : node7856;
																assign node7856 = (inp[10]) ? 4'b0001 : 4'b0101;
														assign node7860 = (inp[14]) ? node7862 : 4'b0001;
															assign node7862 = (inp[11]) ? 4'b0001 : 4'b0000;
													assign node7865 = (inp[10]) ? node7867 : 4'b0101;
														assign node7867 = (inp[11]) ? 4'b0001 : node7868;
															assign node7868 = (inp[14]) ? node7870 : 4'b0000;
																assign node7870 = (inp[1]) ? 4'b0000 : 4'b0101;
										assign node7875 = (inp[7]) ? node7929 : node7876;
											assign node7876 = (inp[1]) ? node7904 : node7877;
												assign node7877 = (inp[14]) ? node7889 : node7878;
													assign node7878 = (inp[13]) ? node7884 : node7879;
														assign node7879 = (inp[12]) ? node7881 : 4'b1000;
															assign node7881 = (inp[10]) ? 4'b1000 : 4'b0000;
														assign node7884 = (inp[10]) ? 4'b0000 : node7885;
															assign node7885 = (inp[12]) ? 4'b1000 : 4'b0000;
													assign node7889 = (inp[11]) ? node7901 : node7890;
														assign node7890 = (inp[13]) ? node7896 : node7891;
															assign node7891 = (inp[12]) ? 4'b0001 : node7892;
																assign node7892 = (inp[10]) ? 4'b1001 : 4'b0001;
															assign node7896 = (inp[10]) ? node7898 : 4'b1001;
																assign node7898 = (inp[12]) ? 4'b1001 : 4'b0001;
														assign node7901 = (inp[10]) ? 4'b0000 : 4'b1000;
												assign node7904 = (inp[13]) ? node7916 : node7905;
													assign node7905 = (inp[10]) ? 4'b1001 : node7906;
														assign node7906 = (inp[12]) ? node7910 : node7907;
															assign node7907 = (inp[14]) ? 4'b1000 : 4'b1001;
															assign node7910 = (inp[14]) ? node7912 : 4'b0001;
																assign node7912 = (inp[11]) ? 4'b0001 : 4'b0000;
													assign node7916 = (inp[14]) ? node7922 : node7917;
														assign node7917 = (inp[12]) ? node7919 : 4'b0001;
															assign node7919 = (inp[10]) ? 4'b0001 : 4'b1001;
														assign node7922 = (inp[11]) ? 4'b0001 : node7923;
															assign node7923 = (inp[12]) ? node7925 : 4'b0000;
																assign node7925 = (inp[10]) ? 4'b0000 : 4'b1000;
											assign node7929 = (inp[13]) ? node7931 : 4'b0101;
												assign node7931 = (inp[10]) ? node7941 : node7932;
													assign node7932 = (inp[12]) ? 4'b0101 : node7933;
														assign node7933 = (inp[1]) ? 4'b0001 : node7934;
															assign node7934 = (inp[11]) ? 4'b0000 : node7935;
																assign node7935 = (inp[14]) ? 4'b0101 : 4'b0000;
													assign node7941 = (inp[1]) ? node7949 : node7942;
														assign node7942 = (inp[14]) ? node7944 : 4'b0000;
															assign node7944 = (inp[11]) ? 4'b0000 : node7945;
																assign node7945 = (inp[12]) ? 4'b0101 : 4'b0001;
														assign node7949 = (inp[12]) ? node7951 : 4'b0001;
															assign node7951 = (inp[11]) ? 4'b0001 : 4'b0000;
									assign node7954 = (inp[1]) ? node8042 : node7955;
										assign node7955 = (inp[11]) ? node8007 : node7956;
											assign node7956 = (inp[14]) ? node7980 : node7957;
												assign node7957 = (inp[13]) ? node7967 : node7958;
													assign node7958 = (inp[12]) ? node7960 : 4'b1000;
														assign node7960 = (inp[10]) ? 4'b1000 : node7961;
															assign node7961 = (inp[4]) ? node7963 : 4'b0000;
																assign node7963 = (inp[7]) ? 4'b0000 : 4'b0100;
													assign node7967 = (inp[7]) ? node7973 : node7968;
														assign node7968 = (inp[12]) ? node7970 : 4'b0100;
															assign node7970 = (inp[10]) ? 4'b0100 : 4'b1100;
														assign node7973 = (inp[12]) ? node7977 : node7974;
															assign node7974 = (inp[4]) ? 4'b0100 : 4'b0000;
															assign node7977 = (inp[10]) ? 4'b0000 : 4'b1000;
												assign node7980 = (inp[4]) ? node7992 : node7981;
													assign node7981 = (inp[13]) ? node7987 : node7982;
														assign node7982 = (inp[10]) ? node7984 : 4'b0001;
															assign node7984 = (inp[12]) ? 4'b0001 : 4'b1001;
														assign node7987 = (inp[10]) ? node7989 : 4'b1001;
															assign node7989 = (inp[12]) ? 4'b1001 : 4'b0001;
													assign node7992 = (inp[7]) ? node8000 : node7993;
														assign node7993 = (inp[13]) ? node7995 : 4'b0101;
															assign node7995 = (inp[10]) ? node7997 : 4'b1101;
																assign node7997 = (inp[12]) ? 4'b1101 : 4'b0101;
														assign node8000 = (inp[10]) ? node8004 : node8001;
															assign node8001 = (inp[13]) ? 4'b1001 : 4'b0001;
															assign node8004 = (inp[13]) ? 4'b0101 : 4'b1001;
											assign node8007 = (inp[13]) ? node8025 : node8008;
												assign node8008 = (inp[12]) ? node8014 : node8009;
													assign node8009 = (inp[7]) ? 4'b1000 : node8010;
														assign node8010 = (inp[4]) ? 4'b1100 : 4'b1000;
													assign node8014 = (inp[10]) ? node8020 : node8015;
														assign node8015 = (inp[7]) ? 4'b0000 : node8016;
															assign node8016 = (inp[4]) ? 4'b0100 : 4'b0000;
														assign node8020 = (inp[14]) ? node8022 : 4'b1000;
															assign node8022 = (inp[4]) ? 4'b1100 : 4'b1000;
												assign node8025 = (inp[12]) ? node8031 : node8026;
													assign node8026 = (inp[7]) ? node8028 : 4'b0100;
														assign node8028 = (inp[4]) ? 4'b0100 : 4'b0000;
													assign node8031 = (inp[10]) ? node8037 : node8032;
														assign node8032 = (inp[7]) ? 4'b1000 : node8033;
															assign node8033 = (inp[4]) ? 4'b1100 : 4'b1000;
														assign node8037 = (inp[7]) ? node8039 : 4'b0100;
															assign node8039 = (inp[4]) ? 4'b0100 : 4'b0000;
										assign node8042 = (inp[13]) ? node8080 : node8043;
											assign node8043 = (inp[14]) ? node8055 : node8044;
												assign node8044 = (inp[4]) ? node8050 : node8045;
													assign node8045 = (inp[12]) ? node8047 : 4'b1001;
														assign node8047 = (inp[10]) ? 4'b1001 : 4'b0001;
													assign node8050 = (inp[7]) ? node8052 : 4'b1101;
														assign node8052 = (inp[12]) ? 4'b0001 : 4'b1001;
												assign node8055 = (inp[11]) ? node8069 : node8056;
													assign node8056 = (inp[7]) ? node8064 : node8057;
														assign node8057 = (inp[4]) ? node8059 : 4'b1000;
															assign node8059 = (inp[10]) ? 4'b1100 : node8060;
																assign node8060 = (inp[12]) ? 4'b0100 : 4'b1100;
														assign node8064 = (inp[10]) ? 4'b1000 : node8065;
															assign node8065 = (inp[12]) ? 4'b0000 : 4'b1000;
													assign node8069 = (inp[10]) ? node8073 : node8070;
														assign node8070 = (inp[12]) ? 4'b0001 : 4'b1001;
														assign node8073 = (inp[12]) ? 4'b1101 : node8074;
															assign node8074 = (inp[4]) ? node8076 : 4'b1001;
																assign node8076 = (inp[7]) ? 4'b1001 : 4'b1101;
											assign node8080 = (inp[10]) ? node8104 : node8081;
												assign node8081 = (inp[12]) ? node8091 : node8082;
													assign node8082 = (inp[14]) ? node8088 : node8083;
														assign node8083 = (inp[7]) ? node8085 : 4'b0101;
															assign node8085 = (inp[11]) ? 4'b0001 : 4'b0101;
														assign node8088 = (inp[11]) ? 4'b0101 : 4'b0100;
													assign node8091 = (inp[4]) ? node8097 : node8092;
														assign node8092 = (inp[11]) ? 4'b1001 : node8093;
															assign node8093 = (inp[14]) ? 4'b1000 : 4'b1001;
														assign node8097 = (inp[7]) ? 4'b1001 : node8098;
															assign node8098 = (inp[14]) ? node8100 : 4'b1101;
																assign node8100 = (inp[11]) ? 4'b1101 : 4'b1100;
												assign node8104 = (inp[7]) ? node8110 : node8105;
													assign node8105 = (inp[14]) ? node8107 : 4'b0101;
														assign node8107 = (inp[11]) ? 4'b0101 : 4'b0100;
													assign node8110 = (inp[4]) ? 4'b0101 : node8111;
														assign node8111 = (inp[14]) ? 4'b0000 : 4'b0001;
						assign node8116 = (inp[3]) ? node8820 : node8117;
							assign node8117 = (inp[4]) ? node8443 : node8118;
								assign node8118 = (inp[13]) ? node8270 : node8119;
									assign node8119 = (inp[0]) ? node8225 : node8120;
										assign node8120 = (inp[10]) ? node8166 : node8121;
											assign node8121 = (inp[11]) ? node8151 : node8122;
												assign node8122 = (inp[2]) ? node8140 : node8123;
													assign node8123 = (inp[12]) ? node8133 : node8124;
														assign node8124 = (inp[1]) ? node8128 : node8125;
															assign node8125 = (inp[14]) ? 4'b1100 : 4'b1101;
															assign node8128 = (inp[7]) ? node8130 : 4'b0001;
																assign node8130 = (inp[14]) ? 4'b1101 : 4'b0100;
														assign node8133 = (inp[1]) ? node8137 : node8134;
															assign node8134 = (inp[14]) ? 4'b0100 : 4'b0101;
															assign node8137 = (inp[14]) ? 4'b1101 : 4'b1100;
													assign node8140 = (inp[12]) ? node8148 : node8141;
														assign node8141 = (inp[14]) ? 4'b1100 : node8142;
															assign node8142 = (inp[1]) ? node8144 : 4'b1100;
																assign node8144 = (inp[7]) ? 4'b1100 : 4'b0000;
														assign node8148 = (inp[1]) ? 4'b1100 : 4'b0100;
												assign node8151 = (inp[1]) ? node8157 : node8152;
													assign node8152 = (inp[2]) ? node8154 : 4'b1100;
														assign node8154 = (inp[12]) ? 4'b0101 : 4'b1101;
													assign node8157 = (inp[2]) ? node8161 : node8158;
														assign node8158 = (inp[7]) ? 4'b0101 : 4'b0001;
														assign node8161 = (inp[14]) ? node8163 : 4'b1101;
															assign node8163 = (inp[7]) ? 4'b1101 : 4'b0001;
											assign node8166 = (inp[7]) ? node8198 : node8167;
												assign node8167 = (inp[2]) ? node8185 : node8168;
													assign node8168 = (inp[12]) ? node8172 : node8169;
														assign node8169 = (inp[1]) ? 4'b0001 : 4'b1001;
														assign node8172 = (inp[14]) ? node8180 : node8173;
															assign node8173 = (inp[1]) ? node8177 : node8174;
																assign node8174 = (inp[11]) ? 4'b1001 : 4'b0001;
																assign node8177 = (inp[11]) ? 4'b0001 : 4'b1001;
															assign node8180 = (inp[11]) ? 4'b1001 : node8181;
																assign node8181 = (inp[1]) ? 4'b1001 : 4'b0001;
													assign node8185 = (inp[1]) ? node8191 : node8186;
														assign node8186 = (inp[14]) ? 4'b0000 : node8187;
															assign node8187 = (inp[11]) ? 4'b1000 : 4'b0001;
														assign node8191 = (inp[11]) ? 4'b1001 : node8192;
															assign node8192 = (inp[14]) ? node8194 : 4'b1000;
																assign node8194 = (inp[12]) ? 4'b0001 : 4'b1001;
												assign node8198 = (inp[1]) ? node8214 : node8199;
													assign node8199 = (inp[2]) ? node8207 : node8200;
														assign node8200 = (inp[11]) ? node8204 : node8201;
															assign node8201 = (inp[14]) ? 4'b0100 : 4'b0101;
															assign node8204 = (inp[12]) ? 4'b0100 : 4'b1100;
														assign node8207 = (inp[12]) ? node8211 : node8208;
															assign node8208 = (inp[11]) ? 4'b0101 : 4'b0100;
															assign node8211 = (inp[11]) ? 4'b1101 : 4'b1100;
													assign node8214 = (inp[2]) ? node8222 : node8215;
														assign node8215 = (inp[11]) ? 4'b0001 : node8216;
															assign node8216 = (inp[12]) ? node8218 : 4'b0001;
																assign node8218 = (inp[14]) ? 4'b0101 : 4'b1100;
														assign node8222 = (inp[11]) ? 4'b0101 : 4'b0100;
										assign node8225 = (inp[2]) ? 4'b0101 : node8226;
											assign node8226 = (inp[1]) ? node8248 : node8227;
												assign node8227 = (inp[14]) ? node8233 : node8228;
													assign node8228 = (inp[12]) ? node8230 : 4'b1100;
														assign node8230 = (inp[10]) ? 4'b1100 : 4'b0100;
													assign node8233 = (inp[11]) ? node8239 : node8234;
														assign node8234 = (inp[10]) ? node8236 : 4'b0101;
															assign node8236 = (inp[7]) ? 4'b1101 : 4'b0000;
														assign node8239 = (inp[12]) ? node8245 : node8240;
															assign node8240 = (inp[7]) ? 4'b1100 : node8241;
																assign node8241 = (inp[10]) ? 4'b0001 : 4'b1100;
															assign node8245 = (inp[10]) ? 4'b1100 : 4'b0100;
												assign node8248 = (inp[7]) ? node8256 : node8249;
													assign node8249 = (inp[10]) ? node8253 : node8250;
														assign node8250 = (inp[11]) ? 4'b0101 : 4'b1101;
														assign node8253 = (inp[11]) ? 4'b0001 : 4'b0000;
													assign node8256 = (inp[10]) ? node8264 : node8257;
														assign node8257 = (inp[12]) ? node8259 : 4'b1101;
															assign node8259 = (inp[14]) ? node8261 : 4'b0101;
																assign node8261 = (inp[11]) ? 4'b0101 : 4'b0100;
														assign node8264 = (inp[14]) ? node8266 : 4'b1101;
															assign node8266 = (inp[12]) ? 4'b1101 : 4'b1100;
									assign node8270 = (inp[1]) ? node8356 : node8271;
										assign node8271 = (inp[0]) ? node8309 : node8272;
											assign node8272 = (inp[2]) ? node8290 : node8273;
												assign node8273 = (inp[11]) ? node8285 : node8274;
													assign node8274 = (inp[12]) ? node8280 : node8275;
														assign node8275 = (inp[10]) ? node8277 : 4'b1001;
															assign node8277 = (inp[7]) ? 4'b1001 : 4'b1101;
														assign node8280 = (inp[7]) ? 4'b0001 : node8281;
															assign node8281 = (inp[10]) ? 4'b0101 : 4'b0001;
													assign node8285 = (inp[7]) ? 4'b1001 : node8286;
														assign node8286 = (inp[10]) ? 4'b1101 : 4'b1001;
												assign node8290 = (inp[10]) ? node8298 : node8291;
													assign node8291 = (inp[11]) ? 4'b0000 : node8292;
														assign node8292 = (inp[7]) ? 4'b0100 : node8293;
															assign node8293 = (inp[12]) ? 4'b1001 : 4'b0000;
													assign node8298 = (inp[14]) ? node8304 : node8299;
														assign node8299 = (inp[11]) ? node8301 : 4'b1001;
															assign node8301 = (inp[12]) ? 4'b1000 : 4'b0100;
														assign node8304 = (inp[12]) ? 4'b1000 : node8305;
															assign node8305 = (inp[11]) ? 4'b0000 : 4'b1000;
											assign node8309 = (inp[7]) ? node8333 : node8310;
												assign node8310 = (inp[2]) ? node8326 : node8311;
													assign node8311 = (inp[11]) ? node8319 : node8312;
														assign node8312 = (inp[12]) ? node8316 : node8313;
															assign node8313 = (inp[10]) ? 4'b0000 : 4'b1000;
															assign node8316 = (inp[10]) ? 4'b1000 : 4'b0000;
														assign node8319 = (inp[12]) ? node8323 : node8320;
															assign node8320 = (inp[10]) ? 4'b0001 : 4'b1001;
															assign node8323 = (inp[10]) ? 4'b1001 : 4'b0001;
													assign node8326 = (inp[11]) ? node8328 : 4'b0101;
														assign node8328 = (inp[10]) ? 4'b0000 : node8329;
															assign node8329 = (inp[12]) ? 4'b0101 : 4'b0000;
												assign node8333 = (inp[2]) ? 4'b0101 : node8334;
													assign node8334 = (inp[10]) ? node8346 : node8335;
														assign node8335 = (inp[12]) ? node8341 : node8336;
															assign node8336 = (inp[14]) ? node8338 : 4'b0100;
																assign node8338 = (inp[11]) ? 4'b0100 : 4'b1101;
															assign node8341 = (inp[11]) ? 4'b1100 : node8342;
																assign node8342 = (inp[14]) ? 4'b1101 : 4'b1100;
														assign node8346 = (inp[12]) ? node8350 : node8347;
															assign node8347 = (inp[14]) ? 4'b0001 : 4'b0000;
															assign node8350 = (inp[14]) ? node8352 : 4'b0100;
																assign node8352 = (inp[11]) ? 4'b0100 : 4'b1101;
										assign node8356 = (inp[11]) ? node8408 : node8357;
											assign node8357 = (inp[0]) ? node8395 : node8358;
												assign node8358 = (inp[12]) ? node8382 : node8359;
													assign node8359 = (inp[2]) ? node8373 : node8360;
														assign node8360 = (inp[14]) ? node8368 : node8361;
															assign node8361 = (inp[7]) ? node8365 : node8362;
																assign node8362 = (inp[10]) ? 4'b0001 : 4'b0101;
																assign node8365 = (inp[10]) ? 4'b0101 : 4'b0001;
															assign node8368 = (inp[7]) ? node8370 : 4'b0000;
																assign node8370 = (inp[10]) ? 4'b0101 : 4'b0001;
														assign node8373 = (inp[14]) ? node8379 : node8374;
															assign node8374 = (inp[7]) ? node8376 : 4'b0100;
																assign node8376 = (inp[10]) ? 4'b0000 : 4'b1000;
															assign node8379 = (inp[10]) ? 4'b0101 : 4'b0001;
													assign node8382 = (inp[2]) ? node8388 : node8383;
														assign node8383 = (inp[14]) ? 4'b1001 : node8384;
															assign node8384 = (inp[10]) ? 4'b1101 : 4'b1001;
														assign node8388 = (inp[14]) ? node8392 : node8389;
															assign node8389 = (inp[10]) ? 4'b0100 : 4'b0000;
															assign node8392 = (inp[10]) ? 4'b1001 : 4'b0001;
												assign node8395 = (inp[2]) ? node8401 : node8396;
													assign node8396 = (inp[10]) ? 4'b0000 : node8397;
														assign node8397 = (inp[7]) ? 4'b1100 : 4'b1000;
													assign node8401 = (inp[7]) ? 4'b0101 : node8402;
														assign node8402 = (inp[12]) ? node8404 : 4'b0000;
															assign node8404 = (inp[10]) ? 4'b0000 : 4'b0101;
											assign node8408 = (inp[10]) ? node8430 : node8409;
												assign node8409 = (inp[0]) ? node8419 : node8410;
													assign node8410 = (inp[7]) ? node8414 : node8411;
														assign node8411 = (inp[2]) ? 4'b0001 : 4'b0101;
														assign node8414 = (inp[12]) ? 4'b0001 : node8415;
															assign node8415 = (inp[2]) ? 4'b1001 : 4'b0001;
													assign node8419 = (inp[2]) ? node8425 : node8420;
														assign node8420 = (inp[7]) ? node8422 : 4'b1001;
															assign node8422 = (inp[12]) ? 4'b1101 : 4'b0101;
														assign node8425 = (inp[12]) ? 4'b0101 : node8426;
															assign node8426 = (inp[7]) ? 4'b0101 : 4'b0001;
												assign node8430 = (inp[2]) ? node8436 : node8431;
													assign node8431 = (inp[7]) ? node8433 : 4'b0001;
														assign node8433 = (inp[0]) ? 4'b0001 : 4'b0101;
													assign node8436 = (inp[7]) ? node8440 : node8437;
														assign node8437 = (inp[0]) ? 4'b0001 : 4'b0101;
														assign node8440 = (inp[0]) ? 4'b0101 : 4'b0001;
								assign node8443 = (inp[1]) ? node8651 : node8444;
									assign node8444 = (inp[7]) ? node8560 : node8445;
										assign node8445 = (inp[0]) ? node8495 : node8446;
											assign node8446 = (inp[2]) ? node8468 : node8447;
												assign node8447 = (inp[10]) ? node8457 : node8448;
													assign node8448 = (inp[12]) ? 4'b1000 : node8449;
														assign node8449 = (inp[11]) ? node8453 : node8450;
															assign node8450 = (inp[13]) ? 4'b1000 : 4'b1001;
															assign node8453 = (inp[13]) ? 4'b0001 : 4'b0000;
													assign node8457 = (inp[11]) ? node8463 : node8458;
														assign node8458 = (inp[13]) ? node8460 : 4'b1001;
															assign node8460 = (inp[12]) ? 4'b0100 : 4'b0001;
														assign node8463 = (inp[13]) ? node8465 : 4'b0100;
															assign node8465 = (inp[12]) ? 4'b0000 : 4'b1000;
												assign node8468 = (inp[11]) ? node8488 : node8469;
													assign node8469 = (inp[12]) ? node8481 : node8470;
														assign node8470 = (inp[13]) ? node8474 : node8471;
															assign node8471 = (inp[10]) ? 4'b1001 : 4'b1101;
															assign node8474 = (inp[14]) ? node8478 : node8475;
																assign node8475 = (inp[10]) ? 4'b1000 : 4'b1001;
																assign node8478 = (inp[10]) ? 4'b0001 : 4'b1001;
														assign node8481 = (inp[10]) ? 4'b0001 : node8482;
															assign node8482 = (inp[14]) ? 4'b0100 : node8483;
																assign node8483 = (inp[13]) ? 4'b0001 : 4'b0101;
													assign node8488 = (inp[10]) ? node8492 : node8489;
														assign node8489 = (inp[13]) ? 4'b1001 : 4'b1100;
														assign node8492 = (inp[13]) ? 4'b1000 : 4'b1001;
											assign node8495 = (inp[10]) ? node8525 : node8496;
												assign node8496 = (inp[12]) ? node8510 : node8497;
													assign node8497 = (inp[13]) ? node8503 : node8498;
														assign node8498 = (inp[2]) ? 4'b1000 : node8499;
															assign node8499 = (inp[11]) ? 4'b1001 : 4'b1000;
														assign node8503 = (inp[14]) ? node8505 : 4'b0000;
															assign node8505 = (inp[11]) ? 4'b0000 : node8506;
																assign node8506 = (inp[2]) ? 4'b1001 : 4'b0000;
													assign node8510 = (inp[13]) ? node8520 : node8511;
														assign node8511 = (inp[14]) ? node8513 : 4'b0000;
															assign node8513 = (inp[11]) ? node8517 : node8514;
																assign node8514 = (inp[2]) ? 4'b0001 : 4'b0000;
																assign node8517 = (inp[2]) ? 4'b0000 : 4'b0001;
														assign node8520 = (inp[2]) ? 4'b1000 : node8521;
															assign node8521 = (inp[11]) ? 4'b0000 : 4'b0100;
												assign node8525 = (inp[2]) ? node8545 : node8526;
													assign node8526 = (inp[12]) ? node8536 : node8527;
														assign node8527 = (inp[13]) ? node8531 : node8528;
															assign node8528 = (inp[14]) ? 4'b0100 : 4'b0101;
															assign node8531 = (inp[11]) ? 4'b0000 : node8532;
																assign node8532 = (inp[14]) ? 4'b1000 : 4'b1001;
														assign node8536 = (inp[11]) ? node8542 : node8537;
															assign node8537 = (inp[14]) ? 4'b1000 : node8538;
																assign node8538 = (inp[13]) ? 4'b1001 : 4'b1000;
															assign node8542 = (inp[13]) ? 4'b1000 : 4'b1001;
													assign node8545 = (inp[13]) ? node8553 : node8546;
														assign node8546 = (inp[11]) ? 4'b1000 : node8547;
															assign node8547 = (inp[14]) ? node8549 : 4'b1000;
																assign node8549 = (inp[12]) ? 4'b0001 : 4'b1001;
														assign node8553 = (inp[14]) ? node8555 : 4'b0000;
															assign node8555 = (inp[11]) ? 4'b0000 : node8556;
																assign node8556 = (inp[12]) ? 4'b1001 : 4'b0001;
										assign node8560 = (inp[2]) ? node8622 : node8561;
											assign node8561 = (inp[11]) ? node8587 : node8562;
												assign node8562 = (inp[0]) ? node8578 : node8563;
													assign node8563 = (inp[10]) ? node8571 : node8564;
														assign node8564 = (inp[12]) ? node8568 : node8565;
															assign node8565 = (inp[13]) ? 4'b0101 : 4'b1101;
															assign node8568 = (inp[13]) ? 4'b1001 : 4'b0101;
														assign node8571 = (inp[13]) ? 4'b0000 : node8572;
															assign node8572 = (inp[14]) ? 4'b1001 : node8573;
																assign node8573 = (inp[12]) ? 4'b1000 : 4'b0000;
													assign node8578 = (inp[10]) ? node8582 : node8579;
														assign node8579 = (inp[12]) ? 4'b0000 : 4'b1000;
														assign node8582 = (inp[12]) ? 4'b1000 : node8583;
															assign node8583 = (inp[13]) ? 4'b0100 : 4'b0000;
												assign node8587 = (inp[0]) ? node8599 : node8588;
													assign node8588 = (inp[13]) ? node8594 : node8589;
														assign node8589 = (inp[12]) ? node8591 : 4'b0000;
															assign node8591 = (inp[14]) ? 4'b0000 : 4'b1101;
														assign node8594 = (inp[12]) ? node8596 : 4'b0001;
															assign node8596 = (inp[10]) ? 4'b0001 : 4'b0100;
													assign node8599 = (inp[13]) ? node8615 : node8600;
														assign node8600 = (inp[14]) ? node8608 : node8601;
															assign node8601 = (inp[12]) ? node8605 : node8602;
																assign node8602 = (inp[10]) ? 4'b0001 : 4'b1001;
																assign node8605 = (inp[10]) ? 4'b1001 : 4'b0001;
															assign node8608 = (inp[10]) ? node8612 : node8609;
																assign node8609 = (inp[12]) ? 4'b0001 : 4'b1001;
																assign node8612 = (inp[12]) ? 4'b1001 : 4'b0001;
														assign node8615 = (inp[12]) ? node8619 : node8616;
															assign node8616 = (inp[10]) ? 4'b0000 : 4'b1001;
															assign node8619 = (inp[10]) ? 4'b1001 : 4'b0001;
											assign node8622 = (inp[0]) ? node8642 : node8623;
												assign node8623 = (inp[13]) ? node8637 : node8624;
													assign node8624 = (inp[10]) ? node8630 : node8625;
														assign node8625 = (inp[11]) ? 4'b1000 : node8626;
															assign node8626 = (inp[12]) ? 4'b0000 : 4'b1001;
														assign node8630 = (inp[11]) ? node8634 : node8631;
															assign node8631 = (inp[14]) ? 4'b0100 : 4'b0101;
															assign node8634 = (inp[12]) ? 4'b0100 : 4'b1100;
													assign node8637 = (inp[11]) ? 4'b1001 : node8638;
														assign node8638 = (inp[12]) ? 4'b0001 : 4'b1001;
												assign node8642 = (inp[13]) ? node8644 : 4'b0101;
													assign node8644 = (inp[10]) ? 4'b0000 : node8645;
														assign node8645 = (inp[12]) ? 4'b0101 : node8646;
															assign node8646 = (inp[11]) ? 4'b0000 : 4'b0101;
									assign node8651 = (inp[11]) ? node8767 : node8652;
										assign node8652 = (inp[2]) ? node8710 : node8653;
											assign node8653 = (inp[10]) ? node8671 : node8654;
												assign node8654 = (inp[0]) ? node8662 : node8655;
													assign node8655 = (inp[13]) ? node8659 : node8656;
														assign node8656 = (inp[14]) ? 4'b0000 : 4'b0001;
														assign node8659 = (inp[12]) ? 4'b0000 : 4'b1000;
													assign node8662 = (inp[13]) ? node8664 : 4'b1000;
														assign node8664 = (inp[7]) ? 4'b1000 : node8665;
															assign node8665 = (inp[14]) ? 4'b0001 : node8666;
																assign node8666 = (inp[12]) ? 4'b0000 : 4'b1000;
												assign node8671 = (inp[0]) ? node8697 : node8672;
													assign node8672 = (inp[13]) ? node8686 : node8673;
														assign node8673 = (inp[14]) ? node8681 : node8674;
															assign node8674 = (inp[7]) ? node8678 : node8675;
																assign node8675 = (inp[12]) ? 4'b0101 : 4'b0000;
																assign node8678 = (inp[12]) ? 4'b0001 : 4'b1001;
															assign node8681 = (inp[12]) ? 4'b0000 : node8682;
																assign node8682 = (inp[7]) ? 4'b1000 : 4'b0000;
														assign node8686 = (inp[12]) ? node8694 : node8687;
															assign node8687 = (inp[7]) ? node8691 : node8688;
																assign node8688 = (inp[14]) ? 4'b1001 : 4'b0000;
																assign node8691 = (inp[14]) ? 4'b0100 : 4'b0000;
															assign node8694 = (inp[14]) ? 4'b1001 : 4'b1000;
													assign node8697 = (inp[13]) ? node8701 : node8698;
														assign node8698 = (inp[7]) ? 4'b0000 : 4'b0100;
														assign node8701 = (inp[14]) ? node8703 : 4'b0000;
															assign node8703 = (inp[7]) ? node8707 : node8704;
																assign node8704 = (inp[12]) ? 4'b1001 : 4'b0001;
																assign node8707 = (inp[12]) ? 4'b0100 : 4'b0001;
											assign node8710 = (inp[12]) ? node8736 : node8711;
												assign node8711 = (inp[14]) ? node8729 : node8712;
													assign node8712 = (inp[7]) ? node8722 : node8713;
														assign node8713 = (inp[13]) ? node8717 : node8714;
															assign node8714 = (inp[0]) ? 4'b1001 : 4'b0001;
															assign node8717 = (inp[10]) ? 4'b0001 : node8718;
																assign node8718 = (inp[0]) ? 4'b0001 : 4'b0101;
														assign node8722 = (inp[13]) ? 4'b0001 : node8723;
															assign node8723 = (inp[0]) ? 4'b0101 : node8724;
																assign node8724 = (inp[10]) ? 4'b0001 : 4'b0100;
													assign node8729 = (inp[13]) ? node8733 : node8730;
														assign node8730 = (inp[0]) ? 4'b0101 : 4'b0001;
														assign node8733 = (inp[10]) ? 4'b0000 : 4'b0001;
												assign node8736 = (inp[0]) ? node8750 : node8737;
													assign node8737 = (inp[13]) ? node8745 : node8738;
														assign node8738 = (inp[10]) ? node8742 : node8739;
															assign node8739 = (inp[14]) ? 4'b1001 : 4'b1000;
															assign node8742 = (inp[7]) ? 4'b0101 : 4'b1001;
														assign node8745 = (inp[14]) ? node8747 : 4'b1001;
															assign node8747 = (inp[10]) ? 4'b1000 : 4'b1001;
													assign node8750 = (inp[7]) ? node8764 : node8751;
														assign node8751 = (inp[14]) ? node8759 : node8752;
															assign node8752 = (inp[13]) ? node8756 : node8753;
																assign node8753 = (inp[10]) ? 4'b1001 : 4'b0001;
																assign node8756 = (inp[10]) ? 4'b0001 : 4'b1001;
															assign node8759 = (inp[10]) ? node8761 : 4'b0000;
																assign node8761 = (inp[13]) ? 4'b0000 : 4'b1000;
														assign node8764 = (inp[13]) ? 4'b0001 : 4'b0101;
										assign node8767 = (inp[10]) ? node8805 : node8768;
											assign node8768 = (inp[2]) ? node8780 : node8769;
												assign node8769 = (inp[12]) ? node8771 : 4'b1001;
													assign node8771 = (inp[13]) ? node8775 : node8772;
														assign node8772 = (inp[0]) ? 4'b1001 : 4'b0001;
														assign node8775 = (inp[0]) ? node8777 : 4'b1001;
															assign node8777 = (inp[7]) ? 4'b1001 : 4'b0001;
												assign node8780 = (inp[7]) ? node8792 : node8781;
													assign node8781 = (inp[0]) ? node8785 : node8782;
														assign node8782 = (inp[12]) ? 4'b0101 : 4'b0001;
														assign node8785 = (inp[13]) ? node8789 : node8786;
															assign node8786 = (inp[12]) ? 4'b0001 : 4'b1001;
															assign node8789 = (inp[14]) ? 4'b1001 : 4'b0001;
													assign node8792 = (inp[0]) ? node8800 : node8793;
														assign node8793 = (inp[12]) ? node8797 : node8794;
															assign node8794 = (inp[13]) ? 4'b0001 : 4'b0101;
															assign node8797 = (inp[13]) ? 4'b0001 : 4'b1001;
														assign node8800 = (inp[12]) ? 4'b0101 : node8801;
															assign node8801 = (inp[13]) ? 4'b0001 : 4'b0101;
											assign node8805 = (inp[13]) ? 4'b0001 : node8806;
												assign node8806 = (inp[0]) ? node8812 : node8807;
													assign node8807 = (inp[7]) ? node8809 : 4'b0001;
														assign node8809 = (inp[2]) ? 4'b0001 : 4'b1001;
													assign node8812 = (inp[7]) ? node8816 : node8813;
														assign node8813 = (inp[2]) ? 4'b1001 : 4'b0101;
														assign node8816 = (inp[2]) ? 4'b0101 : 4'b0001;
							assign node8820 = (inp[4]) ? node9236 : node8821;
								assign node8821 = (inp[1]) ? node9053 : node8822;
									assign node8822 = (inp[0]) ? node8926 : node8823;
										assign node8823 = (inp[7]) ? node8881 : node8824;
											assign node8824 = (inp[2]) ? node8850 : node8825;
												assign node8825 = (inp[13]) ? node8837 : node8826;
													assign node8826 = (inp[10]) ? node8832 : node8827;
														assign node8827 = (inp[11]) ? 4'b0001 : node8828;
															assign node8828 = (inp[14]) ? 4'b1000 : 4'b1001;
														assign node8832 = (inp[11]) ? 4'b1000 : node8833;
															assign node8833 = (inp[14]) ? 4'b1001 : 4'b0000;
													assign node8837 = (inp[10]) ? node8843 : node8838;
														assign node8838 = (inp[12]) ? node8840 : 4'b0000;
															assign node8840 = (inp[11]) ? 4'b0000 : 4'b1000;
														assign node8843 = (inp[11]) ? 4'b1000 : node8844;
															assign node8844 = (inp[12]) ? 4'b1001 : node8845;
																assign node8845 = (inp[14]) ? 4'b0001 : 4'b0000;
												assign node8850 = (inp[11]) ? node8868 : node8851;
													assign node8851 = (inp[14]) ? node8859 : node8852;
														assign node8852 = (inp[13]) ? node8856 : node8853;
															assign node8853 = (inp[10]) ? 4'b0000 : 4'b1000;
															assign node8856 = (inp[10]) ? 4'b1000 : 4'b0001;
														assign node8859 = (inp[12]) ? node8861 : 4'b1001;
															assign node8861 = (inp[13]) ? node8865 : node8862;
																assign node8862 = (inp[10]) ? 4'b0000 : 4'b0001;
																assign node8865 = (inp[10]) ? 4'b0001 : 4'b0000;
													assign node8868 = (inp[10]) ? node8874 : node8869;
														assign node8869 = (inp[12]) ? node8871 : 4'b0001;
															assign node8871 = (inp[13]) ? 4'b0001 : 4'b1000;
														assign node8874 = (inp[12]) ? node8878 : node8875;
															assign node8875 = (inp[13]) ? 4'b0001 : 4'b0000;
															assign node8878 = (inp[13]) ? 4'b0000 : 4'b0001;
											assign node8881 = (inp[10]) ? node8905 : node8882;
												assign node8882 = (inp[13]) ? node8894 : node8883;
													assign node8883 = (inp[11]) ? node8889 : node8884;
														assign node8884 = (inp[14]) ? node8886 : 4'b1000;
															assign node8886 = (inp[2]) ? 4'b0001 : 4'b1000;
														assign node8889 = (inp[12]) ? node8891 : 4'b0000;
															assign node8891 = (inp[2]) ? 4'b1000 : 4'b0000;
													assign node8894 = (inp[11]) ? node8900 : node8895;
														assign node8895 = (inp[14]) ? node8897 : 4'b0001;
															assign node8897 = (inp[12]) ? 4'b0001 : 4'b0000;
														assign node8900 = (inp[2]) ? 4'b1000 : node8901;
															assign node8901 = (inp[12]) ? 4'b0001 : 4'b1001;
												assign node8905 = (inp[2]) ? node8917 : node8906;
													assign node8906 = (inp[11]) ? node8914 : node8907;
														assign node8907 = (inp[13]) ? node8909 : 4'b1001;
															assign node8909 = (inp[12]) ? node8911 : 4'b0001;
																assign node8911 = (inp[14]) ? 4'b0000 : 4'b0001;
														assign node8914 = (inp[13]) ? 4'b1001 : 4'b0001;
													assign node8917 = (inp[11]) ? node8921 : node8918;
														assign node8918 = (inp[13]) ? 4'b1001 : 4'b0000;
														assign node8921 = (inp[13]) ? 4'b0000 : node8922;
															assign node8922 = (inp[12]) ? 4'b0001 : 4'b1001;
										assign node8926 = (inp[11]) ? node9006 : node8927;
											assign node8927 = (inp[2]) ? node8963 : node8928;
												assign node8928 = (inp[12]) ? node8946 : node8929;
													assign node8929 = (inp[10]) ? node8937 : node8930;
														assign node8930 = (inp[7]) ? 4'b1001 : node8931;
															assign node8931 = (inp[13]) ? 4'b0000 : node8932;
																assign node8932 = (inp[14]) ? 4'b1000 : 4'b1001;
														assign node8937 = (inp[14]) ? node8941 : node8938;
															assign node8938 = (inp[7]) ? 4'b1000 : 4'b0000;
															assign node8941 = (inp[13]) ? node8943 : 4'b0000;
																assign node8943 = (inp[7]) ? 4'b0001 : 4'b0000;
													assign node8946 = (inp[14]) ? node8954 : node8947;
														assign node8947 = (inp[13]) ? node8949 : 4'b0001;
															assign node8949 = (inp[7]) ? node8951 : 4'b0000;
																assign node8951 = (inp[10]) ? 4'b0000 : 4'b0001;
														assign node8954 = (inp[13]) ? node8960 : node8955;
															assign node8955 = (inp[7]) ? 4'b0000 : node8956;
																assign node8956 = (inp[10]) ? 4'b0001 : 4'b0000;
															assign node8960 = (inp[10]) ? 4'b0000 : 4'b0001;
												assign node8963 = (inp[14]) ? node8989 : node8964;
													assign node8964 = (inp[13]) ? node8978 : node8965;
														assign node8965 = (inp[7]) ? node8973 : node8966;
															assign node8966 = (inp[10]) ? node8970 : node8967;
																assign node8967 = (inp[12]) ? 4'b0000 : 4'b1000;
																assign node8970 = (inp[12]) ? 4'b1000 : 4'b0000;
															assign node8973 = (inp[12]) ? node8975 : 4'b1000;
																assign node8975 = (inp[10]) ? 4'b1000 : 4'b0000;
														assign node8978 = (inp[12]) ? node8984 : node8979;
															assign node8979 = (inp[7]) ? 4'b0000 : node8980;
																assign node8980 = (inp[10]) ? 4'b0000 : 4'b1000;
															assign node8984 = (inp[10]) ? 4'b1000 : node8985;
																assign node8985 = (inp[7]) ? 4'b1000 : 4'b0000;
													assign node8989 = (inp[13]) ? node8999 : node8990;
														assign node8990 = (inp[7]) ? node8994 : node8991;
															assign node8991 = (inp[12]) ? 4'b0001 : 4'b0000;
															assign node8994 = (inp[10]) ? node8996 : 4'b0001;
																assign node8996 = (inp[12]) ? 4'b0001 : 4'b1001;
														assign node8999 = (inp[7]) ? node9001 : 4'b1000;
															assign node9001 = (inp[10]) ? node9003 : 4'b1001;
																assign node9003 = (inp[12]) ? 4'b1001 : 4'b0000;
											assign node9006 = (inp[13]) ? node9022 : node9007;
												assign node9007 = (inp[2]) ? node9013 : node9008;
													assign node9008 = (inp[10]) ? node9010 : 4'b1000;
														assign node9010 = (inp[7]) ? 4'b1000 : 4'b1001;
													assign node9013 = (inp[10]) ? node9017 : node9014;
														assign node9014 = (inp[12]) ? 4'b0000 : 4'b1000;
														assign node9017 = (inp[12]) ? 4'b1000 : node9018;
															assign node9018 = (inp[7]) ? 4'b1000 : 4'b0001;
												assign node9022 = (inp[2]) ? node9038 : node9023;
													assign node9023 = (inp[12]) ? node9031 : node9024;
														assign node9024 = (inp[7]) ? node9028 : node9025;
															assign node9025 = (inp[10]) ? 4'b1001 : 4'b1000;
															assign node9028 = (inp[10]) ? 4'b1000 : 4'b1001;
														assign node9031 = (inp[7]) ? node9035 : node9032;
															assign node9032 = (inp[10]) ? 4'b0001 : 4'b0000;
															assign node9035 = (inp[10]) ? 4'b1000 : 4'b1001;
													assign node9038 = (inp[7]) ? node9046 : node9039;
														assign node9039 = (inp[12]) ? node9043 : node9040;
															assign node9040 = (inp[10]) ? 4'b0000 : 4'b1001;
															assign node9043 = (inp[10]) ? 4'b1001 : 4'b0001;
														assign node9046 = (inp[10]) ? node9050 : node9047;
															assign node9047 = (inp[12]) ? 4'b1000 : 4'b0000;
															assign node9050 = (inp[12]) ? 4'b0000 : 4'b0001;
									assign node9053 = (inp[11]) ? node9175 : node9054;
										assign node9054 = (inp[10]) ? node9126 : node9055;
											assign node9055 = (inp[7]) ? node9093 : node9056;
												assign node9056 = (inp[2]) ? node9074 : node9057;
													assign node9057 = (inp[12]) ? node9065 : node9058;
														assign node9058 = (inp[0]) ? 4'b0001 : node9059;
															assign node9059 = (inp[13]) ? node9061 : 4'b1001;
																assign node9061 = (inp[14]) ? 4'b1001 : 4'b0000;
														assign node9065 = (inp[0]) ? node9067 : 4'b1001;
															assign node9067 = (inp[13]) ? node9071 : node9068;
																assign node9068 = (inp[14]) ? 4'b1001 : 4'b1000;
																assign node9071 = (inp[14]) ? 4'b1000 : 4'b1001;
													assign node9074 = (inp[12]) ? node9086 : node9075;
														assign node9075 = (inp[14]) ? node9081 : node9076;
															assign node9076 = (inp[13]) ? 4'b1000 : node9077;
																assign node9077 = (inp[0]) ? 4'b1001 : 4'b1000;
															assign node9081 = (inp[13]) ? node9083 : 4'b1000;
																assign node9083 = (inp[0]) ? 4'b1000 : 4'b1001;
														assign node9086 = (inp[13]) ? node9090 : node9087;
															assign node9087 = (inp[0]) ? 4'b0001 : 4'b0000;
															assign node9090 = (inp[0]) ? 4'b1000 : 4'b1001;
												assign node9093 = (inp[0]) ? node9111 : node9094;
													assign node9094 = (inp[13]) ? node9104 : node9095;
														assign node9095 = (inp[2]) ? node9101 : node9096;
															assign node9096 = (inp[14]) ? node9098 : 4'b1000;
																assign node9098 = (inp[12]) ? 4'b0001 : 4'b1001;
															assign node9101 = (inp[14]) ? 4'b0000 : 4'b0001;
														assign node9104 = (inp[14]) ? node9106 : 4'b0000;
															assign node9106 = (inp[2]) ? node9108 : 4'b0000;
																assign node9108 = (inp[12]) ? 4'b1001 : 4'b0001;
													assign node9111 = (inp[13]) ? node9123 : node9112;
														assign node9112 = (inp[12]) ? node9120 : node9113;
															assign node9113 = (inp[14]) ? node9117 : node9114;
																assign node9114 = (inp[2]) ? 4'b1001 : 4'b0000;
																assign node9117 = (inp[2]) ? 4'b1000 : 4'b1001;
															assign node9120 = (inp[2]) ? 4'b0000 : 4'b1000;
														assign node9123 = (inp[12]) ? 4'b1001 : 4'b0001;
											assign node9126 = (inp[13]) ? node9146 : node9127;
												assign node9127 = (inp[2]) ? node9133 : node9128;
													assign node9128 = (inp[14]) ? node9130 : 4'b0001;
														assign node9130 = (inp[0]) ? 4'b0001 : 4'b0000;
													assign node9133 = (inp[7]) ? node9143 : node9134;
														assign node9134 = (inp[12]) ? node9138 : node9135;
															assign node9135 = (inp[14]) ? 4'b0000 : 4'b1000;
															assign node9138 = (inp[0]) ? 4'b0000 : node9139;
																assign node9139 = (inp[14]) ? 4'b0001 : 4'b0000;
														assign node9143 = (inp[0]) ? 4'b1000 : 4'b0000;
												assign node9146 = (inp[0]) ? node9162 : node9147;
													assign node9147 = (inp[12]) ? node9153 : node9148;
														assign node9148 = (inp[14]) ? 4'b1000 : node9149;
															assign node9149 = (inp[2]) ? 4'b1000 : 4'b1001;
														assign node9153 = (inp[2]) ? node9159 : node9154;
															assign node9154 = (inp[14]) ? 4'b0000 : node9155;
																assign node9155 = (inp[7]) ? 4'b0001 : 4'b0000;
															assign node9159 = (inp[7]) ? 4'b1001 : 4'b1000;
													assign node9162 = (inp[2]) ? node9170 : node9163;
														assign node9163 = (inp[12]) ? node9165 : 4'b0000;
															assign node9165 = (inp[7]) ? node9167 : 4'b1000;
																assign node9167 = (inp[14]) ? 4'b1000 : 4'b1001;
														assign node9170 = (inp[7]) ? 4'b0000 : node9171;
															assign node9171 = (inp[14]) ? 4'b0001 : 4'b0000;
										assign node9175 = (inp[13]) ? node9215 : node9176;
											assign node9176 = (inp[2]) ? node9188 : node9177;
												assign node9177 = (inp[7]) ? node9179 : 4'b0001;
													assign node9179 = (inp[0]) ? node9183 : node9180;
														assign node9180 = (inp[10]) ? 4'b1001 : 4'b0001;
														assign node9183 = (inp[10]) ? 4'b0001 : node9184;
															assign node9184 = (inp[14]) ? 4'b1001 : 4'b0001;
												assign node9188 = (inp[12]) ? node9202 : node9189;
													assign node9189 = (inp[10]) ? node9191 : 4'b1001;
														assign node9191 = (inp[14]) ? node9197 : node9192;
															assign node9192 = (inp[7]) ? node9194 : 4'b0001;
																assign node9194 = (inp[0]) ? 4'b1001 : 4'b0001;
															assign node9197 = (inp[0]) ? node9199 : 4'b1001;
																assign node9199 = (inp[7]) ? 4'b1001 : 4'b0001;
													assign node9202 = (inp[10]) ? node9208 : node9203;
														assign node9203 = (inp[0]) ? 4'b0001 : node9204;
															assign node9204 = (inp[7]) ? 4'b0001 : 4'b1001;
														assign node9208 = (inp[7]) ? node9212 : node9209;
															assign node9209 = (inp[0]) ? 4'b0001 : 4'b1001;
															assign node9212 = (inp[0]) ? 4'b1001 : 4'b0001;
											assign node9215 = (inp[10]) ? 4'b0001 : node9216;
												assign node9216 = (inp[0]) ? node9224 : node9217;
													assign node9217 = (inp[12]) ? 4'b0001 : node9218;
														assign node9218 = (inp[2]) ? 4'b0001 : node9219;
															assign node9219 = (inp[7]) ? 4'b1001 : 4'b0001;
													assign node9224 = (inp[2]) ? node9230 : node9225;
														assign node9225 = (inp[7]) ? 4'b0001 : node9226;
															assign node9226 = (inp[12]) ? 4'b1001 : 4'b0001;
														assign node9230 = (inp[12]) ? 4'b1001 : node9231;
															assign node9231 = (inp[7]) ? 4'b0001 : 4'b1001;
								assign node9236 = (inp[13]) ? node9442 : node9237;
									assign node9237 = (inp[1]) ? node9359 : node9238;
										assign node9238 = (inp[0]) ? node9294 : node9239;
											assign node9239 = (inp[2]) ? node9269 : node9240;
												assign node9240 = (inp[7]) ? node9260 : node9241;
													assign node9241 = (inp[14]) ? node9253 : node9242;
														assign node9242 = (inp[12]) ? node9248 : node9243;
															assign node9243 = (inp[10]) ? node9245 : 4'b1000;
																assign node9245 = (inp[11]) ? 4'b0001 : 4'b0000;
															assign node9248 = (inp[10]) ? 4'b0000 : node9249;
																assign node9249 = (inp[11]) ? 4'b0000 : 4'b0001;
														assign node9253 = (inp[11]) ? node9257 : node9254;
															assign node9254 = (inp[10]) ? 4'b0000 : 4'b0001;
															assign node9257 = (inp[10]) ? 4'b0001 : 4'b0000;
													assign node9260 = (inp[11]) ? 4'b0001 : node9261;
														assign node9261 = (inp[14]) ? 4'b0000 : node9262;
															assign node9262 = (inp[10]) ? node9264 : 4'b0001;
																assign node9264 = (inp[12]) ? 4'b0001 : 4'b0000;
												assign node9269 = (inp[12]) ? node9283 : node9270;
													assign node9270 = (inp[10]) ? node9276 : node9271;
														assign node9271 = (inp[7]) ? 4'b1000 : node9272;
															assign node9272 = (inp[11]) ? 4'b0000 : 4'b0001;
														assign node9276 = (inp[7]) ? node9278 : 4'b0001;
															assign node9278 = (inp[11]) ? 4'b0001 : node9279;
																assign node9279 = (inp[14]) ? 4'b0000 : 4'b0001;
													assign node9283 = (inp[11]) ? node9289 : node9284;
														assign node9284 = (inp[7]) ? 4'b1000 : node9285;
															assign node9285 = (inp[10]) ? 4'b0001 : 4'b1000;
														assign node9289 = (inp[7]) ? 4'b0001 : node9290;
															assign node9290 = (inp[10]) ? 4'b1000 : 4'b1001;
											assign node9294 = (inp[12]) ? node9328 : node9295;
												assign node9295 = (inp[10]) ? node9311 : node9296;
													assign node9296 = (inp[2]) ? node9304 : node9297;
														assign node9297 = (inp[11]) ? node9301 : node9298;
															assign node9298 = (inp[7]) ? 4'b1000 : 4'b1001;
															assign node9301 = (inp[14]) ? 4'b0000 : 4'b0001;
														assign node9304 = (inp[7]) ? 4'b1001 : node9305;
															assign node9305 = (inp[14]) ? 4'b1000 : node9306;
																assign node9306 = (inp[11]) ? 4'b1000 : 4'b1001;
													assign node9311 = (inp[7]) ? node9319 : node9312;
														assign node9312 = (inp[2]) ? node9314 : 4'b1000;
															assign node9314 = (inp[11]) ? 4'b0000 : node9315;
																assign node9315 = (inp[14]) ? 4'b1001 : 4'b0000;
														assign node9319 = (inp[2]) ? node9323 : node9320;
															assign node9320 = (inp[11]) ? 4'b0001 : 4'b0000;
															assign node9323 = (inp[11]) ? 4'b1000 : node9324;
																assign node9324 = (inp[14]) ? 4'b0000 : 4'b0001;
												assign node9328 = (inp[2]) ? node9344 : node9329;
													assign node9329 = (inp[7]) ? node9337 : node9330;
														assign node9330 = (inp[10]) ? 4'b0000 : node9331;
															assign node9331 = (inp[11]) ? 4'b0001 : node9332;
																assign node9332 = (inp[14]) ? 4'b1000 : 4'b1001;
														assign node9337 = (inp[10]) ? node9341 : node9338;
															assign node9338 = (inp[11]) ? 4'b0000 : 4'b1000;
															assign node9341 = (inp[11]) ? 4'b1000 : 4'b1001;
													assign node9344 = (inp[10]) ? node9352 : node9345;
														assign node9345 = (inp[7]) ? node9349 : node9346;
															assign node9346 = (inp[11]) ? 4'b1000 : 4'b0000;
															assign node9349 = (inp[11]) ? 4'b0001 : 4'b0000;
														assign node9352 = (inp[11]) ? 4'b0000 : node9353;
															assign node9353 = (inp[7]) ? node9355 : 4'b0001;
																assign node9355 = (inp[14]) ? 4'b0000 : 4'b0001;
										assign node9359 = (inp[11]) ? node9421 : node9360;
											assign node9360 = (inp[10]) ? node9390 : node9361;
												assign node9361 = (inp[12]) ? node9377 : node9362;
													assign node9362 = (inp[7]) ? node9368 : node9363;
														assign node9363 = (inp[0]) ? node9365 : 4'b0000;
															assign node9365 = (inp[14]) ? 4'b0000 : 4'b0001;
														assign node9368 = (inp[0]) ? node9372 : node9369;
															assign node9369 = (inp[14]) ? 4'b1000 : 4'b1001;
															assign node9372 = (inp[14]) ? 4'b1000 : node9373;
																assign node9373 = (inp[2]) ? 4'b0000 : 4'b1000;
													assign node9377 = (inp[7]) ? node9381 : node9378;
														assign node9378 = (inp[0]) ? 4'b1001 : 4'b1000;
														assign node9381 = (inp[0]) ? node9387 : node9382;
															assign node9382 = (inp[2]) ? 4'b0001 : node9383;
																assign node9383 = (inp[14]) ? 4'b0000 : 4'b0001;
															assign node9387 = (inp[14]) ? 4'b0001 : 4'b1000;
												assign node9390 = (inp[12]) ? node9406 : node9391;
													assign node9391 = (inp[7]) ? node9401 : node9392;
														assign node9392 = (inp[0]) ? node9398 : node9393;
															assign node9393 = (inp[14]) ? 4'b0001 : node9394;
																assign node9394 = (inp[2]) ? 4'b0001 : 4'b0000;
															assign node9398 = (inp[2]) ? 4'b0000 : 4'b0001;
														assign node9401 = (inp[0]) ? node9403 : 4'b0000;
															assign node9403 = (inp[14]) ? 4'b0001 : 4'b0000;
													assign node9406 = (inp[14]) ? node9412 : node9407;
														assign node9407 = (inp[0]) ? 4'b1000 : node9408;
															assign node9408 = (inp[7]) ? 4'b0001 : 4'b0000;
														assign node9412 = (inp[2]) ? node9416 : node9413;
															assign node9413 = (inp[0]) ? 4'b0001 : 4'b1000;
															assign node9416 = (inp[0]) ? node9418 : 4'b0001;
																assign node9418 = (inp[7]) ? 4'b0001 : 4'b0000;
											assign node9421 = (inp[10]) ? 4'b0001 : node9422;
												assign node9422 = (inp[12]) ? node9434 : node9423;
													assign node9423 = (inp[2]) ? node9429 : node9424;
														assign node9424 = (inp[7]) ? 4'b0001 : node9425;
															assign node9425 = (inp[0]) ? 4'b1001 : 4'b0001;
														assign node9429 = (inp[0]) ? 4'b0001 : node9430;
															assign node9430 = (inp[7]) ? 4'b1001 : 4'b0001;
													assign node9434 = (inp[0]) ? node9436 : 4'b1001;
														assign node9436 = (inp[7]) ? node9438 : 4'b0001;
															assign node9438 = (inp[2]) ? 4'b1001 : 4'b0001;
									assign node9442 = (inp[10]) ? node9536 : node9443;
										assign node9443 = (inp[1]) ? node9503 : node9444;
											assign node9444 = (inp[14]) ? node9466 : node9445;
												assign node9445 = (inp[11]) ? node9455 : node9446;
													assign node9446 = (inp[0]) ? node9450 : node9447;
														assign node9447 = (inp[7]) ? 4'b0001 : 4'b0000;
														assign node9450 = (inp[7]) ? 4'b0000 : node9451;
															assign node9451 = (inp[12]) ? 4'b0001 : 4'b0000;
													assign node9455 = (inp[12]) ? 4'b0000 : node9456;
														assign node9456 = (inp[7]) ? node9458 : 4'b0000;
															assign node9458 = (inp[2]) ? node9462 : node9459;
																assign node9459 = (inp[0]) ? 4'b0000 : 4'b0001;
																assign node9462 = (inp[0]) ? 4'b0001 : 4'b0000;
												assign node9466 = (inp[2]) ? node9488 : node9467;
													assign node9467 = (inp[0]) ? node9477 : node9468;
														assign node9468 = (inp[12]) ? node9470 : 4'b0001;
															assign node9470 = (inp[11]) ? node9474 : node9471;
																assign node9471 = (inp[7]) ? 4'b0001 : 4'b0000;
																assign node9474 = (inp[7]) ? 4'b0000 : 4'b0001;
														assign node9477 = (inp[12]) ? node9483 : node9478;
															assign node9478 = (inp[11]) ? 4'b0000 : node9479;
																assign node9479 = (inp[7]) ? 4'b0000 : 4'b0001;
															assign node9483 = (inp[11]) ? 4'b0001 : node9484;
																assign node9484 = (inp[7]) ? 4'b0000 : 4'b0001;
													assign node9488 = (inp[0]) ? node9494 : node9489;
														assign node9489 = (inp[7]) ? 4'b0000 : node9490;
															assign node9490 = (inp[12]) ? 4'b0001 : 4'b0000;
														assign node9494 = (inp[7]) ? node9500 : node9495;
															assign node9495 = (inp[11]) ? node9497 : 4'b0000;
																assign node9497 = (inp[12]) ? 4'b0001 : 4'b0000;
															assign node9500 = (inp[12]) ? 4'b0000 : 4'b0001;
											assign node9503 = (inp[11]) ? 4'b0001 : node9504;
												assign node9504 = (inp[7]) ? node9520 : node9505;
													assign node9505 = (inp[0]) ? node9515 : node9506;
														assign node9506 = (inp[14]) ? node9510 : node9507;
															assign node9507 = (inp[12]) ? 4'b0000 : 4'b0001;
															assign node9510 = (inp[12]) ? 4'b0001 : node9511;
																assign node9511 = (inp[2]) ? 4'b0001 : 4'b0000;
														assign node9515 = (inp[12]) ? 4'b0000 : node9516;
															assign node9516 = (inp[14]) ? 4'b0001 : 4'b0000;
													assign node9520 = (inp[2]) ? node9528 : node9521;
														assign node9521 = (inp[0]) ? 4'b0001 : node9522;
															assign node9522 = (inp[14]) ? 4'b0000 : node9523;
																assign node9523 = (inp[12]) ? 4'b0001 : 4'b0000;
														assign node9528 = (inp[0]) ? node9530 : 4'b0001;
															assign node9530 = (inp[12]) ? 4'b0000 : node9531;
																assign node9531 = (inp[14]) ? 4'b0001 : 4'b0000;
										assign node9536 = (inp[11]) ? 4'b0000 : node9537;
											assign node9537 = (inp[1]) ? 4'b0000 : node9538;
												assign node9538 = (inp[2]) ? node9550 : node9539;
													assign node9539 = (inp[14]) ? node9541 : 4'b0000;
														assign node9541 = (inp[0]) ? node9547 : node9542;
															assign node9542 = (inp[12]) ? node9544 : 4'b0001;
																assign node9544 = (inp[7]) ? 4'b0000 : 4'b0001;
															assign node9547 = (inp[7]) ? 4'b0001 : 4'b0000;
													assign node9550 = (inp[7]) ? node9558 : node9551;
														assign node9551 = (inp[0]) ? 4'b0001 : node9552;
															assign node9552 = (inp[12]) ? node9554 : 4'b0001;
																assign node9554 = (inp[14]) ? 4'b0000 : 4'b0001;
														assign node9558 = (inp[12]) ? 4'b0000 : node9559;
															assign node9559 = (inp[0]) ? 4'b0001 : node9560;
																assign node9560 = (inp[14]) ? 4'b0000 : 4'b0001;
				assign node9567 = (inp[0]) ? node11745 : node9568;
					assign node9568 = (inp[6]) ? node10144 : node9569;
						assign node9569 = (inp[2]) ? node10029 : node9570;
							assign node9570 = (inp[5]) ? node9674 : node9571;
								assign node9571 = (inp[3]) ? node9573 : 4'b0011;
									assign node9573 = (inp[7]) ? node9647 : node9574;
										assign node9574 = (inp[4]) ? node9602 : node9575;
											assign node9575 = (inp[13]) ? node9577 : 4'b0011;
												assign node9577 = (inp[12]) ? node9591 : node9578;
													assign node9578 = (inp[1]) ? node9586 : node9579;
														assign node9579 = (inp[14]) ? node9581 : 4'b0000;
															assign node9581 = (inp[11]) ? 4'b0000 : node9582;
																assign node9582 = (inp[10]) ? 4'b0001 : 4'b0011;
														assign node9586 = (inp[11]) ? 4'b0001 : node9587;
															assign node9587 = (inp[14]) ? 4'b0000 : 4'b0001;
													assign node9591 = (inp[10]) ? node9593 : 4'b0011;
														assign node9593 = (inp[11]) ? node9599 : node9594;
															assign node9594 = (inp[1]) ? node9596 : 4'b0011;
																assign node9596 = (inp[14]) ? 4'b0000 : 4'b0001;
															assign node9599 = (inp[1]) ? 4'b0001 : 4'b0000;
											assign node9602 = (inp[1]) ? node9628 : node9603;
												assign node9603 = (inp[11]) ? node9621 : node9604;
													assign node9604 = (inp[14]) ? node9614 : node9605;
														assign node9605 = (inp[10]) ? node9611 : node9606;
															assign node9606 = (inp[13]) ? node9608 : 4'b0000;
																assign node9608 = (inp[12]) ? 4'b1000 : 4'b0000;
															assign node9611 = (inp[13]) ? 4'b0000 : 4'b1000;
														assign node9614 = (inp[13]) ? node9616 : 4'b0001;
															assign node9616 = (inp[10]) ? node9618 : 4'b1001;
																assign node9618 = (inp[12]) ? 4'b1001 : 4'b0001;
													assign node9621 = (inp[13]) ? 4'b0000 : node9622;
														assign node9622 = (inp[10]) ? 4'b1000 : node9623;
															assign node9623 = (inp[12]) ? 4'b0000 : 4'b1000;
												assign node9628 = (inp[13]) ? node9638 : node9629;
													assign node9629 = (inp[14]) ? node9635 : node9630;
														assign node9630 = (inp[10]) ? 4'b1001 : node9631;
															assign node9631 = (inp[12]) ? 4'b0001 : 4'b1001;
														assign node9635 = (inp[11]) ? 4'b1001 : 4'b1000;
													assign node9638 = (inp[14]) ? node9644 : node9639;
														assign node9639 = (inp[12]) ? node9641 : 4'b0001;
															assign node9641 = (inp[10]) ? 4'b0001 : 4'b1001;
														assign node9644 = (inp[11]) ? 4'b1001 : 4'b0000;
										assign node9647 = (inp[13]) ? node9649 : 4'b0011;
											assign node9649 = (inp[4]) ? node9651 : 4'b0011;
												assign node9651 = (inp[12]) ? node9665 : node9652;
													assign node9652 = (inp[1]) ? node9660 : node9653;
														assign node9653 = (inp[14]) ? node9655 : 4'b0000;
															assign node9655 = (inp[11]) ? 4'b0000 : node9656;
																assign node9656 = (inp[10]) ? 4'b0001 : 4'b0011;
														assign node9660 = (inp[14]) ? node9662 : 4'b0001;
															assign node9662 = (inp[11]) ? 4'b0001 : 4'b0000;
													assign node9665 = (inp[10]) ? node9667 : 4'b0011;
														assign node9667 = (inp[1]) ? node9669 : 4'b0011;
															assign node9669 = (inp[14]) ? node9671 : 4'b0001;
																assign node9671 = (inp[11]) ? 4'b0001 : 4'b0000;
								assign node9674 = (inp[1]) ? node9852 : node9675;
									assign node9675 = (inp[11]) ? node9793 : node9676;
										assign node9676 = (inp[14]) ? node9732 : node9677;
											assign node9677 = (inp[13]) ? node9703 : node9678;
												assign node9678 = (inp[12]) ? node9690 : node9679;
													assign node9679 = (inp[3]) ? node9685 : node9680;
														assign node9680 = (inp[7]) ? 4'b1000 : node9681;
															assign node9681 = (inp[4]) ? 4'b1100 : 4'b1000;
														assign node9685 = (inp[4]) ? node9687 : 4'b1100;
															assign node9687 = (inp[7]) ? 4'b1100 : 4'b1000;
													assign node9690 = (inp[10]) ? node9698 : node9691;
														assign node9691 = (inp[3]) ? 4'b0100 : node9692;
															assign node9692 = (inp[4]) ? node9694 : 4'b0000;
																assign node9694 = (inp[7]) ? 4'b0000 : 4'b0100;
														assign node9698 = (inp[3]) ? node9700 : 4'b1000;
															assign node9700 = (inp[7]) ? 4'b1100 : 4'b1000;
												assign node9703 = (inp[10]) ? node9721 : node9704;
													assign node9704 = (inp[12]) ? node9714 : node9705;
														assign node9705 = (inp[4]) ? node9711 : node9706;
															assign node9706 = (inp[7]) ? node9708 : 4'b0000;
																assign node9708 = (inp[3]) ? 4'b0100 : 4'b0000;
															assign node9711 = (inp[3]) ? 4'b0000 : 4'b0100;
														assign node9714 = (inp[7]) ? 4'b1000 : node9715;
															assign node9715 = (inp[3]) ? 4'b1100 : node9716;
																assign node9716 = (inp[4]) ? 4'b1100 : 4'b1000;
													assign node9721 = (inp[3]) ? node9727 : node9722;
														assign node9722 = (inp[4]) ? 4'b0100 : node9723;
															assign node9723 = (inp[7]) ? 4'b0000 : 4'b0100;
														assign node9727 = (inp[7]) ? node9729 : 4'b0000;
															assign node9729 = (inp[4]) ? 4'b0000 : 4'b0100;
											assign node9732 = (inp[13]) ? node9764 : node9733;
												assign node9733 = (inp[3]) ? node9751 : node9734;
													assign node9734 = (inp[4]) ? node9740 : node9735;
														assign node9735 = (inp[12]) ? 4'b0001 : node9736;
															assign node9736 = (inp[10]) ? 4'b1001 : 4'b0001;
														assign node9740 = (inp[7]) ? node9746 : node9741;
															assign node9741 = (inp[10]) ? node9743 : 4'b0101;
																assign node9743 = (inp[12]) ? 4'b0101 : 4'b1101;
															assign node9746 = (inp[12]) ? 4'b0001 : node9747;
																assign node9747 = (inp[10]) ? 4'b1001 : 4'b0001;
													assign node9751 = (inp[10]) ? node9757 : node9752;
														assign node9752 = (inp[7]) ? 4'b0101 : node9753;
															assign node9753 = (inp[4]) ? 4'b0001 : 4'b0101;
														assign node9757 = (inp[12]) ? 4'b0101 : node9758;
															assign node9758 = (inp[4]) ? node9760 : 4'b1101;
																assign node9760 = (inp[7]) ? 4'b1101 : 4'b1001;
												assign node9764 = (inp[12]) ? node9782 : node9765;
													assign node9765 = (inp[10]) ? node9775 : node9766;
														assign node9766 = (inp[3]) ? node9770 : node9767;
															assign node9767 = (inp[4]) ? 4'b1101 : 4'b1001;
															assign node9770 = (inp[4]) ? node9772 : 4'b1101;
																assign node9772 = (inp[7]) ? 4'b1101 : 4'b1001;
														assign node9775 = (inp[3]) ? node9777 : 4'b0101;
															assign node9777 = (inp[7]) ? node9779 : 4'b0001;
																assign node9779 = (inp[4]) ? 4'b0001 : 4'b0101;
													assign node9782 = (inp[3]) ? node9788 : node9783;
														assign node9783 = (inp[4]) ? node9785 : 4'b1001;
															assign node9785 = (inp[7]) ? 4'b1001 : 4'b1101;
														assign node9788 = (inp[7]) ? 4'b1101 : node9789;
															assign node9789 = (inp[4]) ? 4'b1001 : 4'b1101;
										assign node9793 = (inp[13]) ? node9817 : node9794;
											assign node9794 = (inp[3]) ? node9808 : node9795;
												assign node9795 = (inp[10]) ? node9803 : node9796;
													assign node9796 = (inp[12]) ? node9798 : 4'b1000;
														assign node9798 = (inp[7]) ? 4'b0000 : node9799;
															assign node9799 = (inp[4]) ? 4'b0100 : 4'b0000;
													assign node9803 = (inp[7]) ? 4'b1000 : node9804;
														assign node9804 = (inp[4]) ? 4'b1100 : 4'b1000;
												assign node9808 = (inp[12]) ? node9814 : node9809;
													assign node9809 = (inp[7]) ? 4'b1100 : node9810;
														assign node9810 = (inp[4]) ? 4'b1000 : 4'b1100;
													assign node9814 = (inp[10]) ? 4'b1100 : 4'b0100;
											assign node9817 = (inp[10]) ? node9841 : node9818;
												assign node9818 = (inp[12]) ? node9830 : node9819;
													assign node9819 = (inp[3]) ? node9825 : node9820;
														assign node9820 = (inp[4]) ? 4'b0100 : node9821;
															assign node9821 = (inp[7]) ? 4'b0000 : 4'b0100;
														assign node9825 = (inp[7]) ? node9827 : 4'b0000;
															assign node9827 = (inp[4]) ? 4'b0000 : 4'b0100;
													assign node9830 = (inp[3]) ? node9836 : node9831;
														assign node9831 = (inp[7]) ? 4'b1000 : node9832;
															assign node9832 = (inp[4]) ? 4'b1100 : 4'b1000;
														assign node9836 = (inp[4]) ? node9838 : 4'b1100;
															assign node9838 = (inp[7]) ? 4'b1100 : 4'b1000;
												assign node9841 = (inp[3]) ? node9847 : node9842;
													assign node9842 = (inp[7]) ? node9844 : 4'b0100;
														assign node9844 = (inp[4]) ? 4'b0100 : 4'b0000;
													assign node9847 = (inp[7]) ? node9849 : 4'b0000;
														assign node9849 = (inp[4]) ? 4'b0000 : 4'b0100;
									assign node9852 = (inp[11]) ? node9960 : node9853;
										assign node9853 = (inp[14]) ? node9905 : node9854;
											assign node9854 = (inp[13]) ? node9880 : node9855;
												assign node9855 = (inp[10]) ? node9869 : node9856;
													assign node9856 = (inp[12]) ? node9860 : node9857;
														assign node9857 = (inp[4]) ? 4'b1101 : 4'b1001;
														assign node9860 = (inp[3]) ? node9864 : node9861;
															assign node9861 = (inp[4]) ? 4'b0101 : 4'b0001;
															assign node9864 = (inp[7]) ? 4'b0101 : node9865;
																assign node9865 = (inp[4]) ? 4'b0001 : 4'b0101;
													assign node9869 = (inp[3]) ? node9875 : node9870;
														assign node9870 = (inp[7]) ? 4'b1001 : node9871;
															assign node9871 = (inp[4]) ? 4'b1101 : 4'b1001;
														assign node9875 = (inp[4]) ? node9877 : 4'b1101;
															assign node9877 = (inp[7]) ? 4'b1101 : 4'b1001;
												assign node9880 = (inp[12]) ? node9890 : node9881;
													assign node9881 = (inp[3]) ? node9887 : node9882;
														assign node9882 = (inp[4]) ? 4'b0101 : node9883;
															assign node9883 = (inp[7]) ? 4'b0001 : 4'b0101;
														assign node9887 = (inp[4]) ? 4'b0001 : 4'b0101;
													assign node9890 = (inp[10]) ? node9898 : node9891;
														assign node9891 = (inp[3]) ? 4'b1101 : node9892;
															assign node9892 = (inp[7]) ? 4'b1001 : node9893;
																assign node9893 = (inp[4]) ? 4'b1101 : 4'b1001;
														assign node9898 = (inp[3]) ? 4'b0001 : node9899;
															assign node9899 = (inp[4]) ? 4'b0101 : node9900;
																assign node9900 = (inp[7]) ? 4'b0001 : 4'b0101;
											assign node9905 = (inp[13]) ? node9931 : node9906;
												assign node9906 = (inp[3]) ? node9916 : node9907;
													assign node9907 = (inp[12]) ? node9913 : node9908;
														assign node9908 = (inp[4]) ? node9910 : 4'b1000;
															assign node9910 = (inp[7]) ? 4'b1000 : 4'b1100;
														assign node9913 = (inp[10]) ? 4'b1000 : 4'b0000;
													assign node9916 = (inp[7]) ? node9926 : node9917;
														assign node9917 = (inp[4]) ? node9921 : node9918;
															assign node9918 = (inp[10]) ? 4'b1100 : 4'b0100;
															assign node9921 = (inp[10]) ? 4'b1000 : node9922;
																assign node9922 = (inp[12]) ? 4'b0000 : 4'b1000;
														assign node9926 = (inp[12]) ? node9928 : 4'b1100;
															assign node9928 = (inp[10]) ? 4'b1100 : 4'b0100;
												assign node9931 = (inp[10]) ? node9949 : node9932;
													assign node9932 = (inp[12]) ? node9940 : node9933;
														assign node9933 = (inp[3]) ? node9937 : node9934;
															assign node9934 = (inp[7]) ? 4'b0000 : 4'b0100;
															assign node9937 = (inp[4]) ? 4'b0000 : 4'b0100;
														assign node9940 = (inp[4]) ? node9942 : 4'b1100;
															assign node9942 = (inp[7]) ? node9946 : node9943;
																assign node9943 = (inp[3]) ? 4'b1000 : 4'b1100;
																assign node9946 = (inp[3]) ? 4'b1100 : 4'b1000;
													assign node9949 = (inp[3]) ? node9955 : node9950;
														assign node9950 = (inp[7]) ? node9952 : 4'b0100;
															assign node9952 = (inp[4]) ? 4'b0100 : 4'b0000;
														assign node9955 = (inp[7]) ? node9957 : 4'b0000;
															assign node9957 = (inp[4]) ? 4'b0000 : 4'b0100;
										assign node9960 = (inp[13]) ? node9994 : node9961;
											assign node9961 = (inp[3]) ? node9977 : node9962;
												assign node9962 = (inp[10]) ? node9972 : node9963;
													assign node9963 = (inp[12]) ? node9967 : node9964;
														assign node9964 = (inp[7]) ? 4'b1001 : 4'b1101;
														assign node9967 = (inp[14]) ? node9969 : 4'b0001;
															assign node9969 = (inp[4]) ? 4'b0101 : 4'b0001;
													assign node9972 = (inp[4]) ? node9974 : 4'b1001;
														assign node9974 = (inp[7]) ? 4'b1001 : 4'b1101;
												assign node9977 = (inp[12]) ? node9983 : node9978;
													assign node9978 = (inp[7]) ? 4'b1101 : node9979;
														assign node9979 = (inp[4]) ? 4'b1001 : 4'b1101;
													assign node9983 = (inp[10]) ? node9989 : node9984;
														assign node9984 = (inp[7]) ? 4'b0101 : node9985;
															assign node9985 = (inp[4]) ? 4'b0001 : 4'b0101;
														assign node9989 = (inp[7]) ? 4'b1101 : node9990;
															assign node9990 = (inp[4]) ? 4'b1001 : 4'b1101;
											assign node9994 = (inp[10]) ? node10018 : node9995;
												assign node9995 = (inp[12]) ? node10007 : node9996;
													assign node9996 = (inp[3]) ? node10002 : node9997;
														assign node9997 = (inp[4]) ? 4'b0101 : node9998;
															assign node9998 = (inp[14]) ? 4'b0001 : 4'b0101;
														assign node10002 = (inp[4]) ? 4'b0001 : node10003;
															assign node10003 = (inp[7]) ? 4'b0101 : 4'b0001;
													assign node10007 = (inp[3]) ? node10013 : node10008;
														assign node10008 = (inp[7]) ? 4'b1001 : node10009;
															assign node10009 = (inp[4]) ? 4'b1101 : 4'b1001;
														assign node10013 = (inp[7]) ? 4'b1101 : node10014;
															assign node10014 = (inp[4]) ? 4'b1001 : 4'b1101;
												assign node10018 = (inp[3]) ? node10024 : node10019;
													assign node10019 = (inp[7]) ? node10021 : 4'b0101;
														assign node10021 = (inp[4]) ? 4'b0101 : 4'b0001;
													assign node10024 = (inp[7]) ? node10026 : 4'b0001;
														assign node10026 = (inp[4]) ? 4'b0001 : 4'b0101;
							assign node10029 = (inp[3]) ? node10031 : 4'b0011;
								assign node10031 = (inp[5]) ? node10033 : 4'b0011;
									assign node10033 = (inp[4]) ? node10061 : node10034;
										assign node10034 = (inp[13]) ? node10036 : 4'b0011;
											assign node10036 = (inp[7]) ? 4'b0011 : node10037;
												assign node10037 = (inp[10]) ? node10045 : node10038;
													assign node10038 = (inp[12]) ? 4'b0011 : node10039;
														assign node10039 = (inp[1]) ? 4'b0001 : node10040;
															assign node10040 = (inp[14]) ? 4'b0011 : 4'b0000;
													assign node10045 = (inp[14]) ? node10047 : 4'b0001;
														assign node10047 = (inp[12]) ? node10055 : node10048;
															assign node10048 = (inp[1]) ? node10052 : node10049;
																assign node10049 = (inp[11]) ? 4'b0000 : 4'b0001;
																assign node10052 = (inp[11]) ? 4'b0001 : 4'b0000;
															assign node10055 = (inp[11]) ? node10057 : 4'b0000;
																assign node10057 = (inp[1]) ? 4'b0001 : 4'b0000;
										assign node10061 = (inp[7]) ? node10117 : node10062;
											assign node10062 = (inp[1]) ? node10088 : node10063;
												assign node10063 = (inp[11]) ? node10077 : node10064;
													assign node10064 = (inp[14]) ? node10070 : node10065;
														assign node10065 = (inp[13]) ? 4'b0000 : node10066;
															assign node10066 = (inp[10]) ? 4'b1000 : 4'b0000;
														assign node10070 = (inp[13]) ? node10072 : 4'b0001;
															assign node10072 = (inp[10]) ? node10074 : 4'b1001;
																assign node10074 = (inp[12]) ? 4'b1001 : 4'b0001;
													assign node10077 = (inp[13]) ? node10083 : node10078;
														assign node10078 = (inp[12]) ? node10080 : 4'b1000;
															assign node10080 = (inp[10]) ? 4'b1000 : 4'b0000;
														assign node10083 = (inp[12]) ? node10085 : 4'b0000;
															assign node10085 = (inp[10]) ? 4'b0000 : 4'b1000;
												assign node10088 = (inp[14]) ? node10100 : node10089;
													assign node10089 = (inp[13]) ? node10095 : node10090;
														assign node10090 = (inp[12]) ? node10092 : 4'b1001;
															assign node10092 = (inp[10]) ? 4'b1001 : 4'b0001;
														assign node10095 = (inp[10]) ? 4'b0001 : node10096;
															assign node10096 = (inp[12]) ? 4'b1001 : 4'b0001;
													assign node10100 = (inp[11]) ? node10106 : node10101;
														assign node10101 = (inp[13]) ? node10103 : 4'b1000;
															assign node10103 = (inp[10]) ? 4'b0000 : 4'b1000;
														assign node10106 = (inp[13]) ? node10112 : node10107;
															assign node10107 = (inp[10]) ? 4'b1001 : node10108;
																assign node10108 = (inp[12]) ? 4'b0001 : 4'b1001;
															assign node10112 = (inp[12]) ? node10114 : 4'b0001;
																assign node10114 = (inp[10]) ? 4'b0001 : 4'b1001;
											assign node10117 = (inp[13]) ? node10119 : 4'b0011;
												assign node10119 = (inp[12]) ? node10133 : node10120;
													assign node10120 = (inp[1]) ? node10128 : node10121;
														assign node10121 = (inp[14]) ? node10123 : 4'b0000;
															assign node10123 = (inp[11]) ? 4'b0000 : node10124;
																assign node10124 = (inp[10]) ? 4'b0001 : 4'b0011;
														assign node10128 = (inp[11]) ? 4'b0001 : node10129;
															assign node10129 = (inp[14]) ? 4'b0000 : 4'b0001;
													assign node10133 = (inp[10]) ? node10135 : 4'b0011;
														assign node10135 = (inp[1]) ? node10139 : node10136;
															assign node10136 = (inp[11]) ? 4'b0000 : 4'b0011;
															assign node10139 = (inp[11]) ? 4'b0001 : node10140;
																assign node10140 = (inp[14]) ? 4'b0000 : 4'b0001;
						assign node10144 = (inp[5]) ? node10926 : node10145;
							assign node10145 = (inp[1]) ? node10579 : node10146;
								assign node10146 = (inp[14]) ? node10354 : node10147;
									assign node10147 = (inp[13]) ? node10239 : node10148;
										assign node10148 = (inp[3]) ? node10176 : node10149;
											assign node10149 = (inp[7]) ? node10171 : node10150;
												assign node10150 = (inp[4]) ? node10156 : node10151;
													assign node10151 = (inp[10]) ? 4'b1000 : node10152;
														assign node10152 = (inp[12]) ? 4'b0000 : 4'b1000;
													assign node10156 = (inp[2]) ? node10166 : node10157;
														assign node10157 = (inp[12]) ? node10163 : node10158;
															assign node10158 = (inp[10]) ? node10160 : 4'b1100;
																assign node10160 = (inp[11]) ? 4'b0001 : 4'b0000;
															assign node10163 = (inp[10]) ? 4'b1100 : 4'b0100;
														assign node10166 = (inp[10]) ? 4'b1100 : node10167;
															assign node10167 = (inp[12]) ? 4'b0100 : 4'b1100;
												assign node10171 = (inp[12]) ? node10173 : 4'b1000;
													assign node10173 = (inp[10]) ? 4'b1000 : 4'b0000;
											assign node10176 = (inp[11]) ? node10204 : node10177;
												assign node10177 = (inp[7]) ? node10189 : node10178;
													assign node10178 = (inp[12]) ? node10182 : node10179;
														assign node10179 = (inp[4]) ? 4'b0000 : 4'b1000;
														assign node10182 = (inp[10]) ? node10184 : 4'b0000;
															assign node10184 = (inp[2]) ? node10186 : 4'b1100;
																assign node10186 = (inp[4]) ? 4'b1000 : 4'b1100;
													assign node10189 = (inp[4]) ? node10199 : node10190;
														assign node10190 = (inp[2]) ? node10196 : node10191;
															assign node10191 = (inp[10]) ? node10193 : 4'b0000;
																assign node10193 = (inp[12]) ? 4'b1000 : 4'b0000;
															assign node10196 = (inp[12]) ? 4'b0100 : 4'b1100;
														assign node10199 = (inp[12]) ? 4'b0100 : node10200;
															assign node10200 = (inp[10]) ? 4'b0100 : 4'b1100;
												assign node10204 = (inp[2]) ? node10220 : node10205;
													assign node10205 = (inp[4]) ? node10211 : node10206;
														assign node10206 = (inp[7]) ? node10208 : 4'b1001;
															assign node10208 = (inp[12]) ? 4'b1001 : 4'b0001;
														assign node10211 = (inp[7]) ? node10213 : 4'b1101;
															assign node10213 = (inp[10]) ? node10217 : node10214;
																assign node10214 = (inp[12]) ? 4'b0101 : 4'b1101;
																assign node10217 = (inp[12]) ? 4'b1101 : 4'b0101;
													assign node10220 = (inp[7]) ? node10234 : node10221;
														assign node10221 = (inp[4]) ? node10227 : node10222;
															assign node10222 = (inp[12]) ? node10224 : 4'b1100;
																assign node10224 = (inp[10]) ? 4'b1100 : 4'b0100;
															assign node10227 = (inp[10]) ? node10231 : node10228;
																assign node10228 = (inp[12]) ? 4'b0000 : 4'b1000;
																assign node10231 = (inp[12]) ? 4'b1000 : 4'b0001;
														assign node10234 = (inp[12]) ? node10236 : 4'b1100;
															assign node10236 = (inp[10]) ? 4'b1100 : 4'b0100;
										assign node10239 = (inp[12]) ? node10301 : node10240;
											assign node10240 = (inp[3]) ? node10264 : node10241;
												assign node10241 = (inp[2]) ? node10259 : node10242;
													assign node10242 = (inp[10]) ? node10252 : node10243;
														assign node10243 = (inp[7]) ? node10249 : node10244;
															assign node10244 = (inp[4]) ? node10246 : 4'b0100;
																assign node10246 = (inp[11]) ? 4'b1001 : 4'b1000;
															assign node10249 = (inp[4]) ? 4'b0100 : 4'b0000;
														assign node10252 = (inp[7]) ? 4'b0000 : node10253;
															assign node10253 = (inp[4]) ? node10255 : 4'b0100;
																assign node10255 = (inp[11]) ? 4'b0001 : 4'b0000;
													assign node10259 = (inp[4]) ? 4'b0100 : node10260;
														assign node10260 = (inp[7]) ? 4'b0000 : 4'b0100;
												assign node10264 = (inp[4]) ? node10278 : node10265;
													assign node10265 = (inp[10]) ? node10273 : node10266;
														assign node10266 = (inp[2]) ? node10270 : node10267;
															assign node10267 = (inp[11]) ? 4'b1001 : 4'b1000;
															assign node10270 = (inp[7]) ? 4'b0100 : 4'b0000;
														assign node10273 = (inp[11]) ? node10275 : 4'b0100;
															assign node10275 = (inp[2]) ? 4'b0100 : 4'b0101;
													assign node10278 = (inp[10]) ? node10292 : node10279;
														assign node10279 = (inp[2]) ? node10287 : node10280;
															assign node10280 = (inp[7]) ? node10284 : node10281;
																assign node10281 = (inp[11]) ? 4'b0000 : 4'b0001;
																assign node10284 = (inp[11]) ? 4'b1101 : 4'b1100;
															assign node10287 = (inp[7]) ? 4'b0000 : node10288;
																assign node10288 = (inp[11]) ? 4'b1001 : 4'b1000;
														assign node10292 = (inp[2]) ? node10298 : node10293;
															assign node10293 = (inp[7]) ? 4'b0000 : node10294;
																assign node10294 = (inp[11]) ? 4'b0000 : 4'b1001;
															assign node10298 = (inp[11]) ? 4'b0001 : 4'b0000;
											assign node10301 = (inp[10]) ? node10319 : node10302;
												assign node10302 = (inp[3]) ? node10308 : node10303;
													assign node10303 = (inp[4]) ? node10305 : 4'b1000;
														assign node10305 = (inp[7]) ? 4'b1000 : 4'b1100;
													assign node10308 = (inp[2]) ? 4'b1100 : node10309;
														assign node10309 = (inp[7]) ? node10313 : node10310;
															assign node10310 = (inp[4]) ? 4'b0000 : 4'b0100;
															assign node10313 = (inp[11]) ? 4'b0101 : node10314;
																assign node10314 = (inp[4]) ? 4'b0100 : 4'b0000;
												assign node10319 = (inp[3]) ? node10329 : node10320;
													assign node10320 = (inp[7]) ? node10326 : node10321;
														assign node10321 = (inp[4]) ? node10323 : 4'b0100;
															assign node10323 = (inp[2]) ? 4'b0100 : 4'b1001;
														assign node10326 = (inp[4]) ? 4'b0100 : 4'b0000;
													assign node10329 = (inp[2]) ? node10345 : node10330;
														assign node10330 = (inp[11]) ? node10338 : node10331;
															assign node10331 = (inp[4]) ? node10335 : node10332;
																assign node10332 = (inp[7]) ? 4'b1000 : 4'b1100;
																assign node10335 = (inp[7]) ? 4'b1100 : 4'b1001;
															assign node10338 = (inp[4]) ? node10342 : node10339;
																assign node10339 = (inp[7]) ? 4'b1001 : 4'b1101;
																assign node10342 = (inp[7]) ? 4'b1101 : 4'b1000;
														assign node10345 = (inp[7]) ? node10351 : node10346;
															assign node10346 = (inp[4]) ? node10348 : 4'b0000;
																assign node10348 = (inp[11]) ? 4'b1001 : 4'b1000;
															assign node10351 = (inp[4]) ? 4'b0000 : 4'b0100;
									assign node10354 = (inp[11]) ? node10462 : node10355;
										assign node10355 = (inp[3]) ? node10399 : node10356;
											assign node10356 = (inp[13]) ? node10372 : node10357;
												assign node10357 = (inp[10]) ? node10363 : node10358;
													assign node10358 = (inp[4]) ? node10360 : 4'b0001;
														assign node10360 = (inp[7]) ? 4'b0001 : 4'b0101;
													assign node10363 = (inp[12]) ? node10369 : node10364;
														assign node10364 = (inp[7]) ? 4'b1001 : node10365;
															assign node10365 = (inp[4]) ? 4'b1101 : 4'b1001;
														assign node10369 = (inp[4]) ? 4'b0101 : 4'b0001;
												assign node10372 = (inp[10]) ? node10386 : node10373;
													assign node10373 = (inp[2]) ? node10381 : node10374;
														assign node10374 = (inp[4]) ? node10376 : 4'b1001;
															assign node10376 = (inp[12]) ? 4'b0000 : node10377;
																assign node10377 = (inp[7]) ? 4'b1001 : 4'b1000;
														assign node10381 = (inp[7]) ? 4'b1001 : node10382;
															assign node10382 = (inp[4]) ? 4'b1101 : 4'b1001;
													assign node10386 = (inp[12]) ? node10394 : node10387;
														assign node10387 = (inp[7]) ? node10389 : 4'b0101;
															assign node10389 = (inp[4]) ? node10391 : 4'b0001;
																assign node10391 = (inp[2]) ? 4'b0101 : 4'b0000;
														assign node10394 = (inp[4]) ? node10396 : 4'b1001;
															assign node10396 = (inp[7]) ? 4'b1001 : 4'b1101;
											assign node10399 = (inp[2]) ? node10435 : node10400;
												assign node10400 = (inp[4]) ? node10420 : node10401;
													assign node10401 = (inp[7]) ? node10413 : node10402;
														assign node10402 = (inp[13]) ? node10408 : node10403;
															assign node10403 = (inp[10]) ? 4'b0100 : node10404;
																assign node10404 = (inp[12]) ? 4'b0000 : 4'b1000;
															assign node10408 = (inp[12]) ? 4'b1100 : node10409;
																assign node10409 = (inp[10]) ? 4'b0100 : 4'b1100;
														assign node10413 = (inp[10]) ? node10417 : node10414;
															assign node10414 = (inp[12]) ? 4'b0000 : 4'b1000;
															assign node10417 = (inp[12]) ? 4'b1000 : 4'b0000;
													assign node10420 = (inp[7]) ? node10428 : node10421;
														assign node10421 = (inp[13]) ? 4'b1000 : node10422;
															assign node10422 = (inp[10]) ? 4'b1100 : node10423;
																assign node10423 = (inp[12]) ? 4'b0100 : 4'b1100;
														assign node10428 = (inp[12]) ? node10432 : node10429;
															assign node10429 = (inp[10]) ? 4'b0100 : 4'b1100;
															assign node10432 = (inp[10]) ? 4'b1100 : 4'b0100;
												assign node10435 = (inp[7]) ? node10449 : node10436;
													assign node10436 = (inp[4]) ? node10444 : node10437;
														assign node10437 = (inp[10]) ? node10439 : 4'b1101;
															assign node10439 = (inp[13]) ? 4'b0001 : node10440;
																assign node10440 = (inp[12]) ? 4'b0101 : 4'b1101;
														assign node10444 = (inp[10]) ? 4'b0000 : node10445;
															assign node10445 = (inp[13]) ? 4'b0000 : 4'b0001;
													assign node10449 = (inp[13]) ? node10455 : node10450;
														assign node10450 = (inp[4]) ? node10452 : 4'b0101;
															assign node10452 = (inp[12]) ? 4'b0101 : 4'b1101;
														assign node10455 = (inp[12]) ? 4'b1101 : node10456;
															assign node10456 = (inp[10]) ? node10458 : 4'b1101;
																assign node10458 = (inp[4]) ? 4'b0000 : 4'b0101;
										assign node10462 = (inp[2]) ? node10530 : node10463;
											assign node10463 = (inp[3]) ? node10493 : node10464;
												assign node10464 = (inp[13]) ? node10480 : node10465;
													assign node10465 = (inp[12]) ? node10477 : node10466;
														assign node10466 = (inp[10]) ? node10472 : node10467;
															assign node10467 = (inp[4]) ? node10469 : 4'b1000;
																assign node10469 = (inp[7]) ? 4'b1000 : 4'b1100;
															assign node10472 = (inp[4]) ? node10474 : 4'b1000;
																assign node10474 = (inp[7]) ? 4'b1000 : 4'b0001;
														assign node10477 = (inp[10]) ? 4'b1000 : 4'b0000;
													assign node10480 = (inp[4]) ? node10484 : node10481;
														assign node10481 = (inp[7]) ? 4'b0000 : 4'b0100;
														assign node10484 = (inp[10]) ? node10490 : node10485;
															assign node10485 = (inp[7]) ? node10487 : 4'b1001;
																assign node10487 = (inp[12]) ? 4'b1000 : 4'b0100;
															assign node10490 = (inp[12]) ? 4'b1001 : 4'b0001;
												assign node10493 = (inp[4]) ? node10517 : node10494;
													assign node10494 = (inp[13]) ? node10504 : node10495;
														assign node10495 = (inp[10]) ? node10499 : node10496;
															assign node10496 = (inp[12]) ? 4'b0001 : 4'b1001;
															assign node10499 = (inp[12]) ? 4'b1001 : node10500;
																assign node10500 = (inp[7]) ? 4'b0001 : 4'b0101;
														assign node10504 = (inp[7]) ? node10510 : node10505;
															assign node10505 = (inp[10]) ? node10507 : 4'b1101;
																assign node10507 = (inp[12]) ? 4'b1101 : 4'b0101;
															assign node10510 = (inp[10]) ? node10514 : node10511;
																assign node10511 = (inp[12]) ? 4'b0001 : 4'b1001;
																assign node10514 = (inp[12]) ? 4'b1001 : 4'b0101;
													assign node10517 = (inp[13]) ? node10523 : node10518;
														assign node10518 = (inp[10]) ? 4'b0001 : node10519;
															assign node10519 = (inp[12]) ? 4'b0101 : 4'b1101;
														assign node10523 = (inp[12]) ? node10525 : 4'b0000;
															assign node10525 = (inp[7]) ? node10527 : 4'b1000;
																assign node10527 = (inp[10]) ? 4'b1101 : 4'b0101;
											assign node10530 = (inp[13]) ? node10550 : node10531;
												assign node10531 = (inp[3]) ? node10541 : node10532;
													assign node10532 = (inp[4]) ? node10538 : node10533;
														assign node10533 = (inp[12]) ? node10535 : 4'b1000;
															assign node10535 = (inp[10]) ? 4'b1000 : 4'b0000;
														assign node10538 = (inp[7]) ? 4'b1000 : 4'b1100;
													assign node10541 = (inp[12]) ? node10543 : 4'b1100;
														assign node10543 = (inp[10]) ? node10547 : node10544;
															assign node10544 = (inp[7]) ? 4'b0100 : 4'b0000;
															assign node10547 = (inp[7]) ? 4'b1100 : 4'b1000;
												assign node10550 = (inp[3]) ? node10568 : node10551;
													assign node10551 = (inp[12]) ? node10557 : node10552;
														assign node10552 = (inp[7]) ? node10554 : 4'b0100;
															assign node10554 = (inp[4]) ? 4'b0100 : 4'b0000;
														assign node10557 = (inp[10]) ? node10563 : node10558;
															assign node10558 = (inp[7]) ? 4'b1000 : node10559;
																assign node10559 = (inp[4]) ? 4'b1100 : 4'b1000;
															assign node10563 = (inp[7]) ? node10565 : 4'b0100;
																assign node10565 = (inp[4]) ? 4'b0100 : 4'b0000;
													assign node10568 = (inp[4]) ? node10576 : node10569;
														assign node10569 = (inp[12]) ? node10571 : 4'b0000;
															assign node10571 = (inp[10]) ? node10573 : 4'b1100;
																assign node10573 = (inp[7]) ? 4'b0100 : 4'b0000;
														assign node10576 = (inp[7]) ? 4'b0000 : 4'b0001;
								assign node10579 = (inp[11]) ? node10789 : node10580;
									assign node10580 = (inp[14]) ? node10684 : node10581;
										assign node10581 = (inp[2]) ? node10627 : node10582;
											assign node10582 = (inp[3]) ? node10608 : node10583;
												assign node10583 = (inp[4]) ? node10593 : node10584;
													assign node10584 = (inp[13]) ? node10590 : node10585;
														assign node10585 = (inp[12]) ? node10587 : 4'b1001;
															assign node10587 = (inp[10]) ? 4'b1001 : 4'b0001;
														assign node10590 = (inp[10]) ? 4'b0101 : 4'b1001;
													assign node10593 = (inp[10]) ? node10603 : node10594;
														assign node10594 = (inp[7]) ? node10598 : node10595;
															assign node10595 = (inp[13]) ? 4'b1000 : 4'b0101;
															assign node10598 = (inp[13]) ? node10600 : 4'b1001;
																assign node10600 = (inp[12]) ? 4'b1001 : 4'b0101;
														assign node10603 = (inp[13]) ? 4'b0000 : node10604;
															assign node10604 = (inp[7]) ? 4'b1001 : 4'b0000;
												assign node10608 = (inp[10]) ? node10616 : node10609;
													assign node10609 = (inp[4]) ? 4'b1100 : node10610;
														assign node10610 = (inp[7]) ? 4'b1000 : node10611;
															assign node10611 = (inp[13]) ? 4'b1100 : 4'b1000;
													assign node10616 = (inp[4]) ? node10622 : node10617;
														assign node10617 = (inp[13]) ? 4'b0100 : node10618;
															assign node10618 = (inp[7]) ? 4'b0000 : 4'b0100;
														assign node10622 = (inp[7]) ? node10624 : 4'b0000;
															assign node10624 = (inp[13]) ? 4'b0000 : 4'b0100;
											assign node10627 = (inp[13]) ? node10655 : node10628;
												assign node10628 = (inp[3]) ? node10642 : node10629;
													assign node10629 = (inp[4]) ? node10635 : node10630;
														assign node10630 = (inp[12]) ? node10632 : 4'b1001;
															assign node10632 = (inp[10]) ? 4'b1001 : 4'b0001;
														assign node10635 = (inp[7]) ? 4'b1001 : node10636;
															assign node10636 = (inp[12]) ? node10638 : 4'b1101;
																assign node10638 = (inp[10]) ? 4'b1101 : 4'b0101;
													assign node10642 = (inp[12]) ? node10648 : node10643;
														assign node10643 = (inp[7]) ? 4'b1101 : node10644;
															assign node10644 = (inp[4]) ? 4'b1001 : 4'b1101;
														assign node10648 = (inp[10]) ? 4'b1101 : node10649;
															assign node10649 = (inp[7]) ? 4'b0101 : node10650;
																assign node10650 = (inp[4]) ? 4'b0001 : 4'b0101;
												assign node10655 = (inp[10]) ? node10673 : node10656;
													assign node10656 = (inp[12]) ? node10666 : node10657;
														assign node10657 = (inp[3]) ? node10661 : node10658;
															assign node10658 = (inp[4]) ? 4'b0101 : 4'b0001;
															assign node10661 = (inp[7]) ? 4'b0001 : node10662;
																assign node10662 = (inp[4]) ? 4'b1000 : 4'b0001;
														assign node10666 = (inp[3]) ? 4'b1101 : node10667;
															assign node10667 = (inp[7]) ? 4'b1001 : node10668;
																assign node10668 = (inp[4]) ? 4'b1101 : 4'b1001;
													assign node10673 = (inp[3]) ? node10679 : node10674;
														assign node10674 = (inp[4]) ? 4'b0101 : node10675;
															assign node10675 = (inp[7]) ? 4'b0001 : 4'b0101;
														assign node10679 = (inp[4]) ? 4'b0000 : node10680;
															assign node10680 = (inp[7]) ? 4'b0101 : 4'b0001;
										assign node10684 = (inp[10]) ? node10746 : node10685;
											assign node10685 = (inp[3]) ? node10713 : node10686;
												assign node10686 = (inp[4]) ? node10694 : node10687;
													assign node10687 = (inp[12]) ? node10691 : node10688;
														assign node10688 = (inp[13]) ? 4'b0000 : 4'b1000;
														assign node10691 = (inp[13]) ? 4'b1000 : 4'b0000;
													assign node10694 = (inp[7]) ? node10706 : node10695;
														assign node10695 = (inp[2]) ? node10699 : node10696;
															assign node10696 = (inp[13]) ? 4'b1000 : 4'b1100;
															assign node10699 = (inp[12]) ? node10703 : node10700;
																assign node10700 = (inp[13]) ? 4'b0100 : 4'b1100;
																assign node10703 = (inp[13]) ? 4'b1100 : 4'b0100;
														assign node10706 = (inp[12]) ? node10710 : node10707;
															assign node10707 = (inp[13]) ? 4'b0100 : 4'b1000;
															assign node10710 = (inp[13]) ? 4'b1000 : 4'b0000;
												assign node10713 = (inp[2]) ? node10725 : node10714;
													assign node10714 = (inp[4]) ? node10720 : node10715;
														assign node10715 = (inp[7]) ? 4'b1000 : node10716;
															assign node10716 = (inp[13]) ? 4'b1100 : 4'b1000;
														assign node10720 = (inp[13]) ? node10722 : 4'b1100;
															assign node10722 = (inp[7]) ? 4'b1100 : 4'b0001;
													assign node10725 = (inp[4]) ? node10733 : node10726;
														assign node10726 = (inp[13]) ? node10730 : node10727;
															assign node10727 = (inp[12]) ? 4'b0100 : 4'b1100;
															assign node10730 = (inp[12]) ? 4'b1100 : 4'b0100;
														assign node10733 = (inp[7]) ? node10739 : node10734;
															assign node10734 = (inp[12]) ? node10736 : 4'b1000;
																assign node10736 = (inp[13]) ? 4'b1000 : 4'b0000;
															assign node10739 = (inp[13]) ? node10743 : node10740;
																assign node10740 = (inp[12]) ? 4'b0100 : 4'b1100;
																assign node10743 = (inp[12]) ? 4'b1100 : 4'b0000;
											assign node10746 = (inp[13]) ? node10766 : node10747;
												assign node10747 = (inp[3]) ? node10753 : node10748;
													assign node10748 = (inp[4]) ? node10750 : 4'b1000;
														assign node10750 = (inp[7]) ? 4'b1000 : 4'b0000;
													assign node10753 = (inp[2]) ? node10761 : node10754;
														assign node10754 = (inp[7]) ? node10758 : node10755;
															assign node10755 = (inp[4]) ? 4'b0000 : 4'b0100;
															assign node10758 = (inp[4]) ? 4'b0100 : 4'b0000;
														assign node10761 = (inp[4]) ? node10763 : 4'b1100;
															assign node10763 = (inp[7]) ? 4'b1100 : 4'b0000;
												assign node10766 = (inp[4]) ? node10776 : node10767;
													assign node10767 = (inp[3]) ? node10771 : node10768;
														assign node10768 = (inp[7]) ? 4'b0000 : 4'b0100;
														assign node10771 = (inp[7]) ? 4'b0100 : node10772;
															assign node10772 = (inp[2]) ? 4'b0000 : 4'b0100;
													assign node10776 = (inp[2]) ? node10786 : node10777;
														assign node10777 = (inp[3]) ? node10779 : 4'b0000;
															assign node10779 = (inp[7]) ? node10783 : node10780;
																assign node10780 = (inp[12]) ? 4'b1001 : 4'b0001;
																assign node10783 = (inp[12]) ? 4'b0000 : 4'b0001;
														assign node10786 = (inp[3]) ? 4'b0000 : 4'b0100;
									assign node10789 = (inp[10]) ? node10873 : node10790;
										assign node10790 = (inp[3]) ? node10836 : node10791;
											assign node10791 = (inp[7]) ? node10813 : node10792;
												assign node10792 = (inp[4]) ? node10800 : node10793;
													assign node10793 = (inp[12]) ? node10797 : node10794;
														assign node10794 = (inp[13]) ? 4'b0101 : 4'b1001;
														assign node10797 = (inp[13]) ? 4'b1001 : 4'b0001;
													assign node10800 = (inp[2]) ? node10806 : node10801;
														assign node10801 = (inp[13]) ? 4'b1001 : node10802;
															assign node10802 = (inp[12]) ? 4'b0101 : 4'b1101;
														assign node10806 = (inp[13]) ? node10810 : node10807;
															assign node10807 = (inp[12]) ? 4'b0101 : 4'b1101;
															assign node10810 = (inp[12]) ? 4'b1101 : 4'b0101;
												assign node10813 = (inp[4]) ? node10829 : node10814;
													assign node10814 = (inp[14]) ? node10822 : node10815;
														assign node10815 = (inp[12]) ? node10819 : node10816;
															assign node10816 = (inp[13]) ? 4'b0001 : 4'b1001;
															assign node10819 = (inp[13]) ? 4'b1001 : 4'b0001;
														assign node10822 = (inp[12]) ? node10826 : node10823;
															assign node10823 = (inp[13]) ? 4'b0001 : 4'b1001;
															assign node10826 = (inp[13]) ? 4'b1001 : 4'b0001;
													assign node10829 = (inp[12]) ? node10833 : node10830;
														assign node10830 = (inp[13]) ? 4'b0101 : 4'b1001;
														assign node10833 = (inp[13]) ? 4'b1001 : 4'b0001;
											assign node10836 = (inp[2]) ? node10848 : node10837;
												assign node10837 = (inp[4]) ? node10843 : node10838;
													assign node10838 = (inp[13]) ? node10840 : 4'b1001;
														assign node10840 = (inp[7]) ? 4'b1001 : 4'b1101;
													assign node10843 = (inp[7]) ? 4'b1101 : node10844;
														assign node10844 = (inp[13]) ? 4'b1001 : 4'b1101;
												assign node10848 = (inp[7]) ? node10864 : node10849;
													assign node10849 = (inp[4]) ? node10859 : node10850;
														assign node10850 = (inp[14]) ? node10854 : node10851;
															assign node10851 = (inp[12]) ? 4'b0101 : 4'b0001;
															assign node10854 = (inp[13]) ? 4'b1101 : node10855;
																assign node10855 = (inp[12]) ? 4'b0101 : 4'b1101;
														assign node10859 = (inp[13]) ? 4'b1001 : node10860;
															assign node10860 = (inp[12]) ? 4'b0001 : 4'b1001;
													assign node10864 = (inp[12]) ? node10870 : node10865;
														assign node10865 = (inp[13]) ? node10867 : 4'b1101;
															assign node10867 = (inp[4]) ? 4'b0001 : 4'b0101;
														assign node10870 = (inp[13]) ? 4'b1101 : 4'b0101;
										assign node10873 = (inp[13]) ? node10911 : node10874;
											assign node10874 = (inp[3]) ? node10884 : node10875;
												assign node10875 = (inp[7]) ? 4'b1001 : node10876;
													assign node10876 = (inp[2]) ? node10880 : node10877;
														assign node10877 = (inp[4]) ? 4'b0001 : 4'b1001;
														assign node10880 = (inp[4]) ? 4'b1101 : 4'b1001;
												assign node10884 = (inp[2]) ? node10906 : node10885;
													assign node10885 = (inp[12]) ? node10901 : node10886;
														assign node10886 = (inp[14]) ? node10894 : node10887;
															assign node10887 = (inp[4]) ? node10891 : node10888;
																assign node10888 = (inp[7]) ? 4'b0001 : 4'b0101;
																assign node10891 = (inp[7]) ? 4'b0101 : 4'b0001;
															assign node10894 = (inp[4]) ? node10898 : node10895;
																assign node10895 = (inp[7]) ? 4'b0001 : 4'b0101;
																assign node10898 = (inp[7]) ? 4'b0101 : 4'b0001;
														assign node10901 = (inp[7]) ? 4'b0001 : node10902;
															assign node10902 = (inp[4]) ? 4'b0001 : 4'b0101;
													assign node10906 = (inp[4]) ? node10908 : 4'b1101;
														assign node10908 = (inp[7]) ? 4'b1101 : 4'b0001;
											assign node10911 = (inp[4]) ? node10921 : node10912;
												assign node10912 = (inp[3]) ? node10916 : node10913;
													assign node10913 = (inp[7]) ? 4'b0001 : 4'b0101;
													assign node10916 = (inp[7]) ? 4'b0101 : node10917;
														assign node10917 = (inp[2]) ? 4'b0001 : 4'b0101;
												assign node10921 = (inp[2]) ? node10923 : 4'b0001;
													assign node10923 = (inp[3]) ? 4'b0001 : 4'b0101;
							assign node10926 = (inp[3]) ? node11348 : node10927;
								assign node10927 = (inp[11]) ? node11193 : node10928;
									assign node10928 = (inp[4]) ? node11054 : node10929;
										assign node10929 = (inp[2]) ? node11005 : node10930;
											assign node10930 = (inp[13]) ? node10970 : node10931;
												assign node10931 = (inp[7]) ? node10949 : node10932;
													assign node10932 = (inp[10]) ? node10942 : node10933;
														assign node10933 = (inp[14]) ? node10937 : node10934;
															assign node10934 = (inp[12]) ? 4'b1000 : 4'b0100;
															assign node10937 = (inp[1]) ? 4'b1001 : node10938;
																assign node10938 = (inp[12]) ? 4'b0000 : 4'b1000;
														assign node10942 = (inp[1]) ? node10946 : node10943;
															assign node10943 = (inp[14]) ? 4'b0100 : 4'b0101;
															assign node10946 = (inp[14]) ? 4'b0101 : 4'b1100;
													assign node10949 = (inp[10]) ? node10963 : node10950;
														assign node10950 = (inp[12]) ? node10958 : node10951;
															assign node10951 = (inp[1]) ? node10955 : node10952;
																assign node10952 = (inp[14]) ? 4'b1000 : 4'b1001;
																assign node10955 = (inp[14]) ? 4'b1001 : 4'b0000;
															assign node10958 = (inp[1]) ? 4'b1001 : node10959;
																assign node10959 = (inp[14]) ? 4'b0000 : 4'b0001;
														assign node10963 = (inp[1]) ? node10967 : node10964;
															assign node10964 = (inp[14]) ? 4'b0000 : 4'b0001;
															assign node10967 = (inp[14]) ? 4'b0001 : 4'b1000;
												assign node10970 = (inp[10]) ? node10988 : node10971;
													assign node10971 = (inp[12]) ? node10979 : node10972;
														assign node10972 = (inp[1]) ? node10976 : node10973;
															assign node10973 = (inp[14]) ? 4'b0100 : 4'b0101;
															assign node10976 = (inp[7]) ? 4'b0101 : 4'b0001;
														assign node10979 = (inp[1]) ? node10985 : node10980;
															assign node10980 = (inp[7]) ? node10982 : 4'b1101;
																assign node10982 = (inp[14]) ? 4'b1000 : 4'b1001;
															assign node10985 = (inp[14]) ? 4'b0101 : 4'b0100;
													assign node10988 = (inp[7]) ? node10996 : node10989;
														assign node10989 = (inp[12]) ? node10993 : node10990;
															assign node10990 = (inp[1]) ? 4'b0001 : 4'b1001;
															assign node10993 = (inp[1]) ? 4'b1001 : 4'b0001;
														assign node10996 = (inp[1]) ? node11000 : node10997;
															assign node10997 = (inp[14]) ? 4'b1100 : 4'b1101;
															assign node11000 = (inp[12]) ? node11002 : 4'b0001;
																assign node11002 = (inp[14]) ? 4'b1101 : 4'b0100;
											assign node11005 = (inp[10]) ? node11023 : node11006;
												assign node11006 = (inp[13]) ? node11012 : node11007;
													assign node11007 = (inp[12]) ? node11009 : 4'b1000;
														assign node11009 = (inp[1]) ? 4'b1000 : 4'b0000;
													assign node11012 = (inp[7]) ? node11018 : node11013;
														assign node11013 = (inp[1]) ? 4'b1100 : node11014;
															assign node11014 = (inp[12]) ? 4'b0100 : 4'b1100;
														assign node11018 = (inp[14]) ? 4'b1000 : node11019;
															assign node11019 = (inp[12]) ? 4'b0000 : 4'b1000;
												assign node11023 = (inp[12]) ? node11041 : node11024;
													assign node11024 = (inp[1]) ? node11030 : node11025;
														assign node11025 = (inp[13]) ? 4'b0100 : node11026;
															assign node11026 = (inp[7]) ? 4'b0000 : 4'b0100;
														assign node11030 = (inp[14]) ? node11036 : node11031;
															assign node11031 = (inp[7]) ? 4'b0100 : node11032;
																assign node11032 = (inp[13]) ? 4'b0000 : 4'b0100;
															assign node11036 = (inp[13]) ? 4'b0001 : node11037;
																assign node11037 = (inp[7]) ? 4'b0000 : 4'b0100;
													assign node11041 = (inp[1]) ? node11047 : node11042;
														assign node11042 = (inp[7]) ? 4'b1000 : node11043;
															assign node11043 = (inp[13]) ? 4'b1100 : 4'b1000;
														assign node11047 = (inp[13]) ? node11051 : node11048;
															assign node11048 = (inp[7]) ? 4'b0000 : 4'b0100;
															assign node11051 = (inp[14]) ? 4'b0100 : 4'b0000;
										assign node11054 = (inp[1]) ? node11124 : node11055;
											assign node11055 = (inp[12]) ? node11089 : node11056;
												assign node11056 = (inp[13]) ? node11072 : node11057;
													assign node11057 = (inp[10]) ? node11065 : node11058;
														assign node11058 = (inp[2]) ? node11060 : 4'b1001;
															assign node11060 = (inp[7]) ? 4'b1100 : node11061;
																assign node11061 = (inp[14]) ? 4'b1000 : 4'b1001;
														assign node11065 = (inp[2]) ? node11069 : node11066;
															assign node11066 = (inp[14]) ? 4'b1101 : 4'b0000;
															assign node11069 = (inp[14]) ? 4'b0000 : 4'b0001;
													assign node11072 = (inp[10]) ? node11082 : node11073;
														assign node11073 = (inp[7]) ? node11075 : 4'b0100;
															assign node11075 = (inp[14]) ? node11079 : node11076;
																assign node11076 = (inp[2]) ? 4'b0001 : 4'b0000;
																assign node11079 = (inp[2]) ? 4'b0000 : 4'b0001;
														assign node11082 = (inp[2]) ? 4'b1001 : node11083;
															assign node11083 = (inp[14]) ? 4'b0001 : node11084;
																assign node11084 = (inp[7]) ? 4'b1000 : 4'b0000;
												assign node11089 = (inp[13]) ? node11103 : node11090;
													assign node11090 = (inp[2]) ? node11096 : node11091;
														assign node11091 = (inp[7]) ? 4'b0001 : node11092;
															assign node11092 = (inp[10]) ? 4'b0101 : 4'b0001;
														assign node11096 = (inp[14]) ? node11098 : 4'b0001;
															assign node11098 = (inp[7]) ? node11100 : 4'b0000;
																assign node11100 = (inp[10]) ? 4'b0000 : 4'b0100;
													assign node11103 = (inp[2]) ? node11113 : node11104;
														assign node11104 = (inp[14]) ? node11106 : 4'b0000;
															assign node11106 = (inp[10]) ? node11110 : node11107;
																assign node11107 = (inp[7]) ? 4'b0101 : 4'b1001;
																assign node11110 = (inp[7]) ? 4'b0001 : 4'b0000;
														assign node11113 = (inp[14]) ? node11119 : node11114;
															assign node11114 = (inp[7]) ? 4'b1001 : node11115;
																assign node11115 = (inp[10]) ? 4'b0001 : 4'b1001;
															assign node11119 = (inp[10]) ? node11121 : 4'b1000;
																assign node11121 = (inp[7]) ? 4'b1000 : 4'b0001;
											assign node11124 = (inp[12]) ? node11156 : node11125;
												assign node11125 = (inp[13]) ? node11143 : node11126;
													assign node11126 = (inp[2]) ? node11136 : node11127;
														assign node11127 = (inp[7]) ? node11133 : node11128;
															assign node11128 = (inp[10]) ? node11130 : 4'b0101;
																assign node11130 = (inp[14]) ? 4'b1000 : 4'b1001;
															assign node11133 = (inp[10]) ? 4'b0101 : 4'b0001;
														assign node11136 = (inp[14]) ? node11140 : node11137;
															assign node11137 = (inp[10]) ? 4'b1000 : 4'b0000;
															assign node11140 = (inp[10]) ? 4'b1001 : 4'b1100;
													assign node11143 = (inp[2]) ? node11149 : node11144;
														assign node11144 = (inp[10]) ? 4'b0000 : node11145;
															assign node11145 = (inp[14]) ? 4'b1000 : 4'b1001;
														assign node11149 = (inp[14]) ? 4'b0001 : node11150;
															assign node11150 = (inp[7]) ? node11152 : 4'b0001;
																assign node11152 = (inp[10]) ? 4'b0001 : 4'b1000;
												assign node11156 = (inp[2]) ? node11172 : node11157;
													assign node11157 = (inp[13]) ? node11165 : node11158;
														assign node11158 = (inp[10]) ? node11160 : 4'b1001;
															assign node11160 = (inp[7]) ? 4'b1001 : node11161;
																assign node11161 = (inp[14]) ? 4'b0000 : 4'b0001;
														assign node11165 = (inp[14]) ? 4'b1000 : node11166;
															assign node11166 = (inp[10]) ? node11168 : 4'b1001;
																assign node11168 = (inp[7]) ? 4'b1001 : 4'b1000;
													assign node11172 = (inp[14]) ? node11184 : node11173;
														assign node11173 = (inp[7]) ? node11177 : node11174;
															assign node11174 = (inp[13]) ? 4'b1001 : 4'b1000;
															assign node11177 = (inp[13]) ? node11181 : node11178;
																assign node11178 = (inp[10]) ? 4'b1000 : 4'b1100;
																assign node11181 = (inp[10]) ? 4'b0100 : 4'b0000;
														assign node11184 = (inp[10]) ? node11190 : node11185;
															assign node11185 = (inp[13]) ? node11187 : 4'b1100;
																assign node11187 = (inp[7]) ? 4'b0001 : 4'b0101;
															assign node11190 = (inp[13]) ? 4'b1001 : 4'b0001;
									assign node11193 = (inp[1]) ? node11283 : node11194;
										assign node11194 = (inp[13]) ? node11234 : node11195;
											assign node11195 = (inp[2]) ? node11209 : node11196;
												assign node11196 = (inp[4]) ? node11204 : node11197;
													assign node11197 = (inp[10]) ? node11199 : 4'b1000;
														assign node11199 = (inp[12]) ? 4'b0100 : node11200;
															assign node11200 = (inp[7]) ? 4'b1000 : 4'b1100;
													assign node11204 = (inp[7]) ? 4'b1001 : node11205;
														assign node11205 = (inp[12]) ? 4'b0000 : 4'b1001;
												assign node11209 = (inp[4]) ? node11225 : node11210;
													assign node11210 = (inp[7]) ? node11218 : node11211;
														assign node11211 = (inp[12]) ? node11215 : node11212;
															assign node11212 = (inp[10]) ? 4'b0101 : 4'b1001;
															assign node11215 = (inp[10]) ? 4'b1001 : 4'b0001;
														assign node11218 = (inp[10]) ? node11222 : node11219;
															assign node11219 = (inp[12]) ? 4'b0001 : 4'b1001;
															assign node11222 = (inp[12]) ? 4'b1001 : 4'b0001;
													assign node11225 = (inp[10]) ? node11231 : node11226;
														assign node11226 = (inp[7]) ? node11228 : 4'b1000;
															assign node11228 = (inp[12]) ? 4'b0101 : 4'b1101;
														assign node11231 = (inp[12]) ? 4'b0000 : 4'b1000;
											assign node11234 = (inp[10]) ? node11256 : node11235;
												assign node11235 = (inp[7]) ? node11245 : node11236;
													assign node11236 = (inp[2]) ? node11240 : node11237;
														assign node11237 = (inp[4]) ? 4'b1000 : 4'b0100;
														assign node11240 = (inp[4]) ? 4'b0100 : node11241;
															assign node11241 = (inp[12]) ? 4'b0101 : 4'b1101;
													assign node11245 = (inp[2]) ? node11251 : node11246;
														assign node11246 = (inp[4]) ? node11248 : 4'b0100;
															assign node11248 = (inp[12]) ? 4'b0000 : 4'b1000;
														assign node11251 = (inp[4]) ? 4'b0000 : node11252;
															assign node11252 = (inp[12]) ? 4'b0001 : 4'b1001;
												assign node11256 = (inp[7]) ? node11268 : node11257;
													assign node11257 = (inp[4]) ? node11263 : node11258;
														assign node11258 = (inp[12]) ? node11260 : 4'b0000;
															assign node11260 = (inp[2]) ? 4'b1101 : 4'b1001;
														assign node11263 = (inp[12]) ? node11265 : 4'b1001;
															assign node11265 = (inp[2]) ? 4'b1001 : 4'b0001;
													assign node11268 = (inp[12]) ? node11276 : node11269;
														assign node11269 = (inp[4]) ? node11273 : node11270;
															assign node11270 = (inp[2]) ? 4'b0101 : 4'b0100;
															assign node11273 = (inp[2]) ? 4'b0100 : 4'b1000;
														assign node11276 = (inp[2]) ? node11280 : node11277;
															assign node11277 = (inp[4]) ? 4'b1000 : 4'b1100;
															assign node11280 = (inp[4]) ? 4'b1000 : 4'b1001;
										assign node11283 = (inp[13]) ? node11321 : node11284;
											assign node11284 = (inp[12]) ? node11302 : node11285;
												assign node11285 = (inp[10]) ? node11293 : node11286;
													assign node11286 = (inp[2]) ? node11290 : node11287;
														assign node11287 = (inp[7]) ? 4'b0001 : 4'b0101;
														assign node11290 = (inp[4]) ? 4'b0001 : 4'b1001;
													assign node11293 = (inp[4]) ? 4'b1001 : node11294;
														assign node11294 = (inp[7]) ? node11298 : node11295;
															assign node11295 = (inp[14]) ? 4'b1101 : 4'b0101;
															assign node11298 = (inp[2]) ? 4'b0001 : 4'b1001;
												assign node11302 = (inp[4]) ? node11310 : node11303;
													assign node11303 = (inp[10]) ? node11305 : 4'b1001;
														assign node11305 = (inp[2]) ? 4'b0001 : node11306;
															assign node11306 = (inp[7]) ? 4'b1001 : 4'b1101;
													assign node11310 = (inp[10]) ? node11316 : node11311;
														assign node11311 = (inp[2]) ? node11313 : 4'b0101;
															assign node11313 = (inp[7]) ? 4'b1101 : 4'b1001;
														assign node11316 = (inp[2]) ? 4'b1001 : node11317;
															assign node11317 = (inp[7]) ? 4'b0101 : 4'b1001;
											assign node11321 = (inp[10]) ? node11341 : node11322;
												assign node11322 = (inp[4]) ? node11330 : node11323;
													assign node11323 = (inp[2]) ? node11327 : node11324;
														assign node11324 = (inp[7]) ? 4'b1101 : 4'b0001;
														assign node11327 = (inp[7]) ? 4'b1001 : 4'b1101;
													assign node11330 = (inp[2]) ? node11336 : node11331;
														assign node11331 = (inp[12]) ? 4'b1001 : node11332;
															assign node11332 = (inp[7]) ? 4'b0001 : 4'b0101;
														assign node11336 = (inp[12]) ? 4'b0001 : node11337;
															assign node11337 = (inp[14]) ? 4'b1001 : 4'b0001;
												assign node11341 = (inp[4]) ? 4'b0001 : node11342;
													assign node11342 = (inp[7]) ? node11344 : 4'b0001;
														assign node11344 = (inp[2]) ? 4'b0101 : 4'b0001;
								assign node11348 = (inp[4]) ? node11568 : node11349;
									assign node11349 = (inp[1]) ? node11461 : node11350;
										assign node11350 = (inp[11]) ? node11414 : node11351;
											assign node11351 = (inp[12]) ? node11379 : node11352;
												assign node11352 = (inp[13]) ? node11364 : node11353;
													assign node11353 = (inp[2]) ? node11359 : node11354;
														assign node11354 = (inp[14]) ? 4'b1000 : node11355;
															assign node11355 = (inp[10]) ? 4'b1001 : 4'b1000;
														assign node11359 = (inp[10]) ? node11361 : 4'b1001;
															assign node11361 = (inp[14]) ? 4'b1001 : 4'b0000;
													assign node11364 = (inp[10]) ? node11374 : node11365;
														assign node11365 = (inp[2]) ? node11369 : node11366;
															assign node11366 = (inp[7]) ? 4'b1001 : 4'b0001;
															assign node11369 = (inp[7]) ? node11371 : 4'b1000;
																assign node11371 = (inp[14]) ? 4'b0001 : 4'b0000;
														assign node11374 = (inp[2]) ? 4'b0001 : node11375;
															assign node11375 = (inp[7]) ? 4'b1000 : 4'b0000;
												assign node11379 = (inp[10]) ? node11395 : node11380;
													assign node11380 = (inp[14]) ? node11388 : node11381;
														assign node11381 = (inp[13]) ? node11383 : 4'b1000;
															assign node11383 = (inp[2]) ? node11385 : 4'b0000;
																assign node11385 = (inp[7]) ? 4'b0000 : 4'b1000;
														assign node11388 = (inp[13]) ? node11392 : node11389;
															assign node11389 = (inp[2]) ? 4'b0001 : 4'b1000;
															assign node11392 = (inp[7]) ? 4'b1001 : 4'b0001;
													assign node11395 = (inp[13]) ? node11407 : node11396;
														assign node11396 = (inp[7]) ? node11402 : node11397;
															assign node11397 = (inp[2]) ? node11399 : 4'b0001;
																assign node11399 = (inp[14]) ? 4'b1001 : 4'b1000;
															assign node11402 = (inp[2]) ? 4'b0001 : node11403;
																assign node11403 = (inp[14]) ? 4'b0000 : 4'b0001;
														assign node11407 = (inp[14]) ? node11411 : node11408;
															assign node11408 = (inp[7]) ? 4'b0000 : 4'b0001;
															assign node11411 = (inp[2]) ? 4'b1000 : 4'b0000;
											assign node11414 = (inp[12]) ? node11436 : node11415;
												assign node11415 = (inp[2]) ? node11425 : node11416;
													assign node11416 = (inp[13]) ? 4'b0000 : node11417;
														assign node11417 = (inp[10]) ? node11421 : node11418;
															assign node11418 = (inp[7]) ? 4'b0001 : 4'b0000;
															assign node11421 = (inp[7]) ? 4'b0000 : 4'b0001;
													assign node11425 = (inp[10]) ? node11431 : node11426;
														assign node11426 = (inp[13]) ? 4'b0001 : node11427;
															assign node11427 = (inp[7]) ? 4'b1001 : 4'b0000;
														assign node11431 = (inp[13]) ? node11433 : 4'b0000;
															assign node11433 = (inp[7]) ? 4'b1000 : 4'b0001;
												assign node11436 = (inp[2]) ? node11450 : node11437;
													assign node11437 = (inp[7]) ? node11443 : node11438;
														assign node11438 = (inp[13]) ? 4'b1000 : node11439;
															assign node11439 = (inp[10]) ? 4'b0001 : 4'b0000;
														assign node11443 = (inp[10]) ? node11447 : node11444;
															assign node11444 = (inp[13]) ? 4'b0001 : 4'b1001;
															assign node11447 = (inp[13]) ? 4'b1001 : 4'b1000;
													assign node11450 = (inp[10]) ? node11456 : node11451;
														assign node11451 = (inp[13]) ? node11453 : 4'b1001;
															assign node11453 = (inp[7]) ? 4'b0000 : 4'b1001;
														assign node11456 = (inp[13]) ? node11458 : 4'b0000;
															assign node11458 = (inp[7]) ? 4'b0000 : 4'b0001;
										assign node11461 = (inp[11]) ? node11535 : node11462;
											assign node11462 = (inp[10]) ? node11498 : node11463;
												assign node11463 = (inp[2]) ? node11481 : node11464;
													assign node11464 = (inp[13]) ? node11474 : node11465;
														assign node11465 = (inp[12]) ? node11471 : node11466;
															assign node11466 = (inp[14]) ? node11468 : 4'b1000;
																assign node11468 = (inp[7]) ? 4'b1000 : 4'b1001;
															assign node11471 = (inp[7]) ? 4'b0000 : 4'b1000;
														assign node11474 = (inp[7]) ? node11476 : 4'b0000;
															assign node11476 = (inp[14]) ? 4'b1000 : node11477;
																assign node11477 = (inp[12]) ? 4'b0001 : 4'b1001;
													assign node11481 = (inp[13]) ? node11491 : node11482;
														assign node11482 = (inp[14]) ? node11488 : node11483;
															assign node11483 = (inp[12]) ? node11485 : 4'b0001;
																assign node11485 = (inp[7]) ? 4'b1001 : 4'b0001;
															assign node11488 = (inp[12]) ? 4'b0000 : 4'b0001;
														assign node11491 = (inp[12]) ? 4'b0000 : node11492;
															assign node11492 = (inp[7]) ? 4'b1000 : node11493;
																assign node11493 = (inp[14]) ? 4'b0001 : 4'b0000;
												assign node11498 = (inp[7]) ? node11516 : node11499;
													assign node11499 = (inp[12]) ? node11501 : 4'b1001;
														assign node11501 = (inp[14]) ? node11509 : node11502;
															assign node11502 = (inp[13]) ? node11506 : node11503;
																assign node11503 = (inp[2]) ? 4'b0001 : 4'b1001;
																assign node11506 = (inp[2]) ? 4'b1001 : 4'b0001;
															assign node11509 = (inp[13]) ? node11513 : node11510;
																assign node11510 = (inp[2]) ? 4'b0000 : 4'b1001;
																assign node11513 = (inp[2]) ? 4'b1001 : 4'b0001;
													assign node11516 = (inp[14]) ? node11524 : node11517;
														assign node11517 = (inp[2]) ? node11519 : 4'b1000;
															assign node11519 = (inp[13]) ? 4'b0000 : node11520;
																assign node11520 = (inp[12]) ? 4'b0001 : 4'b1001;
														assign node11524 = (inp[13]) ? node11530 : node11525;
															assign node11525 = (inp[2]) ? node11527 : 4'b0001;
																assign node11527 = (inp[12]) ? 4'b0000 : 4'b1000;
															assign node11530 = (inp[2]) ? 4'b1001 : node11531;
																assign node11531 = (inp[12]) ? 4'b0001 : 4'b1001;
											assign node11535 = (inp[10]) ? node11561 : node11536;
												assign node11536 = (inp[13]) ? node11550 : node11537;
													assign node11537 = (inp[7]) ? node11545 : node11538;
														assign node11538 = (inp[2]) ? node11542 : node11539;
															assign node11539 = (inp[12]) ? 4'b1001 : 4'b0001;
															assign node11542 = (inp[12]) ? 4'b0001 : 4'b1001;
														assign node11545 = (inp[2]) ? 4'b0001 : node11546;
															assign node11546 = (inp[12]) ? 4'b1001 : 4'b0001;
													assign node11550 = (inp[12]) ? node11556 : node11551;
														assign node11551 = (inp[2]) ? 4'b1001 : node11552;
															assign node11552 = (inp[7]) ? 4'b0001 : 4'b1001;
														assign node11556 = (inp[7]) ? 4'b1001 : node11557;
															assign node11557 = (inp[2]) ? 4'b0001 : 4'b1001;
												assign node11561 = (inp[2]) ? node11563 : 4'b0001;
													assign node11563 = (inp[7]) ? node11565 : 4'b0001;
														assign node11565 = (inp[13]) ? 4'b0001 : 4'b1001;
									assign node11568 = (inp[13]) ? node11686 : node11569;
										assign node11569 = (inp[1]) ? node11639 : node11570;
											assign node11570 = (inp[2]) ? node11604 : node11571;
												assign node11571 = (inp[7]) ? node11579 : node11572;
													assign node11572 = (inp[11]) ? 4'b0000 : node11573;
														assign node11573 = (inp[14]) ? 4'b0000 : node11574;
															assign node11574 = (inp[10]) ? 4'b0001 : 4'b0000;
													assign node11579 = (inp[14]) ? node11595 : node11580;
														assign node11580 = (inp[10]) ? node11588 : node11581;
															assign node11581 = (inp[12]) ? node11585 : node11582;
																assign node11582 = (inp[11]) ? 4'b0001 : 4'b0000;
																assign node11585 = (inp[11]) ? 4'b1000 : 4'b0000;
															assign node11588 = (inp[12]) ? node11592 : node11589;
																assign node11589 = (inp[11]) ? 4'b1000 : 4'b0000;
																assign node11592 = (inp[11]) ? 4'b0000 : 4'b1000;
														assign node11595 = (inp[12]) ? node11599 : node11596;
															assign node11596 = (inp[10]) ? 4'b0000 : 4'b0001;
															assign node11599 = (inp[11]) ? 4'b1000 : node11600;
																assign node11600 = (inp[10]) ? 4'b0001 : 4'b1001;
												assign node11604 = (inp[10]) ? node11626 : node11605;
													assign node11605 = (inp[14]) ? node11617 : node11606;
														assign node11606 = (inp[12]) ? node11612 : node11607;
															assign node11607 = (inp[11]) ? node11609 : 4'b0000;
																assign node11609 = (inp[7]) ? 4'b1000 : 4'b1001;
															assign node11612 = (inp[11]) ? 4'b0000 : node11613;
																assign node11613 = (inp[7]) ? 4'b1001 : 4'b1000;
														assign node11617 = (inp[11]) ? node11621 : node11618;
															assign node11618 = (inp[7]) ? 4'b1001 : 4'b0000;
															assign node11621 = (inp[7]) ? node11623 : 4'b1001;
																assign node11623 = (inp[12]) ? 4'b0000 : 4'b1000;
													assign node11626 = (inp[11]) ? node11636 : node11627;
														assign node11627 = (inp[14]) ? 4'b0001 : node11628;
															assign node11628 = (inp[7]) ? node11632 : node11629;
																assign node11629 = (inp[12]) ? 4'b0000 : 4'b1000;
																assign node11632 = (inp[12]) ? 4'b1001 : 4'b0001;
														assign node11636 = (inp[12]) ? 4'b0001 : 4'b0000;
											assign node11639 = (inp[11]) ? node11673 : node11640;
												assign node11640 = (inp[7]) ? node11656 : node11641;
													assign node11641 = (inp[14]) ? 4'b0001 : node11642;
														assign node11642 = (inp[12]) ? node11650 : node11643;
															assign node11643 = (inp[10]) ? node11647 : node11644;
																assign node11644 = (inp[2]) ? 4'b1000 : 4'b0001;
																assign node11647 = (inp[2]) ? 4'b0001 : 4'b1000;
															assign node11650 = (inp[2]) ? node11652 : 4'b0000;
																assign node11652 = (inp[10]) ? 4'b0001 : 4'b0000;
													assign node11656 = (inp[2]) ? node11666 : node11657;
														assign node11657 = (inp[14]) ? node11661 : node11658;
															assign node11658 = (inp[10]) ? 4'b0001 : 4'b0000;
															assign node11661 = (inp[10]) ? 4'b0000 : node11662;
																assign node11662 = (inp[12]) ? 4'b1000 : 4'b0001;
														assign node11666 = (inp[12]) ? 4'b0000 : node11667;
															assign node11667 = (inp[14]) ? node11669 : 4'b0000;
																assign node11669 = (inp[10]) ? 4'b1000 : 4'b0000;
												assign node11673 = (inp[10]) ? 4'b0001 : node11674;
													assign node11674 = (inp[12]) ? node11680 : node11675;
														assign node11675 = (inp[2]) ? 4'b0001 : node11676;
															assign node11676 = (inp[7]) ? 4'b0001 : 4'b1001;
														assign node11680 = (inp[7]) ? node11682 : 4'b0001;
															assign node11682 = (inp[2]) ? 4'b1001 : 4'b0001;
										assign node11686 = (inp[10]) ? node11720 : node11687;
											assign node11687 = (inp[11]) ? node11705 : node11688;
												assign node11688 = (inp[12]) ? 4'b0000 : node11689;
													assign node11689 = (inp[7]) ? node11697 : node11690;
														assign node11690 = (inp[1]) ? 4'b0000 : node11691;
															assign node11691 = (inp[2]) ? node11693 : 4'b0000;
																assign node11693 = (inp[14]) ? 4'b0001 : 4'b0000;
														assign node11697 = (inp[2]) ? node11699 : 4'b0001;
															assign node11699 = (inp[1]) ? 4'b0000 : node11700;
																assign node11700 = (inp[14]) ? 4'b0000 : 4'b0001;
												assign node11705 = (inp[1]) ? 4'b0001 : node11706;
													assign node11706 = (inp[14]) ? node11708 : 4'b0000;
														assign node11708 = (inp[12]) ? node11714 : node11709;
															assign node11709 = (inp[2]) ? node11711 : 4'b0000;
																assign node11711 = (inp[7]) ? 4'b0001 : 4'b0000;
															assign node11714 = (inp[7]) ? node11716 : 4'b0001;
																assign node11716 = (inp[2]) ? 4'b0000 : 4'b0001;
											assign node11720 = (inp[11]) ? 4'b0000 : node11721;
												assign node11721 = (inp[1]) ? 4'b0000 : node11722;
													assign node11722 = (inp[12]) ? node11734 : node11723;
														assign node11723 = (inp[7]) ? node11729 : node11724;
															assign node11724 = (inp[14]) ? 4'b0000 : node11725;
																assign node11725 = (inp[2]) ? 4'b0000 : 4'b0001;
															assign node11729 = (inp[14]) ? node11731 : 4'b0000;
																assign node11731 = (inp[2]) ? 4'b0001 : 4'b0000;
														assign node11734 = (inp[7]) ? node11738 : node11735;
															assign node11735 = (inp[2]) ? 4'b0001 : 4'b0000;
															assign node11738 = (inp[2]) ? node11740 : 4'b0001;
																assign node11740 = (inp[14]) ? 4'b0000 : 4'b0001;
					assign node11745 = (inp[6]) ? node11747 : 4'b0001;
						assign node11747 = (inp[2]) ? node12259 : node11748;
							assign node11748 = (inp[5]) ? node11850 : node11749;
								assign node11749 = (inp[3]) ? node11751 : 4'b0001;
									assign node11751 = (inp[7]) ? node11825 : node11752;
										assign node11752 = (inp[4]) ? node11766 : node11753;
											assign node11753 = (inp[13]) ? node11755 : 4'b0001;
												assign node11755 = (inp[1]) ? node11759 : node11756;
													assign node11756 = (inp[14]) ? 4'b0001 : 4'b0000;
													assign node11759 = (inp[14]) ? node11761 : 4'b0001;
														assign node11761 = (inp[11]) ? 4'b0001 : node11762;
															assign node11762 = (inp[12]) ? 4'b0001 : 4'b0000;
											assign node11766 = (inp[1]) ? node11796 : node11767;
												assign node11767 = (inp[11]) ? node11787 : node11768;
													assign node11768 = (inp[14]) ? node11776 : node11769;
														assign node11769 = (inp[13]) ? node11773 : node11770;
															assign node11770 = (inp[10]) ? 4'b1000 : 4'b0000;
															assign node11773 = (inp[12]) ? 4'b1000 : 4'b0000;
														assign node11776 = (inp[13]) ? node11782 : node11777;
															assign node11777 = (inp[10]) ? node11779 : 4'b0001;
																assign node11779 = (inp[12]) ? 4'b0001 : 4'b1001;
															assign node11782 = (inp[10]) ? node11784 : 4'b1001;
																assign node11784 = (inp[12]) ? 4'b1001 : 4'b0001;
													assign node11787 = (inp[13]) ? node11793 : node11788;
														assign node11788 = (inp[12]) ? node11790 : 4'b1000;
															assign node11790 = (inp[10]) ? 4'b1000 : 4'b0000;
														assign node11793 = (inp[12]) ? 4'b1000 : 4'b0000;
												assign node11796 = (inp[11]) ? node11814 : node11797;
													assign node11797 = (inp[14]) ? node11807 : node11798;
														assign node11798 = (inp[12]) ? node11800 : 4'b0001;
															assign node11800 = (inp[10]) ? node11804 : node11801;
																assign node11801 = (inp[13]) ? 4'b1001 : 4'b0001;
																assign node11804 = (inp[13]) ? 4'b0001 : 4'b1001;
														assign node11807 = (inp[13]) ? node11809 : 4'b1000;
															assign node11809 = (inp[12]) ? node11811 : 4'b0000;
																assign node11811 = (inp[10]) ? 4'b0000 : 4'b1000;
													assign node11814 = (inp[13]) ? node11820 : node11815;
														assign node11815 = (inp[12]) ? node11817 : 4'b1001;
															assign node11817 = (inp[10]) ? 4'b1001 : 4'b0001;
														assign node11820 = (inp[12]) ? node11822 : 4'b0001;
															assign node11822 = (inp[10]) ? 4'b0001 : 4'b1001;
										assign node11825 = (inp[4]) ? node11827 : 4'b0001;
											assign node11827 = (inp[13]) ? node11829 : 4'b0001;
												assign node11829 = (inp[1]) ? node11841 : node11830;
													assign node11830 = (inp[10]) ? node11836 : node11831;
														assign node11831 = (inp[11]) ? node11833 : 4'b0001;
															assign node11833 = (inp[12]) ? 4'b0001 : 4'b0000;
														assign node11836 = (inp[14]) ? node11838 : 4'b0000;
															assign node11838 = (inp[11]) ? 4'b0000 : 4'b0001;
													assign node11841 = (inp[14]) ? node11843 : 4'b0001;
														assign node11843 = (inp[11]) ? 4'b0001 : node11844;
															assign node11844 = (inp[10]) ? 4'b0000 : node11845;
																assign node11845 = (inp[12]) ? 4'b0001 : 4'b0000;
								assign node11850 = (inp[13]) ? node12066 : node11851;
									assign node11851 = (inp[11]) ? node11975 : node11852;
										assign node11852 = (inp[12]) ? node11908 : node11853;
											assign node11853 = (inp[3]) ? node11877 : node11854;
												assign node11854 = (inp[7]) ? node11868 : node11855;
													assign node11855 = (inp[10]) ? node11863 : node11856;
														assign node11856 = (inp[14]) ? node11860 : node11857;
															assign node11857 = (inp[1]) ? 4'b1101 : 4'b1100;
															assign node11860 = (inp[1]) ? 4'b1000 : 4'b0001;
														assign node11863 = (inp[4]) ? 4'b0000 : node11864;
															assign node11864 = (inp[1]) ? 4'b1001 : 4'b1000;
													assign node11868 = (inp[14]) ? node11872 : node11869;
														assign node11869 = (inp[1]) ? 4'b1001 : 4'b1000;
														assign node11872 = (inp[1]) ? 4'b1000 : node11873;
															assign node11873 = (inp[10]) ? 4'b1001 : 4'b0001;
												assign node11877 = (inp[4]) ? node11889 : node11878;
													assign node11878 = (inp[10]) ? node11884 : node11879;
														assign node11879 = (inp[14]) ? 4'b1000 : node11880;
															assign node11880 = (inp[7]) ? 4'b1000 : 4'b0000;
														assign node11884 = (inp[7]) ? 4'b0000 : node11885;
															assign node11885 = (inp[14]) ? 4'b1001 : 4'b1000;
													assign node11889 = (inp[14]) ? node11901 : node11890;
														assign node11890 = (inp[10]) ? node11894 : node11891;
															assign node11891 = (inp[1]) ? 4'b0001 : 4'b1001;
															assign node11894 = (inp[7]) ? node11898 : node11895;
																assign node11895 = (inp[1]) ? 4'b0001 : 4'b1001;
																assign node11898 = (inp[1]) ? 4'b1000 : 4'b0000;
														assign node11901 = (inp[10]) ? 4'b0000 : node11902;
															assign node11902 = (inp[7]) ? 4'b0000 : node11903;
																assign node11903 = (inp[1]) ? 4'b1000 : 4'b1001;
											assign node11908 = (inp[4]) ? node11940 : node11909;
												assign node11909 = (inp[3]) ? node11925 : node11910;
													assign node11910 = (inp[10]) ? node11918 : node11911;
														assign node11911 = (inp[14]) ? node11915 : node11912;
															assign node11912 = (inp[1]) ? 4'b0001 : 4'b0000;
															assign node11915 = (inp[1]) ? 4'b0000 : 4'b0001;
														assign node11918 = (inp[1]) ? node11922 : node11919;
															assign node11919 = (inp[14]) ? 4'b0001 : 4'b1000;
															assign node11922 = (inp[14]) ? 4'b1000 : 4'b1001;
													assign node11925 = (inp[1]) ? node11931 : node11926;
														assign node11926 = (inp[10]) ? node11928 : 4'b0000;
															assign node11928 = (inp[7]) ? 4'b1000 : 4'b0001;
														assign node11931 = (inp[10]) ? node11933 : 4'b1000;
															assign node11933 = (inp[14]) ? node11937 : node11934;
																assign node11934 = (inp[7]) ? 4'b0000 : 4'b1000;
																assign node11937 = (inp[7]) ? 4'b0000 : 4'b0001;
												assign node11940 = (inp[7]) ? node11954 : node11941;
													assign node11941 = (inp[3]) ? node11949 : node11942;
														assign node11942 = (inp[1]) ? node11944 : 4'b0101;
															assign node11944 = (inp[10]) ? 4'b0000 : node11945;
																assign node11945 = (inp[14]) ? 4'b0100 : 4'b0101;
														assign node11949 = (inp[10]) ? 4'b0001 : node11950;
															assign node11950 = (inp[1]) ? 4'b0000 : 4'b0001;
													assign node11954 = (inp[3]) ? node11966 : node11955;
														assign node11955 = (inp[10]) ? node11959 : node11956;
															assign node11956 = (inp[1]) ? 4'b0001 : 4'b0000;
															assign node11959 = (inp[1]) ? node11963 : node11960;
																assign node11960 = (inp[14]) ? 4'b0001 : 4'b1000;
																assign node11963 = (inp[14]) ? 4'b1000 : 4'b1001;
														assign node11966 = (inp[10]) ? node11972 : node11967;
															assign node11967 = (inp[14]) ? node11969 : 4'b0001;
																assign node11969 = (inp[1]) ? 4'b0000 : 4'b0001;
															assign node11972 = (inp[1]) ? 4'b0001 : 4'b0000;
										assign node11975 = (inp[1]) ? node12019 : node11976;
											assign node11976 = (inp[3]) ? node11996 : node11977;
												assign node11977 = (inp[12]) ? node11985 : node11978;
													assign node11978 = (inp[4]) ? node11980 : 4'b1000;
														assign node11980 = (inp[10]) ? node11982 : 4'b1100;
															assign node11982 = (inp[7]) ? 4'b1000 : 4'b0001;
													assign node11985 = (inp[10]) ? node11991 : node11986;
														assign node11986 = (inp[4]) ? node11988 : 4'b0000;
															assign node11988 = (inp[7]) ? 4'b0000 : 4'b0100;
														assign node11991 = (inp[4]) ? node11993 : 4'b1000;
															assign node11993 = (inp[7]) ? 4'b1000 : 4'b1100;
												assign node11996 = (inp[4]) ? node12008 : node11997;
													assign node11997 = (inp[12]) ? node12001 : node11998;
														assign node11998 = (inp[10]) ? 4'b1000 : 4'b1001;
														assign node12001 = (inp[7]) ? node12005 : node12002;
															assign node12002 = (inp[10]) ? 4'b0000 : 4'b0001;
															assign node12005 = (inp[10]) ? 4'b1001 : 4'b0001;
													assign node12008 = (inp[10]) ? node12014 : node12009;
														assign node12009 = (inp[12]) ? node12011 : 4'b0001;
															assign node12011 = (inp[7]) ? 4'b1001 : 4'b1000;
														assign node12014 = (inp[7]) ? node12016 : 4'b0001;
															assign node12016 = (inp[12]) ? 4'b0001 : 4'b0000;
											assign node12019 = (inp[3]) ? node12039 : node12020;
												assign node12020 = (inp[12]) ? node12032 : node12021;
													assign node12021 = (inp[10]) ? node12027 : node12022;
														assign node12022 = (inp[4]) ? node12024 : 4'b1001;
															assign node12024 = (inp[7]) ? 4'b1001 : 4'b1101;
														assign node12027 = (inp[7]) ? 4'b1001 : node12028;
															assign node12028 = (inp[4]) ? 4'b0001 : 4'b1001;
													assign node12032 = (inp[10]) ? 4'b1001 : node12033;
														assign node12033 = (inp[4]) ? node12035 : 4'b0001;
															assign node12035 = (inp[7]) ? 4'b0001 : 4'b0101;
												assign node12039 = (inp[4]) ? node12055 : node12040;
													assign node12040 = (inp[14]) ? node12048 : node12041;
														assign node12041 = (inp[7]) ? node12045 : node12042;
															assign node12042 = (inp[10]) ? 4'b1001 : 4'b0001;
															assign node12045 = (inp[10]) ? 4'b0001 : 4'b1001;
														assign node12048 = (inp[12]) ? 4'b1001 : node12049;
															assign node12049 = (inp[7]) ? node12051 : 4'b1001;
																assign node12051 = (inp[10]) ? 4'b0001 : 4'b1001;
													assign node12055 = (inp[10]) ? 4'b0001 : node12056;
														assign node12056 = (inp[14]) ? node12060 : node12057;
															assign node12057 = (inp[7]) ? 4'b0001 : 4'b1001;
															assign node12060 = (inp[12]) ? 4'b0001 : node12061;
																assign node12061 = (inp[7]) ? 4'b1001 : 4'b0001;
									assign node12066 = (inp[3]) ? node12178 : node12067;
										assign node12067 = (inp[10]) ? node12127 : node12068;
											assign node12068 = (inp[12]) ? node12108 : node12069;
												assign node12069 = (inp[1]) ? node12087 : node12070;
													assign node12070 = (inp[14]) ? node12076 : node12071;
														assign node12071 = (inp[4]) ? node12073 : 4'b0100;
															assign node12073 = (inp[7]) ? 4'b0100 : 4'b1001;
														assign node12076 = (inp[11]) ? node12082 : node12077;
															assign node12077 = (inp[7]) ? 4'b1001 : node12078;
																assign node12078 = (inp[4]) ? 4'b1000 : 4'b1001;
															assign node12082 = (inp[7]) ? node12084 : 4'b1001;
																assign node12084 = (inp[4]) ? 4'b0100 : 4'b0000;
													assign node12087 = (inp[11]) ? node12101 : node12088;
														assign node12088 = (inp[14]) ? node12096 : node12089;
															assign node12089 = (inp[7]) ? node12093 : node12090;
																assign node12090 = (inp[4]) ? 4'b1000 : 4'b0101;
																assign node12093 = (inp[4]) ? 4'b0101 : 4'b0001;
															assign node12096 = (inp[7]) ? node12098 : 4'b0100;
																assign node12098 = (inp[4]) ? 4'b0100 : 4'b0000;
														assign node12101 = (inp[4]) ? node12105 : node12102;
															assign node12102 = (inp[7]) ? 4'b0001 : 4'b0101;
															assign node12105 = (inp[7]) ? 4'b0101 : 4'b1001;
												assign node12108 = (inp[4]) ? node12120 : node12109;
													assign node12109 = (inp[1]) ? node12115 : node12110;
														assign node12110 = (inp[14]) ? node12112 : 4'b1000;
															assign node12112 = (inp[11]) ? 4'b1000 : 4'b1001;
														assign node12115 = (inp[11]) ? 4'b1001 : node12116;
															assign node12116 = (inp[14]) ? 4'b1000 : 4'b1001;
													assign node12120 = (inp[1]) ? 4'b1000 : node12121;
														assign node12121 = (inp[7]) ? 4'b1000 : node12122;
															assign node12122 = (inp[11]) ? 4'b0001 : 4'b0000;
											assign node12127 = (inp[7]) ? node12151 : node12128;
												assign node12128 = (inp[4]) ? node12140 : node12129;
													assign node12129 = (inp[1]) ? node12135 : node12130;
														assign node12130 = (inp[14]) ? node12132 : 4'b0100;
															assign node12132 = (inp[11]) ? 4'b0100 : 4'b0101;
														assign node12135 = (inp[14]) ? node12137 : 4'b0101;
															assign node12137 = (inp[11]) ? 4'b0101 : 4'b0100;
													assign node12140 = (inp[11]) ? node12146 : node12141;
														assign node12141 = (inp[1]) ? 4'b0000 : node12142;
															assign node12142 = (inp[12]) ? 4'b1000 : 4'b0000;
														assign node12146 = (inp[12]) ? node12148 : 4'b0001;
															assign node12148 = (inp[1]) ? 4'b0001 : 4'b1001;
												assign node12151 = (inp[1]) ? node12171 : node12152;
													assign node12152 = (inp[14]) ? node12160 : node12153;
														assign node12153 = (inp[4]) ? node12155 : 4'b0000;
															assign node12155 = (inp[11]) ? 4'b0001 : node12156;
																assign node12156 = (inp[12]) ? 4'b0100 : 4'b0000;
														assign node12160 = (inp[12]) ? node12168 : node12161;
															assign node12161 = (inp[4]) ? node12165 : node12162;
																assign node12162 = (inp[11]) ? 4'b0000 : 4'b0001;
																assign node12165 = (inp[11]) ? 4'b0001 : 4'b0000;
															assign node12168 = (inp[11]) ? 4'b0100 : 4'b1001;
													assign node12171 = (inp[11]) ? 4'b0001 : node12172;
														assign node12172 = (inp[12]) ? 4'b0000 : node12173;
															assign node12173 = (inp[14]) ? 4'b0000 : 4'b0001;
										assign node12178 = (inp[4]) ? node12226 : node12179;
											assign node12179 = (inp[10]) ? node12201 : node12180;
												assign node12180 = (inp[1]) ? node12188 : node12181;
													assign node12181 = (inp[7]) ? 4'b0000 : node12182;
														assign node12182 = (inp[11]) ? 4'b0000 : node12183;
															assign node12183 = (inp[12]) ? 4'b1001 : 4'b0000;
													assign node12188 = (inp[14]) ? node12196 : node12189;
														assign node12189 = (inp[11]) ? 4'b0001 : node12190;
															assign node12190 = (inp[12]) ? 4'b0000 : node12191;
																assign node12191 = (inp[7]) ? 4'b1000 : 4'b0001;
														assign node12196 = (inp[11]) ? node12198 : 4'b0001;
															assign node12198 = (inp[12]) ? 4'b0001 : 4'b1001;
												assign node12201 = (inp[1]) ? node12213 : node12202;
													assign node12202 = (inp[7]) ? node12208 : node12203;
														assign node12203 = (inp[11]) ? 4'b1001 : node12204;
															assign node12204 = (inp[12]) ? 4'b0001 : 4'b1001;
														assign node12208 = (inp[14]) ? 4'b1000 : node12209;
															assign node12209 = (inp[11]) ? 4'b0000 : 4'b1001;
													assign node12213 = (inp[11]) ? 4'b0001 : node12214;
														assign node12214 = (inp[12]) ? node12220 : node12215;
															assign node12215 = (inp[7]) ? 4'b0001 : node12216;
																assign node12216 = (inp[14]) ? 4'b0000 : 4'b0001;
															assign node12220 = (inp[14]) ? 4'b1001 : node12221;
																assign node12221 = (inp[7]) ? 4'b0000 : 4'b1001;
											assign node12226 = (inp[10]) ? node12246 : node12227;
												assign node12227 = (inp[7]) ? node12233 : node12228;
													assign node12228 = (inp[1]) ? 4'b0001 : node12229;
														assign node12229 = (inp[12]) ? 4'b0000 : 4'b0001;
													assign node12233 = (inp[12]) ? node12235 : 4'b0000;
														assign node12235 = (inp[1]) ? node12241 : node12236;
															assign node12236 = (inp[11]) ? 4'b0000 : node12237;
																assign node12237 = (inp[14]) ? 4'b0001 : 4'b0000;
															assign node12241 = (inp[11]) ? 4'b0001 : node12242;
																assign node12242 = (inp[14]) ? 4'b0000 : 4'b0001;
												assign node12246 = (inp[14]) ? 4'b0000 : node12247;
													assign node12247 = (inp[11]) ? 4'b0000 : node12248;
														assign node12248 = (inp[1]) ? 4'b0000 : node12249;
															assign node12249 = (inp[12]) ? node12253 : node12250;
																assign node12250 = (inp[7]) ? 4'b0001 : 4'b0000;
																assign node12253 = (inp[7]) ? 4'b0000 : 4'b0001;
							assign node12259 = (inp[3]) ? node12261 : 4'b0001;
								assign node12261 = (inp[5]) ? node12263 : 4'b0001;
									assign node12263 = (inp[4]) ? node12287 : node12264;
										assign node12264 = (inp[13]) ? node12266 : 4'b0001;
											assign node12266 = (inp[7]) ? 4'b0001 : node12267;
												assign node12267 = (inp[1]) ? node12279 : node12268;
													assign node12268 = (inp[14]) ? node12274 : node12269;
														assign node12269 = (inp[10]) ? 4'b0000 : node12270;
															assign node12270 = (inp[12]) ? 4'b0001 : 4'b0000;
														assign node12274 = (inp[11]) ? node12276 : 4'b0001;
															assign node12276 = (inp[12]) ? 4'b0001 : 4'b0000;
													assign node12279 = (inp[11]) ? 4'b0001 : node12280;
														assign node12280 = (inp[10]) ? node12282 : 4'b0001;
															assign node12282 = (inp[14]) ? 4'b0000 : 4'b0001;
										assign node12287 = (inp[7]) ? node12337 : node12288;
											assign node12288 = (inp[1]) ? node12314 : node12289;
												assign node12289 = (inp[13]) ? node12307 : node12290;
													assign node12290 = (inp[14]) ? node12300 : node12291;
														assign node12291 = (inp[11]) ? node12297 : node12292;
															assign node12292 = (inp[12]) ? 4'b1000 : node12293;
																assign node12293 = (inp[10]) ? 4'b0000 : 4'b1000;
															assign node12297 = (inp[10]) ? 4'b1000 : 4'b0000;
														assign node12300 = (inp[11]) ? node12304 : node12301;
															assign node12301 = (inp[10]) ? 4'b0000 : 4'b0001;
															assign node12304 = (inp[12]) ? 4'b0000 : 4'b0001;
													assign node12307 = (inp[11]) ? 4'b0000 : node12308;
														assign node12308 = (inp[14]) ? 4'b0000 : node12309;
															assign node12309 = (inp[12]) ? 4'b0000 : 4'b0001;
												assign node12314 = (inp[11]) ? node12324 : node12315;
													assign node12315 = (inp[10]) ? 4'b0000 : node12316;
														assign node12316 = (inp[13]) ? node12320 : node12317;
															assign node12317 = (inp[12]) ? 4'b0000 : 4'b1000;
															assign node12320 = (inp[12]) ? 4'b0000 : 4'b0001;
													assign node12324 = (inp[14]) ? node12330 : node12325;
														assign node12325 = (inp[12]) ? 4'b0001 : node12326;
															assign node12326 = (inp[10]) ? 4'b0001 : 4'b1001;
														assign node12330 = (inp[12]) ? 4'b0001 : node12331;
															assign node12331 = (inp[10]) ? node12333 : 4'b0001;
																assign node12333 = (inp[13]) ? 4'b0000 : 4'b0001;
											assign node12337 = (inp[13]) ? node12339 : 4'b0001;
												assign node12339 = (inp[10]) ? node12347 : node12340;
													assign node12340 = (inp[12]) ? 4'b0001 : node12341;
														assign node12341 = (inp[1]) ? node12343 : 4'b0000;
															assign node12343 = (inp[11]) ? 4'b0001 : 4'b0000;
													assign node12347 = (inp[12]) ? node12349 : 4'b0000;
														assign node12349 = (inp[14]) ? node12351 : 4'b0000;
															assign node12351 = (inp[11]) ? 4'b0000 : 4'b0001;
		assign node12354 = (inp[9]) ? node18598 : node12355;
			assign node12355 = (inp[15]) ? node15743 : node12356;
				assign node12356 = (inp[6]) ? node13104 : node12357;
					assign node12357 = (inp[0]) ? 4'b1100 : node12358;
						assign node12358 = (inp[2]) ? node12802 : node12359;
							assign node12359 = (inp[1]) ? node12571 : node12360;
								assign node12360 = (inp[13]) ? node12466 : node12361;
									assign node12361 = (inp[10]) ? node12407 : node12362;
										assign node12362 = (inp[3]) ? node12390 : node12363;
											assign node12363 = (inp[5]) ? node12373 : node12364;
												assign node12364 = (inp[7]) ? 4'b1110 : node12365;
													assign node12365 = (inp[4]) ? node12367 : 4'b1110;
														assign node12367 = (inp[14]) ? node12369 : 4'b1001;
															assign node12369 = (inp[11]) ? 4'b1001 : 4'b1000;
												assign node12373 = (inp[14]) ? node12379 : node12374;
													assign node12374 = (inp[7]) ? 4'b1101 : node12375;
														assign node12375 = (inp[4]) ? 4'b1001 : 4'b1101;
													assign node12379 = (inp[11]) ? node12385 : node12380;
														assign node12380 = (inp[7]) ? 4'b1100 : node12381;
															assign node12381 = (inp[4]) ? 4'b1000 : 4'b1100;
														assign node12385 = (inp[4]) ? node12387 : 4'b1101;
															assign node12387 = (inp[7]) ? 4'b1101 : 4'b1001;
											assign node12390 = (inp[14]) ? node12396 : node12391;
												assign node12391 = (inp[4]) ? node12393 : 4'b1001;
													assign node12393 = (inp[7]) ? 4'b1001 : 4'b1101;
												assign node12396 = (inp[11]) ? node12402 : node12397;
													assign node12397 = (inp[7]) ? 4'b1000 : node12398;
														assign node12398 = (inp[4]) ? 4'b1100 : 4'b1000;
													assign node12402 = (inp[7]) ? 4'b1001 : node12403;
														assign node12403 = (inp[4]) ? 4'b1101 : 4'b1001;
										assign node12407 = (inp[12]) ? node12437 : node12408;
											assign node12408 = (inp[14]) ? node12420 : node12409;
												assign node12409 = (inp[3]) ? node12415 : node12410;
													assign node12410 = (inp[7]) ? node12412 : 4'b0001;
														assign node12412 = (inp[5]) ? 4'b0101 : 4'b0001;
													assign node12415 = (inp[4]) ? 4'b0101 : node12416;
														assign node12416 = (inp[7]) ? 4'b0001 : 4'b0101;
												assign node12420 = (inp[11]) ? node12428 : node12421;
													assign node12421 = (inp[3]) ? node12423 : 4'b0000;
														assign node12423 = (inp[7]) ? node12425 : 4'b0100;
															assign node12425 = (inp[4]) ? 4'b0100 : 4'b0000;
													assign node12428 = (inp[3]) ? node12432 : node12429;
														assign node12429 = (inp[4]) ? 4'b0001 : 4'b1110;
														assign node12432 = (inp[4]) ? 4'b0101 : node12433;
															assign node12433 = (inp[7]) ? 4'b0001 : 4'b0101;
											assign node12437 = (inp[3]) ? node12457 : node12438;
												assign node12438 = (inp[5]) ? node12446 : node12439;
													assign node12439 = (inp[4]) ? node12441 : 4'b1110;
														assign node12441 = (inp[7]) ? 4'b1110 : node12442;
															assign node12442 = (inp[11]) ? 4'b1001 : 4'b1000;
													assign node12446 = (inp[4]) ? node12448 : 4'b1101;
														assign node12448 = (inp[7]) ? node12454 : node12449;
															assign node12449 = (inp[14]) ? node12451 : 4'b1001;
																assign node12451 = (inp[11]) ? 4'b1001 : 4'b1000;
															assign node12454 = (inp[14]) ? 4'b1100 : 4'b1101;
												assign node12457 = (inp[11]) ? node12461 : node12458;
													assign node12458 = (inp[14]) ? 4'b1000 : 4'b1001;
													assign node12461 = (inp[4]) ? node12463 : 4'b1001;
														assign node12463 = (inp[7]) ? 4'b1001 : 4'b1101;
									assign node12466 = (inp[3]) ? node12518 : node12467;
										assign node12467 = (inp[4]) ? node12501 : node12468;
											assign node12468 = (inp[7]) ? node12486 : node12469;
												assign node12469 = (inp[14]) ? node12475 : node12470;
													assign node12470 = (inp[12]) ? 4'b0001 : node12471;
														assign node12471 = (inp[10]) ? 4'b1001 : 4'b0001;
													assign node12475 = (inp[11]) ? node12481 : node12476;
														assign node12476 = (inp[10]) ? node12478 : 4'b0000;
															assign node12478 = (inp[12]) ? 4'b0000 : 4'b1000;
														assign node12481 = (inp[12]) ? 4'b0001 : node12482;
															assign node12482 = (inp[10]) ? 4'b1001 : 4'b0001;
												assign node12486 = (inp[5]) ? node12488 : 4'b1110;
													assign node12488 = (inp[12]) ? node12496 : node12489;
														assign node12489 = (inp[10]) ? node12491 : 4'b0101;
															assign node12491 = (inp[14]) ? node12493 : 4'b1101;
																assign node12493 = (inp[11]) ? 4'b1101 : 4'b1100;
														assign node12496 = (inp[11]) ? 4'b0101 : node12497;
															assign node12497 = (inp[14]) ? 4'b0100 : 4'b0101;
											assign node12501 = (inp[14]) ? node12507 : node12502;
												assign node12502 = (inp[12]) ? 4'b0001 : node12503;
													assign node12503 = (inp[10]) ? 4'b1001 : 4'b0001;
												assign node12507 = (inp[11]) ? node12513 : node12508;
													assign node12508 = (inp[10]) ? node12510 : 4'b0000;
														assign node12510 = (inp[12]) ? 4'b0000 : 4'b1000;
													assign node12513 = (inp[10]) ? node12515 : 4'b0001;
														assign node12515 = (inp[12]) ? 4'b0001 : 4'b1001;
										assign node12518 = (inp[12]) ? node12554 : node12519;
											assign node12519 = (inp[10]) ? node12537 : node12520;
												assign node12520 = (inp[14]) ? node12526 : node12521;
													assign node12521 = (inp[4]) ? 4'b0101 : node12522;
														assign node12522 = (inp[7]) ? 4'b0001 : 4'b0101;
													assign node12526 = (inp[11]) ? node12532 : node12527;
														assign node12527 = (inp[7]) ? node12529 : 4'b0100;
															assign node12529 = (inp[4]) ? 4'b0100 : 4'b0000;
														assign node12532 = (inp[4]) ? 4'b0101 : node12533;
															assign node12533 = (inp[7]) ? 4'b0001 : 4'b0101;
												assign node12537 = (inp[14]) ? node12543 : node12538;
													assign node12538 = (inp[4]) ? 4'b1101 : node12539;
														assign node12539 = (inp[7]) ? 4'b1001 : 4'b1101;
													assign node12543 = (inp[11]) ? node12549 : node12544;
														assign node12544 = (inp[4]) ? 4'b1100 : node12545;
															assign node12545 = (inp[7]) ? 4'b1000 : 4'b1100;
														assign node12549 = (inp[4]) ? 4'b1101 : node12550;
															assign node12550 = (inp[7]) ? 4'b1001 : 4'b1101;
											assign node12554 = (inp[11]) ? node12566 : node12555;
												assign node12555 = (inp[14]) ? node12561 : node12556;
													assign node12556 = (inp[7]) ? node12558 : 4'b0101;
														assign node12558 = (inp[4]) ? 4'b0101 : 4'b0001;
													assign node12561 = (inp[4]) ? 4'b0100 : node12562;
														assign node12562 = (inp[7]) ? 4'b0000 : 4'b0100;
												assign node12566 = (inp[7]) ? node12568 : 4'b0101;
													assign node12568 = (inp[4]) ? 4'b0101 : 4'b0001;
								assign node12571 = (inp[14]) ? node12655 : node12572;
									assign node12572 = (inp[13]) ? node12616 : node12573;
										assign node12573 = (inp[12]) ? node12587 : node12574;
											assign node12574 = (inp[3]) ? node12582 : node12575;
												assign node12575 = (inp[7]) ? node12577 : 4'b0000;
													assign node12577 = (inp[4]) ? 4'b0000 : node12578;
														assign node12578 = (inp[5]) ? 4'b0100 : 4'b1110;
												assign node12582 = (inp[7]) ? node12584 : 4'b0100;
													assign node12584 = (inp[4]) ? 4'b0100 : 4'b0000;
											assign node12587 = (inp[10]) ? node12603 : node12588;
												assign node12588 = (inp[3]) ? node12598 : node12589;
													assign node12589 = (inp[7]) ? node12595 : node12590;
														assign node12590 = (inp[4]) ? 4'b1000 : node12591;
															assign node12591 = (inp[5]) ? 4'b1100 : 4'b1110;
														assign node12595 = (inp[5]) ? 4'b1100 : 4'b1110;
													assign node12598 = (inp[7]) ? 4'b1000 : node12599;
														assign node12599 = (inp[4]) ? 4'b1100 : 4'b1000;
												assign node12603 = (inp[3]) ? node12611 : node12604;
													assign node12604 = (inp[7]) ? node12606 : 4'b0000;
														assign node12606 = (inp[4]) ? 4'b0000 : node12607;
															assign node12607 = (inp[5]) ? 4'b0100 : 4'b1110;
													assign node12611 = (inp[7]) ? node12613 : 4'b0100;
														assign node12613 = (inp[4]) ? 4'b0100 : 4'b0000;
										assign node12616 = (inp[10]) ? node12642 : node12617;
											assign node12617 = (inp[12]) ? node12629 : node12618;
												assign node12618 = (inp[3]) ? node12624 : node12619;
													assign node12619 = (inp[7]) ? node12621 : 4'b1000;
														assign node12621 = (inp[4]) ? 4'b1000 : 4'b1100;
													assign node12624 = (inp[7]) ? node12626 : 4'b1100;
														assign node12626 = (inp[4]) ? 4'b1100 : 4'b1000;
												assign node12629 = (inp[3]) ? node12637 : node12630;
													assign node12630 = (inp[7]) ? node12632 : 4'b0000;
														assign node12632 = (inp[4]) ? 4'b0000 : node12633;
															assign node12633 = (inp[5]) ? 4'b0100 : 4'b1110;
													assign node12637 = (inp[4]) ? 4'b0100 : node12638;
														assign node12638 = (inp[7]) ? 4'b0000 : 4'b0100;
											assign node12642 = (inp[3]) ? node12650 : node12643;
												assign node12643 = (inp[7]) ? node12645 : 4'b1000;
													assign node12645 = (inp[4]) ? 4'b1000 : node12646;
														assign node12646 = (inp[5]) ? 4'b1100 : 4'b1110;
												assign node12650 = (inp[7]) ? node12652 : 4'b1100;
													assign node12652 = (inp[4]) ? 4'b1100 : 4'b1000;
									assign node12655 = (inp[11]) ? node12725 : node12656;
										assign node12656 = (inp[13]) ? node12690 : node12657;
											assign node12657 = (inp[3]) ? node12673 : node12658;
												assign node12658 = (inp[4]) ? node12664 : node12659;
													assign node12659 = (inp[5]) ? node12661 : 4'b1110;
														assign node12661 = (inp[12]) ? 4'b1101 : 4'b0101;
													assign node12664 = (inp[12]) ? node12668 : node12665;
														assign node12665 = (inp[10]) ? 4'b0001 : 4'b1001;
														assign node12668 = (inp[7]) ? node12670 : 4'b1001;
															assign node12670 = (inp[5]) ? 4'b1101 : 4'b1110;
												assign node12673 = (inp[12]) ? node12685 : node12674;
													assign node12674 = (inp[10]) ? node12680 : node12675;
														assign node12675 = (inp[7]) ? 4'b1001 : node12676;
															assign node12676 = (inp[4]) ? 4'b1101 : 4'b1001;
														assign node12680 = (inp[7]) ? node12682 : 4'b0101;
															assign node12682 = (inp[5]) ? 4'b0001 : 4'b0101;
													assign node12685 = (inp[7]) ? 4'b1001 : node12686;
														assign node12686 = (inp[4]) ? 4'b1101 : 4'b1001;
											assign node12690 = (inp[12]) ? node12712 : node12691;
												assign node12691 = (inp[10]) ? node12701 : node12692;
													assign node12692 = (inp[3]) ? node12698 : node12693;
														assign node12693 = (inp[7]) ? node12695 : 4'b0001;
															assign node12695 = (inp[5]) ? 4'b0101 : 4'b1110;
														assign node12698 = (inp[7]) ? 4'b0001 : 4'b0101;
													assign node12701 = (inp[3]) ? node12707 : node12702;
														assign node12702 = (inp[7]) ? node12704 : 4'b1001;
															assign node12704 = (inp[5]) ? 4'b1101 : 4'b1110;
														assign node12707 = (inp[7]) ? node12709 : 4'b1101;
															assign node12709 = (inp[4]) ? 4'b1101 : 4'b1001;
												assign node12712 = (inp[3]) ? node12720 : node12713;
													assign node12713 = (inp[7]) ? node12715 : 4'b0001;
														assign node12715 = (inp[5]) ? node12717 : 4'b1110;
															assign node12717 = (inp[4]) ? 4'b0001 : 4'b0101;
													assign node12720 = (inp[7]) ? node12722 : 4'b0101;
														assign node12722 = (inp[4]) ? 4'b0101 : 4'b0001;
										assign node12725 = (inp[3]) ? node12765 : node12726;
											assign node12726 = (inp[7]) ? node12742 : node12727;
												assign node12727 = (inp[13]) ? node12737 : node12728;
													assign node12728 = (inp[12]) ? node12730 : 4'b0000;
														assign node12730 = (inp[10]) ? 4'b0000 : node12731;
															assign node12731 = (inp[4]) ? 4'b1000 : node12732;
																assign node12732 = (inp[5]) ? 4'b1100 : 4'b1110;
													assign node12737 = (inp[12]) ? node12739 : 4'b1000;
														assign node12739 = (inp[10]) ? 4'b1000 : 4'b0000;
												assign node12742 = (inp[4]) ? node12754 : node12743;
													assign node12743 = (inp[5]) ? node12745 : 4'b1110;
														assign node12745 = (inp[12]) ? node12747 : 4'b0100;
															assign node12747 = (inp[10]) ? node12751 : node12748;
																assign node12748 = (inp[13]) ? 4'b0100 : 4'b1100;
																assign node12751 = (inp[13]) ? 4'b1100 : 4'b0100;
													assign node12754 = (inp[13]) ? node12762 : node12755;
														assign node12755 = (inp[12]) ? node12757 : 4'b0000;
															assign node12757 = (inp[10]) ? 4'b0000 : node12758;
																assign node12758 = (inp[5]) ? 4'b1100 : 4'b1110;
														assign node12762 = (inp[10]) ? 4'b1000 : 4'b0000;
											assign node12765 = (inp[4]) ? node12787 : node12766;
												assign node12766 = (inp[7]) ? node12776 : node12767;
													assign node12767 = (inp[13]) ? node12773 : node12768;
														assign node12768 = (inp[12]) ? node12770 : 4'b0100;
															assign node12770 = (inp[10]) ? 4'b0100 : 4'b1000;
														assign node12773 = (inp[12]) ? 4'b0100 : 4'b1100;
													assign node12776 = (inp[13]) ? node12782 : node12777;
														assign node12777 = (inp[10]) ? 4'b0000 : node12778;
															assign node12778 = (inp[12]) ? 4'b1000 : 4'b0000;
														assign node12782 = (inp[5]) ? 4'b1000 : node12783;
															assign node12783 = (inp[12]) ? 4'b0000 : 4'b1000;
												assign node12787 = (inp[13]) ? node12797 : node12788;
													assign node12788 = (inp[5]) ? 4'b0100 : node12789;
														assign node12789 = (inp[12]) ? node12791 : 4'b0100;
															assign node12791 = (inp[10]) ? 4'b0100 : node12792;
																assign node12792 = (inp[7]) ? 4'b1000 : 4'b1100;
													assign node12797 = (inp[10]) ? 4'b1100 : node12798;
														assign node12798 = (inp[12]) ? 4'b0100 : 4'b1100;
							assign node12802 = (inp[5]) ? node12804 : 4'b1110;
								assign node12804 = (inp[3]) ? node12944 : node12805;
									assign node12805 = (inp[4]) ? node12853 : node12806;
										assign node12806 = (inp[7]) ? 4'b1110 : node12807;
											assign node12807 = (inp[13]) ? node12825 : node12808;
												assign node12808 = (inp[12]) ? node12820 : node12809;
													assign node12809 = (inp[10]) ? node12817 : node12810;
														assign node12810 = (inp[1]) ? node12812 : 4'b1110;
															assign node12812 = (inp[11]) ? 4'b0000 : node12813;
																assign node12813 = (inp[14]) ? 4'b1110 : 4'b0000;
														assign node12817 = (inp[1]) ? 4'b0000 : 4'b0001;
													assign node12820 = (inp[10]) ? node12822 : 4'b1110;
														assign node12822 = (inp[1]) ? 4'b0000 : 4'b1110;
												assign node12825 = (inp[12]) ? node12841 : node12826;
													assign node12826 = (inp[1]) ? node12834 : node12827;
														assign node12827 = (inp[10]) ? 4'b1000 : node12828;
															assign node12828 = (inp[14]) ? node12830 : 4'b0001;
																assign node12830 = (inp[11]) ? 4'b0001 : 4'b0000;
														assign node12834 = (inp[11]) ? 4'b1000 : node12835;
															assign node12835 = (inp[14]) ? node12837 : 4'b1000;
																assign node12837 = (inp[10]) ? 4'b1001 : 4'b0001;
													assign node12841 = (inp[1]) ? node12845 : node12842;
														assign node12842 = (inp[11]) ? 4'b0001 : 4'b0000;
														assign node12845 = (inp[11]) ? node12849 : node12846;
															assign node12846 = (inp[14]) ? 4'b0001 : 4'b0000;
															assign node12849 = (inp[10]) ? 4'b1000 : 4'b0000;
										assign node12853 = (inp[13]) ? node12909 : node12854;
											assign node12854 = (inp[7]) ? node12884 : node12855;
												assign node12855 = (inp[1]) ? node12869 : node12856;
													assign node12856 = (inp[10]) ? node12862 : node12857;
														assign node12857 = (inp[11]) ? 4'b1001 : node12858;
															assign node12858 = (inp[14]) ? 4'b1000 : 4'b1001;
														assign node12862 = (inp[12]) ? 4'b1001 : node12863;
															assign node12863 = (inp[14]) ? node12865 : 4'b0001;
																assign node12865 = (inp[11]) ? 4'b0001 : 4'b0000;
													assign node12869 = (inp[11]) ? node12879 : node12870;
														assign node12870 = (inp[14]) ? node12874 : node12871;
															assign node12871 = (inp[12]) ? 4'b1000 : 4'b0000;
															assign node12874 = (inp[12]) ? 4'b1001 : node12875;
																assign node12875 = (inp[10]) ? 4'b0001 : 4'b1001;
														assign node12879 = (inp[12]) ? node12881 : 4'b0000;
															assign node12881 = (inp[10]) ? 4'b0000 : 4'b1000;
												assign node12884 = (inp[12]) ? node12900 : node12885;
													assign node12885 = (inp[10]) ? node12889 : node12886;
														assign node12886 = (inp[1]) ? 4'b0000 : 4'b1110;
														assign node12889 = (inp[1]) ? node12895 : node12890;
															assign node12890 = (inp[11]) ? 4'b0001 : node12891;
																assign node12891 = (inp[14]) ? 4'b0000 : 4'b0001;
															assign node12895 = (inp[11]) ? 4'b0000 : node12896;
																assign node12896 = (inp[14]) ? 4'b0001 : 4'b0000;
													assign node12900 = (inp[10]) ? node12902 : 4'b1110;
														assign node12902 = (inp[1]) ? node12904 : 4'b1110;
															assign node12904 = (inp[14]) ? node12906 : 4'b0000;
																assign node12906 = (inp[11]) ? 4'b0000 : 4'b1110;
											assign node12909 = (inp[1]) ? node12927 : node12910;
												assign node12910 = (inp[10]) ? node12916 : node12911;
													assign node12911 = (inp[14]) ? node12913 : 4'b0001;
														assign node12913 = (inp[11]) ? 4'b0001 : 4'b0000;
													assign node12916 = (inp[12]) ? node12922 : node12917;
														assign node12917 = (inp[14]) ? node12919 : 4'b1001;
															assign node12919 = (inp[7]) ? 4'b1000 : 4'b1001;
														assign node12922 = (inp[14]) ? node12924 : 4'b0001;
															assign node12924 = (inp[11]) ? 4'b0001 : 4'b0000;
												assign node12927 = (inp[11]) ? node12939 : node12928;
													assign node12928 = (inp[14]) ? node12934 : node12929;
														assign node12929 = (inp[12]) ? node12931 : 4'b1000;
															assign node12931 = (inp[10]) ? 4'b1000 : 4'b0000;
														assign node12934 = (inp[10]) ? node12936 : 4'b0001;
															assign node12936 = (inp[12]) ? 4'b0001 : 4'b1001;
													assign node12939 = (inp[12]) ? node12941 : 4'b1000;
														assign node12941 = (inp[10]) ? 4'b1000 : 4'b0000;
									assign node12944 = (inp[1]) ? node13026 : node12945;
										assign node12945 = (inp[13]) ? node12987 : node12946;
											assign node12946 = (inp[12]) ? node12974 : node12947;
												assign node12947 = (inp[10]) ? node12957 : node12948;
													assign node12948 = (inp[4]) ? node12954 : node12949;
														assign node12949 = (inp[11]) ? 4'b1001 : node12950;
															assign node12950 = (inp[14]) ? 4'b1000 : 4'b1001;
														assign node12954 = (inp[7]) ? 4'b1001 : 4'b1101;
													assign node12957 = (inp[7]) ? node12963 : node12958;
														assign node12958 = (inp[11]) ? 4'b0101 : node12959;
															assign node12959 = (inp[14]) ? 4'b0100 : 4'b0101;
														assign node12963 = (inp[4]) ? node12969 : node12964;
															assign node12964 = (inp[11]) ? 4'b0001 : node12965;
																assign node12965 = (inp[14]) ? 4'b0000 : 4'b0001;
															assign node12969 = (inp[14]) ? node12971 : 4'b0101;
																assign node12971 = (inp[11]) ? 4'b0101 : 4'b0100;
												assign node12974 = (inp[11]) ? node12982 : node12975;
													assign node12975 = (inp[14]) ? node12977 : 4'b1001;
														assign node12977 = (inp[4]) ? node12979 : 4'b1000;
															assign node12979 = (inp[7]) ? 4'b1000 : 4'b1100;
													assign node12982 = (inp[7]) ? 4'b1001 : node12983;
														assign node12983 = (inp[4]) ? 4'b1101 : 4'b1001;
											assign node12987 = (inp[14]) ? node13005 : node12988;
												assign node12988 = (inp[12]) ? node13000 : node12989;
													assign node12989 = (inp[10]) ? node12995 : node12990;
														assign node12990 = (inp[7]) ? node12992 : 4'b0101;
															assign node12992 = (inp[4]) ? 4'b0101 : 4'b0001;
														assign node12995 = (inp[7]) ? node12997 : 4'b1101;
															assign node12997 = (inp[4]) ? 4'b1101 : 4'b1001;
													assign node13000 = (inp[4]) ? 4'b0101 : node13001;
														assign node13001 = (inp[7]) ? 4'b0001 : 4'b0101;
												assign node13005 = (inp[11]) ? node13015 : node13006;
													assign node13006 = (inp[7]) ? node13012 : node13007;
														assign node13007 = (inp[10]) ? node13009 : 4'b0100;
															assign node13009 = (inp[12]) ? 4'b0100 : 4'b1100;
														assign node13012 = (inp[4]) ? 4'b0100 : 4'b0000;
													assign node13015 = (inp[12]) ? node13021 : node13016;
														assign node13016 = (inp[4]) ? 4'b1101 : node13017;
															assign node13017 = (inp[10]) ? 4'b1001 : 4'b0001;
														assign node13021 = (inp[7]) ? node13023 : 4'b0101;
															assign node13023 = (inp[4]) ? 4'b0101 : 4'b0001;
										assign node13026 = (inp[4]) ? node13066 : node13027;
											assign node13027 = (inp[7]) ? node13049 : node13028;
												assign node13028 = (inp[11]) ? node13038 : node13029;
													assign node13029 = (inp[14]) ? node13033 : node13030;
														assign node13030 = (inp[13]) ? 4'b1100 : 4'b0100;
														assign node13033 = (inp[13]) ? node13035 : 4'b1001;
															assign node13035 = (inp[10]) ? 4'b1101 : 4'b0101;
													assign node13038 = (inp[13]) ? node13044 : node13039;
														assign node13039 = (inp[10]) ? 4'b0100 : node13040;
															assign node13040 = (inp[12]) ? 4'b1000 : 4'b0100;
														assign node13044 = (inp[12]) ? node13046 : 4'b1100;
															assign node13046 = (inp[10]) ? 4'b1100 : 4'b0100;
												assign node13049 = (inp[14]) ? node13061 : node13050;
													assign node13050 = (inp[13]) ? node13056 : node13051;
														assign node13051 = (inp[10]) ? 4'b0000 : node13052;
															assign node13052 = (inp[12]) ? 4'b1000 : 4'b0000;
														assign node13056 = (inp[10]) ? 4'b1000 : node13057;
															assign node13057 = (inp[12]) ? 4'b0000 : 4'b1000;
													assign node13061 = (inp[11]) ? 4'b1000 : node13062;
														assign node13062 = (inp[13]) ? 4'b0001 : 4'b1001;
											assign node13066 = (inp[14]) ? node13080 : node13067;
												assign node13067 = (inp[13]) ? node13075 : node13068;
													assign node13068 = (inp[12]) ? node13070 : 4'b0100;
														assign node13070 = (inp[10]) ? 4'b0100 : node13071;
															assign node13071 = (inp[7]) ? 4'b1000 : 4'b1100;
													assign node13075 = (inp[10]) ? 4'b1100 : node13076;
														assign node13076 = (inp[12]) ? 4'b0100 : 4'b1100;
												assign node13080 = (inp[11]) ? node13090 : node13081;
													assign node13081 = (inp[13]) ? 4'b0101 : node13082;
														assign node13082 = (inp[12]) ? 4'b1001 : node13083;
															assign node13083 = (inp[10]) ? 4'b0101 : node13084;
																assign node13084 = (inp[7]) ? 4'b1001 : 4'b1101;
													assign node13090 = (inp[13]) ? node13098 : node13091;
														assign node13091 = (inp[12]) ? node13093 : 4'b0100;
															assign node13093 = (inp[10]) ? 4'b0100 : node13094;
																assign node13094 = (inp[7]) ? 4'b1000 : 4'b1100;
														assign node13098 = (inp[12]) ? node13100 : 4'b1100;
															assign node13100 = (inp[10]) ? 4'b1100 : 4'b0100;
					assign node13104 = (inp[5]) ? node14204 : node13105;
						assign node13105 = (inp[0]) ? node13853 : node13106;
							assign node13106 = (inp[11]) ? node13540 : node13107;
								assign node13107 = (inp[10]) ? node13319 : node13108;
									assign node13108 = (inp[13]) ? node13212 : node13109;
										assign node13109 = (inp[4]) ? node13165 : node13110;
											assign node13110 = (inp[3]) ? node13140 : node13111;
												assign node13111 = (inp[12]) ? node13127 : node13112;
													assign node13112 = (inp[1]) ? node13116 : node13113;
														assign node13113 = (inp[14]) ? 4'b1100 : 4'b1101;
														assign node13116 = (inp[14]) ? node13122 : node13117;
															assign node13117 = (inp[7]) ? 4'b0100 : node13118;
																assign node13118 = (inp[2]) ? 4'b0000 : 4'b0001;
															assign node13122 = (inp[2]) ? 4'b1101 : node13123;
																assign node13123 = (inp[7]) ? 4'b1101 : 4'b0001;
													assign node13127 = (inp[7]) ? node13133 : node13128;
														assign node13128 = (inp[1]) ? node13130 : 4'b1100;
															assign node13130 = (inp[14]) ? 4'b1101 : 4'b1100;
														assign node13133 = (inp[1]) ? node13137 : node13134;
															assign node13134 = (inp[14]) ? 4'b1100 : 4'b1101;
															assign node13137 = (inp[14]) ? 4'b1101 : 4'b1100;
												assign node13140 = (inp[2]) ? node13148 : node13141;
													assign node13141 = (inp[1]) ? node13143 : 4'b1101;
														assign node13143 = (inp[14]) ? node13145 : 4'b0001;
															assign node13145 = (inp[12]) ? 4'b1101 : 4'b0101;
													assign node13148 = (inp[12]) ? node13158 : node13149;
														assign node13149 = (inp[1]) ? node13153 : node13150;
															assign node13150 = (inp[7]) ? 4'b1001 : 4'b1000;
															assign node13153 = (inp[14]) ? 4'b1001 : node13154;
																assign node13154 = (inp[7]) ? 4'b0000 : 4'b0001;
														assign node13158 = (inp[14]) ? node13162 : node13159;
															assign node13159 = (inp[1]) ? 4'b1000 : 4'b1001;
															assign node13162 = (inp[1]) ? 4'b1001 : 4'b1000;
											assign node13165 = (inp[1]) ? node13185 : node13166;
												assign node13166 = (inp[7]) ? node13178 : node13167;
													assign node13167 = (inp[3]) ? node13173 : node13168;
														assign node13168 = (inp[14]) ? node13170 : 4'b1001;
															assign node13170 = (inp[2]) ? 4'b1000 : 4'b1001;
														assign node13173 = (inp[14]) ? 4'b1001 : node13174;
															assign node13174 = (inp[12]) ? 4'b1000 : 4'b0000;
													assign node13178 = (inp[3]) ? node13182 : node13179;
														assign node13179 = (inp[14]) ? 4'b1100 : 4'b1101;
														assign node13182 = (inp[2]) ? 4'b1001 : 4'b0000;
												assign node13185 = (inp[12]) ? node13199 : node13186;
													assign node13186 = (inp[7]) ? 4'b0001 : node13187;
														assign node13187 = (inp[3]) ? node13193 : node13188;
															assign node13188 = (inp[2]) ? node13190 : 4'b0101;
																assign node13190 = (inp[14]) ? 4'b1001 : 4'b0000;
															assign node13193 = (inp[2]) ? 4'b0101 : node13194;
																assign node13194 = (inp[14]) ? 4'b0000 : 4'b0001;
													assign node13199 = (inp[3]) ? node13207 : node13200;
														assign node13200 = (inp[2]) ? node13202 : 4'b1001;
															assign node13202 = (inp[14]) ? 4'b1101 : node13203;
																assign node13203 = (inp[7]) ? 4'b1100 : 4'b1000;
														assign node13207 = (inp[2]) ? 4'b1001 : node13208;
															assign node13208 = (inp[14]) ? 4'b0000 : 4'b0001;
										assign node13212 = (inp[3]) ? node13270 : node13213;
											assign node13213 = (inp[2]) ? node13243 : node13214;
												assign node13214 = (inp[4]) ? node13232 : node13215;
													assign node13215 = (inp[7]) ? node13221 : node13216;
														assign node13216 = (inp[14]) ? 4'b1001 : node13217;
															assign node13217 = (inp[1]) ? 4'b0001 : 4'b1001;
														assign node13221 = (inp[12]) ? node13225 : node13222;
															assign node13222 = (inp[1]) ? 4'b0001 : 4'b0101;
															assign node13225 = (inp[1]) ? node13229 : node13226;
																assign node13226 = (inp[14]) ? 4'b0100 : 4'b0101;
																assign node13229 = (inp[14]) ? 4'b0101 : 4'b0100;
													assign node13232 = (inp[7]) ? node13238 : node13233;
														assign node13233 = (inp[12]) ? 4'b1101 : node13234;
															assign node13234 = (inp[1]) ? 4'b0101 : 4'b1101;
														assign node13238 = (inp[12]) ? 4'b1001 : node13239;
															assign node13239 = (inp[1]) ? 4'b0101 : 4'b1001;
												assign node13243 = (inp[7]) ? node13253 : node13244;
													assign node13244 = (inp[1]) ? node13248 : node13245;
														assign node13245 = (inp[14]) ? 4'b0000 : 4'b0001;
														assign node13248 = (inp[14]) ? 4'b0001 : node13249;
															assign node13249 = (inp[12]) ? 4'b0000 : 4'b1000;
													assign node13253 = (inp[4]) ? node13261 : node13254;
														assign node13254 = (inp[1]) ? node13258 : node13255;
															assign node13255 = (inp[14]) ? 4'b0100 : 4'b0101;
															assign node13258 = (inp[12]) ? 4'b0100 : 4'b1100;
														assign node13261 = (inp[1]) ? node13265 : node13262;
															assign node13262 = (inp[14]) ? 4'b0000 : 4'b0001;
															assign node13265 = (inp[14]) ? 4'b0001 : node13266;
																assign node13266 = (inp[12]) ? 4'b0000 : 4'b1000;
											assign node13270 = (inp[4]) ? node13288 : node13271;
												assign node13271 = (inp[1]) ? node13279 : node13272;
													assign node13272 = (inp[2]) ? node13274 : 4'b1101;
														assign node13274 = (inp[7]) ? node13276 : 4'b1001;
															assign node13276 = (inp[14]) ? 4'b0000 : 4'b0001;
													assign node13279 = (inp[12]) ? node13281 : 4'b0001;
														assign node13281 = (inp[7]) ? node13283 : 4'b1001;
															assign node13283 = (inp[2]) ? node13285 : 4'b1101;
																assign node13285 = (inp[14]) ? 4'b0001 : 4'b0000;
												assign node13288 = (inp[7]) ? node13304 : node13289;
													assign node13289 = (inp[2]) ? node13299 : node13290;
														assign node13290 = (inp[1]) ? node13296 : node13291;
															assign node13291 = (inp[14]) ? 4'b0101 : node13292;
																assign node13292 = (inp[12]) ? 4'b0100 : 4'b1100;
															assign node13296 = (inp[14]) ? 4'b1100 : 4'b1101;
														assign node13299 = (inp[1]) ? node13301 : 4'b1101;
															assign node13301 = (inp[12]) ? 4'b1101 : 4'b0101;
													assign node13304 = (inp[2]) ? node13314 : node13305;
														assign node13305 = (inp[1]) ? node13311 : node13306;
															assign node13306 = (inp[14]) ? 4'b0001 : node13307;
																assign node13307 = (inp[12]) ? 4'b0000 : 4'b1000;
															assign node13311 = (inp[12]) ? 4'b1001 : 4'b1000;
														assign node13314 = (inp[12]) ? 4'b1001 : node13315;
															assign node13315 = (inp[1]) ? 4'b0101 : 4'b1001;
									assign node13319 = (inp[1]) ? node13413 : node13320;
										assign node13320 = (inp[4]) ? node13364 : node13321;
											assign node13321 = (inp[7]) ? node13333 : node13322;
												assign node13322 = (inp[2]) ? node13324 : 4'b0001;
													assign node13324 = (inp[3]) ? 4'b0001 : node13325;
														assign node13325 = (inp[14]) ? node13329 : node13326;
															assign node13326 = (inp[13]) ? 4'b1001 : 4'b0001;
															assign node13329 = (inp[13]) ? 4'b1000 : 4'b1100;
												assign node13333 = (inp[3]) ? node13351 : node13334;
													assign node13334 = (inp[14]) ? node13342 : node13335;
														assign node13335 = (inp[12]) ? node13339 : node13336;
															assign node13336 = (inp[13]) ? 4'b1101 : 4'b0101;
															assign node13339 = (inp[13]) ? 4'b0101 : 4'b1101;
														assign node13342 = (inp[12]) ? node13348 : node13343;
															assign node13343 = (inp[2]) ? 4'b1100 : node13344;
																assign node13344 = (inp[13]) ? 4'b0001 : 4'b0100;
															assign node13348 = (inp[13]) ? 4'b0100 : 4'b1100;
													assign node13351 = (inp[2]) ? node13355 : node13352;
														assign node13352 = (inp[13]) ? 4'b0001 : 4'b0101;
														assign node13355 = (inp[13]) ? 4'b0001 : node13356;
															assign node13356 = (inp[12]) ? node13360 : node13357;
																assign node13357 = (inp[14]) ? 4'b0000 : 4'b0001;
																assign node13360 = (inp[14]) ? 4'b1000 : 4'b1001;
											assign node13364 = (inp[13]) ? node13392 : node13365;
												assign node13365 = (inp[7]) ? node13377 : node13366;
													assign node13366 = (inp[3]) ? node13372 : node13367;
														assign node13367 = (inp[2]) ? node13369 : 4'b0101;
															assign node13369 = (inp[12]) ? 4'b1000 : 4'b0000;
														assign node13372 = (inp[2]) ? 4'b0101 : node13373;
															assign node13373 = (inp[12]) ? 4'b0001 : 4'b1000;
													assign node13377 = (inp[3]) ? node13385 : node13378;
														assign node13378 = (inp[2]) ? node13380 : 4'b0001;
															assign node13380 = (inp[12]) ? 4'b1100 : node13381;
																assign node13381 = (inp[14]) ? 4'b0000 : 4'b0001;
														assign node13385 = (inp[2]) ? 4'b0001 : node13386;
															assign node13386 = (inp[14]) ? node13388 : 4'b1000;
																assign node13388 = (inp[12]) ? 4'b0001 : 4'b1001;
												assign node13392 = (inp[3]) ? node13402 : node13393;
													assign node13393 = (inp[2]) ? node13395 : 4'b0101;
														assign node13395 = (inp[14]) ? node13399 : node13396;
															assign node13396 = (inp[12]) ? 4'b0001 : 4'b1001;
															assign node13399 = (inp[12]) ? 4'b0000 : 4'b1000;
													assign node13402 = (inp[14]) ? node13406 : node13403;
														assign node13403 = (inp[2]) ? 4'b0101 : 4'b0100;
														assign node13406 = (inp[2]) ? 4'b0101 : node13407;
															assign node13407 = (inp[12]) ? node13409 : 4'b0101;
																assign node13409 = (inp[7]) ? 4'b1001 : 4'b1101;
										assign node13413 = (inp[12]) ? node13479 : node13414;
											assign node13414 = (inp[13]) ? node13452 : node13415;
												assign node13415 = (inp[2]) ? node13433 : node13416;
													assign node13416 = (inp[4]) ? node13424 : node13417;
														assign node13417 = (inp[7]) ? node13419 : 4'b1001;
															assign node13419 = (inp[3]) ? 4'b1101 : node13420;
																assign node13420 = (inp[14]) ? 4'b0101 : 4'b0100;
														assign node13424 = (inp[3]) ? node13428 : node13425;
															assign node13425 = (inp[7]) ? 4'b1001 : 4'b1101;
															assign node13428 = (inp[7]) ? 4'b0001 : node13429;
																assign node13429 = (inp[14]) ? 4'b0100 : 4'b0101;
													assign node13433 = (inp[3]) ? node13443 : node13434;
														assign node13434 = (inp[14]) ? node13438 : node13435;
															assign node13435 = (inp[4]) ? 4'b0000 : 4'b0100;
															assign node13438 = (inp[7]) ? node13440 : 4'b0001;
																assign node13440 = (inp[4]) ? 4'b0001 : 4'b0101;
														assign node13443 = (inp[7]) ? node13447 : node13444;
															assign node13444 = (inp[4]) ? 4'b1101 : 4'b1001;
															assign node13447 = (inp[4]) ? 4'b1001 : node13448;
																assign node13448 = (inp[14]) ? 4'b0001 : 4'b0000;
												assign node13452 = (inp[4]) ? node13468 : node13453;
													assign node13453 = (inp[2]) ? node13461 : node13454;
														assign node13454 = (inp[14]) ? node13456 : 4'b1001;
															assign node13456 = (inp[7]) ? 4'b1001 : node13457;
																assign node13457 = (inp[3]) ? 4'b1000 : 4'b1001;
														assign node13461 = (inp[3]) ? 4'b1001 : node13462;
															assign node13462 = (inp[7]) ? 4'b1100 : node13463;
																assign node13463 = (inp[14]) ? 4'b1001 : 4'b1000;
													assign node13468 = (inp[3]) ? node13474 : node13469;
														assign node13469 = (inp[2]) ? node13471 : 4'b1101;
															assign node13471 = (inp[14]) ? 4'b1001 : 4'b1000;
														assign node13474 = (inp[2]) ? 4'b1101 : node13475;
															assign node13475 = (inp[14]) ? 4'b1100 : 4'b1101;
											assign node13479 = (inp[3]) ? node13511 : node13480;
												assign node13480 = (inp[2]) ? node13492 : node13481;
													assign node13481 = (inp[4]) ? node13487 : node13482;
														assign node13482 = (inp[13]) ? 4'b0001 : node13483;
															assign node13483 = (inp[14]) ? 4'b1101 : 4'b0100;
														assign node13487 = (inp[13]) ? 4'b0101 : node13488;
															assign node13488 = (inp[7]) ? 4'b0001 : 4'b0101;
													assign node13492 = (inp[14]) ? node13502 : node13493;
														assign node13493 = (inp[13]) ? node13497 : node13494;
															assign node13494 = (inp[4]) ? 4'b0000 : 4'b0100;
															assign node13497 = (inp[4]) ? 4'b1000 : node13498;
																assign node13498 = (inp[7]) ? 4'b1100 : 4'b1000;
														assign node13502 = (inp[13]) ? node13508 : node13503;
															assign node13503 = (inp[4]) ? node13505 : 4'b1101;
																assign node13505 = (inp[7]) ? 4'b1101 : 4'b1001;
															assign node13508 = (inp[4]) ? 4'b0001 : 4'b0101;
												assign node13511 = (inp[4]) ? node13527 : node13512;
													assign node13512 = (inp[13]) ? node13520 : node13513;
														assign node13513 = (inp[2]) ? node13517 : node13514;
															assign node13514 = (inp[7]) ? 4'b0101 : 4'b0001;
															assign node13517 = (inp[14]) ? 4'b1001 : 4'b0001;
														assign node13520 = (inp[14]) ? node13522 : 4'b0001;
															assign node13522 = (inp[2]) ? 4'b0001 : node13523;
																assign node13523 = (inp[7]) ? 4'b0001 : 4'b0000;
													assign node13527 = (inp[13]) ? node13535 : node13528;
														assign node13528 = (inp[2]) ? node13532 : node13529;
															assign node13529 = (inp[14]) ? 4'b1000 : 4'b1001;
															assign node13532 = (inp[7]) ? 4'b0001 : 4'b0101;
														assign node13535 = (inp[14]) ? node13537 : 4'b0101;
															assign node13537 = (inp[2]) ? 4'b0101 : 4'b0100;
								assign node13540 = (inp[1]) ? node13744 : node13541;
									assign node13541 = (inp[3]) ? node13631 : node13542;
										assign node13542 = (inp[2]) ? node13596 : node13543;
											assign node13543 = (inp[4]) ? node13565 : node13544;
												assign node13544 = (inp[13]) ? node13556 : node13545;
													assign node13545 = (inp[7]) ? node13551 : node13546;
														assign node13546 = (inp[12]) ? node13548 : 4'b0000;
															assign node13548 = (inp[10]) ? 4'b0000 : 4'b1101;
														assign node13551 = (inp[10]) ? node13553 : 4'b1101;
															assign node13553 = (inp[12]) ? 4'b1101 : 4'b0101;
													assign node13556 = (inp[12]) ? node13560 : node13557;
														assign node13557 = (inp[10]) ? 4'b1000 : 4'b0000;
														assign node13560 = (inp[10]) ? 4'b0000 : node13561;
															assign node13561 = (inp[7]) ? 4'b0101 : 4'b1000;
												assign node13565 = (inp[7]) ? node13585 : node13566;
													assign node13566 = (inp[14]) ? node13576 : node13567;
														assign node13567 = (inp[12]) ? node13571 : node13568;
															assign node13568 = (inp[10]) ? 4'b1100 : 4'b0100;
															assign node13571 = (inp[10]) ? 4'b0100 : node13572;
																assign node13572 = (inp[13]) ? 4'b1100 : 4'b1000;
														assign node13576 = (inp[13]) ? node13580 : node13577;
															assign node13577 = (inp[12]) ? 4'b0100 : 4'b1100;
															assign node13580 = (inp[10]) ? 4'b0100 : node13581;
																assign node13581 = (inp[12]) ? 4'b1100 : 4'b0100;
													assign node13585 = (inp[10]) ? node13591 : node13586;
														assign node13586 = (inp[12]) ? 4'b1000 : node13587;
															assign node13587 = (inp[13]) ? 4'b0100 : 4'b0000;
														assign node13591 = (inp[12]) ? node13593 : 4'b1100;
															assign node13593 = (inp[13]) ? 4'b0100 : 4'b0000;
											assign node13596 = (inp[13]) ? node13614 : node13597;
												assign node13597 = (inp[7]) ? node13607 : node13598;
													assign node13598 = (inp[4]) ? node13602 : node13599;
														assign node13599 = (inp[10]) ? 4'b0001 : 4'b1101;
														assign node13602 = (inp[12]) ? 4'b1001 : node13603;
															assign node13603 = (inp[10]) ? 4'b0001 : 4'b1001;
													assign node13607 = (inp[12]) ? 4'b1101 : node13608;
														assign node13608 = (inp[10]) ? node13610 : 4'b1101;
															assign node13610 = (inp[4]) ? 4'b0001 : 4'b0101;
												assign node13614 = (inp[10]) ? node13620 : node13615;
													assign node13615 = (inp[7]) ? node13617 : 4'b0001;
														assign node13617 = (inp[4]) ? 4'b0001 : 4'b0101;
													assign node13620 = (inp[12]) ? node13626 : node13621;
														assign node13621 = (inp[14]) ? node13623 : 4'b1001;
															assign node13623 = (inp[4]) ? 4'b1001 : 4'b1101;
														assign node13626 = (inp[4]) ? 4'b0001 : node13627;
															assign node13627 = (inp[7]) ? 4'b0101 : 4'b0001;
										assign node13631 = (inp[2]) ? node13685 : node13632;
											assign node13632 = (inp[4]) ? node13666 : node13633;
												assign node13633 = (inp[7]) ? node13645 : node13634;
													assign node13634 = (inp[10]) ? node13640 : node13635;
														assign node13635 = (inp[12]) ? node13637 : 4'b0000;
															assign node13637 = (inp[13]) ? 4'b1000 : 4'b1100;
														assign node13640 = (inp[13]) ? 4'b0001 : node13641;
															assign node13641 = (inp[14]) ? 4'b0000 : 4'b1000;
													assign node13645 = (inp[13]) ? node13659 : node13646;
														assign node13646 = (inp[14]) ? node13652 : node13647;
															assign node13647 = (inp[10]) ? 4'b0100 : node13648;
																assign node13648 = (inp[12]) ? 4'b1100 : 4'b0100;
															assign node13652 = (inp[12]) ? node13656 : node13653;
																assign node13653 = (inp[10]) ? 4'b1100 : 4'b0100;
																assign node13656 = (inp[10]) ? 4'b0100 : 4'b1100;
														assign node13659 = (inp[10]) ? node13663 : node13660;
															assign node13660 = (inp[12]) ? 4'b1100 : 4'b0000;
															assign node13663 = (inp[12]) ? 4'b0000 : 4'b1000;
												assign node13666 = (inp[13]) ? node13676 : node13667;
													assign node13667 = (inp[12]) ? node13671 : node13668;
														assign node13668 = (inp[10]) ? 4'b1001 : 4'b0001;
														assign node13671 = (inp[7]) ? node13673 : 4'b1001;
															assign node13673 = (inp[10]) ? 4'b1001 : 4'b1000;
													assign node13676 = (inp[10]) ? 4'b0101 : node13677;
														assign node13677 = (inp[12]) ? node13681 : node13678;
															assign node13678 = (inp[7]) ? 4'b1001 : 4'b1101;
															assign node13681 = (inp[7]) ? 4'b0001 : 4'b0101;
											assign node13685 = (inp[4]) ? node13715 : node13686;
												assign node13686 = (inp[7]) ? node13704 : node13687;
													assign node13687 = (inp[13]) ? node13693 : node13688;
														assign node13688 = (inp[10]) ? node13690 : 4'b0000;
															assign node13690 = (inp[12]) ? 4'b0000 : 4'b1000;
														assign node13693 = (inp[14]) ? node13699 : node13694;
															assign node13694 = (inp[12]) ? node13696 : 4'b1000;
																assign node13696 = (inp[10]) ? 4'b0000 : 4'b1000;
															assign node13699 = (inp[12]) ? 4'b1000 : node13700;
																assign node13700 = (inp[10]) ? 4'b1000 : 4'b0000;
													assign node13704 = (inp[13]) ? node13710 : node13705;
														assign node13705 = (inp[14]) ? 4'b1001 : node13706;
															assign node13706 = (inp[10]) ? 4'b0001 : 4'b1001;
														assign node13710 = (inp[12]) ? 4'b0001 : node13711;
															assign node13711 = (inp[10]) ? 4'b1000 : 4'b0000;
												assign node13715 = (inp[13]) ? node13735 : node13716;
													assign node13716 = (inp[7]) ? node13724 : node13717;
														assign node13717 = (inp[10]) ? node13721 : node13718;
															assign node13718 = (inp[12]) ? 4'b1000 : 4'b0100;
															assign node13721 = (inp[12]) ? 4'b0100 : 4'b1100;
														assign node13724 = (inp[14]) ? node13730 : node13725;
															assign node13725 = (inp[12]) ? node13727 : 4'b1000;
																assign node13727 = (inp[10]) ? 4'b0000 : 4'b1000;
															assign node13730 = (inp[12]) ? 4'b0000 : node13731;
																assign node13731 = (inp[10]) ? 4'b1000 : 4'b0000;
													assign node13735 = (inp[10]) ? node13741 : node13736;
														assign node13736 = (inp[12]) ? node13738 : 4'b0100;
															assign node13738 = (inp[7]) ? 4'b1000 : 4'b1100;
														assign node13741 = (inp[12]) ? 4'b0100 : 4'b1100;
									assign node13744 = (inp[10]) ? node13812 : node13745;
										assign node13745 = (inp[4]) ? node13777 : node13746;
											assign node13746 = (inp[7]) ? node13756 : node13747;
												assign node13747 = (inp[2]) ? node13749 : 4'b0000;
													assign node13749 = (inp[3]) ? 4'b0000 : node13750;
														assign node13750 = (inp[13]) ? 4'b0000 : node13751;
															assign node13751 = (inp[12]) ? 4'b1100 : 4'b0000;
												assign node13756 = (inp[3]) ? node13770 : node13757;
													assign node13757 = (inp[2]) ? node13763 : node13758;
														assign node13758 = (inp[13]) ? 4'b0000 : node13759;
															assign node13759 = (inp[12]) ? 4'b1100 : 4'b0100;
														assign node13763 = (inp[13]) ? node13767 : node13764;
															assign node13764 = (inp[12]) ? 4'b1100 : 4'b0100;
															assign node13767 = (inp[12]) ? 4'b0100 : 4'b1100;
													assign node13770 = (inp[2]) ? node13774 : node13771;
														assign node13771 = (inp[13]) ? 4'b0000 : 4'b0100;
														assign node13774 = (inp[12]) ? 4'b1000 : 4'b0000;
											assign node13777 = (inp[13]) ? node13801 : node13778;
												assign node13778 = (inp[7]) ? node13790 : node13779;
													assign node13779 = (inp[2]) ? node13785 : node13780;
														assign node13780 = (inp[3]) ? node13782 : 4'b0100;
															assign node13782 = (inp[12]) ? 4'b0000 : 4'b1000;
														assign node13785 = (inp[3]) ? 4'b0100 : node13786;
															assign node13786 = (inp[12]) ? 4'b1000 : 4'b0000;
													assign node13790 = (inp[2]) ? node13796 : node13791;
														assign node13791 = (inp[3]) ? node13793 : 4'b0000;
															assign node13793 = (inp[12]) ? 4'b0000 : 4'b1000;
														assign node13796 = (inp[3]) ? 4'b0000 : node13797;
															assign node13797 = (inp[12]) ? 4'b1100 : 4'b0000;
												assign node13801 = (inp[2]) ? node13807 : node13802;
													assign node13802 = (inp[3]) ? node13804 : 4'b0100;
														assign node13804 = (inp[12]) ? 4'b1100 : 4'b0100;
													assign node13807 = (inp[3]) ? 4'b0100 : node13808;
														assign node13808 = (inp[12]) ? 4'b0000 : 4'b1000;
										assign node13812 = (inp[13]) ? node13840 : node13813;
											assign node13813 = (inp[2]) ? node13827 : node13814;
												assign node13814 = (inp[4]) ? node13820 : node13815;
													assign node13815 = (inp[7]) ? node13817 : 4'b1000;
														assign node13817 = (inp[3]) ? 4'b1100 : 4'b0100;
													assign node13820 = (inp[3]) ? node13824 : node13821;
														assign node13821 = (inp[7]) ? 4'b1000 : 4'b1100;
														assign node13824 = (inp[7]) ? 4'b0000 : 4'b0100;
												assign node13827 = (inp[3]) ? node13833 : node13828;
													assign node13828 = (inp[4]) ? 4'b0000 : node13829;
														assign node13829 = (inp[7]) ? 4'b0100 : 4'b0000;
													assign node13833 = (inp[4]) ? node13837 : node13834;
														assign node13834 = (inp[7]) ? 4'b0000 : 4'b1000;
														assign node13837 = (inp[7]) ? 4'b1000 : 4'b1100;
											assign node13840 = (inp[4]) ? node13848 : node13841;
												assign node13841 = (inp[3]) ? 4'b1000 : node13842;
													assign node13842 = (inp[2]) ? node13844 : 4'b1000;
														assign node13844 = (inp[7]) ? 4'b1100 : 4'b1000;
												assign node13848 = (inp[3]) ? 4'b1100 : node13849;
													assign node13849 = (inp[2]) ? 4'b1000 : 4'b1100;
							assign node13853 = (inp[2]) ? 4'b1100 : node13854;
								assign node13854 = (inp[1]) ? node14026 : node13855;
									assign node13855 = (inp[11]) ? node13959 : node13856;
										assign node13856 = (inp[14]) ? node13906 : node13857;
											assign node13857 = (inp[3]) ? node13875 : node13858;
												assign node13858 = (inp[7]) ? 4'b1100 : node13859;
													assign node13859 = (inp[13]) ? node13869 : node13860;
														assign node13860 = (inp[4]) ? node13866 : node13861;
															assign node13861 = (inp[10]) ? node13863 : 4'b1100;
																assign node13863 = (inp[12]) ? 4'b1100 : 4'b0001;
															assign node13866 = (inp[12]) ? 4'b1001 : 4'b0001;
														assign node13869 = (inp[12]) ? 4'b0001 : node13870;
															assign node13870 = (inp[10]) ? 4'b1001 : 4'b0001;
												assign node13875 = (inp[4]) ? node13895 : node13876;
													assign node13876 = (inp[7]) ? node13886 : node13877;
														assign node13877 = (inp[10]) ? node13879 : 4'b1001;
															assign node13879 = (inp[12]) ? node13883 : node13880;
																assign node13880 = (inp[13]) ? 4'b1101 : 4'b0101;
																assign node13883 = (inp[13]) ? 4'b0101 : 4'b1001;
														assign node13886 = (inp[13]) ? node13890 : node13887;
															assign node13887 = (inp[12]) ? 4'b1001 : 4'b0001;
															assign node13890 = (inp[12]) ? 4'b0001 : node13891;
																assign node13891 = (inp[10]) ? 4'b1001 : 4'b0001;
													assign node13895 = (inp[13]) ? node13901 : node13896;
														assign node13896 = (inp[10]) ? node13898 : 4'b1001;
															assign node13898 = (inp[12]) ? 4'b1101 : 4'b0101;
														assign node13901 = (inp[12]) ? 4'b0101 : node13902;
															assign node13902 = (inp[10]) ? 4'b1101 : 4'b0101;
											assign node13906 = (inp[13]) ? node13934 : node13907;
												assign node13907 = (inp[10]) ? node13919 : node13908;
													assign node13908 = (inp[3]) ? node13914 : node13909;
														assign node13909 = (inp[4]) ? node13911 : 4'b1100;
															assign node13911 = (inp[7]) ? 4'b1100 : 4'b1000;
														assign node13914 = (inp[4]) ? node13916 : 4'b1000;
															assign node13916 = (inp[7]) ? 4'b1000 : 4'b1100;
													assign node13919 = (inp[12]) ? node13931 : node13920;
														assign node13920 = (inp[3]) ? node13926 : node13921;
															assign node13921 = (inp[4]) ? 4'b0000 : node13922;
																assign node13922 = (inp[7]) ? 4'b1100 : 4'b0000;
															assign node13926 = (inp[7]) ? node13928 : 4'b0100;
																assign node13928 = (inp[4]) ? 4'b0100 : 4'b0000;
														assign node13931 = (inp[4]) ? 4'b1000 : 4'b1100;
												assign node13934 = (inp[10]) ? node13946 : node13935;
													assign node13935 = (inp[3]) ? node13941 : node13936;
														assign node13936 = (inp[7]) ? node13938 : 4'b0000;
															assign node13938 = (inp[4]) ? 4'b0000 : 4'b1100;
														assign node13941 = (inp[4]) ? 4'b0100 : node13942;
															assign node13942 = (inp[7]) ? 4'b0000 : 4'b0100;
													assign node13946 = (inp[12]) ? node13956 : node13947;
														assign node13947 = (inp[3]) ? node13953 : node13948;
															assign node13948 = (inp[7]) ? node13950 : 4'b1000;
																assign node13950 = (inp[4]) ? 4'b1000 : 4'b1100;
															assign node13953 = (inp[7]) ? 4'b1000 : 4'b1100;
														assign node13956 = (inp[3]) ? 4'b0100 : 4'b1100;
										assign node13959 = (inp[3]) ? node13991 : node13960;
											assign node13960 = (inp[4]) ? node13974 : node13961;
												assign node13961 = (inp[7]) ? 4'b1100 : node13962;
													assign node13962 = (inp[13]) ? node13968 : node13963;
														assign node13963 = (inp[12]) ? 4'b1100 : node13964;
															assign node13964 = (inp[10]) ? 4'b0001 : 4'b1100;
														assign node13968 = (inp[12]) ? 4'b0001 : node13969;
															assign node13969 = (inp[14]) ? 4'b0001 : 4'b1001;
												assign node13974 = (inp[13]) ? node13986 : node13975;
													assign node13975 = (inp[7]) ? node13981 : node13976;
														assign node13976 = (inp[10]) ? node13978 : 4'b1001;
															assign node13978 = (inp[12]) ? 4'b1001 : 4'b0001;
														assign node13981 = (inp[10]) ? node13983 : 4'b1100;
															assign node13983 = (inp[12]) ? 4'b1100 : 4'b0001;
													assign node13986 = (inp[12]) ? 4'b0001 : node13987;
														assign node13987 = (inp[10]) ? 4'b1001 : 4'b0001;
											assign node13991 = (inp[13]) ? node14009 : node13992;
												assign node13992 = (inp[12]) ? node14004 : node13993;
													assign node13993 = (inp[10]) ? node13999 : node13994;
														assign node13994 = (inp[4]) ? node13996 : 4'b1001;
															assign node13996 = (inp[7]) ? 4'b1001 : 4'b1101;
														assign node13999 = (inp[7]) ? node14001 : 4'b0101;
															assign node14001 = (inp[4]) ? 4'b0101 : 4'b0001;
													assign node14004 = (inp[7]) ? 4'b1001 : node14005;
														assign node14005 = (inp[4]) ? 4'b1101 : 4'b1001;
												assign node14009 = (inp[4]) ? node14021 : node14010;
													assign node14010 = (inp[7]) ? node14016 : node14011;
														assign node14011 = (inp[10]) ? node14013 : 4'b0101;
															assign node14013 = (inp[12]) ? 4'b0101 : 4'b1101;
														assign node14016 = (inp[12]) ? 4'b0001 : node14017;
															assign node14017 = (inp[10]) ? 4'b1001 : 4'b0001;
													assign node14021 = (inp[12]) ? 4'b0101 : node14022;
														assign node14022 = (inp[10]) ? 4'b1101 : 4'b0101;
									assign node14026 = (inp[14]) ? node14092 : node14027;
										assign node14027 = (inp[3]) ? node14055 : node14028;
											assign node14028 = (inp[4]) ? node14042 : node14029;
												assign node14029 = (inp[7]) ? 4'b1100 : node14030;
													assign node14030 = (inp[13]) ? node14036 : node14031;
														assign node14031 = (inp[10]) ? 4'b0000 : node14032;
															assign node14032 = (inp[12]) ? 4'b1100 : 4'b0000;
														assign node14036 = (inp[12]) ? node14038 : 4'b1000;
															assign node14038 = (inp[10]) ? 4'b1000 : 4'b0000;
												assign node14042 = (inp[13]) ? node14050 : node14043;
													assign node14043 = (inp[12]) ? node14045 : 4'b0000;
														assign node14045 = (inp[10]) ? 4'b0000 : node14046;
															assign node14046 = (inp[7]) ? 4'b1100 : 4'b1000;
													assign node14050 = (inp[12]) ? node14052 : 4'b1000;
														assign node14052 = (inp[10]) ? 4'b1000 : 4'b0000;
											assign node14055 = (inp[4]) ? node14079 : node14056;
												assign node14056 = (inp[7]) ? node14068 : node14057;
													assign node14057 = (inp[13]) ? node14063 : node14058;
														assign node14058 = (inp[10]) ? 4'b0100 : node14059;
															assign node14059 = (inp[12]) ? 4'b1000 : 4'b0100;
														assign node14063 = (inp[10]) ? 4'b1100 : node14064;
															assign node14064 = (inp[12]) ? 4'b0100 : 4'b1100;
													assign node14068 = (inp[13]) ? node14074 : node14069;
														assign node14069 = (inp[10]) ? 4'b0000 : node14070;
															assign node14070 = (inp[12]) ? 4'b1000 : 4'b0000;
														assign node14074 = (inp[12]) ? node14076 : 4'b1000;
															assign node14076 = (inp[10]) ? 4'b1000 : 4'b0000;
												assign node14079 = (inp[13]) ? node14087 : node14080;
													assign node14080 = (inp[12]) ? node14082 : 4'b0100;
														assign node14082 = (inp[10]) ? 4'b0100 : node14083;
															assign node14083 = (inp[11]) ? 4'b1000 : 4'b1100;
													assign node14087 = (inp[12]) ? node14089 : 4'b1100;
														assign node14089 = (inp[10]) ? 4'b1100 : 4'b0100;
										assign node14092 = (inp[11]) ? node14146 : node14093;
											assign node14093 = (inp[13]) ? node14119 : node14094;
												assign node14094 = (inp[3]) ? node14108 : node14095;
													assign node14095 = (inp[7]) ? node14103 : node14096;
														assign node14096 = (inp[4]) ? 4'b1001 : node14097;
															assign node14097 = (inp[10]) ? node14099 : 4'b1100;
																assign node14099 = (inp[12]) ? 4'b1100 : 4'b0001;
														assign node14103 = (inp[10]) ? node14105 : 4'b1100;
															assign node14105 = (inp[12]) ? 4'b1100 : 4'b0001;
													assign node14108 = (inp[7]) ? node14116 : node14109;
														assign node14109 = (inp[4]) ? node14111 : 4'b1001;
															assign node14111 = (inp[12]) ? 4'b1101 : node14112;
																assign node14112 = (inp[10]) ? 4'b0101 : 4'b1101;
														assign node14116 = (inp[12]) ? 4'b1001 : 4'b0001;
												assign node14119 = (inp[3]) ? node14129 : node14120;
													assign node14120 = (inp[7]) ? node14126 : node14121;
														assign node14121 = (inp[10]) ? node14123 : 4'b0001;
															assign node14123 = (inp[12]) ? 4'b0001 : 4'b1001;
														assign node14126 = (inp[4]) ? 4'b0001 : 4'b1100;
													assign node14129 = (inp[12]) ? node14141 : node14130;
														assign node14130 = (inp[10]) ? node14136 : node14131;
															assign node14131 = (inp[7]) ? node14133 : 4'b0101;
																assign node14133 = (inp[4]) ? 4'b0101 : 4'b0001;
															assign node14136 = (inp[4]) ? 4'b1101 : node14137;
																assign node14137 = (inp[7]) ? 4'b1001 : 4'b1101;
														assign node14141 = (inp[4]) ? 4'b0101 : node14142;
															assign node14142 = (inp[7]) ? 4'b0001 : 4'b0101;
											assign node14146 = (inp[13]) ? node14176 : node14147;
												assign node14147 = (inp[12]) ? node14155 : node14148;
													assign node14148 = (inp[10]) ? 4'b1100 : node14149;
														assign node14149 = (inp[4]) ? node14151 : 4'b0000;
															assign node14151 = (inp[3]) ? 4'b0100 : 4'b0000;
													assign node14155 = (inp[10]) ? node14167 : node14156;
														assign node14156 = (inp[3]) ? node14162 : node14157;
															assign node14157 = (inp[7]) ? 4'b1100 : node14158;
																assign node14158 = (inp[4]) ? 4'b1000 : 4'b1100;
															assign node14162 = (inp[4]) ? node14164 : 4'b1000;
																assign node14164 = (inp[7]) ? 4'b1000 : 4'b1100;
														assign node14167 = (inp[7]) ? node14169 : 4'b0000;
															assign node14169 = (inp[3]) ? node14173 : node14170;
																assign node14170 = (inp[4]) ? 4'b0000 : 4'b1100;
																assign node14173 = (inp[4]) ? 4'b0100 : 4'b0000;
												assign node14176 = (inp[3]) ? node14186 : node14177;
													assign node14177 = (inp[4]) ? node14181 : node14178;
														assign node14178 = (inp[7]) ? 4'b1100 : 4'b1000;
														assign node14181 = (inp[12]) ? node14183 : 4'b1000;
															assign node14183 = (inp[10]) ? 4'b1000 : 4'b0000;
													assign node14186 = (inp[7]) ? node14192 : node14187;
														assign node14187 = (inp[12]) ? node14189 : 4'b1100;
															assign node14189 = (inp[10]) ? 4'b1100 : 4'b0100;
														assign node14192 = (inp[4]) ? node14198 : node14193;
															assign node14193 = (inp[10]) ? 4'b1000 : node14194;
																assign node14194 = (inp[12]) ? 4'b0000 : 4'b1000;
															assign node14198 = (inp[12]) ? node14200 : 4'b1100;
																assign node14200 = (inp[10]) ? 4'b1100 : 4'b0100;
						assign node14204 = (inp[3]) ? node14974 : node14205;
							assign node14205 = (inp[4]) ? node14577 : node14206;
								assign node14206 = (inp[7]) ? node14402 : node14207;
									assign node14207 = (inp[1]) ? node14307 : node14208;
										assign node14208 = (inp[2]) ? node14246 : node14209;
											assign node14209 = (inp[0]) ? node14229 : node14210;
												assign node14210 = (inp[13]) ? node14218 : node14211;
													assign node14211 = (inp[11]) ? 4'b0000 : node14212;
														assign node14212 = (inp[12]) ? node14214 : 4'b0000;
															assign node14214 = (inp[10]) ? 4'b1000 : 4'b1101;
													assign node14218 = (inp[12]) ? node14224 : node14219;
														assign node14219 = (inp[10]) ? node14221 : 4'b0100;
															assign node14221 = (inp[11]) ? 4'b0001 : 4'b0100;
														assign node14224 = (inp[11]) ? 4'b0100 : node14225;
															assign node14225 = (inp[10]) ? 4'b1100 : 4'b1000;
												assign node14229 = (inp[11]) ? node14237 : node14230;
													assign node14230 = (inp[10]) ? 4'b0001 : node14231;
														assign node14231 = (inp[13]) ? 4'b1001 : node14232;
															assign node14232 = (inp[14]) ? 4'b1100 : 4'b1101;
													assign node14237 = (inp[10]) ? node14243 : node14238;
														assign node14238 = (inp[12]) ? node14240 : 4'b0000;
															assign node14240 = (inp[13]) ? 4'b1000 : 4'b1101;
														assign node14243 = (inp[12]) ? 4'b0000 : 4'b1000;
											assign node14246 = (inp[13]) ? node14272 : node14247;
												assign node14247 = (inp[0]) ? node14265 : node14248;
													assign node14248 = (inp[10]) ? node14258 : node14249;
														assign node14249 = (inp[12]) ? node14255 : node14250;
															assign node14250 = (inp[11]) ? 4'b0001 : node14251;
																assign node14251 = (inp[14]) ? 4'b1101 : 4'b0000;
															assign node14255 = (inp[11]) ? 4'b1100 : 4'b1101;
														assign node14258 = (inp[11]) ? 4'b1001 : node14259;
															assign node14259 = (inp[12]) ? 4'b0001 : node14260;
																assign node14260 = (inp[14]) ? 4'b1001 : 4'b1000;
													assign node14265 = (inp[10]) ? node14267 : 4'b1100;
														assign node14267 = (inp[12]) ? 4'b1100 : node14268;
															assign node14268 = (inp[11]) ? 4'b0001 : 4'b0000;
												assign node14272 = (inp[11]) ? node14294 : node14273;
													assign node14273 = (inp[10]) ? node14285 : node14274;
														assign node14274 = (inp[12]) ? node14280 : node14275;
															assign node14275 = (inp[14]) ? node14277 : 4'b1000;
																assign node14277 = (inp[0]) ? 4'b0000 : 4'b0001;
															assign node14280 = (inp[14]) ? 4'b0001 : node14281;
																assign node14281 = (inp[0]) ? 4'b0001 : 4'b0000;
														assign node14285 = (inp[0]) ? node14289 : node14286;
															assign node14286 = (inp[14]) ? 4'b1001 : 4'b0100;
															assign node14289 = (inp[12]) ? 4'b0000 : node14290;
																assign node14290 = (inp[14]) ? 4'b1000 : 4'b1001;
													assign node14294 = (inp[12]) ? node14302 : node14295;
														assign node14295 = (inp[10]) ? node14299 : node14296;
															assign node14296 = (inp[0]) ? 4'b0001 : 4'b1001;
															assign node14299 = (inp[0]) ? 4'b1001 : 4'b0101;
														assign node14302 = (inp[0]) ? 4'b0001 : node14303;
															assign node14303 = (inp[10]) ? 4'b0101 : 4'b0001;
										assign node14307 = (inp[11]) ? node14369 : node14308;
											assign node14308 = (inp[0]) ? node14342 : node14309;
												assign node14309 = (inp[13]) ? node14325 : node14310;
													assign node14310 = (inp[14]) ? node14316 : node14311;
														assign node14311 = (inp[2]) ? 4'b0001 : node14312;
															assign node14312 = (inp[12]) ? 4'b0000 : 4'b1000;
														assign node14316 = (inp[12]) ? node14320 : node14317;
															assign node14317 = (inp[2]) ? 4'b0000 : 4'b1000;
															assign node14320 = (inp[2]) ? node14322 : 4'b0000;
																assign node14322 = (inp[10]) ? 4'b1000 : 4'b0000;
													assign node14325 = (inp[2]) ? node14333 : node14326;
														assign node14326 = (inp[10]) ? node14330 : node14327;
															assign node14327 = (inp[12]) ? 4'b0100 : 4'b1100;
															assign node14330 = (inp[14]) ? 4'b0001 : 4'b0000;
														assign node14333 = (inp[10]) ? node14337 : node14334;
															assign node14334 = (inp[14]) ? 4'b1000 : 4'b1001;
															assign node14337 = (inp[14]) ? node14339 : 4'b1101;
																assign node14339 = (inp[12]) ? 4'b0100 : 4'b1100;
												assign node14342 = (inp[2]) ? node14354 : node14343;
													assign node14343 = (inp[10]) ? node14351 : node14344;
														assign node14344 = (inp[12]) ? node14346 : 4'b0001;
															assign node14346 = (inp[13]) ? 4'b1001 : node14347;
																assign node14347 = (inp[14]) ? 4'b1101 : 4'b1100;
														assign node14351 = (inp[12]) ? 4'b0001 : 4'b1001;
													assign node14354 = (inp[14]) ? node14360 : node14355;
														assign node14355 = (inp[13]) ? node14357 : 4'b0000;
															assign node14357 = (inp[10]) ? 4'b1000 : 4'b0000;
														assign node14360 = (inp[10]) ? node14364 : node14361;
															assign node14361 = (inp[13]) ? 4'b0001 : 4'b1100;
															assign node14364 = (inp[13]) ? node14366 : 4'b0001;
																assign node14366 = (inp[12]) ? 4'b0001 : 4'b1001;
											assign node14369 = (inp[0]) ? node14389 : node14370;
												assign node14370 = (inp[13]) ? node14376 : node14371;
													assign node14371 = (inp[10]) ? node14373 : 4'b1000;
														assign node14373 = (inp[2]) ? 4'b0000 : 4'b1000;
													assign node14376 = (inp[12]) ? node14384 : node14377;
														assign node14377 = (inp[10]) ? node14381 : node14378;
															assign node14378 = (inp[2]) ? 4'b0100 : 4'b1100;
															assign node14381 = (inp[2]) ? 4'b1100 : 4'b1000;
														assign node14384 = (inp[2]) ? node14386 : 4'b1100;
															assign node14386 = (inp[10]) ? 4'b1100 : 4'b1000;
												assign node14389 = (inp[10]) ? node14397 : node14390;
													assign node14390 = (inp[2]) ? node14392 : 4'b0000;
														assign node14392 = (inp[13]) ? 4'b0000 : node14393;
															assign node14393 = (inp[12]) ? 4'b1100 : 4'b0000;
													assign node14397 = (inp[13]) ? 4'b1000 : node14398;
														assign node14398 = (inp[2]) ? 4'b0000 : 4'b1000;
									assign node14402 = (inp[0]) ? node14510 : node14403;
										assign node14403 = (inp[13]) ? node14453 : node14404;
											assign node14404 = (inp[10]) ? node14428 : node14405;
												assign node14405 = (inp[1]) ? node14419 : node14406;
													assign node14406 = (inp[11]) ? node14412 : node14407;
														assign node14407 = (inp[2]) ? 4'b1101 : node14408;
															assign node14408 = (inp[14]) ? 4'b1101 : 4'b1100;
														assign node14412 = (inp[2]) ? node14416 : node14413;
															assign node14413 = (inp[12]) ? 4'b1101 : 4'b0101;
															assign node14416 = (inp[12]) ? 4'b1100 : 4'b0100;
													assign node14419 = (inp[11]) ? node14423 : node14420;
														assign node14420 = (inp[14]) ? 4'b0100 : 4'b0101;
														assign node14423 = (inp[2]) ? 4'b0100 : node14424;
															assign node14424 = (inp[12]) ? 4'b0100 : 4'b1100;
												assign node14428 = (inp[11]) ? node14444 : node14429;
													assign node14429 = (inp[2]) ? node14437 : node14430;
														assign node14430 = (inp[1]) ? 4'b0000 : node14431;
															assign node14431 = (inp[14]) ? 4'b0101 : node14432;
																assign node14432 = (inp[12]) ? 4'b1100 : 4'b0000;
														assign node14437 = (inp[1]) ? node14439 : 4'b0101;
															assign node14439 = (inp[12]) ? 4'b0101 : node14440;
																assign node14440 = (inp[14]) ? 4'b0000 : 4'b0001;
													assign node14444 = (inp[2]) ? node14448 : node14445;
														assign node14445 = (inp[1]) ? 4'b1000 : 4'b0000;
														assign node14448 = (inp[1]) ? 4'b0000 : node14449;
															assign node14449 = (inp[12]) ? 4'b0100 : 4'b1100;
											assign node14453 = (inp[2]) ? node14475 : node14454;
												assign node14454 = (inp[10]) ? node14464 : node14455;
													assign node14455 = (inp[1]) ? node14459 : node14456;
														assign node14456 = (inp[12]) ? 4'b1000 : 4'b0000;
														assign node14459 = (inp[12]) ? node14461 : 4'b1000;
															assign node14461 = (inp[11]) ? 4'b1000 : 4'b0000;
													assign node14464 = (inp[1]) ? node14470 : node14465;
														assign node14465 = (inp[11]) ? 4'b0100 : node14466;
															assign node14466 = (inp[12]) ? 4'b1000 : 4'b0100;
														assign node14470 = (inp[12]) ? node14472 : 4'b1100;
															assign node14472 = (inp[11]) ? 4'b1100 : 4'b0100;
												assign node14475 = (inp[1]) ? node14495 : node14476;
													assign node14476 = (inp[14]) ? node14486 : node14477;
														assign node14477 = (inp[11]) ? node14483 : node14478;
															assign node14478 = (inp[12]) ? 4'b0000 : node14479;
																assign node14479 = (inp[10]) ? 4'b0000 : 4'b1000;
															assign node14483 = (inp[12]) ? 4'b0001 : 4'b1001;
														assign node14486 = (inp[11]) ? node14492 : node14487;
															assign node14487 = (inp[12]) ? node14489 : 4'b0001;
																assign node14489 = (inp[10]) ? 4'b1001 : 4'b0001;
															assign node14492 = (inp[10]) ? 4'b0001 : 4'b1001;
													assign node14495 = (inp[14]) ? node14501 : node14496;
														assign node14496 = (inp[11]) ? node14498 : 4'b1001;
															assign node14498 = (inp[12]) ? 4'b1000 : 4'b0000;
														assign node14501 = (inp[11]) ? node14507 : node14502;
															assign node14502 = (inp[10]) ? node14504 : 4'b1000;
																assign node14504 = (inp[12]) ? 4'b0000 : 4'b1000;
															assign node14507 = (inp[10]) ? 4'b1000 : 4'b0000;
										assign node14510 = (inp[2]) ? 4'b1100 : node14511;
											assign node14511 = (inp[13]) ? node14545 : node14512;
												assign node14512 = (inp[10]) ? node14526 : node14513;
													assign node14513 = (inp[1]) ? node14519 : node14514;
														assign node14514 = (inp[14]) ? node14516 : 4'b1101;
															assign node14516 = (inp[11]) ? 4'b1101 : 4'b1100;
														assign node14519 = (inp[14]) ? node14523 : node14520;
															assign node14520 = (inp[12]) ? 4'b1100 : 4'b0100;
															assign node14523 = (inp[11]) ? 4'b1100 : 4'b1101;
													assign node14526 = (inp[12]) ? node14536 : node14527;
														assign node14527 = (inp[1]) ? node14531 : node14528;
															assign node14528 = (inp[14]) ? 4'b0100 : 4'b0101;
															assign node14531 = (inp[11]) ? 4'b0100 : node14532;
																assign node14532 = (inp[14]) ? 4'b0101 : 4'b0100;
														assign node14536 = (inp[1]) ? node14542 : node14537;
															assign node14537 = (inp[11]) ? 4'b1101 : node14538;
																assign node14538 = (inp[14]) ? 4'b1100 : 4'b1101;
															assign node14542 = (inp[14]) ? 4'b1101 : 4'b0100;
												assign node14545 = (inp[11]) ? node14565 : node14546;
													assign node14546 = (inp[10]) ? node14560 : node14547;
														assign node14547 = (inp[12]) ? node14553 : node14548;
															assign node14548 = (inp[1]) ? 4'b0001 : node14549;
																assign node14549 = (inp[14]) ? 4'b0100 : 4'b0101;
															assign node14553 = (inp[14]) ? node14557 : node14554;
																assign node14554 = (inp[1]) ? 4'b0100 : 4'b0101;
																assign node14557 = (inp[1]) ? 4'b0101 : 4'b0100;
														assign node14560 = (inp[12]) ? 4'b0001 : node14561;
															assign node14561 = (inp[1]) ? 4'b1001 : 4'b0001;
													assign node14565 = (inp[10]) ? node14571 : node14566;
														assign node14566 = (inp[1]) ? 4'b0000 : node14567;
															assign node14567 = (inp[12]) ? 4'b0101 : 4'b0000;
														assign node14571 = (inp[12]) ? node14573 : 4'b1000;
															assign node14573 = (inp[14]) ? 4'b1000 : 4'b0000;
								assign node14577 = (inp[11]) ? node14837 : node14578;
									assign node14578 = (inp[2]) ? node14694 : node14579;
										assign node14579 = (inp[10]) ? node14637 : node14580;
											assign node14580 = (inp[12]) ? node14608 : node14581;
												assign node14581 = (inp[0]) ? node14593 : node14582;
													assign node14582 = (inp[1]) ? node14588 : node14583;
														assign node14583 = (inp[14]) ? node14585 : 4'b0001;
															assign node14585 = (inp[13]) ? 4'b0001 : 4'b0000;
														assign node14588 = (inp[7]) ? 4'b1001 : node14589;
															assign node14589 = (inp[13]) ? 4'b1001 : 4'b1000;
													assign node14593 = (inp[1]) ? node14599 : node14594;
														assign node14594 = (inp[7]) ? 4'b1001 : node14595;
															assign node14595 = (inp[13]) ? 4'b0001 : 4'b1001;
														assign node14599 = (inp[13]) ? node14603 : node14600;
															assign node14600 = (inp[7]) ? 4'b0001 : 4'b0101;
															assign node14603 = (inp[7]) ? 4'b0101 : node14604;
																assign node14604 = (inp[14]) ? 4'b1000 : 4'b1001;
												assign node14608 = (inp[14]) ? node14626 : node14609;
													assign node14609 = (inp[13]) ? node14619 : node14610;
														assign node14610 = (inp[0]) ? 4'b1001 : node14611;
															assign node14611 = (inp[7]) ? node14615 : node14612;
																assign node14612 = (inp[1]) ? 4'b1000 : 4'b1001;
																assign node14615 = (inp[1]) ? 4'b1000 : 4'b1100;
														assign node14619 = (inp[0]) ? node14623 : node14620;
															assign node14620 = (inp[7]) ? 4'b0101 : 4'b1001;
															assign node14623 = (inp[7]) ? 4'b1001 : 4'b0000;
													assign node14626 = (inp[0]) ? node14630 : node14627;
														assign node14627 = (inp[13]) ? 4'b1001 : 4'b0001;
														assign node14630 = (inp[7]) ? 4'b1001 : node14631;
															assign node14631 = (inp[1]) ? 4'b1000 : node14632;
																assign node14632 = (inp[13]) ? 4'b0001 : 4'b1001;
											assign node14637 = (inp[13]) ? node14661 : node14638;
												assign node14638 = (inp[7]) ? node14650 : node14639;
													assign node14639 = (inp[1]) ? node14641 : 4'b0101;
														assign node14641 = (inp[12]) ? node14647 : node14642;
															assign node14642 = (inp[0]) ? node14644 : 4'b0001;
																assign node14644 = (inp[14]) ? 4'b0000 : 4'b0001;
															assign node14647 = (inp[0]) ? 4'b0101 : 4'b0001;
													assign node14650 = (inp[1]) ? node14652 : 4'b0001;
														assign node14652 = (inp[0]) ? node14658 : node14653;
															assign node14653 = (inp[14]) ? 4'b1001 : node14654;
																assign node14654 = (inp[12]) ? 4'b1000 : 4'b0100;
															assign node14658 = (inp[12]) ? 4'b0001 : 4'b1001;
												assign node14661 = (inp[12]) ? node14675 : node14662;
													assign node14662 = (inp[14]) ? node14670 : node14663;
														assign node14663 = (inp[1]) ? node14667 : node14664;
															assign node14664 = (inp[0]) ? 4'b0000 : 4'b1001;
															assign node14667 = (inp[0]) ? 4'b1001 : 4'b0001;
														assign node14670 = (inp[1]) ? node14672 : 4'b0001;
															assign node14672 = (inp[0]) ? 4'b1000 : 4'b0000;
													assign node14675 = (inp[0]) ? node14685 : node14676;
														assign node14676 = (inp[14]) ? node14682 : node14677;
															assign node14677 = (inp[7]) ? 4'b0001 : node14678;
																assign node14678 = (inp[1]) ? 4'b0001 : 4'b0000;
															assign node14682 = (inp[1]) ? 4'b0000 : 4'b0001;
														assign node14685 = (inp[14]) ? node14689 : node14686;
															assign node14686 = (inp[1]) ? 4'b0001 : 4'b0000;
															assign node14689 = (inp[7]) ? node14691 : 4'b1001;
																assign node14691 = (inp[1]) ? 4'b0000 : 4'b0101;
										assign node14694 = (inp[0]) ? node14766 : node14695;
											assign node14695 = (inp[1]) ? node14733 : node14696;
												assign node14696 = (inp[12]) ? node14718 : node14697;
													assign node14697 = (inp[13]) ? node14709 : node14698;
														assign node14698 = (inp[14]) ? node14704 : node14699;
															assign node14699 = (inp[7]) ? node14701 : 4'b0000;
																assign node14701 = (inp[10]) ? 4'b0000 : 4'b0100;
															assign node14704 = (inp[7]) ? node14706 : 4'b0000;
																assign node14706 = (inp[10]) ? 4'b0000 : 4'b1001;
														assign node14709 = (inp[7]) ? node14715 : node14710;
															assign node14710 = (inp[10]) ? node14712 : 4'b0100;
																assign node14712 = (inp[14]) ? 4'b1000 : 4'b1001;
															assign node14715 = (inp[10]) ? 4'b0100 : 4'b0000;
													assign node14718 = (inp[13]) ? node14726 : node14719;
														assign node14719 = (inp[14]) ? 4'b0101 : node14720;
															assign node14720 = (inp[7]) ? 4'b1000 : node14721;
																assign node14721 = (inp[10]) ? 4'b1000 : 4'b1100;
														assign node14726 = (inp[14]) ? 4'b1000 : node14727;
															assign node14727 = (inp[10]) ? node14729 : 4'b1000;
																assign node14729 = (inp[7]) ? 4'b1000 : 4'b1001;
												assign node14733 = (inp[12]) ? node14753 : node14734;
													assign node14734 = (inp[13]) ? node14742 : node14735;
														assign node14735 = (inp[7]) ? node14737 : 4'b1000;
															assign node14737 = (inp[10]) ? 4'b1000 : node14738;
																assign node14738 = (inp[14]) ? 4'b0100 : 4'b0101;
														assign node14742 = (inp[14]) ? node14748 : node14743;
															assign node14743 = (inp[7]) ? 4'b1000 : node14744;
																assign node14744 = (inp[10]) ? 4'b1000 : 4'b0000;
															assign node14748 = (inp[10]) ? 4'b0001 : node14749;
																assign node14749 = (inp[7]) ? 4'b1000 : 4'b0001;
													assign node14753 = (inp[10]) ? node14763 : node14754;
														assign node14754 = (inp[13]) ? node14758 : node14755;
															assign node14755 = (inp[7]) ? 4'b0101 : 4'b0000;
															assign node14758 = (inp[7]) ? 4'b0000 : node14759;
																assign node14759 = (inp[14]) ? 4'b0100 : 4'b0000;
														assign node14763 = (inp[13]) ? 4'b0001 : 4'b0000;
											assign node14766 = (inp[13]) ? node14804 : node14767;
												assign node14767 = (inp[7]) ? node14785 : node14768;
													assign node14768 = (inp[12]) ? node14780 : node14769;
														assign node14769 = (inp[10]) ? node14775 : node14770;
															assign node14770 = (inp[1]) ? 4'b0000 : node14771;
																assign node14771 = (inp[14]) ? 4'b1000 : 4'b1001;
															assign node14775 = (inp[1]) ? 4'b0001 : node14776;
																assign node14776 = (inp[14]) ? 4'b0000 : 4'b0001;
														assign node14780 = (inp[1]) ? 4'b1001 : node14781;
															assign node14781 = (inp[14]) ? 4'b1000 : 4'b1001;
													assign node14785 = (inp[10]) ? node14793 : node14786;
														assign node14786 = (inp[12]) ? 4'b1100 : node14787;
															assign node14787 = (inp[14]) ? 4'b1100 : node14788;
																assign node14788 = (inp[1]) ? 4'b0000 : 4'b1100;
														assign node14793 = (inp[12]) ? node14801 : node14794;
															assign node14794 = (inp[14]) ? node14798 : node14795;
																assign node14795 = (inp[1]) ? 4'b0000 : 4'b0001;
																assign node14798 = (inp[1]) ? 4'b0001 : 4'b0000;
															assign node14801 = (inp[14]) ? 4'b1100 : 4'b0000;
												assign node14804 = (inp[10]) ? node14822 : node14805;
													assign node14805 = (inp[7]) ? node14813 : node14806;
														assign node14806 = (inp[12]) ? node14808 : 4'b0001;
															assign node14808 = (inp[14]) ? 4'b0001 : node14809;
																assign node14809 = (inp[1]) ? 4'b0000 : 4'b0001;
														assign node14813 = (inp[1]) ? node14817 : node14814;
															assign node14814 = (inp[14]) ? 4'b0000 : 4'b0001;
															assign node14817 = (inp[14]) ? 4'b0001 : node14818;
																assign node14818 = (inp[12]) ? 4'b0000 : 4'b1000;
													assign node14822 = (inp[12]) ? node14830 : node14823;
														assign node14823 = (inp[14]) ? node14827 : node14824;
															assign node14824 = (inp[1]) ? 4'b1000 : 4'b1001;
															assign node14827 = (inp[1]) ? 4'b1001 : 4'b1000;
														assign node14830 = (inp[14]) ? node14834 : node14831;
															assign node14831 = (inp[1]) ? 4'b1000 : 4'b0001;
															assign node14834 = (inp[1]) ? 4'b0001 : 4'b0000;
									assign node14837 = (inp[1]) ? node14915 : node14838;
										assign node14838 = (inp[0]) ? node14876 : node14839;
											assign node14839 = (inp[13]) ? node14855 : node14840;
												assign node14840 = (inp[2]) ? node14848 : node14841;
													assign node14841 = (inp[10]) ? node14843 : 4'b0001;
														assign node14843 = (inp[12]) ? node14845 : 4'b0000;
															assign node14845 = (inp[7]) ? 4'b0001 : 4'b0101;
													assign node14848 = (inp[7]) ? node14850 : 4'b0000;
														assign node14850 = (inp[10]) ? 4'b0000 : node14851;
															assign node14851 = (inp[12]) ? 4'b1001 : 4'b0101;
												assign node14855 = (inp[10]) ? node14863 : node14856;
													assign node14856 = (inp[2]) ? node14860 : node14857;
														assign node14857 = (inp[12]) ? 4'b0000 : 4'b1000;
														assign node14860 = (inp[7]) ? 4'b0000 : 4'b0100;
													assign node14863 = (inp[7]) ? node14869 : node14864;
														assign node14864 = (inp[12]) ? 4'b1001 : node14865;
															assign node14865 = (inp[2]) ? 4'b0001 : 4'b1001;
														assign node14869 = (inp[12]) ? node14873 : node14870;
															assign node14870 = (inp[2]) ? 4'b0001 : 4'b0100;
															assign node14873 = (inp[2]) ? 4'b0100 : 4'b1000;
											assign node14876 = (inp[13]) ? node14902 : node14877;
												assign node14877 = (inp[2]) ? node14891 : node14878;
													assign node14878 = (inp[7]) ? node14884 : node14879;
														assign node14879 = (inp[10]) ? 4'b0100 : node14880;
															assign node14880 = (inp[12]) ? 4'b1000 : 4'b0100;
														assign node14884 = (inp[10]) ? node14888 : node14885;
															assign node14885 = (inp[12]) ? 4'b1000 : 4'b0000;
															assign node14888 = (inp[12]) ? 4'b0000 : 4'b1000;
													assign node14891 = (inp[7]) ? node14897 : node14892;
														assign node14892 = (inp[10]) ? node14894 : 4'b1001;
															assign node14894 = (inp[12]) ? 4'b1001 : 4'b0001;
														assign node14897 = (inp[10]) ? node14899 : 4'b1100;
															assign node14899 = (inp[12]) ? 4'b1100 : 4'b0001;
												assign node14902 = (inp[2]) ? node14910 : node14903;
													assign node14903 = (inp[10]) ? 4'b0001 : node14904;
														assign node14904 = (inp[7]) ? node14906 : 4'b1001;
															assign node14906 = (inp[14]) ? 4'b1000 : 4'b0100;
													assign node14910 = (inp[10]) ? node14912 : 4'b0001;
														assign node14912 = (inp[12]) ? 4'b0001 : 4'b1001;
										assign node14915 = (inp[10]) ? node14961 : node14916;
											assign node14916 = (inp[2]) ? node14938 : node14917;
												assign node14917 = (inp[12]) ? node14923 : node14918;
													assign node14918 = (inp[7]) ? 4'b0000 : node14919;
														assign node14919 = (inp[13]) ? 4'b0000 : 4'b0100;
													assign node14923 = (inp[0]) ? node14929 : node14924;
														assign node14924 = (inp[13]) ? node14926 : 4'b1000;
															assign node14926 = (inp[7]) ? 4'b0000 : 4'b0100;
														assign node14929 = (inp[14]) ? 4'b0100 : node14930;
															assign node14930 = (inp[7]) ? node14934 : node14931;
																assign node14931 = (inp[13]) ? 4'b1000 : 4'b0100;
																assign node14934 = (inp[13]) ? 4'b0100 : 4'b0000;
												assign node14938 = (inp[7]) ? node14948 : node14939;
													assign node14939 = (inp[13]) ? node14945 : node14940;
														assign node14940 = (inp[12]) ? 4'b1000 : node14941;
															assign node14941 = (inp[0]) ? 4'b0000 : 4'b1000;
														assign node14945 = (inp[12]) ? 4'b0000 : 4'b1000;
													assign node14948 = (inp[13]) ? node14956 : node14949;
														assign node14949 = (inp[12]) ? node14953 : node14950;
															assign node14950 = (inp[0]) ? 4'b0000 : 4'b1100;
															assign node14953 = (inp[0]) ? 4'b1100 : 4'b0100;
														assign node14956 = (inp[0]) ? node14958 : 4'b1000;
															assign node14958 = (inp[12]) ? 4'b0000 : 4'b1000;
											assign node14961 = (inp[13]) ? 4'b1000 : node14962;
												assign node14962 = (inp[0]) ? node14968 : node14963;
													assign node14963 = (inp[7]) ? node14965 : 4'b1000;
														assign node14965 = (inp[2]) ? 4'b1000 : 4'b0100;
													assign node14968 = (inp[7]) ? node14970 : 4'b0000;
														assign node14970 = (inp[2]) ? 4'b0000 : 4'b1000;
							assign node14974 = (inp[4]) ? node15408 : node14975;
								assign node14975 = (inp[11]) ? node15239 : node14976;
									assign node14976 = (inp[2]) ? node15106 : node14977;
										assign node14977 = (inp[10]) ? node15037 : node14978;
											assign node14978 = (inp[1]) ? node15014 : node14979;
												assign node14979 = (inp[0]) ? node14995 : node14980;
													assign node14980 = (inp[14]) ? node14986 : node14981;
														assign node14981 = (inp[13]) ? node14983 : 4'b0000;
															assign node14983 = (inp[7]) ? 4'b0001 : 4'b0000;
														assign node14986 = (inp[7]) ? node14990 : node14987;
															assign node14987 = (inp[13]) ? 4'b0001 : 4'b0000;
															assign node14990 = (inp[13]) ? 4'b0001 : node14991;
																assign node14991 = (inp[12]) ? 4'b1001 : 4'b0001;
													assign node14995 = (inp[12]) ? node15007 : node14996;
														assign node14996 = (inp[14]) ? node15002 : node14997;
															assign node14997 = (inp[7]) ? 4'b0000 : node14998;
																assign node14998 = (inp[13]) ? 4'b1001 : 4'b0000;
															assign node15002 = (inp[7]) ? node15004 : 4'b0000;
																assign node15004 = (inp[13]) ? 4'b0000 : 4'b1001;
														assign node15007 = (inp[7]) ? node15011 : node15008;
															assign node15008 = (inp[14]) ? 4'b0000 : 4'b1000;
															assign node15011 = (inp[13]) ? 4'b1000 : 4'b1001;
												assign node15014 = (inp[14]) ? node15028 : node15015;
													assign node15015 = (inp[7]) ? node15021 : node15016;
														assign node15016 = (inp[12]) ? node15018 : 4'b0000;
															assign node15018 = (inp[13]) ? 4'b0001 : 4'b0000;
														assign node15021 = (inp[0]) ? node15025 : node15022;
															assign node15022 = (inp[13]) ? 4'b0001 : 4'b0000;
															assign node15025 = (inp[13]) ? 4'b0000 : 4'b0001;
													assign node15028 = (inp[0]) ? node15030 : 4'b0000;
														assign node15030 = (inp[7]) ? 4'b0000 : node15031;
															assign node15031 = (inp[13]) ? node15033 : 4'b0000;
																assign node15033 = (inp[12]) ? 4'b1001 : 4'b0001;
											assign node15037 = (inp[13]) ? node15079 : node15038;
												assign node15038 = (inp[0]) ? node15054 : node15039;
													assign node15039 = (inp[1]) ? node15049 : node15040;
														assign node15040 = (inp[7]) ? 4'b0000 : node15041;
															assign node15041 = (inp[12]) ? node15045 : node15042;
																assign node15042 = (inp[14]) ? 4'b1000 : 4'b1001;
																assign node15045 = (inp[14]) ? 4'b0000 : 4'b0001;
														assign node15049 = (inp[14]) ? node15051 : 4'b1000;
															assign node15051 = (inp[7]) ? 4'b1001 : 4'b0001;
													assign node15054 = (inp[14]) ? node15064 : node15055;
														assign node15055 = (inp[7]) ? node15059 : node15056;
															assign node15056 = (inp[1]) ? 4'b0000 : 4'b1000;
															assign node15059 = (inp[1]) ? 4'b1000 : node15060;
																assign node15060 = (inp[12]) ? 4'b1000 : 4'b0000;
														assign node15064 = (inp[7]) ? node15072 : node15065;
															assign node15065 = (inp[1]) ? node15069 : node15066;
																assign node15066 = (inp[12]) ? 4'b1000 : 4'b0000;
																assign node15069 = (inp[12]) ? 4'b0000 : 4'b1000;
															assign node15072 = (inp[1]) ? node15076 : node15073;
																assign node15073 = (inp[12]) ? 4'b0001 : 4'b0000;
																assign node15076 = (inp[12]) ? 4'b0000 : 4'b1000;
												assign node15079 = (inp[1]) ? node15095 : node15080;
													assign node15080 = (inp[0]) ? node15088 : node15081;
														assign node15081 = (inp[7]) ? node15085 : node15082;
															assign node15082 = (inp[14]) ? 4'b0000 : 4'b0001;
															assign node15085 = (inp[12]) ? 4'b0000 : 4'b1000;
														assign node15088 = (inp[7]) ? node15092 : node15089;
															assign node15089 = (inp[12]) ? 4'b0001 : 4'b1001;
															assign node15092 = (inp[14]) ? 4'b1000 : 4'b1001;
													assign node15095 = (inp[0]) ? node15101 : node15096;
														assign node15096 = (inp[7]) ? node15098 : 4'b1001;
															assign node15098 = (inp[14]) ? 4'b1001 : 4'b1000;
														assign node15101 = (inp[7]) ? 4'b0001 : node15102;
															assign node15102 = (inp[14]) ? 4'b0000 : 4'b0001;
										assign node15106 = (inp[13]) ? node15186 : node15107;
											assign node15107 = (inp[10]) ? node15143 : node15108;
												assign node15108 = (inp[12]) ? node15130 : node15109;
													assign node15109 = (inp[7]) ? node15119 : node15110;
														assign node15110 = (inp[0]) ? node15114 : node15111;
															assign node15111 = (inp[1]) ? 4'b1001 : 4'b0001;
															assign node15114 = (inp[1]) ? 4'b0001 : node15115;
																assign node15115 = (inp[14]) ? 4'b1000 : 4'b1001;
														assign node15119 = (inp[1]) ? node15125 : node15120;
															assign node15120 = (inp[14]) ? 4'b0000 : node15121;
																assign node15121 = (inp[0]) ? 4'b1001 : 4'b0001;
															assign node15125 = (inp[14]) ? 4'b1001 : node15126;
																assign node15126 = (inp[0]) ? 4'b0000 : 4'b1000;
													assign node15130 = (inp[14]) ? node15138 : node15131;
														assign node15131 = (inp[1]) ? node15133 : 4'b1001;
															assign node15133 = (inp[7]) ? 4'b1000 : node15134;
																assign node15134 = (inp[0]) ? 4'b1000 : 4'b1001;
														assign node15138 = (inp[1]) ? node15140 : 4'b1000;
															assign node15140 = (inp[0]) ? 4'b1001 : 4'b0001;
												assign node15143 = (inp[14]) ? node15163 : node15144;
													assign node15144 = (inp[7]) ? node15154 : node15145;
														assign node15145 = (inp[12]) ? node15149 : node15146;
															assign node15146 = (inp[0]) ? 4'b0001 : 4'b0000;
															assign node15149 = (inp[1]) ? node15151 : 4'b0001;
																assign node15151 = (inp[0]) ? 4'b0001 : 4'b1001;
														assign node15154 = (inp[1]) ? 4'b0001 : node15155;
															assign node15155 = (inp[12]) ? node15159 : node15156;
																assign node15156 = (inp[0]) ? 4'b0001 : 4'b1001;
																assign node15159 = (inp[0]) ? 4'b1001 : 4'b0001;
													assign node15163 = (inp[12]) ? node15177 : node15164;
														assign node15164 = (inp[0]) ? node15172 : node15165;
															assign node15165 = (inp[7]) ? node15169 : node15166;
																assign node15166 = (inp[1]) ? 4'b1000 : 4'b1001;
																assign node15169 = (inp[1]) ? 4'b0001 : 4'b1001;
															assign node15172 = (inp[7]) ? 4'b0001 : node15173;
																assign node15173 = (inp[1]) ? 4'b1001 : 4'b0001;
														assign node15177 = (inp[7]) ? node15183 : node15178;
															assign node15178 = (inp[1]) ? node15180 : 4'b0001;
																assign node15180 = (inp[0]) ? 4'b0001 : 4'b1000;
															assign node15183 = (inp[0]) ? 4'b1000 : 4'b0001;
											assign node15186 = (inp[0]) ? node15208 : node15187;
												assign node15187 = (inp[10]) ? node15197 : node15188;
													assign node15188 = (inp[1]) ? 4'b0000 : node15189;
														assign node15189 = (inp[7]) ? node15191 : 4'b0000;
															assign node15191 = (inp[14]) ? node15193 : 4'b1000;
																assign node15193 = (inp[12]) ? 4'b0001 : 4'b1001;
													assign node15197 = (inp[14]) ? node15201 : node15198;
														assign node15198 = (inp[12]) ? 4'b1001 : 4'b0001;
														assign node15201 = (inp[12]) ? node15203 : 4'b0000;
															assign node15203 = (inp[7]) ? 4'b0000 : node15204;
																assign node15204 = (inp[1]) ? 4'b1001 : 4'b1000;
												assign node15208 = (inp[7]) ? node15226 : node15209;
													assign node15209 = (inp[10]) ? node15215 : node15210;
														assign node15210 = (inp[12]) ? 4'b1001 : node15211;
															assign node15211 = (inp[1]) ? 4'b0001 : 4'b1001;
														assign node15215 = (inp[1]) ? node15219 : node15216;
															assign node15216 = (inp[14]) ? 4'b0001 : 4'b0000;
															assign node15219 = (inp[14]) ? node15223 : node15220;
																assign node15220 = (inp[12]) ? 4'b0001 : 4'b1001;
																assign node15223 = (inp[12]) ? 4'b0000 : 4'b1000;
													assign node15226 = (inp[10]) ? node15234 : node15227;
														assign node15227 = (inp[14]) ? node15231 : node15228;
															assign node15228 = (inp[1]) ? 4'b0000 : 4'b0001;
															assign node15231 = (inp[1]) ? 4'b0001 : 4'b0000;
														assign node15234 = (inp[1]) ? node15236 : 4'b0001;
															assign node15236 = (inp[12]) ? 4'b0001 : 4'b1001;
									assign node15239 = (inp[1]) ? node15347 : node15240;
										assign node15240 = (inp[7]) ? node15296 : node15241;
											assign node15241 = (inp[0]) ? node15271 : node15242;
												assign node15242 = (inp[2]) ? node15258 : node15243;
													assign node15243 = (inp[13]) ? node15247 : node15244;
														assign node15244 = (inp[10]) ? 4'b1001 : 4'b1000;
														assign node15247 = (inp[14]) ? node15253 : node15248;
															assign node15248 = (inp[12]) ? node15250 : 4'b1001;
																assign node15250 = (inp[10]) ? 4'b1001 : 4'b0001;
															assign node15253 = (inp[10]) ? 4'b0000 : node15254;
																assign node15254 = (inp[12]) ? 4'b0001 : 4'b1001;
													assign node15258 = (inp[12]) ? node15264 : node15259;
														assign node15259 = (inp[13]) ? 4'b1000 : node15260;
															assign node15260 = (inp[10]) ? 4'b0001 : 4'b1000;
														assign node15264 = (inp[10]) ? node15268 : node15265;
															assign node15265 = (inp[13]) ? 4'b1000 : 4'b0000;
															assign node15268 = (inp[13]) ? 4'b0000 : 4'b0001;
												assign node15271 = (inp[13]) ? node15281 : node15272;
													assign node15272 = (inp[2]) ? node15274 : 4'b0000;
														assign node15274 = (inp[12]) ? node15278 : node15275;
															assign node15275 = (inp[10]) ? 4'b1000 : 4'b0000;
															assign node15278 = (inp[10]) ? 4'b0000 : 4'b1001;
													assign node15281 = (inp[12]) ? node15289 : node15282;
														assign node15282 = (inp[10]) ? node15286 : node15283;
															assign node15283 = (inp[2]) ? 4'b0000 : 4'b1001;
															assign node15286 = (inp[2]) ? 4'b0001 : 4'b0000;
														assign node15289 = (inp[2]) ? node15293 : node15290;
															assign node15290 = (inp[10]) ? 4'b1000 : 4'b1001;
															assign node15293 = (inp[10]) ? 4'b0001 : 4'b1000;
											assign node15296 = (inp[13]) ? node15320 : node15297;
												assign node15297 = (inp[10]) ? node15307 : node15298;
													assign node15298 = (inp[0]) ? node15304 : node15299;
														assign node15299 = (inp[12]) ? 4'b0001 : node15300;
															assign node15300 = (inp[2]) ? 4'b0001 : 4'b1001;
														assign node15304 = (inp[2]) ? 4'b1001 : 4'b0001;
													assign node15307 = (inp[12]) ? node15315 : node15308;
														assign node15308 = (inp[2]) ? node15312 : node15309;
															assign node15309 = (inp[0]) ? 4'b0000 : 4'b0001;
															assign node15312 = (inp[0]) ? 4'b0001 : 4'b0000;
														assign node15315 = (inp[0]) ? node15317 : 4'b1000;
															assign node15317 = (inp[2]) ? 4'b1001 : 4'b0000;
												assign node15320 = (inp[2]) ? node15334 : node15321;
													assign node15321 = (inp[10]) ? node15327 : node15322;
														assign node15322 = (inp[12]) ? node15324 : 4'b0000;
															assign node15324 = (inp[0]) ? 4'b0000 : 4'b1000;
														assign node15327 = (inp[0]) ? node15331 : node15328;
															assign node15328 = (inp[12]) ? 4'b0000 : 4'b0001;
															assign node15331 = (inp[12]) ? 4'b1001 : 4'b0000;
													assign node15334 = (inp[0]) ? node15340 : node15335;
														assign node15335 = (inp[10]) ? node15337 : 4'b0001;
															assign node15337 = (inp[12]) ? 4'b0001 : 4'b1001;
														assign node15340 = (inp[10]) ? node15344 : node15341;
															assign node15341 = (inp[12]) ? 4'b0001 : 4'b0000;
															assign node15344 = (inp[12]) ? 4'b0000 : 4'b1000;
										assign node15347 = (inp[13]) ? node15385 : node15348;
											assign node15348 = (inp[2]) ? node15372 : node15349;
												assign node15349 = (inp[10]) ? node15365 : node15350;
													assign node15350 = (inp[14]) ? node15358 : node15351;
														assign node15351 = (inp[12]) ? 4'b1000 : node15352;
															assign node15352 = (inp[7]) ? 4'b1000 : node15353;
																assign node15353 = (inp[0]) ? 4'b1000 : 4'b0000;
														assign node15358 = (inp[12]) ? node15362 : node15359;
															assign node15359 = (inp[0]) ? 4'b1000 : 4'b0000;
															assign node15362 = (inp[0]) ? 4'b0000 : 4'b1000;
													assign node15365 = (inp[0]) ? node15369 : node15366;
														assign node15366 = (inp[7]) ? 4'b0000 : 4'b1000;
														assign node15369 = (inp[7]) ? 4'b1000 : 4'b0000;
												assign node15372 = (inp[0]) ? node15374 : 4'b0000;
													assign node15374 = (inp[14]) ? node15376 : 4'b0000;
														assign node15376 = (inp[10]) ? node15382 : node15377;
															assign node15377 = (inp[12]) ? node15379 : 4'b0000;
																assign node15379 = (inp[7]) ? 4'b1000 : 4'b0000;
															assign node15382 = (inp[7]) ? 4'b0000 : 4'b1000;
											assign node15385 = (inp[10]) ? 4'b1000 : node15386;
												assign node15386 = (inp[0]) ? node15398 : node15387;
													assign node15387 = (inp[7]) ? node15393 : node15388;
														assign node15388 = (inp[2]) ? node15390 : 4'b1000;
															assign node15390 = (inp[12]) ? 4'b0000 : 4'b1000;
														assign node15393 = (inp[2]) ? 4'b1000 : node15394;
															assign node15394 = (inp[12]) ? 4'b1000 : 4'b0000;
													assign node15398 = (inp[14]) ? 4'b0000 : node15399;
														assign node15399 = (inp[7]) ? node15401 : 4'b0000;
															assign node15401 = (inp[2]) ? 4'b0000 : node15402;
																assign node15402 = (inp[12]) ? 4'b0000 : 4'b1000;
								assign node15408 = (inp[13]) ? node15616 : node15409;
									assign node15409 = (inp[11]) ? node15531 : node15410;
										assign node15410 = (inp[1]) ? node15472 : node15411;
											assign node15411 = (inp[10]) ? node15439 : node15412;
												assign node15412 = (inp[14]) ? node15424 : node15413;
													assign node15413 = (inp[0]) ? node15419 : node15414;
														assign node15414 = (inp[12]) ? node15416 : 4'b1000;
															assign node15416 = (inp[2]) ? 4'b0000 : 4'b1000;
														assign node15419 = (inp[2]) ? node15421 : 4'b0000;
															assign node15421 = (inp[7]) ? 4'b0000 : 4'b1000;
													assign node15424 = (inp[7]) ? node15434 : node15425;
														assign node15425 = (inp[0]) ? node15431 : node15426;
															assign node15426 = (inp[12]) ? node15428 : 4'b1000;
																assign node15428 = (inp[2]) ? 4'b0000 : 4'b1000;
															assign node15431 = (inp[2]) ? 4'b1001 : 4'b0000;
														assign node15434 = (inp[2]) ? node15436 : 4'b0001;
															assign node15436 = (inp[0]) ? 4'b1001 : 4'b0001;
												assign node15439 = (inp[2]) ? node15457 : node15440;
													assign node15440 = (inp[14]) ? node15448 : node15441;
														assign node15441 = (inp[7]) ? node15443 : 4'b0000;
															assign node15443 = (inp[0]) ? node15445 : 4'b0001;
																assign node15445 = (inp[12]) ? 4'b0001 : 4'b1001;
														assign node15448 = (inp[7]) ? 4'b0000 : node15449;
															assign node15449 = (inp[0]) ? node15453 : node15450;
																assign node15450 = (inp[12]) ? 4'b0001 : 4'b1001;
																assign node15453 = (inp[12]) ? 4'b1001 : 4'b0001;
													assign node15457 = (inp[12]) ? node15461 : node15458;
														assign node15458 = (inp[14]) ? 4'b0000 : 4'b0001;
														assign node15461 = (inp[7]) ? node15467 : node15462;
															assign node15462 = (inp[0]) ? node15464 : 4'b1000;
																assign node15464 = (inp[14]) ? 4'b0000 : 4'b0001;
															assign node15467 = (inp[14]) ? 4'b0001 : node15468;
																assign node15468 = (inp[0]) ? 4'b1000 : 4'b0000;
											assign node15472 = (inp[7]) ? node15498 : node15473;
												assign node15473 = (inp[0]) ? node15485 : node15474;
													assign node15474 = (inp[10]) ? node15480 : node15475;
														assign node15475 = (inp[2]) ? 4'b0001 : node15476;
															assign node15476 = (inp[14]) ? 4'b0000 : 4'b0001;
														assign node15480 = (inp[2]) ? 4'b0000 : node15481;
															assign node15481 = (inp[12]) ? 4'b0001 : 4'b0000;
													assign node15485 = (inp[14]) ? node15493 : node15486;
														assign node15486 = (inp[2]) ? node15490 : node15487;
															assign node15487 = (inp[12]) ? 4'b0000 : 4'b1000;
															assign node15490 = (inp[10]) ? 4'b0001 : 4'b0000;
														assign node15493 = (inp[2]) ? node15495 : 4'b0001;
															assign node15495 = (inp[10]) ? 4'b0001 : 4'b1000;
												assign node15498 = (inp[0]) ? node15518 : node15499;
													assign node15499 = (inp[12]) ? node15507 : node15500;
														assign node15500 = (inp[2]) ? node15502 : 4'b0001;
															assign node15502 = (inp[10]) ? 4'b0000 : node15503;
																assign node15503 = (inp[14]) ? 4'b0001 : 4'b0000;
														assign node15507 = (inp[10]) ? node15513 : node15508;
															assign node15508 = (inp[2]) ? node15510 : 4'b1000;
																assign node15510 = (inp[14]) ? 4'b1000 : 4'b0000;
															assign node15513 = (inp[2]) ? 4'b0001 : node15514;
																assign node15514 = (inp[14]) ? 4'b0001 : 4'b1000;
													assign node15518 = (inp[10]) ? node15524 : node15519;
														assign node15519 = (inp[2]) ? node15521 : 4'b0000;
															assign node15521 = (inp[14]) ? 4'b0000 : 4'b0001;
														assign node15524 = (inp[12]) ? 4'b0000 : node15525;
															assign node15525 = (inp[2]) ? node15527 : 4'b0000;
																assign node15527 = (inp[14]) ? 4'b1000 : 4'b0000;
										assign node15531 = (inp[1]) ? node15581 : node15532;
											assign node15532 = (inp[2]) ? node15558 : node15533;
												assign node15533 = (inp[10]) ? node15549 : node15534;
													assign node15534 = (inp[12]) ? node15542 : node15535;
														assign node15535 = (inp[0]) ? node15539 : node15536;
															assign node15536 = (inp[7]) ? 4'b1000 : 4'b0000;
															assign node15539 = (inp[7]) ? 4'b1001 : 4'b1000;
														assign node15542 = (inp[7]) ? node15546 : node15543;
															assign node15543 = (inp[0]) ? 4'b1000 : 4'b1001;
															assign node15546 = (inp[0]) ? 4'b0001 : 4'b1000;
													assign node15549 = (inp[0]) ? node15553 : node15550;
														assign node15550 = (inp[7]) ? 4'b0001 : 4'b1000;
														assign node15553 = (inp[12]) ? 4'b0000 : node15554;
															assign node15554 = (inp[14]) ? 4'b1000 : 4'b0000;
												assign node15558 = (inp[10]) ? node15568 : node15559;
													assign node15559 = (inp[0]) ? node15563 : node15560;
														assign node15560 = (inp[7]) ? 4'b0000 : 4'b0001;
														assign node15563 = (inp[7]) ? node15565 : 4'b0000;
															assign node15565 = (inp[12]) ? 4'b1000 : 4'b0001;
													assign node15568 = (inp[0]) ? node15574 : node15569;
														assign node15569 = (inp[14]) ? 4'b1000 : node15570;
															assign node15570 = (inp[12]) ? 4'b0000 : 4'b1000;
														assign node15574 = (inp[14]) ? node15576 : 4'b0000;
															assign node15576 = (inp[7]) ? 4'b0000 : node15577;
																assign node15577 = (inp[12]) ? 4'b0001 : 4'b0000;
											assign node15581 = (inp[10]) ? 4'b0000 : node15582;
												assign node15582 = (inp[2]) ? node15602 : node15583;
													assign node15583 = (inp[12]) ? node15589 : node15584;
														assign node15584 = (inp[0]) ? 4'b0000 : node15585;
															assign node15585 = (inp[7]) ? 4'b1000 : 4'b0000;
														assign node15589 = (inp[14]) ? node15597 : node15590;
															assign node15590 = (inp[0]) ? node15594 : node15591;
																assign node15591 = (inp[7]) ? 4'b0000 : 4'b1000;
																assign node15594 = (inp[7]) ? 4'b1000 : 4'b0000;
															assign node15597 = (inp[0]) ? 4'b0000 : node15598;
																assign node15598 = (inp[7]) ? 4'b0000 : 4'b1000;
													assign node15602 = (inp[7]) ? node15610 : node15603;
														assign node15603 = (inp[12]) ? node15607 : node15604;
															assign node15604 = (inp[0]) ? 4'b0000 : 4'b1000;
															assign node15607 = (inp[0]) ? 4'b1000 : 4'b0000;
														assign node15610 = (inp[0]) ? node15612 : 4'b0000;
															assign node15612 = (inp[12]) ? 4'b0000 : 4'b1000;
									assign node15616 = (inp[10]) ? node15700 : node15617;
										assign node15617 = (inp[1]) ? node15669 : node15618;
											assign node15618 = (inp[12]) ? node15638 : node15619;
												assign node15619 = (inp[7]) ? node15625 : node15620;
													assign node15620 = (inp[0]) ? 4'b0000 : node15621;
														assign node15621 = (inp[2]) ? 4'b0001 : 4'b0000;
													assign node15625 = (inp[0]) ? node15631 : node15626;
														assign node15626 = (inp[2]) ? 4'b0000 : node15627;
															assign node15627 = (inp[11]) ? 4'b0001 : 4'b0000;
														assign node15631 = (inp[2]) ? 4'b0001 : node15632;
															assign node15632 = (inp[14]) ? node15634 : 4'b0000;
																assign node15634 = (inp[11]) ? 4'b0000 : 4'b0001;
												assign node15638 = (inp[7]) ? node15658 : node15639;
													assign node15639 = (inp[0]) ? node15649 : node15640;
														assign node15640 = (inp[14]) ? 4'b0001 : node15641;
															assign node15641 = (inp[2]) ? node15645 : node15642;
																assign node15642 = (inp[11]) ? 4'b0001 : 4'b0000;
																assign node15645 = (inp[11]) ? 4'b0000 : 4'b0001;
														assign node15649 = (inp[2]) ? node15655 : node15650;
															assign node15650 = (inp[14]) ? 4'b0000 : node15651;
																assign node15651 = (inp[11]) ? 4'b0000 : 4'b0001;
															assign node15655 = (inp[11]) ? 4'b0001 : 4'b0000;
													assign node15658 = (inp[0]) ? node15660 : 4'b0000;
														assign node15660 = (inp[14]) ? 4'b0001 : node15661;
															assign node15661 = (inp[11]) ? node15665 : node15662;
																assign node15662 = (inp[2]) ? 4'b0001 : 4'b0000;
																assign node15665 = (inp[2]) ? 4'b0000 : 4'b0001;
											assign node15669 = (inp[11]) ? 4'b0000 : node15670;
												assign node15670 = (inp[0]) ? node15688 : node15671;
													assign node15671 = (inp[12]) ? node15681 : node15672;
														assign node15672 = (inp[14]) ? node15678 : node15673;
															assign node15673 = (inp[7]) ? 4'b0001 : node15674;
																assign node15674 = (inp[2]) ? 4'b0000 : 4'b0001;
															assign node15678 = (inp[7]) ? 4'b0000 : 4'b0001;
														assign node15681 = (inp[14]) ? node15683 : 4'b0000;
															assign node15683 = (inp[2]) ? node15685 : 4'b0001;
																assign node15685 = (inp[7]) ? 4'b0001 : 4'b0000;
													assign node15688 = (inp[7]) ? node15694 : node15689;
														assign node15689 = (inp[2]) ? node15691 : 4'b0000;
															assign node15691 = (inp[14]) ? 4'b0000 : 4'b0001;
														assign node15694 = (inp[12]) ? 4'b0000 : node15695;
															assign node15695 = (inp[2]) ? 4'b0000 : 4'b0001;
										assign node15700 = (inp[11]) ? 4'b0000 : node15701;
											assign node15701 = (inp[1]) ? 4'b0000 : node15702;
												assign node15702 = (inp[2]) ? node15722 : node15703;
													assign node15703 = (inp[14]) ? node15711 : node15704;
														assign node15704 = (inp[7]) ? 4'b0000 : node15705;
															assign node15705 = (inp[0]) ? node15707 : 4'b0000;
																assign node15707 = (inp[12]) ? 4'b0000 : 4'b0001;
														assign node15711 = (inp[7]) ? node15717 : node15712;
															assign node15712 = (inp[12]) ? node15714 : 4'b0000;
																assign node15714 = (inp[0]) ? 4'b0000 : 4'b0001;
															assign node15717 = (inp[12]) ? node15719 : 4'b0001;
																assign node15719 = (inp[0]) ? 4'b0001 : 4'b0000;
													assign node15722 = (inp[12]) ? node15730 : node15723;
														assign node15723 = (inp[0]) ? 4'b0000 : node15724;
															assign node15724 = (inp[14]) ? node15726 : 4'b0001;
																assign node15726 = (inp[7]) ? 4'b0000 : 4'b0001;
														assign node15730 = (inp[0]) ? node15736 : node15731;
															assign node15731 = (inp[14]) ? 4'b0000 : node15732;
																assign node15732 = (inp[7]) ? 4'b0000 : 4'b0001;
															assign node15736 = (inp[7]) ? 4'b0001 : node15737;
																assign node15737 = (inp[14]) ? 4'b0001 : 4'b0000;
				assign node15743 = (inp[0]) ? node17915 : node15744;
					assign node15744 = (inp[6]) ? node16352 : node15745;
						assign node15745 = (inp[5]) ? node15881 : node15746;
							assign node15746 = (inp[3]) ? node15748 : 4'b1010;
								assign node15748 = (inp[2]) ? 4'b1010 : node15749;
									assign node15749 = (inp[4]) ? node15801 : node15750;
										assign node15750 = (inp[7]) ? 4'b1010 : node15751;
											assign node15751 = (inp[13]) ? node15775 : node15752;
												assign node15752 = (inp[12]) ? node15766 : node15753;
													assign node15753 = (inp[10]) ? node15757 : node15754;
														assign node15754 = (inp[1]) ? 4'b0000 : 4'b1010;
														assign node15757 = (inp[1]) ? node15761 : node15758;
															assign node15758 = (inp[11]) ? 4'b0001 : 4'b0000;
															assign node15761 = (inp[11]) ? 4'b0000 : node15762;
																assign node15762 = (inp[14]) ? 4'b0001 : 4'b0000;
													assign node15766 = (inp[10]) ? node15768 : 4'b1010;
														assign node15768 = (inp[1]) ? node15770 : 4'b1010;
															assign node15770 = (inp[11]) ? 4'b0000 : node15771;
																assign node15771 = (inp[14]) ? 4'b1010 : 4'b0000;
												assign node15775 = (inp[1]) ? node15783 : node15776;
													assign node15776 = (inp[11]) ? node15780 : node15777;
														assign node15777 = (inp[14]) ? 4'b0000 : 4'b0001;
														assign node15780 = (inp[12]) ? 4'b0001 : 4'b1001;
													assign node15783 = (inp[10]) ? node15795 : node15784;
														assign node15784 = (inp[12]) ? node15790 : node15785;
															assign node15785 = (inp[11]) ? 4'b1000 : node15786;
																assign node15786 = (inp[14]) ? 4'b0001 : 4'b1000;
															assign node15790 = (inp[11]) ? 4'b0000 : node15791;
																assign node15791 = (inp[14]) ? 4'b0001 : 4'b0000;
														assign node15795 = (inp[11]) ? 4'b1000 : node15796;
															assign node15796 = (inp[14]) ? 4'b1001 : 4'b1000;
										assign node15801 = (inp[1]) ? node15833 : node15802;
											assign node15802 = (inp[13]) ? node15820 : node15803;
												assign node15803 = (inp[7]) ? node15815 : node15804;
													assign node15804 = (inp[14]) ? node15810 : node15805;
														assign node15805 = (inp[10]) ? node15807 : 4'b1001;
															assign node15807 = (inp[12]) ? 4'b1001 : 4'b0001;
														assign node15810 = (inp[11]) ? node15812 : 4'b1000;
															assign node15812 = (inp[10]) ? 4'b0001 : 4'b1001;
													assign node15815 = (inp[10]) ? node15817 : 4'b1010;
														assign node15817 = (inp[11]) ? 4'b1010 : 4'b0001;
												assign node15820 = (inp[12]) ? node15828 : node15821;
													assign node15821 = (inp[10]) ? node15823 : 4'b0001;
														assign node15823 = (inp[14]) ? node15825 : 4'b1001;
															assign node15825 = (inp[11]) ? 4'b1001 : 4'b1000;
													assign node15828 = (inp[11]) ? 4'b0001 : node15829;
														assign node15829 = (inp[14]) ? 4'b0000 : 4'b0001;
											assign node15833 = (inp[11]) ? node15867 : node15834;
												assign node15834 = (inp[14]) ? node15852 : node15835;
													assign node15835 = (inp[10]) ? node15849 : node15836;
														assign node15836 = (inp[7]) ? node15844 : node15837;
															assign node15837 = (inp[12]) ? node15841 : node15838;
																assign node15838 = (inp[13]) ? 4'b1000 : 4'b0000;
																assign node15841 = (inp[13]) ? 4'b0000 : 4'b1000;
															assign node15844 = (inp[13]) ? node15846 : 4'b1010;
																assign node15846 = (inp[12]) ? 4'b0000 : 4'b1000;
														assign node15849 = (inp[13]) ? 4'b1000 : 4'b0000;
													assign node15852 = (inp[13]) ? node15862 : node15853;
														assign node15853 = (inp[7]) ? node15857 : node15854;
															assign node15854 = (inp[10]) ? 4'b0001 : 4'b1001;
															assign node15857 = (inp[12]) ? 4'b1010 : node15858;
																assign node15858 = (inp[10]) ? 4'b0001 : 4'b1010;
														assign node15862 = (inp[10]) ? node15864 : 4'b0001;
															assign node15864 = (inp[12]) ? 4'b0001 : 4'b1001;
												assign node15867 = (inp[13]) ? node15875 : node15868;
													assign node15868 = (inp[12]) ? node15870 : 4'b0000;
														assign node15870 = (inp[10]) ? 4'b0000 : node15871;
															assign node15871 = (inp[7]) ? 4'b1010 : 4'b1000;
													assign node15875 = (inp[12]) ? node15877 : 4'b1000;
														assign node15877 = (inp[10]) ? 4'b1000 : 4'b0000;
							assign node15881 = (inp[2]) ? node16233 : node15882;
								assign node15882 = (inp[1]) ? node16064 : node15883;
									assign node15883 = (inp[14]) ? node15951 : node15884;
										assign node15884 = (inp[13]) ? node15920 : node15885;
											assign node15885 = (inp[12]) ? node15909 : node15886;
												assign node15886 = (inp[10]) ? node15898 : node15887;
													assign node15887 = (inp[3]) ? node15893 : node15888;
														assign node15888 = (inp[4]) ? node15890 : 4'b1001;
															assign node15890 = (inp[11]) ? 4'b1101 : 4'b1001;
														assign node15893 = (inp[4]) ? node15895 : 4'b1101;
															assign node15895 = (inp[7]) ? 4'b1101 : 4'b1001;
													assign node15898 = (inp[3]) ? node15904 : node15899;
														assign node15899 = (inp[7]) ? node15901 : 4'b0101;
															assign node15901 = (inp[4]) ? 4'b0101 : 4'b0001;
														assign node15904 = (inp[4]) ? 4'b0001 : node15905;
															assign node15905 = (inp[7]) ? 4'b0101 : 4'b0001;
												assign node15909 = (inp[3]) ? node15915 : node15910;
													assign node15910 = (inp[4]) ? node15912 : 4'b1001;
														assign node15912 = (inp[7]) ? 4'b1001 : 4'b1101;
													assign node15915 = (inp[7]) ? 4'b1101 : node15916;
														assign node15916 = (inp[4]) ? 4'b1001 : 4'b1101;
											assign node15920 = (inp[12]) ? node15940 : node15921;
												assign node15921 = (inp[10]) ? node15929 : node15922;
													assign node15922 = (inp[3]) ? 4'b0001 : node15923;
														assign node15923 = (inp[4]) ? 4'b0101 : node15924;
															assign node15924 = (inp[7]) ? 4'b0001 : 4'b0101;
													assign node15929 = (inp[3]) ? node15935 : node15930;
														assign node15930 = (inp[7]) ? node15932 : 4'b1101;
															assign node15932 = (inp[4]) ? 4'b1101 : 4'b1001;
														assign node15935 = (inp[4]) ? 4'b1001 : node15936;
															assign node15936 = (inp[7]) ? 4'b1101 : 4'b1001;
												assign node15940 = (inp[3]) ? node15946 : node15941;
													assign node15941 = (inp[7]) ? node15943 : 4'b0101;
														assign node15943 = (inp[4]) ? 4'b0101 : 4'b0001;
													assign node15946 = (inp[7]) ? node15948 : 4'b0001;
														assign node15948 = (inp[4]) ? 4'b0001 : 4'b0101;
										assign node15951 = (inp[11]) ? node16007 : node15952;
											assign node15952 = (inp[13]) ? node15978 : node15953;
												assign node15953 = (inp[12]) ? node15971 : node15954;
													assign node15954 = (inp[10]) ? node15964 : node15955;
														assign node15955 = (inp[7]) ? 4'b1000 : node15956;
															assign node15956 = (inp[4]) ? node15960 : node15957;
																assign node15957 = (inp[3]) ? 4'b1100 : 4'b1000;
																assign node15960 = (inp[3]) ? 4'b1000 : 4'b1100;
														assign node15964 = (inp[3]) ? 4'b0000 : node15965;
															assign node15965 = (inp[7]) ? node15967 : 4'b0100;
																assign node15967 = (inp[4]) ? 4'b0100 : 4'b0000;
													assign node15971 = (inp[3]) ? node15973 : 4'b1000;
														assign node15973 = (inp[7]) ? 4'b1100 : node15974;
															assign node15974 = (inp[4]) ? 4'b1000 : 4'b1100;
												assign node15978 = (inp[10]) ? node15990 : node15979;
													assign node15979 = (inp[3]) ? node15985 : node15980;
														assign node15980 = (inp[4]) ? 4'b0100 : node15981;
															assign node15981 = (inp[7]) ? 4'b0000 : 4'b0100;
														assign node15985 = (inp[7]) ? node15987 : 4'b0000;
															assign node15987 = (inp[4]) ? 4'b0000 : 4'b0100;
													assign node15990 = (inp[12]) ? node16000 : node15991;
														assign node15991 = (inp[3]) ? node15997 : node15992;
															assign node15992 = (inp[7]) ? node15994 : 4'b1100;
																assign node15994 = (inp[4]) ? 4'b1100 : 4'b1000;
															assign node15997 = (inp[4]) ? 4'b1000 : 4'b1100;
														assign node16000 = (inp[4]) ? node16004 : node16001;
															assign node16001 = (inp[3]) ? 4'b0100 : 4'b0000;
															assign node16004 = (inp[3]) ? 4'b0000 : 4'b0100;
											assign node16007 = (inp[13]) ? node16035 : node16008;
												assign node16008 = (inp[12]) ? node16024 : node16009;
													assign node16009 = (inp[10]) ? node16015 : node16010;
														assign node16010 = (inp[3]) ? node16012 : 4'b1001;
															assign node16012 = (inp[4]) ? 4'b1001 : 4'b1101;
														assign node16015 = (inp[3]) ? node16019 : node16016;
															assign node16016 = (inp[7]) ? 4'b0001 : 4'b0101;
															assign node16019 = (inp[4]) ? 4'b0001 : node16020;
																assign node16020 = (inp[7]) ? 4'b0101 : 4'b0001;
													assign node16024 = (inp[4]) ? node16028 : node16025;
														assign node16025 = (inp[3]) ? 4'b1101 : 4'b1001;
														assign node16028 = (inp[3]) ? node16032 : node16029;
															assign node16029 = (inp[7]) ? 4'b1001 : 4'b1101;
															assign node16032 = (inp[7]) ? 4'b1101 : 4'b1001;
												assign node16035 = (inp[10]) ? node16047 : node16036;
													assign node16036 = (inp[3]) ? node16042 : node16037;
														assign node16037 = (inp[4]) ? 4'b0101 : node16038;
															assign node16038 = (inp[7]) ? 4'b0001 : 4'b0101;
														assign node16042 = (inp[4]) ? 4'b0001 : node16043;
															assign node16043 = (inp[7]) ? 4'b0101 : 4'b0001;
													assign node16047 = (inp[12]) ? node16059 : node16048;
														assign node16048 = (inp[3]) ? node16054 : node16049;
															assign node16049 = (inp[7]) ? node16051 : 4'b1101;
																assign node16051 = (inp[4]) ? 4'b1101 : 4'b1001;
															assign node16054 = (inp[7]) ? node16056 : 4'b1001;
																assign node16056 = (inp[4]) ? 4'b1001 : 4'b1101;
														assign node16059 = (inp[3]) ? node16061 : 4'b0101;
															assign node16061 = (inp[7]) ? 4'b0101 : 4'b0001;
									assign node16064 = (inp[14]) ? node16126 : node16065;
										assign node16065 = (inp[13]) ? node16097 : node16066;
											assign node16066 = (inp[10]) ? node16086 : node16067;
												assign node16067 = (inp[12]) ? node16075 : node16068;
													assign node16068 = (inp[3]) ? 4'b0000 : node16069;
														assign node16069 = (inp[7]) ? node16071 : 4'b0100;
															assign node16071 = (inp[11]) ? 4'b0000 : 4'b0100;
													assign node16075 = (inp[3]) ? node16081 : node16076;
														assign node16076 = (inp[7]) ? 4'b1000 : node16077;
															assign node16077 = (inp[11]) ? 4'b1100 : 4'b1000;
														assign node16081 = (inp[4]) ? node16083 : 4'b1100;
															assign node16083 = (inp[7]) ? 4'b1100 : 4'b1000;
												assign node16086 = (inp[3]) ? node16092 : node16087;
													assign node16087 = (inp[7]) ? node16089 : 4'b0100;
														assign node16089 = (inp[4]) ? 4'b0100 : 4'b0000;
													assign node16092 = (inp[7]) ? node16094 : 4'b0000;
														assign node16094 = (inp[4]) ? 4'b0000 : 4'b0100;
											assign node16097 = (inp[12]) ? node16109 : node16098;
												assign node16098 = (inp[3]) ? node16104 : node16099;
													assign node16099 = (inp[7]) ? node16101 : 4'b1100;
														assign node16101 = (inp[4]) ? 4'b1100 : 4'b1000;
													assign node16104 = (inp[4]) ? 4'b1000 : node16105;
														assign node16105 = (inp[7]) ? 4'b1100 : 4'b1000;
												assign node16109 = (inp[10]) ? node16121 : node16110;
													assign node16110 = (inp[3]) ? node16116 : node16111;
														assign node16111 = (inp[7]) ? node16113 : 4'b0100;
															assign node16113 = (inp[4]) ? 4'b0100 : 4'b0000;
														assign node16116 = (inp[4]) ? 4'b0000 : node16117;
															assign node16117 = (inp[7]) ? 4'b0100 : 4'b0000;
													assign node16121 = (inp[3]) ? node16123 : 4'b1100;
														assign node16123 = (inp[4]) ? 4'b1000 : 4'b1100;
										assign node16126 = (inp[11]) ? node16182 : node16127;
											assign node16127 = (inp[13]) ? node16159 : node16128;
												assign node16128 = (inp[10]) ? node16140 : node16129;
													assign node16129 = (inp[3]) ? node16135 : node16130;
														assign node16130 = (inp[7]) ? 4'b1001 : node16131;
															assign node16131 = (inp[12]) ? 4'b1001 : 4'b1101;
														assign node16135 = (inp[4]) ? node16137 : 4'b1101;
															assign node16137 = (inp[7]) ? 4'b1101 : 4'b1001;
													assign node16140 = (inp[12]) ? node16152 : node16141;
														assign node16141 = (inp[3]) ? node16147 : node16142;
															assign node16142 = (inp[4]) ? 4'b0101 : node16143;
																assign node16143 = (inp[7]) ? 4'b0001 : 4'b0101;
															assign node16147 = (inp[7]) ? node16149 : 4'b0001;
																assign node16149 = (inp[4]) ? 4'b0001 : 4'b0101;
														assign node16152 = (inp[3]) ? node16154 : 4'b1001;
															assign node16154 = (inp[7]) ? 4'b1101 : node16155;
																assign node16155 = (inp[4]) ? 4'b1001 : 4'b1101;
												assign node16159 = (inp[10]) ? node16171 : node16160;
													assign node16160 = (inp[3]) ? node16166 : node16161;
														assign node16161 = (inp[7]) ? node16163 : 4'b0101;
															assign node16163 = (inp[12]) ? 4'b0001 : 4'b0101;
														assign node16166 = (inp[4]) ? 4'b0001 : node16167;
															assign node16167 = (inp[7]) ? 4'b0101 : 4'b0001;
													assign node16171 = (inp[12]) ? node16177 : node16172;
														assign node16172 = (inp[3]) ? node16174 : 4'b1101;
															assign node16174 = (inp[4]) ? 4'b1001 : 4'b1101;
														assign node16177 = (inp[4]) ? node16179 : 4'b0001;
															assign node16179 = (inp[3]) ? 4'b0001 : 4'b0101;
											assign node16182 = (inp[13]) ? node16210 : node16183;
												assign node16183 = (inp[12]) ? node16195 : node16184;
													assign node16184 = (inp[3]) ? node16190 : node16185;
														assign node16185 = (inp[4]) ? 4'b0100 : node16186;
															assign node16186 = (inp[7]) ? 4'b0000 : 4'b0100;
														assign node16190 = (inp[4]) ? 4'b0000 : node16191;
															assign node16191 = (inp[10]) ? 4'b0000 : 4'b0100;
													assign node16195 = (inp[10]) ? node16205 : node16196;
														assign node16196 = (inp[4]) ? node16198 : 4'b1100;
															assign node16198 = (inp[7]) ? node16202 : node16199;
																assign node16199 = (inp[3]) ? 4'b1000 : 4'b1100;
																assign node16202 = (inp[3]) ? 4'b1100 : 4'b1000;
														assign node16205 = (inp[7]) ? 4'b0100 : node16206;
															assign node16206 = (inp[3]) ? 4'b0000 : 4'b0100;
												assign node16210 = (inp[3]) ? node16222 : node16211;
													assign node16211 = (inp[10]) ? node16217 : node16212;
														assign node16212 = (inp[12]) ? 4'b0100 : node16213;
															assign node16213 = (inp[7]) ? 4'b1000 : 4'b1100;
														assign node16217 = (inp[4]) ? 4'b1100 : node16218;
															assign node16218 = (inp[7]) ? 4'b1000 : 4'b1100;
													assign node16222 = (inp[10]) ? node16228 : node16223;
														assign node16223 = (inp[12]) ? node16225 : 4'b1000;
															assign node16225 = (inp[4]) ? 4'b0000 : 4'b0100;
														assign node16228 = (inp[4]) ? 4'b1000 : node16229;
															assign node16229 = (inp[7]) ? 4'b1100 : 4'b1000;
								assign node16233 = (inp[3]) ? node16235 : 4'b1010;
									assign node16235 = (inp[7]) ? node16305 : node16236;
										assign node16236 = (inp[1]) ? node16270 : node16237;
											assign node16237 = (inp[13]) ? node16257 : node16238;
												assign node16238 = (inp[4]) ? node16248 : node16239;
													assign node16239 = (inp[10]) ? node16241 : 4'b1010;
														assign node16241 = (inp[12]) ? 4'b1010 : node16242;
															assign node16242 = (inp[14]) ? node16244 : 4'b0001;
																assign node16244 = (inp[11]) ? 4'b0001 : 4'b0000;
													assign node16248 = (inp[12]) ? node16252 : node16249;
														assign node16249 = (inp[10]) ? 4'b0001 : 4'b1000;
														assign node16252 = (inp[14]) ? node16254 : 4'b1001;
															assign node16254 = (inp[11]) ? 4'b1001 : 4'b1000;
												assign node16257 = (inp[11]) ? node16265 : node16258;
													assign node16258 = (inp[14]) ? node16260 : 4'b0001;
														assign node16260 = (inp[10]) ? node16262 : 4'b0000;
															assign node16262 = (inp[12]) ? 4'b0000 : 4'b1000;
													assign node16265 = (inp[12]) ? 4'b0001 : node16266;
														assign node16266 = (inp[10]) ? 4'b1001 : 4'b0001;
											assign node16270 = (inp[11]) ? node16292 : node16271;
												assign node16271 = (inp[14]) ? node16283 : node16272;
													assign node16272 = (inp[13]) ? node16278 : node16273;
														assign node16273 = (inp[10]) ? 4'b0000 : node16274;
															assign node16274 = (inp[12]) ? 4'b1000 : 4'b0000;
														assign node16278 = (inp[12]) ? node16280 : 4'b1000;
															assign node16280 = (inp[10]) ? 4'b1000 : 4'b0000;
													assign node16283 = (inp[13]) ? node16287 : node16284;
														assign node16284 = (inp[4]) ? 4'b1001 : 4'b1010;
														assign node16287 = (inp[10]) ? node16289 : 4'b0001;
															assign node16289 = (inp[12]) ? 4'b0001 : 4'b1001;
												assign node16292 = (inp[13]) ? node16300 : node16293;
													assign node16293 = (inp[10]) ? 4'b0000 : node16294;
														assign node16294 = (inp[12]) ? node16296 : 4'b0000;
															assign node16296 = (inp[4]) ? 4'b1000 : 4'b1010;
													assign node16300 = (inp[12]) ? node16302 : 4'b1000;
														assign node16302 = (inp[10]) ? 4'b1000 : 4'b0000;
										assign node16305 = (inp[4]) ? node16307 : 4'b1010;
											assign node16307 = (inp[13]) ? node16327 : node16308;
												assign node16308 = (inp[12]) ? node16318 : node16309;
													assign node16309 = (inp[10]) ? node16315 : node16310;
														assign node16310 = (inp[1]) ? node16312 : 4'b1010;
															assign node16312 = (inp[11]) ? 4'b0000 : 4'b1010;
														assign node16315 = (inp[1]) ? 4'b0000 : 4'b0001;
													assign node16318 = (inp[1]) ? node16320 : 4'b1010;
														assign node16320 = (inp[10]) ? node16322 : 4'b1010;
															assign node16322 = (inp[14]) ? node16324 : 4'b0000;
																assign node16324 = (inp[11]) ? 4'b0000 : 4'b1010;
												assign node16327 = (inp[12]) ? node16339 : node16328;
													assign node16328 = (inp[11]) ? 4'b1000 : node16329;
														assign node16329 = (inp[10]) ? node16335 : node16330;
															assign node16330 = (inp[14]) ? node16332 : 4'b1000;
																assign node16332 = (inp[1]) ? 4'b0001 : 4'b0000;
															assign node16335 = (inp[1]) ? 4'b1001 : 4'b1000;
													assign node16339 = (inp[1]) ? node16345 : node16340;
														assign node16340 = (inp[11]) ? 4'b0001 : node16341;
															assign node16341 = (inp[14]) ? 4'b0000 : 4'b0001;
														assign node16345 = (inp[10]) ? 4'b1000 : node16346;
															assign node16346 = (inp[11]) ? 4'b0000 : node16347;
																assign node16347 = (inp[14]) ? 4'b0001 : 4'b0000;
						assign node16352 = (inp[5]) ? node17132 : node16353;
							assign node16353 = (inp[1]) ? node16763 : node16354;
								assign node16354 = (inp[13]) ? node16524 : node16355;
									assign node16355 = (inp[10]) ? node16409 : node16356;
										assign node16356 = (inp[3]) ? node16378 : node16357;
											assign node16357 = (inp[14]) ? node16363 : node16358;
												assign node16358 = (inp[7]) ? 4'b1001 : node16359;
													assign node16359 = (inp[4]) ? 4'b1101 : 4'b1001;
												assign node16363 = (inp[11]) ? node16369 : node16364;
													assign node16364 = (inp[4]) ? node16366 : 4'b1000;
														assign node16366 = (inp[7]) ? 4'b1000 : 4'b1100;
													assign node16369 = (inp[7]) ? 4'b1001 : node16370;
														assign node16370 = (inp[4]) ? node16372 : 4'b1001;
															assign node16372 = (inp[2]) ? 4'b1101 : node16373;
																assign node16373 = (inp[12]) ? 4'b1101 : 4'b0000;
											assign node16378 = (inp[11]) ? node16390 : node16379;
												assign node16379 = (inp[4]) ? node16385 : node16380;
													assign node16380 = (inp[2]) ? node16382 : 4'b1001;
														assign node16382 = (inp[14]) ? 4'b1100 : 4'b1101;
													assign node16385 = (inp[2]) ? node16387 : 4'b1101;
														assign node16387 = (inp[7]) ? 4'b1101 : 4'b1000;
												assign node16390 = (inp[2]) ? node16402 : node16391;
													assign node16391 = (inp[12]) ? node16399 : node16392;
														assign node16392 = (inp[7]) ? node16396 : node16393;
															assign node16393 = (inp[4]) ? 4'b0000 : 4'b0100;
															assign node16396 = (inp[4]) ? 4'b0100 : 4'b0000;
														assign node16399 = (inp[4]) ? 4'b1100 : 4'b1000;
													assign node16402 = (inp[4]) ? node16404 : 4'b1101;
														assign node16404 = (inp[7]) ? 4'b1101 : node16405;
															assign node16405 = (inp[12]) ? 4'b1001 : 4'b0000;
										assign node16409 = (inp[12]) ? node16471 : node16410;
											assign node16410 = (inp[11]) ? node16448 : node16411;
												assign node16411 = (inp[14]) ? node16429 : node16412;
													assign node16412 = (inp[3]) ? node16422 : node16413;
														assign node16413 = (inp[4]) ? node16417 : node16414;
															assign node16414 = (inp[7]) ? 4'b0001 : 4'b0101;
															assign node16417 = (inp[7]) ? 4'b0101 : node16418;
																assign node16418 = (inp[2]) ? 4'b0101 : 4'b0001;
														assign node16422 = (inp[2]) ? 4'b0001 : node16423;
															assign node16423 = (inp[4]) ? 4'b0001 : node16424;
																assign node16424 = (inp[7]) ? 4'b0001 : 4'b0101;
													assign node16429 = (inp[2]) ? node16437 : node16430;
														assign node16430 = (inp[7]) ? node16432 : 4'b0001;
															assign node16432 = (inp[4]) ? 4'b0100 : node16433;
																assign node16433 = (inp[3]) ? 4'b0001 : 4'b0000;
														assign node16437 = (inp[3]) ? node16443 : node16438;
															assign node16438 = (inp[7]) ? node16440 : 4'b0100;
																assign node16440 = (inp[4]) ? 4'b0100 : 4'b0000;
															assign node16443 = (inp[4]) ? node16445 : 4'b0100;
																assign node16445 = (inp[7]) ? 4'b0000 : 4'b0001;
												assign node16448 = (inp[2]) ? node16464 : node16449;
													assign node16449 = (inp[3]) ? node16457 : node16450;
														assign node16450 = (inp[7]) ? node16454 : node16451;
															assign node16451 = (inp[4]) ? 4'b1000 : 4'b0101;
															assign node16454 = (inp[4]) ? 4'b0101 : 4'b0001;
														assign node16457 = (inp[7]) ? node16461 : node16458;
															assign node16458 = (inp[4]) ? 4'b1000 : 4'b1100;
															assign node16461 = (inp[4]) ? 4'b1100 : 4'b1000;
													assign node16464 = (inp[3]) ? node16466 : 4'b0101;
														assign node16466 = (inp[7]) ? node16468 : 4'b1000;
															assign node16468 = (inp[4]) ? 4'b0001 : 4'b0101;
											assign node16471 = (inp[3]) ? node16495 : node16472;
												assign node16472 = (inp[14]) ? node16484 : node16473;
													assign node16473 = (inp[4]) ? node16475 : 4'b1001;
														assign node16475 = (inp[2]) ? node16481 : node16476;
															assign node16476 = (inp[7]) ? 4'b1001 : node16477;
																assign node16477 = (inp[11]) ? 4'b0000 : 4'b0001;
															assign node16481 = (inp[7]) ? 4'b1001 : 4'b1101;
													assign node16484 = (inp[11]) ? node16492 : node16485;
														assign node16485 = (inp[4]) ? node16487 : 4'b1000;
															assign node16487 = (inp[2]) ? node16489 : 4'b0001;
																assign node16489 = (inp[7]) ? 4'b1000 : 4'b1100;
														assign node16492 = (inp[7]) ? 4'b1001 : 4'b1101;
												assign node16495 = (inp[2]) ? node16513 : node16496;
													assign node16496 = (inp[11]) ? node16506 : node16497;
														assign node16497 = (inp[14]) ? 4'b0101 : node16498;
															assign node16498 = (inp[7]) ? node16502 : node16499;
																assign node16499 = (inp[4]) ? 4'b0001 : 4'b0101;
																assign node16502 = (inp[4]) ? 4'b0101 : 4'b0001;
														assign node16506 = (inp[7]) ? node16510 : node16507;
															assign node16507 = (inp[4]) ? 4'b0000 : 4'b0100;
															assign node16510 = (inp[4]) ? 4'b0100 : 4'b0000;
													assign node16513 = (inp[4]) ? node16519 : node16514;
														assign node16514 = (inp[14]) ? node16516 : 4'b1101;
															assign node16516 = (inp[11]) ? 4'b1101 : 4'b1100;
														assign node16519 = (inp[7]) ? 4'b1101 : node16520;
															assign node16520 = (inp[11]) ? 4'b0000 : 4'b0001;
									assign node16524 = (inp[12]) ? node16646 : node16525;
										assign node16525 = (inp[10]) ? node16595 : node16526;
											assign node16526 = (inp[3]) ? node16566 : node16527;
												assign node16527 = (inp[2]) ? node16553 : node16528;
													assign node16528 = (inp[14]) ? node16538 : node16529;
														assign node16529 = (inp[7]) ? node16535 : node16530;
															assign node16530 = (inp[11]) ? node16532 : 4'b1001;
																assign node16532 = (inp[4]) ? 4'b0000 : 4'b0101;
															assign node16535 = (inp[4]) ? 4'b0101 : 4'b0001;
														assign node16538 = (inp[7]) ? node16546 : node16539;
															assign node16539 = (inp[4]) ? node16543 : node16540;
																assign node16540 = (inp[11]) ? 4'b0101 : 4'b0100;
																assign node16543 = (inp[11]) ? 4'b0000 : 4'b1001;
															assign node16546 = (inp[4]) ? node16550 : node16547;
																assign node16547 = (inp[11]) ? 4'b0001 : 4'b0000;
																assign node16550 = (inp[11]) ? 4'b0000 : 4'b0100;
													assign node16553 = (inp[7]) ? node16559 : node16554;
														assign node16554 = (inp[14]) ? node16556 : 4'b0101;
															assign node16556 = (inp[11]) ? 4'b0101 : 4'b0100;
														assign node16559 = (inp[4]) ? 4'b0101 : node16560;
															assign node16560 = (inp[14]) ? node16562 : 4'b0001;
																assign node16562 = (inp[11]) ? 4'b0001 : 4'b0000;
												assign node16566 = (inp[11]) ? node16584 : node16567;
													assign node16567 = (inp[2]) ? node16577 : node16568;
														assign node16568 = (inp[7]) ? node16574 : node16569;
															assign node16569 = (inp[4]) ? node16571 : 4'b1101;
																assign node16571 = (inp[14]) ? 4'b0001 : 4'b1000;
															assign node16574 = (inp[4]) ? 4'b1101 : 4'b1001;
														assign node16577 = (inp[7]) ? 4'b0000 : node16578;
															assign node16578 = (inp[4]) ? 4'b1001 : node16579;
																assign node16579 = (inp[14]) ? 4'b0000 : 4'b0001;
													assign node16584 = (inp[4]) ? node16590 : node16585;
														assign node16585 = (inp[2]) ? node16587 : 4'b0100;
															assign node16587 = (inp[7]) ? 4'b0101 : 4'b0001;
														assign node16590 = (inp[2]) ? 4'b0000 : node16591;
															assign node16591 = (inp[7]) ? 4'b0000 : 4'b1001;
											assign node16595 = (inp[4]) ? node16627 : node16596;
												assign node16596 = (inp[14]) ? node16608 : node16597;
													assign node16597 = (inp[3]) ? node16601 : node16598;
														assign node16598 = (inp[7]) ? 4'b1001 : 4'b1101;
														assign node16601 = (inp[2]) ? node16605 : node16602;
															assign node16602 = (inp[11]) ? 4'b1100 : 4'b0101;
															assign node16605 = (inp[7]) ? 4'b1101 : 4'b1001;
													assign node16608 = (inp[11]) ? node16618 : node16609;
														assign node16609 = (inp[3]) ? node16613 : node16610;
															assign node16610 = (inp[7]) ? 4'b1000 : 4'b1100;
															assign node16613 = (inp[2]) ? node16615 : 4'b0101;
																assign node16615 = (inp[7]) ? 4'b1100 : 4'b1000;
														assign node16618 = (inp[2]) ? node16622 : node16619;
															assign node16619 = (inp[3]) ? 4'b1100 : 4'b1101;
															assign node16622 = (inp[3]) ? node16624 : 4'b1101;
																assign node16624 = (inp[7]) ? 4'b1101 : 4'b1001;
												assign node16627 = (inp[2]) ? node16637 : node16628;
													assign node16628 = (inp[3]) ? node16632 : node16629;
														assign node16629 = (inp[11]) ? 4'b1000 : 4'b0001;
														assign node16632 = (inp[14]) ? 4'b0001 : node16633;
															assign node16633 = (inp[11]) ? 4'b0001 : 4'b0000;
													assign node16637 = (inp[3]) ? node16643 : node16638;
														assign node16638 = (inp[14]) ? node16640 : 4'b1101;
															assign node16640 = (inp[11]) ? 4'b1101 : 4'b1100;
														assign node16643 = (inp[11]) ? 4'b1000 : 4'b0001;
										assign node16646 = (inp[10]) ? node16708 : node16647;
											assign node16647 = (inp[3]) ? node16675 : node16648;
												assign node16648 = (inp[14]) ? node16658 : node16649;
													assign node16649 = (inp[7]) ? node16655 : node16650;
														assign node16650 = (inp[4]) ? node16652 : 4'b0101;
															assign node16652 = (inp[2]) ? 4'b0101 : 4'b1001;
														assign node16655 = (inp[4]) ? 4'b0101 : 4'b0001;
													assign node16658 = (inp[11]) ? node16668 : node16659;
														assign node16659 = (inp[2]) ? 4'b0100 : node16660;
															assign node16660 = (inp[4]) ? node16664 : node16661;
																assign node16661 = (inp[7]) ? 4'b0000 : 4'b0100;
																assign node16664 = (inp[7]) ? 4'b0100 : 4'b1001;
														assign node16668 = (inp[7]) ? node16672 : node16669;
															assign node16669 = (inp[4]) ? 4'b1000 : 4'b0101;
															assign node16672 = (inp[4]) ? 4'b0101 : 4'b0001;
												assign node16675 = (inp[2]) ? node16691 : node16676;
													assign node16676 = (inp[11]) ? node16684 : node16677;
														assign node16677 = (inp[4]) ? node16681 : node16678;
															assign node16678 = (inp[7]) ? 4'b1001 : 4'b1101;
															assign node16681 = (inp[7]) ? 4'b1101 : 4'b0001;
														assign node16684 = (inp[4]) ? node16688 : node16685;
															assign node16685 = (inp[7]) ? 4'b1000 : 4'b1100;
															assign node16688 = (inp[7]) ? 4'b1100 : 4'b0001;
													assign node16691 = (inp[4]) ? node16699 : node16692;
														assign node16692 = (inp[7]) ? 4'b0101 : node16693;
															assign node16693 = (inp[11]) ? 4'b0001 : node16694;
																assign node16694 = (inp[14]) ? 4'b0000 : 4'b0001;
														assign node16699 = (inp[7]) ? node16703 : node16700;
															assign node16700 = (inp[11]) ? 4'b1000 : 4'b1001;
															assign node16703 = (inp[14]) ? node16705 : 4'b0001;
																assign node16705 = (inp[11]) ? 4'b0001 : 4'b0000;
											assign node16708 = (inp[4]) ? node16730 : node16709;
												assign node16709 = (inp[3]) ? node16721 : node16710;
													assign node16710 = (inp[7]) ? node16716 : node16711;
														assign node16711 = (inp[11]) ? 4'b0101 : node16712;
															assign node16712 = (inp[14]) ? 4'b0100 : 4'b0101;
														assign node16716 = (inp[14]) ? node16718 : 4'b0001;
															assign node16718 = (inp[11]) ? 4'b0001 : 4'b0000;
													assign node16721 = (inp[11]) ? node16725 : node16722;
														assign node16722 = (inp[2]) ? 4'b0100 : 4'b0101;
														assign node16725 = (inp[2]) ? node16727 : 4'b0100;
															assign node16727 = (inp[7]) ? 4'b0101 : 4'b0001;
												assign node16730 = (inp[3]) ? node16740 : node16731;
													assign node16731 = (inp[2]) ? node16735 : node16732;
														assign node16732 = (inp[11]) ? 4'b0000 : 4'b0001;
														assign node16735 = (inp[11]) ? 4'b0101 : node16736;
															assign node16736 = (inp[14]) ? 4'b0100 : 4'b0101;
													assign node16740 = (inp[14]) ? node16754 : node16741;
														assign node16741 = (inp[7]) ? node16747 : node16742;
															assign node16742 = (inp[11]) ? 4'b0001 : node16743;
																assign node16743 = (inp[2]) ? 4'b0001 : 4'b0000;
															assign node16747 = (inp[11]) ? node16751 : node16748;
																assign node16748 = (inp[2]) ? 4'b0001 : 4'b0000;
																assign node16751 = (inp[2]) ? 4'b0000 : 4'b0001;
														assign node16754 = (inp[11]) ? node16760 : node16755;
															assign node16755 = (inp[7]) ? 4'b0001 : node16756;
																assign node16756 = (inp[2]) ? 4'b0001 : 4'b1001;
															assign node16760 = (inp[2]) ? 4'b0000 : 4'b0001;
								assign node16763 = (inp[11]) ? node16993 : node16764;
									assign node16764 = (inp[14]) ? node16884 : node16765;
										assign node16765 = (inp[3]) ? node16821 : node16766;
											assign node16766 = (inp[7]) ? node16796 : node16767;
												assign node16767 = (inp[2]) ? node16785 : node16768;
													assign node16768 = (inp[4]) ? node16776 : node16769;
														assign node16769 = (inp[10]) ? 4'b1100 : node16770;
															assign node16770 = (inp[12]) ? node16772 : 4'b0100;
																assign node16772 = (inp[13]) ? 4'b0100 : 4'b1000;
														assign node16776 = (inp[12]) ? node16780 : node16777;
															assign node16777 = (inp[10]) ? 4'b1001 : 4'b0001;
															assign node16780 = (inp[10]) ? 4'b0001 : node16781;
																assign node16781 = (inp[13]) ? 4'b1001 : 4'b1100;
													assign node16785 = (inp[13]) ? node16791 : node16786;
														assign node16786 = (inp[12]) ? node16788 : 4'b0100;
															assign node16788 = (inp[4]) ? 4'b1100 : 4'b0100;
														assign node16791 = (inp[10]) ? 4'b1100 : node16792;
															assign node16792 = (inp[12]) ? 4'b0100 : 4'b1100;
												assign node16796 = (inp[4]) ? node16808 : node16797;
													assign node16797 = (inp[13]) ? node16803 : node16798;
														assign node16798 = (inp[12]) ? node16800 : 4'b0000;
															assign node16800 = (inp[10]) ? 4'b0000 : 4'b1000;
														assign node16803 = (inp[10]) ? 4'b1000 : node16804;
															assign node16804 = (inp[12]) ? 4'b0000 : 4'b1000;
													assign node16808 = (inp[2]) ? node16814 : node16809;
														assign node16809 = (inp[13]) ? node16811 : 4'b0100;
															assign node16811 = (inp[12]) ? 4'b0100 : 4'b0001;
														assign node16814 = (inp[12]) ? node16818 : node16815;
															assign node16815 = (inp[13]) ? 4'b1100 : 4'b0100;
															assign node16818 = (inp[13]) ? 4'b0100 : 4'b1000;
											assign node16821 = (inp[2]) ? node16851 : node16822;
												assign node16822 = (inp[4]) ? node16838 : node16823;
													assign node16823 = (inp[13]) ? node16833 : node16824;
														assign node16824 = (inp[7]) ? 4'b1001 : node16825;
															assign node16825 = (inp[10]) ? node16829 : node16826;
																assign node16826 = (inp[12]) ? 4'b1001 : 4'b0101;
																assign node16829 = (inp[12]) ? 4'b0101 : 4'b1101;
														assign node16833 = (inp[10]) ? node16835 : 4'b0101;
															assign node16835 = (inp[12]) ? 4'b0101 : 4'b1101;
													assign node16838 = (inp[7]) ? node16846 : node16839;
														assign node16839 = (inp[13]) ? node16841 : 4'b0001;
															assign node16841 = (inp[10]) ? node16843 : 4'b1001;
																assign node16843 = (inp[12]) ? 4'b0001 : 4'b1001;
														assign node16846 = (inp[13]) ? 4'b0001 : node16847;
															assign node16847 = (inp[10]) ? 4'b1101 : 4'b0101;
												assign node16851 = (inp[4]) ? node16867 : node16852;
													assign node16852 = (inp[7]) ? node16860 : node16853;
														assign node16853 = (inp[13]) ? 4'b1000 : node16854;
															assign node16854 = (inp[10]) ? 4'b0000 : node16855;
																assign node16855 = (inp[12]) ? 4'b1100 : 4'b0000;
														assign node16860 = (inp[13]) ? 4'b1100 : node16861;
															assign node16861 = (inp[12]) ? node16863 : 4'b0100;
																assign node16863 = (inp[10]) ? 4'b0100 : 4'b1100;
													assign node16867 = (inp[10]) ? node16877 : node16868;
														assign node16868 = (inp[12]) ? node16874 : node16869;
															assign node16869 = (inp[13]) ? 4'b0001 : node16870;
																assign node16870 = (inp[7]) ? 4'b0000 : 4'b0001;
															assign node16874 = (inp[13]) ? 4'b0000 : 4'b1000;
														assign node16877 = (inp[12]) ? node16879 : 4'b1001;
															assign node16879 = (inp[13]) ? 4'b0001 : node16880;
																assign node16880 = (inp[7]) ? 4'b0000 : 4'b0001;
										assign node16884 = (inp[13]) ? node16932 : node16885;
											assign node16885 = (inp[3]) ? node16907 : node16886;
												assign node16886 = (inp[10]) ? node16892 : node16887;
													assign node16887 = (inp[7]) ? 4'b1001 : node16888;
														assign node16888 = (inp[4]) ? 4'b1101 : 4'b1001;
													assign node16892 = (inp[12]) ? node16902 : node16893;
														assign node16893 = (inp[2]) ? node16899 : node16894;
															assign node16894 = (inp[4]) ? node16896 : 4'b0101;
																assign node16896 = (inp[7]) ? 4'b0101 : 4'b1001;
															assign node16899 = (inp[7]) ? 4'b0001 : 4'b0101;
														assign node16902 = (inp[7]) ? 4'b1001 : node16903;
															assign node16903 = (inp[4]) ? 4'b0001 : 4'b1001;
												assign node16907 = (inp[2]) ? node16923 : node16908;
													assign node16908 = (inp[12]) ? node16916 : node16909;
														assign node16909 = (inp[4]) ? node16911 : 4'b1101;
															assign node16911 = (inp[10]) ? 4'b0000 : node16912;
																assign node16912 = (inp[7]) ? 4'b0101 : 4'b0001;
														assign node16916 = (inp[10]) ? node16918 : 4'b1101;
															assign node16918 = (inp[7]) ? node16920 : 4'b0101;
																assign node16920 = (inp[4]) ? 4'b0101 : 4'b0001;
													assign node16923 = (inp[4]) ? node16925 : 4'b1101;
														assign node16925 = (inp[7]) ? 4'b1101 : node16926;
															assign node16926 = (inp[12]) ? 4'b1001 : node16927;
																assign node16927 = (inp[10]) ? 4'b1001 : 4'b0001;
											assign node16932 = (inp[4]) ? node16960 : node16933;
												assign node16933 = (inp[10]) ? node16945 : node16934;
													assign node16934 = (inp[3]) ? node16938 : node16935;
														assign node16935 = (inp[7]) ? 4'b0001 : 4'b0101;
														assign node16938 = (inp[12]) ? node16940 : 4'b0101;
															assign node16940 = (inp[2]) ? node16942 : 4'b1101;
																assign node16942 = (inp[7]) ? 4'b0101 : 4'b0001;
													assign node16945 = (inp[12]) ? node16953 : node16946;
														assign node16946 = (inp[7]) ? 4'b1101 : node16947;
															assign node16947 = (inp[2]) ? node16949 : 4'b1101;
																assign node16949 = (inp[3]) ? 4'b1001 : 4'b1101;
														assign node16953 = (inp[2]) ? node16955 : 4'b0101;
															assign node16955 = (inp[3]) ? node16957 : 4'b0101;
																assign node16957 = (inp[7]) ? 4'b0101 : 4'b0001;
												assign node16960 = (inp[3]) ? node16974 : node16961;
													assign node16961 = (inp[2]) ? node16969 : node16962;
														assign node16962 = (inp[10]) ? node16966 : node16963;
															assign node16963 = (inp[12]) ? 4'b0101 : 4'b0001;
															assign node16966 = (inp[12]) ? 4'b0001 : 4'b1001;
														assign node16969 = (inp[10]) ? node16971 : 4'b0101;
															assign node16971 = (inp[12]) ? 4'b0101 : 4'b1101;
													assign node16974 = (inp[2]) ? node16984 : node16975;
														assign node16975 = (inp[10]) ? node16981 : node16976;
															assign node16976 = (inp[7]) ? node16978 : 4'b1000;
																assign node16978 = (inp[12]) ? 4'b1101 : 4'b0001;
															assign node16981 = (inp[12]) ? 4'b0000 : 4'b1000;
														assign node16984 = (inp[7]) ? node16990 : node16985;
															assign node16985 = (inp[12]) ? node16987 : 4'b1001;
																assign node16987 = (inp[10]) ? 4'b0001 : 4'b1001;
															assign node16990 = (inp[10]) ? 4'b1001 : 4'b0001;
									assign node16993 = (inp[10]) ? node17091 : node16994;
										assign node16994 = (inp[2]) ? node17030 : node16995;
											assign node16995 = (inp[4]) ? node17017 : node16996;
												assign node16996 = (inp[7]) ? node17006 : node16997;
													assign node16997 = (inp[3]) ? 4'b0100 : node16998;
														assign node16998 = (inp[13]) ? node17002 : node16999;
															assign node16999 = (inp[12]) ? 4'b1000 : 4'b0100;
															assign node17002 = (inp[12]) ? 4'b0100 : 4'b1100;
													assign node17006 = (inp[3]) ? node17014 : node17007;
														assign node17007 = (inp[13]) ? node17011 : node17008;
															assign node17008 = (inp[12]) ? 4'b1000 : 4'b0000;
															assign node17011 = (inp[12]) ? 4'b0000 : 4'b1000;
														assign node17014 = (inp[13]) ? 4'b0100 : 4'b0000;
												assign node17017 = (inp[7]) ? node17023 : node17018;
													assign node17018 = (inp[14]) ? node17020 : 4'b0000;
														assign node17020 = (inp[13]) ? 4'b1000 : 4'b0000;
													assign node17023 = (inp[13]) ? 4'b0000 : node17024;
														assign node17024 = (inp[12]) ? node17026 : 4'b0100;
															assign node17026 = (inp[3]) ? 4'b0100 : 4'b1000;
											assign node17030 = (inp[3]) ? node17068 : node17031;
												assign node17031 = (inp[7]) ? node17045 : node17032;
													assign node17032 = (inp[4]) ? node17040 : node17033;
														assign node17033 = (inp[13]) ? node17037 : node17034;
															assign node17034 = (inp[12]) ? 4'b1000 : 4'b0100;
															assign node17037 = (inp[12]) ? 4'b0100 : 4'b1100;
														assign node17040 = (inp[12]) ? node17042 : 4'b0100;
															assign node17042 = (inp[13]) ? 4'b0100 : 4'b1100;
													assign node17045 = (inp[4]) ? node17061 : node17046;
														assign node17046 = (inp[14]) ? node17054 : node17047;
															assign node17047 = (inp[12]) ? node17051 : node17048;
																assign node17048 = (inp[13]) ? 4'b1000 : 4'b0000;
																assign node17051 = (inp[13]) ? 4'b0000 : 4'b1000;
															assign node17054 = (inp[13]) ? node17058 : node17055;
																assign node17055 = (inp[12]) ? 4'b1000 : 4'b0000;
																assign node17058 = (inp[12]) ? 4'b0000 : 4'b1000;
														assign node17061 = (inp[12]) ? node17065 : node17062;
															assign node17062 = (inp[13]) ? 4'b1100 : 4'b0100;
															assign node17065 = (inp[13]) ? 4'b0100 : 4'b1000;
												assign node17068 = (inp[4]) ? node17084 : node17069;
													assign node17069 = (inp[7]) ? node17077 : node17070;
														assign node17070 = (inp[13]) ? node17074 : node17071;
															assign node17071 = (inp[12]) ? 4'b1100 : 4'b0000;
															assign node17074 = (inp[12]) ? 4'b0000 : 4'b1000;
														assign node17077 = (inp[13]) ? node17081 : node17078;
															assign node17078 = (inp[12]) ? 4'b1100 : 4'b0100;
															assign node17081 = (inp[12]) ? 4'b0100 : 4'b1100;
													assign node17084 = (inp[12]) ? node17086 : 4'b0000;
														assign node17086 = (inp[13]) ? 4'b0000 : node17087;
															assign node17087 = (inp[14]) ? 4'b0000 : 4'b1100;
										assign node17091 = (inp[13]) ? node17117 : node17092;
											assign node17092 = (inp[3]) ? node17102 : node17093;
												assign node17093 = (inp[7]) ? node17099 : node17094;
													assign node17094 = (inp[4]) ? node17096 : 4'b0100;
														assign node17096 = (inp[2]) ? 4'b0100 : 4'b1000;
													assign node17099 = (inp[4]) ? 4'b0100 : 4'b0000;
												assign node17102 = (inp[2]) ? node17110 : node17103;
													assign node17103 = (inp[4]) ? node17107 : node17104;
														assign node17104 = (inp[7]) ? 4'b1000 : 4'b1100;
														assign node17107 = (inp[7]) ? 4'b1100 : 4'b0000;
													assign node17110 = (inp[4]) ? node17114 : node17111;
														assign node17111 = (inp[7]) ? 4'b0100 : 4'b0000;
														assign node17114 = (inp[7]) ? 4'b0000 : 4'b1000;
											assign node17117 = (inp[4]) ? node17127 : node17118;
												assign node17118 = (inp[7]) ? node17124 : node17119;
													assign node17119 = (inp[2]) ? node17121 : 4'b1100;
														assign node17121 = (inp[14]) ? 4'b1100 : 4'b1000;
													assign node17124 = (inp[3]) ? 4'b1100 : 4'b1000;
												assign node17127 = (inp[3]) ? 4'b1000 : node17128;
													assign node17128 = (inp[2]) ? 4'b1100 : 4'b1000;
							assign node17132 = (inp[3]) ? node17510 : node17133;
								assign node17133 = (inp[4]) ? node17325 : node17134;
									assign node17134 = (inp[11]) ? node17252 : node17135;
										assign node17135 = (inp[2]) ? node17205 : node17136;
											assign node17136 = (inp[13]) ? node17170 : node17137;
												assign node17137 = (inp[7]) ? node17155 : node17138;
													assign node17138 = (inp[1]) ? node17148 : node17139;
														assign node17139 = (inp[14]) ? node17143 : node17140;
															assign node17140 = (inp[10]) ? 4'b1100 : 4'b0100;
															assign node17143 = (inp[10]) ? node17145 : 4'b1001;
																assign node17145 = (inp[12]) ? 4'b0101 : 4'b1101;
														assign node17148 = (inp[14]) ? node17150 : 4'b0101;
															assign node17150 = (inp[12]) ? node17152 : 4'b0100;
																assign node17152 = (inp[10]) ? 4'b1100 : 4'b0100;
													assign node17155 = (inp[12]) ? node17165 : node17156;
														assign node17156 = (inp[1]) ? node17160 : node17157;
															assign node17157 = (inp[14]) ? 4'b1001 : 4'b0000;
															assign node17160 = (inp[14]) ? node17162 : 4'b0001;
																assign node17162 = (inp[10]) ? 4'b0100 : 4'b0000;
														assign node17165 = (inp[1]) ? node17167 : 4'b1000;
															assign node17167 = (inp[14]) ? 4'b1000 : 4'b1001;
												assign node17170 = (inp[10]) ? node17190 : node17171;
													assign node17171 = (inp[7]) ? node17181 : node17172;
														assign node17172 = (inp[12]) ? node17176 : node17173;
															assign node17173 = (inp[1]) ? 4'b1000 : 4'b0000;
															assign node17176 = (inp[1]) ? 4'b0000 : node17177;
																assign node17177 = (inp[14]) ? 4'b0101 : 4'b0100;
														assign node17181 = (inp[1]) ? node17187 : node17182;
															assign node17182 = (inp[12]) ? node17184 : 4'b1100;
																assign node17184 = (inp[14]) ? 4'b0101 : 4'b0100;
															assign node17187 = (inp[14]) ? 4'b1100 : 4'b1101;
													assign node17190 = (inp[14]) ? node17198 : node17191;
														assign node17191 = (inp[12]) ? node17195 : node17192;
															assign node17192 = (inp[1]) ? 4'b1000 : 4'b0000;
															assign node17195 = (inp[1]) ? 4'b0000 : 4'b1000;
														assign node17198 = (inp[12]) ? node17202 : node17199;
															assign node17199 = (inp[1]) ? 4'b1000 : 4'b0000;
															assign node17202 = (inp[7]) ? 4'b1101 : 4'b1000;
											assign node17205 = (inp[10]) ? node17219 : node17206;
												assign node17206 = (inp[12]) ? node17214 : node17207;
													assign node17207 = (inp[1]) ? node17209 : 4'b1001;
														assign node17209 = (inp[7]) ? node17211 : 4'b0101;
															assign node17211 = (inp[13]) ? 4'b0101 : 4'b0001;
													assign node17214 = (inp[13]) ? node17216 : 4'b1001;
														assign node17216 = (inp[7]) ? 4'b1001 : 4'b1101;
												assign node17219 = (inp[12]) ? node17239 : node17220;
													assign node17220 = (inp[1]) ? node17230 : node17221;
														assign node17221 = (inp[14]) ? 4'b0001 : node17222;
															assign node17222 = (inp[7]) ? node17226 : node17223;
																assign node17223 = (inp[13]) ? 4'b0000 : 4'b0101;
																assign node17226 = (inp[13]) ? 4'b0101 : 4'b0001;
														assign node17230 = (inp[14]) ? node17232 : 4'b1001;
															assign node17232 = (inp[7]) ? node17236 : node17233;
																assign node17233 = (inp[13]) ? 4'b1000 : 4'b1101;
																assign node17236 = (inp[13]) ? 4'b1101 : 4'b1001;
													assign node17239 = (inp[7]) ? node17249 : node17240;
														assign node17240 = (inp[13]) ? node17242 : 4'b0101;
															assign node17242 = (inp[14]) ? node17246 : node17243;
																assign node17243 = (inp[1]) ? 4'b0001 : 4'b0000;
																assign node17246 = (inp[1]) ? 4'b0000 : 4'b0101;
														assign node17249 = (inp[13]) ? 4'b0101 : 4'b0001;
										assign node17252 = (inp[1]) ? node17290 : node17253;
											assign node17253 = (inp[2]) ? node17271 : node17254;
												assign node17254 = (inp[13]) ? node17264 : node17255;
													assign node17255 = (inp[12]) ? node17261 : node17256;
														assign node17256 = (inp[7]) ? 4'b0001 : node17257;
															assign node17257 = (inp[10]) ? 4'b1101 : 4'b0101;
														assign node17261 = (inp[10]) ? 4'b1101 : 4'b1001;
													assign node17264 = (inp[7]) ? node17266 : 4'b0000;
														assign node17266 = (inp[10]) ? 4'b0000 : node17267;
															assign node17267 = (inp[12]) ? 4'b0101 : 4'b1101;
												assign node17271 = (inp[10]) ? node17283 : node17272;
													assign node17272 = (inp[12]) ? node17278 : node17273;
														assign node17273 = (inp[7]) ? node17275 : 4'b0100;
															assign node17275 = (inp[13]) ? 4'b0100 : 4'b0000;
														assign node17278 = (inp[7]) ? 4'b1000 : node17279;
															assign node17279 = (inp[13]) ? 4'b1100 : 4'b1000;
													assign node17283 = (inp[7]) ? node17287 : node17284;
														assign node17284 = (inp[13]) ? 4'b0001 : 4'b0100;
														assign node17287 = (inp[13]) ? 4'b0100 : 4'b0000;
											assign node17290 = (inp[10]) ? node17314 : node17291;
												assign node17291 = (inp[2]) ? node17305 : node17292;
													assign node17292 = (inp[13]) ? node17300 : node17293;
														assign node17293 = (inp[7]) ? node17297 : node17294;
															assign node17294 = (inp[12]) ? 4'b0100 : 4'b1100;
															assign node17297 = (inp[12]) ? 4'b0000 : 4'b1000;
														assign node17300 = (inp[7]) ? node17302 : 4'b1000;
															assign node17302 = (inp[12]) ? 4'b1100 : 4'b0100;
													assign node17305 = (inp[7]) ? node17311 : node17306;
														assign node17306 = (inp[14]) ? node17308 : 4'b0100;
															assign node17308 = (inp[12]) ? 4'b0100 : 4'b0000;
														assign node17311 = (inp[13]) ? 4'b0100 : 4'b0000;
												assign node17314 = (inp[13]) ? node17320 : node17315;
													assign node17315 = (inp[2]) ? node17317 : 4'b0100;
														assign node17317 = (inp[7]) ? 4'b1000 : 4'b1100;
													assign node17320 = (inp[7]) ? node17322 : 4'b1000;
														assign node17322 = (inp[2]) ? 4'b1100 : 4'b1000;
									assign node17325 = (inp[1]) ? node17427 : node17326;
										assign node17326 = (inp[11]) ? node17394 : node17327;
											assign node17327 = (inp[10]) ? node17359 : node17328;
												assign node17328 = (inp[14]) ? node17346 : node17329;
													assign node17329 = (inp[2]) ? node17337 : node17330;
														assign node17330 = (inp[13]) ? node17334 : node17331;
															assign node17331 = (inp[12]) ? 4'b1000 : 4'b0100;
															assign node17334 = (inp[12]) ? 4'b0001 : 4'b1001;
														assign node17337 = (inp[12]) ? node17343 : node17338;
															assign node17338 = (inp[13]) ? node17340 : 4'b0000;
																assign node17340 = (inp[7]) ? 4'b1000 : 4'b0000;
															assign node17343 = (inp[7]) ? 4'b0000 : 4'b0100;
													assign node17346 = (inp[2]) ? node17356 : node17347;
														assign node17347 = (inp[13]) ? node17353 : node17348;
															assign node17348 = (inp[12]) ? 4'b1000 : node17349;
																assign node17349 = (inp[7]) ? 4'b0000 : 4'b0100;
															assign node17353 = (inp[12]) ? 4'b0000 : 4'b1000;
														assign node17356 = (inp[12]) ? 4'b1101 : 4'b1001;
												assign node17359 = (inp[12]) ? node17373 : node17360;
													assign node17360 = (inp[2]) ? node17368 : node17361;
														assign node17361 = (inp[13]) ? node17365 : node17362;
															assign node17362 = (inp[7]) ? 4'b0100 : 4'b0000;
															assign node17365 = (inp[7]) ? 4'b1000 : 4'b1001;
														assign node17368 = (inp[13]) ? 4'b0000 : node17369;
															assign node17369 = (inp[14]) ? 4'b1001 : 4'b1000;
													assign node17373 = (inp[13]) ? node17381 : node17374;
														assign node17374 = (inp[14]) ? node17376 : 4'b1000;
															assign node17376 = (inp[2]) ? 4'b0001 : node17377;
																assign node17377 = (inp[7]) ? 4'b1000 : 4'b0000;
														assign node17381 = (inp[14]) ? node17389 : node17382;
															assign node17382 = (inp[2]) ? node17386 : node17383;
																assign node17383 = (inp[7]) ? 4'b1001 : 4'b0001;
																assign node17386 = (inp[7]) ? 4'b0100 : 4'b1000;
															assign node17389 = (inp[7]) ? node17391 : 4'b1000;
																assign node17391 = (inp[2]) ? 4'b1001 : 4'b1000;
											assign node17394 = (inp[13]) ? node17412 : node17395;
												assign node17395 = (inp[2]) ? node17405 : node17396;
													assign node17396 = (inp[10]) ? node17400 : node17397;
														assign node17397 = (inp[7]) ? 4'b0000 : 4'b0100;
														assign node17400 = (inp[7]) ? 4'b0100 : node17401;
															assign node17401 = (inp[12]) ? 4'b0001 : 4'b1001;
													assign node17405 = (inp[10]) ? 4'b1001 : node17406;
														assign node17406 = (inp[12]) ? node17408 : 4'b0001;
															assign node17408 = (inp[7]) ? 4'b1100 : 4'b1001;
												assign node17412 = (inp[2]) ? node17420 : node17413;
													assign node17413 = (inp[10]) ? node17415 : 4'b1001;
														assign node17415 = (inp[12]) ? node17417 : 4'b0000;
															assign node17417 = (inp[7]) ? 4'b1001 : 4'b1000;
													assign node17420 = (inp[10]) ? 4'b0000 : node17421;
														assign node17421 = (inp[7]) ? node17423 : 4'b0000;
															assign node17423 = (inp[12]) ? 4'b0001 : 4'b1001;
										assign node17427 = (inp[11]) ? node17483 : node17428;
											assign node17428 = (inp[13]) ? node17458 : node17429;
												assign node17429 = (inp[2]) ? node17445 : node17430;
													assign node17430 = (inp[12]) ? node17436 : node17431;
														assign node17431 = (inp[10]) ? 4'b0000 : node17432;
															assign node17432 = (inp[7]) ? 4'b1000 : 4'b1100;
														assign node17436 = (inp[7]) ? node17442 : node17437;
															assign node17437 = (inp[10]) ? node17439 : 4'b0100;
																assign node17439 = (inp[14]) ? 4'b1001 : 4'b1000;
															assign node17442 = (inp[10]) ? 4'b0100 : 4'b0000;
													assign node17445 = (inp[14]) ? node17451 : node17446;
														assign node17446 = (inp[7]) ? node17448 : 4'b0101;
															assign node17448 = (inp[10]) ? 4'b1001 : 4'b0001;
														assign node17451 = (inp[10]) ? node17453 : 4'b0000;
															assign node17453 = (inp[12]) ? 4'b1000 : node17454;
																assign node17454 = (inp[7]) ? 4'b0000 : 4'b0100;
												assign node17458 = (inp[2]) ? node17468 : node17459;
													assign node17459 = (inp[10]) ? 4'b0001 : node17460;
														assign node17460 = (inp[14]) ? node17464 : node17461;
															assign node17461 = (inp[7]) ? 4'b0000 : 4'b0100;
															assign node17464 = (inp[12]) ? 4'b1001 : 4'b0101;
													assign node17468 = (inp[12]) ? node17476 : node17469;
														assign node17469 = (inp[14]) ? 4'b1000 : node17470;
															assign node17470 = (inp[10]) ? 4'b1000 : node17471;
																assign node17471 = (inp[7]) ? 4'b1001 : 4'b1000;
														assign node17476 = (inp[10]) ? 4'b0000 : node17477;
															assign node17477 = (inp[14]) ? node17479 : 4'b1001;
																assign node17479 = (inp[7]) ? 4'b1000 : 4'b0000;
											assign node17483 = (inp[13]) ? node17501 : node17484;
												assign node17484 = (inp[10]) ? node17496 : node17485;
													assign node17485 = (inp[12]) ? node17491 : node17486;
														assign node17486 = (inp[2]) ? 4'b1000 : node17487;
															assign node17487 = (inp[7]) ? 4'b1000 : 4'b0000;
														assign node17491 = (inp[2]) ? 4'b0000 : node17492;
															assign node17492 = (inp[7]) ? 4'b1000 : 4'b1100;
													assign node17496 = (inp[7]) ? 4'b0000 : node17497;
														assign node17497 = (inp[2]) ? 4'b0100 : 4'b0000;
												assign node17501 = (inp[10]) ? 4'b1000 : node17502;
													assign node17502 = (inp[2]) ? 4'b1000 : node17503;
														assign node17503 = (inp[7]) ? node17505 : 4'b0000;
															assign node17505 = (inp[12]) ? 4'b0000 : 4'b1000;
								assign node17510 = (inp[1]) ? node17754 : node17511;
									assign node17511 = (inp[4]) ? node17637 : node17512;
										assign node17512 = (inp[7]) ? node17572 : node17513;
											assign node17513 = (inp[10]) ? node17545 : node17514;
												assign node17514 = (inp[11]) ? node17534 : node17515;
													assign node17515 = (inp[12]) ? node17525 : node17516;
														assign node17516 = (inp[14]) ? node17520 : node17517;
															assign node17517 = (inp[2]) ? 4'b0001 : 4'b0000;
															assign node17520 = (inp[13]) ? 4'b1000 : node17521;
																assign node17521 = (inp[2]) ? 4'b0000 : 4'b0001;
														assign node17525 = (inp[14]) ? node17529 : node17526;
															assign node17526 = (inp[2]) ? 4'b1001 : 4'b0000;
															assign node17529 = (inp[13]) ? 4'b1000 : node17530;
																assign node17530 = (inp[2]) ? 4'b1000 : 4'b1001;
													assign node17534 = (inp[13]) ? node17540 : node17535;
														assign node17535 = (inp[2]) ? 4'b0001 : node17536;
															assign node17536 = (inp[14]) ? 4'b0001 : 4'b1001;
														assign node17540 = (inp[12]) ? node17542 : 4'b0000;
															assign node17542 = (inp[2]) ? 4'b0000 : 4'b0001;
												assign node17545 = (inp[12]) ? node17561 : node17546;
													assign node17546 = (inp[2]) ? node17556 : node17547;
														assign node17547 = (inp[14]) ? node17553 : node17548;
															assign node17548 = (inp[11]) ? 4'b1000 : node17549;
																assign node17549 = (inp[13]) ? 4'b1000 : 4'b0000;
															assign node17553 = (inp[13]) ? 4'b1001 : 4'b1000;
														assign node17556 = (inp[11]) ? node17558 : 4'b0000;
															assign node17558 = (inp[13]) ? 4'b1000 : 4'b0000;
													assign node17561 = (inp[13]) ? node17565 : node17562;
														assign node17562 = (inp[11]) ? 4'b0001 : 4'b0000;
														assign node17565 = (inp[2]) ? node17569 : node17566;
															assign node17566 = (inp[11]) ? 4'b0000 : 4'b0001;
															assign node17569 = (inp[11]) ? 4'b1000 : 4'b0000;
											assign node17572 = (inp[10]) ? node17608 : node17573;
												assign node17573 = (inp[11]) ? node17597 : node17574;
													assign node17574 = (inp[12]) ? node17590 : node17575;
														assign node17575 = (inp[14]) ? node17583 : node17576;
															assign node17576 = (inp[2]) ? node17580 : node17577;
																assign node17577 = (inp[13]) ? 4'b0000 : 4'b0001;
																assign node17580 = (inp[13]) ? 4'b0001 : 4'b0000;
															assign node17583 = (inp[2]) ? node17587 : node17584;
																assign node17584 = (inp[13]) ? 4'b0000 : 4'b0001;
																assign node17587 = (inp[13]) ? 4'b0001 : 4'b0000;
														assign node17590 = (inp[13]) ? node17594 : node17591;
															assign node17591 = (inp[2]) ? 4'b1000 : 4'b1001;
															assign node17594 = (inp[14]) ? 4'b0000 : 4'b0001;
													assign node17597 = (inp[12]) ? node17603 : node17598;
														assign node17598 = (inp[2]) ? 4'b1000 : node17599;
															assign node17599 = (inp[13]) ? 4'b0001 : 4'b1000;
														assign node17603 = (inp[13]) ? node17605 : 4'b0000;
															assign node17605 = (inp[2]) ? 4'b0000 : 4'b0001;
												assign node17608 = (inp[13]) ? node17620 : node17609;
													assign node17609 = (inp[11]) ? node17615 : node17610;
														assign node17610 = (inp[2]) ? node17612 : 4'b0000;
															assign node17612 = (inp[14]) ? 4'b0000 : 4'b0001;
														assign node17615 = (inp[2]) ? node17617 : 4'b0001;
															assign node17617 = (inp[12]) ? 4'b0001 : 4'b1001;
													assign node17620 = (inp[12]) ? node17628 : node17621;
														assign node17621 = (inp[2]) ? node17625 : node17622;
															assign node17622 = (inp[11]) ? 4'b0001 : 4'b1001;
															assign node17625 = (inp[11]) ? 4'b1001 : 4'b1000;
														assign node17628 = (inp[2]) ? node17632 : node17629;
															assign node17629 = (inp[11]) ? 4'b0001 : 4'b1001;
															assign node17632 = (inp[11]) ? 4'b1001 : node17633;
																assign node17633 = (inp[14]) ? 4'b0001 : 4'b0000;
										assign node17637 = (inp[13]) ? node17701 : node17638;
											assign node17638 = (inp[10]) ? node17668 : node17639;
												assign node17639 = (inp[7]) ? node17653 : node17640;
													assign node17640 = (inp[11]) ? node17646 : node17641;
														assign node17641 = (inp[12]) ? 4'b0001 : node17642;
															assign node17642 = (inp[2]) ? 4'b0001 : 4'b1001;
														assign node17646 = (inp[12]) ? node17650 : node17647;
															assign node17647 = (inp[2]) ? 4'b0001 : 4'b1001;
															assign node17650 = (inp[2]) ? 4'b1000 : 4'b0001;
													assign node17653 = (inp[2]) ? node17661 : node17654;
														assign node17654 = (inp[12]) ? 4'b0000 : node17655;
															assign node17655 = (inp[11]) ? 4'b1000 : node17656;
																assign node17656 = (inp[14]) ? 4'b1000 : 4'b1001;
														assign node17661 = (inp[12]) ? node17665 : node17662;
															assign node17662 = (inp[14]) ? 4'b0000 : 4'b0001;
															assign node17665 = (inp[11]) ? 4'b1001 : 4'b0001;
												assign node17668 = (inp[12]) ? node17680 : node17669;
													assign node17669 = (inp[2]) ? node17675 : node17670;
														assign node17670 = (inp[7]) ? node17672 : 4'b0000;
															assign node17672 = (inp[11]) ? 4'b0000 : 4'b0001;
														assign node17675 = (inp[7]) ? node17677 : 4'b0001;
															assign node17677 = (inp[11]) ? 4'b0000 : 4'b1000;
													assign node17680 = (inp[7]) ? node17686 : node17681;
														assign node17681 = (inp[11]) ? 4'b0001 : node17682;
															assign node17682 = (inp[2]) ? 4'b1000 : 4'b0001;
														assign node17686 = (inp[14]) ? node17694 : node17687;
															assign node17687 = (inp[2]) ? node17691 : node17688;
																assign node17688 = (inp[11]) ? 4'b0000 : 4'b0001;
																assign node17691 = (inp[11]) ? 4'b0001 : 4'b0000;
															assign node17694 = (inp[2]) ? node17698 : node17695;
																assign node17695 = (inp[11]) ? 4'b0000 : 4'b0001;
																assign node17698 = (inp[11]) ? 4'b0001 : 4'b0000;
											assign node17701 = (inp[10]) ? node17735 : node17702;
												assign node17702 = (inp[2]) ? node17720 : node17703;
													assign node17703 = (inp[14]) ? node17713 : node17704;
														assign node17704 = (inp[7]) ? node17706 : 4'b0000;
															assign node17706 = (inp[11]) ? node17710 : node17707;
																assign node17707 = (inp[12]) ? 4'b0000 : 4'b0001;
																assign node17710 = (inp[12]) ? 4'b0001 : 4'b0000;
														assign node17713 = (inp[7]) ? node17717 : node17714;
															assign node17714 = (inp[11]) ? 4'b0000 : 4'b0001;
															assign node17717 = (inp[11]) ? 4'b0001 : 4'b0000;
													assign node17720 = (inp[7]) ? node17726 : node17721;
														assign node17721 = (inp[12]) ? 4'b0001 : node17722;
															assign node17722 = (inp[11]) ? 4'b0000 : 4'b0001;
														assign node17726 = (inp[11]) ? node17732 : node17727;
															assign node17727 = (inp[14]) ? node17729 : 4'b0000;
																assign node17729 = (inp[12]) ? 4'b0001 : 4'b0000;
															assign node17732 = (inp[12]) ? 4'b0000 : 4'b0001;
												assign node17735 = (inp[11]) ? 4'b0000 : node17736;
													assign node17736 = (inp[12]) ? node17744 : node17737;
														assign node17737 = (inp[7]) ? node17739 : 4'b0000;
															assign node17739 = (inp[14]) ? node17741 : 4'b0000;
																assign node17741 = (inp[2]) ? 4'b0001 : 4'b0000;
														assign node17744 = (inp[14]) ? node17748 : node17745;
															assign node17745 = (inp[2]) ? 4'b0001 : 4'b0000;
															assign node17748 = (inp[2]) ? node17750 : 4'b0001;
																assign node17750 = (inp[7]) ? 4'b0000 : 4'b0001;
									assign node17754 = (inp[4]) ? node17852 : node17755;
										assign node17755 = (inp[11]) ? node17815 : node17756;
											assign node17756 = (inp[10]) ? node17796 : node17757;
												assign node17757 = (inp[2]) ? node17775 : node17758;
													assign node17758 = (inp[12]) ? node17766 : node17759;
														assign node17759 = (inp[7]) ? 4'b0000 : node17760;
															assign node17760 = (inp[13]) ? 4'b1001 : node17761;
																assign node17761 = (inp[14]) ? 4'b0000 : 4'b0001;
														assign node17766 = (inp[13]) ? node17772 : node17767;
															assign node17767 = (inp[7]) ? 4'b1001 : node17768;
																assign node17768 = (inp[14]) ? 4'b1000 : 4'b1001;
															assign node17772 = (inp[7]) ? 4'b1000 : 4'b0001;
													assign node17775 = (inp[12]) ? node17787 : node17776;
														assign node17776 = (inp[13]) ? node17782 : node17777;
															assign node17777 = (inp[14]) ? node17779 : 4'b1000;
																assign node17779 = (inp[7]) ? 4'b1000 : 4'b1001;
															assign node17782 = (inp[7]) ? 4'b1001 : node17783;
																assign node17783 = (inp[14]) ? 4'b1000 : 4'b1001;
														assign node17787 = (inp[14]) ? node17791 : node17788;
															assign node17788 = (inp[7]) ? 4'b0000 : 4'b1000;
															assign node17791 = (inp[7]) ? 4'b1001 : node17792;
																assign node17792 = (inp[13]) ? 4'b0000 : 4'b0001;
												assign node17796 = (inp[2]) ? node17806 : node17797;
													assign node17797 = (inp[12]) ? node17799 : 4'b0000;
														assign node17799 = (inp[13]) ? node17801 : 4'b0000;
															assign node17801 = (inp[7]) ? node17803 : 4'b1000;
																assign node17803 = (inp[14]) ? 4'b1000 : 4'b1001;
													assign node17806 = (inp[13]) ? node17810 : node17807;
														assign node17807 = (inp[7]) ? 4'b1001 : 4'b0001;
														assign node17810 = (inp[12]) ? 4'b0000 : node17811;
															assign node17811 = (inp[14]) ? 4'b0001 : 4'b0000;
											assign node17815 = (inp[10]) ? node17843 : node17816;
												assign node17816 = (inp[13]) ? node17836 : node17817;
													assign node17817 = (inp[7]) ? node17825 : node17818;
														assign node17818 = (inp[12]) ? node17822 : node17819;
															assign node17819 = (inp[2]) ? 4'b0000 : 4'b1000;
															assign node17822 = (inp[2]) ? 4'b1000 : 4'b0000;
														assign node17825 = (inp[14]) ? node17831 : node17826;
															assign node17826 = (inp[2]) ? 4'b1000 : node17827;
																assign node17827 = (inp[12]) ? 4'b0000 : 4'b1000;
															assign node17831 = (inp[12]) ? 4'b1000 : node17832;
																assign node17832 = (inp[2]) ? 4'b0000 : 4'b1000;
													assign node17836 = (inp[2]) ? node17838 : 4'b0000;
														assign node17838 = (inp[7]) ? 4'b0000 : node17839;
															assign node17839 = (inp[14]) ? 4'b0000 : 4'b1000;
												assign node17843 = (inp[13]) ? 4'b1000 : node17844;
													assign node17844 = (inp[7]) ? node17848 : node17845;
														assign node17845 = (inp[2]) ? 4'b1000 : 4'b0000;
														assign node17848 = (inp[2]) ? 4'b0000 : 4'b1000;
										assign node17852 = (inp[11]) ? node17896 : node17853;
											assign node17853 = (inp[13]) ? node17881 : node17854;
												assign node17854 = (inp[7]) ? node17868 : node17855;
													assign node17855 = (inp[14]) ? node17857 : 4'b0000;
														assign node17857 = (inp[12]) ? node17863 : node17858;
															assign node17858 = (inp[2]) ? 4'b0000 : node17859;
																assign node17859 = (inp[10]) ? 4'b0000 : 4'b1000;
															assign node17863 = (inp[2]) ? 4'b1000 : node17864;
																assign node17864 = (inp[10]) ? 4'b0000 : 4'b1000;
													assign node17868 = (inp[12]) ? node17874 : node17869;
														assign node17869 = (inp[10]) ? 4'b0001 : node17870;
															assign node17870 = (inp[2]) ? 4'b1001 : 4'b1000;
														assign node17874 = (inp[14]) ? node17876 : 4'b0001;
															assign node17876 = (inp[10]) ? 4'b0001 : node17877;
																assign node17877 = (inp[2]) ? 4'b0001 : 4'b0000;
												assign node17881 = (inp[10]) ? 4'b0000 : node17882;
													assign node17882 = (inp[12]) ? node17888 : node17883;
														assign node17883 = (inp[14]) ? 4'b0000 : node17884;
															assign node17884 = (inp[2]) ? 4'b0001 : 4'b0000;
														assign node17888 = (inp[7]) ? node17890 : 4'b0001;
															assign node17890 = (inp[2]) ? node17892 : 4'b0000;
																assign node17892 = (inp[14]) ? 4'b0000 : 4'b0001;
											assign node17896 = (inp[10]) ? 4'b0000 : node17897;
												assign node17897 = (inp[13]) ? 4'b0000 : node17898;
													assign node17898 = (inp[12]) ? node17904 : node17899;
														assign node17899 = (inp[7]) ? node17901 : 4'b0000;
															assign node17901 = (inp[2]) ? 4'b1000 : 4'b0000;
														assign node17904 = (inp[14]) ? node17908 : node17905;
															assign node17905 = (inp[2]) ? 4'b1000 : 4'b0000;
															assign node17908 = (inp[7]) ? node17910 : 4'b1000;
																assign node17910 = (inp[2]) ? 4'b0000 : 4'b1000;
					assign node17915 = (inp[6]) ? node17917 : 4'b1000;
						assign node17917 = (inp[5]) ? node18035 : node17918;
							assign node17918 = (inp[2]) ? 4'b1000 : node17919;
								assign node17919 = (inp[3]) ? node17921 : 4'b1000;
									assign node17921 = (inp[7]) ? node17987 : node17922;
										assign node17922 = (inp[1]) ? node17954 : node17923;
											assign node17923 = (inp[13]) ? node17941 : node17924;
												assign node17924 = (inp[4]) ? node17930 : node17925;
													assign node17925 = (inp[11]) ? node17927 : 4'b1000;
														assign node17927 = (inp[12]) ? 4'b1000 : 4'b0001;
													assign node17930 = (inp[14]) ? node17936 : node17931;
														assign node17931 = (inp[12]) ? 4'b1001 : node17932;
															assign node17932 = (inp[10]) ? 4'b0001 : 4'b1001;
														assign node17936 = (inp[11]) ? 4'b1001 : node17937;
															assign node17937 = (inp[10]) ? 4'b0000 : 4'b1000;
												assign node17941 = (inp[10]) ? node17947 : node17942;
													assign node17942 = (inp[14]) ? node17944 : 4'b0001;
														assign node17944 = (inp[11]) ? 4'b0001 : 4'b0000;
													assign node17947 = (inp[12]) ? 4'b0001 : node17948;
														assign node17948 = (inp[14]) ? node17950 : 4'b1001;
															assign node17950 = (inp[11]) ? 4'b1001 : 4'b1000;
											assign node17954 = (inp[11]) ? node17976 : node17955;
												assign node17955 = (inp[14]) ? node17963 : node17956;
													assign node17956 = (inp[13]) ? 4'b1000 : node17957;
														assign node17957 = (inp[10]) ? 4'b0000 : node17958;
															assign node17958 = (inp[12]) ? 4'b1000 : 4'b0000;
													assign node17963 = (inp[13]) ? node17971 : node17964;
														assign node17964 = (inp[10]) ? node17968 : node17965;
															assign node17965 = (inp[4]) ? 4'b1001 : 4'b1000;
															assign node17968 = (inp[12]) ? 4'b1001 : 4'b0001;
														assign node17971 = (inp[12]) ? 4'b0001 : node17972;
															assign node17972 = (inp[10]) ? 4'b1001 : 4'b0001;
												assign node17976 = (inp[13]) ? node17982 : node17977;
													assign node17977 = (inp[12]) ? node17979 : 4'b0000;
														assign node17979 = (inp[10]) ? 4'b0000 : 4'b1000;
													assign node17982 = (inp[12]) ? node17984 : 4'b1000;
														assign node17984 = (inp[10]) ? 4'b1000 : 4'b0000;
										assign node17987 = (inp[4]) ? node17989 : 4'b1000;
											assign node17989 = (inp[13]) ? node18011 : node17990;
												assign node17990 = (inp[10]) ? node18000 : node17991;
													assign node17991 = (inp[1]) ? node17993 : 4'b1000;
														assign node17993 = (inp[12]) ? 4'b1000 : node17994;
															assign node17994 = (inp[11]) ? 4'b0000 : node17995;
																assign node17995 = (inp[14]) ? 4'b1000 : 4'b0000;
													assign node18000 = (inp[12]) ? node18008 : node18001;
														assign node18001 = (inp[14]) ? node18003 : 4'b0001;
															assign node18003 = (inp[11]) ? 4'b0000 : node18004;
																assign node18004 = (inp[1]) ? 4'b0001 : 4'b0000;
														assign node18008 = (inp[1]) ? 4'b0000 : 4'b1000;
												assign node18011 = (inp[1]) ? node18025 : node18012;
													assign node18012 = (inp[14]) ? node18018 : node18013;
														assign node18013 = (inp[10]) ? node18015 : 4'b0001;
															assign node18015 = (inp[11]) ? 4'b0001 : 4'b1001;
														assign node18018 = (inp[11]) ? 4'b0001 : node18019;
															assign node18019 = (inp[12]) ? 4'b0000 : node18020;
																assign node18020 = (inp[10]) ? 4'b1000 : 4'b0000;
													assign node18025 = (inp[12]) ? node18031 : node18026;
														assign node18026 = (inp[11]) ? 4'b1000 : node18027;
															assign node18027 = (inp[14]) ? 4'b1001 : 4'b1000;
														assign node18031 = (inp[10]) ? 4'b1000 : 4'b0000;
							assign node18035 = (inp[2]) ? node18447 : node18036;
								assign node18036 = (inp[3]) ? node18250 : node18037;
									assign node18037 = (inp[1]) ? node18145 : node18038;
										assign node18038 = (inp[13]) ? node18092 : node18039;
											assign node18039 = (inp[10]) ? node18057 : node18040;
												assign node18040 = (inp[11]) ? node18052 : node18041;
													assign node18041 = (inp[14]) ? node18047 : node18042;
														assign node18042 = (inp[7]) ? 4'b1001 : node18043;
															assign node18043 = (inp[4]) ? 4'b1101 : 4'b1001;
														assign node18047 = (inp[4]) ? node18049 : 4'b1000;
															assign node18049 = (inp[7]) ? 4'b1000 : 4'b1100;
													assign node18052 = (inp[4]) ? node18054 : 4'b1001;
														assign node18054 = (inp[7]) ? 4'b1001 : 4'b1101;
												assign node18057 = (inp[12]) ? node18083 : node18058;
													assign node18058 = (inp[14]) ? node18068 : node18059;
														assign node18059 = (inp[4]) ? node18063 : node18060;
															assign node18060 = (inp[7]) ? 4'b0001 : 4'b0101;
															assign node18063 = (inp[7]) ? 4'b0101 : node18064;
																assign node18064 = (inp[11]) ? 4'b1000 : 4'b0001;
														assign node18068 = (inp[11]) ? node18076 : node18069;
															assign node18069 = (inp[4]) ? node18073 : node18070;
																assign node18070 = (inp[7]) ? 4'b0000 : 4'b0100;
																assign node18073 = (inp[7]) ? 4'b0100 : 4'b0001;
															assign node18076 = (inp[4]) ? node18080 : node18077;
																assign node18077 = (inp[7]) ? 4'b0001 : 4'b0101;
																assign node18080 = (inp[7]) ? 4'b0101 : 4'b1000;
													assign node18083 = (inp[14]) ? node18085 : 4'b1001;
														assign node18085 = (inp[7]) ? node18089 : node18086;
															assign node18086 = (inp[4]) ? 4'b0000 : 4'b1000;
															assign node18089 = (inp[11]) ? 4'b1001 : 4'b1000;
											assign node18092 = (inp[4]) ? node18120 : node18093;
												assign node18093 = (inp[7]) ? node18111 : node18094;
													assign node18094 = (inp[12]) ? node18106 : node18095;
														assign node18095 = (inp[10]) ? node18101 : node18096;
															assign node18096 = (inp[14]) ? node18098 : 4'b0101;
																assign node18098 = (inp[11]) ? 4'b0101 : 4'b0100;
															assign node18101 = (inp[11]) ? 4'b1101 : node18102;
																assign node18102 = (inp[14]) ? 4'b1100 : 4'b1101;
														assign node18106 = (inp[11]) ? 4'b0101 : node18107;
															assign node18107 = (inp[14]) ? 4'b0100 : 4'b0101;
													assign node18111 = (inp[12]) ? node18115 : node18112;
														assign node18112 = (inp[10]) ? 4'b1001 : 4'b0001;
														assign node18115 = (inp[11]) ? 4'b0001 : node18116;
															assign node18116 = (inp[14]) ? 4'b0000 : 4'b0001;
												assign node18120 = (inp[11]) ? node18130 : node18121;
													assign node18121 = (inp[7]) ? node18125 : node18122;
														assign node18122 = (inp[10]) ? 4'b0001 : 4'b1001;
														assign node18125 = (inp[10]) ? 4'b0001 : node18126;
															assign node18126 = (inp[14]) ? 4'b0100 : 4'b0101;
													assign node18130 = (inp[7]) ? node18138 : node18131;
														assign node18131 = (inp[12]) ? node18135 : node18132;
															assign node18132 = (inp[10]) ? 4'b1000 : 4'b0000;
															assign node18135 = (inp[10]) ? 4'b0000 : 4'b1000;
														assign node18138 = (inp[10]) ? node18142 : node18139;
															assign node18139 = (inp[14]) ? 4'b0101 : 4'b0000;
															assign node18142 = (inp[14]) ? 4'b1000 : 4'b0000;
										assign node18145 = (inp[11]) ? node18213 : node18146;
											assign node18146 = (inp[14]) ? node18178 : node18147;
												assign node18147 = (inp[4]) ? node18165 : node18148;
													assign node18148 = (inp[7]) ? node18158 : node18149;
														assign node18149 = (inp[13]) ? node18155 : node18150;
															assign node18150 = (inp[12]) ? node18152 : 4'b0100;
																assign node18152 = (inp[10]) ? 4'b0100 : 4'b1000;
															assign node18155 = (inp[10]) ? 4'b1100 : 4'b0100;
														assign node18158 = (inp[13]) ? 4'b1000 : node18159;
															assign node18159 = (inp[12]) ? node18161 : 4'b0000;
																assign node18161 = (inp[10]) ? 4'b0000 : 4'b1000;
													assign node18165 = (inp[10]) ? node18175 : node18166;
														assign node18166 = (inp[13]) ? node18172 : node18167;
															assign node18167 = (inp[12]) ? node18169 : 4'b0100;
																assign node18169 = (inp[7]) ? 4'b1000 : 4'b1100;
															assign node18172 = (inp[7]) ? 4'b0100 : 4'b0001;
														assign node18175 = (inp[12]) ? 4'b0001 : 4'b1001;
												assign node18178 = (inp[13]) ? node18190 : node18179;
													assign node18179 = (inp[7]) ? node18185 : node18180;
														assign node18180 = (inp[4]) ? node18182 : 4'b1001;
															assign node18182 = (inp[10]) ? 4'b1001 : 4'b1101;
														assign node18185 = (inp[12]) ? 4'b1001 : node18186;
															assign node18186 = (inp[4]) ? 4'b0101 : 4'b0001;
													assign node18190 = (inp[4]) ? node18200 : node18191;
														assign node18191 = (inp[7]) ? node18197 : node18192;
															assign node18192 = (inp[10]) ? node18194 : 4'b0101;
																assign node18194 = (inp[12]) ? 4'b0101 : 4'b1101;
															assign node18197 = (inp[12]) ? 4'b0001 : 4'b1001;
														assign node18200 = (inp[7]) ? node18208 : node18201;
															assign node18201 = (inp[10]) ? node18205 : node18202;
																assign node18202 = (inp[12]) ? 4'b1001 : 4'b0001;
																assign node18205 = (inp[12]) ? 4'b0001 : 4'b1001;
															assign node18208 = (inp[12]) ? node18210 : 4'b0001;
																assign node18210 = (inp[10]) ? 4'b0001 : 4'b0101;
											assign node18213 = (inp[10]) ? node18237 : node18214;
												assign node18214 = (inp[4]) ? node18230 : node18215;
													assign node18215 = (inp[7]) ? node18223 : node18216;
														assign node18216 = (inp[13]) ? node18220 : node18217;
															assign node18217 = (inp[12]) ? 4'b1000 : 4'b0100;
															assign node18220 = (inp[12]) ? 4'b0100 : 4'b1100;
														assign node18223 = (inp[13]) ? node18227 : node18224;
															assign node18224 = (inp[12]) ? 4'b1000 : 4'b0000;
															assign node18227 = (inp[12]) ? 4'b0000 : 4'b1000;
													assign node18230 = (inp[13]) ? 4'b0000 : node18231;
														assign node18231 = (inp[7]) ? node18233 : 4'b0000;
															assign node18233 = (inp[14]) ? 4'b0100 : 4'b1000;
												assign node18237 = (inp[13]) ? node18245 : node18238;
													assign node18238 = (inp[7]) ? node18242 : node18239;
														assign node18239 = (inp[4]) ? 4'b1000 : 4'b0100;
														assign node18242 = (inp[4]) ? 4'b0100 : 4'b0000;
													assign node18245 = (inp[4]) ? 4'b1000 : node18246;
														assign node18246 = (inp[7]) ? 4'b1000 : 4'b1100;
									assign node18250 = (inp[4]) ? node18364 : node18251;
										assign node18251 = (inp[11]) ? node18321 : node18252;
											assign node18252 = (inp[13]) ? node18282 : node18253;
												assign node18253 = (inp[7]) ? node18271 : node18254;
													assign node18254 = (inp[1]) ? node18262 : node18255;
														assign node18255 = (inp[14]) ? 4'b1001 : node18256;
															assign node18256 = (inp[12]) ? 4'b1001 : node18257;
																assign node18257 = (inp[10]) ? 4'b1000 : 4'b0000;
														assign node18262 = (inp[14]) ? node18266 : node18263;
															assign node18263 = (inp[10]) ? 4'b1001 : 4'b0001;
															assign node18266 = (inp[12]) ? node18268 : 4'b0000;
																assign node18268 = (inp[10]) ? 4'b1000 : 4'b0000;
													assign node18271 = (inp[10]) ? node18277 : node18272;
														assign node18272 = (inp[1]) ? node18274 : 4'b1001;
															assign node18274 = (inp[12]) ? 4'b1001 : 4'b0001;
														assign node18277 = (inp[14]) ? node18279 : 4'b0001;
															assign node18279 = (inp[12]) ? 4'b0001 : 4'b0000;
												assign node18282 = (inp[14]) ? node18302 : node18283;
													assign node18283 = (inp[12]) ? node18291 : node18284;
														assign node18284 = (inp[1]) ? node18288 : node18285;
															assign node18285 = (inp[10]) ? 4'b0000 : 4'b1000;
															assign node18288 = (inp[10]) ? 4'b1000 : 4'b1001;
														assign node18291 = (inp[7]) ? node18297 : node18292;
															assign node18292 = (inp[1]) ? 4'b0000 : node18293;
																assign node18293 = (inp[10]) ? 4'b1000 : 4'b0000;
															assign node18297 = (inp[1]) ? node18299 : 4'b0000;
																assign node18299 = (inp[10]) ? 4'b0000 : 4'b1001;
													assign node18302 = (inp[7]) ? node18308 : node18303;
														assign node18303 = (inp[1]) ? 4'b0001 : node18304;
															assign node18304 = (inp[12]) ? 4'b0001 : 4'b0000;
														assign node18308 = (inp[1]) ? node18316 : node18309;
															assign node18309 = (inp[12]) ? node18313 : node18310;
																assign node18310 = (inp[10]) ? 4'b0000 : 4'b0001;
																assign node18313 = (inp[10]) ? 4'b1001 : 4'b0001;
															assign node18316 = (inp[10]) ? node18318 : 4'b1000;
																assign node18318 = (inp[12]) ? 4'b0000 : 4'b1000;
											assign node18321 = (inp[1]) ? node18349 : node18322;
												assign node18322 = (inp[13]) ? node18338 : node18323;
													assign node18323 = (inp[7]) ? node18331 : node18324;
														assign node18324 = (inp[12]) ? node18328 : node18325;
															assign node18325 = (inp[10]) ? 4'b1001 : 4'b0001;
															assign node18328 = (inp[10]) ? 4'b1001 : 4'b1000;
														assign node18331 = (inp[10]) ? node18335 : node18332;
															assign node18332 = (inp[12]) ? 4'b1000 : 4'b0000;
															assign node18335 = (inp[12]) ? 4'b0000 : 4'b1000;
													assign node18338 = (inp[7]) ? node18344 : node18339;
														assign node18339 = (inp[10]) ? node18341 : 4'b0000;
															assign node18341 = (inp[12]) ? 4'b0000 : 4'b0001;
														assign node18344 = (inp[10]) ? 4'b0000 : node18345;
															assign node18345 = (inp[12]) ? 4'b0001 : 4'b1001;
												assign node18349 = (inp[13]) ? node18357 : node18350;
													assign node18350 = (inp[10]) ? 4'b0000 : node18351;
														assign node18351 = (inp[7]) ? 4'b0000 : node18352;
															assign node18352 = (inp[12]) ? 4'b0000 : 4'b1000;
													assign node18357 = (inp[12]) ? 4'b1000 : node18358;
														assign node18358 = (inp[10]) ? 4'b1000 : node18359;
															assign node18359 = (inp[7]) ? 4'b0000 : 4'b1000;
										assign node18364 = (inp[13]) ? node18414 : node18365;
											assign node18365 = (inp[7]) ? node18395 : node18366;
												assign node18366 = (inp[11]) ? node18384 : node18367;
													assign node18367 = (inp[12]) ? node18375 : node18368;
														assign node18368 = (inp[14]) ? node18370 : 4'b0001;
															assign node18370 = (inp[1]) ? 4'b0000 : node18371;
																assign node18371 = (inp[10]) ? 4'b0000 : 4'b0001;
														assign node18375 = (inp[10]) ? node18381 : node18376;
															assign node18376 = (inp[1]) ? 4'b1001 : node18377;
																assign node18377 = (inp[14]) ? 4'b1000 : 4'b1001;
															assign node18381 = (inp[14]) ? 4'b0001 : 4'b0000;
													assign node18384 = (inp[12]) ? node18390 : node18385;
														assign node18385 = (inp[10]) ? node18387 : 4'b1000;
															assign node18387 = (inp[1]) ? 4'b0000 : 4'b0001;
														assign node18390 = (inp[10]) ? node18392 : 4'b0000;
															assign node18392 = (inp[1]) ? 4'b0000 : 4'b1000;
												assign node18395 = (inp[1]) ? node18407 : node18396;
													assign node18396 = (inp[11]) ? 4'b0001 : node18397;
														assign node18397 = (inp[14]) ? node18403 : node18398;
															assign node18398 = (inp[12]) ? 4'b0001 : node18399;
																assign node18399 = (inp[10]) ? 4'b0000 : 4'b0001;
															assign node18403 = (inp[12]) ? 4'b1000 : 4'b1001;
													assign node18407 = (inp[10]) ? 4'b0000 : node18408;
														assign node18408 = (inp[11]) ? 4'b0000 : node18409;
															assign node18409 = (inp[14]) ? 4'b0001 : 4'b1000;
											assign node18414 = (inp[11]) ? node18440 : node18415;
												assign node18415 = (inp[10]) ? node18431 : node18416;
													assign node18416 = (inp[7]) ? node18424 : node18417;
														assign node18417 = (inp[12]) ? 4'b0000 : node18418;
															assign node18418 = (inp[1]) ? 4'b0001 : node18419;
																assign node18419 = (inp[14]) ? 4'b0000 : 4'b0001;
														assign node18424 = (inp[12]) ? 4'b0001 : node18425;
															assign node18425 = (inp[1]) ? 4'b0000 : node18426;
																assign node18426 = (inp[14]) ? 4'b0001 : 4'b0000;
													assign node18431 = (inp[1]) ? 4'b0000 : node18432;
														assign node18432 = (inp[7]) ? 4'b0000 : node18433;
															assign node18433 = (inp[12]) ? node18435 : 4'b0001;
																assign node18435 = (inp[14]) ? 4'b0000 : 4'b0001;
												assign node18440 = (inp[7]) ? 4'b0000 : node18441;
													assign node18441 = (inp[10]) ? 4'b0000 : node18442;
														assign node18442 = (inp[1]) ? 4'b0000 : 4'b0001;
								assign node18447 = (inp[3]) ? node18449 : 4'b1000;
									assign node18449 = (inp[4]) ? node18507 : node18450;
										assign node18450 = (inp[7]) ? 4'b1000 : node18451;
											assign node18451 = (inp[13]) ? node18475 : node18452;
												assign node18452 = (inp[1]) ? node18458 : node18453;
													assign node18453 = (inp[12]) ? 4'b1000 : node18454;
														assign node18454 = (inp[10]) ? 4'b0001 : 4'b1000;
													assign node18458 = (inp[12]) ? node18470 : node18459;
														assign node18459 = (inp[10]) ? node18465 : node18460;
															assign node18460 = (inp[14]) ? node18462 : 4'b0000;
																assign node18462 = (inp[11]) ? 4'b0000 : 4'b1000;
															assign node18465 = (inp[14]) ? node18467 : 4'b0000;
																assign node18467 = (inp[11]) ? 4'b0000 : 4'b0001;
														assign node18470 = (inp[10]) ? node18472 : 4'b1000;
															assign node18472 = (inp[14]) ? 4'b1000 : 4'b0000;
												assign node18475 = (inp[1]) ? node18489 : node18476;
													assign node18476 = (inp[14]) ? node18482 : node18477;
														assign node18477 = (inp[12]) ? 4'b0001 : node18478;
															assign node18478 = (inp[10]) ? 4'b1001 : 4'b0001;
														assign node18482 = (inp[11]) ? 4'b0001 : node18483;
															assign node18483 = (inp[12]) ? 4'b0000 : node18484;
																assign node18484 = (inp[10]) ? 4'b1000 : 4'b0000;
													assign node18489 = (inp[14]) ? node18495 : node18490;
														assign node18490 = (inp[10]) ? 4'b1000 : node18491;
															assign node18491 = (inp[12]) ? 4'b0000 : 4'b1000;
														assign node18495 = (inp[11]) ? node18501 : node18496;
															assign node18496 = (inp[12]) ? 4'b0001 : node18497;
																assign node18497 = (inp[10]) ? 4'b1001 : 4'b0001;
															assign node18501 = (inp[10]) ? 4'b1000 : node18502;
																assign node18502 = (inp[12]) ? 4'b0000 : 4'b1000;
										assign node18507 = (inp[13]) ? node18561 : node18508;
											assign node18508 = (inp[10]) ? node18532 : node18509;
												assign node18509 = (inp[1]) ? node18521 : node18510;
													assign node18510 = (inp[7]) ? 4'b1000 : node18511;
														assign node18511 = (inp[12]) ? node18515 : node18512;
															assign node18512 = (inp[11]) ? 4'b0000 : 4'b1001;
															assign node18515 = (inp[11]) ? 4'b1001 : node18516;
																assign node18516 = (inp[14]) ? 4'b1000 : 4'b1001;
													assign node18521 = (inp[12]) ? node18527 : node18522;
														assign node18522 = (inp[11]) ? 4'b0000 : node18523;
															assign node18523 = (inp[7]) ? 4'b0000 : 4'b0001;
														assign node18527 = (inp[7]) ? 4'b1000 : node18528;
															assign node18528 = (inp[11]) ? 4'b0000 : 4'b1000;
												assign node18532 = (inp[11]) ? node18554 : node18533;
													assign node18533 = (inp[7]) ? node18541 : node18534;
														assign node18534 = (inp[14]) ? node18536 : 4'b0001;
															assign node18536 = (inp[12]) ? 4'b0001 : node18537;
																assign node18537 = (inp[1]) ? 4'b0000 : 4'b0001;
														assign node18541 = (inp[12]) ? node18549 : node18542;
															assign node18542 = (inp[14]) ? node18546 : node18543;
																assign node18543 = (inp[1]) ? 4'b0000 : 4'b0001;
																assign node18546 = (inp[1]) ? 4'b0001 : 4'b0000;
															assign node18549 = (inp[14]) ? 4'b1000 : node18550;
																assign node18550 = (inp[1]) ? 4'b0000 : 4'b1000;
													assign node18554 = (inp[1]) ? 4'b0000 : node18555;
														assign node18555 = (inp[7]) ? 4'b0001 : node18556;
															assign node18556 = (inp[12]) ? 4'b0000 : 4'b1000;
											assign node18561 = (inp[11]) ? node18589 : node18562;
												assign node18562 = (inp[14]) ? node18572 : node18563;
													assign node18563 = (inp[1]) ? 4'b0000 : node18564;
														assign node18564 = (inp[7]) ? 4'b0001 : node18565;
															assign node18565 = (inp[12]) ? 4'b0000 : node18566;
																assign node18566 = (inp[10]) ? 4'b0001 : 4'b0000;
													assign node18572 = (inp[10]) ? node18582 : node18573;
														assign node18573 = (inp[7]) ? 4'b0001 : node18574;
															assign node18574 = (inp[12]) ? node18578 : node18575;
																assign node18575 = (inp[1]) ? 4'b0001 : 4'b0000;
																assign node18578 = (inp[1]) ? 4'b0000 : 4'b0001;
														assign node18582 = (inp[7]) ? node18584 : 4'b0000;
															assign node18584 = (inp[1]) ? 4'b0000 : node18585;
																assign node18585 = (inp[12]) ? 4'b0001 : 4'b0000;
												assign node18589 = (inp[7]) ? node18591 : 4'b0000;
													assign node18591 = (inp[10]) ? 4'b0000 : node18592;
														assign node18592 = (inp[1]) ? 4'b0000 : node18593;
															assign node18593 = (inp[12]) ? 4'b0001 : 4'b0000;
			assign node18598 = (inp[15]) ? node21858 : node18599;
				assign node18599 = (inp[6]) ? node19375 : node18600;
					assign node18600 = (inp[0]) ? 4'b0100 : node18601;
						assign node18601 = (inp[2]) ? node19109 : node18602;
							assign node18602 = (inp[3]) ? node18894 : node18603;
								assign node18603 = (inp[5]) ? node18709 : node18604;
									assign node18604 = (inp[4]) ? node18632 : node18605;
										assign node18605 = (inp[7]) ? 4'b0110 : node18606;
											assign node18606 = (inp[13]) ? node18608 : 4'b0110;
												assign node18608 = (inp[12]) ? node18624 : node18609;
													assign node18609 = (inp[10]) ? node18617 : node18610;
														assign node18610 = (inp[1]) ? node18612 : 4'b0110;
															assign node18612 = (inp[14]) ? node18614 : 4'b0000;
																assign node18614 = (inp[11]) ? 4'b0000 : 4'b0110;
														assign node18617 = (inp[1]) ? 4'b0000 : node18618;
															assign node18618 = (inp[11]) ? 4'b0001 : node18619;
																assign node18619 = (inp[14]) ? 4'b0000 : 4'b0001;
													assign node18624 = (inp[1]) ? node18626 : 4'b0110;
														assign node18626 = (inp[10]) ? node18628 : 4'b0110;
															assign node18628 = (inp[14]) ? 4'b0110 : 4'b0000;
										assign node18632 = (inp[7]) ? node18688 : node18633;
											assign node18633 = (inp[1]) ? node18661 : node18634;
												assign node18634 = (inp[14]) ? node18646 : node18635;
													assign node18635 = (inp[13]) ? node18641 : node18636;
														assign node18636 = (inp[10]) ? node18638 : 4'b0001;
															assign node18638 = (inp[12]) ? 4'b0001 : 4'b1001;
														assign node18641 = (inp[12]) ? 4'b1001 : node18642;
															assign node18642 = (inp[10]) ? 4'b0001 : 4'b1001;
													assign node18646 = (inp[11]) ? node18656 : node18647;
														assign node18647 = (inp[13]) ? node18651 : node18648;
															assign node18648 = (inp[10]) ? 4'b1000 : 4'b0000;
															assign node18651 = (inp[10]) ? node18653 : 4'b1000;
																assign node18653 = (inp[12]) ? 4'b1000 : 4'b0000;
														assign node18656 = (inp[10]) ? 4'b0001 : node18657;
															assign node18657 = (inp[13]) ? 4'b1001 : 4'b0001;
												assign node18661 = (inp[11]) ? node18679 : node18662;
													assign node18662 = (inp[14]) ? node18670 : node18663;
														assign node18663 = (inp[13]) ? 4'b0000 : node18664;
															assign node18664 = (inp[12]) ? node18666 : 4'b1000;
																assign node18666 = (inp[10]) ? 4'b1000 : 4'b0000;
														assign node18670 = (inp[13]) ? node18676 : node18671;
															assign node18671 = (inp[12]) ? 4'b0001 : node18672;
																assign node18672 = (inp[10]) ? 4'b1001 : 4'b0001;
															assign node18676 = (inp[12]) ? 4'b1001 : 4'b0001;
													assign node18679 = (inp[13]) ? node18685 : node18680;
														assign node18680 = (inp[12]) ? node18682 : 4'b1000;
															assign node18682 = (inp[10]) ? 4'b1000 : 4'b0000;
														assign node18685 = (inp[10]) ? 4'b0000 : 4'b1000;
											assign node18688 = (inp[13]) ? node18690 : 4'b0110;
												assign node18690 = (inp[12]) ? node18702 : node18691;
													assign node18691 = (inp[10]) ? node18695 : node18692;
														assign node18692 = (inp[1]) ? 4'b0000 : 4'b0110;
														assign node18695 = (inp[1]) ? 4'b0000 : node18696;
															assign node18696 = (inp[14]) ? node18698 : 4'b0001;
																assign node18698 = (inp[11]) ? 4'b0001 : 4'b0000;
													assign node18702 = (inp[14]) ? 4'b0110 : node18703;
														assign node18703 = (inp[10]) ? node18705 : 4'b0110;
															assign node18705 = (inp[1]) ? 4'b0000 : 4'b0110;
									assign node18709 = (inp[1]) ? node18799 : node18710;
										assign node18710 = (inp[14]) ? node18748 : node18711;
											assign node18711 = (inp[7]) ? node18735 : node18712;
												assign node18712 = (inp[4]) ? node18724 : node18713;
													assign node18713 = (inp[13]) ? node18719 : node18714;
														assign node18714 = (inp[10]) ? node18716 : 4'b0101;
															assign node18716 = (inp[12]) ? 4'b0101 : 4'b1101;
														assign node18719 = (inp[12]) ? 4'b1101 : node18720;
															assign node18720 = (inp[10]) ? 4'b0001 : 4'b1101;
													assign node18724 = (inp[13]) ? node18730 : node18725;
														assign node18725 = (inp[10]) ? node18727 : 4'b0001;
															assign node18727 = (inp[12]) ? 4'b0001 : 4'b1001;
														assign node18730 = (inp[12]) ? 4'b1001 : node18731;
															assign node18731 = (inp[10]) ? 4'b0001 : 4'b1001;
												assign node18735 = (inp[13]) ? node18741 : node18736;
													assign node18736 = (inp[10]) ? node18738 : 4'b0101;
														assign node18738 = (inp[12]) ? 4'b0101 : 4'b1101;
													assign node18741 = (inp[12]) ? 4'b1101 : node18742;
														assign node18742 = (inp[10]) ? node18744 : 4'b1101;
															assign node18744 = (inp[4]) ? 4'b0001 : 4'b0101;
											assign node18748 = (inp[11]) ? node18772 : node18749;
												assign node18749 = (inp[13]) ? node18761 : node18750;
													assign node18750 = (inp[10]) ? node18756 : node18751;
														assign node18751 = (inp[7]) ? 4'b0100 : node18752;
															assign node18752 = (inp[4]) ? 4'b0000 : 4'b0100;
														assign node18756 = (inp[12]) ? 4'b0100 : node18757;
															assign node18757 = (inp[4]) ? 4'b1000 : 4'b1100;
													assign node18761 = (inp[12]) ? 4'b1100 : node18762;
														assign node18762 = (inp[10]) ? node18766 : node18763;
															assign node18763 = (inp[7]) ? 4'b1100 : 4'b1000;
															assign node18766 = (inp[4]) ? 4'b0000 : node18767;
																assign node18767 = (inp[7]) ? 4'b0100 : 4'b0000;
												assign node18772 = (inp[4]) ? node18784 : node18773;
													assign node18773 = (inp[13]) ? node18777 : node18774;
														assign node18774 = (inp[10]) ? 4'b1101 : 4'b0101;
														assign node18777 = (inp[10]) ? node18779 : 4'b1101;
															assign node18779 = (inp[12]) ? 4'b1101 : node18780;
																assign node18780 = (inp[7]) ? 4'b0101 : 4'b0001;
													assign node18784 = (inp[7]) ? node18794 : node18785;
														assign node18785 = (inp[10]) ? node18787 : 4'b1001;
															assign node18787 = (inp[12]) ? node18791 : node18788;
																assign node18788 = (inp[13]) ? 4'b0001 : 4'b1001;
																assign node18791 = (inp[13]) ? 4'b1001 : 4'b0001;
														assign node18794 = (inp[10]) ? 4'b0001 : node18795;
															assign node18795 = (inp[13]) ? 4'b1101 : 4'b0101;
										assign node18799 = (inp[7]) ? node18853 : node18800;
											assign node18800 = (inp[4]) ? node18824 : node18801;
												assign node18801 = (inp[13]) ? node18811 : node18802;
													assign node18802 = (inp[10]) ? 4'b1100 : node18803;
														assign node18803 = (inp[12]) ? 4'b0100 : node18804;
															assign node18804 = (inp[11]) ? 4'b1100 : node18805;
																assign node18805 = (inp[14]) ? 4'b0101 : 4'b1100;
													assign node18811 = (inp[12]) ? node18817 : node18812;
														assign node18812 = (inp[11]) ? 4'b0000 : node18813;
															assign node18813 = (inp[14]) ? 4'b0001 : 4'b0000;
														assign node18817 = (inp[10]) ? node18819 : 4'b1100;
															assign node18819 = (inp[14]) ? node18821 : 4'b0000;
																assign node18821 = (inp[11]) ? 4'b0000 : 4'b1101;
												assign node18824 = (inp[14]) ? node18836 : node18825;
													assign node18825 = (inp[13]) ? node18831 : node18826;
														assign node18826 = (inp[12]) ? node18828 : 4'b1000;
															assign node18828 = (inp[10]) ? 4'b1000 : 4'b0000;
														assign node18831 = (inp[10]) ? 4'b0000 : node18832;
															assign node18832 = (inp[12]) ? 4'b1000 : 4'b0000;
													assign node18836 = (inp[11]) ? node18846 : node18837;
														assign node18837 = (inp[10]) ? node18839 : 4'b0001;
															assign node18839 = (inp[13]) ? node18843 : node18840;
																assign node18840 = (inp[12]) ? 4'b0001 : 4'b1001;
																assign node18843 = (inp[12]) ? 4'b1001 : 4'b0001;
														assign node18846 = (inp[13]) ? node18848 : 4'b1000;
															assign node18848 = (inp[10]) ? 4'b0000 : node18849;
																assign node18849 = (inp[12]) ? 4'b1000 : 4'b0000;
											assign node18853 = (inp[11]) ? node18877 : node18854;
												assign node18854 = (inp[14]) ? node18864 : node18855;
													assign node18855 = (inp[4]) ? node18861 : node18856;
														assign node18856 = (inp[12]) ? 4'b0100 : node18857;
															assign node18857 = (inp[13]) ? 4'b0100 : 4'b1100;
														assign node18861 = (inp[13]) ? 4'b0000 : 4'b0100;
													assign node18864 = (inp[13]) ? node18870 : node18865;
														assign node18865 = (inp[12]) ? 4'b0101 : node18866;
															assign node18866 = (inp[10]) ? 4'b1101 : 4'b0101;
														assign node18870 = (inp[10]) ? node18872 : 4'b1101;
															assign node18872 = (inp[12]) ? 4'b1101 : node18873;
																assign node18873 = (inp[4]) ? 4'b0001 : 4'b0101;
												assign node18877 = (inp[13]) ? node18883 : node18878;
													assign node18878 = (inp[12]) ? node18880 : 4'b1100;
														assign node18880 = (inp[10]) ? 4'b1100 : 4'b0100;
													assign node18883 = (inp[4]) ? node18889 : node18884;
														assign node18884 = (inp[10]) ? 4'b0100 : node18885;
															assign node18885 = (inp[12]) ? 4'b1100 : 4'b0100;
														assign node18889 = (inp[12]) ? node18891 : 4'b0000;
															assign node18891 = (inp[10]) ? 4'b0000 : 4'b1100;
								assign node18894 = (inp[4]) ? node18986 : node18895;
									assign node18895 = (inp[1]) ? node18937 : node18896;
										assign node18896 = (inp[11]) ? node18924 : node18897;
											assign node18897 = (inp[14]) ? node18911 : node18898;
												assign node18898 = (inp[13]) ? node18904 : node18899;
													assign node18899 = (inp[12]) ? 4'b0001 : node18900;
														assign node18900 = (inp[10]) ? 4'b1001 : 4'b0001;
													assign node18904 = (inp[12]) ? 4'b1001 : node18905;
														assign node18905 = (inp[10]) ? node18907 : 4'b1001;
															assign node18907 = (inp[7]) ? 4'b0001 : 4'b0101;
												assign node18911 = (inp[13]) ? node18917 : node18912;
													assign node18912 = (inp[12]) ? 4'b0000 : node18913;
														assign node18913 = (inp[10]) ? 4'b1000 : 4'b0000;
													assign node18917 = (inp[10]) ? node18919 : 4'b1000;
														assign node18919 = (inp[12]) ? 4'b1000 : node18920;
															assign node18920 = (inp[7]) ? 4'b0000 : 4'b0100;
											assign node18924 = (inp[13]) ? node18930 : node18925;
												assign node18925 = (inp[12]) ? 4'b0001 : node18926;
													assign node18926 = (inp[10]) ? 4'b1001 : 4'b0001;
												assign node18930 = (inp[12]) ? 4'b1001 : node18931;
													assign node18931 = (inp[10]) ? node18933 : 4'b1001;
														assign node18933 = (inp[7]) ? 4'b0001 : 4'b0101;
										assign node18937 = (inp[14]) ? node18955 : node18938;
											assign node18938 = (inp[13]) ? node18944 : node18939;
												assign node18939 = (inp[12]) ? node18941 : 4'b1000;
													assign node18941 = (inp[10]) ? 4'b1000 : 4'b0000;
												assign node18944 = (inp[7]) ? node18950 : node18945;
													assign node18945 = (inp[12]) ? node18947 : 4'b0100;
														assign node18947 = (inp[10]) ? 4'b0100 : 4'b1000;
													assign node18950 = (inp[12]) ? node18952 : 4'b0000;
														assign node18952 = (inp[10]) ? 4'b0000 : 4'b1000;
											assign node18955 = (inp[11]) ? node18969 : node18956;
												assign node18956 = (inp[13]) ? node18962 : node18957;
													assign node18957 = (inp[12]) ? 4'b0001 : node18958;
														assign node18958 = (inp[10]) ? 4'b1001 : 4'b0001;
													assign node18962 = (inp[10]) ? node18964 : 4'b1001;
														assign node18964 = (inp[7]) ? node18966 : 4'b0101;
															assign node18966 = (inp[5]) ? 4'b0001 : 4'b1001;
												assign node18969 = (inp[13]) ? node18975 : node18970;
													assign node18970 = (inp[12]) ? node18972 : 4'b1000;
														assign node18972 = (inp[10]) ? 4'b1000 : 4'b0000;
													assign node18975 = (inp[7]) ? node18981 : node18976;
														assign node18976 = (inp[10]) ? 4'b0100 : node18977;
															assign node18977 = (inp[12]) ? 4'b1000 : 4'b0100;
														assign node18981 = (inp[10]) ? 4'b0000 : node18982;
															assign node18982 = (inp[12]) ? 4'b1000 : 4'b0000;
									assign node18986 = (inp[7]) ? node19050 : node18987;
										assign node18987 = (inp[1]) ? node19021 : node18988;
											assign node18988 = (inp[14]) ? node19000 : node18989;
												assign node18989 = (inp[13]) ? node18995 : node18990;
													assign node18990 = (inp[12]) ? 4'b0101 : node18991;
														assign node18991 = (inp[10]) ? 4'b1101 : 4'b0101;
													assign node18995 = (inp[10]) ? node18997 : 4'b1101;
														assign node18997 = (inp[12]) ? 4'b1101 : 4'b0101;
												assign node19000 = (inp[11]) ? node19012 : node19001;
													assign node19001 = (inp[13]) ? node19007 : node19002;
														assign node19002 = (inp[10]) ? node19004 : 4'b0100;
															assign node19004 = (inp[12]) ? 4'b0100 : 4'b1100;
														assign node19007 = (inp[12]) ? 4'b1100 : node19008;
															assign node19008 = (inp[10]) ? 4'b0100 : 4'b1100;
													assign node19012 = (inp[13]) ? node19018 : node19013;
														assign node19013 = (inp[12]) ? 4'b0101 : node19014;
															assign node19014 = (inp[10]) ? 4'b1101 : 4'b0101;
														assign node19018 = (inp[10]) ? 4'b0101 : 4'b1101;
											assign node19021 = (inp[11]) ? node19039 : node19022;
												assign node19022 = (inp[14]) ? node19028 : node19023;
													assign node19023 = (inp[13]) ? 4'b0100 : node19024;
														assign node19024 = (inp[12]) ? 4'b0100 : 4'b1100;
													assign node19028 = (inp[13]) ? node19034 : node19029;
														assign node19029 = (inp[10]) ? node19031 : 4'b0101;
															assign node19031 = (inp[12]) ? 4'b0101 : 4'b1101;
														assign node19034 = (inp[10]) ? node19036 : 4'b1101;
															assign node19036 = (inp[12]) ? 4'b1101 : 4'b0101;
												assign node19039 = (inp[13]) ? node19045 : node19040;
													assign node19040 = (inp[12]) ? node19042 : 4'b1100;
														assign node19042 = (inp[10]) ? 4'b1100 : 4'b0100;
													assign node19045 = (inp[12]) ? node19047 : 4'b0100;
														assign node19047 = (inp[10]) ? 4'b0100 : 4'b1100;
										assign node19050 = (inp[1]) ? node19080 : node19051;
											assign node19051 = (inp[13]) ? node19063 : node19052;
												assign node19052 = (inp[14]) ? node19058 : node19053;
													assign node19053 = (inp[12]) ? 4'b0001 : node19054;
														assign node19054 = (inp[10]) ? 4'b1001 : 4'b0001;
													assign node19058 = (inp[11]) ? 4'b0001 : node19059;
														assign node19059 = (inp[10]) ? 4'b1000 : 4'b0000;
												assign node19063 = (inp[10]) ? node19069 : node19064;
													assign node19064 = (inp[14]) ? node19066 : 4'b1001;
														assign node19066 = (inp[5]) ? 4'b1001 : 4'b1000;
													assign node19069 = (inp[12]) ? node19075 : node19070;
														assign node19070 = (inp[14]) ? node19072 : 4'b0101;
															assign node19072 = (inp[11]) ? 4'b0101 : 4'b0100;
														assign node19075 = (inp[5]) ? node19077 : 4'b1001;
															assign node19077 = (inp[14]) ? 4'b1000 : 4'b1001;
											assign node19080 = (inp[13]) ? node19096 : node19081;
												assign node19081 = (inp[12]) ? node19089 : node19082;
													assign node19082 = (inp[11]) ? 4'b1000 : node19083;
														assign node19083 = (inp[14]) ? node19085 : 4'b1000;
															assign node19085 = (inp[10]) ? 4'b1001 : 4'b0001;
													assign node19089 = (inp[11]) ? node19093 : node19090;
														assign node19090 = (inp[14]) ? 4'b0001 : 4'b0000;
														assign node19093 = (inp[10]) ? 4'b1000 : 4'b0000;
												assign node19096 = (inp[12]) ? node19102 : node19097;
													assign node19097 = (inp[14]) ? node19099 : 4'b0100;
														assign node19099 = (inp[11]) ? 4'b0100 : 4'b0101;
													assign node19102 = (inp[10]) ? 4'b0100 : node19103;
														assign node19103 = (inp[11]) ? 4'b1000 : node19104;
															assign node19104 = (inp[14]) ? 4'b1001 : 4'b1000;
							assign node19109 = (inp[5]) ? node19111 : 4'b0110;
								assign node19111 = (inp[3]) ? node19199 : node19112;
									assign node19112 = (inp[7]) ? node19180 : node19113;
										assign node19113 = (inp[4]) ? node19129 : node19114;
											assign node19114 = (inp[13]) ? node19116 : 4'b0110;
												assign node19116 = (inp[10]) ? node19122 : node19117;
													assign node19117 = (inp[1]) ? node19119 : 4'b0110;
														assign node19119 = (inp[11]) ? 4'b0000 : 4'b0110;
													assign node19122 = (inp[1]) ? node19124 : 4'b0001;
														assign node19124 = (inp[11]) ? 4'b0000 : node19125;
															assign node19125 = (inp[12]) ? 4'b0110 : 4'b0000;
											assign node19129 = (inp[1]) ? node19151 : node19130;
												assign node19130 = (inp[14]) ? node19142 : node19131;
													assign node19131 = (inp[13]) ? node19137 : node19132;
														assign node19132 = (inp[12]) ? 4'b0001 : node19133;
															assign node19133 = (inp[11]) ? 4'b1001 : 4'b0001;
														assign node19137 = (inp[12]) ? 4'b1001 : node19138;
															assign node19138 = (inp[10]) ? 4'b0001 : 4'b1001;
													assign node19142 = (inp[11]) ? 4'b1001 : node19143;
														assign node19143 = (inp[13]) ? 4'b1000 : node19144;
															assign node19144 = (inp[12]) ? 4'b0000 : node19145;
																assign node19145 = (inp[10]) ? 4'b1000 : 4'b0000;
												assign node19151 = (inp[14]) ? node19165 : node19152;
													assign node19152 = (inp[13]) ? node19158 : node19153;
														assign node19153 = (inp[12]) ? node19155 : 4'b1000;
															assign node19155 = (inp[10]) ? 4'b1000 : 4'b0000;
														assign node19158 = (inp[11]) ? 4'b0000 : node19159;
															assign node19159 = (inp[12]) ? node19161 : 4'b0000;
																assign node19161 = (inp[10]) ? 4'b0000 : 4'b1000;
													assign node19165 = (inp[11]) ? node19173 : node19166;
														assign node19166 = (inp[13]) ? 4'b1001 : node19167;
															assign node19167 = (inp[10]) ? node19169 : 4'b0001;
																assign node19169 = (inp[12]) ? 4'b0001 : 4'b1001;
														assign node19173 = (inp[13]) ? node19177 : node19174;
															assign node19174 = (inp[12]) ? 4'b0000 : 4'b1000;
															assign node19177 = (inp[12]) ? 4'b1000 : 4'b0000;
										assign node19180 = (inp[13]) ? node19182 : 4'b0110;
											assign node19182 = (inp[4]) ? node19184 : 4'b0110;
												assign node19184 = (inp[1]) ? node19190 : node19185;
													assign node19185 = (inp[10]) ? node19187 : 4'b0110;
														assign node19187 = (inp[12]) ? 4'b0110 : 4'b0001;
													assign node19190 = (inp[11]) ? 4'b0000 : node19191;
														assign node19191 = (inp[14]) ? 4'b0110 : node19192;
															assign node19192 = (inp[12]) ? node19194 : 4'b0000;
																assign node19194 = (inp[10]) ? 4'b0000 : 4'b0110;
									assign node19199 = (inp[1]) ? node19281 : node19200;
										assign node19200 = (inp[7]) ? node19246 : node19201;
											assign node19201 = (inp[4]) ? node19231 : node19202;
												assign node19202 = (inp[14]) ? node19214 : node19203;
													assign node19203 = (inp[13]) ? node19209 : node19204;
														assign node19204 = (inp[12]) ? 4'b0001 : node19205;
															assign node19205 = (inp[10]) ? 4'b1001 : 4'b0001;
														assign node19209 = (inp[12]) ? 4'b1001 : node19210;
															assign node19210 = (inp[10]) ? 4'b0101 : 4'b1001;
													assign node19214 = (inp[11]) ? node19222 : node19215;
														assign node19215 = (inp[12]) ? node19219 : node19216;
															assign node19216 = (inp[13]) ? 4'b0100 : 4'b1000;
															assign node19219 = (inp[13]) ? 4'b1000 : 4'b0000;
														assign node19222 = (inp[10]) ? node19224 : 4'b1001;
															assign node19224 = (inp[13]) ? node19228 : node19225;
																assign node19225 = (inp[12]) ? 4'b0001 : 4'b1001;
																assign node19228 = (inp[12]) ? 4'b1001 : 4'b0101;
												assign node19231 = (inp[13]) ? node19239 : node19232;
													assign node19232 = (inp[12]) ? 4'b0101 : node19233;
														assign node19233 = (inp[10]) ? node19235 : 4'b0101;
															assign node19235 = (inp[14]) ? 4'b1100 : 4'b1101;
													assign node19239 = (inp[12]) ? 4'b1101 : node19240;
														assign node19240 = (inp[10]) ? node19242 : 4'b1101;
															assign node19242 = (inp[14]) ? 4'b0100 : 4'b0101;
											assign node19246 = (inp[13]) ? node19262 : node19247;
												assign node19247 = (inp[11]) ? node19257 : node19248;
													assign node19248 = (inp[14]) ? node19252 : node19249;
														assign node19249 = (inp[10]) ? 4'b1001 : 4'b0001;
														assign node19252 = (inp[10]) ? node19254 : 4'b0000;
															assign node19254 = (inp[12]) ? 4'b0000 : 4'b1000;
													assign node19257 = (inp[12]) ? 4'b0001 : node19258;
														assign node19258 = (inp[10]) ? 4'b1001 : 4'b0001;
												assign node19262 = (inp[11]) ? node19274 : node19263;
													assign node19263 = (inp[14]) ? node19269 : node19264;
														assign node19264 = (inp[12]) ? 4'b1001 : node19265;
															assign node19265 = (inp[4]) ? 4'b1001 : 4'b0001;
														assign node19269 = (inp[10]) ? node19271 : 4'b1000;
															assign node19271 = (inp[12]) ? 4'b1000 : 4'b0000;
													assign node19274 = (inp[12]) ? 4'b1001 : node19275;
														assign node19275 = (inp[10]) ? node19277 : 4'b1001;
															assign node19277 = (inp[4]) ? 4'b0101 : 4'b0001;
										assign node19281 = (inp[4]) ? node19323 : node19282;
											assign node19282 = (inp[11]) ? node19310 : node19283;
												assign node19283 = (inp[14]) ? node19295 : node19284;
													assign node19284 = (inp[13]) ? node19290 : node19285;
														assign node19285 = (inp[10]) ? 4'b1000 : node19286;
															assign node19286 = (inp[12]) ? 4'b0000 : 4'b1000;
														assign node19290 = (inp[12]) ? 4'b1000 : node19291;
															assign node19291 = (inp[7]) ? 4'b0000 : 4'b0100;
													assign node19295 = (inp[10]) ? node19299 : node19296;
														assign node19296 = (inp[13]) ? 4'b1001 : 4'b0001;
														assign node19299 = (inp[7]) ? node19303 : node19300;
															assign node19300 = (inp[13]) ? 4'b0101 : 4'b0001;
															assign node19303 = (inp[12]) ? node19307 : node19304;
																assign node19304 = (inp[13]) ? 4'b0001 : 4'b1001;
																assign node19307 = (inp[13]) ? 4'b1001 : 4'b0001;
												assign node19310 = (inp[13]) ? node19316 : node19311;
													assign node19311 = (inp[10]) ? 4'b1000 : node19312;
														assign node19312 = (inp[12]) ? 4'b0000 : 4'b1000;
													assign node19316 = (inp[7]) ? 4'b0000 : node19317;
														assign node19317 = (inp[12]) ? node19319 : 4'b0100;
															assign node19319 = (inp[10]) ? 4'b0100 : 4'b1000;
											assign node19323 = (inp[7]) ? node19351 : node19324;
												assign node19324 = (inp[14]) ? node19336 : node19325;
													assign node19325 = (inp[13]) ? node19331 : node19326;
														assign node19326 = (inp[10]) ? 4'b1100 : node19327;
															assign node19327 = (inp[12]) ? 4'b0100 : 4'b1100;
														assign node19331 = (inp[10]) ? 4'b0100 : node19332;
															assign node19332 = (inp[12]) ? 4'b1100 : 4'b0100;
													assign node19336 = (inp[11]) ? node19344 : node19337;
														assign node19337 = (inp[13]) ? node19339 : 4'b0101;
															assign node19339 = (inp[12]) ? 4'b1101 : node19340;
																assign node19340 = (inp[10]) ? 4'b0101 : 4'b1101;
														assign node19344 = (inp[12]) ? node19346 : 4'b0100;
															assign node19346 = (inp[10]) ? node19348 : 4'b1100;
																assign node19348 = (inp[13]) ? 4'b0100 : 4'b1100;
												assign node19351 = (inp[13]) ? node19361 : node19352;
													assign node19352 = (inp[12]) ? node19354 : 4'b1000;
														assign node19354 = (inp[10]) ? 4'b1000 : node19355;
															assign node19355 = (inp[11]) ? 4'b0000 : node19356;
																assign node19356 = (inp[14]) ? 4'b0001 : 4'b0000;
													assign node19361 = (inp[12]) ? node19367 : node19362;
														assign node19362 = (inp[10]) ? node19364 : 4'b0100;
															assign node19364 = (inp[14]) ? 4'b0101 : 4'b0100;
														assign node19367 = (inp[10]) ? 4'b0100 : node19368;
															assign node19368 = (inp[11]) ? 4'b1000 : node19369;
																assign node19369 = (inp[14]) ? 4'b1001 : 4'b1000;
					assign node19375 = (inp[5]) ? node20395 : node19376;
						assign node19376 = (inp[0]) ? node20088 : node19377;
							assign node19377 = (inp[11]) ? node19769 : node19378;
								assign node19378 = (inp[4]) ? node19550 : node19379;
									assign node19379 = (inp[3]) ? node19471 : node19380;
										assign node19380 = (inp[13]) ? node19412 : node19381;
											assign node19381 = (inp[12]) ? node19403 : node19382;
												assign node19382 = (inp[10]) ? node19390 : node19383;
													assign node19383 = (inp[1]) ? node19387 : node19384;
														assign node19384 = (inp[14]) ? 4'b0100 : 4'b0101;
														assign node19387 = (inp[14]) ? 4'b0101 : 4'b1100;
													assign node19390 = (inp[2]) ? node19398 : node19391;
														assign node19391 = (inp[7]) ? node19395 : node19392;
															assign node19392 = (inp[1]) ? 4'b0001 : 4'b1100;
															assign node19395 = (inp[1]) ? 4'b1100 : 4'b1101;
														assign node19398 = (inp[1]) ? 4'b1100 : node19399;
															assign node19399 = (inp[14]) ? 4'b1100 : 4'b1101;
												assign node19403 = (inp[14]) ? node19409 : node19404;
													assign node19404 = (inp[1]) ? node19406 : 4'b0101;
														assign node19406 = (inp[10]) ? 4'b1100 : 4'b0100;
													assign node19409 = (inp[1]) ? 4'b0101 : 4'b0100;
											assign node19412 = (inp[12]) ? node19444 : node19413;
												assign node19413 = (inp[7]) ? node19431 : node19414;
													assign node19414 = (inp[10]) ? node19424 : node19415;
														assign node19415 = (inp[2]) ? node19419 : node19416;
															assign node19416 = (inp[1]) ? 4'b1001 : 4'b0001;
															assign node19419 = (inp[14]) ? 4'b1101 : node19420;
																assign node19420 = (inp[1]) ? 4'b0000 : 4'b1101;
														assign node19424 = (inp[14]) ? 4'b0001 : node19425;
															assign node19425 = (inp[1]) ? node19427 : 4'b0001;
																assign node19427 = (inp[2]) ? 4'b0000 : 4'b0001;
													assign node19431 = (inp[10]) ? node19437 : node19432;
														assign node19432 = (inp[14]) ? node19434 : 4'b0100;
															assign node19434 = (inp[1]) ? 4'b1101 : 4'b1100;
														assign node19437 = (inp[1]) ? node19441 : node19438;
															assign node19438 = (inp[14]) ? 4'b0100 : 4'b0101;
															assign node19441 = (inp[2]) ? 4'b0100 : 4'b0001;
												assign node19444 = (inp[2]) ? node19454 : node19445;
													assign node19445 = (inp[7]) ? node19449 : node19446;
														assign node19446 = (inp[10]) ? 4'b1001 : 4'b0001;
														assign node19449 = (inp[14]) ? 4'b1101 : node19450;
															assign node19450 = (inp[1]) ? 4'b1100 : 4'b1101;
													assign node19454 = (inp[10]) ? node19462 : node19455;
														assign node19455 = (inp[7]) ? 4'b1100 : node19456;
															assign node19456 = (inp[14]) ? node19458 : 4'b1100;
																assign node19458 = (inp[1]) ? 4'b1101 : 4'b1100;
														assign node19462 = (inp[1]) ? node19466 : node19463;
															assign node19463 = (inp[14]) ? 4'b1100 : 4'b1101;
															assign node19466 = (inp[14]) ? 4'b1101 : node19467;
																assign node19467 = (inp[7]) ? 4'b0100 : 4'b0000;
										assign node19471 = (inp[2]) ? node19505 : node19472;
											assign node19472 = (inp[7]) ? node19492 : node19473;
												assign node19473 = (inp[13]) ? node19485 : node19474;
													assign node19474 = (inp[10]) ? node19480 : node19475;
														assign node19475 = (inp[12]) ? 4'b0101 : node19476;
															assign node19476 = (inp[1]) ? 4'b1101 : 4'b0101;
														assign node19480 = (inp[1]) ? node19482 : 4'b1101;
															assign node19482 = (inp[12]) ? 4'b1101 : 4'b0001;
													assign node19485 = (inp[10]) ? 4'b1001 : node19486;
														assign node19486 = (inp[1]) ? node19488 : 4'b0001;
															assign node19488 = (inp[12]) ? 4'b0001 : 4'b1001;
												assign node19492 = (inp[10]) ? node19498 : node19493;
													assign node19493 = (inp[1]) ? node19495 : 4'b0101;
														assign node19495 = (inp[12]) ? 4'b0101 : 4'b1101;
													assign node19498 = (inp[12]) ? 4'b1101 : node19499;
														assign node19499 = (inp[1]) ? node19501 : 4'b1101;
															assign node19501 = (inp[13]) ? 4'b0001 : 4'b0101;
											assign node19505 = (inp[13]) ? node19523 : node19506;
												assign node19506 = (inp[14]) ? node19516 : node19507;
													assign node19507 = (inp[1]) ? node19511 : node19508;
														assign node19508 = (inp[10]) ? 4'b1001 : 4'b0001;
														assign node19511 = (inp[12]) ? node19513 : 4'b1000;
															assign node19513 = (inp[10]) ? 4'b1000 : 4'b0000;
													assign node19516 = (inp[1]) ? 4'b0001 : node19517;
														assign node19517 = (inp[12]) ? 4'b0000 : node19518;
															assign node19518 = (inp[10]) ? 4'b1000 : 4'b0000;
												assign node19523 = (inp[7]) ? node19531 : node19524;
													assign node19524 = (inp[10]) ? 4'b1001 : node19525;
														assign node19525 = (inp[1]) ? node19527 : 4'b0001;
															assign node19527 = (inp[12]) ? 4'b0001 : 4'b1001;
													assign node19531 = (inp[10]) ? node19541 : node19532;
														assign node19532 = (inp[14]) ? node19538 : node19533;
															assign node19533 = (inp[1]) ? node19535 : 4'b1001;
																assign node19535 = (inp[12]) ? 4'b1000 : 4'b0000;
															assign node19538 = (inp[1]) ? 4'b1001 : 4'b1000;
														assign node19541 = (inp[1]) ? node19545 : node19542;
															assign node19542 = (inp[12]) ? 4'b1000 : 4'b0000;
															assign node19545 = (inp[14]) ? node19547 : 4'b0000;
																assign node19547 = (inp[12]) ? 4'b1001 : 4'b0001;
									assign node19550 = (inp[13]) ? node19656 : node19551;
										assign node19551 = (inp[10]) ? node19603 : node19552;
											assign node19552 = (inp[1]) ? node19574 : node19553;
												assign node19553 = (inp[7]) ? node19567 : node19554;
													assign node19554 = (inp[14]) ? node19562 : node19555;
														assign node19555 = (inp[3]) ? node19557 : 4'b0001;
															assign node19557 = (inp[2]) ? 4'b0001 : node19558;
																assign node19558 = (inp[12]) ? 4'b0000 : 4'b1000;
														assign node19562 = (inp[3]) ? 4'b0001 : node19563;
															assign node19563 = (inp[2]) ? 4'b0000 : 4'b0001;
													assign node19567 = (inp[2]) ? node19569 : 4'b0001;
														assign node19569 = (inp[3]) ? 4'b0001 : node19570;
															assign node19570 = (inp[14]) ? 4'b0100 : 4'b0101;
												assign node19574 = (inp[12]) ? node19584 : node19575;
													assign node19575 = (inp[2]) ? node19577 : 4'b1001;
														assign node19577 = (inp[3]) ? 4'b1001 : node19578;
															assign node19578 = (inp[14]) ? node19580 : 4'b1100;
																assign node19580 = (inp[7]) ? 4'b0101 : 4'b0001;
													assign node19584 = (inp[7]) ? node19596 : node19585;
														assign node19585 = (inp[2]) ? node19591 : node19586;
															assign node19586 = (inp[3]) ? node19588 : 4'b0001;
																assign node19588 = (inp[14]) ? 4'b1000 : 4'b1001;
															assign node19591 = (inp[3]) ? 4'b0001 : node19592;
																assign node19592 = (inp[14]) ? 4'b0001 : 4'b0000;
														assign node19596 = (inp[2]) ? node19598 : 4'b0001;
															assign node19598 = (inp[3]) ? 4'b0001 : node19599;
																assign node19599 = (inp[14]) ? 4'b0101 : 4'b0100;
											assign node19603 = (inp[2]) ? node19625 : node19604;
												assign node19604 = (inp[3]) ? node19612 : node19605;
													assign node19605 = (inp[12]) ? 4'b1001 : node19606;
														assign node19606 = (inp[1]) ? node19608 : 4'b1001;
															assign node19608 = (inp[14]) ? 4'b0001 : 4'b0101;
													assign node19612 = (inp[14]) ? node19618 : node19613;
														assign node19613 = (inp[1]) ? node19615 : 4'b0000;
															assign node19615 = (inp[12]) ? 4'b0001 : 4'b1001;
														assign node19618 = (inp[1]) ? node19622 : node19619;
															assign node19619 = (inp[12]) ? 4'b1001 : 4'b0001;
															assign node19622 = (inp[12]) ? 4'b0000 : 4'b1000;
												assign node19625 = (inp[3]) ? node19649 : node19626;
													assign node19626 = (inp[7]) ? node19638 : node19627;
														assign node19627 = (inp[12]) ? node19633 : node19628;
															assign node19628 = (inp[1]) ? 4'b1001 : node19629;
																assign node19629 = (inp[14]) ? 4'b1000 : 4'b1001;
															assign node19633 = (inp[1]) ? 4'b0001 : node19634;
																assign node19634 = (inp[14]) ? 4'b0000 : 4'b0001;
														assign node19638 = (inp[12]) ? node19646 : node19639;
															assign node19639 = (inp[1]) ? node19643 : node19640;
																assign node19640 = (inp[14]) ? 4'b1100 : 4'b1101;
																assign node19643 = (inp[14]) ? 4'b1101 : 4'b1100;
															assign node19646 = (inp[1]) ? 4'b0101 : 4'b0100;
													assign node19649 = (inp[1]) ? node19651 : 4'b1001;
														assign node19651 = (inp[12]) ? 4'b1001 : node19652;
															assign node19652 = (inp[7]) ? 4'b0001 : 4'b0101;
										assign node19656 = (inp[7]) ? node19714 : node19657;
											assign node19657 = (inp[2]) ? node19677 : node19658;
												assign node19658 = (inp[3]) ? node19666 : node19659;
													assign node19659 = (inp[10]) ? node19661 : 4'b0101;
														assign node19661 = (inp[1]) ? node19663 : 4'b1101;
															assign node19663 = (inp[12]) ? 4'b1101 : 4'b0101;
													assign node19666 = (inp[1]) ? 4'b0100 : node19667;
														assign node19667 = (inp[14]) ? node19673 : node19668;
															assign node19668 = (inp[12]) ? 4'b1000 : node19669;
																assign node19669 = (inp[10]) ? 4'b1100 : 4'b0100;
															assign node19673 = (inp[10]) ? 4'b1101 : 4'b1001;
												assign node19677 = (inp[3]) ? node19703 : node19678;
													assign node19678 = (inp[12]) ? node19692 : node19679;
														assign node19679 = (inp[10]) ? node19685 : node19680;
															assign node19680 = (inp[14]) ? 4'b1001 : node19681;
																assign node19681 = (inp[1]) ? 4'b0000 : 4'b1001;
															assign node19685 = (inp[14]) ? node19689 : node19686;
																assign node19686 = (inp[1]) ? 4'b0000 : 4'b0001;
																assign node19689 = (inp[1]) ? 4'b0001 : 4'b0000;
														assign node19692 = (inp[10]) ? node19698 : node19693;
															assign node19693 = (inp[1]) ? 4'b1000 : node19694;
																assign node19694 = (inp[14]) ? 4'b1000 : 4'b1001;
															assign node19698 = (inp[14]) ? node19700 : 4'b0000;
																assign node19700 = (inp[1]) ? 4'b1001 : 4'b1000;
													assign node19703 = (inp[10]) ? node19709 : node19704;
														assign node19704 = (inp[1]) ? node19706 : 4'b0101;
															assign node19706 = (inp[12]) ? 4'b0101 : 4'b1101;
														assign node19709 = (inp[1]) ? node19711 : 4'b1101;
															assign node19711 = (inp[12]) ? 4'b1101 : 4'b0101;
											assign node19714 = (inp[2]) ? node19740 : node19715;
												assign node19715 = (inp[3]) ? node19723 : node19716;
													assign node19716 = (inp[10]) ? 4'b1001 : node19717;
														assign node19717 = (inp[1]) ? node19719 : 4'b0001;
															assign node19719 = (inp[12]) ? 4'b0001 : 4'b1001;
													assign node19723 = (inp[1]) ? node19733 : node19724;
														assign node19724 = (inp[14]) ? node19730 : node19725;
															assign node19725 = (inp[12]) ? 4'b1000 : node19726;
																assign node19726 = (inp[10]) ? 4'b1000 : 4'b0000;
															assign node19730 = (inp[12]) ? 4'b0001 : 4'b1001;
														assign node19733 = (inp[14]) ? node19737 : node19734;
															assign node19734 = (inp[10]) ? 4'b1001 : 4'b0001;
															assign node19737 = (inp[10]) ? 4'b0100 : 4'b0000;
												assign node19740 = (inp[3]) ? node19758 : node19741;
													assign node19741 = (inp[12]) ? node19751 : node19742;
														assign node19742 = (inp[10]) ? node19746 : node19743;
															assign node19743 = (inp[14]) ? 4'b1100 : 4'b1101;
															assign node19746 = (inp[14]) ? 4'b0001 : node19747;
																assign node19747 = (inp[1]) ? 4'b0000 : 4'b0001;
														assign node19751 = (inp[14]) ? node19755 : node19752;
															assign node19752 = (inp[1]) ? 4'b1100 : 4'b1101;
															assign node19755 = (inp[1]) ? 4'b1101 : 4'b1100;
													assign node19758 = (inp[10]) ? node19764 : node19759;
														assign node19759 = (inp[1]) ? node19761 : 4'b0001;
															assign node19761 = (inp[12]) ? 4'b0001 : 4'b1001;
														assign node19764 = (inp[12]) ? 4'b1001 : node19765;
															assign node19765 = (inp[1]) ? 4'b0101 : 4'b1001;
								assign node19769 = (inp[1]) ? node19953 : node19770;
									assign node19770 = (inp[3]) ? node19860 : node19771;
										assign node19771 = (inp[2]) ? node19827 : node19772;
											assign node19772 = (inp[4]) ? node19792 : node19773;
												assign node19773 = (inp[13]) ? node19781 : node19774;
													assign node19774 = (inp[10]) ? node19776 : 4'b0101;
														assign node19776 = (inp[12]) ? 4'b0101 : node19777;
															assign node19777 = (inp[7]) ? 4'b1101 : 4'b0000;
													assign node19781 = (inp[7]) ? node19787 : node19782;
														assign node19782 = (inp[12]) ? 4'b1000 : node19783;
															assign node19783 = (inp[10]) ? 4'b0000 : 4'b1000;
														assign node19787 = (inp[10]) ? node19789 : 4'b1101;
															assign node19789 = (inp[12]) ? 4'b1101 : 4'b0000;
												assign node19792 = (inp[13]) ? node19812 : node19793;
													assign node19793 = (inp[7]) ? node19801 : node19794;
														assign node19794 = (inp[12]) ? node19798 : node19795;
															assign node19795 = (inp[10]) ? 4'b0100 : 4'b1000;
															assign node19798 = (inp[10]) ? 4'b1000 : 4'b0000;
														assign node19801 = (inp[14]) ? node19807 : node19802;
															assign node19802 = (inp[12]) ? 4'b0000 : node19803;
																assign node19803 = (inp[10]) ? 4'b0000 : 4'b1000;
															assign node19807 = (inp[12]) ? node19809 : 4'b0000;
																assign node19809 = (inp[10]) ? 4'b1000 : 4'b0000;
													assign node19812 = (inp[7]) ? node19820 : node19813;
														assign node19813 = (inp[10]) ? node19817 : node19814;
															assign node19814 = (inp[12]) ? 4'b0100 : 4'b1100;
															assign node19817 = (inp[12]) ? 4'b1100 : 4'b0100;
														assign node19820 = (inp[12]) ? node19824 : node19821;
															assign node19821 = (inp[10]) ? 4'b0100 : 4'b1000;
															assign node19824 = (inp[10]) ? 4'b1000 : 4'b0000;
											assign node19827 = (inp[13]) ? node19841 : node19828;
												assign node19828 = (inp[10]) ? node19834 : node19829;
													assign node19829 = (inp[4]) ? node19831 : 4'b0101;
														assign node19831 = (inp[7]) ? 4'b0101 : 4'b0001;
													assign node19834 = (inp[12]) ? node19836 : 4'b1101;
														assign node19836 = (inp[7]) ? 4'b0101 : node19837;
															assign node19837 = (inp[4]) ? 4'b0001 : 4'b0101;
												assign node19841 = (inp[7]) ? node19853 : node19842;
													assign node19842 = (inp[4]) ? node19848 : node19843;
														assign node19843 = (inp[12]) ? 4'b1101 : node19844;
															assign node19844 = (inp[10]) ? 4'b0001 : 4'b1101;
														assign node19848 = (inp[10]) ? node19850 : 4'b1001;
															assign node19850 = (inp[14]) ? 4'b0001 : 4'b1001;
													assign node19853 = (inp[10]) ? node19855 : 4'b1101;
														assign node19855 = (inp[12]) ? 4'b1101 : node19856;
															assign node19856 = (inp[4]) ? 4'b0001 : 4'b0101;
										assign node19860 = (inp[2]) ? node19908 : node19861;
											assign node19861 = (inp[4]) ? node19887 : node19862;
												assign node19862 = (inp[13]) ? node19872 : node19863;
													assign node19863 = (inp[12]) ? node19869 : node19864;
														assign node19864 = (inp[10]) ? node19866 : 4'b1100;
															assign node19866 = (inp[7]) ? 4'b0100 : 4'b0000;
														assign node19869 = (inp[10]) ? 4'b1100 : 4'b0100;
													assign node19872 = (inp[7]) ? node19880 : node19873;
														assign node19873 = (inp[10]) ? node19877 : node19874;
															assign node19874 = (inp[12]) ? 4'b0000 : 4'b1000;
															assign node19877 = (inp[12]) ? 4'b1000 : 4'b0000;
														assign node19880 = (inp[10]) ? node19884 : node19881;
															assign node19881 = (inp[12]) ? 4'b0100 : 4'b1100;
															assign node19884 = (inp[12]) ? 4'b1100 : 4'b0000;
												assign node19887 = (inp[13]) ? node19897 : node19888;
													assign node19888 = (inp[10]) ? 4'b0001 : node19889;
														assign node19889 = (inp[12]) ? node19893 : node19890;
															assign node19890 = (inp[7]) ? 4'b1000 : 4'b1001;
															assign node19893 = (inp[7]) ? 4'b0000 : 4'b0001;
													assign node19897 = (inp[7]) ? node19903 : node19898;
														assign node19898 = (inp[12]) ? node19900 : 4'b0101;
															assign node19900 = (inp[10]) ? 4'b1101 : 4'b1001;
														assign node19903 = (inp[10]) ? 4'b1001 : node19904;
															assign node19904 = (inp[12]) ? 4'b1001 : 4'b0001;
											assign node19908 = (inp[4]) ? node19930 : node19909;
												assign node19909 = (inp[13]) ? node19917 : node19910;
													assign node19910 = (inp[10]) ? node19912 : 4'b0001;
														assign node19912 = (inp[12]) ? 4'b0001 : node19913;
															assign node19913 = (inp[7]) ? 4'b1001 : 4'b0000;
													assign node19917 = (inp[7]) ? node19927 : node19918;
														assign node19918 = (inp[14]) ? node19924 : node19919;
															assign node19919 = (inp[12]) ? 4'b0000 : node19920;
																assign node19920 = (inp[10]) ? 4'b0000 : 4'b1000;
															assign node19924 = (inp[12]) ? 4'b1000 : 4'b0000;
														assign node19927 = (inp[10]) ? 4'b0000 : 4'b1001;
												assign node19930 = (inp[7]) ? node19944 : node19931;
													assign node19931 = (inp[13]) ? node19939 : node19932;
														assign node19932 = (inp[10]) ? node19936 : node19933;
															assign node19933 = (inp[12]) ? 4'b0000 : 4'b1000;
															assign node19936 = (inp[12]) ? 4'b1000 : 4'b0100;
														assign node19939 = (inp[12]) ? 4'b0100 : node19940;
															assign node19940 = (inp[10]) ? 4'b0100 : 4'b1100;
													assign node19944 = (inp[12]) ? node19950 : node19945;
														assign node19945 = (inp[10]) ? node19947 : 4'b1000;
															assign node19947 = (inp[13]) ? 4'b0100 : 4'b0000;
														assign node19950 = (inp[10]) ? 4'b1000 : 4'b0000;
									assign node19953 = (inp[10]) ? node20037 : node19954;
										assign node19954 = (inp[4]) ? node19994 : node19955;
											assign node19955 = (inp[3]) ? node19971 : node19956;
												assign node19956 = (inp[13]) ? node19960 : node19957;
													assign node19957 = (inp[12]) ? 4'b0100 : 4'b1100;
													assign node19960 = (inp[12]) ? node19966 : node19961;
														assign node19961 = (inp[7]) ? 4'b0100 : node19962;
															assign node19962 = (inp[2]) ? 4'b0000 : 4'b1000;
														assign node19966 = (inp[7]) ? 4'b1100 : node19967;
															assign node19967 = (inp[2]) ? 4'b1100 : 4'b1000;
												assign node19971 = (inp[2]) ? node19977 : node19972;
													assign node19972 = (inp[7]) ? 4'b1100 : node19973;
														assign node19973 = (inp[13]) ? 4'b1000 : 4'b1100;
													assign node19977 = (inp[7]) ? node19983 : node19978;
														assign node19978 = (inp[12]) ? node19980 : 4'b1000;
															assign node19980 = (inp[13]) ? 4'b1000 : 4'b0000;
														assign node19983 = (inp[14]) ? node19989 : node19984;
															assign node19984 = (inp[13]) ? node19986 : 4'b1000;
																assign node19986 = (inp[12]) ? 4'b1000 : 4'b0000;
															assign node19989 = (inp[12]) ? 4'b0000 : node19990;
																assign node19990 = (inp[13]) ? 4'b0000 : 4'b1000;
											assign node19994 = (inp[13]) ? node20010 : node19995;
												assign node19995 = (inp[2]) ? node20001 : node19996;
													assign node19996 = (inp[3]) ? node19998 : 4'b1000;
														assign node19998 = (inp[12]) ? 4'b1000 : 4'b0000;
													assign node20001 = (inp[3]) ? 4'b1000 : node20002;
														assign node20002 = (inp[7]) ? node20006 : node20003;
															assign node20003 = (inp[12]) ? 4'b0000 : 4'b1000;
															assign node20006 = (inp[12]) ? 4'b0100 : 4'b1100;
												assign node20010 = (inp[7]) ? node20022 : node20011;
													assign node20011 = (inp[3]) ? node20017 : node20012;
														assign node20012 = (inp[2]) ? node20014 : 4'b1100;
															assign node20014 = (inp[12]) ? 4'b1000 : 4'b0000;
														assign node20017 = (inp[2]) ? 4'b1100 : node20018;
															assign node20018 = (inp[12]) ? 4'b0100 : 4'b1100;
													assign node20022 = (inp[14]) ? node20030 : node20023;
														assign node20023 = (inp[3]) ? node20027 : node20024;
															assign node20024 = (inp[12]) ? 4'b1000 : 4'b0000;
															assign node20027 = (inp[2]) ? 4'b1000 : 4'b0000;
														assign node20030 = (inp[12]) ? node20032 : 4'b1000;
															assign node20032 = (inp[2]) ? 4'b1000 : node20033;
																assign node20033 = (inp[3]) ? 4'b0000 : 4'b1000;
										assign node20037 = (inp[13]) ? node20075 : node20038;
											assign node20038 = (inp[7]) ? node20062 : node20039;
												assign node20039 = (inp[4]) ? node20045 : node20040;
													assign node20040 = (inp[2]) ? node20042 : 4'b0000;
														assign node20042 = (inp[3]) ? 4'b0000 : 4'b1100;
													assign node20045 = (inp[12]) ? node20053 : node20046;
														assign node20046 = (inp[2]) ? node20050 : node20047;
															assign node20047 = (inp[3]) ? 4'b1000 : 4'b0100;
															assign node20050 = (inp[3]) ? 4'b0100 : 4'b1000;
														assign node20053 = (inp[14]) ? 4'b0100 : node20054;
															assign node20054 = (inp[2]) ? node20058 : node20055;
																assign node20055 = (inp[3]) ? 4'b1000 : 4'b0100;
																assign node20058 = (inp[3]) ? 4'b0100 : 4'b1000;
												assign node20062 = (inp[4]) ? node20068 : node20063;
													assign node20063 = (inp[3]) ? node20065 : 4'b1100;
														assign node20065 = (inp[2]) ? 4'b1000 : 4'b0100;
													assign node20068 = (inp[2]) ? node20072 : node20069;
														assign node20069 = (inp[3]) ? 4'b1000 : 4'b0000;
														assign node20072 = (inp[3]) ? 4'b0000 : 4'b1100;
											assign node20075 = (inp[4]) ? node20083 : node20076;
												assign node20076 = (inp[2]) ? node20078 : 4'b0000;
													assign node20078 = (inp[3]) ? 4'b0000 : node20079;
														assign node20079 = (inp[7]) ? 4'b0100 : 4'b0000;
												assign node20083 = (inp[3]) ? 4'b0100 : node20084;
													assign node20084 = (inp[2]) ? 4'b0000 : 4'b0100;
							assign node20088 = (inp[2]) ? 4'b0100 : node20089;
								assign node20089 = (inp[3]) ? node20203 : node20090;
									assign node20090 = (inp[4]) ? node20118 : node20091;
										assign node20091 = (inp[13]) ? node20093 : 4'b0100;
											assign node20093 = (inp[7]) ? 4'b0100 : node20094;
												assign node20094 = (inp[10]) ? node20102 : node20095;
													assign node20095 = (inp[11]) ? node20097 : 4'b0100;
														assign node20097 = (inp[1]) ? node20099 : 4'b0100;
															assign node20099 = (inp[14]) ? 4'b0000 : 4'b0100;
													assign node20102 = (inp[12]) ? node20114 : node20103;
														assign node20103 = (inp[1]) ? node20109 : node20104;
															assign node20104 = (inp[11]) ? 4'b0001 : node20105;
																assign node20105 = (inp[14]) ? 4'b0000 : 4'b0001;
															assign node20109 = (inp[11]) ? 4'b0000 : node20110;
																assign node20110 = (inp[14]) ? 4'b0001 : 4'b0000;
														assign node20114 = (inp[1]) ? 4'b0000 : 4'b0100;
										assign node20118 = (inp[7]) ? node20176 : node20119;
											assign node20119 = (inp[1]) ? node20145 : node20120;
												assign node20120 = (inp[11]) ? node20134 : node20121;
													assign node20121 = (inp[14]) ? node20127 : node20122;
														assign node20122 = (inp[12]) ? node20124 : 4'b1001;
															assign node20124 = (inp[13]) ? 4'b1001 : 4'b0001;
														assign node20127 = (inp[13]) ? node20131 : node20128;
															assign node20128 = (inp[10]) ? 4'b1000 : 4'b0000;
															assign node20131 = (inp[12]) ? 4'b1000 : 4'b0000;
													assign node20134 = (inp[13]) ? node20140 : node20135;
														assign node20135 = (inp[12]) ? 4'b0001 : node20136;
															assign node20136 = (inp[10]) ? 4'b1001 : 4'b0001;
														assign node20140 = (inp[10]) ? node20142 : 4'b1001;
															assign node20142 = (inp[12]) ? 4'b1001 : 4'b0001;
												assign node20145 = (inp[11]) ? node20165 : node20146;
													assign node20146 = (inp[14]) ? node20156 : node20147;
														assign node20147 = (inp[10]) ? 4'b0000 : node20148;
															assign node20148 = (inp[12]) ? node20152 : node20149;
																assign node20149 = (inp[13]) ? 4'b0000 : 4'b1000;
																assign node20152 = (inp[13]) ? 4'b1000 : 4'b0000;
														assign node20156 = (inp[13]) ? node20162 : node20157;
															assign node20157 = (inp[10]) ? node20159 : 4'b0001;
																assign node20159 = (inp[12]) ? 4'b0001 : 4'b1001;
															assign node20162 = (inp[12]) ? 4'b1001 : 4'b0001;
													assign node20165 = (inp[13]) ? node20171 : node20166;
														assign node20166 = (inp[12]) ? node20168 : 4'b1000;
															assign node20168 = (inp[10]) ? 4'b1000 : 4'b0000;
														assign node20171 = (inp[12]) ? node20173 : 4'b0000;
															assign node20173 = (inp[10]) ? 4'b0000 : 4'b1000;
											assign node20176 = (inp[13]) ? node20178 : 4'b0100;
												assign node20178 = (inp[12]) ? node20196 : node20179;
													assign node20179 = (inp[10]) ? node20187 : node20180;
														assign node20180 = (inp[1]) ? node20182 : 4'b0100;
															assign node20182 = (inp[11]) ? 4'b0000 : node20183;
																assign node20183 = (inp[14]) ? 4'b0100 : 4'b0000;
														assign node20187 = (inp[1]) ? node20191 : node20188;
															assign node20188 = (inp[11]) ? 4'b0001 : 4'b0000;
															assign node20191 = (inp[14]) ? node20193 : 4'b0000;
																assign node20193 = (inp[11]) ? 4'b0000 : 4'b0001;
													assign node20196 = (inp[10]) ? node20198 : 4'b0100;
														assign node20198 = (inp[1]) ? node20200 : 4'b0100;
															assign node20200 = (inp[11]) ? 4'b0000 : 4'b0100;
									assign node20203 = (inp[1]) ? node20301 : node20204;
										assign node20204 = (inp[11]) ? node20264 : node20205;
											assign node20205 = (inp[14]) ? node20235 : node20206;
												assign node20206 = (inp[4]) ? node20218 : node20207;
													assign node20207 = (inp[13]) ? node20213 : node20208;
														assign node20208 = (inp[10]) ? node20210 : 4'b0001;
															assign node20210 = (inp[12]) ? 4'b0001 : 4'b1001;
														assign node20213 = (inp[12]) ? 4'b1001 : node20214;
															assign node20214 = (inp[10]) ? 4'b0001 : 4'b1001;
													assign node20218 = (inp[7]) ? node20224 : node20219;
														assign node20219 = (inp[13]) ? 4'b1101 : node20220;
															assign node20220 = (inp[12]) ? 4'b0101 : 4'b1101;
														assign node20224 = (inp[13]) ? node20230 : node20225;
															assign node20225 = (inp[10]) ? node20227 : 4'b0001;
																assign node20227 = (inp[12]) ? 4'b0001 : 4'b1001;
															assign node20230 = (inp[12]) ? 4'b1001 : node20231;
																assign node20231 = (inp[10]) ? 4'b0101 : 4'b1001;
												assign node20235 = (inp[13]) ? node20249 : node20236;
													assign node20236 = (inp[10]) ? node20242 : node20237;
														assign node20237 = (inp[4]) ? node20239 : 4'b0000;
															assign node20239 = (inp[7]) ? 4'b0000 : 4'b0100;
														assign node20242 = (inp[12]) ? 4'b0000 : node20243;
															assign node20243 = (inp[7]) ? 4'b1000 : node20244;
																assign node20244 = (inp[4]) ? 4'b1100 : 4'b1000;
													assign node20249 = (inp[12]) ? node20259 : node20250;
														assign node20250 = (inp[10]) ? node20254 : node20251;
															assign node20251 = (inp[7]) ? 4'b1000 : 4'b1100;
															assign node20254 = (inp[4]) ? 4'b0100 : node20255;
																assign node20255 = (inp[7]) ? 4'b0000 : 4'b0100;
														assign node20259 = (inp[7]) ? 4'b1000 : node20260;
															assign node20260 = (inp[4]) ? 4'b1100 : 4'b1000;
											assign node20264 = (inp[4]) ? node20278 : node20265;
												assign node20265 = (inp[13]) ? node20271 : node20266;
													assign node20266 = (inp[10]) ? node20268 : 4'b0001;
														assign node20268 = (inp[12]) ? 4'b0001 : 4'b1001;
													assign node20271 = (inp[10]) ? node20273 : 4'b1001;
														assign node20273 = (inp[12]) ? 4'b1001 : node20274;
															assign node20274 = (inp[7]) ? 4'b0001 : 4'b0101;
												assign node20278 = (inp[7]) ? node20290 : node20279;
													assign node20279 = (inp[13]) ? node20285 : node20280;
														assign node20280 = (inp[10]) ? node20282 : 4'b0101;
															assign node20282 = (inp[12]) ? 4'b0101 : 4'b1101;
														assign node20285 = (inp[10]) ? node20287 : 4'b1101;
															assign node20287 = (inp[12]) ? 4'b1101 : 4'b0101;
													assign node20290 = (inp[13]) ? node20296 : node20291;
														assign node20291 = (inp[10]) ? node20293 : 4'b0001;
															assign node20293 = (inp[12]) ? 4'b0001 : 4'b1001;
														assign node20296 = (inp[12]) ? 4'b1001 : node20297;
															assign node20297 = (inp[10]) ? 4'b0101 : 4'b1001;
										assign node20301 = (inp[14]) ? node20337 : node20302;
											assign node20302 = (inp[13]) ? node20318 : node20303;
												assign node20303 = (inp[12]) ? node20309 : node20304;
													assign node20304 = (inp[7]) ? 4'b1000 : node20305;
														assign node20305 = (inp[4]) ? 4'b1100 : 4'b1000;
													assign node20309 = (inp[10]) ? node20315 : node20310;
														assign node20310 = (inp[4]) ? node20312 : 4'b0000;
															assign node20312 = (inp[7]) ? 4'b0000 : 4'b0100;
														assign node20315 = (inp[4]) ? 4'b1100 : 4'b1000;
												assign node20318 = (inp[7]) ? node20326 : node20319;
													assign node20319 = (inp[12]) ? node20321 : 4'b0100;
														assign node20321 = (inp[10]) ? 4'b0100 : node20322;
															assign node20322 = (inp[4]) ? 4'b1100 : 4'b1000;
													assign node20326 = (inp[4]) ? node20332 : node20327;
														assign node20327 = (inp[12]) ? node20329 : 4'b0000;
															assign node20329 = (inp[10]) ? 4'b0000 : 4'b1000;
														assign node20332 = (inp[10]) ? 4'b0100 : node20333;
															assign node20333 = (inp[12]) ? 4'b1000 : 4'b0100;
											assign node20337 = (inp[11]) ? node20369 : node20338;
												assign node20338 = (inp[4]) ? node20350 : node20339;
													assign node20339 = (inp[13]) ? node20345 : node20340;
														assign node20340 = (inp[10]) ? node20342 : 4'b0001;
															assign node20342 = (inp[12]) ? 4'b0001 : 4'b1001;
														assign node20345 = (inp[12]) ? 4'b1001 : node20346;
															assign node20346 = (inp[10]) ? 4'b0101 : 4'b1001;
													assign node20350 = (inp[7]) ? node20360 : node20351;
														assign node20351 = (inp[13]) ? node20357 : node20352;
															assign node20352 = (inp[12]) ? 4'b0101 : node20353;
																assign node20353 = (inp[10]) ? 4'b1101 : 4'b0101;
															assign node20357 = (inp[12]) ? 4'b1101 : 4'b0101;
														assign node20360 = (inp[13]) ? node20366 : node20361;
															assign node20361 = (inp[12]) ? 4'b0001 : node20362;
																assign node20362 = (inp[10]) ? 4'b1001 : 4'b0001;
															assign node20366 = (inp[12]) ? 4'b1001 : 4'b0101;
												assign node20369 = (inp[13]) ? node20381 : node20370;
													assign node20370 = (inp[10]) ? node20376 : node20371;
														assign node20371 = (inp[12]) ? 4'b0000 : node20372;
															assign node20372 = (inp[4]) ? 4'b1100 : 4'b1000;
														assign node20376 = (inp[4]) ? node20378 : 4'b1000;
															assign node20378 = (inp[7]) ? 4'b1000 : 4'b1100;
													assign node20381 = (inp[7]) ? node20383 : 4'b0100;
														assign node20383 = (inp[4]) ? node20389 : node20384;
															assign node20384 = (inp[12]) ? node20386 : 4'b0000;
																assign node20386 = (inp[10]) ? 4'b0000 : 4'b1000;
															assign node20389 = (inp[12]) ? node20391 : 4'b0100;
																assign node20391 = (inp[10]) ? 4'b0100 : 4'b1000;
						assign node20395 = (inp[3]) ? node21105 : node20396;
							assign node20396 = (inp[4]) ? node20716 : node20397;
								assign node20397 = (inp[0]) ? node20591 : node20398;
									assign node20398 = (inp[13]) ? node20486 : node20399;
										assign node20399 = (inp[10]) ? node20435 : node20400;
											assign node20400 = (inp[11]) ? node20420 : node20401;
												assign node20401 = (inp[2]) ? node20415 : node20402;
													assign node20402 = (inp[1]) ? node20408 : node20403;
														assign node20403 = (inp[14]) ? 4'b0101 : node20404;
															assign node20404 = (inp[12]) ? 4'b0100 : 4'b1100;
														assign node20408 = (inp[14]) ? 4'b1100 : node20409;
															assign node20409 = (inp[7]) ? 4'b1101 : node20410;
																assign node20410 = (inp[12]) ? 4'b1101 : 4'b0000;
													assign node20415 = (inp[1]) ? node20417 : 4'b0101;
														assign node20417 = (inp[12]) ? 4'b0101 : 4'b1101;
												assign node20420 = (inp[2]) ? node20430 : node20421;
													assign node20421 = (inp[1]) ? node20425 : node20422;
														assign node20422 = (inp[12]) ? 4'b0101 : 4'b1101;
														assign node20425 = (inp[7]) ? node20427 : 4'b0000;
															assign node20427 = (inp[12]) ? 4'b1100 : 4'b0100;
													assign node20430 = (inp[12]) ? node20432 : 4'b1100;
														assign node20432 = (inp[1]) ? 4'b1100 : 4'b0100;
											assign node20435 = (inp[7]) ? node20467 : node20436;
												assign node20436 = (inp[2]) ? node20448 : node20437;
													assign node20437 = (inp[1]) ? node20443 : node20438;
														assign node20438 = (inp[12]) ? node20440 : 4'b1000;
															assign node20440 = (inp[11]) ? 4'b1000 : 4'b0000;
														assign node20443 = (inp[12]) ? node20445 : 4'b0000;
															assign node20445 = (inp[11]) ? 4'b0000 : 4'b1000;
													assign node20448 = (inp[1]) ? node20458 : node20449;
														assign node20449 = (inp[14]) ? node20453 : node20450;
															assign node20450 = (inp[11]) ? 4'b0001 : 4'b0000;
															assign node20453 = (inp[12]) ? node20455 : 4'b0001;
																assign node20455 = (inp[11]) ? 4'b0001 : 4'b1101;
														assign node20458 = (inp[12]) ? node20464 : node20459;
															assign node20459 = (inp[11]) ? 4'b1000 : node20460;
																assign node20460 = (inp[14]) ? 4'b1000 : 4'b1001;
															assign node20464 = (inp[14]) ? 4'b0000 : 4'b1000;
												assign node20467 = (inp[2]) ? node20479 : node20468;
													assign node20468 = (inp[1]) ? node20474 : node20469;
														assign node20469 = (inp[14]) ? 4'b0101 : node20470;
															assign node20470 = (inp[11]) ? 4'b0101 : 4'b0100;
														assign node20474 = (inp[11]) ? 4'b0000 : node20475;
															assign node20475 = (inp[12]) ? 4'b0101 : 4'b0000;
													assign node20479 = (inp[11]) ? node20481 : 4'b1101;
														assign node20481 = (inp[12]) ? node20483 : 4'b0100;
															assign node20483 = (inp[1]) ? 4'b0100 : 4'b1100;
										assign node20486 = (inp[2]) ? node20534 : node20487;
											assign node20487 = (inp[1]) ? node20505 : node20488;
												assign node20488 = (inp[12]) ? node20494 : node20489;
													assign node20489 = (inp[7]) ? 4'b1000 : node20490;
														assign node20490 = (inp[10]) ? 4'b1100 : 4'b1000;
													assign node20494 = (inp[11]) ? node20500 : node20495;
														assign node20495 = (inp[7]) ? 4'b0000 : node20496;
															assign node20496 = (inp[10]) ? 4'b0100 : 4'b0000;
														assign node20500 = (inp[10]) ? node20502 : 4'b1000;
															assign node20502 = (inp[7]) ? 4'b1000 : 4'b1100;
												assign node20505 = (inp[12]) ? node20521 : node20506;
													assign node20506 = (inp[14]) ? 4'b0100 : node20507;
														assign node20507 = (inp[11]) ? node20515 : node20508;
															assign node20508 = (inp[7]) ? node20512 : node20509;
																assign node20509 = (inp[10]) ? 4'b0000 : 4'b0100;
																assign node20512 = (inp[10]) ? 4'b0100 : 4'b0000;
															assign node20515 = (inp[7]) ? node20517 : 4'b0100;
																assign node20517 = (inp[10]) ? 4'b0100 : 4'b0000;
													assign node20521 = (inp[11]) ? node20527 : node20522;
														assign node20522 = (inp[10]) ? node20524 : 4'b1000;
															assign node20524 = (inp[7]) ? 4'b1000 : 4'b1100;
														assign node20527 = (inp[10]) ? node20531 : node20528;
															assign node20528 = (inp[7]) ? 4'b0000 : 4'b0100;
															assign node20531 = (inp[7]) ? 4'b0100 : 4'b0000;
											assign node20534 = (inp[1]) ? node20564 : node20535;
												assign node20535 = (inp[10]) ? node20557 : node20536;
													assign node20536 = (inp[7]) ? node20548 : node20537;
														assign node20537 = (inp[12]) ? node20543 : node20538;
															assign node20538 = (inp[14]) ? node20540 : 4'b0000;
																assign node20540 = (inp[11]) ? 4'b0001 : 4'b1001;
															assign node20543 = (inp[11]) ? 4'b1001 : node20544;
																assign node20544 = (inp[14]) ? 4'b1001 : 4'b1000;
														assign node20548 = (inp[12]) ? node20554 : node20549;
															assign node20549 = (inp[11]) ? 4'b0001 : node20550;
																assign node20550 = (inp[14]) ? 4'b0101 : 4'b0000;
															assign node20554 = (inp[11]) ? 4'b0100 : 4'b0101;
													assign node20557 = (inp[11]) ? 4'b1001 : node20558;
														assign node20558 = (inp[14]) ? node20560 : 4'b1000;
															assign node20560 = (inp[7]) ? 4'b0001 : 4'b1001;
												assign node20564 = (inp[14]) ? node20580 : node20565;
													assign node20565 = (inp[11]) ? node20573 : node20566;
														assign node20566 = (inp[10]) ? node20568 : 4'b0001;
															assign node20568 = (inp[12]) ? 4'b1001 : node20569;
																assign node20569 = (inp[7]) ? 4'b0001 : 4'b0101;
														assign node20573 = (inp[10]) ? node20577 : node20574;
															assign node20574 = (inp[12]) ? 4'b0000 : 4'b1000;
															assign node20577 = (inp[7]) ? 4'b0000 : 4'b0100;
													assign node20580 = (inp[10]) ? node20586 : node20581;
														assign node20581 = (inp[11]) ? node20583 : 4'b0000;
															assign node20583 = (inp[12]) ? 4'b0000 : 4'b1000;
														assign node20586 = (inp[12]) ? 4'b1000 : node20587;
															assign node20587 = (inp[7]) ? 4'b0000 : 4'b0100;
									assign node20591 = (inp[2]) ? node20699 : node20592;
										assign node20592 = (inp[13]) ? node20642 : node20593;
											assign node20593 = (inp[1]) ? node20617 : node20594;
												assign node20594 = (inp[14]) ? node20604 : node20595;
													assign node20595 = (inp[10]) ? node20597 : 4'b0101;
														assign node20597 = (inp[12]) ? 4'b0101 : node20598;
															assign node20598 = (inp[11]) ? node20600 : 4'b1101;
																assign node20600 = (inp[7]) ? 4'b1101 : 4'b0000;
													assign node20604 = (inp[11]) ? node20610 : node20605;
														assign node20605 = (inp[12]) ? 4'b0100 : node20606;
															assign node20606 = (inp[10]) ? 4'b1100 : 4'b0100;
														assign node20610 = (inp[10]) ? node20612 : 4'b0101;
															assign node20612 = (inp[7]) ? node20614 : 4'b0000;
																assign node20614 = (inp[12]) ? 4'b0101 : 4'b1101;
												assign node20617 = (inp[11]) ? node20631 : node20618;
													assign node20618 = (inp[14]) ? node20626 : node20619;
														assign node20619 = (inp[12]) ? node20623 : node20620;
															assign node20620 = (inp[10]) ? 4'b0001 : 4'b1100;
															assign node20623 = (inp[10]) ? 4'b1100 : 4'b0100;
														assign node20626 = (inp[12]) ? 4'b0101 : node20627;
															assign node20627 = (inp[10]) ? 4'b0001 : 4'b0101;
													assign node20631 = (inp[7]) ? node20637 : node20632;
														assign node20632 = (inp[10]) ? 4'b0000 : node20633;
															assign node20633 = (inp[12]) ? 4'b0100 : 4'b1100;
														assign node20637 = (inp[10]) ? 4'b1100 : node20638;
															assign node20638 = (inp[12]) ? 4'b0100 : 4'b1100;
											assign node20642 = (inp[11]) ? node20682 : node20643;
												assign node20643 = (inp[7]) ? node20663 : node20644;
													assign node20644 = (inp[14]) ? node20656 : node20645;
														assign node20645 = (inp[10]) ? node20651 : node20646;
															assign node20646 = (inp[1]) ? node20648 : 4'b0001;
																assign node20648 = (inp[12]) ? 4'b0001 : 4'b1001;
															assign node20651 = (inp[1]) ? node20653 : 4'b1001;
																assign node20653 = (inp[12]) ? 4'b1001 : 4'b0001;
														assign node20656 = (inp[12]) ? 4'b1001 : node20657;
															assign node20657 = (inp[10]) ? node20659 : 4'b1001;
																assign node20659 = (inp[1]) ? 4'b0001 : 4'b1001;
													assign node20663 = (inp[12]) ? node20673 : node20664;
														assign node20664 = (inp[10]) ? node20668 : node20665;
															assign node20665 = (inp[14]) ? 4'b1101 : 4'b0100;
															assign node20668 = (inp[1]) ? 4'b0001 : node20669;
																assign node20669 = (inp[14]) ? 4'b0100 : 4'b0101;
														assign node20673 = (inp[1]) ? node20677 : node20674;
															assign node20674 = (inp[14]) ? 4'b1100 : 4'b1101;
															assign node20677 = (inp[14]) ? 4'b1101 : node20678;
																assign node20678 = (inp[10]) ? 4'b0100 : 4'b1100;
												assign node20682 = (inp[10]) ? node20694 : node20683;
													assign node20683 = (inp[7]) ? node20689 : node20684;
														assign node20684 = (inp[1]) ? 4'b1000 : node20685;
															assign node20685 = (inp[12]) ? 4'b0000 : 4'b1000;
														assign node20689 = (inp[1]) ? node20691 : 4'b1101;
															assign node20691 = (inp[12]) ? 4'b1100 : 4'b0100;
													assign node20694 = (inp[12]) ? node20696 : 4'b0000;
														assign node20696 = (inp[1]) ? 4'b0000 : 4'b1000;
										assign node20699 = (inp[7]) ? 4'b0100 : node20700;
											assign node20700 = (inp[13]) ? node20702 : 4'b0100;
												assign node20702 = (inp[12]) ? node20710 : node20703;
													assign node20703 = (inp[10]) ? node20707 : node20704;
														assign node20704 = (inp[1]) ? 4'b0000 : 4'b0100;
														assign node20707 = (inp[1]) ? 4'b0000 : 4'b0001;
													assign node20710 = (inp[1]) ? node20712 : 4'b0100;
														assign node20712 = (inp[10]) ? 4'b0000 : 4'b0100;
								assign node20716 = (inp[2]) ? node20910 : node20717;
									assign node20717 = (inp[11]) ? node20831 : node20718;
										assign node20718 = (inp[10]) ? node20772 : node20719;
											assign node20719 = (inp[0]) ? node20755 : node20720;
												assign node20720 = (inp[13]) ? node20742 : node20721;
													assign node20721 = (inp[7]) ? node20731 : node20722;
														assign node20722 = (inp[14]) ? node20726 : node20723;
															assign node20723 = (inp[1]) ? 4'b0000 : 4'b0001;
															assign node20726 = (inp[1]) ? node20728 : 4'b0000;
																assign node20728 = (inp[12]) ? 4'b1001 : 4'b0001;
														assign node20731 = (inp[1]) ? node20735 : node20732;
															assign node20732 = (inp[12]) ? 4'b0100 : 4'b1100;
															assign node20735 = (inp[12]) ? node20739 : node20736;
																assign node20736 = (inp[14]) ? 4'b0001 : 4'b0000;
																assign node20739 = (inp[14]) ? 4'b1100 : 4'b0000;
													assign node20742 = (inp[1]) ? 4'b0001 : node20743;
														assign node20743 = (inp[7]) ? node20747 : node20744;
															assign node20744 = (inp[12]) ? 4'b0001 : 4'b1001;
															assign node20747 = (inp[12]) ? node20751 : node20748;
																assign node20748 = (inp[14]) ? 4'b0100 : 4'b0101;
																assign node20751 = (inp[14]) ? 4'b1000 : 4'b1001;
												assign node20755 = (inp[12]) ? node20763 : node20756;
													assign node20756 = (inp[1]) ? node20758 : 4'b0001;
														assign node20758 = (inp[13]) ? node20760 : 4'b1001;
															assign node20760 = (inp[14]) ? 4'b0000 : 4'b0001;
													assign node20763 = (inp[7]) ? 4'b0001 : node20764;
														assign node20764 = (inp[1]) ? node20768 : node20765;
															assign node20765 = (inp[13]) ? 4'b0101 : 4'b0001;
															assign node20768 = (inp[14]) ? 4'b0000 : 4'b0001;
											assign node20772 = (inp[7]) ? node20804 : node20773;
												assign node20773 = (inp[1]) ? node20789 : node20774;
													assign node20774 = (inp[0]) ? node20784 : node20775;
														assign node20775 = (inp[12]) ? node20779 : node20776;
															assign node20776 = (inp[14]) ? 4'b1000 : 4'b0000;
															assign node20779 = (inp[13]) ? 4'b1001 : node20780;
																assign node20780 = (inp[14]) ? 4'b1000 : 4'b1001;
														assign node20784 = (inp[13]) ? node20786 : 4'b1001;
															assign node20786 = (inp[14]) ? 4'b1001 : 4'b1000;
													assign node20789 = (inp[13]) ? node20797 : node20790;
														assign node20790 = (inp[0]) ? 4'b1001 : node20791;
															assign node20791 = (inp[14]) ? 4'b0101 : node20792;
																assign node20792 = (inp[12]) ? 4'b0100 : 4'b1100;
														assign node20797 = (inp[14]) ? node20799 : 4'b1001;
															assign node20799 = (inp[0]) ? node20801 : 4'b1000;
																assign node20801 = (inp[12]) ? 4'b1000 : 4'b0000;
												assign node20804 = (inp[12]) ? node20820 : node20805;
													assign node20805 = (inp[1]) ? node20815 : node20806;
														assign node20806 = (inp[13]) ? node20812 : node20807;
															assign node20807 = (inp[14]) ? node20809 : 4'b1001;
																assign node20809 = (inp[0]) ? 4'b1001 : 4'b1000;
															assign node20812 = (inp[0]) ? 4'b1001 : 4'b0001;
														assign node20815 = (inp[0]) ? 4'b0001 : node20816;
															assign node20816 = (inp[13]) ? 4'b1001 : 4'b0001;
													assign node20820 = (inp[13]) ? 4'b1001 : node20821;
														assign node20821 = (inp[1]) ? node20827 : node20822;
															assign node20822 = (inp[14]) ? node20824 : 4'b1001;
																assign node20824 = (inp[0]) ? 4'b1001 : 4'b1000;
															assign node20827 = (inp[0]) ? 4'b1001 : 4'b0001;
										assign node20831 = (inp[10]) ? node20867 : node20832;
											assign node20832 = (inp[1]) ? node20854 : node20833;
												assign node20833 = (inp[13]) ? node20841 : node20834;
													assign node20834 = (inp[0]) ? node20838 : node20835;
														assign node20835 = (inp[7]) ? 4'b1100 : 4'b1001;
														assign node20838 = (inp[12]) ? 4'b0000 : 4'b1000;
													assign node20841 = (inp[12]) ? node20847 : node20842;
														assign node20842 = (inp[0]) ? node20844 : 4'b0000;
															assign node20844 = (inp[14]) ? 4'b0001 : 4'b1000;
														assign node20847 = (inp[0]) ? node20851 : node20848;
															assign node20848 = (inp[7]) ? 4'b0101 : 4'b1000;
															assign node20851 = (inp[7]) ? 4'b0000 : 4'b0100;
												assign node20854 = (inp[12]) ? node20856 : 4'b1000;
													assign node20856 = (inp[7]) ? 4'b1000 : node20857;
														assign node20857 = (inp[14]) ? node20859 : 4'b1000;
															assign node20859 = (inp[13]) ? node20863 : node20860;
																assign node20860 = (inp[0]) ? 4'b1000 : 4'b0000;
																assign node20863 = (inp[0]) ? 4'b0000 : 4'b1000;
											assign node20867 = (inp[1]) ? node20897 : node20868;
												assign node20868 = (inp[12]) ? node20884 : node20869;
													assign node20869 = (inp[0]) ? node20877 : node20870;
														assign node20870 = (inp[7]) ? node20874 : node20871;
															assign node20871 = (inp[13]) ? 4'b0001 : 4'b0101;
															assign node20874 = (inp[14]) ? 4'b0001 : 4'b1000;
														assign node20877 = (inp[13]) ? node20881 : node20878;
															assign node20878 = (inp[7]) ? 4'b0000 : 4'b0100;
															assign node20881 = (inp[14]) ? 4'b0100 : 4'b1001;
													assign node20884 = (inp[7]) ? node20892 : node20885;
														assign node20885 = (inp[13]) ? node20889 : node20886;
															assign node20886 = (inp[0]) ? 4'b1000 : 4'b1001;
															assign node20889 = (inp[0]) ? 4'b1001 : 4'b0001;
														assign node20892 = (inp[0]) ? 4'b1000 : node20893;
															assign node20893 = (inp[13]) ? 4'b0000 : 4'b1001;
												assign node20897 = (inp[0]) ? node20903 : node20898;
													assign node20898 = (inp[13]) ? 4'b0000 : node20899;
														assign node20899 = (inp[7]) ? 4'b1000 : 4'b0000;
													assign node20903 = (inp[12]) ? 4'b0000 : node20904;
														assign node20904 = (inp[7]) ? 4'b0000 : node20905;
															assign node20905 = (inp[13]) ? 4'b0000 : 4'b0100;
									assign node20910 = (inp[7]) ? node21030 : node20911;
										assign node20911 = (inp[1]) ? node20967 : node20912;
											assign node20912 = (inp[11]) ? node20944 : node20913;
												assign node20913 = (inp[14]) ? node20933 : node20914;
													assign node20914 = (inp[0]) ? node20926 : node20915;
														assign node20915 = (inp[10]) ? node20921 : node20916;
															assign node20916 = (inp[13]) ? 4'b1000 : node20917;
																assign node20917 = (inp[12]) ? 4'b0100 : 4'b1100;
															assign node20921 = (inp[13]) ? 4'b0001 : node20922;
																assign node20922 = (inp[12]) ? 4'b0000 : 4'b1000;
														assign node20926 = (inp[12]) ? node20930 : node20927;
															assign node20927 = (inp[13]) ? 4'b0001 : 4'b1001;
															assign node20930 = (inp[13]) ? 4'b1001 : 4'b0001;
													assign node20933 = (inp[10]) ? node20939 : node20934;
														assign node20934 = (inp[13]) ? 4'b1000 : node20935;
															assign node20935 = (inp[0]) ? 4'b0000 : 4'b0101;
														assign node20939 = (inp[12]) ? 4'b0000 : node20940;
															assign node20940 = (inp[13]) ? 4'b0000 : 4'b1000;
												assign node20944 = (inp[0]) ? node20956 : node20945;
													assign node20945 = (inp[10]) ? node20951 : node20946;
														assign node20946 = (inp[13]) ? 4'b1000 : node20947;
															assign node20947 = (inp[12]) ? 4'b0101 : 4'b1101;
														assign node20951 = (inp[13]) ? node20953 : 4'b1000;
															assign node20953 = (inp[12]) ? 4'b0001 : 4'b1001;
													assign node20956 = (inp[13]) ? node20962 : node20957;
														assign node20957 = (inp[12]) ? 4'b0001 : node20958;
															assign node20958 = (inp[10]) ? 4'b1001 : 4'b0001;
														assign node20962 = (inp[10]) ? node20964 : 4'b1001;
															assign node20964 = (inp[12]) ? 4'b1001 : 4'b0001;
											assign node20967 = (inp[11]) ? node21013 : node20968;
												assign node20968 = (inp[14]) ? node20990 : node20969;
													assign node20969 = (inp[13]) ? node20981 : node20970;
														assign node20970 = (inp[10]) ? node20976 : node20971;
															assign node20971 = (inp[0]) ? node20973 : 4'b0000;
																assign node20973 = (inp[12]) ? 4'b0000 : 4'b1000;
															assign node20976 = (inp[12]) ? 4'b1000 : node20977;
																assign node20977 = (inp[0]) ? 4'b1000 : 4'b0000;
														assign node20981 = (inp[12]) ? node20987 : node20982;
															assign node20982 = (inp[10]) ? 4'b0000 : node20983;
																assign node20983 = (inp[0]) ? 4'b0000 : 4'b0100;
															assign node20987 = (inp[10]) ? 4'b0000 : 4'b1000;
													assign node20990 = (inp[0]) ? node21004 : node20991;
														assign node20991 = (inp[10]) ? node20999 : node20992;
															assign node20992 = (inp[12]) ? node20996 : node20993;
																assign node20993 = (inp[13]) ? 4'b0100 : 4'b0000;
																assign node20996 = (inp[13]) ? 4'b1000 : 4'b1100;
															assign node20999 = (inp[13]) ? 4'b1001 : node21000;
																assign node21000 = (inp[12]) ? 4'b1000 : 4'b0000;
														assign node21004 = (inp[13]) ? node21010 : node21005;
															assign node21005 = (inp[12]) ? 4'b0001 : node21006;
																assign node21006 = (inp[10]) ? 4'b1001 : 4'b0001;
															assign node21010 = (inp[10]) ? 4'b0001 : 4'b1001;
												assign node21013 = (inp[0]) ? node21021 : node21014;
													assign node21014 = (inp[13]) ? node21016 : 4'b0000;
														assign node21016 = (inp[10]) ? 4'b0000 : node21017;
															assign node21017 = (inp[12]) ? 4'b0100 : 4'b0000;
													assign node21021 = (inp[13]) ? node21025 : node21022;
														assign node21022 = (inp[12]) ? 4'b0000 : 4'b1000;
														assign node21025 = (inp[12]) ? node21027 : 4'b0000;
															assign node21027 = (inp[10]) ? 4'b0000 : 4'b1000;
										assign node21030 = (inp[0]) ? node21080 : node21031;
											assign node21031 = (inp[13]) ? node21069 : node21032;
												assign node21032 = (inp[1]) ? node21056 : node21033;
													assign node21033 = (inp[10]) ? node21047 : node21034;
														assign node21034 = (inp[12]) ? node21042 : node21035;
															assign node21035 = (inp[14]) ? node21039 : node21036;
																assign node21036 = (inp[11]) ? 4'b1001 : 4'b1000;
																assign node21039 = (inp[11]) ? 4'b1001 : 4'b0001;
															assign node21042 = (inp[14]) ? 4'b0001 : node21043;
																assign node21043 = (inp[11]) ? 4'b0001 : 4'b0000;
														assign node21047 = (inp[14]) ? node21051 : node21048;
															assign node21048 = (inp[11]) ? 4'b0101 : 4'b0100;
															assign node21051 = (inp[12]) ? node21053 : 4'b0101;
																assign node21053 = (inp[11]) ? 4'b0101 : 4'b1001;
													assign node21056 = (inp[10]) ? node21062 : node21057;
														assign node21057 = (inp[11]) ? node21059 : 4'b1000;
															assign node21059 = (inp[12]) ? 4'b1000 : 4'b0100;
														assign node21062 = (inp[12]) ? node21064 : 4'b0000;
															assign node21064 = (inp[11]) ? 4'b0000 : node21065;
																assign node21065 = (inp[14]) ? 4'b0100 : 4'b0101;
												assign node21069 = (inp[1]) ? node21075 : node21070;
													assign node21070 = (inp[12]) ? node21072 : 4'b1000;
														assign node21072 = (inp[11]) ? 4'b1000 : 4'b0000;
													assign node21075 = (inp[11]) ? 4'b0000 : node21076;
														assign node21076 = (inp[12]) ? 4'b1000 : 4'b0000;
											assign node21080 = (inp[13]) ? node21082 : 4'b0100;
												assign node21082 = (inp[10]) ? node21090 : node21083;
													assign node21083 = (inp[1]) ? node21085 : 4'b0100;
														assign node21085 = (inp[12]) ? 4'b0100 : node21086;
															assign node21086 = (inp[11]) ? 4'b0000 : 4'b0100;
													assign node21090 = (inp[12]) ? node21098 : node21091;
														assign node21091 = (inp[1]) ? node21093 : 4'b0001;
															assign node21093 = (inp[14]) ? node21095 : 4'b0000;
																assign node21095 = (inp[11]) ? 4'b0000 : 4'b0001;
														assign node21098 = (inp[1]) ? node21100 : 4'b0100;
															assign node21100 = (inp[14]) ? node21102 : 4'b0000;
																assign node21102 = (inp[11]) ? 4'b0000 : 4'b0100;
							assign node21105 = (inp[4]) ? node21511 : node21106;
								assign node21106 = (inp[11]) ? node21356 : node21107;
									assign node21107 = (inp[2]) ? node21211 : node21108;
										assign node21108 = (inp[13]) ? node21154 : node21109;
											assign node21109 = (inp[10]) ? node21131 : node21110;
												assign node21110 = (inp[14]) ? node21116 : node21111;
													assign node21111 = (inp[1]) ? node21113 : 4'b1000;
														assign node21113 = (inp[7]) ? 4'b1001 : 4'b1000;
													assign node21116 = (inp[1]) ? node21122 : node21117;
														assign node21117 = (inp[12]) ? 4'b0001 : node21118;
															assign node21118 = (inp[0]) ? 4'b0001 : 4'b1001;
														assign node21122 = (inp[0]) ? node21126 : node21123;
															assign node21123 = (inp[7]) ? 4'b0000 : 4'b1000;
															assign node21126 = (inp[7]) ? 4'b1000 : node21127;
																assign node21127 = (inp[12]) ? 4'b1000 : 4'b0000;
												assign node21131 = (inp[1]) ? node21143 : node21132;
													assign node21132 = (inp[0]) ? node21134 : 4'b1000;
														assign node21134 = (inp[7]) ? node21138 : node21135;
															assign node21135 = (inp[12]) ? 4'b0000 : 4'b1000;
															assign node21138 = (inp[14]) ? node21140 : 4'b0000;
																assign node21140 = (inp[12]) ? 4'b1001 : 4'b0001;
													assign node21143 = (inp[12]) ? node21149 : node21144;
														assign node21144 = (inp[14]) ? node21146 : 4'b0000;
															assign node21146 = (inp[0]) ? 4'b0000 : 4'b0001;
														assign node21149 = (inp[7]) ? 4'b0001 : node21150;
															assign node21150 = (inp[0]) ? 4'b1000 : 4'b0000;
											assign node21154 = (inp[1]) ? node21182 : node21155;
												assign node21155 = (inp[0]) ? node21171 : node21156;
													assign node21156 = (inp[7]) ? node21162 : node21157;
														assign node21157 = (inp[10]) ? node21159 : 4'b1001;
															assign node21159 = (inp[12]) ? 4'b1000 : 4'b0000;
														assign node21162 = (inp[10]) ? node21166 : node21163;
															assign node21163 = (inp[14]) ? 4'b0000 : 4'b0001;
															assign node21166 = (inp[14]) ? node21168 : 4'b0000;
																assign node21168 = (inp[12]) ? 4'b1001 : 4'b0000;
													assign node21171 = (inp[14]) ? 4'b0000 : node21172;
														assign node21172 = (inp[10]) ? 4'b0001 : node21173;
															assign node21173 = (inp[7]) ? node21177 : node21174;
																assign node21174 = (inp[12]) ? 4'b0000 : 4'b0001;
																assign node21177 = (inp[12]) ? 4'b0000 : 4'b1000;
												assign node21182 = (inp[0]) ? node21196 : node21183;
													assign node21183 = (inp[10]) ? node21191 : node21184;
														assign node21184 = (inp[12]) ? node21188 : node21185;
															assign node21185 = (inp[7]) ? 4'b0001 : 4'b1001;
															assign node21188 = (inp[7]) ? 4'b1001 : 4'b1000;
														assign node21191 = (inp[14]) ? 4'b0001 : node21192;
															assign node21192 = (inp[7]) ? 4'b1000 : 4'b0001;
													assign node21196 = (inp[14]) ? node21206 : node21197;
														assign node21197 = (inp[12]) ? node21201 : node21198;
															assign node21198 = (inp[10]) ? 4'b0000 : 4'b1000;
															assign node21201 = (inp[7]) ? 4'b1000 : node21202;
																assign node21202 = (inp[10]) ? 4'b1001 : 4'b1000;
														assign node21206 = (inp[10]) ? 4'b1001 : node21207;
															assign node21207 = (inp[7]) ? 4'b1000 : 4'b1001;
										assign node21211 = (inp[7]) ? node21275 : node21212;
											assign node21212 = (inp[12]) ? node21246 : node21213;
												assign node21213 = (inp[14]) ? node21229 : node21214;
													assign node21214 = (inp[10]) ? node21222 : node21215;
														assign node21215 = (inp[1]) ? 4'b1000 : node21216;
															assign node21216 = (inp[13]) ? 4'b0000 : node21217;
																assign node21217 = (inp[0]) ? 4'b0001 : 4'b1001;
														assign node21222 = (inp[1]) ? node21224 : 4'b1001;
															assign node21224 = (inp[13]) ? node21226 : 4'b0001;
																assign node21226 = (inp[0]) ? 4'b0001 : 4'b1001;
													assign node21229 = (inp[13]) ? node21239 : node21230;
														assign node21230 = (inp[0]) ? node21236 : node21231;
															assign node21231 = (inp[1]) ? node21233 : 4'b0001;
																assign node21233 = (inp[10]) ? 4'b0000 : 4'b0001;
															assign node21236 = (inp[1]) ? 4'b0001 : 4'b0000;
														assign node21239 = (inp[10]) ? node21243 : node21240;
															assign node21240 = (inp[1]) ? 4'b1000 : 4'b0001;
															assign node21243 = (inp[1]) ? 4'b0000 : 4'b1000;
												assign node21246 = (inp[10]) ? node21256 : node21247;
													assign node21247 = (inp[0]) ? 4'b0001 : node21248;
														assign node21248 = (inp[13]) ? node21250 : 4'b0001;
															assign node21250 = (inp[14]) ? 4'b1001 : node21251;
																assign node21251 = (inp[1]) ? 4'b1000 : 4'b0000;
													assign node21256 = (inp[1]) ? node21270 : node21257;
														assign node21257 = (inp[14]) ? node21263 : node21258;
															assign node21258 = (inp[13]) ? 4'b0001 : node21259;
																assign node21259 = (inp[0]) ? 4'b0001 : 4'b1001;
															assign node21263 = (inp[13]) ? node21267 : node21264;
																assign node21264 = (inp[0]) ? 4'b0000 : 4'b1001;
																assign node21267 = (inp[0]) ? 4'b1001 : 4'b0000;
														assign node21270 = (inp[0]) ? node21272 : 4'b0001;
															assign node21272 = (inp[13]) ? 4'b1001 : 4'b0001;
											assign node21275 = (inp[10]) ? node21319 : node21276;
												assign node21276 = (inp[0]) ? node21300 : node21277;
													assign node21277 = (inp[12]) ? node21291 : node21278;
														assign node21278 = (inp[1]) ? node21284 : node21279;
															assign node21279 = (inp[13]) ? 4'b0000 : node21280;
																assign node21280 = (inp[14]) ? 4'b1000 : 4'b1001;
															assign node21284 = (inp[14]) ? node21288 : node21285;
																assign node21285 = (inp[13]) ? 4'b0001 : 4'b0000;
																assign node21288 = (inp[13]) ? 4'b0000 : 4'b0001;
														assign node21291 = (inp[1]) ? node21297 : node21292;
															assign node21292 = (inp[13]) ? node21294 : 4'b0000;
																assign node21294 = (inp[14]) ? 4'b0001 : 4'b0000;
															assign node21297 = (inp[14]) ? 4'b1000 : 4'b0000;
													assign node21300 = (inp[13]) ? node21308 : node21301;
														assign node21301 = (inp[1]) ? node21305 : node21302;
															assign node21302 = (inp[14]) ? 4'b0000 : 4'b0001;
															assign node21305 = (inp[14]) ? 4'b0001 : 4'b1000;
														assign node21308 = (inp[12]) ? node21314 : node21309;
															assign node21309 = (inp[14]) ? node21311 : 4'b0000;
																assign node21311 = (inp[1]) ? 4'b1001 : 4'b1000;
															assign node21314 = (inp[14]) ? node21316 : 4'b1001;
																assign node21316 = (inp[1]) ? 4'b1001 : 4'b1000;
												assign node21319 = (inp[0]) ? node21333 : node21320;
													assign node21320 = (inp[13]) ? node21326 : node21321;
														assign node21321 = (inp[12]) ? 4'b1001 : node21322;
															assign node21322 = (inp[1]) ? 4'b1001 : 4'b0001;
														assign node21326 = (inp[1]) ? node21328 : 4'b1000;
															assign node21328 = (inp[14]) ? node21330 : 4'b1000;
																assign node21330 = (inp[12]) ? 4'b0001 : 4'b1001;
													assign node21333 = (inp[13]) ? node21345 : node21334;
														assign node21334 = (inp[12]) ? node21340 : node21335;
															assign node21335 = (inp[1]) ? node21337 : 4'b1000;
																assign node21337 = (inp[14]) ? 4'b1001 : 4'b1000;
															assign node21340 = (inp[14]) ? node21342 : 4'b1000;
																assign node21342 = (inp[1]) ? 4'b0001 : 4'b0000;
														assign node21345 = (inp[12]) ? node21351 : node21346;
															assign node21346 = (inp[1]) ? 4'b0001 : node21347;
																assign node21347 = (inp[14]) ? 4'b0000 : 4'b0001;
															assign node21351 = (inp[1]) ? 4'b0000 : node21352;
																assign node21352 = (inp[14]) ? 4'b1000 : 4'b1001;
									assign node21356 = (inp[1]) ? node21450 : node21357;
										assign node21357 = (inp[7]) ? node21401 : node21358;
											assign node21358 = (inp[10]) ? node21378 : node21359;
												assign node21359 = (inp[0]) ? node21367 : node21360;
													assign node21360 = (inp[2]) ? 4'b0000 : node21361;
														assign node21361 = (inp[12]) ? 4'b0000 : node21362;
															assign node21362 = (inp[13]) ? 4'b0001 : 4'b0000;
													assign node21367 = (inp[13]) ? node21373 : node21368;
														assign node21368 = (inp[2]) ? 4'b0001 : node21369;
															assign node21369 = (inp[12]) ? 4'b0001 : 4'b1001;
														assign node21373 = (inp[2]) ? node21375 : 4'b0001;
															assign node21375 = (inp[12]) ? 4'b0000 : 4'b1000;
												assign node21378 = (inp[0]) ? node21390 : node21379;
													assign node21379 = (inp[2]) ? node21383 : node21380;
														assign node21380 = (inp[12]) ? 4'b0001 : 4'b1001;
														assign node21383 = (inp[13]) ? node21387 : node21384;
															assign node21384 = (inp[12]) ? 4'b0000 : 4'b1000;
															assign node21387 = (inp[12]) ? 4'b1001 : 4'b0000;
													assign node21390 = (inp[2]) ? node21396 : node21391;
														assign node21391 = (inp[13]) ? node21393 : 4'b1000;
															assign node21393 = (inp[12]) ? 4'b0000 : 4'b1000;
														assign node21396 = (inp[12]) ? node21398 : 4'b0000;
															assign node21398 = (inp[13]) ? 4'b1000 : 4'b0001;
											assign node21401 = (inp[13]) ? node21425 : node21402;
												assign node21402 = (inp[10]) ? node21414 : node21403;
													assign node21403 = (inp[0]) ? node21409 : node21404;
														assign node21404 = (inp[2]) ? 4'b1001 : node21405;
															assign node21405 = (inp[12]) ? 4'b1001 : 4'b0001;
														assign node21409 = (inp[2]) ? 4'b0001 : node21410;
															assign node21410 = (inp[12]) ? 4'b0001 : 4'b1001;
													assign node21414 = (inp[0]) ? node21420 : node21415;
														assign node21415 = (inp[2]) ? node21417 : 4'b0000;
															assign node21417 = (inp[12]) ? 4'b0000 : 4'b1000;
														assign node21420 = (inp[2]) ? node21422 : 4'b0001;
															assign node21422 = (inp[12]) ? 4'b0001 : 4'b1001;
												assign node21425 = (inp[2]) ? node21437 : node21426;
													assign node21426 = (inp[0]) ? node21432 : node21427;
														assign node21427 = (inp[10]) ? 4'b1000 : node21428;
															assign node21428 = (inp[12]) ? 4'b0000 : 4'b1000;
														assign node21432 = (inp[10]) ? node21434 : 4'b1000;
															assign node21434 = (inp[12]) ? 4'b0001 : 4'b1001;
													assign node21437 = (inp[10]) ? node21443 : node21438;
														assign node21438 = (inp[0]) ? 4'b1001 : node21439;
															assign node21439 = (inp[12]) ? 4'b0001 : 4'b1001;
														assign node21443 = (inp[0]) ? node21447 : node21444;
															assign node21444 = (inp[12]) ? 4'b0000 : 4'b0001;
															assign node21447 = (inp[12]) ? 4'b1001 : 4'b0000;
										assign node21450 = (inp[2]) ? node21476 : node21451;
											assign node21451 = (inp[7]) ? node21461 : node21452;
												assign node21452 = (inp[10]) ? 4'b0000 : node21453;
													assign node21453 = (inp[0]) ? node21455 : 4'b0000;
														assign node21455 = (inp[12]) ? node21457 : 4'b0000;
															assign node21457 = (inp[13]) ? 4'b1000 : 4'b0000;
												assign node21461 = (inp[13]) ? node21469 : node21462;
													assign node21462 = (inp[0]) ? node21466 : node21463;
														assign node21463 = (inp[10]) ? 4'b1000 : 4'b0000;
														assign node21466 = (inp[10]) ? 4'b0000 : 4'b1000;
													assign node21469 = (inp[10]) ? 4'b0000 : node21470;
														assign node21470 = (inp[12]) ? 4'b0000 : node21471;
															assign node21471 = (inp[0]) ? 4'b0000 : 4'b1000;
											assign node21476 = (inp[13]) ? node21502 : node21477;
												assign node21477 = (inp[12]) ? node21493 : node21478;
													assign node21478 = (inp[10]) ? node21480 : 4'b1000;
														assign node21480 = (inp[14]) ? node21488 : node21481;
															assign node21481 = (inp[7]) ? node21485 : node21482;
																assign node21482 = (inp[0]) ? 4'b0000 : 4'b1000;
																assign node21485 = (inp[0]) ? 4'b1000 : 4'b0000;
															assign node21488 = (inp[0]) ? node21490 : 4'b1000;
																assign node21490 = (inp[7]) ? 4'b1000 : 4'b0000;
													assign node21493 = (inp[0]) ? node21497 : node21494;
														assign node21494 = (inp[7]) ? 4'b0000 : 4'b1000;
														assign node21497 = (inp[10]) ? node21499 : 4'b0000;
															assign node21499 = (inp[7]) ? 4'b1000 : 4'b0000;
												assign node21502 = (inp[0]) ? node21504 : 4'b0000;
													assign node21504 = (inp[10]) ? 4'b0000 : node21505;
														assign node21505 = (inp[12]) ? 4'b1000 : node21506;
															assign node21506 = (inp[7]) ? 4'b0000 : 4'b1000;
								assign node21511 = (inp[13]) ? node21709 : node21512;
									assign node21512 = (inp[11]) ? node21642 : node21513;
										assign node21513 = (inp[10]) ? node21575 : node21514;
											assign node21514 = (inp[7]) ? node21544 : node21515;
												assign node21515 = (inp[1]) ? node21529 : node21516;
													assign node21516 = (inp[14]) ? node21526 : node21517;
														assign node21517 = (inp[0]) ? node21521 : node21518;
															assign node21518 = (inp[2]) ? 4'b1000 : 4'b0000;
															assign node21521 = (inp[12]) ? node21523 : 4'b1000;
																assign node21523 = (inp[2]) ? 4'b0000 : 4'b1000;
														assign node21526 = (inp[0]) ? 4'b0001 : 4'b0000;
													assign node21529 = (inp[0]) ? node21535 : node21530;
														assign node21530 = (inp[12]) ? node21532 : 4'b1001;
															assign node21532 = (inp[2]) ? 4'b1000 : 4'b0001;
														assign node21535 = (inp[2]) ? node21541 : node21536;
															assign node21536 = (inp[14]) ? 4'b1000 : node21537;
																assign node21537 = (inp[12]) ? 4'b1000 : 4'b0000;
															assign node21541 = (inp[14]) ? 4'b1000 : 4'b1001;
												assign node21544 = (inp[0]) ? node21560 : node21545;
													assign node21545 = (inp[14]) ? node21551 : node21546;
														assign node21546 = (inp[2]) ? node21548 : 4'b0000;
															assign node21548 = (inp[12]) ? 4'b1001 : 4'b0000;
														assign node21551 = (inp[1]) ? node21557 : node21552;
															assign node21552 = (inp[12]) ? 4'b1001 : node21553;
																assign node21553 = (inp[2]) ? 4'b1001 : 4'b0001;
															assign node21557 = (inp[12]) ? 4'b0000 : 4'b1000;
													assign node21560 = (inp[12]) ? node21568 : node21561;
														assign node21561 = (inp[2]) ? node21565 : node21562;
															assign node21562 = (inp[14]) ? 4'b1000 : 4'b1001;
															assign node21565 = (inp[1]) ? 4'b1001 : 4'b0001;
														assign node21568 = (inp[14]) ? node21570 : 4'b0001;
															assign node21570 = (inp[1]) ? node21572 : 4'b0001;
																assign node21572 = (inp[2]) ? 4'b0001 : 4'b0000;
											assign node21575 = (inp[1]) ? node21607 : node21576;
												assign node21576 = (inp[7]) ? node21588 : node21577;
													assign node21577 = (inp[2]) ? node21583 : node21578;
														assign node21578 = (inp[14]) ? node21580 : 4'b0001;
															assign node21580 = (inp[12]) ? 4'b1000 : 4'b0001;
														assign node21583 = (inp[0]) ? node21585 : 4'b0000;
															assign node21585 = (inp[12]) ? 4'b0000 : 4'b1000;
													assign node21588 = (inp[2]) ? node21598 : node21589;
														assign node21589 = (inp[12]) ? node21595 : node21590;
															assign node21590 = (inp[0]) ? node21592 : 4'b1000;
																assign node21592 = (inp[14]) ? 4'b0000 : 4'b0001;
															assign node21595 = (inp[0]) ? 4'b1000 : 4'b0000;
														assign node21598 = (inp[14]) ? node21602 : node21599;
															assign node21599 = (inp[0]) ? 4'b0000 : 4'b0001;
															assign node21602 = (inp[0]) ? node21604 : 4'b1001;
																assign node21604 = (inp[12]) ? 4'b1001 : 4'b0001;
												assign node21607 = (inp[12]) ? node21625 : node21608;
													assign node21608 = (inp[7]) ? node21620 : node21609;
														assign node21609 = (inp[0]) ? node21615 : node21610;
															assign node21610 = (inp[2]) ? 4'b0000 : node21611;
																assign node21611 = (inp[14]) ? 4'b0000 : 4'b0001;
															assign node21615 = (inp[14]) ? 4'b1000 : node21616;
																assign node21616 = (inp[2]) ? 4'b1000 : 4'b0000;
														assign node21620 = (inp[2]) ? node21622 : 4'b0001;
															assign node21622 = (inp[0]) ? 4'b0000 : 4'b0001;
													assign node21625 = (inp[7]) ? node21637 : node21626;
														assign node21626 = (inp[0]) ? node21632 : node21627;
															assign node21627 = (inp[14]) ? node21629 : 4'b0001;
																assign node21629 = (inp[2]) ? 4'b0000 : 4'b0001;
															assign node21632 = (inp[2]) ? node21634 : 4'b0000;
																assign node21634 = (inp[14]) ? 4'b0001 : 4'b0000;
														assign node21637 = (inp[0]) ? 4'b0001 : node21638;
															assign node21638 = (inp[14]) ? 4'b0001 : 4'b1000;
										assign node21642 = (inp[1]) ? node21682 : node21643;
											assign node21643 = (inp[0]) ? node21663 : node21644;
												assign node21644 = (inp[10]) ? node21654 : node21645;
													assign node21645 = (inp[2]) ? node21649 : node21646;
														assign node21646 = (inp[7]) ? 4'b0000 : 4'b0001;
														assign node21649 = (inp[7]) ? node21651 : 4'b1000;
															assign node21651 = (inp[12]) ? 4'b0001 : 4'b1001;
													assign node21654 = (inp[7]) ? node21660 : node21655;
														assign node21655 = (inp[2]) ? node21657 : 4'b0000;
															assign node21657 = (inp[12]) ? 4'b0001 : 4'b0000;
														assign node21660 = (inp[12]) ? 4'b0000 : 4'b1000;
												assign node21663 = (inp[10]) ? node21673 : node21664;
													assign node21664 = (inp[7]) ? node21670 : node21665;
														assign node21665 = (inp[2]) ? node21667 : 4'b0000;
															assign node21667 = (inp[12]) ? 4'b0001 : 4'b1001;
														assign node21670 = (inp[14]) ? 4'b0000 : 4'b1000;
													assign node21673 = (inp[14]) ? 4'b0001 : node21674;
														assign node21674 = (inp[12]) ? node21678 : node21675;
															assign node21675 = (inp[2]) ? 4'b0001 : 4'b0000;
															assign node21678 = (inp[2]) ? 4'b1000 : 4'b0001;
											assign node21682 = (inp[10]) ? 4'b0000 : node21683;
												assign node21683 = (inp[2]) ? node21697 : node21684;
													assign node21684 = (inp[14]) ? 4'b0000 : node21685;
														assign node21685 = (inp[7]) ? node21691 : node21686;
															assign node21686 = (inp[12]) ? 4'b0000 : node21687;
																assign node21687 = (inp[0]) ? 4'b1000 : 4'b0000;
															assign node21691 = (inp[12]) ? node21693 : 4'b0000;
																assign node21693 = (inp[0]) ? 4'b0000 : 4'b1000;
													assign node21697 = (inp[12]) ? node21703 : node21698;
														assign node21698 = (inp[7]) ? node21700 : 4'b0000;
															assign node21700 = (inp[0]) ? 4'b0000 : 4'b1000;
														assign node21703 = (inp[7]) ? node21705 : 4'b1000;
															assign node21705 = (inp[0]) ? 4'b1000 : 4'b0000;
									assign node21709 = (inp[11]) ? node21819 : node21710;
										assign node21710 = (inp[10]) ? node21780 : node21711;
											assign node21711 = (inp[12]) ? node21743 : node21712;
												assign node21712 = (inp[0]) ? node21728 : node21713;
													assign node21713 = (inp[14]) ? node21721 : node21714;
														assign node21714 = (inp[7]) ? 4'b0000 : node21715;
															assign node21715 = (inp[1]) ? 4'b0000 : node21716;
																assign node21716 = (inp[2]) ? 4'b0001 : 4'b0000;
														assign node21721 = (inp[2]) ? 4'b0000 : node21722;
															assign node21722 = (inp[7]) ? node21724 : 4'b0000;
																assign node21724 = (inp[1]) ? 4'b0001 : 4'b0000;
													assign node21728 = (inp[2]) ? node21736 : node21729;
														assign node21729 = (inp[14]) ? 4'b0000 : node21730;
															assign node21730 = (inp[7]) ? node21732 : 4'b0000;
																assign node21732 = (inp[1]) ? 4'b0000 : 4'b0001;
														assign node21736 = (inp[7]) ? node21740 : node21737;
															assign node21737 = (inp[14]) ? 4'b0001 : 4'b0000;
															assign node21740 = (inp[14]) ? 4'b0000 : 4'b0001;
												assign node21743 = (inp[7]) ? node21761 : node21744;
													assign node21744 = (inp[0]) ? node21750 : node21745;
														assign node21745 = (inp[14]) ? node21747 : 4'b0001;
															assign node21747 = (inp[1]) ? 4'b0000 : 4'b0001;
														assign node21750 = (inp[14]) ? node21756 : node21751;
															assign node21751 = (inp[2]) ? 4'b0000 : node21752;
																assign node21752 = (inp[1]) ? 4'b0001 : 4'b0000;
															assign node21756 = (inp[1]) ? 4'b0001 : node21757;
																assign node21757 = (inp[2]) ? 4'b0001 : 4'b0000;
													assign node21761 = (inp[0]) ? node21769 : node21762;
														assign node21762 = (inp[2]) ? node21764 : 4'b0000;
															assign node21764 = (inp[14]) ? node21766 : 4'b0000;
																assign node21766 = (inp[1]) ? 4'b0000 : 4'b0001;
														assign node21769 = (inp[1]) ? node21775 : node21770;
															assign node21770 = (inp[14]) ? 4'b0000 : node21771;
																assign node21771 = (inp[2]) ? 4'b0000 : 4'b0001;
															assign node21775 = (inp[2]) ? 4'b0001 : node21776;
																assign node21776 = (inp[14]) ? 4'b0000 : 4'b0001;
											assign node21780 = (inp[1]) ? 4'b0000 : node21781;
												assign node21781 = (inp[12]) ? node21799 : node21782;
													assign node21782 = (inp[2]) ? node21794 : node21783;
														assign node21783 = (inp[7]) ? node21789 : node21784;
															assign node21784 = (inp[0]) ? node21786 : 4'b0001;
																assign node21786 = (inp[14]) ? 4'b0001 : 4'b0000;
															assign node21789 = (inp[0]) ? node21791 : 4'b0000;
																assign node21791 = (inp[14]) ? 4'b0000 : 4'b0001;
														assign node21794 = (inp[7]) ? node21796 : 4'b0000;
															assign node21796 = (inp[14]) ? 4'b0001 : 4'b0000;
													assign node21799 = (inp[2]) ? node21805 : node21800;
														assign node21800 = (inp[14]) ? 4'b0000 : node21801;
															assign node21801 = (inp[7]) ? 4'b0000 : 4'b0001;
														assign node21805 = (inp[14]) ? node21811 : node21806;
															assign node21806 = (inp[7]) ? node21808 : 4'b0000;
																assign node21808 = (inp[0]) ? 4'b0000 : 4'b0001;
															assign node21811 = (inp[0]) ? node21815 : node21812;
																assign node21812 = (inp[7]) ? 4'b0000 : 4'b0001;
																assign node21815 = (inp[7]) ? 4'b0001 : 4'b0000;
										assign node21819 = (inp[1]) ? 4'b0000 : node21820;
											assign node21820 = (inp[10]) ? 4'b0000 : node21821;
												assign node21821 = (inp[0]) ? node21843 : node21822;
													assign node21822 = (inp[12]) ? node21828 : node21823;
														assign node21823 = (inp[2]) ? node21825 : 4'b0000;
															assign node21825 = (inp[7]) ? 4'b0001 : 4'b0000;
														assign node21828 = (inp[14]) ? node21836 : node21829;
															assign node21829 = (inp[2]) ? node21833 : node21830;
																assign node21830 = (inp[7]) ? 4'b0001 : 4'b0000;
																assign node21833 = (inp[7]) ? 4'b0000 : 4'b0001;
															assign node21836 = (inp[2]) ? node21840 : node21837;
																assign node21837 = (inp[7]) ? 4'b0001 : 4'b0000;
																assign node21840 = (inp[7]) ? 4'b0000 : 4'b0001;
													assign node21843 = (inp[14]) ? node21845 : 4'b0000;
														assign node21845 = (inp[7]) ? node21851 : node21846;
															assign node21846 = (inp[2]) ? 4'b0000 : node21847;
																assign node21847 = (inp[12]) ? 4'b0000 : 4'b0001;
															assign node21851 = (inp[2]) ? node21853 : 4'b0000;
																assign node21853 = (inp[12]) ? 4'b0001 : 4'b0000;
				assign node21858 = (inp[0]) ? node23842 : node21859;
					assign node21859 = (inp[6]) ? node22421 : node21860;
						assign node21860 = (inp[5]) ? node21982 : node21861;
							assign node21861 = (inp[3]) ? node21863 : 4'b0010;
								assign node21863 = (inp[2]) ? 4'b0010 : node21864;
									assign node21864 = (inp[4]) ? node21892 : node21865;
										assign node21865 = (inp[7]) ? 4'b0010 : node21866;
											assign node21866 = (inp[13]) ? node21868 : 4'b0010;
												assign node21868 = (inp[12]) ? node21882 : node21869;
													assign node21869 = (inp[10]) ? node21873 : node21870;
														assign node21870 = (inp[1]) ? 4'b0000 : 4'b0010;
														assign node21873 = (inp[1]) ? node21879 : node21874;
															assign node21874 = (inp[14]) ? node21876 : 4'b0001;
																assign node21876 = (inp[11]) ? 4'b0001 : 4'b0000;
															assign node21879 = (inp[14]) ? 4'b0001 : 4'b0000;
													assign node21882 = (inp[10]) ? node21884 : 4'b0010;
														assign node21884 = (inp[1]) ? node21886 : 4'b0010;
															assign node21886 = (inp[14]) ? node21888 : 4'b0000;
																assign node21888 = (inp[11]) ? 4'b0000 : 4'b0010;
										assign node21892 = (inp[7]) ? node21954 : node21893;
											assign node21893 = (inp[1]) ? node21923 : node21894;
												assign node21894 = (inp[14]) ? node21906 : node21895;
													assign node21895 = (inp[13]) ? node21901 : node21896;
														assign node21896 = (inp[12]) ? 4'b0001 : node21897;
															assign node21897 = (inp[10]) ? 4'b1001 : 4'b0001;
														assign node21901 = (inp[10]) ? node21903 : 4'b1001;
															assign node21903 = (inp[12]) ? 4'b1001 : 4'b0001;
													assign node21906 = (inp[11]) ? node21918 : node21907;
														assign node21907 = (inp[13]) ? node21913 : node21908;
															assign node21908 = (inp[10]) ? node21910 : 4'b0000;
																assign node21910 = (inp[12]) ? 4'b0000 : 4'b1000;
															assign node21913 = (inp[10]) ? node21915 : 4'b1000;
																assign node21915 = (inp[12]) ? 4'b1000 : 4'b0000;
														assign node21918 = (inp[13]) ? node21920 : 4'b0001;
															assign node21920 = (inp[12]) ? 4'b1001 : 4'b0001;
												assign node21923 = (inp[14]) ? node21935 : node21924;
													assign node21924 = (inp[13]) ? node21930 : node21925;
														assign node21925 = (inp[12]) ? node21927 : 4'b1000;
															assign node21927 = (inp[10]) ? 4'b1000 : 4'b0000;
														assign node21930 = (inp[10]) ? 4'b0000 : node21931;
															assign node21931 = (inp[12]) ? 4'b1000 : 4'b0000;
													assign node21935 = (inp[11]) ? node21947 : node21936;
														assign node21936 = (inp[13]) ? node21942 : node21937;
															assign node21937 = (inp[10]) ? node21939 : 4'b0001;
																assign node21939 = (inp[12]) ? 4'b0001 : 4'b1001;
															assign node21942 = (inp[10]) ? node21944 : 4'b1001;
																assign node21944 = (inp[12]) ? 4'b1001 : 4'b0001;
														assign node21947 = (inp[13]) ? 4'b0000 : node21948;
															assign node21948 = (inp[12]) ? node21950 : 4'b1000;
																assign node21950 = (inp[10]) ? 4'b1000 : 4'b0000;
											assign node21954 = (inp[13]) ? node21956 : 4'b0010;
												assign node21956 = (inp[10]) ? node21964 : node21957;
													assign node21957 = (inp[11]) ? node21959 : 4'b0010;
														assign node21959 = (inp[12]) ? 4'b0010 : node21960;
															assign node21960 = (inp[1]) ? 4'b0000 : 4'b0010;
													assign node21964 = (inp[12]) ? node21974 : node21965;
														assign node21965 = (inp[1]) ? node21971 : node21966;
															assign node21966 = (inp[14]) ? node21968 : 4'b0001;
																assign node21968 = (inp[11]) ? 4'b0001 : 4'b0000;
															assign node21971 = (inp[14]) ? 4'b0001 : 4'b0000;
														assign node21974 = (inp[1]) ? node21976 : 4'b0010;
															assign node21976 = (inp[11]) ? 4'b0000 : node21977;
																assign node21977 = (inp[14]) ? 4'b0010 : 4'b0000;
							assign node21982 = (inp[2]) ? node22316 : node21983;
								assign node21983 = (inp[1]) ? node22153 : node21984;
									assign node21984 = (inp[13]) ? node22068 : node21985;
										assign node21985 = (inp[3]) ? node22029 : node21986;
											assign node21986 = (inp[12]) ? node22012 : node21987;
												assign node21987 = (inp[10]) ? node21997 : node21988;
													assign node21988 = (inp[11]) ? node21992 : node21989;
														assign node21989 = (inp[14]) ? 4'b0000 : 4'b0001;
														assign node21992 = (inp[4]) ? node21994 : 4'b0001;
															assign node21994 = (inp[7]) ? 4'b0001 : 4'b0101;
													assign node21997 = (inp[7]) ? node22007 : node21998;
														assign node21998 = (inp[4]) ? node22002 : node21999;
															assign node21999 = (inp[11]) ? 4'b1001 : 4'b1000;
															assign node22002 = (inp[14]) ? node22004 : 4'b1101;
																assign node22004 = (inp[11]) ? 4'b1101 : 4'b1100;
														assign node22007 = (inp[14]) ? node22009 : 4'b1001;
															assign node22009 = (inp[11]) ? 4'b1001 : 4'b1000;
												assign node22012 = (inp[11]) ? node22024 : node22013;
													assign node22013 = (inp[14]) ? node22019 : node22014;
														assign node22014 = (inp[4]) ? node22016 : 4'b0001;
															assign node22016 = (inp[7]) ? 4'b0001 : 4'b0101;
														assign node22019 = (inp[4]) ? node22021 : 4'b0000;
															assign node22021 = (inp[7]) ? 4'b0000 : 4'b0100;
													assign node22024 = (inp[4]) ? node22026 : 4'b0001;
														assign node22026 = (inp[7]) ? 4'b0001 : 4'b0101;
											assign node22029 = (inp[10]) ? node22047 : node22030;
												assign node22030 = (inp[11]) ? node22042 : node22031;
													assign node22031 = (inp[14]) ? node22037 : node22032;
														assign node22032 = (inp[4]) ? node22034 : 4'b0101;
															assign node22034 = (inp[7]) ? 4'b0101 : 4'b0001;
														assign node22037 = (inp[4]) ? node22039 : 4'b0100;
															assign node22039 = (inp[7]) ? 4'b0100 : 4'b0000;
													assign node22042 = (inp[4]) ? node22044 : 4'b0101;
														assign node22044 = (inp[7]) ? 4'b0101 : 4'b0001;
												assign node22047 = (inp[12]) ? node22059 : node22048;
													assign node22048 = (inp[4]) ? node22050 : 4'b1101;
														assign node22050 = (inp[7]) ? node22054 : node22051;
															assign node22051 = (inp[11]) ? 4'b1001 : 4'b1000;
															assign node22054 = (inp[14]) ? node22056 : 4'b1101;
																assign node22056 = (inp[11]) ? 4'b1101 : 4'b1100;
													assign node22059 = (inp[7]) ? node22063 : node22060;
														assign node22060 = (inp[14]) ? 4'b0000 : 4'b0001;
														assign node22063 = (inp[14]) ? node22065 : 4'b0101;
															assign node22065 = (inp[11]) ? 4'b0101 : 4'b0100;
										assign node22068 = (inp[14]) ? node22106 : node22069;
											assign node22069 = (inp[12]) ? node22095 : node22070;
												assign node22070 = (inp[10]) ? node22088 : node22071;
													assign node22071 = (inp[11]) ? node22079 : node22072;
														assign node22072 = (inp[7]) ? 4'b1001 : node22073;
															assign node22073 = (inp[3]) ? 4'b1001 : node22074;
																assign node22074 = (inp[4]) ? 4'b1101 : 4'b1001;
														assign node22079 = (inp[4]) ? node22083 : node22080;
															assign node22080 = (inp[3]) ? 4'b1101 : 4'b1001;
															assign node22083 = (inp[3]) ? 4'b1001 : node22084;
																assign node22084 = (inp[7]) ? 4'b1001 : 4'b1101;
													assign node22088 = (inp[3]) ? 4'b0001 : node22089;
														assign node22089 = (inp[7]) ? node22091 : 4'b0101;
															assign node22091 = (inp[4]) ? 4'b0101 : 4'b0001;
												assign node22095 = (inp[3]) ? node22101 : node22096;
													assign node22096 = (inp[4]) ? node22098 : 4'b1001;
														assign node22098 = (inp[7]) ? 4'b1001 : 4'b1101;
													assign node22101 = (inp[7]) ? 4'b1101 : node22102;
														assign node22102 = (inp[4]) ? 4'b1001 : 4'b1101;
											assign node22106 = (inp[11]) ? node22130 : node22107;
												assign node22107 = (inp[10]) ? node22119 : node22108;
													assign node22108 = (inp[3]) ? node22114 : node22109;
														assign node22109 = (inp[4]) ? node22111 : 4'b1000;
															assign node22111 = (inp[7]) ? 4'b1000 : 4'b1100;
														assign node22114 = (inp[4]) ? node22116 : 4'b1100;
															assign node22116 = (inp[7]) ? 4'b1100 : 4'b1000;
													assign node22119 = (inp[12]) ? node22123 : node22120;
														assign node22120 = (inp[3]) ? 4'b0000 : 4'b0100;
														assign node22123 = (inp[3]) ? 4'b1100 : node22124;
															assign node22124 = (inp[4]) ? node22126 : 4'b1000;
																assign node22126 = (inp[7]) ? 4'b1000 : 4'b1100;
												assign node22130 = (inp[12]) ? node22142 : node22131;
													assign node22131 = (inp[10]) ? node22139 : node22132;
														assign node22132 = (inp[7]) ? 4'b1001 : node22133;
															assign node22133 = (inp[3]) ? 4'b1101 : node22134;
																assign node22134 = (inp[4]) ? 4'b1101 : 4'b1001;
														assign node22139 = (inp[3]) ? 4'b0001 : 4'b0101;
													assign node22142 = (inp[3]) ? node22148 : node22143;
														assign node22143 = (inp[4]) ? node22145 : 4'b1001;
															assign node22145 = (inp[7]) ? 4'b1001 : 4'b1101;
														assign node22148 = (inp[4]) ? node22150 : 4'b1101;
															assign node22150 = (inp[7]) ? 4'b1101 : 4'b1001;
									assign node22153 = (inp[14]) ? node22217 : node22154;
										assign node22154 = (inp[13]) ? node22188 : node22155;
											assign node22155 = (inp[3]) ? node22173 : node22156;
												assign node22156 = (inp[10]) ? node22168 : node22157;
													assign node22157 = (inp[12]) ? node22163 : node22158;
														assign node22158 = (inp[7]) ? 4'b1000 : node22159;
															assign node22159 = (inp[4]) ? 4'b1100 : 4'b1000;
														assign node22163 = (inp[7]) ? 4'b0000 : node22164;
															assign node22164 = (inp[4]) ? 4'b0100 : 4'b0000;
													assign node22168 = (inp[4]) ? node22170 : 4'b1000;
														assign node22170 = (inp[7]) ? 4'b1000 : 4'b1100;
												assign node22173 = (inp[7]) ? node22183 : node22174;
													assign node22174 = (inp[4]) ? 4'b1000 : node22175;
														assign node22175 = (inp[11]) ? node22177 : 4'b1100;
															assign node22177 = (inp[12]) ? node22179 : 4'b1100;
																assign node22179 = (inp[10]) ? 4'b1100 : 4'b0100;
													assign node22183 = (inp[10]) ? 4'b1100 : node22184;
														assign node22184 = (inp[12]) ? 4'b0100 : 4'b1100;
											assign node22188 = (inp[10]) ? node22206 : node22189;
												assign node22189 = (inp[12]) ? node22201 : node22190;
													assign node22190 = (inp[3]) ? node22196 : node22191;
														assign node22191 = (inp[7]) ? node22193 : 4'b0100;
															assign node22193 = (inp[4]) ? 4'b0100 : 4'b0000;
														assign node22196 = (inp[7]) ? node22198 : 4'b0000;
															assign node22198 = (inp[11]) ? 4'b0100 : 4'b0000;
													assign node22201 = (inp[3]) ? 4'b1100 : node22202;
														assign node22202 = (inp[7]) ? 4'b1000 : 4'b1100;
												assign node22206 = (inp[3]) ? node22212 : node22207;
													assign node22207 = (inp[7]) ? node22209 : 4'b0100;
														assign node22209 = (inp[4]) ? 4'b0100 : 4'b0000;
													assign node22212 = (inp[7]) ? node22214 : 4'b0000;
														assign node22214 = (inp[4]) ? 4'b0000 : 4'b0100;
										assign node22217 = (inp[11]) ? node22273 : node22218;
											assign node22218 = (inp[13]) ? node22244 : node22219;
												assign node22219 = (inp[3]) ? node22229 : node22220;
													assign node22220 = (inp[10]) ? node22226 : node22221;
														assign node22221 = (inp[4]) ? node22223 : 4'b0001;
															assign node22223 = (inp[7]) ? 4'b0001 : 4'b0101;
														assign node22226 = (inp[12]) ? 4'b0001 : 4'b1001;
													assign node22229 = (inp[7]) ? node22239 : node22230;
														assign node22230 = (inp[4]) ? node22234 : node22231;
															assign node22231 = (inp[12]) ? 4'b0101 : 4'b1101;
															assign node22234 = (inp[10]) ? node22236 : 4'b0001;
																assign node22236 = (inp[12]) ? 4'b0001 : 4'b1001;
														assign node22239 = (inp[12]) ? 4'b0101 : node22240;
															assign node22240 = (inp[10]) ? 4'b1101 : 4'b0101;
												assign node22244 = (inp[12]) ? node22262 : node22245;
													assign node22245 = (inp[10]) ? node22255 : node22246;
														assign node22246 = (inp[3]) ? node22250 : node22247;
															assign node22247 = (inp[4]) ? 4'b1101 : 4'b1001;
															assign node22250 = (inp[4]) ? node22252 : 4'b1101;
																assign node22252 = (inp[7]) ? 4'b1101 : 4'b1001;
														assign node22255 = (inp[3]) ? node22257 : 4'b0101;
															assign node22257 = (inp[7]) ? node22259 : 4'b0001;
																assign node22259 = (inp[4]) ? 4'b0001 : 4'b0101;
													assign node22262 = (inp[3]) ? node22268 : node22263;
														assign node22263 = (inp[7]) ? 4'b1001 : node22264;
															assign node22264 = (inp[4]) ? 4'b1101 : 4'b1001;
														assign node22268 = (inp[7]) ? 4'b1101 : node22269;
															assign node22269 = (inp[4]) ? 4'b1001 : 4'b1101;
											assign node22273 = (inp[13]) ? node22295 : node22274;
												assign node22274 = (inp[12]) ? node22284 : node22275;
													assign node22275 = (inp[3]) ? node22281 : node22276;
														assign node22276 = (inp[7]) ? 4'b1000 : node22277;
															assign node22277 = (inp[4]) ? 4'b1100 : 4'b1000;
														assign node22281 = (inp[7]) ? 4'b1100 : 4'b1000;
													assign node22284 = (inp[10]) ? node22292 : node22285;
														assign node22285 = (inp[3]) ? 4'b0100 : node22286;
															assign node22286 = (inp[4]) ? node22288 : 4'b0000;
																assign node22288 = (inp[7]) ? 4'b0000 : 4'b0100;
														assign node22292 = (inp[4]) ? 4'b1100 : 4'b1000;
												assign node22295 = (inp[3]) ? node22305 : node22296;
													assign node22296 = (inp[4]) ? 4'b0100 : node22297;
														assign node22297 = (inp[10]) ? node22301 : node22298;
															assign node22298 = (inp[12]) ? 4'b1000 : 4'b0000;
															assign node22301 = (inp[7]) ? 4'b0000 : 4'b0100;
													assign node22305 = (inp[4]) ? node22311 : node22306;
														assign node22306 = (inp[7]) ? node22308 : 4'b0000;
															assign node22308 = (inp[10]) ? 4'b0100 : 4'b1100;
														assign node22311 = (inp[12]) ? node22313 : 4'b0000;
															assign node22313 = (inp[7]) ? 4'b0000 : 4'b1000;
								assign node22316 = (inp[3]) ? node22318 : 4'b0010;
									assign node22318 = (inp[4]) ? node22338 : node22319;
										assign node22319 = (inp[7]) ? 4'b0010 : node22320;
											assign node22320 = (inp[13]) ? node22322 : 4'b0010;
												assign node22322 = (inp[12]) ? node22328 : node22323;
													assign node22323 = (inp[1]) ? 4'b0000 : node22324;
														assign node22324 = (inp[10]) ? 4'b0001 : 4'b0010;
													assign node22328 = (inp[1]) ? node22330 : 4'b0010;
														assign node22330 = (inp[10]) ? node22332 : 4'b0010;
															assign node22332 = (inp[11]) ? 4'b0000 : node22333;
																assign node22333 = (inp[14]) ? 4'b0010 : 4'b0000;
										assign node22338 = (inp[7]) ? node22402 : node22339;
											assign node22339 = (inp[1]) ? node22369 : node22340;
												assign node22340 = (inp[11]) ? node22358 : node22341;
													assign node22341 = (inp[14]) ? node22349 : node22342;
														assign node22342 = (inp[13]) ? node22346 : node22343;
															assign node22343 = (inp[12]) ? 4'b0001 : 4'b1001;
															assign node22346 = (inp[12]) ? 4'b1001 : 4'b0001;
														assign node22349 = (inp[10]) ? node22351 : 4'b0000;
															assign node22351 = (inp[12]) ? node22355 : node22352;
																assign node22352 = (inp[13]) ? 4'b0000 : 4'b1000;
																assign node22355 = (inp[13]) ? 4'b1000 : 4'b0000;
													assign node22358 = (inp[13]) ? node22364 : node22359;
														assign node22359 = (inp[10]) ? node22361 : 4'b0001;
															assign node22361 = (inp[12]) ? 4'b0001 : 4'b1001;
														assign node22364 = (inp[10]) ? node22366 : 4'b1001;
															assign node22366 = (inp[12]) ? 4'b1001 : 4'b0001;
												assign node22369 = (inp[11]) ? node22391 : node22370;
													assign node22370 = (inp[14]) ? node22380 : node22371;
														assign node22371 = (inp[13]) ? node22377 : node22372;
															assign node22372 = (inp[12]) ? node22374 : 4'b1000;
																assign node22374 = (inp[10]) ? 4'b1000 : 4'b0000;
															assign node22377 = (inp[12]) ? 4'b1000 : 4'b0000;
														assign node22380 = (inp[13]) ? node22386 : node22381;
															assign node22381 = (inp[10]) ? node22383 : 4'b0001;
																assign node22383 = (inp[12]) ? 4'b0001 : 4'b1001;
															assign node22386 = (inp[10]) ? node22388 : 4'b1001;
																assign node22388 = (inp[12]) ? 4'b1001 : 4'b0001;
													assign node22391 = (inp[13]) ? node22397 : node22392;
														assign node22392 = (inp[10]) ? 4'b1000 : node22393;
															assign node22393 = (inp[12]) ? 4'b0000 : 4'b1000;
														assign node22397 = (inp[12]) ? node22399 : 4'b0000;
															assign node22399 = (inp[10]) ? 4'b0000 : 4'b1000;
											assign node22402 = (inp[13]) ? node22404 : 4'b0010;
												assign node22404 = (inp[12]) ? node22416 : node22405;
													assign node22405 = (inp[10]) ? node22413 : node22406;
														assign node22406 = (inp[11]) ? 4'b0000 : node22407;
															assign node22407 = (inp[14]) ? 4'b0010 : node22408;
																assign node22408 = (inp[1]) ? 4'b0000 : 4'b0010;
														assign node22413 = (inp[1]) ? 4'b0000 : 4'b0001;
													assign node22416 = (inp[10]) ? node22418 : 4'b0010;
														assign node22418 = (inp[1]) ? 4'b0000 : 4'b0010;
						assign node22421 = (inp[5]) ? node23101 : node22422;
							assign node22422 = (inp[11]) ? node22834 : node22423;
								assign node22423 = (inp[3]) ? node22623 : node22424;
									assign node22424 = (inp[4]) ? node22492 : node22425;
										assign node22425 = (inp[13]) ? node22451 : node22426;
											assign node22426 = (inp[10]) ? node22436 : node22427;
												assign node22427 = (inp[1]) ? node22431 : node22428;
													assign node22428 = (inp[14]) ? 4'b0000 : 4'b0001;
													assign node22431 = (inp[14]) ? 4'b0001 : node22432;
														assign node22432 = (inp[12]) ? 4'b0000 : 4'b1000;
												assign node22436 = (inp[12]) ? node22444 : node22437;
													assign node22437 = (inp[14]) ? node22441 : node22438;
														assign node22438 = (inp[1]) ? 4'b1000 : 4'b1001;
														assign node22441 = (inp[1]) ? 4'b1001 : 4'b1000;
													assign node22444 = (inp[1]) ? node22448 : node22445;
														assign node22445 = (inp[14]) ? 4'b0000 : 4'b0001;
														assign node22448 = (inp[14]) ? 4'b0001 : 4'b1000;
											assign node22451 = (inp[12]) ? node22483 : node22452;
												assign node22452 = (inp[10]) ? node22462 : node22453;
													assign node22453 = (inp[1]) ? node22457 : node22454;
														assign node22454 = (inp[14]) ? 4'b1000 : 4'b1001;
														assign node22457 = (inp[14]) ? 4'b1001 : node22458;
															assign node22458 = (inp[7]) ? 4'b0000 : 4'b0100;
													assign node22462 = (inp[7]) ? node22476 : node22463;
														assign node22463 = (inp[2]) ? node22469 : node22464;
															assign node22464 = (inp[1]) ? 4'b0101 : node22465;
																assign node22465 = (inp[14]) ? 4'b0100 : 4'b0101;
															assign node22469 = (inp[1]) ? node22473 : node22470;
																assign node22470 = (inp[14]) ? 4'b0100 : 4'b0101;
																assign node22473 = (inp[14]) ? 4'b0101 : 4'b0100;
														assign node22476 = (inp[1]) ? node22480 : node22477;
															assign node22477 = (inp[14]) ? 4'b0000 : 4'b0001;
															assign node22480 = (inp[14]) ? 4'b0001 : 4'b0000;
												assign node22483 = (inp[1]) ? node22487 : node22484;
													assign node22484 = (inp[14]) ? 4'b1000 : 4'b1001;
													assign node22487 = (inp[14]) ? 4'b1001 : node22488;
														assign node22488 = (inp[10]) ? 4'b0000 : 4'b1000;
										assign node22492 = (inp[7]) ? node22556 : node22493;
											assign node22493 = (inp[13]) ? node22521 : node22494;
												assign node22494 = (inp[12]) ? node22512 : node22495;
													assign node22495 = (inp[10]) ? node22503 : node22496;
														assign node22496 = (inp[14]) ? node22500 : node22497;
															assign node22497 = (inp[1]) ? 4'b1100 : 4'b0101;
															assign node22500 = (inp[1]) ? 4'b0101 : 4'b0100;
														assign node22503 = (inp[2]) ? node22507 : node22504;
															assign node22504 = (inp[14]) ? 4'b1100 : 4'b0001;
															assign node22507 = (inp[14]) ? 4'b1101 : node22508;
																assign node22508 = (inp[1]) ? 4'b1100 : 4'b1101;
													assign node22512 = (inp[14]) ? node22518 : node22513;
														assign node22513 = (inp[1]) ? node22515 : 4'b0101;
															assign node22515 = (inp[10]) ? 4'b1100 : 4'b0100;
														assign node22518 = (inp[1]) ? 4'b0101 : 4'b0100;
												assign node22521 = (inp[2]) ? node22533 : node22522;
													assign node22522 = (inp[10]) ? node22528 : node22523;
														assign node22523 = (inp[1]) ? node22525 : 4'b0001;
															assign node22525 = (inp[12]) ? 4'b0001 : 4'b1001;
														assign node22528 = (inp[12]) ? 4'b1001 : node22529;
															assign node22529 = (inp[1]) ? 4'b0001 : 4'b1001;
													assign node22533 = (inp[12]) ? node22543 : node22534;
														assign node22534 = (inp[10]) ? node22540 : node22535;
															assign node22535 = (inp[1]) ? 4'b0100 : node22536;
																assign node22536 = (inp[14]) ? 4'b1100 : 4'b1101;
															assign node22540 = (inp[1]) ? 4'b0101 : 4'b0100;
														assign node22543 = (inp[10]) ? node22551 : node22544;
															assign node22544 = (inp[14]) ? node22548 : node22545;
																assign node22545 = (inp[1]) ? 4'b1100 : 4'b1101;
																assign node22548 = (inp[1]) ? 4'b1101 : 4'b1100;
															assign node22551 = (inp[1]) ? node22553 : 4'b1101;
																assign node22553 = (inp[14]) ? 4'b1101 : 4'b0100;
											assign node22556 = (inp[13]) ? node22592 : node22557;
												assign node22557 = (inp[12]) ? node22571 : node22558;
													assign node22558 = (inp[10]) ? node22566 : node22559;
														assign node22559 = (inp[1]) ? node22563 : node22560;
															assign node22560 = (inp[14]) ? 4'b0000 : 4'b0001;
															assign node22563 = (inp[14]) ? 4'b0001 : 4'b1000;
														assign node22566 = (inp[14]) ? 4'b1001 : node22567;
															assign node22567 = (inp[1]) ? 4'b1000 : 4'b1001;
													assign node22571 = (inp[2]) ? node22579 : node22572;
														assign node22572 = (inp[14]) ? node22576 : node22573;
															assign node22573 = (inp[1]) ? 4'b0000 : 4'b0001;
															assign node22576 = (inp[1]) ? 4'b0001 : 4'b0000;
														assign node22579 = (inp[10]) ? node22587 : node22580;
															assign node22580 = (inp[14]) ? node22584 : node22581;
																assign node22581 = (inp[1]) ? 4'b0000 : 4'b0001;
																assign node22584 = (inp[1]) ? 4'b0001 : 4'b0000;
															assign node22587 = (inp[14]) ? node22589 : 4'b1000;
																assign node22589 = (inp[1]) ? 4'b0001 : 4'b0000;
												assign node22592 = (inp[10]) ? node22602 : node22593;
													assign node22593 = (inp[14]) ? node22599 : node22594;
														assign node22594 = (inp[1]) ? node22596 : 4'b1001;
															assign node22596 = (inp[12]) ? 4'b1000 : 4'b0100;
														assign node22599 = (inp[1]) ? 4'b1001 : 4'b1000;
													assign node22602 = (inp[2]) ? node22614 : node22603;
														assign node22603 = (inp[12]) ? node22609 : node22604;
															assign node22604 = (inp[1]) ? 4'b0001 : node22605;
																assign node22605 = (inp[14]) ? 4'b0100 : 4'b0101;
															assign node22609 = (inp[1]) ? 4'b0100 : node22610;
																assign node22610 = (inp[14]) ? 4'b1000 : 4'b1001;
														assign node22614 = (inp[12]) ? 4'b0100 : node22615;
															assign node22615 = (inp[1]) ? node22619 : node22616;
																assign node22616 = (inp[14]) ? 4'b0100 : 4'b0101;
																assign node22619 = (inp[14]) ? 4'b0101 : 4'b0100;
									assign node22623 = (inp[2]) ? node22697 : node22624;
										assign node22624 = (inp[10]) ? node22660 : node22625;
											assign node22625 = (inp[4]) ? node22643 : node22626;
												assign node22626 = (inp[13]) ? node22632 : node22627;
													assign node22627 = (inp[12]) ? 4'b0001 : node22628;
														assign node22628 = (inp[1]) ? 4'b1001 : 4'b0001;
													assign node22632 = (inp[7]) ? node22638 : node22633;
														assign node22633 = (inp[1]) ? node22635 : 4'b0101;
															assign node22635 = (inp[12]) ? 4'b0101 : 4'b1101;
														assign node22638 = (inp[12]) ? 4'b0001 : node22639;
															assign node22639 = (inp[1]) ? 4'b1001 : 4'b0001;
												assign node22643 = (inp[7]) ? node22655 : node22644;
													assign node22644 = (inp[13]) ? node22646 : 4'b0101;
														assign node22646 = (inp[12]) ? 4'b0001 : node22647;
															assign node22647 = (inp[14]) ? node22651 : node22648;
																assign node22648 = (inp[1]) ? 4'b0001 : 4'b0000;
																assign node22651 = (inp[1]) ? 4'b0000 : 4'b0001;
													assign node22655 = (inp[12]) ? 4'b0101 : node22656;
														assign node22656 = (inp[1]) ? 4'b1101 : 4'b0101;
											assign node22660 = (inp[1]) ? node22676 : node22661;
												assign node22661 = (inp[4]) ? node22667 : node22662;
													assign node22662 = (inp[7]) ? 4'b1001 : node22663;
														assign node22663 = (inp[13]) ? 4'b1101 : 4'b1001;
													assign node22667 = (inp[13]) ? node22669 : 4'b1101;
														assign node22669 = (inp[7]) ? 4'b1101 : node22670;
															assign node22670 = (inp[14]) ? node22672 : 4'b1000;
																assign node22672 = (inp[12]) ? 4'b0001 : 4'b1001;
												assign node22676 = (inp[12]) ? node22690 : node22677;
													assign node22677 = (inp[4]) ? node22683 : node22678;
														assign node22678 = (inp[7]) ? node22680 : 4'b0101;
															assign node22680 = (inp[13]) ? 4'b0101 : 4'b0001;
														assign node22683 = (inp[13]) ? node22687 : node22684;
															assign node22684 = (inp[7]) ? 4'b0101 : 4'b0001;
															assign node22687 = (inp[14]) ? 4'b0000 : 4'b0001;
													assign node22690 = (inp[4]) ? 4'b1101 : node22691;
														assign node22691 = (inp[7]) ? 4'b1001 : node22692;
															assign node22692 = (inp[13]) ? 4'b1101 : 4'b1001;
										assign node22697 = (inp[7]) ? node22771 : node22698;
											assign node22698 = (inp[4]) ? node22744 : node22699;
												assign node22699 = (inp[13]) ? node22719 : node22700;
													assign node22700 = (inp[10]) ? node22710 : node22701;
														assign node22701 = (inp[14]) ? node22707 : node22702;
															assign node22702 = (inp[1]) ? node22704 : 4'b0101;
																assign node22704 = (inp[12]) ? 4'b0100 : 4'b1100;
															assign node22707 = (inp[1]) ? 4'b0101 : 4'b0100;
														assign node22710 = (inp[14]) ? node22714 : node22711;
															assign node22711 = (inp[1]) ? 4'b1100 : 4'b1101;
															assign node22714 = (inp[1]) ? 4'b0101 : node22715;
																assign node22715 = (inp[12]) ? 4'b0100 : 4'b1100;
													assign node22719 = (inp[12]) ? node22731 : node22720;
														assign node22720 = (inp[10]) ? node22724 : node22721;
															assign node22721 = (inp[14]) ? 4'b1100 : 4'b0000;
															assign node22724 = (inp[14]) ? node22728 : node22725;
																assign node22725 = (inp[1]) ? 4'b0000 : 4'b0001;
																assign node22728 = (inp[1]) ? 4'b0001 : 4'b0000;
														assign node22731 = (inp[10]) ? node22739 : node22732;
															assign node22732 = (inp[14]) ? node22736 : node22733;
																assign node22733 = (inp[1]) ? 4'b1100 : 4'b1101;
																assign node22736 = (inp[1]) ? 4'b1101 : 4'b1100;
															assign node22739 = (inp[14]) ? node22741 : 4'b0000;
																assign node22741 = (inp[1]) ? 4'b1101 : 4'b1100;
												assign node22744 = (inp[13]) ? node22760 : node22745;
													assign node22745 = (inp[14]) ? node22753 : node22746;
														assign node22746 = (inp[1]) ? node22750 : node22747;
															assign node22747 = (inp[10]) ? 4'b1001 : 4'b0001;
															assign node22750 = (inp[10]) ? 4'b0001 : 4'b1000;
														assign node22753 = (inp[1]) ? 4'b0001 : node22754;
															assign node22754 = (inp[10]) ? node22756 : 4'b0000;
																assign node22756 = (inp[12]) ? 4'b0000 : 4'b1000;
													assign node22760 = (inp[10]) ? node22766 : node22761;
														assign node22761 = (inp[12]) ? 4'b0001 : node22762;
															assign node22762 = (inp[1]) ? 4'b1001 : 4'b0001;
														assign node22766 = (inp[12]) ? 4'b1001 : node22767;
															assign node22767 = (inp[1]) ? 4'b0001 : 4'b1001;
											assign node22771 = (inp[13]) ? node22805 : node22772;
												assign node22772 = (inp[12]) ? node22792 : node22773;
													assign node22773 = (inp[10]) ? node22785 : node22774;
														assign node22774 = (inp[4]) ? node22780 : node22775;
															assign node22775 = (inp[14]) ? node22777 : 4'b0101;
																assign node22777 = (inp[1]) ? 4'b0101 : 4'b0100;
															assign node22780 = (inp[1]) ? 4'b1100 : node22781;
																assign node22781 = (inp[14]) ? 4'b0100 : 4'b0101;
														assign node22785 = (inp[1]) ? node22789 : node22786;
															assign node22786 = (inp[14]) ? 4'b1100 : 4'b1101;
															assign node22789 = (inp[14]) ? 4'b1101 : 4'b1100;
													assign node22792 = (inp[10]) ? node22798 : node22793;
														assign node22793 = (inp[1]) ? node22795 : 4'b0101;
															assign node22795 = (inp[14]) ? 4'b0101 : 4'b0100;
														assign node22798 = (inp[14]) ? node22802 : node22799;
															assign node22799 = (inp[1]) ? 4'b1100 : 4'b0101;
															assign node22802 = (inp[1]) ? 4'b0101 : 4'b0100;
												assign node22805 = (inp[12]) ? node22825 : node22806;
													assign node22806 = (inp[10]) ? node22816 : node22807;
														assign node22807 = (inp[14]) ? node22813 : node22808;
															assign node22808 = (inp[1]) ? node22810 : 4'b1101;
																assign node22810 = (inp[4]) ? 4'b0000 : 4'b0100;
															assign node22813 = (inp[1]) ? 4'b1101 : 4'b1100;
														assign node22816 = (inp[4]) ? node22822 : node22817;
															assign node22817 = (inp[14]) ? 4'b0101 : node22818;
																assign node22818 = (inp[1]) ? 4'b0100 : 4'b0101;
															assign node22822 = (inp[14]) ? 4'b0000 : 4'b0001;
													assign node22825 = (inp[14]) ? node22831 : node22826;
														assign node22826 = (inp[1]) ? node22828 : 4'b1101;
															assign node22828 = (inp[10]) ? 4'b0000 : 4'b1100;
														assign node22831 = (inp[1]) ? 4'b1101 : 4'b1100;
								assign node22834 = (inp[1]) ? node22974 : node22835;
									assign node22835 = (inp[3]) ? node22889 : node22836;
										assign node22836 = (inp[13]) ? node22858 : node22837;
											assign node22837 = (inp[12]) ? node22853 : node22838;
												assign node22838 = (inp[10]) ? node22844 : node22839;
													assign node22839 = (inp[7]) ? 4'b0001 : node22840;
														assign node22840 = (inp[4]) ? 4'b0101 : 4'b0001;
													assign node22844 = (inp[4]) ? node22846 : 4'b1001;
														assign node22846 = (inp[2]) ? node22850 : node22847;
															assign node22847 = (inp[7]) ? 4'b1001 : 4'b0000;
															assign node22850 = (inp[7]) ? 4'b1001 : 4'b1101;
												assign node22853 = (inp[4]) ? node22855 : 4'b0001;
													assign node22855 = (inp[7]) ? 4'b0001 : 4'b0101;
											assign node22858 = (inp[10]) ? node22870 : node22859;
												assign node22859 = (inp[7]) ? 4'b1001 : node22860;
													assign node22860 = (inp[2]) ? node22866 : node22861;
														assign node22861 = (inp[4]) ? node22863 : 4'b1001;
															assign node22863 = (inp[12]) ? 4'b0000 : 4'b1000;
														assign node22866 = (inp[4]) ? 4'b1101 : 4'b1001;
												assign node22870 = (inp[12]) ? node22882 : node22871;
													assign node22871 = (inp[2]) ? node22877 : node22872;
														assign node22872 = (inp[4]) ? 4'b0000 : node22873;
															assign node22873 = (inp[7]) ? 4'b0001 : 4'b0101;
														assign node22877 = (inp[7]) ? node22879 : 4'b0101;
															assign node22879 = (inp[4]) ? 4'b0101 : 4'b0001;
													assign node22882 = (inp[4]) ? node22884 : 4'b1001;
														assign node22884 = (inp[7]) ? 4'b1001 : node22885;
															assign node22885 = (inp[2]) ? 4'b1101 : 4'b1000;
										assign node22889 = (inp[2]) ? node22935 : node22890;
											assign node22890 = (inp[4]) ? node22912 : node22891;
												assign node22891 = (inp[7]) ? node22903 : node22892;
													assign node22892 = (inp[12]) ? node22896 : node22893;
														assign node22893 = (inp[10]) ? 4'b0100 : 4'b1100;
														assign node22896 = (inp[13]) ? node22900 : node22897;
															assign node22897 = (inp[10]) ? 4'b1000 : 4'b0000;
															assign node22900 = (inp[10]) ? 4'b1100 : 4'b0100;
													assign node22903 = (inp[10]) ? node22907 : node22904;
														assign node22904 = (inp[12]) ? 4'b0000 : 4'b1000;
														assign node22907 = (inp[12]) ? 4'b1000 : node22908;
															assign node22908 = (inp[13]) ? 4'b0100 : 4'b0000;
												assign node22912 = (inp[7]) ? node22926 : node22913;
													assign node22913 = (inp[13]) ? node22921 : node22914;
														assign node22914 = (inp[10]) ? node22918 : node22915;
															assign node22915 = (inp[12]) ? 4'b0100 : 4'b1100;
															assign node22918 = (inp[12]) ? 4'b1100 : 4'b0000;
														assign node22921 = (inp[10]) ? 4'b1001 : node22922;
															assign node22922 = (inp[12]) ? 4'b0000 : 4'b0001;
													assign node22926 = (inp[10]) ? node22930 : node22927;
														assign node22927 = (inp[12]) ? 4'b0100 : 4'b1100;
														assign node22930 = (inp[12]) ? 4'b1100 : node22931;
															assign node22931 = (inp[13]) ? 4'b0000 : 4'b0100;
											assign node22935 = (inp[4]) ? node22949 : node22936;
												assign node22936 = (inp[13]) ? node22942 : node22937;
													assign node22937 = (inp[10]) ? node22939 : 4'b0101;
														assign node22939 = (inp[12]) ? 4'b0101 : 4'b1101;
													assign node22942 = (inp[10]) ? node22944 : 4'b1101;
														assign node22944 = (inp[12]) ? 4'b1101 : node22945;
															assign node22945 = (inp[7]) ? 4'b0101 : 4'b0001;
												assign node22949 = (inp[7]) ? node22963 : node22950;
													assign node22950 = (inp[13]) ? node22956 : node22951;
														assign node22951 = (inp[12]) ? 4'b0001 : node22952;
															assign node22952 = (inp[10]) ? 4'b0000 : 4'b0001;
														assign node22956 = (inp[10]) ? node22960 : node22957;
															assign node22957 = (inp[12]) ? 4'b0000 : 4'b1000;
															assign node22960 = (inp[12]) ? 4'b1000 : 4'b0000;
													assign node22963 = (inp[13]) ? node22969 : node22964;
														assign node22964 = (inp[10]) ? node22966 : 4'b0101;
															assign node22966 = (inp[12]) ? 4'b0101 : 4'b1101;
														assign node22969 = (inp[12]) ? 4'b1101 : node22970;
															assign node22970 = (inp[10]) ? 4'b0000 : 4'b1101;
									assign node22974 = (inp[13]) ? node23032 : node22975;
										assign node22975 = (inp[3]) ? node23001 : node22976;
											assign node22976 = (inp[12]) ? node22986 : node22977;
												assign node22977 = (inp[7]) ? 4'b1000 : node22978;
													assign node22978 = (inp[4]) ? node22980 : 4'b1000;
														assign node22980 = (inp[10]) ? node22982 : 4'b1100;
															assign node22982 = (inp[2]) ? 4'b1100 : 4'b0000;
												assign node22986 = (inp[10]) ? node22992 : node22987;
													assign node22987 = (inp[4]) ? node22989 : 4'b0000;
														assign node22989 = (inp[7]) ? 4'b0000 : 4'b0100;
													assign node22992 = (inp[4]) ? node22994 : 4'b1000;
														assign node22994 = (inp[2]) ? node22998 : node22995;
															assign node22995 = (inp[7]) ? 4'b1000 : 4'b0000;
															assign node22998 = (inp[7]) ? 4'b1000 : 4'b1100;
											assign node23001 = (inp[7]) ? node23019 : node23002;
												assign node23002 = (inp[4]) ? node23012 : node23003;
													assign node23003 = (inp[2]) ? node23007 : node23004;
														assign node23004 = (inp[10]) ? 4'b0100 : 4'b1000;
														assign node23007 = (inp[10]) ? 4'b1100 : node23008;
															assign node23008 = (inp[12]) ? 4'b0100 : 4'b1100;
													assign node23012 = (inp[10]) ? 4'b0000 : node23013;
														assign node23013 = (inp[2]) ? node23015 : 4'b1100;
															assign node23015 = (inp[12]) ? 4'b0000 : 4'b1000;
												assign node23019 = (inp[2]) ? node23027 : node23020;
													assign node23020 = (inp[4]) ? node23024 : node23021;
														assign node23021 = (inp[10]) ? 4'b0000 : 4'b1000;
														assign node23024 = (inp[10]) ? 4'b0100 : 4'b1100;
													assign node23027 = (inp[12]) ? node23029 : 4'b1100;
														assign node23029 = (inp[10]) ? 4'b1100 : 4'b0100;
										assign node23032 = (inp[10]) ? node23076 : node23033;
											assign node23033 = (inp[12]) ? node23055 : node23034;
												assign node23034 = (inp[3]) ? node23042 : node23035;
													assign node23035 = (inp[2]) ? 4'b0100 : node23036;
														assign node23036 = (inp[7]) ? node23038 : 4'b1000;
															assign node23038 = (inp[4]) ? 4'b0100 : 4'b0000;
													assign node23042 = (inp[2]) ? node23050 : node23043;
														assign node23043 = (inp[4]) ? node23047 : node23044;
															assign node23044 = (inp[7]) ? 4'b1000 : 4'b1100;
															assign node23047 = (inp[7]) ? 4'b1100 : 4'b1000;
														assign node23050 = (inp[7]) ? 4'b0000 : node23051;
															assign node23051 = (inp[4]) ? 4'b1000 : 4'b0000;
												assign node23055 = (inp[3]) ? node23063 : node23056;
													assign node23056 = (inp[2]) ? node23058 : 4'b1000;
														assign node23058 = (inp[7]) ? 4'b1000 : node23059;
															assign node23059 = (inp[4]) ? 4'b1100 : 4'b1000;
													assign node23063 = (inp[2]) ? node23071 : node23064;
														assign node23064 = (inp[7]) ? node23068 : node23065;
															assign node23065 = (inp[4]) ? 4'b0000 : 4'b1100;
															assign node23068 = (inp[4]) ? 4'b1100 : 4'b1000;
														assign node23071 = (inp[4]) ? node23073 : 4'b1100;
															assign node23073 = (inp[7]) ? 4'b1100 : 4'b1000;
											assign node23076 = (inp[4]) ? node23096 : node23077;
												assign node23077 = (inp[2]) ? node23083 : node23078;
													assign node23078 = (inp[3]) ? 4'b0100 : node23079;
														assign node23079 = (inp[7]) ? 4'b0000 : 4'b0100;
													assign node23083 = (inp[12]) ? node23089 : node23084;
														assign node23084 = (inp[3]) ? node23086 : 4'b0000;
															assign node23086 = (inp[7]) ? 4'b0100 : 4'b0000;
														assign node23089 = (inp[7]) ? node23093 : node23090;
															assign node23090 = (inp[3]) ? 4'b0000 : 4'b0100;
															assign node23093 = (inp[3]) ? 4'b0100 : 4'b0000;
												assign node23096 = (inp[3]) ? 4'b0000 : node23097;
													assign node23097 = (inp[2]) ? 4'b0100 : 4'b0000;
							assign node23101 = (inp[3]) ? node23475 : node23102;
								assign node23102 = (inp[11]) ? node23332 : node23103;
									assign node23103 = (inp[4]) ? node23215 : node23104;
										assign node23104 = (inp[2]) ? node23180 : node23105;
											assign node23105 = (inp[13]) ? node23137 : node23106;
												assign node23106 = (inp[10]) ? node23114 : node23107;
													assign node23107 = (inp[1]) ? node23111 : node23108;
														assign node23108 = (inp[14]) ? 4'b0001 : 4'b1000;
														assign node23111 = (inp[14]) ? 4'b1000 : 4'b1001;
													assign node23114 = (inp[7]) ? node23126 : node23115;
														assign node23115 = (inp[1]) ? node23121 : node23116;
															assign node23116 = (inp[14]) ? node23118 : 4'b0100;
																assign node23118 = (inp[12]) ? 4'b1001 : 4'b0101;
															assign node23121 = (inp[12]) ? 4'b0100 : node23122;
																assign node23122 = (inp[14]) ? 4'b1100 : 4'b1101;
														assign node23126 = (inp[12]) ? node23132 : node23127;
															assign node23127 = (inp[1]) ? 4'b1001 : node23128;
																assign node23128 = (inp[14]) ? 4'b0001 : 4'b0000;
															assign node23132 = (inp[14]) ? 4'b0000 : node23133;
																assign node23133 = (inp[1]) ? 4'b0001 : 4'b0000;
												assign node23137 = (inp[7]) ? node23157 : node23138;
													assign node23138 = (inp[10]) ? node23150 : node23139;
														assign node23139 = (inp[1]) ? node23145 : node23140;
															assign node23140 = (inp[14]) ? 4'b1101 : node23141;
																assign node23141 = (inp[12]) ? 4'b1100 : 4'b0100;
															assign node23145 = (inp[12]) ? node23147 : 4'b0000;
																assign node23147 = (inp[14]) ? 4'b0100 : 4'b0101;
														assign node23150 = (inp[12]) ? node23154 : node23151;
															assign node23151 = (inp[1]) ? 4'b0000 : 4'b1000;
															assign node23154 = (inp[1]) ? 4'b1000 : 4'b0000;
													assign node23157 = (inp[1]) ? node23169 : node23158;
														assign node23158 = (inp[14]) ? node23164 : node23159;
															assign node23159 = (inp[12]) ? node23161 : 4'b0100;
																assign node23161 = (inp[10]) ? 4'b1100 : 4'b1000;
															assign node23164 = (inp[10]) ? node23166 : 4'b1001;
																assign node23166 = (inp[12]) ? 4'b0101 : 4'b1101;
														assign node23169 = (inp[14]) ? node23173 : node23170;
															assign node23170 = (inp[10]) ? 4'b1101 : 4'b0101;
															assign node23173 = (inp[12]) ? node23177 : node23174;
																assign node23174 = (inp[10]) ? 4'b0000 : 4'b0100;
																assign node23177 = (inp[10]) ? 4'b1100 : 4'b0100;
											assign node23180 = (inp[13]) ? node23194 : node23181;
												assign node23181 = (inp[10]) ? node23187 : node23182;
													assign node23182 = (inp[12]) ? 4'b0001 : node23183;
														assign node23183 = (inp[1]) ? 4'b1001 : 4'b0001;
													assign node23187 = (inp[1]) ? node23189 : 4'b1001;
														assign node23189 = (inp[14]) ? 4'b1001 : node23190;
															assign node23190 = (inp[7]) ? 4'b0001 : 4'b0101;
												assign node23194 = (inp[7]) ? node23208 : node23195;
													assign node23195 = (inp[10]) ? node23201 : node23196;
														assign node23196 = (inp[12]) ? 4'b0101 : node23197;
															assign node23197 = (inp[1]) ? 4'b1101 : 4'b0101;
														assign node23201 = (inp[1]) ? node23203 : 4'b1101;
															assign node23203 = (inp[12]) ? 4'b1101 : node23204;
																assign node23204 = (inp[14]) ? 4'b0000 : 4'b0001;
													assign node23208 = (inp[10]) ? node23210 : 4'b0001;
														assign node23210 = (inp[12]) ? 4'b1001 : node23211;
															assign node23211 = (inp[1]) ? 4'b0101 : 4'b1001;
										assign node23215 = (inp[2]) ? node23267 : node23216;
											assign node23216 = (inp[13]) ? node23244 : node23217;
												assign node23217 = (inp[10]) ? node23227 : node23218;
													assign node23218 = (inp[12]) ? node23224 : node23219;
														assign node23219 = (inp[1]) ? node23221 : 4'b1000;
															assign node23221 = (inp[7]) ? 4'b0000 : 4'b0100;
														assign node23224 = (inp[1]) ? 4'b1000 : 4'b0000;
													assign node23227 = (inp[12]) ? node23237 : node23228;
														assign node23228 = (inp[1]) ? node23232 : node23229;
															assign node23229 = (inp[7]) ? 4'b1000 : 4'b1100;
															assign node23232 = (inp[7]) ? 4'b0100 : node23233;
																assign node23233 = (inp[14]) ? 4'b0001 : 4'b1000;
														assign node23237 = (inp[7]) ? node23241 : node23238;
															assign node23238 = (inp[1]) ? 4'b0000 : 4'b0100;
															assign node23241 = (inp[1]) ? 4'b1000 : 4'b0000;
												assign node23244 = (inp[1]) ? node23260 : node23245;
													assign node23245 = (inp[14]) ? node23253 : node23246;
														assign node23246 = (inp[7]) ? node23250 : node23247;
															assign node23247 = (inp[12]) ? 4'b1001 : 4'b0001;
															assign node23250 = (inp[10]) ? 4'b0001 : 4'b0100;
														assign node23253 = (inp[12]) ? node23255 : 4'b0000;
															assign node23255 = (inp[10]) ? 4'b0100 : node23256;
																assign node23256 = (inp[7]) ? 4'b0100 : 4'b1000;
													assign node23260 = (inp[14]) ? node23264 : node23261;
														assign node23261 = (inp[10]) ? 4'b1001 : 4'b1000;
														assign node23264 = (inp[12]) ? 4'b0001 : 4'b1001;
											assign node23267 = (inp[10]) ? node23301 : node23268;
												assign node23268 = (inp[13]) ? node23284 : node23269;
													assign node23269 = (inp[7]) ? node23279 : node23270;
														assign node23270 = (inp[1]) ? node23276 : node23271;
															assign node23271 = (inp[14]) ? 4'b0001 : node23272;
																assign node23272 = (inp[12]) ? 4'b0000 : 4'b1000;
															assign node23276 = (inp[14]) ? 4'b1000 : 4'b1001;
														assign node23279 = (inp[1]) ? node23281 : 4'b0101;
															assign node23281 = (inp[12]) ? 4'b0101 : 4'b1101;
													assign node23284 = (inp[1]) ? node23292 : node23285;
														assign node23285 = (inp[14]) ? 4'b1001 : node23286;
															assign node23286 = (inp[12]) ? 4'b1000 : node23287;
																assign node23287 = (inp[7]) ? 4'b0000 : 4'b0100;
														assign node23292 = (inp[14]) ? node23298 : node23293;
															assign node23293 = (inp[7]) ? 4'b0001 : node23294;
																assign node23294 = (inp[12]) ? 4'b0101 : 4'b0000;
															assign node23298 = (inp[7]) ? 4'b0000 : 4'b0100;
												assign node23301 = (inp[13]) ? node23317 : node23302;
													assign node23302 = (inp[12]) ? node23310 : node23303;
														assign node23303 = (inp[1]) ? node23307 : node23304;
															assign node23304 = (inp[14]) ? 4'b0001 : 4'b0000;
															assign node23307 = (inp[14]) ? 4'b1000 : 4'b1001;
														assign node23310 = (inp[14]) ? node23314 : node23311;
															assign node23311 = (inp[1]) ? 4'b0001 : 4'b0000;
															assign node23314 = (inp[1]) ? 4'b0000 : 4'b1001;
													assign node23317 = (inp[7]) ? node23325 : node23318;
														assign node23318 = (inp[1]) ? node23322 : node23319;
															assign node23319 = (inp[12]) ? 4'b0000 : 4'b1000;
															assign node23322 = (inp[12]) ? 4'b1000 : 4'b0000;
														assign node23325 = (inp[14]) ? node23329 : node23326;
															assign node23326 = (inp[1]) ? 4'b0000 : 4'b1000;
															assign node23329 = (inp[1]) ? 4'b1000 : 4'b1001;
									assign node23332 = (inp[1]) ? node23412 : node23333;
										assign node23333 = (inp[4]) ? node23373 : node23334;
											assign node23334 = (inp[2]) ? node23352 : node23335;
												assign node23335 = (inp[13]) ? node23343 : node23336;
													assign node23336 = (inp[10]) ? node23340 : node23337;
														assign node23337 = (inp[12]) ? 4'b0001 : 4'b1001;
														assign node23340 = (inp[7]) ? 4'b0001 : 4'b0101;
													assign node23343 = (inp[10]) ? node23349 : node23344;
														assign node23344 = (inp[12]) ? node23346 : 4'b0101;
															assign node23346 = (inp[7]) ? 4'b1001 : 4'b1101;
														assign node23349 = (inp[7]) ? 4'b1101 : 4'b1000;
												assign node23352 = (inp[13]) ? node23360 : node23353;
													assign node23353 = (inp[12]) ? node23357 : node23354;
														assign node23354 = (inp[10]) ? 4'b0000 : 4'b1000;
														assign node23357 = (inp[10]) ? 4'b1000 : 4'b0000;
													assign node23360 = (inp[7]) ? node23366 : node23361;
														assign node23361 = (inp[12]) ? node23363 : 4'b1100;
															assign node23363 = (inp[10]) ? 4'b1100 : 4'b0100;
														assign node23366 = (inp[12]) ? node23370 : node23367;
															assign node23367 = (inp[10]) ? 4'b0100 : 4'b1000;
															assign node23370 = (inp[10]) ? 4'b1000 : 4'b0000;
											assign node23373 = (inp[13]) ? node23391 : node23374;
												assign node23374 = (inp[2]) ? node23384 : node23375;
													assign node23375 = (inp[7]) ? 4'b1000 : node23376;
														assign node23376 = (inp[12]) ? node23380 : node23377;
															assign node23377 = (inp[10]) ? 4'b0001 : 4'b1000;
															assign node23380 = (inp[10]) ? 4'b1100 : 4'b1000;
													assign node23384 = (inp[10]) ? 4'b0001 : node23385;
														assign node23385 = (inp[7]) ? node23387 : 4'b1001;
															assign node23387 = (inp[12]) ? 4'b0100 : 4'b1100;
												assign node23391 = (inp[10]) ? node23401 : node23392;
													assign node23392 = (inp[12]) ? node23398 : node23393;
														assign node23393 = (inp[7]) ? 4'b0001 : node23394;
															assign node23394 = (inp[2]) ? 4'b0101 : 4'b0001;
														assign node23398 = (inp[2]) ? 4'b1001 : 4'b0001;
													assign node23401 = (inp[7]) ? node23407 : node23402;
														assign node23402 = (inp[12]) ? node23404 : 4'b1000;
															assign node23404 = (inp[2]) ? 4'b1000 : 4'b0000;
														assign node23407 = (inp[12]) ? node23409 : 4'b1001;
															assign node23409 = (inp[2]) ? 4'b1001 : 4'b0001;
										assign node23412 = (inp[13]) ? node23444 : node23413;
											assign node23413 = (inp[2]) ? node23429 : node23414;
												assign node23414 = (inp[10]) ? node23422 : node23415;
													assign node23415 = (inp[7]) ? 4'b0000 : node23416;
														assign node23416 = (inp[12]) ? node23418 : 4'b0100;
															assign node23418 = (inp[4]) ? 4'b0100 : 4'b1000;
													assign node23422 = (inp[7]) ? node23426 : node23423;
														assign node23423 = (inp[4]) ? 4'b1000 : 4'b1100;
														assign node23426 = (inp[4]) ? 4'b0100 : 4'b1000;
												assign node23429 = (inp[7]) ? node23435 : node23430;
													assign node23430 = (inp[4]) ? 4'b1000 : node23431;
														assign node23431 = (inp[10]) ? 4'b0100 : 4'b1000;
													assign node23435 = (inp[10]) ? node23441 : node23436;
														assign node23436 = (inp[4]) ? node23438 : 4'b1000;
															assign node23438 = (inp[12]) ? 4'b1100 : 4'b0000;
														assign node23441 = (inp[4]) ? 4'b1000 : 4'b0000;
											assign node23444 = (inp[10]) ? node23468 : node23445;
												assign node23445 = (inp[4]) ? node23455 : node23446;
													assign node23446 = (inp[2]) ? node23452 : node23447;
														assign node23447 = (inp[7]) ? node23449 : 4'b0000;
															assign node23449 = (inp[12]) ? 4'b0100 : 4'b1100;
														assign node23452 = (inp[7]) ? 4'b1000 : 4'b1100;
													assign node23455 = (inp[7]) ? node23461 : node23456;
														assign node23456 = (inp[2]) ? 4'b0000 : node23457;
															assign node23457 = (inp[12]) ? 4'b1000 : 4'b0100;
														assign node23461 = (inp[12]) ? node23465 : node23462;
															assign node23462 = (inp[2]) ? 4'b1000 : 4'b0000;
															assign node23465 = (inp[2]) ? 4'b0000 : 4'b1000;
												assign node23468 = (inp[4]) ? 4'b0000 : node23469;
													assign node23469 = (inp[7]) ? node23471 : 4'b0000;
														assign node23471 = (inp[2]) ? 4'b0100 : 4'b0000;
								assign node23475 = (inp[1]) ? node23689 : node23476;
									assign node23476 = (inp[13]) ? node23592 : node23477;
										assign node23477 = (inp[2]) ? node23541 : node23478;
											assign node23478 = (inp[12]) ? node23508 : node23479;
												assign node23479 = (inp[14]) ? node23499 : node23480;
													assign node23480 = (inp[7]) ? node23490 : node23481;
														assign node23481 = (inp[4]) ? node23485 : node23482;
															assign node23482 = (inp[11]) ? 4'b0000 : 4'b1000;
															assign node23485 = (inp[11]) ? 4'b0001 : node23486;
																assign node23486 = (inp[10]) ? 4'b0000 : 4'b0001;
														assign node23490 = (inp[10]) ? node23494 : node23491;
															assign node23491 = (inp[4]) ? 4'b0001 : 4'b1001;
															assign node23494 = (inp[11]) ? 4'b1001 : node23495;
																assign node23495 = (inp[4]) ? 4'b1001 : 4'b1000;
													assign node23499 = (inp[4]) ? 4'b0001 : node23500;
														assign node23500 = (inp[11]) ? node23502 : 4'b0001;
															assign node23502 = (inp[10]) ? 4'b0000 : node23503;
																assign node23503 = (inp[7]) ? 4'b0000 : 4'b0001;
												assign node23508 = (inp[11]) ? node23528 : node23509;
													assign node23509 = (inp[4]) ? node23515 : node23510;
														assign node23510 = (inp[14]) ? 4'b0001 : node23511;
															assign node23511 = (inp[10]) ? 4'b0000 : 4'b0001;
														assign node23515 = (inp[10]) ? node23521 : node23516;
															assign node23516 = (inp[7]) ? 4'b1000 : node23517;
																assign node23517 = (inp[14]) ? 4'b1000 : 4'b1001;
															assign node23521 = (inp[14]) ? node23525 : node23522;
																assign node23522 = (inp[7]) ? 4'b0001 : 4'b0000;
																assign node23525 = (inp[7]) ? 4'b0000 : 4'b1001;
													assign node23528 = (inp[7]) ? node23534 : node23529;
														assign node23529 = (inp[10]) ? node23531 : 4'b1000;
															assign node23531 = (inp[4]) ? 4'b1000 : 4'b0000;
														assign node23534 = (inp[4]) ? node23538 : node23535;
															assign node23535 = (inp[10]) ? 4'b1001 : 4'b1000;
															assign node23538 = (inp[10]) ? 4'b0001 : 4'b1001;
											assign node23541 = (inp[4]) ? node23561 : node23542;
												assign node23542 = (inp[10]) ? node23548 : node23543;
													assign node23543 = (inp[11]) ? 4'b1000 : node23544;
														assign node23544 = (inp[12]) ? 4'b0000 : 4'b1000;
													assign node23548 = (inp[11]) ? node23556 : node23549;
														assign node23549 = (inp[14]) ? node23551 : 4'b1001;
															assign node23551 = (inp[12]) ? node23553 : 4'b1000;
																assign node23553 = (inp[7]) ? 4'b0000 : 4'b1000;
														assign node23556 = (inp[12]) ? node23558 : 4'b0001;
															assign node23558 = (inp[7]) ? 4'b1000 : 4'b1001;
												assign node23561 = (inp[10]) ? node23573 : node23562;
													assign node23562 = (inp[11]) ? node23568 : node23563;
														assign node23563 = (inp[14]) ? 4'b1000 : node23564;
															assign node23564 = (inp[7]) ? 4'b1000 : 4'b1001;
														assign node23568 = (inp[7]) ? 4'b0001 : node23569;
															assign node23569 = (inp[12]) ? 4'b0000 : 4'b1000;
													assign node23573 = (inp[7]) ? node23583 : node23574;
														assign node23574 = (inp[12]) ? node23578 : node23575;
															assign node23575 = (inp[11]) ? 4'b1000 : 4'b0000;
															assign node23578 = (inp[14]) ? 4'b0000 : node23579;
																assign node23579 = (inp[11]) ? 4'b0000 : 4'b0001;
														assign node23583 = (inp[12]) ? node23587 : node23584;
															assign node23584 = (inp[11]) ? 4'b0001 : 4'b0000;
															assign node23587 = (inp[11]) ? 4'b1000 : node23588;
																assign node23588 = (inp[14]) ? 4'b0001 : 4'b1000;
										assign node23592 = (inp[4]) ? node23644 : node23593;
											assign node23593 = (inp[7]) ? node23615 : node23594;
												assign node23594 = (inp[11]) ? node23612 : node23595;
													assign node23595 = (inp[2]) ? node23607 : node23596;
														assign node23596 = (inp[12]) ? node23602 : node23597;
															assign node23597 = (inp[10]) ? 4'b0000 : node23598;
																assign node23598 = (inp[14]) ? 4'b0000 : 4'b0001;
															assign node23602 = (inp[14]) ? 4'b0001 : node23603;
																assign node23603 = (inp[10]) ? 4'b0000 : 4'b0001;
														assign node23607 = (inp[14]) ? 4'b1001 : node23608;
															assign node23608 = (inp[10]) ? 4'b1000 : 4'b1001;
													assign node23612 = (inp[2]) ? 4'b0000 : 4'b1001;
												assign node23615 = (inp[12]) ? node23633 : node23616;
													assign node23616 = (inp[10]) ? node23624 : node23617;
														assign node23617 = (inp[11]) ? 4'b0000 : node23618;
															assign node23618 = (inp[2]) ? node23620 : 4'b1000;
																assign node23620 = (inp[14]) ? 4'b0000 : 4'b0001;
														assign node23624 = (inp[14]) ? 4'b0001 : node23625;
															assign node23625 = (inp[11]) ? node23629 : node23626;
																assign node23626 = (inp[2]) ? 4'b0000 : 4'b0001;
																assign node23629 = (inp[2]) ? 4'b0001 : 4'b0000;
													assign node23633 = (inp[2]) ? node23641 : node23634;
														assign node23634 = (inp[11]) ? node23638 : node23635;
															assign node23635 = (inp[10]) ? 4'b0001 : 4'b1000;
															assign node23638 = (inp[10]) ? 4'b1000 : 4'b0000;
														assign node23641 = (inp[11]) ? 4'b0001 : 4'b1001;
											assign node23644 = (inp[11]) ? node23672 : node23645;
												assign node23645 = (inp[12]) ? node23663 : node23646;
													assign node23646 = (inp[7]) ? node23654 : node23647;
														assign node23647 = (inp[10]) ? node23649 : 4'b0001;
															assign node23649 = (inp[14]) ? node23651 : 4'b0001;
																assign node23651 = (inp[2]) ? 4'b0000 : 4'b0001;
														assign node23654 = (inp[14]) ? node23660 : node23655;
															assign node23655 = (inp[2]) ? 4'b0000 : node23656;
																assign node23656 = (inp[10]) ? 4'b0001 : 4'b0000;
															assign node23660 = (inp[10]) ? 4'b0000 : 4'b0001;
													assign node23663 = (inp[7]) ? node23669 : node23664;
														assign node23664 = (inp[2]) ? 4'b0000 : node23665;
															assign node23665 = (inp[10]) ? 4'b0000 : 4'b0001;
														assign node23669 = (inp[2]) ? 4'b0001 : 4'b0000;
												assign node23672 = (inp[10]) ? 4'b0000 : node23673;
													assign node23673 = (inp[14]) ? node23681 : node23674;
														assign node23674 = (inp[12]) ? node23676 : 4'b0000;
															assign node23676 = (inp[7]) ? node23678 : 4'b0000;
																assign node23678 = (inp[2]) ? 4'b0001 : 4'b0000;
														assign node23681 = (inp[12]) ? node23685 : node23682;
															assign node23682 = (inp[2]) ? 4'b0000 : 4'b0001;
															assign node23685 = (inp[2]) ? 4'b0001 : 4'b0000;
									assign node23689 = (inp[11]) ? node23795 : node23690;
										assign node23690 = (inp[4]) ? node23754 : node23691;
											assign node23691 = (inp[10]) ? node23723 : node23692;
												assign node23692 = (inp[13]) ? node23710 : node23693;
													assign node23693 = (inp[2]) ? node23703 : node23694;
														assign node23694 = (inp[7]) ? 4'b0001 : node23695;
															assign node23695 = (inp[14]) ? node23699 : node23696;
																assign node23696 = (inp[12]) ? 4'b0001 : 4'b1001;
																assign node23699 = (inp[12]) ? 4'b0000 : 4'b1000;
														assign node23703 = (inp[12]) ? node23705 : 4'b0000;
															assign node23705 = (inp[14]) ? 4'b1000 : node23706;
																assign node23706 = (inp[7]) ? 4'b1000 : 4'b0000;
													assign node23710 = (inp[14]) ? node23718 : node23711;
														assign node23711 = (inp[2]) ? 4'b0001 : node23712;
															assign node23712 = (inp[12]) ? 4'b0000 : node23713;
																assign node23713 = (inp[7]) ? 4'b1000 : 4'b0001;
														assign node23718 = (inp[12]) ? 4'b0001 : node23719;
															assign node23719 = (inp[7]) ? 4'b0001 : 4'b0000;
												assign node23723 = (inp[7]) ? node23735 : node23724;
													assign node23724 = (inp[12]) ? node23726 : 4'b1000;
														assign node23726 = (inp[14]) ? node23728 : 4'b1000;
															assign node23728 = (inp[13]) ? node23732 : node23729;
																assign node23729 = (inp[2]) ? 4'b0001 : 4'b1000;
																assign node23732 = (inp[2]) ? 4'b1000 : 4'b0000;
													assign node23735 = (inp[13]) ? node23745 : node23736;
														assign node23736 = (inp[2]) ? node23740 : node23737;
															assign node23737 = (inp[14]) ? 4'b0000 : 4'b0001;
															assign node23740 = (inp[14]) ? 4'b0001 : node23741;
																assign node23741 = (inp[12]) ? 4'b0000 : 4'b1000;
														assign node23745 = (inp[14]) ? node23749 : node23746;
															assign node23746 = (inp[2]) ? 4'b1001 : 4'b0001;
															assign node23749 = (inp[2]) ? 4'b1000 : node23750;
																assign node23750 = (inp[12]) ? 4'b0000 : 4'b1000;
											assign node23754 = (inp[10]) ? node23782 : node23755;
												assign node23755 = (inp[7]) ? node23771 : node23756;
													assign node23756 = (inp[12]) ? node23762 : node23757;
														assign node23757 = (inp[13]) ? 4'b0001 : node23758;
															assign node23758 = (inp[14]) ? 4'b0000 : 4'b0001;
														assign node23762 = (inp[2]) ? node23766 : node23763;
															assign node23763 = (inp[14]) ? 4'b0001 : 4'b0000;
															assign node23766 = (inp[13]) ? 4'b0000 : node23767;
																assign node23767 = (inp[14]) ? 4'b0000 : 4'b0001;
													assign node23771 = (inp[12]) ? node23777 : node23772;
														assign node23772 = (inp[2]) ? 4'b0001 : node23773;
															assign node23773 = (inp[13]) ? 4'b0001 : 4'b0000;
														assign node23777 = (inp[13]) ? node23779 : 4'b1001;
															assign node23779 = (inp[14]) ? 4'b0001 : 4'b0000;
												assign node23782 = (inp[13]) ? 4'b0000 : node23783;
													assign node23783 = (inp[7]) ? node23789 : node23784;
														assign node23784 = (inp[2]) ? 4'b0000 : node23785;
															assign node23785 = (inp[14]) ? 4'b0000 : 4'b0001;
														assign node23789 = (inp[14]) ? 4'b0001 : node23790;
															assign node23790 = (inp[2]) ? 4'b0001 : 4'b1000;
										assign node23795 = (inp[10]) ? node23831 : node23796;
											assign node23796 = (inp[4]) ? node23818 : node23797;
												assign node23797 = (inp[13]) ? node23807 : node23798;
													assign node23798 = (inp[2]) ? node23802 : node23799;
														assign node23799 = (inp[12]) ? 4'b1000 : 4'b0000;
														assign node23802 = (inp[12]) ? 4'b0000 : node23803;
															assign node23803 = (inp[7]) ? 4'b0000 : 4'b1000;
													assign node23807 = (inp[12]) ? node23813 : node23808;
														assign node23808 = (inp[7]) ? node23810 : 4'b1000;
															assign node23810 = (inp[2]) ? 4'b1000 : 4'b0000;
														assign node23813 = (inp[7]) ? 4'b1000 : node23814;
															assign node23814 = (inp[2]) ? 4'b0000 : 4'b1000;
												assign node23818 = (inp[13]) ? 4'b0000 : node23819;
													assign node23819 = (inp[2]) ? node23825 : node23820;
														assign node23820 = (inp[7]) ? 4'b0000 : node23821;
															assign node23821 = (inp[12]) ? 4'b0000 : 4'b1000;
														assign node23825 = (inp[7]) ? node23827 : 4'b0000;
															assign node23827 = (inp[12]) ? 4'b1000 : 4'b0000;
											assign node23831 = (inp[7]) ? node23833 : 4'b0000;
												assign node23833 = (inp[12]) ? node23835 : 4'b0000;
													assign node23835 = (inp[4]) ? 4'b0000 : node23836;
														assign node23836 = (inp[2]) ? node23838 : 4'b0000;
															assign node23838 = (inp[13]) ? 4'b0000 : 4'b1000;
					assign node23842 = (inp[6]) ? node23844 : 4'b0000;
						assign node23844 = (inp[2]) ? node24310 : node23845;
							assign node23845 = (inp[5]) ? node23935 : node23846;
								assign node23846 = (inp[3]) ? node23848 : 4'b0000;
									assign node23848 = (inp[4]) ? node23860 : node23849;
										assign node23849 = (inp[12]) ? 4'b0000 : node23850;
											assign node23850 = (inp[1]) ? 4'b0000 : node23851;
												assign node23851 = (inp[7]) ? 4'b0000 : node23852;
													assign node23852 = (inp[10]) ? node23854 : 4'b0000;
														assign node23854 = (inp[13]) ? 4'b0001 : 4'b0000;
										assign node23860 = (inp[7]) ? node23920 : node23861;
											assign node23861 = (inp[1]) ? node23893 : node23862;
												assign node23862 = (inp[14]) ? node23874 : node23863;
													assign node23863 = (inp[13]) ? node23869 : node23864;
														assign node23864 = (inp[10]) ? node23866 : 4'b0001;
															assign node23866 = (inp[12]) ? 4'b0001 : 4'b1001;
														assign node23869 = (inp[10]) ? node23871 : 4'b1001;
															assign node23871 = (inp[12]) ? 4'b1001 : 4'b0001;
													assign node23874 = (inp[11]) ? node23884 : node23875;
														assign node23875 = (inp[13]) ? node23881 : node23876;
															assign node23876 = (inp[12]) ? 4'b0000 : node23877;
																assign node23877 = (inp[10]) ? 4'b1000 : 4'b0000;
															assign node23881 = (inp[12]) ? 4'b1000 : 4'b0000;
														assign node23884 = (inp[13]) ? node23890 : node23885;
															assign node23885 = (inp[10]) ? node23887 : 4'b0001;
																assign node23887 = (inp[12]) ? 4'b0001 : 4'b1001;
															assign node23890 = (inp[12]) ? 4'b1001 : 4'b0001;
												assign node23893 = (inp[14]) ? node23905 : node23894;
													assign node23894 = (inp[13]) ? node23900 : node23895;
														assign node23895 = (inp[10]) ? 4'b1000 : node23896;
															assign node23896 = (inp[12]) ? 4'b0000 : 4'b1000;
														assign node23900 = (inp[10]) ? 4'b0000 : node23901;
															assign node23901 = (inp[12]) ? 4'b1000 : 4'b0000;
													assign node23905 = (inp[11]) ? node23915 : node23906;
														assign node23906 = (inp[12]) ? 4'b0001 : node23907;
															assign node23907 = (inp[10]) ? node23911 : node23908;
																assign node23908 = (inp[13]) ? 4'b1001 : 4'b0001;
																assign node23911 = (inp[13]) ? 4'b0001 : 4'b1001;
														assign node23915 = (inp[13]) ? 4'b0000 : node23916;
															assign node23916 = (inp[12]) ? 4'b0000 : 4'b1000;
											assign node23920 = (inp[13]) ? node23922 : 4'b0000;
												assign node23922 = (inp[12]) ? 4'b0000 : node23923;
													assign node23923 = (inp[10]) ? node23925 : 4'b0000;
														assign node23925 = (inp[11]) ? 4'b0000 : node23926;
															assign node23926 = (inp[14]) ? node23930 : node23927;
																assign node23927 = (inp[1]) ? 4'b0000 : 4'b0001;
																assign node23930 = (inp[1]) ? 4'b0001 : 4'b0000;
								assign node23935 = (inp[1]) ? node24145 : node23936;
									assign node23936 = (inp[3]) ? node24036 : node23937;
										assign node23937 = (inp[13]) ? node23979 : node23938;
											assign node23938 = (inp[7]) ? node23964 : node23939;
												assign node23939 = (inp[4]) ? node23949 : node23940;
													assign node23940 = (inp[11]) ? node23944 : node23941;
														assign node23941 = (inp[14]) ? 4'b0000 : 4'b0001;
														assign node23944 = (inp[12]) ? 4'b0001 : node23945;
															assign node23945 = (inp[10]) ? 4'b1001 : 4'b0001;
													assign node23949 = (inp[12]) ? node23959 : node23950;
														assign node23950 = (inp[10]) ? node23956 : node23951;
															assign node23951 = (inp[11]) ? 4'b0101 : node23952;
																assign node23952 = (inp[14]) ? 4'b0100 : 4'b0101;
															assign node23956 = (inp[11]) ? 4'b0000 : 4'b1100;
														assign node23959 = (inp[14]) ? node23961 : 4'b0101;
															assign node23961 = (inp[11]) ? 4'b0101 : 4'b0100;
												assign node23964 = (inp[11]) ? node23974 : node23965;
													assign node23965 = (inp[14]) ? node23969 : node23966;
														assign node23966 = (inp[12]) ? 4'b0001 : 4'b1001;
														assign node23969 = (inp[10]) ? node23971 : 4'b0000;
															assign node23971 = (inp[12]) ? 4'b0000 : 4'b1000;
													assign node23974 = (inp[10]) ? node23976 : 4'b0001;
														assign node23976 = (inp[12]) ? 4'b0001 : 4'b1001;
											assign node23979 = (inp[12]) ? node24013 : node23980;
												assign node23980 = (inp[10]) ? node23994 : node23981;
													assign node23981 = (inp[11]) ? node23989 : node23982;
														assign node23982 = (inp[4]) ? node23986 : node23983;
															assign node23983 = (inp[14]) ? 4'b1000 : 4'b1001;
															assign node23986 = (inp[7]) ? 4'b1001 : 4'b0001;
														assign node23989 = (inp[7]) ? 4'b1001 : node23990;
															assign node23990 = (inp[4]) ? 4'b1000 : 4'b1001;
													assign node23994 = (inp[4]) ? node24006 : node23995;
														assign node23995 = (inp[7]) ? node24001 : node23996;
															assign node23996 = (inp[14]) ? node23998 : 4'b0101;
																assign node23998 = (inp[11]) ? 4'b0101 : 4'b0100;
															assign node24001 = (inp[14]) ? node24003 : 4'b0001;
																assign node24003 = (inp[11]) ? 4'b0001 : 4'b0000;
														assign node24006 = (inp[11]) ? 4'b0000 : node24007;
															assign node24007 = (inp[7]) ? node24009 : 4'b1001;
																assign node24009 = (inp[14]) ? 4'b0100 : 4'b0101;
												assign node24013 = (inp[14]) ? node24021 : node24014;
													assign node24014 = (inp[4]) ? node24016 : 4'b1001;
														assign node24016 = (inp[7]) ? 4'b1001 : node24017;
															assign node24017 = (inp[11]) ? 4'b0000 : 4'b0001;
													assign node24021 = (inp[4]) ? node24025 : node24022;
														assign node24022 = (inp[11]) ? 4'b1001 : 4'b1000;
														assign node24025 = (inp[7]) ? node24033 : node24026;
															assign node24026 = (inp[10]) ? node24030 : node24027;
																assign node24027 = (inp[11]) ? 4'b0000 : 4'b0001;
																assign node24030 = (inp[11]) ? 4'b1000 : 4'b1001;
															assign node24033 = (inp[11]) ? 4'b1001 : 4'b1000;
										assign node24036 = (inp[4]) ? node24086 : node24037;
											assign node24037 = (inp[10]) ? node24061 : node24038;
												assign node24038 = (inp[11]) ? node24050 : node24039;
													assign node24039 = (inp[13]) ? node24041 : 4'b0001;
														assign node24041 = (inp[14]) ? node24047 : node24042;
															assign node24042 = (inp[12]) ? node24044 : 4'b0000;
																assign node24044 = (inp[7]) ? 4'b0001 : 4'b1000;
															assign node24047 = (inp[7]) ? 4'b0001 : 4'b1001;
													assign node24050 = (inp[13]) ? node24054 : node24051;
														assign node24051 = (inp[12]) ? 4'b0000 : 4'b1000;
														assign node24054 = (inp[7]) ? node24058 : node24055;
															assign node24055 = (inp[12]) ? 4'b1001 : 4'b0001;
															assign node24058 = (inp[12]) ? 4'b0000 : 4'b0001;
												assign node24061 = (inp[7]) ? node24073 : node24062;
													assign node24062 = (inp[13]) ? node24070 : node24063;
														assign node24063 = (inp[14]) ? node24067 : node24064;
															assign node24064 = (inp[11]) ? 4'b0001 : 4'b0000;
															assign node24067 = (inp[12]) ? 4'b1001 : 4'b0001;
														assign node24070 = (inp[12]) ? 4'b0000 : 4'b1000;
													assign node24073 = (inp[12]) ? node24081 : node24074;
														assign node24074 = (inp[11]) ? node24078 : node24075;
															assign node24075 = (inp[13]) ? 4'b1000 : 4'b1001;
															assign node24078 = (inp[13]) ? 4'b1001 : 4'b0000;
														assign node24081 = (inp[13]) ? node24083 : 4'b1001;
															assign node24083 = (inp[11]) ? 4'b1001 : 4'b0001;
											assign node24086 = (inp[13]) ? node24118 : node24087;
												assign node24087 = (inp[10]) ? node24101 : node24088;
													assign node24088 = (inp[7]) ? node24096 : node24089;
														assign node24089 = (inp[12]) ? 4'b1001 : node24090;
															assign node24090 = (inp[11]) ? 4'b0000 : node24091;
																assign node24091 = (inp[14]) ? 4'b1000 : 4'b1001;
														assign node24096 = (inp[12]) ? node24098 : 4'b1000;
															assign node24098 = (inp[11]) ? 4'b1000 : 4'b0000;
													assign node24101 = (inp[11]) ? node24113 : node24102;
														assign node24102 = (inp[14]) ? node24108 : node24103;
															assign node24103 = (inp[7]) ? 4'b0001 : node24104;
																assign node24104 = (inp[12]) ? 4'b0000 : 4'b1000;
															assign node24108 = (inp[7]) ? node24110 : 4'b0001;
																assign node24110 = (inp[12]) ? 4'b1000 : 4'b0001;
														assign node24113 = (inp[7]) ? node24115 : 4'b0000;
															assign node24115 = (inp[12]) ? 4'b0000 : 4'b1000;
												assign node24118 = (inp[10]) ? node24136 : node24119;
													assign node24119 = (inp[14]) ? node24129 : node24120;
														assign node24120 = (inp[7]) ? node24124 : node24121;
															assign node24121 = (inp[11]) ? 4'b0001 : 4'b0000;
															assign node24124 = (inp[11]) ? node24126 : 4'b0001;
																assign node24126 = (inp[12]) ? 4'b0000 : 4'b0001;
														assign node24129 = (inp[7]) ? node24133 : node24130;
															assign node24130 = (inp[12]) ? 4'b0001 : 4'b0000;
															assign node24133 = (inp[12]) ? 4'b0000 : 4'b0001;
													assign node24136 = (inp[11]) ? 4'b0000 : node24137;
														assign node24137 = (inp[14]) ? node24139 : 4'b0000;
															assign node24139 = (inp[7]) ? node24141 : 4'b0001;
																assign node24141 = (inp[12]) ? 4'b0000 : 4'b0001;
									assign node24145 = (inp[11]) ? node24253 : node24146;
										assign node24146 = (inp[3]) ? node24208 : node24147;
											assign node24147 = (inp[14]) ? node24183 : node24148;
												assign node24148 = (inp[4]) ? node24162 : node24149;
													assign node24149 = (inp[13]) ? node24155 : node24150;
														assign node24150 = (inp[10]) ? 4'b1000 : node24151;
															assign node24151 = (inp[12]) ? 4'b0000 : 4'b1000;
														assign node24155 = (inp[10]) ? 4'b0100 : node24156;
															assign node24156 = (inp[12]) ? 4'b1000 : node24157;
																assign node24157 = (inp[7]) ? 4'b0000 : 4'b0100;
													assign node24162 = (inp[12]) ? node24172 : node24163;
														assign node24163 = (inp[10]) ? 4'b0001 : node24164;
															assign node24164 = (inp[7]) ? node24168 : node24165;
																assign node24165 = (inp[13]) ? 4'b1001 : 4'b1100;
																assign node24168 = (inp[13]) ? 4'b0100 : 4'b1000;
														assign node24172 = (inp[13]) ? node24178 : node24173;
															assign node24173 = (inp[10]) ? node24175 : 4'b0100;
																assign node24175 = (inp[7]) ? 4'b1000 : 4'b1100;
															assign node24178 = (inp[7]) ? node24180 : 4'b1001;
																assign node24180 = (inp[10]) ? 4'b0100 : 4'b1000;
												assign node24183 = (inp[13]) ? node24199 : node24184;
													assign node24184 = (inp[4]) ? node24190 : node24185;
														assign node24185 = (inp[10]) ? node24187 : 4'b0001;
															assign node24187 = (inp[12]) ? 4'b0001 : 4'b1001;
														assign node24190 = (inp[7]) ? node24196 : node24191;
															assign node24191 = (inp[10]) ? node24193 : 4'b0101;
																assign node24193 = (inp[12]) ? 4'b0101 : 4'b0001;
															assign node24196 = (inp[10]) ? 4'b1001 : 4'b0001;
													assign node24199 = (inp[10]) ? node24201 : 4'b1001;
														assign node24201 = (inp[12]) ? 4'b1001 : node24202;
															assign node24202 = (inp[4]) ? 4'b0001 : node24203;
																assign node24203 = (inp[7]) ? 4'b0001 : 4'b0101;
											assign node24208 = (inp[13]) ? node24240 : node24209;
												assign node24209 = (inp[4]) ? node24223 : node24210;
													assign node24210 = (inp[12]) ? node24216 : node24211;
														assign node24211 = (inp[10]) ? node24213 : 4'b1001;
															assign node24213 = (inp[7]) ? 4'b0001 : 4'b1001;
														assign node24216 = (inp[7]) ? node24220 : node24217;
															assign node24217 = (inp[14]) ? 4'b0000 : 4'b0001;
															assign node24220 = (inp[10]) ? 4'b1001 : 4'b0001;
													assign node24223 = (inp[7]) ? node24229 : node24224;
														assign node24224 = (inp[10]) ? node24226 : 4'b0001;
															assign node24226 = (inp[14]) ? 4'b0001 : 4'b0000;
														assign node24229 = (inp[12]) ? node24235 : node24230;
															assign node24230 = (inp[10]) ? 4'b0000 : node24231;
																assign node24231 = (inp[14]) ? 4'b0001 : 4'b0000;
															assign node24235 = (inp[14]) ? 4'b1000 : node24236;
																assign node24236 = (inp[10]) ? 4'b0001 : 4'b0000;
												assign node24240 = (inp[4]) ? 4'b0000 : node24241;
													assign node24241 = (inp[12]) ? node24247 : node24242;
														assign node24242 = (inp[7]) ? node24244 : 4'b0000;
															assign node24244 = (inp[14]) ? 4'b0000 : 4'b0001;
														assign node24247 = (inp[14]) ? 4'b1000 : node24248;
															assign node24248 = (inp[10]) ? 4'b1001 : 4'b0001;
										assign node24253 = (inp[13]) ? node24287 : node24254;
											assign node24254 = (inp[3]) ? node24272 : node24255;
												assign node24255 = (inp[12]) ? node24263 : node24256;
													assign node24256 = (inp[7]) ? 4'b1000 : node24257;
														assign node24257 = (inp[4]) ? node24259 : 4'b1000;
															assign node24259 = (inp[10]) ? 4'b0000 : 4'b1100;
													assign node24263 = (inp[10]) ? node24267 : node24264;
														assign node24264 = (inp[4]) ? 4'b0100 : 4'b0000;
														assign node24267 = (inp[4]) ? node24269 : 4'b1000;
															assign node24269 = (inp[7]) ? 4'b1000 : 4'b0000;
												assign node24272 = (inp[10]) ? node24282 : node24273;
													assign node24273 = (inp[7]) ? node24277 : node24274;
														assign node24274 = (inp[12]) ? 4'b1000 : 4'b0000;
														assign node24277 = (inp[4]) ? node24279 : 4'b1000;
															assign node24279 = (inp[12]) ? 4'b0000 : 4'b1000;
													assign node24282 = (inp[7]) ? 4'b0000 : node24283;
														assign node24283 = (inp[4]) ? 4'b0000 : 4'b1000;
											assign node24287 = (inp[10]) ? node24303 : node24288;
												assign node24288 = (inp[3]) ? node24296 : node24289;
													assign node24289 = (inp[12]) ? 4'b1000 : node24290;
														assign node24290 = (inp[4]) ? 4'b0100 : node24291;
															assign node24291 = (inp[7]) ? 4'b0000 : 4'b0100;
													assign node24296 = (inp[7]) ? node24298 : 4'b0000;
														assign node24298 = (inp[4]) ? 4'b0000 : node24299;
															assign node24299 = (inp[12]) ? 4'b0000 : 4'b1000;
												assign node24303 = (inp[7]) ? 4'b0000 : node24304;
													assign node24304 = (inp[4]) ? 4'b0000 : node24305;
														assign node24305 = (inp[3]) ? 4'b0000 : 4'b0100;
							assign node24310 = (inp[5]) ? node24312 : 4'b0000;
								assign node24312 = (inp[3]) ? node24314 : 4'b0000;
									assign node24314 = (inp[7]) ? node24380 : node24315;
										assign node24315 = (inp[4]) ? node24325 : node24316;
											assign node24316 = (inp[13]) ? node24318 : 4'b0000;
												assign node24318 = (inp[10]) ? node24320 : 4'b0000;
													assign node24320 = (inp[12]) ? 4'b0000 : node24321;
														assign node24321 = (inp[1]) ? 4'b0000 : 4'b0001;
											assign node24325 = (inp[11]) ? node24361 : node24326;
												assign node24326 = (inp[13]) ? node24346 : node24327;
													assign node24327 = (inp[12]) ? node24337 : node24328;
														assign node24328 = (inp[1]) ? node24334 : node24329;
															assign node24329 = (inp[10]) ? node24331 : 4'b0001;
																assign node24331 = (inp[14]) ? 4'b1000 : 4'b1001;
															assign node24334 = (inp[10]) ? 4'b0001 : 4'b1000;
														assign node24337 = (inp[1]) ? node24341 : node24338;
															assign node24338 = (inp[14]) ? 4'b0000 : 4'b0001;
															assign node24341 = (inp[10]) ? 4'b1000 : node24342;
																assign node24342 = (inp[14]) ? 4'b0001 : 4'b0000;
													assign node24346 = (inp[1]) ? node24356 : node24347;
														assign node24347 = (inp[12]) ? node24351 : node24348;
															assign node24348 = (inp[14]) ? 4'b0001 : 4'b0000;
															assign node24351 = (inp[10]) ? node24353 : 4'b0001;
																assign node24353 = (inp[14]) ? 4'b0000 : 4'b0001;
														assign node24356 = (inp[14]) ? 4'b0000 : node24357;
															assign node24357 = (inp[12]) ? 4'b0001 : 4'b0000;
												assign node24361 = (inp[1]) ? node24373 : node24362;
													assign node24362 = (inp[13]) ? node24368 : node24363;
														assign node24363 = (inp[10]) ? node24365 : 4'b0001;
															assign node24365 = (inp[12]) ? 4'b0001 : 4'b0000;
														assign node24368 = (inp[10]) ? 4'b0000 : node24369;
															assign node24369 = (inp[12]) ? 4'b0000 : 4'b0001;
													assign node24373 = (inp[13]) ? 4'b0000 : node24374;
														assign node24374 = (inp[12]) ? 4'b0000 : node24375;
															assign node24375 = (inp[10]) ? 4'b0000 : 4'b1000;
										assign node24380 = (inp[13]) ? node24382 : 4'b0000;
											assign node24382 = (inp[14]) ? 4'b0000 : node24383;
												assign node24383 = (inp[11]) ? 4'b0000 : node24384;
													assign node24384 = (inp[4]) ? node24386 : 4'b0000;
														assign node24386 = (inp[10]) ? node24388 : 4'b0000;
															assign node24388 = (inp[1]) ? 4'b0000 : node24389;
																assign node24389 = (inp[12]) ? 4'b0000 : 4'b0001;

endmodule