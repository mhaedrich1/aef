module dtc_split33_bm61 (
	input  wire [12-1:0] inp,
	output wire [11-1:0] outp
);

	wire [11-1:0] node1;
	wire [11-1:0] node2;
	wire [11-1:0] node3;
	wire [11-1:0] node4;
	wire [11-1:0] node5;
	wire [11-1:0] node6;
	wire [11-1:0] node7;
	wire [11-1:0] node8;
	wire [11-1:0] node9;
	wire [11-1:0] node10;
	wire [11-1:0] node13;
	wire [11-1:0] node17;
	wire [11-1:0] node18;
	wire [11-1:0] node19;
	wire [11-1:0] node22;
	wire [11-1:0] node23;
	wire [11-1:0] node27;
	wire [11-1:0] node30;
	wire [11-1:0] node31;
	wire [11-1:0] node32;
	wire [11-1:0] node33;
	wire [11-1:0] node36;
	wire [11-1:0] node37;
	wire [11-1:0] node41;
	wire [11-1:0] node42;
	wire [11-1:0] node45;
	wire [11-1:0] node46;
	wire [11-1:0] node50;
	wire [11-1:0] node51;
	wire [11-1:0] node54;
	wire [11-1:0] node55;
	wire [11-1:0] node59;
	wire [11-1:0] node60;
	wire [11-1:0] node61;
	wire [11-1:0] node62;
	wire [11-1:0] node63;
	wire [11-1:0] node67;
	wire [11-1:0] node68;
	wire [11-1:0] node70;
	wire [11-1:0] node73;
	wire [11-1:0] node76;
	wire [11-1:0] node77;
	wire [11-1:0] node79;
	wire [11-1:0] node82;
	wire [11-1:0] node84;
	wire [11-1:0] node87;
	wire [11-1:0] node88;
	wire [11-1:0] node89;
	wire [11-1:0] node91;
	wire [11-1:0] node92;
	wire [11-1:0] node95;
	wire [11-1:0] node98;
	wire [11-1:0] node99;
	wire [11-1:0] node103;
	wire [11-1:0] node104;
	wire [11-1:0] node105;
	wire [11-1:0] node108;
	wire [11-1:0] node112;
	wire [11-1:0] node113;
	wire [11-1:0] node114;
	wire [11-1:0] node115;
	wire [11-1:0] node117;
	wire [11-1:0] node119;
	wire [11-1:0] node120;
	wire [11-1:0] node124;
	wire [11-1:0] node125;
	wire [11-1:0] node128;
	wire [11-1:0] node129;
	wire [11-1:0] node131;
	wire [11-1:0] node134;
	wire [11-1:0] node136;
	wire [11-1:0] node139;
	wire [11-1:0] node140;
	wire [11-1:0] node141;
	wire [11-1:0] node144;
	wire [11-1:0] node147;
	wire [11-1:0] node148;
	wire [11-1:0] node152;
	wire [11-1:0] node153;
	wire [11-1:0] node154;
	wire [11-1:0] node155;
	wire [11-1:0] node156;
	wire [11-1:0] node159;
	wire [11-1:0] node162;
	wire [11-1:0] node165;
	wire [11-1:0] node167;
	wire [11-1:0] node170;
	wire [11-1:0] node171;
	wire [11-1:0] node172;
	wire [11-1:0] node174;
	wire [11-1:0] node177;
	wire [11-1:0] node180;
	wire [11-1:0] node181;
	wire [11-1:0] node184;
	wire [11-1:0] node186;
	wire [11-1:0] node188;
	wire [11-1:0] node191;
	wire [11-1:0] node192;
	wire [11-1:0] node193;
	wire [11-1:0] node194;
	wire [11-1:0] node195;
	wire [11-1:0] node196;
	wire [11-1:0] node197;
	wire [11-1:0] node200;
	wire [11-1:0] node204;
	wire [11-1:0] node205;
	wire [11-1:0] node207;
	wire [11-1:0] node208;
	wire [11-1:0] node212;
	wire [11-1:0] node215;
	wire [11-1:0] node216;
	wire [11-1:0] node217;
	wire [11-1:0] node218;
	wire [11-1:0] node221;
	wire [11-1:0] node224;
	wire [11-1:0] node226;
	wire [11-1:0] node227;
	wire [11-1:0] node231;
	wire [11-1:0] node232;
	wire [11-1:0] node233;
	wire [11-1:0] node236;
	wire [11-1:0] node240;
	wire [11-1:0] node241;
	wire [11-1:0] node242;
	wire [11-1:0] node243;
	wire [11-1:0] node244;
	wire [11-1:0] node245;
	wire [11-1:0] node249;
	wire [11-1:0] node252;
	wire [11-1:0] node254;
	wire [11-1:0] node257;
	wire [11-1:0] node258;
	wire [11-1:0] node260;
	wire [11-1:0] node263;
	wire [11-1:0] node264;
	wire [11-1:0] node268;
	wire [11-1:0] node270;
	wire [11-1:0] node271;
	wire [11-1:0] node272;
	wire [11-1:0] node274;
	wire [11-1:0] node278;
	wire [11-1:0] node280;
	wire [11-1:0] node281;
	wire [11-1:0] node284;
	wire [11-1:0] node287;
	wire [11-1:0] node288;
	wire [11-1:0] node289;
	wire [11-1:0] node290;
	wire [11-1:0] node292;
	wire [11-1:0] node294;
	wire [11-1:0] node297;
	wire [11-1:0] node298;
	wire [11-1:0] node301;
	wire [11-1:0] node302;
	wire [11-1:0] node303;
	wire [11-1:0] node307;
	wire [11-1:0] node310;
	wire [11-1:0] node311;
	wire [11-1:0] node312;
	wire [11-1:0] node315;
	wire [11-1:0] node318;
	wire [11-1:0] node319;
	wire [11-1:0] node320;
	wire [11-1:0] node324;
	wire [11-1:0] node327;
	wire [11-1:0] node328;
	wire [11-1:0] node329;
	wire [11-1:0] node330;
	wire [11-1:0] node333;
	wire [11-1:0] node334;
	wire [11-1:0] node336;
	wire [11-1:0] node340;
	wire [11-1:0] node341;
	wire [11-1:0] node344;
	wire [11-1:0] node346;
	wire [11-1:0] node347;
	wire [11-1:0] node351;
	wire [11-1:0] node352;
	wire [11-1:0] node353;
	wire [11-1:0] node354;
	wire [11-1:0] node358;
	wire [11-1:0] node360;
	wire [11-1:0] node363;
	wire [11-1:0] node364;
	wire [11-1:0] node365;
	wire [11-1:0] node368;
	wire [11-1:0] node372;
	wire [11-1:0] node373;
	wire [11-1:0] node374;
	wire [11-1:0] node375;
	wire [11-1:0] node376;
	wire [11-1:0] node377;
	wire [11-1:0] node380;
	wire [11-1:0] node381;
	wire [11-1:0] node385;
	wire [11-1:0] node386;
	wire [11-1:0] node387;
	wire [11-1:0] node390;
	wire [11-1:0] node391;
	wire [11-1:0] node395;
	wire [11-1:0] node396;
	wire [11-1:0] node399;
	wire [11-1:0] node402;
	wire [11-1:0] node403;
	wire [11-1:0] node404;
	wire [11-1:0] node405;
	wire [11-1:0] node408;
	wire [11-1:0] node409;
	wire [11-1:0] node413;
	wire [11-1:0] node414;
	wire [11-1:0] node415;
	wire [11-1:0] node417;
	wire [11-1:0] node421;
	wire [11-1:0] node424;
	wire [11-1:0] node425;
	wire [11-1:0] node428;
	wire [11-1:0] node430;
	wire [11-1:0] node432;
	wire [11-1:0] node433;
	wire [11-1:0] node437;
	wire [11-1:0] node438;
	wire [11-1:0] node439;
	wire [11-1:0] node440;
	wire [11-1:0] node441;
	wire [11-1:0] node444;
	wire [11-1:0] node445;
	wire [11-1:0] node449;
	wire [11-1:0] node450;
	wire [11-1:0] node453;
	wire [11-1:0] node456;
	wire [11-1:0] node457;
	wire [11-1:0] node458;
	wire [11-1:0] node459;
	wire [11-1:0] node461;
	wire [11-1:0] node465;
	wire [11-1:0] node467;
	wire [11-1:0] node470;
	wire [11-1:0] node471;
	wire [11-1:0] node472;
	wire [11-1:0] node477;
	wire [11-1:0] node478;
	wire [11-1:0] node479;
	wire [11-1:0] node480;
	wire [11-1:0] node483;
	wire [11-1:0] node486;
	wire [11-1:0] node487;
	wire [11-1:0] node488;
	wire [11-1:0] node492;
	wire [11-1:0] node493;
	wire [11-1:0] node495;
	wire [11-1:0] node498;
	wire [11-1:0] node500;
	wire [11-1:0] node503;
	wire [11-1:0] node504;
	wire [11-1:0] node505;
	wire [11-1:0] node508;
	wire [11-1:0] node509;
	wire [11-1:0] node512;
	wire [11-1:0] node515;
	wire [11-1:0] node516;
	wire [11-1:0] node518;
	wire [11-1:0] node520;
	wire [11-1:0] node523;
	wire [11-1:0] node525;
	wire [11-1:0] node528;
	wire [11-1:0] node529;
	wire [11-1:0] node530;
	wire [11-1:0] node531;
	wire [11-1:0] node532;
	wire [11-1:0] node534;
	wire [11-1:0] node536;
	wire [11-1:0] node538;
	wire [11-1:0] node541;
	wire [11-1:0] node542;
	wire [11-1:0] node544;
	wire [11-1:0] node547;
	wire [11-1:0] node549;
	wire [11-1:0] node552;
	wire [11-1:0] node553;
	wire [11-1:0] node554;
	wire [11-1:0] node556;
	wire [11-1:0] node559;
	wire [11-1:0] node560;
	wire [11-1:0] node561;
	wire [11-1:0] node565;
	wire [11-1:0] node568;
	wire [11-1:0] node569;
	wire [11-1:0] node572;
	wire [11-1:0] node575;
	wire [11-1:0] node576;
	wire [11-1:0] node577;
	wire [11-1:0] node579;
	wire [11-1:0] node582;
	wire [11-1:0] node583;
	wire [11-1:0] node586;
	wire [11-1:0] node589;
	wire [11-1:0] node590;
	wire [11-1:0] node593;
	wire [11-1:0] node594;
	wire [11-1:0] node597;
	wire [11-1:0] node598;
	wire [11-1:0] node600;
	wire [11-1:0] node603;
	wire [11-1:0] node606;
	wire [11-1:0] node607;
	wire [11-1:0] node608;
	wire [11-1:0] node609;
	wire [11-1:0] node610;
	wire [11-1:0] node613;
	wire [11-1:0] node616;
	wire [11-1:0] node617;
	wire [11-1:0] node620;
	wire [11-1:0] node622;
	wire [11-1:0] node625;
	wire [11-1:0] node626;
	wire [11-1:0] node627;
	wire [11-1:0] node628;
	wire [11-1:0] node632;
	wire [11-1:0] node633;
	wire [11-1:0] node636;
	wire [11-1:0] node637;
	wire [11-1:0] node641;
	wire [11-1:0] node642;
	wire [11-1:0] node643;
	wire [11-1:0] node647;
	wire [11-1:0] node648;
	wire [11-1:0] node650;
	wire [11-1:0] node654;
	wire [11-1:0] node655;
	wire [11-1:0] node656;
	wire [11-1:0] node657;
	wire [11-1:0] node660;
	wire [11-1:0] node663;
	wire [11-1:0] node664;
	wire [11-1:0] node665;
	wire [11-1:0] node669;
	wire [11-1:0] node671;
	wire [11-1:0] node673;
	wire [11-1:0] node676;
	wire [11-1:0] node677;
	wire [11-1:0] node678;
	wire [11-1:0] node680;
	wire [11-1:0] node683;
	wire [11-1:0] node686;
	wire [11-1:0] node687;
	wire [11-1:0] node688;
	wire [11-1:0] node691;
	wire [11-1:0] node694;
	wire [11-1:0] node695;
	wire [11-1:0] node699;
	wire [11-1:0] node700;
	wire [11-1:0] node701;
	wire [11-1:0] node702;
	wire [11-1:0] node703;
	wire [11-1:0] node704;
	wire [11-1:0] node705;
	wire [11-1:0] node706;
	wire [11-1:0] node710;
	wire [11-1:0] node711;
	wire [11-1:0] node714;
	wire [11-1:0] node717;
	wire [11-1:0] node718;
	wire [11-1:0] node719;
	wire [11-1:0] node720;
	wire [11-1:0] node724;
	wire [11-1:0] node726;
	wire [11-1:0] node729;
	wire [11-1:0] node730;
	wire [11-1:0] node732;
	wire [11-1:0] node735;
	wire [11-1:0] node738;
	wire [11-1:0] node739;
	wire [11-1:0] node740;
	wire [11-1:0] node741;
	wire [11-1:0] node744;
	wire [11-1:0] node745;
	wire [11-1:0] node749;
	wire [11-1:0] node750;
	wire [11-1:0] node752;
	wire [11-1:0] node755;
	wire [11-1:0] node758;
	wire [11-1:0] node759;
	wire [11-1:0] node760;
	wire [11-1:0] node763;
	wire [11-1:0] node764;
	wire [11-1:0] node767;
	wire [11-1:0] node770;
	wire [11-1:0] node771;
	wire [11-1:0] node774;
	wire [11-1:0] node776;
	wire [11-1:0] node779;
	wire [11-1:0] node780;
	wire [11-1:0] node781;
	wire [11-1:0] node782;
	wire [11-1:0] node783;
	wire [11-1:0] node784;
	wire [11-1:0] node785;
	wire [11-1:0] node788;
	wire [11-1:0] node792;
	wire [11-1:0] node793;
	wire [11-1:0] node796;
	wire [11-1:0] node798;
	wire [11-1:0] node801;
	wire [11-1:0] node802;
	wire [11-1:0] node804;
	wire [11-1:0] node807;
	wire [11-1:0] node808;
	wire [11-1:0] node812;
	wire [11-1:0] node813;
	wire [11-1:0] node814;
	wire [11-1:0] node816;
	wire [11-1:0] node819;
	wire [11-1:0] node821;
	wire [11-1:0] node822;
	wire [11-1:0] node826;
	wire [11-1:0] node827;
	wire [11-1:0] node828;
	wire [11-1:0] node831;
	wire [11-1:0] node834;
	wire [11-1:0] node837;
	wire [11-1:0] node838;
	wire [11-1:0] node839;
	wire [11-1:0] node840;
	wire [11-1:0] node843;
	wire [11-1:0] node846;
	wire [11-1:0] node849;
	wire [11-1:0] node850;
	wire [11-1:0] node851;
	wire [11-1:0] node852;
	wire [11-1:0] node857;
	wire [11-1:0] node858;
	wire [11-1:0] node859;
	wire [11-1:0] node864;
	wire [11-1:0] node865;
	wire [11-1:0] node866;
	wire [11-1:0] node867;
	wire [11-1:0] node868;
	wire [11-1:0] node869;
	wire [11-1:0] node870;
	wire [11-1:0] node874;
	wire [11-1:0] node876;
	wire [11-1:0] node877;
	wire [11-1:0] node880;
	wire [11-1:0] node883;
	wire [11-1:0] node884;
	wire [11-1:0] node885;
	wire [11-1:0] node889;
	wire [11-1:0] node890;
	wire [11-1:0] node892;
	wire [11-1:0] node896;
	wire [11-1:0] node897;
	wire [11-1:0] node898;
	wire [11-1:0] node899;
	wire [11-1:0] node903;
	wire [11-1:0] node904;
	wire [11-1:0] node908;
	wire [11-1:0] node909;
	wire [11-1:0] node910;
	wire [11-1:0] node914;
	wire [11-1:0] node916;
	wire [11-1:0] node919;
	wire [11-1:0] node920;
	wire [11-1:0] node921;
	wire [11-1:0] node922;
	wire [11-1:0] node923;
	wire [11-1:0] node926;
	wire [11-1:0] node927;
	wire [11-1:0] node931;
	wire [11-1:0] node933;
	wire [11-1:0] node936;
	wire [11-1:0] node937;
	wire [11-1:0] node940;
	wire [11-1:0] node942;
	wire [11-1:0] node945;
	wire [11-1:0] node946;
	wire [11-1:0] node947;
	wire [11-1:0] node950;
	wire [11-1:0] node951;
	wire [11-1:0] node953;
	wire [11-1:0] node957;
	wire [11-1:0] node959;
	wire [11-1:0] node960;
	wire [11-1:0] node964;
	wire [11-1:0] node965;
	wire [11-1:0] node966;
	wire [11-1:0] node967;
	wire [11-1:0] node968;
	wire [11-1:0] node969;
	wire [11-1:0] node973;
	wire [11-1:0] node976;
	wire [11-1:0] node978;
	wire [11-1:0] node979;
	wire [11-1:0] node983;
	wire [11-1:0] node984;
	wire [11-1:0] node985;
	wire [11-1:0] node986;
	wire [11-1:0] node989;
	wire [11-1:0] node990;
	wire [11-1:0] node994;
	wire [11-1:0] node995;
	wire [11-1:0] node997;
	wire [11-1:0] node1000;
	wire [11-1:0] node1001;
	wire [11-1:0] node1005;
	wire [11-1:0] node1006;
	wire [11-1:0] node1009;
	wire [11-1:0] node1010;
	wire [11-1:0] node1014;
	wire [11-1:0] node1015;
	wire [11-1:0] node1016;
	wire [11-1:0] node1019;
	wire [11-1:0] node1020;
	wire [11-1:0] node1021;
	wire [11-1:0] node1025;
	wire [11-1:0] node1026;
	wire [11-1:0] node1029;
	wire [11-1:0] node1032;
	wire [11-1:0] node1033;
	wire [11-1:0] node1034;
	wire [11-1:0] node1035;
	wire [11-1:0] node1039;
	wire [11-1:0] node1040;
	wire [11-1:0] node1044;
	wire [11-1:0] node1045;
	wire [11-1:0] node1048;
	wire [11-1:0] node1049;
	wire [11-1:0] node1050;
	wire [11-1:0] node1055;
	wire [11-1:0] node1056;
	wire [11-1:0] node1057;
	wire [11-1:0] node1058;
	wire [11-1:0] node1059;
	wire [11-1:0] node1060;
	wire [11-1:0] node1061;
	wire [11-1:0] node1064;
	wire [11-1:0] node1067;
	wire [11-1:0] node1068;
	wire [11-1:0] node1069;
	wire [11-1:0] node1072;
	wire [11-1:0] node1075;
	wire [11-1:0] node1076;
	wire [11-1:0] node1080;
	wire [11-1:0] node1081;
	wire [11-1:0] node1083;
	wire [11-1:0] node1084;
	wire [11-1:0] node1086;
	wire [11-1:0] node1089;
	wire [11-1:0] node1092;
	wire [11-1:0] node1093;
	wire [11-1:0] node1095;
	wire [11-1:0] node1097;
	wire [11-1:0] node1101;
	wire [11-1:0] node1102;
	wire [11-1:0] node1103;
	wire [11-1:0] node1104;
	wire [11-1:0] node1106;
	wire [11-1:0] node1109;
	wire [11-1:0] node1110;
	wire [11-1:0] node1114;
	wire [11-1:0] node1116;
	wire [11-1:0] node1119;
	wire [11-1:0] node1120;
	wire [11-1:0] node1121;
	wire [11-1:0] node1123;
	wire [11-1:0] node1126;
	wire [11-1:0] node1127;
	wire [11-1:0] node1130;
	wire [11-1:0] node1133;
	wire [11-1:0] node1135;
	wire [11-1:0] node1138;
	wire [11-1:0] node1139;
	wire [11-1:0] node1140;
	wire [11-1:0] node1141;
	wire [11-1:0] node1142;
	wire [11-1:0] node1145;
	wire [11-1:0] node1147;
	wire [11-1:0] node1150;
	wire [11-1:0] node1151;
	wire [11-1:0] node1153;
	wire [11-1:0] node1156;
	wire [11-1:0] node1157;
	wire [11-1:0] node1160;
	wire [11-1:0] node1163;
	wire [11-1:0] node1164;
	wire [11-1:0] node1165;
	wire [11-1:0] node1168;
	wire [11-1:0] node1171;
	wire [11-1:0] node1174;
	wire [11-1:0] node1175;
	wire [11-1:0] node1176;
	wire [11-1:0] node1177;
	wire [11-1:0] node1180;
	wire [11-1:0] node1182;
	wire [11-1:0] node1185;
	wire [11-1:0] node1187;
	wire [11-1:0] node1189;
	wire [11-1:0] node1192;
	wire [11-1:0] node1193;
	wire [11-1:0] node1194;
	wire [11-1:0] node1196;
	wire [11-1:0] node1199;
	wire [11-1:0] node1200;
	wire [11-1:0] node1204;
	wire [11-1:0] node1205;
	wire [11-1:0] node1208;
	wire [11-1:0] node1211;
	wire [11-1:0] node1212;
	wire [11-1:0] node1213;
	wire [11-1:0] node1214;
	wire [11-1:0] node1215;
	wire [11-1:0] node1216;
	wire [11-1:0] node1217;
	wire [11-1:0] node1219;
	wire [11-1:0] node1222;
	wire [11-1:0] node1224;
	wire [11-1:0] node1227;
	wire [11-1:0] node1229;
	wire [11-1:0] node1232;
	wire [11-1:0] node1233;
	wire [11-1:0] node1234;
	wire [11-1:0] node1237;
	wire [11-1:0] node1241;
	wire [11-1:0] node1242;
	wire [11-1:0] node1243;
	wire [11-1:0] node1244;
	wire [11-1:0] node1247;
	wire [11-1:0] node1249;
	wire [11-1:0] node1252;
	wire [11-1:0] node1254;
	wire [11-1:0] node1257;
	wire [11-1:0] node1259;
	wire [11-1:0] node1260;
	wire [11-1:0] node1263;
	wire [11-1:0] node1266;
	wire [11-1:0] node1267;
	wire [11-1:0] node1268;
	wire [11-1:0] node1269;
	wire [11-1:0] node1270;
	wire [11-1:0] node1271;
	wire [11-1:0] node1276;
	wire [11-1:0] node1277;
	wire [11-1:0] node1280;
	wire [11-1:0] node1283;
	wire [11-1:0] node1285;
	wire [11-1:0] node1286;
	wire [11-1:0] node1289;
	wire [11-1:0] node1292;
	wire [11-1:0] node1293;
	wire [11-1:0] node1294;
	wire [11-1:0] node1295;
	wire [11-1:0] node1298;
	wire [11-1:0] node1301;
	wire [11-1:0] node1303;
	wire [11-1:0] node1306;
	wire [11-1:0] node1307;
	wire [11-1:0] node1308;
	wire [11-1:0] node1313;
	wire [11-1:0] node1314;
	wire [11-1:0] node1315;
	wire [11-1:0] node1316;
	wire [11-1:0] node1317;
	wire [11-1:0] node1320;
	wire [11-1:0] node1323;
	wire [11-1:0] node1326;
	wire [11-1:0] node1327;
	wire [11-1:0] node1328;
	wire [11-1:0] node1329;
	wire [11-1:0] node1334;
	wire [11-1:0] node1337;
	wire [11-1:0] node1338;
	wire [11-1:0] node1339;
	wire [11-1:0] node1340;
	wire [11-1:0] node1343;
	wire [11-1:0] node1346;
	wire [11-1:0] node1347;
	wire [11-1:0] node1351;
	wire [11-1:0] node1352;
	wire [11-1:0] node1353;
	wire [11-1:0] node1356;
	wire [11-1:0] node1357;
	wire [11-1:0] node1358;
	wire [11-1:0] node1361;
	wire [11-1:0] node1365;
	wire [11-1:0] node1368;
	wire [11-1:0] node1369;
	wire [11-1:0] node1370;
	wire [11-1:0] node1371;
	wire [11-1:0] node1372;
	wire [11-1:0] node1373;
	wire [11-1:0] node1374;
	wire [11-1:0] node1375;
	wire [11-1:0] node1376;
	wire [11-1:0] node1377;
	wire [11-1:0] node1380;
	wire [11-1:0] node1383;
	wire [11-1:0] node1385;
	wire [11-1:0] node1388;
	wire [11-1:0] node1389;
	wire [11-1:0] node1392;
	wire [11-1:0] node1395;
	wire [11-1:0] node1396;
	wire [11-1:0] node1398;
	wire [11-1:0] node1399;
	wire [11-1:0] node1402;
	wire [11-1:0] node1405;
	wire [11-1:0] node1406;
	wire [11-1:0] node1407;
	wire [11-1:0] node1411;
	wire [11-1:0] node1414;
	wire [11-1:0] node1415;
	wire [11-1:0] node1416;
	wire [11-1:0] node1417;
	wire [11-1:0] node1418;
	wire [11-1:0] node1421;
	wire [11-1:0] node1424;
	wire [11-1:0] node1426;
	wire [11-1:0] node1429;
	wire [11-1:0] node1430;
	wire [11-1:0] node1431;
	wire [11-1:0] node1435;
	wire [11-1:0] node1436;
	wire [11-1:0] node1440;
	wire [11-1:0] node1441;
	wire [11-1:0] node1442;
	wire [11-1:0] node1445;
	wire [11-1:0] node1448;
	wire [11-1:0] node1449;
	wire [11-1:0] node1453;
	wire [11-1:0] node1454;
	wire [11-1:0] node1455;
	wire [11-1:0] node1456;
	wire [11-1:0] node1457;
	wire [11-1:0] node1459;
	wire [11-1:0] node1462;
	wire [11-1:0] node1463;
	wire [11-1:0] node1466;
	wire [11-1:0] node1469;
	wire [11-1:0] node1470;
	wire [11-1:0] node1472;
	wire [11-1:0] node1476;
	wire [11-1:0] node1477;
	wire [11-1:0] node1478;
	wire [11-1:0] node1479;
	wire [11-1:0] node1484;
	wire [11-1:0] node1485;
	wire [11-1:0] node1488;
	wire [11-1:0] node1491;
	wire [11-1:0] node1492;
	wire [11-1:0] node1493;
	wire [11-1:0] node1496;
	wire [11-1:0] node1497;
	wire [11-1:0] node1498;
	wire [11-1:0] node1500;
	wire [11-1:0] node1503;
	wire [11-1:0] node1506;
	wire [11-1:0] node1507;
	wire [11-1:0] node1510;
	wire [11-1:0] node1513;
	wire [11-1:0] node1514;
	wire [11-1:0] node1515;
	wire [11-1:0] node1516;
	wire [11-1:0] node1519;
	wire [11-1:0] node1521;
	wire [11-1:0] node1524;
	wire [11-1:0] node1525;
	wire [11-1:0] node1528;
	wire [11-1:0] node1530;
	wire [11-1:0] node1533;
	wire [11-1:0] node1535;
	wire [11-1:0] node1536;
	wire [11-1:0] node1540;
	wire [11-1:0] node1541;
	wire [11-1:0] node1542;
	wire [11-1:0] node1543;
	wire [11-1:0] node1544;
	wire [11-1:0] node1545;
	wire [11-1:0] node1546;
	wire [11-1:0] node1550;
	wire [11-1:0] node1553;
	wire [11-1:0] node1554;
	wire [11-1:0] node1557;
	wire [11-1:0] node1560;
	wire [11-1:0] node1561;
	wire [11-1:0] node1562;
	wire [11-1:0] node1565;
	wire [11-1:0] node1566;
	wire [11-1:0] node1569;
	wire [11-1:0] node1573;
	wire [11-1:0] node1574;
	wire [11-1:0] node1575;
	wire [11-1:0] node1576;
	wire [11-1:0] node1577;
	wire [11-1:0] node1580;
	wire [11-1:0] node1583;
	wire [11-1:0] node1585;
	wire [11-1:0] node1588;
	wire [11-1:0] node1590;
	wire [11-1:0] node1591;
	wire [11-1:0] node1594;
	wire [11-1:0] node1597;
	wire [11-1:0] node1598;
	wire [11-1:0] node1599;
	wire [11-1:0] node1602;
	wire [11-1:0] node1605;
	wire [11-1:0] node1607;
	wire [11-1:0] node1610;
	wire [11-1:0] node1611;
	wire [11-1:0] node1612;
	wire [11-1:0] node1613;
	wire [11-1:0] node1614;
	wire [11-1:0] node1617;
	wire [11-1:0] node1618;
	wire [11-1:0] node1622;
	wire [11-1:0] node1624;
	wire [11-1:0] node1626;
	wire [11-1:0] node1629;
	wire [11-1:0] node1630;
	wire [11-1:0] node1631;
	wire [11-1:0] node1632;
	wire [11-1:0] node1633;
	wire [11-1:0] node1639;
	wire [11-1:0] node1642;
	wire [11-1:0] node1643;
	wire [11-1:0] node1644;
	wire [11-1:0] node1645;
	wire [11-1:0] node1646;
	wire [11-1:0] node1650;
	wire [11-1:0] node1651;
	wire [11-1:0] node1652;
	wire [11-1:0] node1657;
	wire [11-1:0] node1659;
	wire [11-1:0] node1660;
	wire [11-1:0] node1662;
	wire [11-1:0] node1666;
	wire [11-1:0] node1667;
	wire [11-1:0] node1668;
	wire [11-1:0] node1672;
	wire [11-1:0] node1673;
	wire [11-1:0] node1676;
	wire [11-1:0] node1679;
	wire [11-1:0] node1680;
	wire [11-1:0] node1681;
	wire [11-1:0] node1682;
	wire [11-1:0] node1683;
	wire [11-1:0] node1684;
	wire [11-1:0] node1685;
	wire [11-1:0] node1688;
	wire [11-1:0] node1691;
	wire [11-1:0] node1692;
	wire [11-1:0] node1694;
	wire [11-1:0] node1695;
	wire [11-1:0] node1698;
	wire [11-1:0] node1702;
	wire [11-1:0] node1704;
	wire [11-1:0] node1705;
	wire [11-1:0] node1708;
	wire [11-1:0] node1709;
	wire [11-1:0] node1711;
	wire [11-1:0] node1715;
	wire [11-1:0] node1716;
	wire [11-1:0] node1717;
	wire [11-1:0] node1718;
	wire [11-1:0] node1720;
	wire [11-1:0] node1723;
	wire [11-1:0] node1724;
	wire [11-1:0] node1728;
	wire [11-1:0] node1729;
	wire [11-1:0] node1732;
	wire [11-1:0] node1733;
	wire [11-1:0] node1737;
	wire [11-1:0] node1738;
	wire [11-1:0] node1739;
	wire [11-1:0] node1742;
	wire [11-1:0] node1744;
	wire [11-1:0] node1747;
	wire [11-1:0] node1750;
	wire [11-1:0] node1751;
	wire [11-1:0] node1752;
	wire [11-1:0] node1753;
	wire [11-1:0] node1754;
	wire [11-1:0] node1755;
	wire [11-1:0] node1759;
	wire [11-1:0] node1761;
	wire [11-1:0] node1764;
	wire [11-1:0] node1765;
	wire [11-1:0] node1766;
	wire [11-1:0] node1768;
	wire [11-1:0] node1772;
	wire [11-1:0] node1775;
	wire [11-1:0] node1776;
	wire [11-1:0] node1777;
	wire [11-1:0] node1780;
	wire [11-1:0] node1783;
	wire [11-1:0] node1784;
	wire [11-1:0] node1787;
	wire [11-1:0] node1789;
	wire [11-1:0] node1792;
	wire [11-1:0] node1793;
	wire [11-1:0] node1794;
	wire [11-1:0] node1797;
	wire [11-1:0] node1798;
	wire [11-1:0] node1801;
	wire [11-1:0] node1804;
	wire [11-1:0] node1806;
	wire [11-1:0] node1808;
	wire [11-1:0] node1810;
	wire [11-1:0] node1813;
	wire [11-1:0] node1814;
	wire [11-1:0] node1815;
	wire [11-1:0] node1816;
	wire [11-1:0] node1817;
	wire [11-1:0] node1818;
	wire [11-1:0] node1819;
	wire [11-1:0] node1822;
	wire [11-1:0] node1825;
	wire [11-1:0] node1828;
	wire [11-1:0] node1830;
	wire [11-1:0] node1832;
	wire [11-1:0] node1835;
	wire [11-1:0] node1836;
	wire [11-1:0] node1839;
	wire [11-1:0] node1840;
	wire [11-1:0] node1841;
	wire [11-1:0] node1843;
	wire [11-1:0] node1848;
	wire [11-1:0] node1849;
	wire [11-1:0] node1850;
	wire [11-1:0] node1853;
	wire [11-1:0] node1854;
	wire [11-1:0] node1857;
	wire [11-1:0] node1860;
	wire [11-1:0] node1861;
	wire [11-1:0] node1862;
	wire [11-1:0] node1865;
	wire [11-1:0] node1867;
	wire [11-1:0] node1870;
	wire [11-1:0] node1872;
	wire [11-1:0] node1875;
	wire [11-1:0] node1876;
	wire [11-1:0] node1877;
	wire [11-1:0] node1878;
	wire [11-1:0] node1879;
	wire [11-1:0] node1880;
	wire [11-1:0] node1883;
	wire [11-1:0] node1885;
	wire [11-1:0] node1888;
	wire [11-1:0] node1889;
	wire [11-1:0] node1892;
	wire [11-1:0] node1895;
	wire [11-1:0] node1896;
	wire [11-1:0] node1897;
	wire [11-1:0] node1901;
	wire [11-1:0] node1902;
	wire [11-1:0] node1904;
	wire [11-1:0] node1907;
	wire [11-1:0] node1910;
	wire [11-1:0] node1911;
	wire [11-1:0] node1912;
	wire [11-1:0] node1913;
	wire [11-1:0] node1914;
	wire [11-1:0] node1917;
	wire [11-1:0] node1920;
	wire [11-1:0] node1922;
	wire [11-1:0] node1926;
	wire [11-1:0] node1927;
	wire [11-1:0] node1928;
	wire [11-1:0] node1932;
	wire [11-1:0] node1933;
	wire [11-1:0] node1936;
	wire [11-1:0] node1939;
	wire [11-1:0] node1940;
	wire [11-1:0] node1941;
	wire [11-1:0] node1942;
	wire [11-1:0] node1943;
	wire [11-1:0] node1946;
	wire [11-1:0] node1949;
	wire [11-1:0] node1951;
	wire [11-1:0] node1954;
	wire [11-1:0] node1955;
	wire [11-1:0] node1958;
	wire [11-1:0] node1959;
	wire [11-1:0] node1962;
	wire [11-1:0] node1963;
	wire [11-1:0] node1967;
	wire [11-1:0] node1968;
	wire [11-1:0] node1970;
	wire [11-1:0] node1973;
	wire [11-1:0] node1974;
	wire [11-1:0] node1977;
	wire [11-1:0] node1978;
	wire [11-1:0] node1982;
	wire [11-1:0] node1983;
	wire [11-1:0] node1984;
	wire [11-1:0] node1985;
	wire [11-1:0] node1986;
	wire [11-1:0] node1987;
	wire [11-1:0] node1988;
	wire [11-1:0] node1989;
	wire [11-1:0] node1990;
	wire [11-1:0] node1993;
	wire [11-1:0] node1996;
	wire [11-1:0] node1999;
	wire [11-1:0] node2000;
	wire [11-1:0] node2003;
	wire [11-1:0] node2005;
	wire [11-1:0] node2008;
	wire [11-1:0] node2009;
	wire [11-1:0] node2010;
	wire [11-1:0] node2012;
	wire [11-1:0] node2015;
	wire [11-1:0] node2018;
	wire [11-1:0] node2019;
	wire [11-1:0] node2023;
	wire [11-1:0] node2024;
	wire [11-1:0] node2025;
	wire [11-1:0] node2026;
	wire [11-1:0] node2028;
	wire [11-1:0] node2032;
	wire [11-1:0] node2033;
	wire [11-1:0] node2035;
	wire [11-1:0] node2038;
	wire [11-1:0] node2039;
	wire [11-1:0] node2043;
	wire [11-1:0] node2044;
	wire [11-1:0] node2045;
	wire [11-1:0] node2046;
	wire [11-1:0] node2050;
	wire [11-1:0] node2053;
	wire [11-1:0] node2054;
	wire [11-1:0] node2057;
	wire [11-1:0] node2060;
	wire [11-1:0] node2061;
	wire [11-1:0] node2062;
	wire [11-1:0] node2063;
	wire [11-1:0] node2064;
	wire [11-1:0] node2068;
	wire [11-1:0] node2069;
	wire [11-1:0] node2072;
	wire [11-1:0] node2075;
	wire [11-1:0] node2076;
	wire [11-1:0] node2077;
	wire [11-1:0] node2078;
	wire [11-1:0] node2082;
	wire [11-1:0] node2083;
	wire [11-1:0] node2086;
	wire [11-1:0] node2089;
	wire [11-1:0] node2091;
	wire [11-1:0] node2093;
	wire [11-1:0] node2096;
	wire [11-1:0] node2097;
	wire [11-1:0] node2098;
	wire [11-1:0] node2099;
	wire [11-1:0] node2102;
	wire [11-1:0] node2103;
	wire [11-1:0] node2106;
	wire [11-1:0] node2109;
	wire [11-1:0] node2110;
	wire [11-1:0] node2111;
	wire [11-1:0] node2115;
	wire [11-1:0] node2116;
	wire [11-1:0] node2118;
	wire [11-1:0] node2121;
	wire [11-1:0] node2123;
	wire [11-1:0] node2126;
	wire [11-1:0] node2127;
	wire [11-1:0] node2128;
	wire [11-1:0] node2131;
	wire [11-1:0] node2133;
	wire [11-1:0] node2136;
	wire [11-1:0] node2138;
	wire [11-1:0] node2141;
	wire [11-1:0] node2142;
	wire [11-1:0] node2143;
	wire [11-1:0] node2144;
	wire [11-1:0] node2145;
	wire [11-1:0] node2146;
	wire [11-1:0] node2147;
	wire [11-1:0] node2150;
	wire [11-1:0] node2153;
	wire [11-1:0] node2156;
	wire [11-1:0] node2157;
	wire [11-1:0] node2158;
	wire [11-1:0] node2161;
	wire [11-1:0] node2164;
	wire [11-1:0] node2167;
	wire [11-1:0] node2168;
	wire [11-1:0] node2169;
	wire [11-1:0] node2170;
	wire [11-1:0] node2174;
	wire [11-1:0] node2177;
	wire [11-1:0] node2178;
	wire [11-1:0] node2179;
	wire [11-1:0] node2182;
	wire [11-1:0] node2185;
	wire [11-1:0] node2188;
	wire [11-1:0] node2189;
	wire [11-1:0] node2190;
	wire [11-1:0] node2191;
	wire [11-1:0] node2192;
	wire [11-1:0] node2194;
	wire [11-1:0] node2198;
	wire [11-1:0] node2199;
	wire [11-1:0] node2200;
	wire [11-1:0] node2204;
	wire [11-1:0] node2207;
	wire [11-1:0] node2209;
	wire [11-1:0] node2212;
	wire [11-1:0] node2213;
	wire [11-1:0] node2214;
	wire [11-1:0] node2217;
	wire [11-1:0] node2218;
	wire [11-1:0] node2221;
	wire [11-1:0] node2224;
	wire [11-1:0] node2225;
	wire [11-1:0] node2226;
	wire [11-1:0] node2227;
	wire [11-1:0] node2231;
	wire [11-1:0] node2234;
	wire [11-1:0] node2235;
	wire [11-1:0] node2239;
	wire [11-1:0] node2240;
	wire [11-1:0] node2241;
	wire [11-1:0] node2242;
	wire [11-1:0] node2243;
	wire [11-1:0] node2244;
	wire [11-1:0] node2248;
	wire [11-1:0] node2249;
	wire [11-1:0] node2252;
	wire [11-1:0] node2253;
	wire [11-1:0] node2256;
	wire [11-1:0] node2259;
	wire [11-1:0] node2260;
	wire [11-1:0] node2263;
	wire [11-1:0] node2264;
	wire [11-1:0] node2268;
	wire [11-1:0] node2269;
	wire [11-1:0] node2270;
	wire [11-1:0] node2273;
	wire [11-1:0] node2275;
	wire [11-1:0] node2277;
	wire [11-1:0] node2280;
	wire [11-1:0] node2281;
	wire [11-1:0] node2282;
	wire [11-1:0] node2286;
	wire [11-1:0] node2287;
	wire [11-1:0] node2289;
	wire [11-1:0] node2293;
	wire [11-1:0] node2294;
	wire [11-1:0] node2295;
	wire [11-1:0] node2297;
	wire [11-1:0] node2300;
	wire [11-1:0] node2301;
	wire [11-1:0] node2302;
	wire [11-1:0] node2305;
	wire [11-1:0] node2307;
	wire [11-1:0] node2310;
	wire [11-1:0] node2311;
	wire [11-1:0] node2315;
	wire [11-1:0] node2316;
	wire [11-1:0] node2317;
	wire [11-1:0] node2320;
	wire [11-1:0] node2322;
	wire [11-1:0] node2325;
	wire [11-1:0] node2326;
	wire [11-1:0] node2327;
	wire [11-1:0] node2329;
	wire [11-1:0] node2333;
	wire [11-1:0] node2336;
	wire [11-1:0] node2337;
	wire [11-1:0] node2338;
	wire [11-1:0] node2339;
	wire [11-1:0] node2340;
	wire [11-1:0] node2341;
	wire [11-1:0] node2342;
	wire [11-1:0] node2344;
	wire [11-1:0] node2347;
	wire [11-1:0] node2348;
	wire [11-1:0] node2351;
	wire [11-1:0] node2354;
	wire [11-1:0] node2355;
	wire [11-1:0] node2356;
	wire [11-1:0] node2361;
	wire [11-1:0] node2362;
	wire [11-1:0] node2363;
	wire [11-1:0] node2366;
	wire [11-1:0] node2368;
	wire [11-1:0] node2370;
	wire [11-1:0] node2373;
	wire [11-1:0] node2374;
	wire [11-1:0] node2375;
	wire [11-1:0] node2378;
	wire [11-1:0] node2381;
	wire [11-1:0] node2382;
	wire [11-1:0] node2385;
	wire [11-1:0] node2388;
	wire [11-1:0] node2389;
	wire [11-1:0] node2390;
	wire [11-1:0] node2391;
	wire [11-1:0] node2392;
	wire [11-1:0] node2394;
	wire [11-1:0] node2397;
	wire [11-1:0] node2400;
	wire [11-1:0] node2403;
	wire [11-1:0] node2404;
	wire [11-1:0] node2405;
	wire [11-1:0] node2407;
	wire [11-1:0] node2410;
	wire [11-1:0] node2413;
	wire [11-1:0] node2415;
	wire [11-1:0] node2418;
	wire [11-1:0] node2419;
	wire [11-1:0] node2420;
	wire [11-1:0] node2421;
	wire [11-1:0] node2424;
	wire [11-1:0] node2427;
	wire [11-1:0] node2429;
	wire [11-1:0] node2431;
	wire [11-1:0] node2434;
	wire [11-1:0] node2436;
	wire [11-1:0] node2437;
	wire [11-1:0] node2440;
	wire [11-1:0] node2442;
	wire [11-1:0] node2445;
	wire [11-1:0] node2446;
	wire [11-1:0] node2447;
	wire [11-1:0] node2448;
	wire [11-1:0] node2449;
	wire [11-1:0] node2450;
	wire [11-1:0] node2451;
	wire [11-1:0] node2455;
	wire [11-1:0] node2459;
	wire [11-1:0] node2460;
	wire [11-1:0] node2463;
	wire [11-1:0] node2465;
	wire [11-1:0] node2468;
	wire [11-1:0] node2469;
	wire [11-1:0] node2470;
	wire [11-1:0] node2472;
	wire [11-1:0] node2475;
	wire [11-1:0] node2476;
	wire [11-1:0] node2479;
	wire [11-1:0] node2482;
	wire [11-1:0] node2483;
	wire [11-1:0] node2485;
	wire [11-1:0] node2488;
	wire [11-1:0] node2491;
	wire [11-1:0] node2492;
	wire [11-1:0] node2493;
	wire [11-1:0] node2496;
	wire [11-1:0] node2497;
	wire [11-1:0] node2500;
	wire [11-1:0] node2501;
	wire [11-1:0] node2503;
	wire [11-1:0] node2507;
	wire [11-1:0] node2508;
	wire [11-1:0] node2509;
	wire [11-1:0] node2510;
	wire [11-1:0] node2511;
	wire [11-1:0] node2514;
	wire [11-1:0] node2518;
	wire [11-1:0] node2520;
	wire [11-1:0] node2522;
	wire [11-1:0] node2525;
	wire [11-1:0] node2526;
	wire [11-1:0] node2527;
	wire [11-1:0] node2531;
	wire [11-1:0] node2532;
	wire [11-1:0] node2535;
	wire [11-1:0] node2538;
	wire [11-1:0] node2539;
	wire [11-1:0] node2540;
	wire [11-1:0] node2541;
	wire [11-1:0] node2542;
	wire [11-1:0] node2543;
	wire [11-1:0] node2546;
	wire [11-1:0] node2549;
	wire [11-1:0] node2551;
	wire [11-1:0] node2554;
	wire [11-1:0] node2555;
	wire [11-1:0] node2556;
	wire [11-1:0] node2557;
	wire [11-1:0] node2561;
	wire [11-1:0] node2564;
	wire [11-1:0] node2565;
	wire [11-1:0] node2566;
	wire [11-1:0] node2571;
	wire [11-1:0] node2572;
	wire [11-1:0] node2573;
	wire [11-1:0] node2575;
	wire [11-1:0] node2576;
	wire [11-1:0] node2580;
	wire [11-1:0] node2583;
	wire [11-1:0] node2584;
	wire [11-1:0] node2585;
	wire [11-1:0] node2589;
	wire [11-1:0] node2591;
	wire [11-1:0] node2594;
	wire [11-1:0] node2595;
	wire [11-1:0] node2596;
	wire [11-1:0] node2597;
	wire [11-1:0] node2598;
	wire [11-1:0] node2600;
	wire [11-1:0] node2603;
	wire [11-1:0] node2606;
	wire [11-1:0] node2607;
	wire [11-1:0] node2610;
	wire [11-1:0] node2611;
	wire [11-1:0] node2615;
	wire [11-1:0] node2616;
	wire [11-1:0] node2618;
	wire [11-1:0] node2620;
	wire [11-1:0] node2623;
	wire [11-1:0] node2624;
	wire [11-1:0] node2625;
	wire [11-1:0] node2628;
	wire [11-1:0] node2632;
	wire [11-1:0] node2633;
	wire [11-1:0] node2634;
	wire [11-1:0] node2635;
	wire [11-1:0] node2638;
	wire [11-1:0] node2639;
	wire [11-1:0] node2643;
	wire [11-1:0] node2644;
	wire [11-1:0] node2645;
	wire [11-1:0] node2648;
	wire [11-1:0] node2650;
	wire [11-1:0] node2654;
	wire [11-1:0] node2655;
	wire [11-1:0] node2656;
	wire [11-1:0] node2658;
	wire [11-1:0] node2661;
	wire [11-1:0] node2664;
	wire [11-1:0] node2665;
	wire [11-1:0] node2668;

	assign outp = (inp[1]) ? node1368 : node1;
		assign node1 = (inp[7]) ? node699 : node2;
			assign node2 = (inp[2]) ? node372 : node3;
				assign node3 = (inp[0]) ? node191 : node4;
					assign node4 = (inp[4]) ? node112 : node5;
						assign node5 = (inp[9]) ? node59 : node6;
							assign node6 = (inp[5]) ? node30 : node7;
								assign node7 = (inp[6]) ? node17 : node8;
									assign node8 = (inp[11]) ? 11'b11111101001 : node9;
										assign node9 = (inp[3]) ? node13 : node10;
											assign node10 = (inp[8]) ? 11'b11001101011 : 11'b01001101011;
											assign node13 = (inp[10]) ? 11'b01100101111 : 11'b11001101011;
									assign node17 = (inp[3]) ? node27 : node18;
										assign node18 = (inp[8]) ? node22 : node19;
											assign node19 = (inp[10]) ? 11'b11000100010 : 11'b01010000010;
											assign node22 = (inp[11]) ? 11'b11110101000 : node23;
												assign node23 = (inp[10]) ? 11'b11011001010 : 11'b01000101010;
										assign node27 = (inp[10]) ? 11'b01010111110 : 11'b11101111000;
								assign node30 = (inp[6]) ? node50 : node31;
									assign node31 = (inp[8]) ? node41 : node32;
										assign node32 = (inp[10]) ? node36 : node33;
											assign node33 = (inp[3]) ? 11'b11001111010 : 11'b01001111010;
											assign node36 = (inp[11]) ? 11'b11101111000 : node37;
												assign node37 = (inp[3]) ? 11'b01100111110 : 11'b11100111010;
										assign node41 = (inp[11]) ? node45 : node42;
											assign node42 = (inp[3]) ? 11'b11000011011 : 11'b01000011011;
											assign node45 = (inp[3]) ? 11'b11010001010 : node46;
												assign node46 = (inp[10]) ? 11'b11010011010 : 11'b01001011010;
									assign node50 = (inp[10]) ? node54 : node51;
										assign node51 = (inp[8]) ? 11'b01000111011 : 11'b01001011011;
										assign node54 = (inp[11]) ? 11'b01001001111 : node55;
											assign node55 = (inp[3]) ? 11'b01110011101 : 11'b11101011001;
							assign node59 = (inp[10]) ? node87 : node60;
								assign node60 = (inp[3]) ? node76 : node61;
									assign node61 = (inp[5]) ? node67 : node62;
										assign node62 = (inp[11]) ? 11'b01101011010 : node63;
											assign node63 = (inp[6]) ? 11'b01000100000 : 11'b01001101011;
										assign node67 = (inp[6]) ? node73 : node68;
											assign node68 = (inp[8]) ? node70 : 11'b01110101000;
												assign node70 = (inp[11]) ? 11'b01001101010 : 11'b01010111010;
											assign node73 = (inp[8]) ? 11'b01010101001 : 11'b01111001011;
									assign node76 = (inp[5]) ? node82 : node77;
										assign node77 = (inp[6]) ? node79 : 11'b11111101111;
											assign node79 = (inp[11]) ? 11'b11111001110 : 11'b11100001100;
										assign node82 = (inp[6]) ? node84 : 11'b11011111100;
											assign node84 = (inp[8]) ? 11'b11100111111 : 11'b11010011111;
								assign node87 = (inp[5]) ? node103 : node88;
									assign node88 = (inp[8]) ? node98 : node89;
										assign node89 = (inp[3]) ? node91 : 11'b11110111101;
											assign node91 = (inp[11]) ? node95 : node92;
												assign node92 = (inp[6]) ? 11'b01010110100 : 11'b01000111111;
												assign node95 = (inp[6]) ? 11'b01001111111 : 11'b01010111111;
										assign node98 = (inp[11]) ? 11'b11001111101 : node99;
											assign node99 = (inp[3]) ? 11'b01111011110 : 11'b11001011110;
									assign node103 = (inp[3]) ? 11'b01101101100 : node104;
										assign node104 = (inp[8]) ? node108 : node105;
											assign node105 = (inp[11]) ? 11'b11100001101 : 11'b11111101111;
											assign node108 = (inp[11]) ? 11'b11110101110 : 11'b11000101100;
						assign node112 = (inp[5]) ? node152 : node113;
							assign node113 = (inp[6]) ? node139 : node114;
								assign node114 = (inp[10]) ? node124 : node115;
									assign node115 = (inp[3]) ? node117 : 11'b01000011111;
										assign node117 = (inp[9]) ? node119 : 11'b11001001111;
											assign node119 = (inp[11]) ? 11'b11011011011 : node120;
												assign node120 = (inp[8]) ? 11'b11011011011 : 11'b11101011011;
									assign node124 = (inp[11]) ? node128 : node125;
										assign node125 = (inp[3]) ? 11'b01010001011 : 11'b11100001011;
										assign node128 = (inp[3]) ? node134 : node129;
											assign node129 = (inp[9]) ? node131 : 11'b11111011101;
												assign node131 = (inp[8]) ? 11'b11111011011 : 11'b11110011011;
											assign node134 = (inp[8]) ? node136 : 11'b01110011011;
												assign node136 = (inp[9]) ? 11'b01111011011 : 11'b01101011011;
								assign node139 = (inp[8]) ? node147 : node140;
									assign node140 = (inp[9]) ? node144 : node141;
										assign node141 = (inp[10]) ? 11'b11110111111 : 11'b01011101111;
										assign node144 = (inp[3]) ? 11'b11011011001 : 11'b11100011011;
									assign node147 = (inp[3]) ? 11'b01001101000 : node148;
										assign node148 = (inp[10]) ? 11'b11110011100 : 11'b01010011100;
							assign node152 = (inp[11]) ? node170 : node153;
								assign node153 = (inp[9]) ? node165 : node154;
									assign node154 = (inp[10]) ? node162 : node155;
										assign node155 = (inp[8]) ? node159 : node156;
											assign node156 = (inp[3]) ? 11'b11111011110 : 11'b01011011110;
											assign node159 = (inp[6]) ? 11'b01111011101 : 11'b01111111100;
										assign node162 = (inp[6]) ? 11'b01011111001 : 11'b01010011010;
									assign node165 = (inp[6]) ? node167 : 11'b11001011000;
										assign node167 = (inp[10]) ? 11'b01111001011 : 11'b11101001001;
								assign node170 = (inp[10]) ? node180 : node171;
									assign node171 = (inp[9]) ? node177 : node172;
										assign node172 = (inp[8]) ? node174 : 11'b11111111100;
											assign node174 = (inp[6]) ? 11'b11100111101 : 11'b11101111100;
										assign node177 = (inp[8]) ? 11'b11101001000 : 11'b11101101000;
									assign node180 = (inp[3]) ? node184 : node181;
										assign node181 = (inp[8]) ? 11'b11110101100 : 11'b11001001100;
										assign node184 = (inp[8]) ? node186 : 11'b01110101000;
											assign node186 = (inp[6]) ? node188 : 11'b01110101000;
												assign node188 = (inp[9]) ? 11'b01110001001 : 11'b01111001011;
					assign node191 = (inp[3]) ? node287 : node192;
						assign node192 = (inp[11]) ? node240 : node193;
							assign node193 = (inp[6]) ? node215 : node194;
								assign node194 = (inp[5]) ? node204 : node195;
									assign node195 = (inp[9]) ? 11'b01001011011 : node196;
										assign node196 = (inp[8]) ? node200 : node197;
											assign node197 = (inp[4]) ? 11'b01001001001 : 11'b01001101001;
											assign node200 = (inp[4]) ? 11'b01100101001 : 11'b01101101101;
									assign node204 = (inp[4]) ? node212 : node205;
										assign node205 = (inp[9]) ? node207 : 11'b01100001001;
											assign node207 = (inp[10]) ? 11'b01100111000 : node208;
												assign node208 = (inp[8]) ? 11'b01110101100 : 11'b01001101100;
										assign node212 = (inp[8]) ? 11'b01010101010 : 11'b01010011100;
								assign node215 = (inp[5]) ? node231 : node216;
									assign node216 = (inp[8]) ? node224 : node217;
										assign node217 = (inp[4]) ? node221 : node218;
											assign node218 = (inp[9]) ? 11'b01011100110 : 11'b01010100100;
											assign node221 = (inp[10]) ? 11'b01011010100 : 11'b01110010110;
										assign node224 = (inp[10]) ? node226 : 11'b01110101000;
											assign node226 = (inp[4]) ? 11'b01111111110 : node227;
												assign node227 = (inp[9]) ? 11'b01101011000 : 11'b01111001100;
									assign node231 = (inp[8]) ? 11'b01110101001 : node232;
										assign node232 = (inp[4]) ? node236 : node233;
											assign node233 = (inp[9]) ? 11'b01011101111 : 11'b01011001001;
											assign node236 = (inp[9]) ? 11'b01111011001 : 11'b01001111111;
							assign node240 = (inp[9]) ? node268 : node241;
								assign node241 = (inp[10]) ? node257 : node242;
									assign node242 = (inp[6]) ? node252 : node243;
										assign node243 = (inp[5]) ? node249 : node244;
											assign node244 = (inp[8]) ? 11'b01100011011 : node245;
												assign node245 = (inp[4]) ? 11'b01011011001 : 11'b01001111001;
											assign node249 = (inp[4]) ? 11'b01101011010 : 11'b01001111010;
										assign node252 = (inp[8]) ? node254 : 11'b01010010000;
											assign node254 = (inp[4]) ? 11'b01100011000 : 11'b01110011001;
									assign node257 = (inp[5]) ? node263 : node258;
										assign node258 = (inp[8]) ? node260 : 11'b01100101111;
											assign node260 = (inp[6]) ? 11'b01011001100 : 11'b01111111111;
										assign node263 = (inp[4]) ? 11'b01110101100 : node264;
											assign node264 = (inp[8]) ? 11'b01110011100 : 11'b01010111110;
								assign node268 = (inp[10]) ? node270 : 11'b01001001110;
									assign node270 = (inp[8]) ? node278 : node271;
										assign node271 = (inp[5]) ? 11'b01100001011 : node272;
											assign node272 = (inp[4]) ? node274 : 11'b01000101001;
												assign node274 = (inp[6]) ? 11'b01100001001 : 11'b01110001001;
										assign node278 = (inp[6]) ? node280 : 11'b01101101011;
											assign node280 = (inp[5]) ? node284 : node281;
												assign node281 = (inp[4]) ? 11'b01001101001 : 11'b01110001010;
												assign node284 = (inp[4]) ? 11'b01000001011 : 11'b01001101001;
						assign node287 = (inp[10]) ? node327 : node288;
							assign node288 = (inp[5]) ? node310 : node289;
								assign node289 = (inp[4]) ? node297 : node290;
									assign node290 = (inp[6]) ? node292 : 11'b01101111001;
										assign node292 = (inp[9]) ? node294 : 11'b01001001000;
											assign node294 = (inp[11]) ? 11'b01101011010 : 11'b01011011010;
									assign node297 = (inp[9]) ? node301 : node298;
										assign node298 = (inp[11]) ? 11'b01111011001 : 11'b01001011001;
										assign node301 = (inp[6]) ? node307 : node302;
											assign node302 = (inp[11]) ? 11'b01110001001 : node303;
												assign node303 = (inp[8]) ? 11'b01111001001 : 11'b01101001001;
											assign node307 = (inp[8]) ? 11'b01111101011 : 11'b01110001011;
								assign node310 = (inp[4]) ? node318 : node311;
									assign node311 = (inp[9]) ? node315 : node312;
										assign node312 = (inp[11]) ? 11'b01100001011 : 11'b01100001001;
										assign node315 = (inp[6]) ? 11'b01100111001 : 11'b01101111000;
									assign node318 = (inp[8]) ? node324 : node319;
										assign node319 = (inp[6]) ? 11'b01001111000 : node320;
											assign node320 = (inp[9]) ? 11'b01001001010 : 11'b01001011010;
										assign node324 = (inp[9]) ? 11'b01010001010 : 11'b01010111010;
							assign node327 = (inp[4]) ? node351 : node328;
								assign node328 = (inp[9]) ? node340 : node329;
									assign node329 = (inp[11]) ? node333 : node330;
										assign node330 = (inp[8]) ? 11'b01010001010 : 11'b01000101001;
										assign node333 = (inp[6]) ? 11'b01111001001 : node334;
											assign node334 = (inp[5]) ? node336 : 11'b01110101011;
												assign node336 = (inp[8]) ? 11'b01101101000 : 11'b01110101010;
									assign node340 = (inp[5]) ? node344 : node341;
										assign node341 = (inp[11]) ? 11'b01011101001 : 11'b01000100000;
										assign node344 = (inp[11]) ? node346 : 11'b01011101010;
											assign node346 = (inp[6]) ? 11'b01001101010 : node347;
												assign node347 = (inp[8]) ? 11'b01001101010 : 11'b01000101010;
								assign node351 = (inp[5]) ? node363 : node352;
									assign node352 = (inp[9]) ? node358 : node353;
										assign node353 = (inp[8]) ? 11'b01000001010 : node354;
											assign node354 = (inp[6]) ? 11'b01011001011 : 11'b01010001001;
										assign node358 = (inp[8]) ? node360 : 11'b01000001001;
											assign node360 = (inp[6]) ? 11'b01001101001 : 11'b01001001001;
									assign node363 = (inp[6]) ? 11'b01001001011 : node364;
										assign node364 = (inp[8]) ? node368 : node365;
											assign node365 = (inp[11]) ? 11'b01000001000 : 11'b01000001010;
											assign node368 = (inp[9]) ? 11'b01001001000 : 11'b01001001010;
				assign node372 = (inp[0]) ? node528 : node373;
					assign node373 = (inp[8]) ? node437 : node374;
						assign node374 = (inp[5]) ? node402 : node375;
							assign node375 = (inp[6]) ? node385 : node376;
								assign node376 = (inp[9]) ? node380 : node377;
									assign node377 = (inp[11]) ? 11'b01100010111 : 11'b01110001110;
									assign node380 = (inp[10]) ? 11'b11011000001 : node381;
										assign node381 = (inp[3]) ? 11'b11011100111 : 11'b01110110101;
								assign node385 = (inp[10]) ? node395 : node386;
									assign node386 = (inp[4]) ? node390 : node387;
										assign node387 = (inp[3]) ? 11'b11101001011 : 11'b01011011000;
										assign node390 = (inp[9]) ? 11'b11110111000 : node391;
											assign node391 = (inp[11]) ? 11'b01110001100 : 11'b01100101100;
									assign node395 = (inp[3]) ? node399 : node396;
										assign node396 = (inp[9]) ? 11'b11111111110 : 11'b11011111110;
										assign node399 = (inp[9]) ? 11'b01011111010 : 11'b01011101010;
							assign node402 = (inp[9]) ? node424 : node403;
								assign node403 = (inp[10]) ? node413 : node404;
									assign node404 = (inp[4]) ? node408 : node405;
										assign node405 = (inp[6]) ? 11'b01110110001 : 11'b01100010011;
										assign node408 = (inp[6]) ? 11'b01111011100 : node409;
											assign node409 = (inp[11]) ? 11'b01101110110 : 11'b11000110110;
									assign node413 = (inp[4]) ? node421 : node414;
										assign node414 = (inp[3]) ? 11'b01001010101 : node415;
											assign node415 = (inp[11]) ? node417 : 11'b11000111000;
												assign node417 = (inp[6]) ? 11'b11001110011 : 11'b11000010000;
										assign node421 = (inp[3]) ? 11'b01000000011 : 11'b11100000101;
								assign node424 = (inp[4]) ? node428 : node425;
									assign node425 = (inp[6]) ? 11'b11100011110 : 11'b01110000110;
									assign node428 = (inp[6]) ? node430 : 11'b11101100000;
										assign node430 = (inp[11]) ? node432 : 11'b11101100011;
											assign node432 = (inp[3]) ? 11'b11011000011 : node433;
												assign node433 = (inp[10]) ? 11'b11111000001 : 11'b01111000111;
						assign node437 = (inp[4]) ? node477 : node438;
							assign node438 = (inp[9]) ? node456 : node439;
								assign node439 = (inp[3]) ? node449 : node440;
									assign node440 = (inp[10]) ? node444 : node441;
										assign node441 = (inp[6]) ? 11'b01111110010 : 11'b01101110011;
										assign node444 = (inp[5]) ? 11'b11001110001 : node445;
											assign node445 = (inp[6]) ? 11'b11101100001 : 11'b11111000010;
									assign node449 = (inp[6]) ? node453 : node450;
										assign node450 = (inp[11]) ? 11'b01111010101 : 11'b01010110101;
										assign node453 = (inp[5]) ? 11'b11111100010 : 11'b11011010001;
								assign node456 = (inp[11]) ? node470 : node457;
									assign node457 = (inp[6]) ? node465 : node458;
										assign node458 = (inp[5]) ? 11'b01000000111 : node459;
											assign node459 = (inp[10]) ? node461 : 11'b01110000010;
												assign node461 = (inp[3]) ? 11'b01011010100 : 11'b11101010100;
										assign node465 = (inp[5]) ? node467 : 11'b11111110111;
											assign node467 = (inp[10]) ? 11'b11101000100 : 11'b11100010100;
									assign node470 = (inp[5]) ? 11'b11011010110 : node471;
										assign node471 = (inp[3]) ? 11'b11000000101 : node472;
											assign node472 = (inp[6]) ? 11'b01000010001 : 11'b01001010011;
							assign node477 = (inp[5]) ? node503 : node478;
								assign node478 = (inp[10]) ? node486 : node479;
									assign node479 = (inp[11]) ? node483 : node480;
										assign node480 = (inp[3]) ? 11'b11100100111 : 11'b01000000100;
										assign node483 = (inp[9]) ? 11'b11111110000 : 11'b11110100100;
									assign node486 = (inp[3]) ? node492 : node487;
										assign node487 = (inp[11]) ? 11'b11000110011 : node488;
											assign node488 = (inp[6]) ? 11'b11110000011 : 11'b11111100011;
										assign node492 = (inp[9]) ? node498 : node493;
											assign node493 = (inp[11]) ? node495 : 11'b01100100001;
												assign node495 = (inp[6]) ? 11'b01011110010 : 11'b01000010001;
											assign node498 = (inp[11]) ? node500 : 11'b01010010011;
												assign node500 = (inp[6]) ? 11'b01010110010 : 11'b01010110011;
								assign node503 = (inp[11]) ? node515 : node504;
									assign node504 = (inp[9]) ? node508 : node505;
										assign node505 = (inp[6]) ? 11'b11110000100 : 11'b11111000111;
										assign node508 = (inp[6]) ? node512 : node509;
											assign node509 = (inp[3]) ? 11'b11000000001 : 11'b01010010101;
											assign node512 = (inp[10]) ? 11'b01010100000 : 11'b01011110110;
									assign node515 = (inp[10]) ? node523 : node516;
										assign node516 = (inp[9]) ? node518 : 11'b11010010110;
											assign node518 = (inp[3]) ? node520 : 11'b01011000110;
												assign node520 = (inp[6]) ? 11'b11010000010 : 11'b11011000000;
										assign node523 = (inp[3]) ? node525 : 11'b11010000000;
											assign node525 = (inp[6]) ? 11'b01011000000 : 11'b01011000010;
					assign node528 = (inp[3]) ? node606 : node529;
						assign node529 = (inp[5]) ? node575 : node530;
							assign node530 = (inp[6]) ? node552 : node531;
								assign node531 = (inp[11]) ? node541 : node532;
									assign node532 = (inp[4]) ? node534 : 11'b01001100101;
										assign node534 = (inp[8]) ? node536 : 11'b01010110111;
											assign node536 = (inp[10]) ? node538 : 11'b01000110101;
												assign node538 = (inp[9]) ? 11'b01011110001 : 11'b01101110101;
									assign node541 = (inp[4]) ? node547 : node542;
										assign node542 = (inp[10]) ? node544 : 11'b01010010001;
											assign node544 = (inp[8]) ? 11'b01101010111 : 11'b01001100011;
										assign node547 = (inp[8]) ? node549 : 11'b01101100111;
											assign node549 = (inp[9]) ? 11'b01111100111 : 11'b01010000111;
								assign node552 = (inp[8]) ? node568 : node553;
									assign node553 = (inp[9]) ? node559 : node554;
										assign node554 = (inp[11]) ? node556 : 11'b01011001001;
											assign node556 = (inp[4]) ? 11'b01001111010 : 11'b01010011110;
										assign node559 = (inp[10]) ? node565 : node560;
											assign node560 = (inp[11]) ? 11'b01101011100 : node561;
												assign node561 = (inp[4]) ? 11'b01110111100 : 11'b01011101110;
											assign node565 = (inp[4]) ? 11'b01101011010 : 11'b01001111000;
									assign node568 = (inp[9]) ? node572 : node569;
										assign node569 = (inp[4]) ? 11'b01110100011 : 11'b01110000001;
										assign node572 = (inp[4]) ? 11'b01000010001 : 11'b01101110011;
							assign node575 = (inp[10]) ? node589 : node576;
								assign node576 = (inp[11]) ? node582 : node577;
									assign node577 = (inp[9]) ? node579 : 11'b01110100010;
										assign node579 = (inp[4]) ? 11'b01101110100 : 11'b01110000100;
									assign node582 = (inp[8]) ? node586 : node583;
										assign node583 = (inp[4]) ? 11'b01101110000 : 11'b01011010010;
										assign node586 = (inp[4]) ? 11'b01011010000 : 11'b01110110000;
								assign node589 = (inp[9]) ? node593 : node590;
									assign node590 = (inp[4]) ? 11'b01010110100 : 11'b01000010110;
									assign node593 = (inp[8]) ? node597 : node594;
										assign node594 = (inp[11]) ? 11'b01100100001 : 11'b01101110010;
										assign node597 = (inp[11]) ? node603 : node598;
											assign node598 = (inp[4]) ? node600 : 11'b01011010010;
												assign node600 = (inp[6]) ? 11'b01000110010 : 11'b01011110010;
											assign node603 = (inp[4]) ? 11'b01000000010 : 11'b01011000010;
						assign node606 = (inp[8]) ? node654 : node607;
							assign node607 = (inp[6]) ? node625 : node608;
								assign node608 = (inp[10]) ? node616 : node609;
									assign node609 = (inp[5]) ? node613 : node610;
										assign node610 = (inp[11]) ? 11'b01011000001 : 11'b01011001000;
										assign node613 = (inp[4]) ? 11'b01010100000 : 11'b01110000010;
									assign node616 = (inp[4]) ? node620 : node617;
										assign node617 = (inp[11]) ? 11'b01100000001 : 11'b01000001000;
										assign node620 = (inp[9]) ? node622 : 11'b01010100011;
											assign node622 = (inp[11]) ? 11'b01001000001 : 11'b01000000001;
								assign node625 = (inp[5]) ? node641 : node626;
									assign node626 = (inp[4]) ? node632 : node627;
										assign node627 = (inp[10]) ? 11'b01101001010 : node628;
											assign node628 = (inp[11]) ? 11'b01111011000 : 11'b01011001001;
										assign node632 = (inp[10]) ? node636 : node633;
											assign node633 = (inp[11]) ? 11'b01101101010 : 11'b01011111010;
											assign node636 = (inp[11]) ? 11'b01010101000 : node637;
												assign node637 = (inp[9]) ? 11'b01001001000 : 11'b01101101000;
									assign node641 = (inp[11]) ? node647 : node642;
										assign node642 = (inp[10]) ? 11'b01110001010 : node643;
											assign node643 = (inp[4]) ? 11'b01011100001 : 11'b01110011000;
										assign node647 = (inp[10]) ? 11'b01010000001 : node648;
											assign node648 = (inp[9]) ? node650 : 11'b01111100011;
												assign node650 = (inp[4]) ? 11'b01001000011 : 11'b01000110011;
							assign node654 = (inp[5]) ? node676 : node655;
								assign node655 = (inp[10]) ? node663 : node656;
									assign node656 = (inp[11]) ? node660 : node657;
										assign node657 = (inp[9]) ? 11'b01000110001 : 11'b01011110011;
										assign node660 = (inp[4]) ? 11'b01101100001 : 11'b01001000001;
									assign node663 = (inp[6]) ? node669 : node664;
										assign node664 = (inp[11]) ? 11'b01011000001 : node665;
											assign node665 = (inp[9]) ? 11'b01000000010 : 11'b01010000000;
										assign node669 = (inp[11]) ? node671 : 11'b01001100011;
											assign node671 = (inp[4]) ? node673 : 11'b01011100000;
												assign node673 = (inp[9]) ? 11'b01000100000 : 11'b01001100000;
								assign node676 = (inp[9]) ? node686 : node677;
									assign node677 = (inp[6]) ? node683 : node678;
										assign node678 = (inp[10]) ? node680 : 11'b01100100000;
											assign node680 = (inp[4]) ? 11'b01100000011 : 11'b01010100011;
										assign node683 = (inp[10]) ? 11'b01101100000 : 11'b01100010010;
									assign node686 = (inp[4]) ? node694 : node687;
										assign node687 = (inp[11]) ? node691 : node688;
											assign node688 = (inp[10]) ? 11'b01011000000 : 11'b01111010010;
											assign node691 = (inp[6]) ? 11'b01001010010 : 11'b01000110010;
										assign node694 = (inp[10]) ? 11'b01000000000 : node695;
											assign node695 = (inp[11]) ? 11'b01000000010 : 11'b01000100010;
			assign node699 = (inp[6]) ? node1055 : node700;
				assign node700 = (inp[2]) ? node864 : node701;
					assign node701 = (inp[8]) ? node779 : node702;
						assign node702 = (inp[5]) ? node738 : node703;
							assign node703 = (inp[0]) ? node717 : node704;
								assign node704 = (inp[11]) ? node710 : node705;
									assign node705 = (inp[4]) ? 11'b01010100111 : node706;
										assign node706 = (inp[3]) ? 11'b01011110101 : 11'b11011110101;
									assign node710 = (inp[4]) ? node714 : node711;
										assign node711 = (inp[3]) ? 11'b11111100111 : 11'b01011000011;
										assign node714 = (inp[3]) ? 11'b01101110011 : 11'b01001110111;
								assign node717 = (inp[3]) ? node729 : node718;
									assign node718 = (inp[10]) ? node724 : node719;
										assign node719 = (inp[9]) ? 11'b01100010101 : node720;
											assign node720 = (inp[11]) ? 11'b01001010001 : 11'b01001100001;
										assign node724 = (inp[11]) ? node726 : 11'b01001010111;
											assign node726 = (inp[4]) ? 11'b01111100111 : 11'b01011100011;
									assign node729 = (inp[10]) ? node735 : node730;
										assign node730 = (inp[9]) ? node732 : 11'b01000110011;
											assign node732 = (inp[11]) ? 11'b01110100011 : 11'b01100000011;
										assign node735 = (inp[4]) ? 11'b01000100001 : 11'b01100000001;
							assign node738 = (inp[11]) ? node758 : node739;
								assign node739 = (inp[4]) ? node749 : node740;
									assign node740 = (inp[10]) ? node744 : node741;
										assign node741 = (inp[9]) ? 11'b01101010011 : 11'b01001000011;
										assign node744 = (inp[3]) ? 11'b01011000001 : node745;
											assign node745 = (inp[9]) ? 11'b01101010001 : 11'b01101000101;
									assign node749 = (inp[9]) ? node755 : node750;
										assign node750 = (inp[0]) ? node752 : 11'b11000000111;
											assign node752 = (inp[3]) ? 11'b01110010011 : 11'b01010010101;
										assign node755 = (inp[3]) ? 11'b01110100010 : 11'b11010110010;
								assign node758 = (inp[4]) ? node770 : node759;
									assign node759 = (inp[10]) ? node763 : node760;
										assign node760 = (inp[0]) ? 11'b01101100000 : 11'b11111100000;
										assign node763 = (inp[9]) ? node767 : node764;
											assign node764 = (inp[0]) ? 11'b01011110100 : 11'b01001100100;
											assign node767 = (inp[0]) ? 11'b01111000000 : 11'b01011000100;
									assign node770 = (inp[10]) ? node774 : node771;
										assign node771 = (inp[9]) ? 11'b01111000100 : 11'b01101010000;
										assign node774 = (inp[9]) ? node776 : 11'b01011000010;
											assign node776 = (inp[0]) ? 11'b01110000010 : 11'b01100000000;
						assign node779 = (inp[5]) ? node837 : node780;
							assign node780 = (inp[11]) ? node812 : node781;
								assign node781 = (inp[0]) ? node801 : node782;
									assign node782 = (inp[9]) ? node792 : node783;
										assign node783 = (inp[10]) ? 11'b11110110100 : node784;
											assign node784 = (inp[3]) ? node788 : node785;
												assign node785 = (inp[4]) ? 11'b01111100110 : 11'b01010000010;
												assign node788 = (inp[4]) ? 11'b11011100100 : 11'b11111100010;
										assign node792 = (inp[10]) ? node796 : node793;
											assign node793 = (inp[3]) ? 11'b11100100100 : 11'b01100100100;
											assign node796 = (inp[3]) ? node798 : 11'b11000110100;
												assign node798 = (inp[4]) ? 11'b01110010010 : 11'b01101110110;
									assign node801 = (inp[4]) ? node807 : node802;
										assign node802 = (inp[3]) ? node804 : 11'b01100000000;
											assign node804 = (inp[10]) ? 11'b01001100000 : 11'b01001100010;
										assign node807 = (inp[9]) ? 11'b01011010110 : node808;
											assign node808 = (inp[3]) ? 11'b01000110010 : 11'b01101100010;
								assign node812 = (inp[4]) ? node826 : node813;
									assign node813 = (inp[0]) ? node819 : node814;
										assign node814 = (inp[3]) ? node816 : 11'b01010000000;
											assign node816 = (inp[10]) ? 11'b01110010100 : 11'b11110000110;
										assign node819 = (inp[10]) ? node821 : 11'b01100010000;
											assign node821 = (inp[9]) ? 11'b00011101011 : node822;
												assign node822 = (inp[3]) ? 11'b01111000010 : 11'b01111010100;
									assign node826 = (inp[0]) ? node834 : node827;
										assign node827 = (inp[10]) ? node831 : node828;
											assign node828 = (inp[3]) ? 11'b10000111001 : 11'b00010111111;
											assign node831 = (inp[9]) ? 11'b10101111001 : 11'b00110111001;
										assign node834 = (inp[3]) ? 11'b00111101011 : 11'b00100101101;
							assign node837 = (inp[0]) ? node849 : node838;
								assign node838 = (inp[4]) ? node846 : node839;
									assign node839 = (inp[10]) ? node843 : node840;
										assign node840 = (inp[11]) ? 11'b10001101001 : 11'b10010111001;
										assign node843 = (inp[3]) ? 11'b00010101111 : 11'b10000111001;
									assign node846 = (inp[3]) ? 11'b10001011111 : 11'b00110111101;
								assign node849 = (inp[10]) ? node857 : node850;
									assign node850 = (inp[9]) ? 11'b00001111111 : node851;
										assign node851 = (inp[4]) ? 11'b00111011001 : node852;
											assign node852 = (inp[11]) ? 11'b00110101011 : 11'b00100101011;
									assign node857 = (inp[9]) ? 11'b00001101001 : node858;
										assign node858 = (inp[3]) ? 11'b00011001001 : node859;
											assign node859 = (inp[11]) ? 11'b00011001101 : 11'b00010101101;
					assign node864 = (inp[0]) ? node964 : node865;
						assign node865 = (inp[8]) ? node919 : node866;
							assign node866 = (inp[11]) ? node896 : node867;
								assign node867 = (inp[4]) ? node883 : node868;
									assign node868 = (inp[9]) ? node874 : node869;
										assign node869 = (inp[5]) ? 11'b00110111010 : node870;
											assign node870 = (inp[3]) ? 11'b10111001011 : 11'b00111001011;
										assign node874 = (inp[3]) ? node876 : 11'b10010101110;
											assign node876 = (inp[10]) ? node880 : node877;
												assign node877 = (inp[5]) ? 11'b10101111110 : 11'b10110001101;
												assign node880 = (inp[5]) ? 11'b00110101100 : 11'b00101111110;
									assign node883 = (inp[9]) ? node889 : node884;
										assign node884 = (inp[10]) ? 11'b10111001100 : node885;
											assign node885 = (inp[3]) ? 11'b10110101100 : 11'b00100111110;
										assign node889 = (inp[5]) ? 11'b10110001000 : node890;
											assign node890 = (inp[3]) ? node892 : 11'b00011101100;
												assign node892 = (inp[10]) ? 11'b00010111000 : 11'b10001111010;
								assign node896 = (inp[5]) ? node908 : node897;
									assign node897 = (inp[3]) ? node903 : node898;
										assign node898 = (inp[9]) ? 11'b00100011110 : node899;
											assign node899 = (inp[10]) ? 11'b10101001000 : 11'b00101001100;
										assign node903 = (inp[9]) ? 11'b10111111010 : node904;
											assign node904 = (inp[4]) ? 11'b00000011000 : 11'b10100111000;
									assign node908 = (inp[10]) ? node914 : node909;
										assign node909 = (inp[9]) ? 11'b00000001010 : node910;
											assign node910 = (inp[4]) ? 11'b00110111111 : 11'b00111011000;
										assign node914 = (inp[4]) ? node916 : 11'b00101101111;
											assign node916 = (inp[9]) ? 11'b10110101011 : 11'b10100101111;
							assign node919 = (inp[5]) ? node945 : node920;
								assign node920 = (inp[3]) ? node936 : node921;
									assign node921 = (inp[10]) ? node931 : node922;
										assign node922 = (inp[4]) ? node926 : node923;
											assign node923 = (inp[9]) ? 11'b00101001001 : 11'b00111101001;
											assign node926 = (inp[9]) ? 11'b00111011101 : node927;
												assign node927 = (inp[11]) ? 11'b00000101101 : 11'b00011001101;
										assign node931 = (inp[11]) ? node933 : 11'b10101001001;
											assign node933 = (inp[4]) ? 11'b10001011111 : 11'b10101111101;
									assign node936 = (inp[11]) ? node940 : node937;
										assign node937 = (inp[9]) ? 11'b10010001101 : 11'b10000101001;
										assign node940 = (inp[10]) ? node942 : 11'b10000111011;
											assign node942 = (inp[4]) ? 11'b00000011011 : 11'b00010111111;
								assign node945 = (inp[9]) ? node957 : node946;
									assign node946 = (inp[11]) ? node950 : node947;
										assign node947 = (inp[3]) ? 11'b10101011001 : 11'b10011011011;
										assign node950 = (inp[4]) ? 11'b10000011100 : node951;
											assign node951 = (inp[3]) ? node953 : 11'b10110111000;
												assign node953 = (inp[10]) ? 11'b00101001110 : 11'b10100101000;
									assign node957 = (inp[3]) ? node959 : 11'b00011001100;
										assign node959 = (inp[10]) ? 11'b00011101100 : node960;
											assign node960 = (inp[4]) ? 11'b10011101010 : 11'b10110011111;
						assign node964 = (inp[3]) ? node1014 : node965;
							assign node965 = (inp[8]) ? node983 : node966;
								assign node966 = (inp[9]) ? node976 : node967;
									assign node967 = (inp[5]) ? node973 : node968;
										assign node968 = (inp[11]) ? 11'b00001011100 : node969;
											assign node969 = (inp[4]) ? 11'b00000101010 : 11'b00010001111;
										assign node973 = (inp[4]) ? 11'b00011011110 : 11'b00011011010;
									assign node976 = (inp[10]) ? node978 : 11'b00110011110;
										assign node978 = (inp[11]) ? 11'b00111101011 : node979;
											assign node979 = (inp[5]) ? 11'b00100111010 : 11'b00110111010;
								assign node983 = (inp[11]) ? node1005 : node984;
									assign node984 = (inp[10]) ? node994 : node985;
										assign node985 = (inp[9]) ? node989 : node986;
											assign node986 = (inp[5]) ? 11'b00101001011 : 11'b00100101001;
											assign node989 = (inp[4]) ? 11'b00000011111 : node990;
												assign node990 = (inp[5]) ? 11'b00100001101 : 11'b00110001111;
										assign node994 = (inp[9]) ? node1000 : node995;
											assign node995 = (inp[4]) ? node997 : 11'b00001001101;
												assign node997 = (inp[5]) ? 11'b00110111100 : 11'b00100011111;
											assign node1000 = (inp[5]) ? 11'b00001111010 : node1001;
												assign node1001 = (inp[4]) ? 11'b00011111001 : 11'b00110011001;
									assign node1005 = (inp[9]) ? node1009 : node1006;
										assign node1006 = (inp[4]) ? 11'b00010011000 : 11'b00110111000;
										assign node1009 = (inp[10]) ? 11'b00010001011 : node1010;
											assign node1010 = (inp[5]) ? 11'b00011011110 : 11'b00111001101;
							assign node1014 = (inp[4]) ? node1032 : node1015;
								assign node1015 = (inp[8]) ? node1019 : node1016;
									assign node1016 = (inp[11]) ? 11'b00011001010 : 11'b00001101010;
									assign node1019 = (inp[9]) ? node1025 : node1020;
										assign node1020 = (inp[5]) ? 11'b00010001011 : node1021;
											assign node1021 = (inp[10]) ? 11'b00011001001 : 11'b00011001011;
										assign node1025 = (inp[10]) ? node1029 : node1026;
											assign node1026 = (inp[11]) ? 11'b00111111011 : 11'b00110011001;
											assign node1029 = (inp[11]) ? 11'b00010101001 : 11'b00011101000;
								assign node1032 = (inp[5]) ? node1044 : node1033;
									assign node1033 = (inp[8]) ? node1039 : node1034;
										assign node1034 = (inp[10]) ? 11'b00101101010 : node1035;
											assign node1035 = (inp[9]) ? 11'b00101101010 : 11'b00101011000;
										assign node1039 = (inp[9]) ? 11'b00101101011 : node1040;
											assign node1040 = (inp[10]) ? 11'b00110001001 : 11'b00011011001;
									assign node1044 = (inp[8]) ? node1048 : node1045;
										assign node1045 = (inp[10]) ? 11'b00011101011 : 11'b00010001010;
										assign node1048 = (inp[11]) ? 11'b00001001010 : node1049;
											assign node1049 = (inp[9]) ? 11'b00001101000 : node1050;
												assign node1050 = (inp[10]) ? 11'b00100101010 : 11'b00100111010;
				assign node1055 = (inp[0]) ? node1211 : node1056;
					assign node1056 = (inp[8]) ? node1138 : node1057;
						assign node1057 = (inp[5]) ? node1101 : node1058;
							assign node1058 = (inp[2]) ? node1080 : node1059;
								assign node1059 = (inp[9]) ? node1067 : node1060;
									assign node1060 = (inp[11]) ? node1064 : node1061;
										assign node1061 = (inp[4]) ? 11'b00011101110 : 11'b10001101000;
										assign node1064 = (inp[4]) ? 11'b10110001100 : 11'b10000001010;
									assign node1067 = (inp[4]) ? node1075 : node1068;
										assign node1068 = (inp[10]) ? node1072 : node1069;
											assign node1069 = (inp[11]) ? 11'b00101011000 : 11'b00010101000;
											assign node1072 = (inp[11]) ? 11'b00010011100 : 11'b00001111100;
										assign node1075 = (inp[11]) ? 11'b00100110011 : node1076;
											assign node1076 = (inp[10]) ? 11'b00101011000 : 11'b10101011010;
								assign node1080 = (inp[4]) ? node1092 : node1081;
									assign node1081 = (inp[11]) ? node1083 : 11'b10101000010;
										assign node1083 = (inp[9]) ? node1089 : node1084;
											assign node1084 = (inp[3]) ? node1086 : 11'b10110100011;
												assign node1086 = (inp[10]) ? 11'b00100110101 : 11'b10111110001;
											assign node1089 = (inp[10]) ? 11'b10011010101 : 11'b10000100101;
									assign node1092 = (inp[11]) ? 11'b10000010101 : node1093;
										assign node1093 = (inp[3]) ? node1095 : 11'b00000100101;
											assign node1095 = (inp[10]) ? node1097 : 11'b10010110001;
												assign node1097 = (inp[9]) ? 11'b00001110001 : 11'b00000100011;
							assign node1101 = (inp[9]) ? node1119 : node1102;
								assign node1102 = (inp[10]) ? node1114 : node1103;
									assign node1103 = (inp[3]) ? node1109 : node1104;
										assign node1104 = (inp[2]) ? node1106 : 11'b00010110101;
											assign node1106 = (inp[11]) ? 11'b00110010111 : 11'b00110010011;
										assign node1109 = (inp[11]) ? 11'b10110000011 : node1110;
											assign node1110 = (inp[4]) ? 11'b10111010101 : 11'b10110010001;
									assign node1114 = (inp[2]) ? node1116 : 11'b10000100101;
										assign node1116 = (inp[11]) ? 11'b10111000111 : 11'b10100100111;
								assign node1119 = (inp[4]) ? node1133 : node1120;
									assign node1120 = (inp[10]) ? node1126 : node1121;
										assign node1121 = (inp[3]) ? node1123 : 11'b00000110011;
											assign node1123 = (inp[2]) ? 11'b10101010111 : 11'b10001110101;
										assign node1126 = (inp[3]) ? node1130 : node1127;
											assign node1127 = (inp[2]) ? 11'b10001000101 : 11'b10111100111;
											assign node1130 = (inp[11]) ? 11'b00001100101 : 11'b00111100101;
									assign node1133 = (inp[11]) ? node1135 : 11'b10101110001;
										assign node1135 = (inp[10]) ? 11'b10100000011 : 11'b10001000001;
						assign node1138 = (inp[4]) ? node1174 : node1139;
							assign node1139 = (inp[3]) ? node1163 : node1140;
								assign node1140 = (inp[10]) ? node1150 : node1141;
									assign node1141 = (inp[5]) ? node1145 : node1142;
										assign node1142 = (inp[9]) ? 11'b00001000001 : 11'b00010100011;
										assign node1145 = (inp[2]) ? node1147 : 11'b00000110010;
											assign node1147 = (inp[11]) ? 11'b00100000010 : 11'b00110110010;
									assign node1150 = (inp[9]) ? node1156 : node1151;
										assign node1151 = (inp[2]) ? node1153 : 11'b10100010010;
											assign node1153 = (inp[11]) ? 11'b10001000000 : 11'b10111100010;
										assign node1156 = (inp[2]) ? node1160 : node1157;
											assign node1157 = (inp[11]) ? 11'b10001110110 : 11'b10010010101;
											assign node1160 = (inp[11]) ? 11'b10110010100 : 11'b10100110110;
								assign node1163 = (inp[10]) ? node1171 : node1164;
									assign node1164 = (inp[11]) ? node1168 : node1165;
										assign node1165 = (inp[9]) ? 11'b10001010100 : 11'b10111110000;
										assign node1168 = (inp[9]) ? 11'b10110110110 : 11'b10010100000;
									assign node1171 = (inp[2]) ? 11'b00010100100 : 11'b00001100100;
							assign node1174 = (inp[3]) ? node1192 : node1175;
								assign node1175 = (inp[11]) ? node1185 : node1176;
									assign node1176 = (inp[10]) ? node1180 : node1177;
										assign node1177 = (inp[9]) ? 11'b00011100100 : 11'b00000100110;
										assign node1180 = (inp[5]) ? node1182 : 11'b10101010111;
											assign node1182 = (inp[2]) ? 11'b10101100110 : 11'b10010000100;
									assign node1185 = (inp[2]) ? node1187 : 11'b10110110100;
										assign node1187 = (inp[10]) ? node1189 : 11'b00101010100;
											assign node1189 = (inp[9]) ? 11'b10000010000 : 11'b10001010100;
								assign node1192 = (inp[10]) ? node1204 : node1193;
									assign node1193 = (inp[9]) ? node1199 : node1194;
										assign node1194 = (inp[2]) ? node1196 : 11'b10000010110;
											assign node1196 = (inp[11]) ? 11'b10001010100 : 11'b10101110100;
										assign node1199 = (inp[11]) ? 11'b10011010010 : node1200;
											assign node1200 = (inp[5]) ? 11'b10000100000 : 11'b10100110010;
									assign node1204 = (inp[11]) ? node1208 : node1205;
										assign node1205 = (inp[9]) ? 11'b00101110010 : 11'b00101110000;
										assign node1208 = (inp[9]) ? 11'b00101010010 : 11'b00101000010;
					assign node1211 = (inp[3]) ? node1313 : node1212;
						assign node1212 = (inp[8]) ? node1266 : node1213;
							assign node1213 = (inp[5]) ? node1241 : node1214;
								assign node1214 = (inp[2]) ? node1232 : node1215;
									assign node1215 = (inp[9]) ? node1227 : node1216;
										assign node1216 = (inp[11]) ? node1222 : node1217;
											assign node1217 = (inp[10]) ? node1219 : 11'b00011101000;
												assign node1219 = (inp[4]) ? 11'b00010111100 : 11'b00011101100;
											assign node1222 = (inp[10]) ? node1224 : 11'b00000011010;
												assign node1224 = (inp[4]) ? 11'b00101100101 : 11'b00010011100;
										assign node1227 = (inp[4]) ? node1229 : 11'b00111011110;
											assign node1229 = (inp[11]) ? 11'b00100100011 : 11'b00111011010;
									assign node1232 = (inp[9]) ? 11'b00100110101 : node1233;
										assign node1233 = (inp[10]) ? node1237 : node1234;
											assign node1234 = (inp[11]) ? 11'b00001110011 : 11'b00011100011;
											assign node1237 = (inp[4]) ? 11'b00000110111 : 11'b00001000100;
								assign node1241 = (inp[4]) ? node1257 : node1242;
									assign node1242 = (inp[10]) ? node1252 : node1243;
										assign node1243 = (inp[11]) ? node1247 : node1244;
											assign node1244 = (inp[9]) ? 11'b00010100101 : 11'b00011100011;
											assign node1247 = (inp[9]) ? node1249 : 11'b00000110001;
												assign node1249 = (inp[2]) ? 11'b00101010111 : 11'b00101110111;
										assign node1252 = (inp[2]) ? node1254 : 11'b00111010011;
											assign node1254 = (inp[9]) ? 11'b00100000011 : 11'b00100000111;
									assign node1257 = (inp[9]) ? node1259 : 11'b00101000011;
										assign node1259 = (inp[2]) ? node1263 : node1260;
											assign node1260 = (inp[10]) ? 11'b00111010001 : 11'b00100010101;
											assign node1263 = (inp[10]) ? 11'b00101110001 : 11'b00111110101;
							assign node1266 = (inp[5]) ? node1292 : node1267;
								assign node1267 = (inp[2]) ? node1283 : node1268;
									assign node1268 = (inp[11]) ? node1276 : node1269;
										assign node1269 = (inp[4]) ? 11'b00000010101 : node1270;
											assign node1270 = (inp[9]) ? 11'b00101000101 : node1271;
												assign node1271 = (inp[10]) ? 11'b00111000101 : 11'b00110100001;
										assign node1276 = (inp[10]) ? node1280 : node1277;
											assign node1277 = (inp[4]) ? 11'b00111000110 : 11'b00010110110;
											assign node1280 = (inp[4]) ? 11'b00010100100 : 11'b00111100000;
									assign node1283 = (inp[4]) ? node1285 : 11'b00100110000;
										assign node1285 = (inp[9]) ? node1289 : node1286;
											assign node1286 = (inp[10]) ? 11'b00111110100 : 11'b00110100000;
											assign node1289 = (inp[10]) ? 11'b00000110000 : 11'b00011110100;
								assign node1292 = (inp[9]) ? node1306 : node1293;
									assign node1293 = (inp[10]) ? node1301 : node1294;
										assign node1294 = (inp[4]) ? node1298 : node1295;
											assign node1295 = (inp[2]) ? 11'b00111100010 : 11'b00110000010;
											assign node1298 = (inp[11]) ? 11'b00011010010 : 11'b00000000000;
										assign node1301 = (inp[11]) ? node1303 : 11'b00000000110;
											assign node1303 = (inp[4]) ? 11'b00001000110 : 11'b00101110100;
									assign node1306 = (inp[2]) ? 11'b00000010110 : node1307;
										assign node1307 = (inp[10]) ? 11'b00010110010 : node1308;
											assign node1308 = (inp[4]) ? 11'b00001110110 : 11'b00011110100;
						assign node1313 = (inp[10]) ? node1337 : node1314;
							assign node1314 = (inp[11]) ? node1326 : node1315;
								assign node1315 = (inp[4]) ? node1323 : node1316;
									assign node1316 = (inp[9]) ? node1320 : node1317;
										assign node1317 = (inp[8]) ? 11'b00011100010 : 11'b00011000010;
										assign node1320 = (inp[8]) ? 11'b00000110010 : 11'b00010010010;
									assign node1323 = (inp[9]) ? 11'b00011100000 : 11'b00001010001;
								assign node1326 = (inp[8]) ? node1334 : node1327;
									assign node1327 = (inp[2]) ? 11'b00110100001 : node1328;
										assign node1328 = (inp[5]) ? 11'b00011110011 : node1329;
											assign node1329 = (inp[9]) ? 11'b00110100001 : 11'b00111110011;
									assign node1334 = (inp[5]) ? 11'b00010110010 : 11'b00100110000;
							assign node1337 = (inp[5]) ? node1351 : node1338;
								assign node1338 = (inp[8]) ? node1346 : node1339;
									assign node1339 = (inp[9]) ? node1343 : node1340;
										assign node1340 = (inp[4]) ? 11'b00100101010 : 11'b00000101010;
										assign node1343 = (inp[4]) ? 11'b00001001000 : 11'b00010001000;
									assign node1346 = (inp[9]) ? 11'b00011100010 : node1347;
										assign node1347 = (inp[11]) ? 11'b00111000000 : 11'b00111100010;
								assign node1351 = (inp[8]) ? node1365 : node1352;
									assign node1352 = (inp[2]) ? node1356 : node1353;
										assign node1353 = (inp[4]) ? 11'b00011100001 : 11'b00000100011;
										assign node1356 = (inp[9]) ? 11'b00000000001 : node1357;
											assign node1357 = (inp[11]) ? node1361 : node1358;
												assign node1358 = (inp[4]) ? 11'b00111100011 : 11'b00000000001;
												assign node1361 = (inp[4]) ? 11'b00011000001 : 11'b00111000001;
									assign node1365 = (inp[9]) ? 11'b00000100000 : 11'b00101100000;
		assign node1368 = (inp[7]) ? node1982 : node1369;
			assign node1369 = (inp[6]) ? node1679 : node1370;
				assign node1370 = (inp[8]) ? node1540 : node1371;
					assign node1371 = (inp[0]) ? node1453 : node1372;
						assign node1372 = (inp[9]) ? node1414 : node1373;
							assign node1373 = (inp[2]) ? node1395 : node1374;
								assign node1374 = (inp[11]) ? node1388 : node1375;
									assign node1375 = (inp[5]) ? node1383 : node1376;
										assign node1376 = (inp[3]) ? node1380 : node1377;
											assign node1377 = (inp[4]) ? 11'b00001101111 : 11'b00001101011;
											assign node1380 = (inp[10]) ? 11'b00001101101 : 11'b10001101001;
										assign node1383 = (inp[3]) ? node1385 : 11'b10011101101;
											assign node1385 = (inp[4]) ? 11'b00011111011 : 11'b00101111111;
									assign node1388 = (inp[5]) ? node1392 : node1389;
										assign node1389 = (inp[10]) ? 11'b00111011001 : 11'b10111001101;
										assign node1392 = (inp[4]) ? 11'b00000011111 : 11'b00011001111;
								assign node1395 = (inp[11]) ? node1405 : node1396;
									assign node1396 = (inp[5]) ? node1398 : 11'b10101001000;
										assign node1398 = (inp[10]) ? node1402 : node1399;
											assign node1399 = (inp[3]) ? 11'b10100011011 : 11'b00101011001;
											assign node1402 = (inp[3]) ? 11'b00000011111 : 11'b10010011001;
									assign node1405 = (inp[5]) ? node1411 : node1406;
										assign node1406 = (inp[10]) ? 11'b10000111111 : node1407;
											assign node1407 = (inp[3]) ? 11'b10110111001 : 11'b00110101101;
										assign node1411 = (inp[3]) ? 11'b00101101101 : 11'b00101111001;
							assign node1414 = (inp[4]) ? node1440 : node1415;
								assign node1415 = (inp[2]) ? node1429 : node1416;
									assign node1416 = (inp[11]) ? node1424 : node1417;
										assign node1417 = (inp[10]) ? node1421 : node1418;
											assign node1418 = (inp[3]) ? 11'b10000101101 : 11'b00000101011;
											assign node1421 = (inp[3]) ? 11'b00010101111 : 11'b10100101101;
										assign node1424 = (inp[3]) ? node1426 : 11'b00100011011;
											assign node1426 = (inp[10]) ? 11'b00000001101 : 11'b10100001101;
									assign node1429 = (inp[5]) ? node1435 : node1430;
										assign node1430 = (inp[11]) ? 11'b00100111111 : node1431;
											assign node1431 = (inp[3]) ? 11'b00110011110 : 11'b10110011100;
										assign node1435 = (inp[3]) ? 11'b10100111101 : node1436;
											assign node1436 = (inp[11]) ? 11'b10010101111 : 11'b10001001111;
								assign node1440 = (inp[3]) ? node1448 : node1441;
									assign node1441 = (inp[10]) ? node1445 : node1442;
										assign node1442 = (inp[2]) ? 11'b00001101111 : 11'b00011001111;
										assign node1445 = (inp[2]) ? 11'b10011011011 : 11'b10100101011;
									assign node1448 = (inp[10]) ? 11'b00110001001 : node1449;
										assign node1449 = (inp[11]) ? 11'b10001101001 : 11'b10100111001;
						assign node1453 = (inp[3]) ? node1491 : node1454;
							assign node1454 = (inp[9]) ? node1476 : node1455;
								assign node1455 = (inp[10]) ? node1469 : node1456;
									assign node1456 = (inp[11]) ? node1462 : node1457;
										assign node1457 = (inp[2]) ? node1459 : 11'b00001101011;
											assign node1459 = (inp[4]) ? 11'b00000001000 : 11'b00000001011;
										assign node1462 = (inp[5]) ? node1466 : node1463;
											assign node1463 = (inp[2]) ? 11'b00010111001 : 11'b00001011011;
											assign node1466 = (inp[4]) ? 11'b00101111011 : 11'b00000111001;
									assign node1469 = (inp[4]) ? 11'b00100101101 : node1470;
										assign node1470 = (inp[11]) ? node1472 : 11'b00001101111;
											assign node1472 = (inp[2]) ? 11'b00001111101 : 11'b00001011111;
								assign node1476 = (inp[11]) ? node1484 : node1477;
									assign node1477 = (inp[2]) ? 11'b00111111011 : node1478;
										assign node1478 = (inp[5]) ? 11'b00100111001 : node1479;
											assign node1479 = (inp[4]) ? 11'b00100111011 : 11'b00000111011;
									assign node1484 = (inp[4]) ? node1488 : node1485;
										assign node1485 = (inp[2]) ? 11'b00111111111 : 11'b00111011101;
										assign node1488 = (inp[10]) ? 11'b00111001011 : 11'b00001001111;
							assign node1491 = (inp[10]) ? node1513 : node1492;
								assign node1492 = (inp[2]) ? node1496 : node1493;
									assign node1493 = (inp[5]) ? 11'b00111111001 : 11'b00001111001;
									assign node1496 = (inp[11]) ? node1506 : node1497;
										assign node1497 = (inp[5]) ? node1503 : node1498;
											assign node1498 = (inp[4]) ? node1500 : 11'b00010011000;
												assign node1500 = (inp[9]) ? 11'b00110101011 : 11'b00011111011;
											assign node1503 = (inp[4]) ? 11'b00010001001 : 11'b00110001001;
										assign node1506 = (inp[5]) ? node1510 : node1507;
											assign node1507 = (inp[4]) ? 11'b00101001001 : 11'b00111111001;
											assign node1510 = (inp[4]) ? 11'b00011111001 : 11'b00000111001;
								assign node1513 = (inp[9]) ? node1533 : node1514;
									assign node1514 = (inp[4]) ? node1524 : node1515;
										assign node1515 = (inp[5]) ? node1519 : node1516;
											assign node1516 = (inp[11]) ? 11'b00101001001 : 11'b00001001000;
											assign node1519 = (inp[2]) ? node1521 : 11'b00001101001;
												assign node1521 = (inp[11]) ? 11'b00110101011 : 11'b00000001011;
										assign node1524 = (inp[11]) ? node1528 : node1525;
											assign node1525 = (inp[2]) ? 11'b00110001001 : 11'b00111101001;
											assign node1528 = (inp[5]) ? node1530 : 11'b00011001011;
												assign node1530 = (inp[2]) ? 11'b00011101011 : 11'b00011001011;
									assign node1533 = (inp[11]) ? node1535 : 11'b00000101001;
										assign node1535 = (inp[4]) ? 11'b00001001001 : node1536;
											assign node1536 = (inp[5]) ? 11'b00000101001 : 11'b00010001001;
					assign node1540 = (inp[0]) ? node1610 : node1541;
						assign node1541 = (inp[11]) ? node1573 : node1542;
							assign node1542 = (inp[5]) ? node1560 : node1543;
								assign node1543 = (inp[9]) ? node1553 : node1544;
									assign node1544 = (inp[3]) ? node1550 : node1545;
										assign node1545 = (inp[2]) ? 11'b00100101011 : node1546;
											assign node1546 = (inp[10]) ? 11'b10100111100 : 11'b00100101100;
										assign node1550 = (inp[4]) ? 11'b00011101010 : 11'b10010101001;
									assign node1553 = (inp[10]) ? node1557 : node1554;
										assign node1554 = (inp[4]) ? 11'b00011001111 : 11'b10001001111;
										assign node1557 = (inp[2]) ? 11'b00010011111 : 11'b10010111110;
								assign node1560 = (inp[10]) ? 11'b00101011010 : node1561;
									assign node1561 = (inp[3]) ? node1565 : node1562;
										assign node1562 = (inp[2]) ? 11'b00100111000 : 11'b00100111110;
										assign node1565 = (inp[4]) ? node1569 : node1566;
											assign node1566 = (inp[2]) ? 11'b10101111100 : 11'b10001111110;
											assign node1569 = (inp[2]) ? 11'b10100111110 : 11'b10010111110;
							assign node1573 = (inp[3]) ? node1597 : node1574;
								assign node1574 = (inp[10]) ? node1588 : node1575;
									assign node1575 = (inp[4]) ? node1583 : node1576;
										assign node1576 = (inp[5]) ? node1580 : node1577;
											assign node1577 = (inp[2]) ? 11'b00101001001 : 11'b00111011000;
											assign node1580 = (inp[2]) ? 11'b00100001000 : 11'b00000101000;
										assign node1583 = (inp[9]) ? node1585 : 11'b00001011110;
											assign node1585 = (inp[5]) ? 11'b00100001110 : 11'b00100111110;
									assign node1588 = (inp[2]) ? node1590 : 11'b10110101100;
										assign node1590 = (inp[5]) ? node1594 : node1591;
											assign node1591 = (inp[9]) ? 11'b10111111110 : 11'b10000001011;
											assign node1594 = (inp[4]) ? 11'b10001001100 : 11'b10001001110;
								assign node1597 = (inp[10]) ? node1605 : node1598;
									assign node1598 = (inp[9]) ? node1602 : node1599;
										assign node1599 = (inp[5]) ? 11'b10011011100 : 11'b10010001100;
										assign node1602 = (inp[2]) ? 11'b10110111000 : 11'b10011011000;
									assign node1605 = (inp[5]) ? node1607 : 11'b00110011101;
										assign node1607 = (inp[4]) ? 11'b00110001000 : 11'b00111001110;
						assign node1610 = (inp[3]) ? node1642 : node1611;
							assign node1611 = (inp[2]) ? node1629 : node1612;
								assign node1612 = (inp[11]) ? node1622 : node1613;
									assign node1613 = (inp[4]) ? node1617 : node1614;
										assign node1614 = (inp[5]) ? 11'b00100001010 : 11'b00111101110;
										assign node1617 = (inp[10]) ? 11'b00001111000 : node1618;
											assign node1618 = (inp[9]) ? 11'b00011111110 : 11'b00011101000;
									assign node1622 = (inp[9]) ? node1624 : 11'b00001011000;
										assign node1624 = (inp[5]) ? node1626 : 11'b00001011100;
											assign node1626 = (inp[4]) ? 11'b00000001100 : 11'b00000111110;
								assign node1629 = (inp[4]) ? node1639 : node1630;
									assign node1630 = (inp[5]) ? 11'b00101101100 : node1631;
										assign node1631 = (inp[11]) ? 11'b00111011001 : node1632;
											assign node1632 = (inp[9]) ? 11'b00111011001 : node1633;
												assign node1633 = (inp[10]) ? 11'b00101001111 : 11'b00100101011;
									assign node1639 = (inp[10]) ? 11'b00111011110 : 11'b00001011111;
							assign node1642 = (inp[10]) ? node1666 : node1643;
								assign node1643 = (inp[4]) ? node1657 : node1644;
									assign node1644 = (inp[9]) ? node1650 : node1645;
										assign node1645 = (inp[2]) ? 11'b00010101001 : node1646;
											assign node1646 = (inp[5]) ? 11'b00100001000 : 11'b00000001001;
										assign node1650 = (inp[2]) ? 11'b00001011010 : node1651;
											assign node1651 = (inp[11]) ? 11'b00010111000 : node1652;
												assign node1652 = (inp[5]) ? 11'b00101111010 : 11'b00011111000;
									assign node1657 = (inp[9]) ? node1659 : 11'b00101111010;
										assign node1659 = (inp[5]) ? 11'b00001001010 : node1660;
											assign node1660 = (inp[11]) ? node1662 : 11'b00101001001;
												assign node1662 = (inp[2]) ? 11'b00100101000 : 11'b00111001000;
								assign node1666 = (inp[11]) ? node1672 : node1667;
									assign node1667 = (inp[5]) ? 11'b00001001000 : node1668;
										assign node1668 = (inp[2]) ? 11'b00000001011 : 11'b00000101000;
									assign node1672 = (inp[4]) ? node1676 : node1673;
										assign node1673 = (inp[5]) ? 11'b00100001010 : 11'b00111001010;
										assign node1676 = (inp[2]) ? 11'b00000101010 : 11'b00000001000;
				assign node1679 = (inp[0]) ? node1813 : node1680;
					assign node1680 = (inp[2]) ? node1750 : node1681;
						assign node1681 = (inp[8]) ? node1715 : node1682;
							assign node1682 = (inp[11]) ? node1702 : node1683;
								assign node1683 = (inp[4]) ? node1691 : node1684;
									assign node1684 = (inp[10]) ? node1688 : node1685;
										assign node1685 = (inp[5]) ? 11'b10011011010 : 11'b00001101010;
										assign node1688 = (inp[3]) ? 11'b00000001110 : 11'b10000111110;
									assign node1691 = (inp[5]) ? 11'b10001110001 : node1692;
										assign node1692 = (inp[9]) ? node1694 : 11'b10010101100;
											assign node1694 = (inp[3]) ? node1698 : node1695;
												assign node1695 = (inp[10]) ? 11'b10101101010 : 11'b00101101100;
												assign node1698 = (inp[10]) ? 11'b00111111000 : 11'b10111111010;
								assign node1702 = (inp[5]) ? node1704 : 11'b00000011110;
									assign node1704 = (inp[9]) ? node1708 : node1705;
										assign node1705 = (inp[10]) ? 11'b10110110011 : 11'b00011110001;
										assign node1708 = (inp[3]) ? 11'b00011100111 : node1709;
											assign node1709 = (inp[10]) ? node1711 : 11'b00110100011;
												assign node1711 = (inp[4]) ? 11'b10000100011 : 11'b10100100101;
							assign node1715 = (inp[5]) ? node1737 : node1716;
								assign node1716 = (inp[11]) ? node1728 : node1717;
									assign node1717 = (inp[4]) ? node1723 : node1718;
										assign node1718 = (inp[3]) ? node1720 : 11'b10010100001;
											assign node1720 = (inp[9]) ? 11'b10101000101 : 11'b00101000111;
										assign node1723 = (inp[3]) ? 11'b10010010001 : node1724;
											assign node1724 = (inp[9]) ? 11'b00110000111 : 11'b10110010101;
									assign node1728 = (inp[4]) ? node1732 : node1729;
										assign node1729 = (inp[10]) ? 11'b10010010101 : 11'b00011000001;
										assign node1732 = (inp[10]) ? 11'b00111110001 : node1733;
											assign node1733 = (inp[3]) ? 11'b10001110001 : 11'b00011110101;
								assign node1737 = (inp[11]) ? node1747 : node1738;
									assign node1738 = (inp[4]) ? node1742 : node1739;
										assign node1739 = (inp[10]) ? 11'b10110110001 : 11'b00001110001;
										assign node1742 = (inp[10]) ? node1744 : 11'b10011110101;
											assign node1744 = (inp[3]) ? 11'b00001110011 : 11'b10001100111;
									assign node1747 = (inp[9]) ? 11'b10100000011 : 11'b10110000111;
						assign node1750 = (inp[8]) ? node1792 : node1751;
							assign node1751 = (inp[4]) ? node1775 : node1752;
								assign node1752 = (inp[9]) ? node1764 : node1753;
									assign node1753 = (inp[11]) ? node1759 : node1754;
										assign node1754 = (inp[10]) ? 11'b10000110010 : node1755;
											assign node1755 = (inp[3]) ? 11'b10100110010 : 11'b00101110000;
										assign node1759 = (inp[5]) ? node1761 : 11'b10101100000;
											assign node1761 = (inp[10]) ? 11'b00100000110 : 11'b00110010000;
									assign node1764 = (inp[5]) ? node1772 : node1765;
										assign node1765 = (inp[11]) ? 11'b10000110100 : node1766;
											assign node1766 = (inp[10]) ? node1768 : 11'b10101000101;
												assign node1768 = (inp[3]) ? 11'b00110010111 : 11'b10110010111;
										assign node1772 = (inp[3]) ? 11'b00100100100 : 11'b10000100100;
								assign node1775 = (inp[9]) ? node1783 : node1776;
									assign node1776 = (inp[10]) ? node1780 : node1777;
										assign node1777 = (inp[5]) ? 11'b00101010100 : 11'b10100000101;
										assign node1780 = (inp[5]) ? 11'b10111000100 : 11'b10011110110;
									assign node1783 = (inp[5]) ? node1787 : node1784;
										assign node1784 = (inp[11]) ? 11'b10111110010 : 11'b00011110000;
										assign node1787 = (inp[3]) ? node1789 : 11'b10110000000;
											assign node1789 = (inp[11]) ? 11'b10010000010 : 11'b00010000010;
							assign node1792 = (inp[5]) ? node1804 : node1793;
								assign node1793 = (inp[11]) ? node1797 : node1794;
									assign node1794 = (inp[3]) ? 11'b10000000010 : 11'b00000100110;
									assign node1797 = (inp[9]) ? node1801 : node1798;
										assign node1798 = (inp[3]) ? 11'b10010110000 : 11'b00110100000;
										assign node1801 = (inp[3]) ? 11'b00001110110 : 11'b10010110010;
								assign node1804 = (inp[10]) ? node1806 : 11'b00101010000;
									assign node1806 = (inp[9]) ? node1808 : 11'b10001010010;
										assign node1808 = (inp[4]) ? node1810 : 11'b10011000100;
											assign node1810 = (inp[11]) ? 11'b10010000000 : 11'b10010010000;
					assign node1813 = (inp[2]) ? node1875 : node1814;
						assign node1814 = (inp[8]) ? node1848 : node1815;
							assign node1815 = (inp[5]) ? node1835 : node1816;
								assign node1816 = (inp[11]) ? node1828 : node1817;
									assign node1817 = (inp[3]) ? node1825 : node1818;
										assign node1818 = (inp[9]) ? node1822 : node1819;
											assign node1819 = (inp[10]) ? 11'b00011111110 : 11'b00010101010;
											assign node1822 = (inp[10]) ? 11'b00010111000 : 11'b00111111100;
										assign node1825 = (inp[10]) ? 11'b00001101010 : 11'b00000111000;
									assign node1828 = (inp[3]) ? node1830 : 11'b00101001100;
										assign node1830 = (inp[4]) ? node1832 : 11'b00100101010;
											assign node1832 = (inp[9]) ? 11'b00110001010 : 11'b00111011000;
								assign node1835 = (inp[11]) ? node1839 : node1836;
									assign node1836 = (inp[10]) ? 11'b00111001100 : 11'b00101001010;
									assign node1839 = (inp[9]) ? 11'b00100100001 : node1840;
										assign node1840 = (inp[10]) ? 11'b00011100001 : node1841;
											assign node1841 = (inp[3]) ? node1843 : 11'b00011110001;
												assign node1843 = (inp[4]) ? 11'b00001110001 : 11'b00100100011;
							assign node1848 = (inp[10]) ? node1860 : node1849;
								assign node1849 = (inp[11]) ? node1853 : node1850;
									assign node1850 = (inp[4]) ? 11'b00110000011 : 11'b00100100111;
									assign node1853 = (inp[4]) ? node1857 : node1854;
										assign node1854 = (inp[5]) ? 11'b00110110011 : 11'b00010010111;
										assign node1857 = (inp[5]) ? 11'b00011010001 : 11'b00111100101;
								assign node1860 = (inp[4]) ? node1870 : node1861;
									assign node1861 = (inp[3]) ? node1865 : node1862;
										assign node1862 = (inp[5]) ? 11'b00011110011 : 11'b00101010011;
										assign node1865 = (inp[9]) ? node1867 : 11'b00101000011;
											assign node1867 = (inp[11]) ? 11'b00010000011 : 11'b00001000001;
									assign node1870 = (inp[9]) ? node1872 : 11'b00000000111;
										assign node1872 = (inp[3]) ? 11'b00001000011 : 11'b00001100011;
						assign node1875 = (inp[5]) ? node1939 : node1876;
							assign node1876 = (inp[11]) ? node1910 : node1877;
								assign node1877 = (inp[8]) ? node1895 : node1878;
									assign node1878 = (inp[10]) ? node1888 : node1879;
										assign node1879 = (inp[9]) ? node1883 : node1880;
											assign node1880 = (inp[4]) ? 11'b00010000001 : 11'b00011000011;
											assign node1883 = (inp[4]) ? node1885 : 11'b00011010001;
												assign node1885 = (inp[3]) ? 11'b00111100010 : 11'b00111110110;
										assign node1888 = (inp[9]) ? node1892 : node1889;
											assign node1889 = (inp[4]) ? 11'b00000010111 : 11'b00001000101;
											assign node1892 = (inp[3]) ? 11'b00000000011 : 11'b00000010011;
									assign node1895 = (inp[9]) ? node1901 : node1896;
										assign node1896 = (inp[3]) ? 11'b00011100010 : node1897;
											assign node1897 = (inp[10]) ? 11'b00110000100 : 11'b00111100000;
										assign node1901 = (inp[4]) ? node1907 : node1902;
											assign node1902 = (inp[3]) ? node1904 : 11'b00101110000;
												assign node1904 = (inp[10]) ? 11'b00001100010 : 11'b00001110000;
											assign node1907 = (inp[3]) ? 11'b00000100010 : 11'b00000110010;
								assign node1910 = (inp[9]) ? node1926 : node1911;
									assign node1911 = (inp[10]) ? 11'b00000100000 : node1912;
										assign node1912 = (inp[3]) ? node1920 : node1913;
											assign node1913 = (inp[8]) ? node1917 : node1914;
												assign node1914 = (inp[4]) ? 11'b00000110000 : 11'b00001110010;
												assign node1917 = (inp[4]) ? 11'b00101110000 : 11'b00100110000;
											assign node1920 = (inp[4]) ? node1922 : 11'b00000100000;
												assign node1922 = (inp[8]) ? 11'b00100110010 : 11'b00100110000;
									assign node1926 = (inp[10]) ? node1932 : node1927;
										assign node1927 = (inp[3]) ? 11'b00110110000 : node1928;
											assign node1928 = (inp[8]) ? 11'b00011110100 : 11'b00011100100;
										assign node1932 = (inp[4]) ? node1936 : node1933;
											assign node1933 = (inp[3]) ? 11'b00011100000 : 11'b00111100010;
											assign node1936 = (inp[3]) ? 11'b00000100000 : 11'b00000100010;
							assign node1939 = (inp[10]) ? node1967 : node1940;
								assign node1940 = (inp[11]) ? node1954 : node1941;
									assign node1941 = (inp[4]) ? node1949 : node1942;
										assign node1942 = (inp[8]) ? node1946 : node1943;
											assign node1943 = (inp[9]) ? 11'b00110110000 : 11'b00010100010;
											assign node1946 = (inp[3]) ? 11'b00111010010 : 11'b00111000010;
										assign node1949 = (inp[3]) ? node1951 : 11'b00111010100;
											assign node1951 = (inp[8]) ? 11'b00100010010 : 11'b00101010000;
									assign node1954 = (inp[3]) ? node1958 : node1955;
										assign node1955 = (inp[4]) ? 11'b00111010010 : 11'b00000010000;
										assign node1958 = (inp[4]) ? node1962 : node1959;
											assign node1959 = (inp[9]) ? 11'b00001010010 : 11'b00101000010;
											assign node1962 = (inp[9]) ? 11'b00000000010 : node1963;
												assign node1963 = (inp[8]) ? 11'b00000010010 : 11'b00011010010;
								assign node1967 = (inp[11]) ? node1973 : node1968;
									assign node1968 = (inp[3]) ? node1970 : 11'b00110110000;
										assign node1970 = (inp[8]) ? 11'b00100000000 : 11'b00000000010;
									assign node1973 = (inp[4]) ? node1977 : node1974;
										assign node1974 = (inp[8]) ? 11'b00001000000 : 11'b00101000010;
										assign node1977 = (inp[8]) ? 11'b00000000000 : node1978;
											assign node1978 = (inp[9]) ? 11'b00000000000 : 11'b00011000000;
			assign node1982 = (inp[6]) ? node2336 : node1983;
				assign node1983 = (inp[2]) ? node2141 : node1984;
					assign node1984 = (inp[5]) ? node2060 : node1985;
						assign node1985 = (inp[10]) ? node2023 : node1986;
							assign node1986 = (inp[0]) ? node2008 : node1987;
								assign node1987 = (inp[11]) ? node1999 : node1988;
									assign node1988 = (inp[4]) ? node1996 : node1989;
										assign node1989 = (inp[8]) ? node1993 : node1990;
											assign node1990 = (inp[3]) ? 11'b10011100111 : 11'b00011100011;
											assign node1993 = (inp[3]) ? 11'b10110000011 : 11'b00010000011;
										assign node1996 = (inp[8]) ? 11'b00111100101 : 11'b00110100111;
									assign node1999 = (inp[8]) ? node2003 : node2000;
										assign node2000 = (inp[4]) ? 11'b00001100101 : 11'b00011100011;
										assign node2003 = (inp[4]) ? node2005 : 11'b00100110011;
											assign node2005 = (inp[3]) ? 11'b10001110011 : 11'b00011110111;
								assign node2008 = (inp[9]) ? node2018 : node2009;
									assign node2009 = (inp[8]) ? node2015 : node2010;
										assign node2010 = (inp[4]) ? node2012 : 11'b00001100011;
											assign node2012 = (inp[3]) ? 11'b00000110011 : 11'b00000100011;
										assign node2015 = (inp[3]) ? 11'b00010100001 : 11'b00111110011;
									assign node2018 = (inp[3]) ? 11'b00100100011 : node2019;
										assign node2019 = (inp[11]) ? 11'b00101110111 : 11'b00100110111;
							assign node2023 = (inp[8]) ? node2043 : node2024;
								assign node2024 = (inp[4]) ? node2032 : node2025;
									assign node2025 = (inp[0]) ? 11'b00011100001 : node2026;
										assign node2026 = (inp[9]) ? node2028 : 11'b10011100001;
											assign node2028 = (inp[11]) ? 11'b10111110101 : 11'b00011110101;
									assign node2032 = (inp[0]) ? node2038 : node2033;
										assign node2033 = (inp[11]) ? node2035 : 11'b10010110101;
											assign node2035 = (inp[3]) ? 11'b00100110001 : 11'b10100110011;
										assign node2038 = (inp[3]) ? 11'b00000100001 : node2039;
											assign node2039 = (inp[11]) ? 11'b00110100001 : 11'b00100110001;
								assign node2043 = (inp[0]) ? node2053 : node2044;
									assign node2044 = (inp[11]) ? node2050 : node2045;
										assign node2045 = (inp[9]) ? 11'b10001110111 : node2046;
											assign node2046 = (inp[3]) ? 11'b00001100011 : 11'b10010000001;
										assign node2050 = (inp[9]) ? 11'b00111110111 : 11'b00000110111;
									assign node2053 = (inp[9]) ? node2057 : node2054;
										assign node2054 = (inp[11]) ? 11'b00001100101 : 11'b00101110111;
										assign node2057 = (inp[3]) ? 11'b00001100001 : 11'b00011100001;
						assign node2060 = (inp[11]) ? node2096 : node2061;
							assign node2061 = (inp[8]) ? node2075 : node2062;
								assign node2062 = (inp[3]) ? node2068 : node2063;
									assign node2063 = (inp[0]) ? 11'b00110010101 : node2064;
										assign node2064 = (inp[9]) ? 11'b00011010001 : 11'b00001010101;
									assign node2068 = (inp[4]) ? node2072 : node2069;
										assign node2069 = (inp[9]) ? 11'b00101010011 : 11'b00101000011;
										assign node2072 = (inp[0]) ? 11'b00110000001 : 11'b00000010011;
								assign node2075 = (inp[4]) ? node2089 : node2076;
									assign node2076 = (inp[9]) ? node2082 : node2077;
										assign node2077 = (inp[10]) ? 11'b00010100001 : node2078;
											assign node2078 = (inp[3]) ? 11'b10010110011 : 11'b00011110001;
										assign node2082 = (inp[10]) ? node2086 : node2083;
											assign node2083 = (inp[0]) ? 11'b00100110001 : 11'b00000110001;
											assign node2086 = (inp[3]) ? 11'b00010100011 : 11'b00000110011;
									assign node2089 = (inp[0]) ? node2091 : 11'b00111010111;
										assign node2091 = (inp[9]) ? node2093 : 11'b00110110001;
											assign node2093 = (inp[10]) ? 11'b00001000001 : 11'b00011000001;
							assign node2096 = (inp[4]) ? node2126 : node2097;
								assign node2097 = (inp[10]) ? node2109 : node2098;
									assign node2098 = (inp[9]) ? node2102 : node2099;
										assign node2099 = (inp[0]) ? 11'b00101010011 : 11'b00011010011;
										assign node2102 = (inp[0]) ? node2106 : node2103;
											assign node2103 = (inp[8]) ? 11'b00011000001 : 11'b00101000011;
											assign node2106 = (inp[3]) ? 11'b00011010001 : 11'b00111010101;
									assign node2109 = (inp[9]) ? node2115 : node2110;
										assign node2110 = (inp[3]) ? 11'b00011000101 : node2111;
											assign node2111 = (inp[0]) ? 11'b00011010111 : 11'b10001010011;
										assign node2115 = (inp[0]) ? node2121 : node2116;
											assign node2116 = (inp[8]) ? node2118 : 11'b10101000101;
												assign node2118 = (inp[3]) ? 11'b00100000111 : 11'b10100000111;
											assign node2121 = (inp[3]) ? node2123 : 11'b00111000011;
												assign node2123 = (inp[8]) ? 11'b00000000011 : 11'b00001000011;
								assign node2126 = (inp[3]) ? node2136 : node2127;
									assign node2127 = (inp[8]) ? node2131 : node2128;
										assign node2128 = (inp[9]) ? 11'b00110000001 : 11'b00101000101;
										assign node2131 = (inp[0]) ? node2133 : 11'b00110010101;
											assign node2133 = (inp[10]) ? 11'b00010000111 : 11'b00000000111;
									assign node2136 = (inp[0]) ? node2138 : 11'b10110000001;
										assign node2138 = (inp[10]) ? 11'b00000000001 : 11'b00010000001;
					assign node2141 = (inp[0]) ? node2239 : node2142;
						assign node2142 = (inp[8]) ? node2188 : node2143;
							assign node2143 = (inp[5]) ? node2167 : node2144;
								assign node2144 = (inp[11]) ? node2156 : node2145;
									assign node2145 = (inp[4]) ? node2153 : node2146;
										assign node2146 = (inp[10]) ? node2150 : node2147;
											assign node2147 = (inp[9]) ? 11'b10111000111 : 11'b00111000011;
											assign node2150 = (inp[9]) ? 11'b00101010111 : 11'b00101000101;
										assign node2153 = (inp[10]) ? 11'b10000000001 : 11'b10000010011;
									assign node2156 = (inp[10]) ? node2164 : node2157;
										assign node2157 = (inp[4]) ? node2161 : node2158;
											assign node2158 = (inp[9]) ? 11'b00000010001 : 11'b00110000011;
											assign node2161 = (inp[3]) ? 11'b10111110010 : 11'b00101100110;
										assign node2164 = (inp[3]) ? 11'b00111110110 : 11'b10011110110;
								assign node2167 = (inp[11]) ? node2177 : node2168;
									assign node2168 = (inp[10]) ? node2174 : node2169;
										assign node2169 = (inp[3]) ? 11'b10110110010 : node2170;
											assign node2170 = (inp[9]) ? 11'b00010110100 : 11'b00100110110;
										assign node2174 = (inp[9]) ? 11'b10101110010 : 11'b10110100100;
									assign node2177 = (inp[9]) ? node2185 : node2178;
										assign node2178 = (inp[10]) ? node2182 : node2179;
											assign node2179 = (inp[3]) ? 11'b10001110100 : 11'b00111110100;
											assign node2182 = (inp[3]) ? 11'b00010100010 : 11'b10011110000;
										assign node2185 = (inp[4]) ? 11'b00100100110 : 11'b00101100100;
							assign node2188 = (inp[11]) ? node2212 : node2189;
								assign node2189 = (inp[3]) ? node2207 : node2190;
									assign node2190 = (inp[10]) ? node2198 : node2191;
										assign node2191 = (inp[4]) ? 11'b00011000110 : node2192;
											assign node2192 = (inp[5]) ? node2194 : 11'b00110100010;
												assign node2194 = (inp[9]) ? 11'b00101010010 : 11'b00110010000;
										assign node2198 = (inp[4]) ? node2204 : node2199;
											assign node2199 = (inp[5]) ? 11'b10011010010 : node2200;
												assign node2200 = (inp[9]) ? 11'b10111010110 : 11'b10100100010;
											assign node2204 = (inp[5]) ? 11'b10101000110 : 11'b10101000010;
									assign node2207 = (inp[10]) ? node2209 : 11'b10011000000;
										assign node2209 = (inp[5]) ? 11'b00001010110 : 11'b00011010010;
								assign node2212 = (inp[10]) ? node2224 : node2213;
									assign node2213 = (inp[3]) ? node2217 : node2214;
										assign node2214 = (inp[4]) ? 11'b00000000100 : 11'b00110010010;
										assign node2217 = (inp[4]) ? node2221 : node2218;
											assign node2218 = (inp[9]) ? 11'b10000000110 : 11'b10100000010;
											assign node2221 = (inp[9]) ? 11'b10100010010 : 11'b10000010110;
									assign node2224 = (inp[3]) ? node2234 : node2225;
										assign node2225 = (inp[5]) ? node2231 : node2226;
											assign node2226 = (inp[9]) ? 11'b10100010110 : node2227;
												assign node2227 = (inp[4]) ? 11'b10000010100 : 11'b10011000000;
											assign node2231 = (inp[9]) ? 11'b10010000100 : 11'b10010000110;
										assign node2234 = (inp[5]) ? 11'b00100000110 : node2235;
											assign node2235 = (inp[4]) ? 11'b00000010000 : 11'b00010010100;
						assign node2239 = (inp[8]) ? node2293 : node2240;
							assign node2240 = (inp[5]) ? node2268 : node2241;
								assign node2241 = (inp[11]) ? node2259 : node2242;
									assign node2242 = (inp[4]) ? node2248 : node2243;
										assign node2243 = (inp[3]) ? 11'b00001000011 : node2244;
											assign node2244 = (inp[10]) ? 11'b00011010011 : 11'b00001000011;
										assign node2248 = (inp[10]) ? node2252 : node2249;
											assign node2249 = (inp[3]) ? 11'b00011010001 : 11'b00001000001;
											assign node2252 = (inp[3]) ? node2256 : node2253;
												assign node2253 = (inp[9]) ? 11'b00110010001 : 11'b00010010111;
												assign node2256 = (inp[9]) ? 11'b00000000001 : 11'b00100000011;
									assign node2259 = (inp[3]) ? node2263 : node2260;
										assign node2260 = (inp[4]) ? 11'b00001100110 : 11'b00001100010;
										assign node2263 = (inp[4]) ? 11'b00011100010 : node2264;
											assign node2264 = (inp[10]) ? 11'b00100000001 : 11'b00010000011;
								assign node2268 = (inp[3]) ? node2280 : node2269;
									assign node2269 = (inp[10]) ? node2273 : node2270;
										assign node2270 = (inp[11]) ? 11'b00101110000 : 11'b00001100000;
										assign node2273 = (inp[9]) ? node2275 : 11'b00110100110;
											assign node2275 = (inp[11]) ? node2277 : 11'b00111110010;
												assign node2277 = (inp[4]) ? 11'b00110100000 : 11'b00111100000;
									assign node2280 = (inp[9]) ? node2286 : node2281;
										assign node2281 = (inp[11]) ? 11'b00010110010 : node2282;
											assign node2282 = (inp[4]) ? 11'b00100110010 : 11'b00000100010;
										assign node2286 = (inp[11]) ? 11'b00001110010 : node2287;
											assign node2287 = (inp[4]) ? node2289 : 11'b00010100010;
												assign node2289 = (inp[10]) ? 11'b00001100010 : 11'b00011100010;
							assign node2293 = (inp[11]) ? node2315 : node2294;
								assign node2294 = (inp[3]) ? node2300 : node2295;
									assign node2295 = (inp[4]) ? node2297 : 11'b00101000110;
										assign node2297 = (inp[5]) ? 11'b00001000000 : 11'b00101000010;
									assign node2300 = (inp[10]) ? node2310 : node2301;
										assign node2301 = (inp[9]) ? node2305 : node2302;
											assign node2302 = (inp[4]) ? 11'b00011010000 : 11'b00010100010;
											assign node2305 = (inp[4]) ? node2307 : 11'b00111010000;
												assign node2307 = (inp[5]) ? 11'b00001000000 : 11'b00101000010;
										assign node2310 = (inp[4]) ? 11'b00101000010 : node2311;
											assign node2311 = (inp[5]) ? 11'b00011000010 : 11'b00001000010;
								assign node2315 = (inp[10]) ? node2325 : node2316;
									assign node2316 = (inp[3]) ? node2320 : node2317;
										assign node2317 = (inp[5]) ? 11'b00010010100 : 11'b00000010110;
										assign node2320 = (inp[5]) ? node2322 : 11'b00001000000;
											assign node2322 = (inp[4]) ? 11'b00000000000 : 11'b00000010000;
									assign node2325 = (inp[4]) ? node2333 : node2326;
										assign node2326 = (inp[5]) ? 11'b00100000010 : node2327;
											assign node2327 = (inp[3]) ? node2329 : 11'b00100000010;
												assign node2329 = (inp[9]) ? 11'b00010000000 : 11'b00110000010;
										assign node2333 = (inp[3]) ? 11'b00000000010 : 11'b00010000110;
				assign node2336 = (inp[2]) ? node2538 : node2337;
					assign node2337 = (inp[8]) ? node2445 : node2338;
						assign node2338 = (inp[11]) ? node2388 : node2339;
							assign node2339 = (inp[0]) ? node2361 : node2340;
								assign node2340 = (inp[3]) ? node2354 : node2341;
									assign node2341 = (inp[10]) ? node2347 : node2342;
										assign node2342 = (inp[5]) ? node2344 : 11'b00111100100;
											assign node2344 = (inp[4]) ? 11'b00001110100 : 11'b00001110010;
										assign node2347 = (inp[5]) ? node2351 : node2348;
											assign node2348 = (inp[4]) ? 11'b10111100000 : 11'b10011110100;
											assign node2351 = (inp[9]) ? 11'b10101100110 : 11'b10111110010;
									assign node2354 = (inp[9]) ? 11'b00011100100 : node2355;
										assign node2355 = (inp[5]) ? 11'b00101110110 : node2356;
											assign node2356 = (inp[4]) ? 11'b10001100110 : 11'b00001100110;
								assign node2361 = (inp[3]) ? node2373 : node2362;
									assign node2362 = (inp[9]) ? node2366 : node2363;
										assign node2363 = (inp[5]) ? 11'b00111100110 : 11'b00011100110;
										assign node2366 = (inp[10]) ? node2368 : 11'b00011100110;
											assign node2368 = (inp[5]) ? node2370 : 11'b00111110000;
												assign node2370 = (inp[4]) ? 11'b00111110010 : 11'b00111110000;
									assign node2373 = (inp[10]) ? node2381 : node2374;
										assign node2374 = (inp[9]) ? node2378 : node2375;
											assign node2375 = (inp[4]) ? 11'b00111110000 : 11'b00100100000;
											assign node2378 = (inp[4]) ? 11'b00101100000 : 11'b00001110000;
										assign node2381 = (inp[9]) ? node2385 : node2382;
											assign node2382 = (inp[5]) ? 11'b00111100010 : 11'b00101100010;
											assign node2385 = (inp[5]) ? 11'b00001100010 : 11'b00001100000;
							assign node2388 = (inp[9]) ? node2418 : node2389;
								assign node2389 = (inp[10]) ? node2403 : node2390;
									assign node2390 = (inp[3]) ? node2400 : node2391;
										assign node2391 = (inp[5]) ? node2397 : node2392;
											assign node2392 = (inp[0]) ? node2394 : 11'b00001100000;
												assign node2394 = (inp[4]) ? 11'b00000110000 : 11'b00010110010;
											assign node2397 = (inp[4]) ? 11'b00010110110 : 11'b00011110000;
										assign node2400 = (inp[4]) ? 11'b00000110010 : 11'b10010110010;
									assign node2403 = (inp[5]) ? node2413 : node2404;
										assign node2404 = (inp[4]) ? node2410 : node2405;
											assign node2405 = (inp[0]) ? node2407 : 11'b00010110110;
												assign node2407 = (inp[3]) ? 11'b00100100010 : 11'b00010110110;
											assign node2410 = (inp[0]) ? 11'b00100100110 : 11'b10100110110;
										assign node2413 = (inp[4]) ? node2415 : 11'b00011100100;
											assign node2415 = (inp[0]) ? 11'b00010100000 : 11'b00110100000;
								assign node2418 = (inp[5]) ? node2434 : node2419;
									assign node2419 = (inp[3]) ? node2427 : node2420;
										assign node2420 = (inp[10]) ? node2424 : node2421;
											assign node2421 = (inp[0]) ? 11'b00110110100 : 11'b00100110010;
											assign node2424 = (inp[4]) ? 11'b10110110000 : 11'b10100110100;
										assign node2427 = (inp[4]) ? node2429 : 11'b00100110000;
											assign node2429 = (inp[0]) ? node2431 : 11'b00100110000;
												assign node2431 = (inp[10]) ? 11'b00000100000 : 11'b00110100000;
									assign node2434 = (inp[4]) ? node2436 : 11'b00000100110;
										assign node2436 = (inp[3]) ? node2440 : node2437;
											assign node2437 = (inp[0]) ? 11'b00100100100 : 11'b00000100100;
											assign node2440 = (inp[10]) ? node2442 : 11'b10110100000;
												assign node2442 = (inp[0]) ? 11'b00000100000 : 11'b00100100000;
						assign node2445 = (inp[5]) ? node2491 : node2446;
							assign node2446 = (inp[11]) ? node2468 : node2447;
								assign node2447 = (inp[4]) ? node2459 : node2448;
									assign node2448 = (inp[0]) ? 11'b00100110000 : node2449;
										assign node2449 = (inp[3]) ? node2455 : node2450;
											assign node2450 = (inp[10]) ? 11'b10000100010 : node2451;
												assign node2451 = (inp[9]) ? 11'b00000100010 : 11'b00010100010;
											assign node2455 = (inp[10]) ? 11'b00110100110 : 11'b10100100010;
									assign node2459 = (inp[9]) ? node2463 : node2460;
										assign node2460 = (inp[10]) ? 11'b00111010110 : 11'b00110100100;
										assign node2463 = (inp[3]) ? node2465 : 11'b00011010010;
											assign node2465 = (inp[10]) ? 11'b00101010010 : 11'b10001010010;
								assign node2468 = (inp[0]) ? node2482 : node2469;
									assign node2469 = (inp[9]) ? node2475 : node2470;
										assign node2470 = (inp[4]) ? node2472 : 11'b10111010000;
											assign node2472 = (inp[10]) ? 11'b10111010110 : 11'b10001000110;
										assign node2475 = (inp[3]) ? node2479 : node2476;
											assign node2476 = (inp[4]) ? 11'b10101010000 : 11'b00111010000;
											assign node2479 = (inp[4]) ? 11'b00101010000 : 11'b10101000100;
									assign node2482 = (inp[10]) ? node2488 : node2483;
										assign node2483 = (inp[9]) ? node2485 : 11'b00111010000;
											assign node2485 = (inp[3]) ? 11'b00111000000 : 11'b00111000100;
										assign node2488 = (inp[3]) ? 11'b00111000000 : 11'b00001000000;
							assign node2491 = (inp[10]) ? node2507 : node2492;
								assign node2492 = (inp[11]) ? node2496 : node2493;
									assign node2493 = (inp[3]) ? 11'b10011010000 : 11'b00111000000;
									assign node2496 = (inp[0]) ? node2500 : node2497;
										assign node2497 = (inp[3]) ? 11'b10110010100 : 11'b00000010000;
										assign node2500 = (inp[4]) ? 11'b00010010000 : node2501;
											assign node2501 = (inp[9]) ? node2503 : 11'b00110010010;
												assign node2503 = (inp[3]) ? 11'b00010010010 : 11'b00010010110;
								assign node2507 = (inp[4]) ? node2525 : node2508;
									assign node2508 = (inp[3]) ? node2518 : node2509;
										assign node2509 = (inp[0]) ? 11'b00010010010 : node2510;
											assign node2510 = (inp[9]) ? node2514 : node2511;
												assign node2511 = (inp[11]) ? 11'b10010010010 : 11'b10101010000;
												assign node2514 = (inp[11]) ? 11'b10100000110 : 11'b10000000110;
										assign node2518 = (inp[11]) ? node2520 : 11'b00110010110;
											assign node2520 = (inp[0]) ? node2522 : 11'b00100000110;
												assign node2522 = (inp[9]) ? 11'b00000000010 : 11'b00100000010;
									assign node2525 = (inp[3]) ? node2531 : node2526;
										assign node2526 = (inp[9]) ? 11'b00000000000 : node2527;
											assign node2527 = (inp[11]) ? 11'b10100000100 : 11'b10010000100;
										assign node2531 = (inp[11]) ? node2535 : node2532;
											assign node2532 = (inp[9]) ? 11'b00100000000 : 11'b00010010000;
											assign node2535 = (inp[0]) ? 11'b00000000000 : 11'b00100000000;
					assign node2538 = (inp[0]) ? node2594 : node2539;
						assign node2539 = (inp[11]) ? node2571 : node2540;
							assign node2540 = (inp[4]) ? node2554 : node2541;
								assign node2541 = (inp[10]) ? node2549 : node2542;
									assign node2542 = (inp[8]) ? node2546 : node2543;
										assign node2543 = (inp[3]) ? 11'b10111010000 : 11'b00111010000;
										assign node2546 = (inp[3]) ? 11'b10110010000 : 11'b00110010000;
									assign node2549 = (inp[9]) ? node2551 : 11'b10010010000;
										assign node2551 = (inp[8]) ? 11'b00010000100 : 11'b00110000110;
								assign node2554 = (inp[8]) ? node2564 : node2555;
									assign node2555 = (inp[5]) ? node2561 : node2556;
										assign node2556 = (inp[9]) ? 11'b10011010000 : node2557;
											assign node2557 = (inp[10]) ? 11'b10101010100 : 11'b10111000100;
										assign node2561 = (inp[3]) ? 11'b10000010110 : 11'b00100010110;
									assign node2564 = (inp[5]) ? 11'b00000000000 : node2565;
										assign node2565 = (inp[9]) ? 11'b10100010010 : node2566;
											assign node2566 = (inp[10]) ? 11'b00110000010 : 11'b10110000110;
							assign node2571 = (inp[5]) ? node2583 : node2572;
								assign node2572 = (inp[8]) ? node2580 : node2573;
									assign node2573 = (inp[10]) ? node2575 : 11'b10001000110;
										assign node2575 = (inp[9]) ? 11'b00001010000 : node2576;
											assign node2576 = (inp[3]) ? 11'b00101010110 : 11'b10001010110;
									assign node2580 = (inp[9]) ? 11'b00100010100 : 11'b10000010100;
								assign node2583 = (inp[9]) ? node2589 : node2584;
									assign node2584 = (inp[10]) ? 11'b10010010000 : node2585;
										assign node2585 = (inp[8]) ? 11'b00000010100 : 11'b00100010010;
									assign node2589 = (inp[4]) ? node2591 : 11'b10000000100;
										assign node2591 = (inp[8]) ? 11'b10000000000 : 11'b00000000000;
						assign node2594 = (inp[3]) ? node2632 : node2595;
							assign node2595 = (inp[5]) ? node2615 : node2596;
								assign node2596 = (inp[8]) ? node2606 : node2597;
									assign node2597 = (inp[4]) ? node2603 : node2598;
										assign node2598 = (inp[9]) ? node2600 : 11'b00001010000;
											assign node2600 = (inp[10]) ? 11'b00001010010 : 11'b00101010110;
										assign node2603 = (inp[10]) ? 11'b00101010000 : 11'b00011000100;
									assign node2606 = (inp[11]) ? node2610 : node2607;
										assign node2607 = (inp[4]) ? 11'b00010010110 : 11'b00110000010;
										assign node2610 = (inp[10]) ? 11'b00000000000 : node2611;
											assign node2611 = (inp[4]) ? 11'b00100010000 : 11'b00100010010;
								assign node2615 = (inp[11]) ? node2623 : node2616;
									assign node2616 = (inp[9]) ? node2618 : 11'b00110000000;
										assign node2618 = (inp[4]) ? node2620 : 11'b00010010000;
											assign node2620 = (inp[10]) ? 11'b00000010000 : 11'b00000010100;
									assign node2623 = (inp[4]) ? 11'b00110000100 : node2624;
										assign node2624 = (inp[10]) ? node2628 : node2625;
											assign node2625 = (inp[9]) ? 11'b00100010100 : 11'b00000010010;
											assign node2628 = (inp[8]) ? 11'b00100010100 : 11'b00010010100;
							assign node2632 = (inp[11]) ? node2654 : node2633;
								assign node2633 = (inp[10]) ? node2643 : node2634;
									assign node2634 = (inp[9]) ? node2638 : node2635;
										assign node2635 = (inp[8]) ? 11'b00010000010 : 11'b00100010010;
										assign node2638 = (inp[5]) ? 11'b00010000010 : node2639;
											assign node2639 = (inp[8]) ? 11'b00000010010 : 11'b00011010010;
									assign node2643 = (inp[8]) ? 11'b00010000000 : node2644;
										assign node2644 = (inp[4]) ? node2648 : node2645;
											assign node2645 = (inp[5]) ? 11'b00001000000 : 11'b00001000010;
											assign node2648 = (inp[5]) ? node2650 : 11'b00101000000;
												assign node2650 = (inp[9]) ? 11'b00000000010 : 11'b00110000010;
								assign node2654 = (inp[9]) ? node2664 : node2655;
									assign node2655 = (inp[4]) ? node2661 : node2656;
										assign node2656 = (inp[5]) ? node2658 : 11'b00110000000;
											assign node2658 = (inp[8]) ? 11'b00100000000 : 11'b00110000000;
										assign node2661 = (inp[8]) ? 11'b00000000000 : 11'b00010000000;
									assign node2664 = (inp[5]) ? node2668 : node2665;
										assign node2665 = (inp[8]) ? 11'b00000000000 : 11'b00011000010;
										assign node2668 = (inp[10]) ? 11'b00000000000 : 11'b00000010000;

endmodule