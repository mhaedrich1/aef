module dtc_split125_bm25 (
	input  wire [14-1:0] inp,
	output wire [14-1:0] outp
);

	wire [14-1:0] node1;
	wire [14-1:0] node2;
	wire [14-1:0] node3;
	wire [14-1:0] node4;
	wire [14-1:0] node5;
	wire [14-1:0] node6;
	wire [14-1:0] node7;
	wire [14-1:0] node8;
	wire [14-1:0] node9;
	wire [14-1:0] node10;
	wire [14-1:0] node11;
	wire [14-1:0] node15;
	wire [14-1:0] node18;
	wire [14-1:0] node21;
	wire [14-1:0] node22;
	wire [14-1:0] node25;
	wire [14-1:0] node28;
	wire [14-1:0] node29;
	wire [14-1:0] node30;
	wire [14-1:0] node32;
	wire [14-1:0] node33;
	wire [14-1:0] node38;
	wire [14-1:0] node39;
	wire [14-1:0] node40;
	wire [14-1:0] node41;
	wire [14-1:0] node45;
	wire [14-1:0] node46;
	wire [14-1:0] node48;
	wire [14-1:0] node53;
	wire [14-1:0] node54;
	wire [14-1:0] node55;
	wire [14-1:0] node56;
	wire [14-1:0] node57;
	wire [14-1:0] node58;
	wire [14-1:0] node59;
	wire [14-1:0] node64;
	wire [14-1:0] node65;
	wire [14-1:0] node67;
	wire [14-1:0] node71;
	wire [14-1:0] node72;
	wire [14-1:0] node76;
	wire [14-1:0] node77;
	wire [14-1:0] node78;
	wire [14-1:0] node82;
	wire [14-1:0] node84;
	wire [14-1:0] node85;
	wire [14-1:0] node89;
	wire [14-1:0] node90;
	wire [14-1:0] node91;
	wire [14-1:0] node92;
	wire [14-1:0] node95;
	wire [14-1:0] node98;
	wire [14-1:0] node99;
	wire [14-1:0] node101;
	wire [14-1:0] node105;
	wire [14-1:0] node106;
	wire [14-1:0] node109;
	wire [14-1:0] node111;
	wire [14-1:0] node114;
	wire [14-1:0] node115;
	wire [14-1:0] node116;
	wire [14-1:0] node117;
	wire [14-1:0] node118;
	wire [14-1:0] node119;
	wire [14-1:0] node120;
	wire [14-1:0] node123;
	wire [14-1:0] node127;
	wire [14-1:0] node129;
	wire [14-1:0] node130;
	wire [14-1:0] node131;
	wire [14-1:0] node133;
	wire [14-1:0] node138;
	wire [14-1:0] node139;
	wire [14-1:0] node142;
	wire [14-1:0] node143;
	wire [14-1:0] node147;
	wire [14-1:0] node148;
	wire [14-1:0] node149;
	wire [14-1:0] node152;
	wire [14-1:0] node153;
	wire [14-1:0] node157;
	wire [14-1:0] node160;
	wire [14-1:0] node161;
	wire [14-1:0] node162;
	wire [14-1:0] node163;
	wire [14-1:0] node166;
	wire [14-1:0] node168;
	wire [14-1:0] node171;
	wire [14-1:0] node172;
	wire [14-1:0] node174;
	wire [14-1:0] node175;
	wire [14-1:0] node178;
	wire [14-1:0] node181;
	wire [14-1:0] node184;
	wire [14-1:0] node185;
	wire [14-1:0] node187;
	wire [14-1:0] node189;
	wire [14-1:0] node192;
	wire [14-1:0] node195;
	wire [14-1:0] node196;
	wire [14-1:0] node197;
	wire [14-1:0] node198;
	wire [14-1:0] node199;
	wire [14-1:0] node200;
	wire [14-1:0] node201;
	wire [14-1:0] node205;
	wire [14-1:0] node208;
	wire [14-1:0] node209;
	wire [14-1:0] node210;
	wire [14-1:0] node212;
	wire [14-1:0] node215;
	wire [14-1:0] node217;
	wire [14-1:0] node219;
	wire [14-1:0] node222;
	wire [14-1:0] node225;
	wire [14-1:0] node226;
	wire [14-1:0] node227;
	wire [14-1:0] node229;
	wire [14-1:0] node232;
	wire [14-1:0] node235;
	wire [14-1:0] node236;
	wire [14-1:0] node240;
	wire [14-1:0] node241;
	wire [14-1:0] node242;
	wire [14-1:0] node243;
	wire [14-1:0] node245;
	wire [14-1:0] node249;
	wire [14-1:0] node250;
	wire [14-1:0] node252;
	wire [14-1:0] node253;
	wire [14-1:0] node254;
	wire [14-1:0] node256;
	wire [14-1:0] node262;
	wire [14-1:0] node263;
	wire [14-1:0] node264;
	wire [14-1:0] node266;
	wire [14-1:0] node269;
	wire [14-1:0] node270;
	wire [14-1:0] node273;
	wire [14-1:0] node276;
	wire [14-1:0] node277;
	wire [14-1:0] node279;
	wire [14-1:0] node283;
	wire [14-1:0] node284;
	wire [14-1:0] node285;
	wire [14-1:0] node286;
	wire [14-1:0] node287;
	wire [14-1:0] node288;
	wire [14-1:0] node292;
	wire [14-1:0] node293;
	wire [14-1:0] node295;
	wire [14-1:0] node296;
	wire [14-1:0] node298;
	wire [14-1:0] node303;
	wire [14-1:0] node304;
	wire [14-1:0] node305;
	wire [14-1:0] node308;
	wire [14-1:0] node309;
	wire [14-1:0] node313;
	wire [14-1:0] node316;
	wire [14-1:0] node317;
	wire [14-1:0] node320;
	wire [14-1:0] node321;
	wire [14-1:0] node323;
	wire [14-1:0] node324;
	wire [14-1:0] node328;
	wire [14-1:0] node329;
	wire [14-1:0] node333;
	wire [14-1:0] node334;
	wire [14-1:0] node335;
	wire [14-1:0] node336;
	wire [14-1:0] node339;
	wire [14-1:0] node342;
	wire [14-1:0] node343;
	wire [14-1:0] node344;
	wire [14-1:0] node346;
	wire [14-1:0] node350;
	wire [14-1:0] node353;
	wire [14-1:0] node354;
	wire [14-1:0] node355;
	wire [14-1:0] node358;
	wire [14-1:0] node359;
	wire [14-1:0] node361;
	wire [14-1:0] node363;
	wire [14-1:0] node367;
	wire [14-1:0] node368;
	wire [14-1:0] node370;
	wire [14-1:0] node371;
	wire [14-1:0] node372;
	wire [14-1:0] node377;
	wire [14-1:0] node379;
	wire [14-1:0] node380;
	wire [14-1:0] node384;
	wire [14-1:0] node385;
	wire [14-1:0] node386;
	wire [14-1:0] node387;
	wire [14-1:0] node388;
	wire [14-1:0] node389;
	wire [14-1:0] node390;
	wire [14-1:0] node392;
	wire [14-1:0] node395;
	wire [14-1:0] node396;
	wire [14-1:0] node397;
	wire [14-1:0] node402;
	wire [14-1:0] node403;
	wire [14-1:0] node406;
	wire [14-1:0] node409;
	wire [14-1:0] node410;
	wire [14-1:0] node411;
	wire [14-1:0] node412;
	wire [14-1:0] node413;
	wire [14-1:0] node417;
	wire [14-1:0] node420;
	wire [14-1:0] node423;
	wire [14-1:0] node424;
	wire [14-1:0] node426;
	wire [14-1:0] node427;
	wire [14-1:0] node430;
	wire [14-1:0] node433;
	wire [14-1:0] node435;
	wire [14-1:0] node438;
	wire [14-1:0] node439;
	wire [14-1:0] node440;
	wire [14-1:0] node441;
	wire [14-1:0] node444;
	wire [14-1:0] node445;
	wire [14-1:0] node449;
	wire [14-1:0] node450;
	wire [14-1:0] node453;
	wire [14-1:0] node456;
	wire [14-1:0] node457;
	wire [14-1:0] node458;
	wire [14-1:0] node461;
	wire [14-1:0] node462;
	wire [14-1:0] node466;
	wire [14-1:0] node467;
	wire [14-1:0] node469;
	wire [14-1:0] node472;
	wire [14-1:0] node474;
	wire [14-1:0] node477;
	wire [14-1:0] node478;
	wire [14-1:0] node479;
	wire [14-1:0] node480;
	wire [14-1:0] node481;
	wire [14-1:0] node483;
	wire [14-1:0] node486;
	wire [14-1:0] node489;
	wire [14-1:0] node490;
	wire [14-1:0] node491;
	wire [14-1:0] node495;
	wire [14-1:0] node497;
	wire [14-1:0] node498;
	wire [14-1:0] node502;
	wire [14-1:0] node503;
	wire [14-1:0] node504;
	wire [14-1:0] node506;
	wire [14-1:0] node507;
	wire [14-1:0] node511;
	wire [14-1:0] node513;
	wire [14-1:0] node514;
	wire [14-1:0] node518;
	wire [14-1:0] node519;
	wire [14-1:0] node523;
	wire [14-1:0] node524;
	wire [14-1:0] node525;
	wire [14-1:0] node526;
	wire [14-1:0] node528;
	wire [14-1:0] node531;
	wire [14-1:0] node532;
	wire [14-1:0] node536;
	wire [14-1:0] node537;
	wire [14-1:0] node539;
	wire [14-1:0] node542;
	wire [14-1:0] node545;
	wire [14-1:0] node546;
	wire [14-1:0] node547;
	wire [14-1:0] node548;
	wire [14-1:0] node550;
	wire [14-1:0] node554;
	wire [14-1:0] node556;
	wire [14-1:0] node559;
	wire [14-1:0] node560;
	wire [14-1:0] node563;
	wire [14-1:0] node565;
	wire [14-1:0] node568;
	wire [14-1:0] node569;
	wire [14-1:0] node570;
	wire [14-1:0] node571;
	wire [14-1:0] node572;
	wire [14-1:0] node573;
	wire [14-1:0] node574;
	wire [14-1:0] node578;
	wire [14-1:0] node581;
	wire [14-1:0] node582;
	wire [14-1:0] node583;
	wire [14-1:0] node584;
	wire [14-1:0] node589;
	wire [14-1:0] node591;
	wire [14-1:0] node592;
	wire [14-1:0] node593;
	wire [14-1:0] node598;
	wire [14-1:0] node599;
	wire [14-1:0] node600;
	wire [14-1:0] node602;
	wire [14-1:0] node603;
	wire [14-1:0] node607;
	wire [14-1:0] node610;
	wire [14-1:0] node612;
	wire [14-1:0] node615;
	wire [14-1:0] node616;
	wire [14-1:0] node617;
	wire [14-1:0] node618;
	wire [14-1:0] node619;
	wire [14-1:0] node624;
	wire [14-1:0] node625;
	wire [14-1:0] node628;
	wire [14-1:0] node629;
	wire [14-1:0] node631;
	wire [14-1:0] node635;
	wire [14-1:0] node636;
	wire [14-1:0] node638;
	wire [14-1:0] node640;
	wire [14-1:0] node643;
	wire [14-1:0] node644;
	wire [14-1:0] node647;
	wire [14-1:0] node650;
	wire [14-1:0] node651;
	wire [14-1:0] node652;
	wire [14-1:0] node653;
	wire [14-1:0] node654;
	wire [14-1:0] node657;
	wire [14-1:0] node658;
	wire [14-1:0] node660;
	wire [14-1:0] node664;
	wire [14-1:0] node665;
	wire [14-1:0] node667;
	wire [14-1:0] node668;
	wire [14-1:0] node673;
	wire [14-1:0] node674;
	wire [14-1:0] node675;
	wire [14-1:0] node678;
	wire [14-1:0] node681;
	wire [14-1:0] node682;
	wire [14-1:0] node684;
	wire [14-1:0] node686;
	wire [14-1:0] node689;
	wire [14-1:0] node690;
	wire [14-1:0] node694;
	wire [14-1:0] node695;
	wire [14-1:0] node696;
	wire [14-1:0] node697;
	wire [14-1:0] node700;
	wire [14-1:0] node702;
	wire [14-1:0] node705;
	wire [14-1:0] node706;
	wire [14-1:0] node708;
	wire [14-1:0] node712;
	wire [14-1:0] node713;
	wire [14-1:0] node714;
	wire [14-1:0] node716;
	wire [14-1:0] node718;
	wire [14-1:0] node721;
	wire [14-1:0] node723;
	wire [14-1:0] node726;
	wire [14-1:0] node727;
	wire [14-1:0] node728;
	wire [14-1:0] node730;
	wire [14-1:0] node734;
	wire [14-1:0] node735;
	wire [14-1:0] node739;
	wire [14-1:0] node740;
	wire [14-1:0] node741;
	wire [14-1:0] node742;
	wire [14-1:0] node743;
	wire [14-1:0] node744;
	wire [14-1:0] node745;
	wire [14-1:0] node747;
	wire [14-1:0] node748;
	wire [14-1:0] node752;
	wire [14-1:0] node753;
	wire [14-1:0] node754;
	wire [14-1:0] node755;
	wire [14-1:0] node759;
	wire [14-1:0] node762;
	wire [14-1:0] node765;
	wire [14-1:0] node766;
	wire [14-1:0] node767;
	wire [14-1:0] node768;
	wire [14-1:0] node769;
	wire [14-1:0] node772;
	wire [14-1:0] node777;
	wire [14-1:0] node778;
	wire [14-1:0] node779;
	wire [14-1:0] node783;
	wire [14-1:0] node786;
	wire [14-1:0] node787;
	wire [14-1:0] node788;
	wire [14-1:0] node789;
	wire [14-1:0] node792;
	wire [14-1:0] node794;
	wire [14-1:0] node797;
	wire [14-1:0] node798;
	wire [14-1:0] node800;
	wire [14-1:0] node803;
	wire [14-1:0] node804;
	wire [14-1:0] node808;
	wire [14-1:0] node809;
	wire [14-1:0] node811;
	wire [14-1:0] node814;
	wire [14-1:0] node815;
	wire [14-1:0] node818;
	wire [14-1:0] node820;
	wire [14-1:0] node823;
	wire [14-1:0] node824;
	wire [14-1:0] node825;
	wire [14-1:0] node826;
	wire [14-1:0] node827;
	wire [14-1:0] node829;
	wire [14-1:0] node831;
	wire [14-1:0] node834;
	wire [14-1:0] node837;
	wire [14-1:0] node839;
	wire [14-1:0] node841;
	wire [14-1:0] node843;
	wire [14-1:0] node846;
	wire [14-1:0] node847;
	wire [14-1:0] node848;
	wire [14-1:0] node849;
	wire [14-1:0] node853;
	wire [14-1:0] node855;
	wire [14-1:0] node858;
	wire [14-1:0] node859;
	wire [14-1:0] node863;
	wire [14-1:0] node864;
	wire [14-1:0] node865;
	wire [14-1:0] node866;
	wire [14-1:0] node868;
	wire [14-1:0] node871;
	wire [14-1:0] node872;
	wire [14-1:0] node873;
	wire [14-1:0] node876;
	wire [14-1:0] node879;
	wire [14-1:0] node880;
	wire [14-1:0] node884;
	wire [14-1:0] node886;
	wire [14-1:0] node887;
	wire [14-1:0] node889;
	wire [14-1:0] node892;
	wire [14-1:0] node895;
	wire [14-1:0] node896;
	wire [14-1:0] node897;
	wire [14-1:0] node900;
	wire [14-1:0] node902;
	wire [14-1:0] node903;
	wire [14-1:0] node907;
	wire [14-1:0] node908;
	wire [14-1:0] node909;
	wire [14-1:0] node911;
	wire [14-1:0] node915;
	wire [14-1:0] node917;
	wire [14-1:0] node918;
	wire [14-1:0] node922;
	wire [14-1:0] node923;
	wire [14-1:0] node924;
	wire [14-1:0] node925;
	wire [14-1:0] node926;
	wire [14-1:0] node927;
	wire [14-1:0] node928;
	wire [14-1:0] node932;
	wire [14-1:0] node935;
	wire [14-1:0] node936;
	wire [14-1:0] node937;
	wire [14-1:0] node939;
	wire [14-1:0] node943;
	wire [14-1:0] node944;
	wire [14-1:0] node945;
	wire [14-1:0] node950;
	wire [14-1:0] node951;
	wire [14-1:0] node952;
	wire [14-1:0] node953;
	wire [14-1:0] node954;
	wire [14-1:0] node955;
	wire [14-1:0] node960;
	wire [14-1:0] node962;
	wire [14-1:0] node965;
	wire [14-1:0] node966;
	wire [14-1:0] node970;
	wire [14-1:0] node971;
	wire [14-1:0] node974;
	wire [14-1:0] node976;
	wire [14-1:0] node978;
	wire [14-1:0] node981;
	wire [14-1:0] node982;
	wire [14-1:0] node983;
	wire [14-1:0] node984;
	wire [14-1:0] node985;
	wire [14-1:0] node989;
	wire [14-1:0] node992;
	wire [14-1:0] node993;
	wire [14-1:0] node994;
	wire [14-1:0] node997;
	wire [14-1:0] node1000;
	wire [14-1:0] node1001;
	wire [14-1:0] node1003;
	wire [14-1:0] node1005;
	wire [14-1:0] node1006;
	wire [14-1:0] node1011;
	wire [14-1:0] node1012;
	wire [14-1:0] node1013;
	wire [14-1:0] node1016;
	wire [14-1:0] node1017;
	wire [14-1:0] node1021;
	wire [14-1:0] node1023;
	wire [14-1:0] node1025;
	wire [14-1:0] node1028;
	wire [14-1:0] node1029;
	wire [14-1:0] node1030;
	wire [14-1:0] node1031;
	wire [14-1:0] node1032;
	wire [14-1:0] node1033;
	wire [14-1:0] node1036;
	wire [14-1:0] node1037;
	wire [14-1:0] node1040;
	wire [14-1:0] node1044;
	wire [14-1:0] node1046;
	wire [14-1:0] node1049;
	wire [14-1:0] node1050;
	wire [14-1:0] node1051;
	wire [14-1:0] node1052;
	wire [14-1:0] node1055;
	wire [14-1:0] node1057;
	wire [14-1:0] node1061;
	wire [14-1:0] node1062;
	wire [14-1:0] node1066;
	wire [14-1:0] node1067;
	wire [14-1:0] node1068;
	wire [14-1:0] node1069;
	wire [14-1:0] node1073;
	wire [14-1:0] node1075;
	wire [14-1:0] node1077;
	wire [14-1:0] node1080;
	wire [14-1:0] node1081;
	wire [14-1:0] node1082;
	wire [14-1:0] node1083;
	wire [14-1:0] node1087;
	wire [14-1:0] node1088;
	wire [14-1:0] node1089;
	wire [14-1:0] node1094;
	wire [14-1:0] node1095;
	wire [14-1:0] node1098;
	wire [14-1:0] node1100;
	wire [14-1:0] node1102;
	wire [14-1:0] node1105;
	wire [14-1:0] node1106;
	wire [14-1:0] node1107;
	wire [14-1:0] node1108;
	wire [14-1:0] node1109;
	wire [14-1:0] node1110;
	wire [14-1:0] node1111;
	wire [14-1:0] node1114;
	wire [14-1:0] node1116;
	wire [14-1:0] node1119;
	wire [14-1:0] node1120;
	wire [14-1:0] node1122;
	wire [14-1:0] node1124;
	wire [14-1:0] node1127;
	wire [14-1:0] node1130;
	wire [14-1:0] node1131;
	wire [14-1:0] node1132;
	wire [14-1:0] node1135;
	wire [14-1:0] node1138;
	wire [14-1:0] node1139;
	wire [14-1:0] node1142;
	wire [14-1:0] node1145;
	wire [14-1:0] node1146;
	wire [14-1:0] node1147;
	wire [14-1:0] node1148;
	wire [14-1:0] node1150;
	wire [14-1:0] node1153;
	wire [14-1:0] node1156;
	wire [14-1:0] node1158;
	wire [14-1:0] node1160;
	wire [14-1:0] node1163;
	wire [14-1:0] node1164;
	wire [14-1:0] node1165;
	wire [14-1:0] node1168;
	wire [14-1:0] node1171;
	wire [14-1:0] node1172;
	wire [14-1:0] node1176;
	wire [14-1:0] node1177;
	wire [14-1:0] node1178;
	wire [14-1:0] node1179;
	wire [14-1:0] node1180;
	wire [14-1:0] node1181;
	wire [14-1:0] node1185;
	wire [14-1:0] node1187;
	wire [14-1:0] node1190;
	wire [14-1:0] node1191;
	wire [14-1:0] node1195;
	wire [14-1:0] node1196;
	wire [14-1:0] node1197;
	wire [14-1:0] node1200;
	wire [14-1:0] node1203;
	wire [14-1:0] node1204;
	wire [14-1:0] node1205;
	wire [14-1:0] node1207;
	wire [14-1:0] node1211;
	wire [14-1:0] node1214;
	wire [14-1:0] node1215;
	wire [14-1:0] node1216;
	wire [14-1:0] node1217;
	wire [14-1:0] node1220;
	wire [14-1:0] node1222;
	wire [14-1:0] node1223;
	wire [14-1:0] node1227;
	wire [14-1:0] node1228;
	wire [14-1:0] node1231;
	wire [14-1:0] node1234;
	wire [14-1:0] node1235;
	wire [14-1:0] node1237;
	wire [14-1:0] node1240;
	wire [14-1:0] node1242;
	wire [14-1:0] node1245;
	wire [14-1:0] node1246;
	wire [14-1:0] node1247;
	wire [14-1:0] node1248;
	wire [14-1:0] node1249;
	wire [14-1:0] node1250;
	wire [14-1:0] node1254;
	wire [14-1:0] node1255;
	wire [14-1:0] node1256;
	wire [14-1:0] node1260;
	wire [14-1:0] node1263;
	wire [14-1:0] node1264;
	wire [14-1:0] node1265;
	wire [14-1:0] node1266;
	wire [14-1:0] node1269;
	wire [14-1:0] node1272;
	wire [14-1:0] node1274;
	wire [14-1:0] node1276;
	wire [14-1:0] node1278;
	wire [14-1:0] node1281;
	wire [14-1:0] node1282;
	wire [14-1:0] node1283;
	wire [14-1:0] node1287;
	wire [14-1:0] node1289;
	wire [14-1:0] node1292;
	wire [14-1:0] node1293;
	wire [14-1:0] node1294;
	wire [14-1:0] node1297;
	wire [14-1:0] node1299;
	wire [14-1:0] node1302;
	wire [14-1:0] node1303;
	wire [14-1:0] node1304;
	wire [14-1:0] node1307;
	wire [14-1:0] node1308;
	wire [14-1:0] node1309;
	wire [14-1:0] node1314;
	wire [14-1:0] node1315;
	wire [14-1:0] node1316;
	wire [14-1:0] node1319;
	wire [14-1:0] node1322;
	wire [14-1:0] node1325;
	wire [14-1:0] node1326;
	wire [14-1:0] node1327;
	wire [14-1:0] node1328;
	wire [14-1:0] node1329;
	wire [14-1:0] node1330;
	wire [14-1:0] node1332;
	wire [14-1:0] node1333;
	wire [14-1:0] node1339;
	wire [14-1:0] node1340;
	wire [14-1:0] node1342;
	wire [14-1:0] node1343;
	wire [14-1:0] node1347;
	wire [14-1:0] node1348;
	wire [14-1:0] node1350;
	wire [14-1:0] node1354;
	wire [14-1:0] node1355;
	wire [14-1:0] node1356;
	wire [14-1:0] node1357;
	wire [14-1:0] node1361;
	wire [14-1:0] node1364;
	wire [14-1:0] node1365;
	wire [14-1:0] node1368;
	wire [14-1:0] node1369;
	wire [14-1:0] node1373;
	wire [14-1:0] node1374;
	wire [14-1:0] node1375;
	wire [14-1:0] node1377;
	wire [14-1:0] node1379;
	wire [14-1:0] node1380;
	wire [14-1:0] node1382;
	wire [14-1:0] node1386;
	wire [14-1:0] node1387;
	wire [14-1:0] node1389;
	wire [14-1:0] node1392;
	wire [14-1:0] node1393;
	wire [14-1:0] node1396;
	wire [14-1:0] node1398;
	wire [14-1:0] node1401;
	wire [14-1:0] node1402;
	wire [14-1:0] node1403;
	wire [14-1:0] node1404;
	wire [14-1:0] node1407;
	wire [14-1:0] node1411;
	wire [14-1:0] node1412;
	wire [14-1:0] node1415;
	wire [14-1:0] node1416;
	wire [14-1:0] node1418;
	wire [14-1:0] node1421;
	wire [14-1:0] node1422;
	wire [14-1:0] node1426;
	wire [14-1:0] node1427;
	wire [14-1:0] node1428;
	wire [14-1:0] node1429;
	wire [14-1:0] node1430;
	wire [14-1:0] node1431;
	wire [14-1:0] node1432;
	wire [14-1:0] node1433;
	wire [14-1:0] node1434;
	wire [14-1:0] node1435;
	wire [14-1:0] node1438;
	wire [14-1:0] node1439;
	wire [14-1:0] node1443;
	wire [14-1:0] node1444;
	wire [14-1:0] node1447;
	wire [14-1:0] node1450;
	wire [14-1:0] node1451;
	wire [14-1:0] node1452;
	wire [14-1:0] node1454;
	wire [14-1:0] node1458;
	wire [14-1:0] node1461;
	wire [14-1:0] node1462;
	wire [14-1:0] node1464;
	wire [14-1:0] node1465;
	wire [14-1:0] node1469;
	wire [14-1:0] node1470;
	wire [14-1:0] node1472;
	wire [14-1:0] node1473;
	wire [14-1:0] node1478;
	wire [14-1:0] node1479;
	wire [14-1:0] node1480;
	wire [14-1:0] node1481;
	wire [14-1:0] node1482;
	wire [14-1:0] node1486;
	wire [14-1:0] node1489;
	wire [14-1:0] node1490;
	wire [14-1:0] node1493;
	wire [14-1:0] node1495;
	wire [14-1:0] node1498;
	wire [14-1:0] node1499;
	wire [14-1:0] node1500;
	wire [14-1:0] node1502;
	wire [14-1:0] node1504;
	wire [14-1:0] node1507;
	wire [14-1:0] node1509;
	wire [14-1:0] node1510;
	wire [14-1:0] node1514;
	wire [14-1:0] node1515;
	wire [14-1:0] node1517;
	wire [14-1:0] node1519;
	wire [14-1:0] node1522;
	wire [14-1:0] node1523;
	wire [14-1:0] node1527;
	wire [14-1:0] node1528;
	wire [14-1:0] node1529;
	wire [14-1:0] node1530;
	wire [14-1:0] node1532;
	wire [14-1:0] node1533;
	wire [14-1:0] node1536;
	wire [14-1:0] node1537;
	wire [14-1:0] node1541;
	wire [14-1:0] node1542;
	wire [14-1:0] node1543;
	wire [14-1:0] node1544;
	wire [14-1:0] node1549;
	wire [14-1:0] node1550;
	wire [14-1:0] node1554;
	wire [14-1:0] node1555;
	wire [14-1:0] node1556;
	wire [14-1:0] node1558;
	wire [14-1:0] node1561;
	wire [14-1:0] node1562;
	wire [14-1:0] node1565;
	wire [14-1:0] node1568;
	wire [14-1:0] node1569;
	wire [14-1:0] node1570;
	wire [14-1:0] node1574;
	wire [14-1:0] node1577;
	wire [14-1:0] node1578;
	wire [14-1:0] node1579;
	wire [14-1:0] node1580;
	wire [14-1:0] node1584;
	wire [14-1:0] node1585;
	wire [14-1:0] node1589;
	wire [14-1:0] node1590;
	wire [14-1:0] node1591;
	wire [14-1:0] node1592;
	wire [14-1:0] node1595;
	wire [14-1:0] node1598;
	wire [14-1:0] node1599;
	wire [14-1:0] node1603;
	wire [14-1:0] node1604;
	wire [14-1:0] node1607;
	wire [14-1:0] node1610;
	wire [14-1:0] node1611;
	wire [14-1:0] node1612;
	wire [14-1:0] node1613;
	wire [14-1:0] node1614;
	wire [14-1:0] node1615;
	wire [14-1:0] node1616;
	wire [14-1:0] node1619;
	wire [14-1:0] node1622;
	wire [14-1:0] node1624;
	wire [14-1:0] node1625;
	wire [14-1:0] node1629;
	wire [14-1:0] node1630;
	wire [14-1:0] node1633;
	wire [14-1:0] node1635;
	wire [14-1:0] node1636;
	wire [14-1:0] node1640;
	wire [14-1:0] node1641;
	wire [14-1:0] node1642;
	wire [14-1:0] node1644;
	wire [14-1:0] node1645;
	wire [14-1:0] node1649;
	wire [14-1:0] node1650;
	wire [14-1:0] node1652;
	wire [14-1:0] node1656;
	wire [14-1:0] node1658;
	wire [14-1:0] node1661;
	wire [14-1:0] node1662;
	wire [14-1:0] node1663;
	wire [14-1:0] node1665;
	wire [14-1:0] node1667;
	wire [14-1:0] node1670;
	wire [14-1:0] node1671;
	wire [14-1:0] node1672;
	wire [14-1:0] node1676;
	wire [14-1:0] node1679;
	wire [14-1:0] node1680;
	wire [14-1:0] node1681;
	wire [14-1:0] node1682;
	wire [14-1:0] node1686;
	wire [14-1:0] node1688;
	wire [14-1:0] node1691;
	wire [14-1:0] node1694;
	wire [14-1:0] node1695;
	wire [14-1:0] node1696;
	wire [14-1:0] node1697;
	wire [14-1:0] node1698;
	wire [14-1:0] node1699;
	wire [14-1:0] node1700;
	wire [14-1:0] node1706;
	wire [14-1:0] node1707;
	wire [14-1:0] node1709;
	wire [14-1:0] node1713;
	wire [14-1:0] node1714;
	wire [14-1:0] node1717;
	wire [14-1:0] node1718;
	wire [14-1:0] node1720;
	wire [14-1:0] node1722;
	wire [14-1:0] node1726;
	wire [14-1:0] node1727;
	wire [14-1:0] node1728;
	wire [14-1:0] node1729;
	wire [14-1:0] node1730;
	wire [14-1:0] node1735;
	wire [14-1:0] node1736;
	wire [14-1:0] node1737;
	wire [14-1:0] node1739;
	wire [14-1:0] node1743;
	wire [14-1:0] node1746;
	wire [14-1:0] node1747;
	wire [14-1:0] node1748;
	wire [14-1:0] node1751;
	wire [14-1:0] node1752;
	wire [14-1:0] node1756;
	wire [14-1:0] node1757;
	wire [14-1:0] node1759;
	wire [14-1:0] node1762;
	wire [14-1:0] node1765;
	wire [14-1:0] node1766;
	wire [14-1:0] node1767;
	wire [14-1:0] node1768;
	wire [14-1:0] node1769;
	wire [14-1:0] node1770;
	wire [14-1:0] node1771;
	wire [14-1:0] node1772;
	wire [14-1:0] node1773;
	wire [14-1:0] node1775;
	wire [14-1:0] node1781;
	wire [14-1:0] node1782;
	wire [14-1:0] node1784;
	wire [14-1:0] node1787;
	wire [14-1:0] node1790;
	wire [14-1:0] node1791;
	wire [14-1:0] node1792;
	wire [14-1:0] node1793;
	wire [14-1:0] node1794;
	wire [14-1:0] node1799;
	wire [14-1:0] node1800;
	wire [14-1:0] node1802;
	wire [14-1:0] node1805;
	wire [14-1:0] node1808;
	wire [14-1:0] node1809;
	wire [14-1:0] node1810;
	wire [14-1:0] node1814;
	wire [14-1:0] node1817;
	wire [14-1:0] node1818;
	wire [14-1:0] node1819;
	wire [14-1:0] node1820;
	wire [14-1:0] node1823;
	wire [14-1:0] node1826;
	wire [14-1:0] node1827;
	wire [14-1:0] node1831;
	wire [14-1:0] node1832;
	wire [14-1:0] node1833;
	wire [14-1:0] node1834;
	wire [14-1:0] node1836;
	wire [14-1:0] node1840;
	wire [14-1:0] node1842;
	wire [14-1:0] node1843;
	wire [14-1:0] node1845;
	wire [14-1:0] node1849;
	wire [14-1:0] node1850;
	wire [14-1:0] node1852;
	wire [14-1:0] node1855;
	wire [14-1:0] node1858;
	wire [14-1:0] node1859;
	wire [14-1:0] node1860;
	wire [14-1:0] node1861;
	wire [14-1:0] node1862;
	wire [14-1:0] node1863;
	wire [14-1:0] node1866;
	wire [14-1:0] node1869;
	wire [14-1:0] node1870;
	wire [14-1:0] node1874;
	wire [14-1:0] node1875;
	wire [14-1:0] node1879;
	wire [14-1:0] node1880;
	wire [14-1:0] node1881;
	wire [14-1:0] node1882;
	wire [14-1:0] node1885;
	wire [14-1:0] node1886;
	wire [14-1:0] node1890;
	wire [14-1:0] node1893;
	wire [14-1:0] node1895;
	wire [14-1:0] node1896;
	wire [14-1:0] node1900;
	wire [14-1:0] node1901;
	wire [14-1:0] node1902;
	wire [14-1:0] node1903;
	wire [14-1:0] node1905;
	wire [14-1:0] node1909;
	wire [14-1:0] node1910;
	wire [14-1:0] node1913;
	wire [14-1:0] node1915;
	wire [14-1:0] node1918;
	wire [14-1:0] node1919;
	wire [14-1:0] node1921;
	wire [14-1:0] node1923;
	wire [14-1:0] node1924;
	wire [14-1:0] node1928;
	wire [14-1:0] node1929;
	wire [14-1:0] node1931;
	wire [14-1:0] node1934;
	wire [14-1:0] node1936;
	wire [14-1:0] node1938;
	wire [14-1:0] node1941;
	wire [14-1:0] node1942;
	wire [14-1:0] node1943;
	wire [14-1:0] node1944;
	wire [14-1:0] node1945;
	wire [14-1:0] node1946;
	wire [14-1:0] node1947;
	wire [14-1:0] node1952;
	wire [14-1:0] node1953;
	wire [14-1:0] node1954;
	wire [14-1:0] node1957;
	wire [14-1:0] node1960;
	wire [14-1:0] node1962;
	wire [14-1:0] node1965;
	wire [14-1:0] node1966;
	wire [14-1:0] node1967;
	wire [14-1:0] node1969;
	wire [14-1:0] node1970;
	wire [14-1:0] node1974;
	wire [14-1:0] node1977;
	wire [14-1:0] node1978;
	wire [14-1:0] node1979;
	wire [14-1:0] node1983;
	wire [14-1:0] node1985;
	wire [14-1:0] node1988;
	wire [14-1:0] node1989;
	wire [14-1:0] node1990;
	wire [14-1:0] node1991;
	wire [14-1:0] node1992;
	wire [14-1:0] node1996;
	wire [14-1:0] node1999;
	wire [14-1:0] node2000;
	wire [14-1:0] node2002;
	wire [14-1:0] node2005;
	wire [14-1:0] node2006;
	wire [14-1:0] node2010;
	wire [14-1:0] node2011;
	wire [14-1:0] node2012;
	wire [14-1:0] node2016;
	wire [14-1:0] node2017;
	wire [14-1:0] node2020;
	wire [14-1:0] node2021;
	wire [14-1:0] node2025;
	wire [14-1:0] node2026;
	wire [14-1:0] node2027;
	wire [14-1:0] node2028;
	wire [14-1:0] node2029;
	wire [14-1:0] node2030;
	wire [14-1:0] node2032;
	wire [14-1:0] node2033;
	wire [14-1:0] node2038;
	wire [14-1:0] node2040;
	wire [14-1:0] node2041;
	wire [14-1:0] node2045;
	wire [14-1:0] node2046;
	wire [14-1:0] node2047;
	wire [14-1:0] node2049;
	wire [14-1:0] node2053;
	wire [14-1:0] node2056;
	wire [14-1:0] node2057;
	wire [14-1:0] node2058;
	wire [14-1:0] node2060;
	wire [14-1:0] node2061;
	wire [14-1:0] node2065;
	wire [14-1:0] node2066;
	wire [14-1:0] node2068;
	wire [14-1:0] node2072;
	wire [14-1:0] node2073;
	wire [14-1:0] node2076;
	wire [14-1:0] node2077;
	wire [14-1:0] node2080;
	wire [14-1:0] node2083;
	wire [14-1:0] node2084;
	wire [14-1:0] node2085;
	wire [14-1:0] node2086;
	wire [14-1:0] node2087;
	wire [14-1:0] node2088;
	wire [14-1:0] node2093;
	wire [14-1:0] node2094;
	wire [14-1:0] node2096;
	wire [14-1:0] node2100;
	wire [14-1:0] node2101;
	wire [14-1:0] node2102;
	wire [14-1:0] node2105;
	wire [14-1:0] node2106;
	wire [14-1:0] node2110;
	wire [14-1:0] node2113;
	wire [14-1:0] node2114;
	wire [14-1:0] node2115;
	wire [14-1:0] node2117;
	wire [14-1:0] node2120;
	wire [14-1:0] node2121;
	wire [14-1:0] node2123;
	wire [14-1:0] node2127;
	wire [14-1:0] node2128;
	wire [14-1:0] node2131;
	wire [14-1:0] node2133;
	wire [14-1:0] node2134;
	wire [14-1:0] node2138;
	wire [14-1:0] node2139;
	wire [14-1:0] node2140;
	wire [14-1:0] node2141;
	wire [14-1:0] node2142;
	wire [14-1:0] node2143;
	wire [14-1:0] node2144;
	wire [14-1:0] node2145;
	wire [14-1:0] node2148;
	wire [14-1:0] node2151;
	wire [14-1:0] node2152;
	wire [14-1:0] node2154;
	wire [14-1:0] node2155;
	wire [14-1:0] node2159;
	wire [14-1:0] node2162;
	wire [14-1:0] node2163;
	wire [14-1:0] node2164;
	wire [14-1:0] node2168;
	wire [14-1:0] node2169;
	wire [14-1:0] node2170;
	wire [14-1:0] node2171;
	wire [14-1:0] node2175;
	wire [14-1:0] node2177;
	wire [14-1:0] node2180;
	wire [14-1:0] node2183;
	wire [14-1:0] node2184;
	wire [14-1:0] node2185;
	wire [14-1:0] node2186;
	wire [14-1:0] node2189;
	wire [14-1:0] node2190;
	wire [14-1:0] node2192;
	wire [14-1:0] node2196;
	wire [14-1:0] node2197;
	wire [14-1:0] node2199;
	wire [14-1:0] node2200;
	wire [14-1:0] node2205;
	wire [14-1:0] node2206;
	wire [14-1:0] node2209;
	wire [14-1:0] node2210;
	wire [14-1:0] node2211;
	wire [14-1:0] node2214;
	wire [14-1:0] node2217;
	wire [14-1:0] node2219;
	wire [14-1:0] node2222;
	wire [14-1:0] node2223;
	wire [14-1:0] node2224;
	wire [14-1:0] node2225;
	wire [14-1:0] node2226;
	wire [14-1:0] node2227;
	wire [14-1:0] node2231;
	wire [14-1:0] node2232;
	wire [14-1:0] node2236;
	wire [14-1:0] node2237;
	wire [14-1:0] node2238;
	wire [14-1:0] node2240;
	wire [14-1:0] node2245;
	wire [14-1:0] node2246;
	wire [14-1:0] node2247;
	wire [14-1:0] node2249;
	wire [14-1:0] node2250;
	wire [14-1:0] node2251;
	wire [14-1:0] node2256;
	wire [14-1:0] node2259;
	wire [14-1:0] node2260;
	wire [14-1:0] node2261;
	wire [14-1:0] node2264;
	wire [14-1:0] node2265;
	wire [14-1:0] node2267;
	wire [14-1:0] node2271;
	wire [14-1:0] node2272;
	wire [14-1:0] node2273;
	wire [14-1:0] node2277;
	wire [14-1:0] node2280;
	wire [14-1:0] node2281;
	wire [14-1:0] node2282;
	wire [14-1:0] node2284;
	wire [14-1:0] node2287;
	wire [14-1:0] node2288;
	wire [14-1:0] node2291;
	wire [14-1:0] node2293;
	wire [14-1:0] node2296;
	wire [14-1:0] node2297;
	wire [14-1:0] node2298;
	wire [14-1:0] node2301;
	wire [14-1:0] node2304;
	wire [14-1:0] node2305;
	wire [14-1:0] node2308;
	wire [14-1:0] node2311;
	wire [14-1:0] node2312;
	wire [14-1:0] node2313;
	wire [14-1:0] node2314;
	wire [14-1:0] node2315;
	wire [14-1:0] node2316;
	wire [14-1:0] node2317;
	wire [14-1:0] node2321;
	wire [14-1:0] node2322;
	wire [14-1:0] node2326;
	wire [14-1:0] node2327;
	wire [14-1:0] node2329;
	wire [14-1:0] node2330;
	wire [14-1:0] node2334;
	wire [14-1:0] node2335;
	wire [14-1:0] node2339;
	wire [14-1:0] node2340;
	wire [14-1:0] node2341;
	wire [14-1:0] node2343;
	wire [14-1:0] node2344;
	wire [14-1:0] node2348;
	wire [14-1:0] node2350;
	wire [14-1:0] node2353;
	wire [14-1:0] node2354;
	wire [14-1:0] node2357;
	wire [14-1:0] node2360;
	wire [14-1:0] node2361;
	wire [14-1:0] node2362;
	wire [14-1:0] node2363;
	wire [14-1:0] node2364;
	wire [14-1:0] node2366;
	wire [14-1:0] node2370;
	wire [14-1:0] node2373;
	wire [14-1:0] node2374;
	wire [14-1:0] node2376;
	wire [14-1:0] node2379;
	wire [14-1:0] node2382;
	wire [14-1:0] node2383;
	wire [14-1:0] node2384;
	wire [14-1:0] node2385;
	wire [14-1:0] node2389;
	wire [14-1:0] node2390;
	wire [14-1:0] node2392;
	wire [14-1:0] node2395;
	wire [14-1:0] node2398;
	wire [14-1:0] node2399;
	wire [14-1:0] node2401;
	wire [14-1:0] node2403;
	wire [14-1:0] node2406;
	wire [14-1:0] node2409;
	wire [14-1:0] node2410;
	wire [14-1:0] node2411;
	wire [14-1:0] node2412;
	wire [14-1:0] node2413;
	wire [14-1:0] node2416;
	wire [14-1:0] node2418;
	wire [14-1:0] node2421;
	wire [14-1:0] node2423;
	wire [14-1:0] node2425;
	wire [14-1:0] node2426;
	wire [14-1:0] node2428;
	wire [14-1:0] node2432;
	wire [14-1:0] node2433;
	wire [14-1:0] node2435;
	wire [14-1:0] node2436;
	wire [14-1:0] node2440;
	wire [14-1:0] node2441;
	wire [14-1:0] node2444;
	wire [14-1:0] node2445;
	wire [14-1:0] node2449;
	wire [14-1:0] node2450;
	wire [14-1:0] node2451;
	wire [14-1:0] node2453;
	wire [14-1:0] node2455;
	wire [14-1:0] node2458;
	wire [14-1:0] node2460;
	wire [14-1:0] node2462;
	wire [14-1:0] node2463;
	wire [14-1:0] node2467;
	wire [14-1:0] node2468;
	wire [14-1:0] node2469;
	wire [14-1:0] node2472;
	wire [14-1:0] node2474;
	wire [14-1:0] node2477;
	wire [14-1:0] node2478;
	wire [14-1:0] node2479;
	wire [14-1:0] node2483;
	wire [14-1:0] node2484;
	wire [14-1:0] node2485;
	wire [14-1:0] node2490;
	wire [14-1:0] node2491;
	wire [14-1:0] node2492;
	wire [14-1:0] node2493;
	wire [14-1:0] node2494;
	wire [14-1:0] node2495;
	wire [14-1:0] node2496;
	wire [14-1:0] node2497;
	wire [14-1:0] node2501;
	wire [14-1:0] node2502;
	wire [14-1:0] node2504;
	wire [14-1:0] node2508;
	wire [14-1:0] node2510;
	wire [14-1:0] node2511;
	wire [14-1:0] node2515;
	wire [14-1:0] node2516;
	wire [14-1:0] node2517;
	wire [14-1:0] node2518;
	wire [14-1:0] node2521;
	wire [14-1:0] node2523;
	wire [14-1:0] node2526;
	wire [14-1:0] node2528;
	wire [14-1:0] node2531;
	wire [14-1:0] node2532;
	wire [14-1:0] node2535;
	wire [14-1:0] node2536;
	wire [14-1:0] node2540;
	wire [14-1:0] node2541;
	wire [14-1:0] node2542;
	wire [14-1:0] node2543;
	wire [14-1:0] node2545;
	wire [14-1:0] node2546;
	wire [14-1:0] node2550;
	wire [14-1:0] node2553;
	wire [14-1:0] node2554;
	wire [14-1:0] node2557;
	wire [14-1:0] node2560;
	wire [14-1:0] node2561;
	wire [14-1:0] node2563;
	wire [14-1:0] node2564;
	wire [14-1:0] node2568;
	wire [14-1:0] node2569;
	wire [14-1:0] node2570;
	wire [14-1:0] node2571;
	wire [14-1:0] node2574;
	wire [14-1:0] node2577;
	wire [14-1:0] node2580;
	wire [14-1:0] node2581;
	wire [14-1:0] node2584;
	wire [14-1:0] node2587;
	wire [14-1:0] node2588;
	wire [14-1:0] node2589;
	wire [14-1:0] node2590;
	wire [14-1:0] node2592;
	wire [14-1:0] node2594;
	wire [14-1:0] node2595;
	wire [14-1:0] node2599;
	wire [14-1:0] node2600;
	wire [14-1:0] node2602;
	wire [14-1:0] node2604;
	wire [14-1:0] node2607;
	wire [14-1:0] node2608;
	wire [14-1:0] node2612;
	wire [14-1:0] node2613;
	wire [14-1:0] node2614;
	wire [14-1:0] node2617;
	wire [14-1:0] node2619;
	wire [14-1:0] node2620;
	wire [14-1:0] node2621;
	wire [14-1:0] node2623;
	wire [14-1:0] node2626;
	wire [14-1:0] node2627;
	wire [14-1:0] node2632;
	wire [14-1:0] node2633;
	wire [14-1:0] node2636;
	wire [14-1:0] node2638;
	wire [14-1:0] node2639;
	wire [14-1:0] node2643;
	wire [14-1:0] node2644;
	wire [14-1:0] node2645;
	wire [14-1:0] node2646;
	wire [14-1:0] node2649;
	wire [14-1:0] node2651;
	wire [14-1:0] node2652;
	wire [14-1:0] node2656;
	wire [14-1:0] node2657;
	wire [14-1:0] node2658;
	wire [14-1:0] node2660;
	wire [14-1:0] node2663;
	wire [14-1:0] node2667;
	wire [14-1:0] node2668;
	wire [14-1:0] node2669;
	wire [14-1:0] node2670;
	wire [14-1:0] node2674;
	wire [14-1:0] node2675;
	wire [14-1:0] node2679;
	wire [14-1:0] node2680;
	wire [14-1:0] node2682;
	wire [14-1:0] node2684;
	wire [14-1:0] node2687;
	wire [14-1:0] node2690;
	wire [14-1:0] node2691;
	wire [14-1:0] node2692;
	wire [14-1:0] node2693;
	wire [14-1:0] node2694;
	wire [14-1:0] node2695;
	wire [14-1:0] node2697;
	wire [14-1:0] node2698;
	wire [14-1:0] node2702;
	wire [14-1:0] node2703;
	wire [14-1:0] node2707;
	wire [14-1:0] node2708;
	wire [14-1:0] node2709;
	wire [14-1:0] node2710;
	wire [14-1:0] node2715;
	wire [14-1:0] node2716;
	wire [14-1:0] node2720;
	wire [14-1:0] node2721;
	wire [14-1:0] node2723;
	wire [14-1:0] node2727;
	wire [14-1:0] node2728;
	wire [14-1:0] node2729;
	wire [14-1:0] node2730;
	wire [14-1:0] node2733;
	wire [14-1:0] node2734;
	wire [14-1:0] node2735;
	wire [14-1:0] node2739;
	wire [14-1:0] node2742;
	wire [14-1:0] node2743;
	wire [14-1:0] node2744;
	wire [14-1:0] node2746;
	wire [14-1:0] node2750;
	wire [14-1:0] node2752;
	wire [14-1:0] node2755;
	wire [14-1:0] node2756;
	wire [14-1:0] node2757;
	wire [14-1:0] node2760;
	wire [14-1:0] node2762;
	wire [14-1:0] node2764;
	wire [14-1:0] node2767;
	wire [14-1:0] node2769;
	wire [14-1:0] node2770;
	wire [14-1:0] node2773;
	wire [14-1:0] node2775;
	wire [14-1:0] node2776;
	wire [14-1:0] node2778;
	wire [14-1:0] node2782;
	wire [14-1:0] node2783;
	wire [14-1:0] node2784;
	wire [14-1:0] node2785;
	wire [14-1:0] node2786;
	wire [14-1:0] node2790;
	wire [14-1:0] node2791;
	wire [14-1:0] node2794;
	wire [14-1:0] node2795;
	wire [14-1:0] node2797;
	wire [14-1:0] node2800;
	wire [14-1:0] node2801;
	wire [14-1:0] node2805;
	wire [14-1:0] node2806;
	wire [14-1:0] node2807;
	wire [14-1:0] node2809;
	wire [14-1:0] node2813;
	wire [14-1:0] node2814;
	wire [14-1:0] node2817;
	wire [14-1:0] node2820;
	wire [14-1:0] node2821;
	wire [14-1:0] node2823;
	wire [14-1:0] node2824;
	wire [14-1:0] node2825;
	wire [14-1:0] node2826;
	wire [14-1:0] node2831;
	wire [14-1:0] node2833;
	wire [14-1:0] node2834;
	wire [14-1:0] node2836;
	wire [14-1:0] node2840;
	wire [14-1:0] node2841;
	wire [14-1:0] node2842;
	wire [14-1:0] node2844;
	wire [14-1:0] node2847;
	wire [14-1:0] node2849;
	wire [14-1:0] node2852;
	wire [14-1:0] node2853;
	wire [14-1:0] node2854;
	wire [14-1:0] node2858;
	wire [14-1:0] node2859;
	wire [14-1:0] node2861;

	assign outp = (inp[8]) ? node1426 : node1;
		assign node1 = (inp[7]) ? node739 : node2;
			assign node2 = (inp[5]) ? node384 : node3;
				assign node3 = (inp[4]) ? node195 : node4;
					assign node4 = (inp[9]) ? node114 : node5;
						assign node5 = (inp[3]) ? node53 : node6;
							assign node6 = (inp[0]) ? node28 : node7;
								assign node7 = (inp[13]) ? node21 : node8;
									assign node8 = (inp[11]) ? node18 : node9;
										assign node9 = (inp[12]) ? node15 : node10;
											assign node10 = (inp[6]) ? 14'b01111111111111 : node11;
												assign node11 = (inp[10]) ? 14'b01111111111111 : 14'b11111111111111;
											assign node15 = (inp[6]) ? 14'b00011111111111 : 14'b00111111111111;
										assign node18 = (inp[10]) ? 14'b00001111111111 : 14'b00011111111111;
									assign node21 = (inp[12]) ? node25 : node22;
										assign node22 = (inp[10]) ? 14'b00001111111111 : 14'b00011111111111;
										assign node25 = (inp[2]) ? 14'b00000111111111 : 14'b00001111111111;
								assign node28 = (inp[6]) ? node38 : node29;
									assign node29 = (inp[13]) ? 14'b00001111111111 : node30;
										assign node30 = (inp[2]) ? node32 : 14'b00011111111111;
											assign node32 = (inp[10]) ? 14'b00001111111111 : node33;
												assign node33 = (inp[12]) ? 14'b00001111111111 : 14'b00011111111111;
									assign node38 = (inp[1]) ? 14'b00000111111111 : node39;
										assign node39 = (inp[2]) ? node45 : node40;
											assign node40 = (inp[11]) ? 14'b00001111111111 : node41;
												assign node41 = (inp[12]) ? 14'b00001111111111 : 14'b00011111111111;
											assign node45 = (inp[12]) ? 14'b00000111111111 : node46;
												assign node46 = (inp[13]) ? node48 : 14'b00001111111111;
													assign node48 = (inp[10]) ? 14'b00000111111111 : 14'b00001111111111;
							assign node53 = (inp[11]) ? node89 : node54;
								assign node54 = (inp[6]) ? node76 : node55;
									assign node55 = (inp[0]) ? node71 : node56;
										assign node56 = (inp[12]) ? node64 : node57;
											assign node57 = (inp[1]) ? 14'b00001111111111 : node58;
												assign node58 = (inp[2]) ? 14'b00111111111111 : node59;
													assign node59 = (inp[13]) ? 14'b00111111111111 : 14'b01111111111111;
											assign node64 = (inp[10]) ? 14'b00001111111111 : node65;
												assign node65 = (inp[2]) ? node67 : 14'b00011111111111;
													assign node67 = (inp[1]) ? 14'b00001111111111 : 14'b00011111111111;
										assign node71 = (inp[10]) ? 14'b00001111111111 : node72;
											assign node72 = (inp[12]) ? 14'b00000111111111 : 14'b00001111111111;
									assign node76 = (inp[2]) ? node82 : node77;
										assign node77 = (inp[12]) ? 14'b00000111111111 : node78;
											assign node78 = (inp[0]) ? 14'b00001111111111 : 14'b00011111111111;
										assign node82 = (inp[12]) ? node84 : 14'b00000111111111;
											assign node84 = (inp[0]) ? 14'b00000011111111 : node85;
												assign node85 = (inp[1]) ? 14'b00000011111111 : 14'b00000111111111;
								assign node89 = (inp[2]) ? node105 : node90;
									assign node90 = (inp[12]) ? node98 : node91;
										assign node91 = (inp[13]) ? node95 : node92;
											assign node92 = (inp[6]) ? 14'b00001111111111 : 14'b00011111111111;
											assign node95 = (inp[6]) ? 14'b00001111111111 : 14'b00000111111111;
										assign node98 = (inp[0]) ? 14'b00000011111111 : node99;
											assign node99 = (inp[1]) ? node101 : 14'b00000111111111;
												assign node101 = (inp[6]) ? 14'b00000001111111 : 14'b00000111111111;
									assign node105 = (inp[13]) ? node109 : node106;
										assign node106 = (inp[10]) ? 14'b00000011111111 : 14'b00001111111111;
										assign node109 = (inp[0]) ? node111 : 14'b00000011111111;
											assign node111 = (inp[12]) ? 14'b00000001111111 : 14'b00000000111111;
						assign node114 = (inp[10]) ? node160 : node115;
							assign node115 = (inp[0]) ? node147 : node116;
								assign node116 = (inp[13]) ? node138 : node117;
									assign node117 = (inp[1]) ? node127 : node118;
										assign node118 = (inp[2]) ? 14'b00001111111111 : node119;
											assign node119 = (inp[6]) ? node123 : node120;
												assign node120 = (inp[3]) ? 14'b00111111111111 : 14'b01111111111111;
												assign node123 = (inp[11]) ? 14'b00001111111111 : 14'b00011111111111;
										assign node127 = (inp[12]) ? node129 : 14'b00001111111111;
											assign node129 = (inp[2]) ? 14'b00000011111111 : node130;
												assign node130 = (inp[3]) ? 14'b00000111111111 : node131;
													assign node131 = (inp[11]) ? node133 : 14'b00001111111111;
														assign node133 = (inp[6]) ? 14'b00000111111111 : 14'b00001111111111;
									assign node138 = (inp[11]) ? node142 : node139;
										assign node139 = (inp[12]) ? 14'b00000111111111 : 14'b00001111111111;
										assign node142 = (inp[2]) ? 14'b00000001111111 : node143;
											assign node143 = (inp[3]) ? 14'b00000011111111 : 14'b00000111111111;
								assign node147 = (inp[6]) ? node157 : node148;
									assign node148 = (inp[13]) ? node152 : node149;
										assign node149 = (inp[2]) ? 14'b00000011111111 : 14'b00000111111111;
										assign node152 = (inp[11]) ? 14'b00000111111111 : node153;
											assign node153 = (inp[3]) ? 14'b00000111111111 : 14'b00001111111111;
									assign node157 = (inp[1]) ? 14'b00000001111111 : 14'b00000011111111;
							assign node160 = (inp[2]) ? node184 : node161;
								assign node161 = (inp[12]) ? node171 : node162;
									assign node162 = (inp[1]) ? node166 : node163;
										assign node163 = (inp[13]) ? 14'b00001111111111 : 14'b00000111111111;
										assign node166 = (inp[13]) ? node168 : 14'b00000111111111;
											assign node168 = (inp[3]) ? 14'b00000011111111 : 14'b00000111111111;
									assign node171 = (inp[11]) ? node181 : node172;
										assign node172 = (inp[3]) ? node174 : 14'b00000111111111;
											assign node174 = (inp[0]) ? node178 : node175;
												assign node175 = (inp[1]) ? 14'b00000011111111 : 14'b00000111111111;
												assign node178 = (inp[6]) ? 14'b00000001111111 : 14'b00000011111111;
										assign node181 = (inp[6]) ? 14'b00000000111111 : 14'b00000011111111;
								assign node184 = (inp[1]) ? node192 : node185;
									assign node185 = (inp[12]) ? node187 : 14'b00000111111111;
										assign node187 = (inp[6]) ? node189 : 14'b00000011111111;
											assign node189 = (inp[13]) ? 14'b00000000011111 : 14'b00000001111111;
									assign node192 = (inp[12]) ? 14'b00000000111111 : 14'b00000001111111;
					assign node195 = (inp[3]) ? node283 : node196;
						assign node196 = (inp[12]) ? node240 : node197;
							assign node197 = (inp[2]) ? node225 : node198;
								assign node198 = (inp[0]) ? node208 : node199;
									assign node199 = (inp[1]) ? node205 : node200;
										assign node200 = (inp[10]) ? 14'b00001111111111 : node201;
											assign node201 = (inp[6]) ? 14'b00011111111111 : 14'b00111111111111;
										assign node205 = (inp[6]) ? 14'b00000111111111 : 14'b00001111111111;
									assign node208 = (inp[11]) ? node222 : node209;
										assign node209 = (inp[10]) ? node215 : node210;
											assign node210 = (inp[9]) ? node212 : 14'b00001111111111;
												assign node212 = (inp[1]) ? 14'b00000111111111 : 14'b00001111111111;
											assign node215 = (inp[13]) ? node217 : 14'b00001111111111;
												assign node217 = (inp[6]) ? node219 : 14'b00000111111111;
													assign node219 = (inp[9]) ? 14'b00000011111111 : 14'b00000111111111;
										assign node222 = (inp[10]) ? 14'b00000001111111 : 14'b00000111111111;
								assign node225 = (inp[1]) ? node235 : node226;
									assign node226 = (inp[10]) ? node232 : node227;
										assign node227 = (inp[0]) ? node229 : 14'b00000111111111;
											assign node229 = (inp[9]) ? 14'b00000111111111 : 14'b00001111111111;
										assign node232 = (inp[13]) ? 14'b00000011111111 : 14'b00000111111111;
									assign node235 = (inp[13]) ? 14'b00000011111111 : node236;
										assign node236 = (inp[11]) ? 14'b00000011111111 : 14'b00000111111111;
							assign node240 = (inp[13]) ? node262 : node241;
								assign node241 = (inp[6]) ? node249 : node242;
									assign node242 = (inp[1]) ? 14'b00001111111111 : node243;
										assign node243 = (inp[9]) ? node245 : 14'b00000111111111;
											assign node245 = (inp[11]) ? 14'b00000001111111 : 14'b00000111111111;
									assign node249 = (inp[0]) ? 14'b00000011111111 : node250;
										assign node250 = (inp[2]) ? node252 : 14'b00000111111111;
											assign node252 = (inp[10]) ? 14'b00000011111111 : node253;
												assign node253 = (inp[9]) ? 14'b00000011111111 : node254;
													assign node254 = (inp[1]) ? node256 : 14'b00000111111111;
														assign node256 = (inp[11]) ? 14'b00000011111111 : 14'b00000111111111;
								assign node262 = (inp[1]) ? node276 : node263;
									assign node263 = (inp[10]) ? node269 : node264;
										assign node264 = (inp[2]) ? node266 : 14'b00000111111111;
											assign node266 = (inp[6]) ? 14'b00000001111111 : 14'b00000111111111;
										assign node269 = (inp[9]) ? node273 : node270;
											assign node270 = (inp[11]) ? 14'b00000011111111 : 14'b00000111111111;
											assign node273 = (inp[11]) ? 14'b00000000111111 : 14'b00000001111111;
									assign node276 = (inp[10]) ? 14'b00000001111111 : node277;
										assign node277 = (inp[2]) ? node279 : 14'b00000011111111;
											assign node279 = (inp[11]) ? 14'b00000001111111 : 14'b00000000111111;
						assign node283 = (inp[9]) ? node333 : node284;
							assign node284 = (inp[1]) ? node316 : node285;
								assign node285 = (inp[6]) ? node303 : node286;
									assign node286 = (inp[10]) ? node292 : node287;
										assign node287 = (inp[0]) ? 14'b00000111111111 : node288;
											assign node288 = (inp[13]) ? 14'b00001111111111 : 14'b00000111111111;
										assign node292 = (inp[11]) ? 14'b00000000111111 : node293;
											assign node293 = (inp[0]) ? node295 : 14'b00000111111111;
												assign node295 = (inp[13]) ? 14'b00000001111111 : node296;
													assign node296 = (inp[2]) ? node298 : 14'b00000111111111;
														assign node298 = (inp[12]) ? 14'b00000011111111 : 14'b00000111111111;
									assign node303 = (inp[12]) ? node313 : node304;
										assign node304 = (inp[2]) ? node308 : node305;
											assign node305 = (inp[0]) ? 14'b00000111111111 : 14'b00000011111111;
											assign node308 = (inp[11]) ? 14'b00000001111111 : node309;
												assign node309 = (inp[0]) ? 14'b00000011111111 : 14'b00000111111111;
										assign node313 = (inp[2]) ? 14'b00000000111111 : 14'b00000001111111;
								assign node316 = (inp[0]) ? node320 : node317;
									assign node317 = (inp[2]) ? 14'b00000111111111 : 14'b00000011111111;
									assign node320 = (inp[6]) ? node328 : node321;
										assign node321 = (inp[12]) ? node323 : 14'b00000011111111;
											assign node323 = (inp[13]) ? 14'b00000001111111 : node324;
												assign node324 = (inp[11]) ? 14'b00000001111111 : 14'b00000011111111;
										assign node328 = (inp[10]) ? 14'b00000001111111 : node329;
											assign node329 = (inp[11]) ? 14'b00000000111111 : 14'b00000001111111;
							assign node333 = (inp[10]) ? node353 : node334;
								assign node334 = (inp[0]) ? node342 : node335;
									assign node335 = (inp[1]) ? node339 : node336;
										assign node336 = (inp[2]) ? 14'b00001111111111 : 14'b00000111111111;
										assign node339 = (inp[12]) ? 14'b00000001111111 : 14'b00000011111111;
									assign node342 = (inp[13]) ? node350 : node343;
										assign node343 = (inp[1]) ? 14'b00000001111111 : node344;
											assign node344 = (inp[6]) ? node346 : 14'b00000011111111;
												assign node346 = (inp[12]) ? 14'b00000011111111 : 14'b00000001111111;
										assign node350 = (inp[6]) ? 14'b00000000011111 : 14'b00000000111111;
								assign node353 = (inp[12]) ? node367 : node354;
									assign node354 = (inp[13]) ? node358 : node355;
										assign node355 = (inp[1]) ? 14'b00000001111111 : 14'b00000111111111;
										assign node358 = (inp[1]) ? 14'b00000000111111 : node359;
											assign node359 = (inp[11]) ? node361 : 14'b00000001111111;
												assign node361 = (inp[0]) ? node363 : 14'b00000001111111;
													assign node363 = (inp[6]) ? 14'b00000000111111 : 14'b00000001111111;
									assign node367 = (inp[11]) ? node377 : node368;
										assign node368 = (inp[0]) ? node370 : 14'b00000011111111;
											assign node370 = (inp[2]) ? 14'b00000000111111 : node371;
												assign node371 = (inp[6]) ? 14'b00000000111111 : node372;
													assign node372 = (inp[13]) ? 14'b00000000111111 : 14'b00000001111111;
										assign node377 = (inp[1]) ? node379 : 14'b00000000111111;
											assign node379 = (inp[13]) ? 14'b00000000011111 : node380;
												assign node380 = (inp[2]) ? 14'b00000000011111 : 14'b00000000111111;
				assign node384 = (inp[2]) ? node568 : node385;
					assign node385 = (inp[12]) ? node477 : node386;
						assign node386 = (inp[4]) ? node438 : node387;
							assign node387 = (inp[0]) ? node409 : node388;
								assign node388 = (inp[13]) ? node402 : node389;
									assign node389 = (inp[9]) ? node395 : node390;
										assign node390 = (inp[3]) ? node392 : 14'b00011111111111;
											assign node392 = (inp[1]) ? 14'b00011111111111 : 14'b00111111111111;
										assign node395 = (inp[10]) ? 14'b00000111111111 : node396;
											assign node396 = (inp[6]) ? 14'b00001111111111 : node397;
												assign node397 = (inp[11]) ? 14'b00001111111111 : 14'b00111111111111;
									assign node402 = (inp[11]) ? node406 : node403;
										assign node403 = (inp[3]) ? 14'b00000111111111 : 14'b00001111111111;
										assign node406 = (inp[10]) ? 14'b00000011111111 : 14'b00000111111111;
								assign node409 = (inp[6]) ? node423 : node410;
									assign node410 = (inp[1]) ? node420 : node411;
										assign node411 = (inp[13]) ? node417 : node412;
											assign node412 = (inp[3]) ? 14'b00001111111111 : node413;
												assign node413 = (inp[9]) ? 14'b00001111111111 : 14'b00111111111111;
											assign node417 = (inp[11]) ? 14'b00000111111111 : 14'b00001111111111;
										assign node420 = (inp[11]) ? 14'b00000111111111 : 14'b00000011111111;
									assign node423 = (inp[9]) ? node433 : node424;
										assign node424 = (inp[3]) ? node426 : 14'b00000111111111;
											assign node426 = (inp[1]) ? node430 : node427;
												assign node427 = (inp[11]) ? 14'b00000001111111 : 14'b00000011111111;
												assign node430 = (inp[11]) ? 14'b00000011111111 : 14'b00000111111111;
										assign node433 = (inp[13]) ? node435 : 14'b00000011111111;
											assign node435 = (inp[1]) ? 14'b00000001111111 : 14'b00000011111111;
							assign node438 = (inp[10]) ? node456 : node439;
								assign node439 = (inp[13]) ? node449 : node440;
									assign node440 = (inp[1]) ? node444 : node441;
										assign node441 = (inp[11]) ? 14'b00000111111111 : 14'b00001111111111;
										assign node444 = (inp[9]) ? 14'b00000011111111 : node445;
											assign node445 = (inp[0]) ? 14'b00000111111111 : 14'b00001111111111;
									assign node449 = (inp[6]) ? node453 : node450;
										assign node450 = (inp[1]) ? 14'b00000011111111 : 14'b00000111111111;
										assign node453 = (inp[3]) ? 14'b00000001111111 : 14'b00000011111111;
								assign node456 = (inp[0]) ? node466 : node457;
									assign node457 = (inp[13]) ? node461 : node458;
										assign node458 = (inp[6]) ? 14'b00000011111111 : 14'b00000111111111;
										assign node461 = (inp[1]) ? 14'b00000001111111 : node462;
											assign node462 = (inp[9]) ? 14'b00000011111111 : 14'b00000001111111;
									assign node466 = (inp[9]) ? node472 : node467;
										assign node467 = (inp[1]) ? node469 : 14'b00000011111111;
											assign node469 = (inp[3]) ? 14'b00000001111111 : 14'b00000011111111;
										assign node472 = (inp[3]) ? node474 : 14'b00000001111111;
											assign node474 = (inp[1]) ? 14'b00000000111111 : 14'b00000001111111;
						assign node477 = (inp[4]) ? node523 : node478;
							assign node478 = (inp[0]) ? node502 : node479;
								assign node479 = (inp[13]) ? node489 : node480;
									assign node480 = (inp[11]) ? node486 : node481;
										assign node481 = (inp[6]) ? node483 : 14'b00000111111111;
											assign node483 = (inp[10]) ? 14'b00000111111111 : 14'b00001111111111;
										assign node486 = (inp[10]) ? 14'b00000001111111 : 14'b00000111111111;
									assign node489 = (inp[10]) ? node495 : node490;
										assign node490 = (inp[11]) ? 14'b00000011111111 : node491;
											assign node491 = (inp[1]) ? 14'b00000011111111 : 14'b00000111111111;
										assign node495 = (inp[9]) ? node497 : 14'b00000111111111;
											assign node497 = (inp[6]) ? 14'b00000001111111 : node498;
												assign node498 = (inp[1]) ? 14'b00000001111111 : 14'b00000011111111;
								assign node502 = (inp[11]) ? node518 : node503;
									assign node503 = (inp[9]) ? node511 : node504;
										assign node504 = (inp[3]) ? node506 : 14'b00000111111111;
											assign node506 = (inp[1]) ? 14'b00000011111111 : node507;
												assign node507 = (inp[13]) ? 14'b00000011111111 : 14'b00000111111111;
										assign node511 = (inp[3]) ? node513 : 14'b00000011111111;
											assign node513 = (inp[6]) ? 14'b00000001111111 : node514;
												assign node514 = (inp[10]) ? 14'b00000001111111 : 14'b00000011111111;
									assign node518 = (inp[3]) ? 14'b00000001111111 : node519;
										assign node519 = (inp[10]) ? 14'b00000001111111 : 14'b00000011111111;
							assign node523 = (inp[6]) ? node545 : node524;
								assign node524 = (inp[3]) ? node536 : node525;
									assign node525 = (inp[1]) ? node531 : node526;
										assign node526 = (inp[0]) ? node528 : 14'b00001111111111;
											assign node528 = (inp[11]) ? 14'b00000011111111 : 14'b00000111111111;
										assign node531 = (inp[13]) ? 14'b00000001111111 : node532;
											assign node532 = (inp[0]) ? 14'b00000011111111 : 14'b00000111111111;
									assign node536 = (inp[11]) ? node542 : node537;
										assign node537 = (inp[9]) ? node539 : 14'b00000011111111;
											assign node539 = (inp[1]) ? 14'b00000001111111 : 14'b00000011111111;
										assign node542 = (inp[9]) ? 14'b00000000111111 : 14'b00000001111111;
								assign node545 = (inp[11]) ? node559 : node546;
									assign node546 = (inp[10]) ? node554 : node547;
										assign node547 = (inp[3]) ? 14'b00000001111111 : node548;
											assign node548 = (inp[0]) ? node550 : 14'b00000011111111;
												assign node550 = (inp[1]) ? 14'b00000001111111 : 14'b00000011111111;
										assign node554 = (inp[1]) ? node556 : 14'b00000001111111;
											assign node556 = (inp[3]) ? 14'b00000000111111 : 14'b00000001111111;
									assign node559 = (inp[3]) ? node563 : node560;
										assign node560 = (inp[0]) ? 14'b00000000111111 : 14'b00000001111111;
										assign node563 = (inp[13]) ? node565 : 14'b00000000011111;
											assign node565 = (inp[1]) ? 14'b00000000001111 : 14'b00000000011111;
					assign node568 = (inp[10]) ? node650 : node569;
						assign node569 = (inp[13]) ? node615 : node570;
							assign node570 = (inp[11]) ? node598 : node571;
								assign node571 = (inp[6]) ? node581 : node572;
									assign node572 = (inp[3]) ? node578 : node573;
										assign node573 = (inp[9]) ? 14'b00000111111111 : node574;
											assign node574 = (inp[1]) ? 14'b00001111111111 : 14'b00011111111111;
										assign node578 = (inp[9]) ? 14'b00000011111111 : 14'b00000111111111;
									assign node581 = (inp[12]) ? node589 : node582;
										assign node582 = (inp[4]) ? 14'b00000011111111 : node583;
											assign node583 = (inp[0]) ? 14'b00000011111111 : node584;
												assign node584 = (inp[1]) ? 14'b00000111111111 : 14'b00001111111111;
										assign node589 = (inp[1]) ? node591 : 14'b00000011111111;
											assign node591 = (inp[9]) ? 14'b00000001111111 : node592;
												assign node592 = (inp[0]) ? 14'b00000001111111 : node593;
													assign node593 = (inp[3]) ? 14'b00000011111111 : 14'b00000111111111;
								assign node598 = (inp[3]) ? node610 : node599;
									assign node599 = (inp[6]) ? node607 : node600;
										assign node600 = (inp[0]) ? node602 : 14'b00000111111111;
											assign node602 = (inp[4]) ? 14'b00000001111111 : node603;
												assign node603 = (inp[1]) ? 14'b00000011111111 : 14'b00000111111111;
										assign node607 = (inp[1]) ? 14'b00000001111111 : 14'b00000011111111;
									assign node610 = (inp[9]) ? node612 : 14'b00000001111111;
										assign node612 = (inp[1]) ? 14'b00000000111111 : 14'b00000001111111;
							assign node615 = (inp[3]) ? node635 : node616;
								assign node616 = (inp[1]) ? node624 : node617;
									assign node617 = (inp[0]) ? 14'b00000001111111 : node618;
										assign node618 = (inp[9]) ? 14'b00000011111111 : node619;
											assign node619 = (inp[11]) ? 14'b00000111111111 : 14'b00000011111111;
									assign node624 = (inp[4]) ? node628 : node625;
										assign node625 = (inp[9]) ? 14'b00000001111111 : 14'b00000011111111;
										assign node628 = (inp[12]) ? 14'b00000000111111 : node629;
											assign node629 = (inp[9]) ? node631 : 14'b00000011111111;
												assign node631 = (inp[0]) ? 14'b00000000111111 : 14'b00000001111111;
								assign node635 = (inp[12]) ? node643 : node636;
									assign node636 = (inp[11]) ? node638 : 14'b00000001111111;
										assign node638 = (inp[0]) ? node640 : 14'b00000001111111;
											assign node640 = (inp[4]) ? 14'b00000000111111 : 14'b00000001111111;
									assign node643 = (inp[9]) ? node647 : node644;
										assign node644 = (inp[1]) ? 14'b00000000011111 : 14'b00000001111111;
										assign node647 = (inp[0]) ? 14'b00000000011111 : 14'b00000000001111;
						assign node650 = (inp[1]) ? node694 : node651;
							assign node651 = (inp[9]) ? node673 : node652;
								assign node652 = (inp[13]) ? node664 : node653;
									assign node653 = (inp[0]) ? node657 : node654;
										assign node654 = (inp[12]) ? 14'b00000011111111 : 14'b00000111111111;
										assign node657 = (inp[4]) ? 14'b00000001111111 : node658;
											assign node658 = (inp[6]) ? node660 : 14'b00000011111111;
												assign node660 = (inp[3]) ? 14'b00000001111111 : 14'b00000011111111;
									assign node664 = (inp[6]) ? 14'b00000001111111 : node665;
										assign node665 = (inp[12]) ? node667 : 14'b00000011111111;
											assign node667 = (inp[3]) ? 14'b00000000111111 : node668;
												assign node668 = (inp[0]) ? 14'b00000001111111 : 14'b00000011111111;
								assign node673 = (inp[6]) ? node681 : node674;
									assign node674 = (inp[0]) ? node678 : node675;
										assign node675 = (inp[12]) ? 14'b00000001111111 : 14'b00000011111111;
										assign node678 = (inp[4]) ? 14'b00000000111111 : 14'b00000001111111;
									assign node681 = (inp[11]) ? node689 : node682;
										assign node682 = (inp[3]) ? node684 : 14'b00000001111111;
											assign node684 = (inp[0]) ? node686 : 14'b00000000111111;
												assign node686 = (inp[12]) ? 14'b00000000111111 : 14'b00000001111111;
										assign node689 = (inp[4]) ? 14'b00000000111111 : node690;
											assign node690 = (inp[0]) ? 14'b00000000011111 : 14'b00000000111111;
							assign node694 = (inp[12]) ? node712 : node695;
								assign node695 = (inp[13]) ? node705 : node696;
									assign node696 = (inp[3]) ? node700 : node697;
										assign node697 = (inp[11]) ? 14'b00000001111111 : 14'b00000011111111;
										assign node700 = (inp[9]) ? node702 : 14'b00000001111111;
											assign node702 = (inp[0]) ? 14'b00000000111111 : 14'b00000001111111;
									assign node705 = (inp[0]) ? 14'b00000000011111 : node706;
										assign node706 = (inp[6]) ? node708 : 14'b00000001111111;
											assign node708 = (inp[11]) ? 14'b00000000011111 : 14'b00000000111111;
								assign node712 = (inp[6]) ? node726 : node713;
									assign node713 = (inp[3]) ? node721 : node714;
										assign node714 = (inp[9]) ? node716 : 14'b00000011111111;
											assign node716 = (inp[4]) ? node718 : 14'b00000001111111;
												assign node718 = (inp[0]) ? 14'b00000000111111 : 14'b00000001111111;
										assign node721 = (inp[0]) ? node723 : 14'b00000000111111;
											assign node723 = (inp[9]) ? 14'b00000000011111 : 14'b00000000111111;
									assign node726 = (inp[9]) ? node734 : node727;
										assign node727 = (inp[0]) ? 14'b00000000011111 : node728;
											assign node728 = (inp[11]) ? node730 : 14'b00000000111111;
												assign node730 = (inp[3]) ? 14'b00000000011111 : 14'b00000000111111;
										assign node734 = (inp[0]) ? 14'b00000000001111 : node735;
											assign node735 = (inp[13]) ? 14'b00000000011111 : 14'b00000000001111;
			assign node739 = (inp[0]) ? node1105 : node740;
				assign node740 = (inp[1]) ? node922 : node741;
					assign node741 = (inp[3]) ? node823 : node742;
						assign node742 = (inp[6]) ? node786 : node743;
							assign node743 = (inp[2]) ? node765 : node744;
								assign node744 = (inp[10]) ? node752 : node745;
									assign node745 = (inp[9]) ? node747 : 14'b00001111111111;
										assign node747 = (inp[4]) ? 14'b00001111111111 : node748;
											assign node748 = (inp[11]) ? 14'b00001111111111 : 14'b00011111111111;
									assign node752 = (inp[5]) ? node762 : node753;
										assign node753 = (inp[4]) ? node759 : node754;
											assign node754 = (inp[9]) ? 14'b00001111111111 : node755;
												assign node755 = (inp[11]) ? 14'b00011111111111 : 14'b00001111111111;
											assign node759 = (inp[13]) ? 14'b00000111111111 : 14'b00001111111111;
										assign node762 = (inp[12]) ? 14'b00000011111111 : 14'b00000111111111;
								assign node765 = (inp[12]) ? node777 : node766;
									assign node766 = (inp[13]) ? 14'b00000111111111 : node767;
										assign node767 = (inp[5]) ? 14'b00000011111111 : node768;
											assign node768 = (inp[4]) ? node772 : node769;
												assign node769 = (inp[11]) ? 14'b00001111111111 : 14'b00011111111111;
												assign node772 = (inp[11]) ? 14'b00000111111111 : 14'b00001111111111;
									assign node777 = (inp[4]) ? node783 : node778;
										assign node778 = (inp[5]) ? 14'b00000111111111 : node779;
											assign node779 = (inp[10]) ? 14'b00000111111111 : 14'b00000011111111;
										assign node783 = (inp[5]) ? 14'b00000000111111 : 14'b00000011111111;
							assign node786 = (inp[13]) ? node808 : node787;
								assign node787 = (inp[10]) ? node797 : node788;
									assign node788 = (inp[12]) ? node792 : node789;
										assign node789 = (inp[9]) ? 14'b00000111111111 : 14'b00001111111111;
										assign node792 = (inp[9]) ? node794 : 14'b00000111111111;
											assign node794 = (inp[2]) ? 14'b00000011111111 : 14'b00000111111111;
									assign node797 = (inp[12]) ? node803 : node798;
										assign node798 = (inp[9]) ? node800 : 14'b00000111111111;
											assign node800 = (inp[2]) ? 14'b00000111111111 : 14'b00000011111111;
										assign node803 = (inp[2]) ? 14'b00000011111111 : node804;
											assign node804 = (inp[5]) ? 14'b00000000111111 : 14'b00001111111111;
								assign node808 = (inp[12]) ? node814 : node809;
									assign node809 = (inp[5]) ? node811 : 14'b00000011111111;
										assign node811 = (inp[11]) ? 14'b00000000111111 : 14'b00000011111111;
									assign node814 = (inp[9]) ? node818 : node815;
										assign node815 = (inp[11]) ? 14'b00000001111111 : 14'b00000011111111;
										assign node818 = (inp[2]) ? node820 : 14'b00000001111111;
											assign node820 = (inp[10]) ? 14'b00000000011111 : 14'b00000000111111;
						assign node823 = (inp[5]) ? node863 : node824;
							assign node824 = (inp[6]) ? node846 : node825;
								assign node825 = (inp[10]) ? node837 : node826;
									assign node826 = (inp[9]) ? node834 : node827;
										assign node827 = (inp[12]) ? node829 : 14'b00011111111111;
											assign node829 = (inp[13]) ? node831 : 14'b00000111111111;
												assign node831 = (inp[2]) ? 14'b00000111111111 : 14'b00001111111111;
										assign node834 = (inp[12]) ? 14'b00000011111111 : 14'b00000111111111;
									assign node837 = (inp[13]) ? node839 : 14'b00000111111111;
										assign node839 = (inp[4]) ? node841 : 14'b00000011111111;
											assign node841 = (inp[2]) ? node843 : 14'b00000001111111;
												assign node843 = (inp[11]) ? 14'b00000001111111 : 14'b00000011111111;
								assign node846 = (inp[4]) ? node858 : node847;
									assign node847 = (inp[2]) ? node853 : node848;
										assign node848 = (inp[9]) ? 14'b00000011111111 : node849;
											assign node849 = (inp[12]) ? 14'b00000011111111 : 14'b00000111111111;
										assign node853 = (inp[12]) ? node855 : 14'b00000011111111;
											assign node855 = (inp[13]) ? 14'b00000001111111 : 14'b00000011111111;
									assign node858 = (inp[12]) ? 14'b00000001111111 : node859;
										assign node859 = (inp[9]) ? 14'b00000011111111 : 14'b00000001111111;
							assign node863 = (inp[13]) ? node895 : node864;
								assign node864 = (inp[10]) ? node884 : node865;
									assign node865 = (inp[11]) ? node871 : node866;
										assign node866 = (inp[4]) ? node868 : 14'b00000111111111;
											assign node868 = (inp[9]) ? 14'b00000011111111 : 14'b00000111111111;
										assign node871 = (inp[9]) ? node879 : node872;
											assign node872 = (inp[4]) ? node876 : node873;
												assign node873 = (inp[2]) ? 14'b00000111111111 : 14'b00000011111111;
												assign node876 = (inp[12]) ? 14'b00000001111111 : 14'b00000011111111;
											assign node879 = (inp[2]) ? 14'b00000001111111 : node880;
												assign node880 = (inp[4]) ? 14'b00000001111111 : 14'b00000011111111;
									assign node884 = (inp[6]) ? node886 : 14'b00000011111111;
										assign node886 = (inp[9]) ? node892 : node887;
											assign node887 = (inp[4]) ? node889 : 14'b00000001111111;
												assign node889 = (inp[2]) ? 14'b00000000111111 : 14'b00000001111111;
											assign node892 = (inp[11]) ? 14'b00000000011111 : 14'b00000000111111;
								assign node895 = (inp[11]) ? node907 : node896;
									assign node896 = (inp[4]) ? node900 : node897;
										assign node897 = (inp[6]) ? 14'b00000000011111 : 14'b00000011111111;
										assign node900 = (inp[12]) ? node902 : 14'b00000001111111;
											assign node902 = (inp[10]) ? 14'b00000000111111 : node903;
												assign node903 = (inp[9]) ? 14'b00000000111111 : 14'b00000001111111;
									assign node907 = (inp[4]) ? node915 : node908;
										assign node908 = (inp[6]) ? 14'b00000000111111 : node909;
											assign node909 = (inp[2]) ? node911 : 14'b00000001111111;
												assign node911 = (inp[9]) ? 14'b00000000111111 : 14'b00000001111111;
										assign node915 = (inp[10]) ? node917 : 14'b00000000111111;
											assign node917 = (inp[2]) ? 14'b00000000011111 : node918;
												assign node918 = (inp[12]) ? 14'b00000000011111 : 14'b00000000111111;
					assign node922 = (inp[12]) ? node1028 : node923;
						assign node923 = (inp[6]) ? node981 : node924;
							assign node924 = (inp[3]) ? node950 : node925;
								assign node925 = (inp[13]) ? node935 : node926;
									assign node926 = (inp[4]) ? node932 : node927;
										assign node927 = (inp[2]) ? 14'b00000111111111 : node928;
											assign node928 = (inp[5]) ? 14'b00000011111111 : 14'b00000111111111;
										assign node932 = (inp[11]) ? 14'b00000011111111 : 14'b00000111111111;
									assign node935 = (inp[10]) ? node943 : node936;
										assign node936 = (inp[9]) ? 14'b00000001111111 : node937;
											assign node937 = (inp[2]) ? node939 : 14'b00000111111111;
												assign node939 = (inp[4]) ? 14'b00000011111111 : 14'b00000111111111;
										assign node943 = (inp[4]) ? 14'b00000000111111 : node944;
											assign node944 = (inp[9]) ? 14'b00000001111111 : node945;
												assign node945 = (inp[11]) ? 14'b00000001111111 : 14'b00000011111111;
								assign node950 = (inp[10]) ? node970 : node951;
									assign node951 = (inp[2]) ? node965 : node952;
										assign node952 = (inp[9]) ? node960 : node953;
											assign node953 = (inp[5]) ? 14'b00000011111111 : node954;
												assign node954 = (inp[4]) ? 14'b00000111111111 : node955;
													assign node955 = (inp[11]) ? 14'b00000111111111 : 14'b00001111111111;
											assign node960 = (inp[11]) ? node962 : 14'b00000011111111;
												assign node962 = (inp[4]) ? 14'b00000001111111 : 14'b00000011111111;
										assign node965 = (inp[13]) ? 14'b00000001111111 : node966;
											assign node966 = (inp[5]) ? 14'b00000001111111 : 14'b00000011111111;
									assign node970 = (inp[11]) ? node974 : node971;
										assign node971 = (inp[9]) ? 14'b00000001111111 : 14'b00000011111111;
										assign node974 = (inp[5]) ? node976 : 14'b00000001111111;
											assign node976 = (inp[4]) ? node978 : 14'b00000001111111;
												assign node978 = (inp[13]) ? 14'b00000000111111 : 14'b00000001111111;
							assign node981 = (inp[9]) ? node1011 : node982;
								assign node982 = (inp[3]) ? node992 : node983;
									assign node983 = (inp[10]) ? node989 : node984;
										assign node984 = (inp[11]) ? 14'b00000011111111 : node985;
											assign node985 = (inp[5]) ? 14'b00001111111111 : 14'b00000111111111;
										assign node989 = (inp[5]) ? 14'b00000011111111 : 14'b00000001111111;
									assign node992 = (inp[13]) ? node1000 : node993;
										assign node993 = (inp[2]) ? node997 : node994;
											assign node994 = (inp[10]) ? 14'b00000011111111 : 14'b00000111111111;
											assign node997 = (inp[5]) ? 14'b00000000111111 : 14'b00000001111111;
										assign node1000 = (inp[2]) ? 14'b00000000111111 : node1001;
											assign node1001 = (inp[11]) ? node1003 : 14'b00000001111111;
												assign node1003 = (inp[10]) ? node1005 : 14'b00000001111111;
													assign node1005 = (inp[4]) ? 14'b00000000111111 : node1006;
														assign node1006 = (inp[5]) ? 14'b00000000111111 : 14'b00000001111111;
								assign node1011 = (inp[13]) ? node1021 : node1012;
									assign node1012 = (inp[11]) ? node1016 : node1013;
										assign node1013 = (inp[5]) ? 14'b00000001111111 : 14'b00000011111111;
										assign node1016 = (inp[2]) ? 14'b00000000111111 : node1017;
											assign node1017 = (inp[4]) ? 14'b00000000111111 : 14'b00000001111111;
									assign node1021 = (inp[3]) ? node1023 : 14'b00000000111111;
										assign node1023 = (inp[10]) ? node1025 : 14'b00000000111111;
											assign node1025 = (inp[11]) ? 14'b00000000011111 : 14'b00000000001111;
						assign node1028 = (inp[11]) ? node1066 : node1029;
							assign node1029 = (inp[5]) ? node1049 : node1030;
								assign node1030 = (inp[2]) ? node1044 : node1031;
									assign node1031 = (inp[3]) ? 14'b00000011111111 : node1032;
										assign node1032 = (inp[4]) ? node1036 : node1033;
											assign node1033 = (inp[13]) ? 14'b00001111111111 : 14'b00000111111111;
											assign node1036 = (inp[10]) ? node1040 : node1037;
												assign node1037 = (inp[9]) ? 14'b00000011111111 : 14'b00000111111111;
												assign node1040 = (inp[9]) ? 14'b00000000111111 : 14'b00000011111111;
									assign node1044 = (inp[4]) ? node1046 : 14'b00000011111111;
										assign node1046 = (inp[9]) ? 14'b00000000111111 : 14'b00000001111111;
								assign node1049 = (inp[6]) ? node1061 : node1050;
									assign node1050 = (inp[13]) ? 14'b00000000111111 : node1051;
										assign node1051 = (inp[4]) ? node1055 : node1052;
											assign node1052 = (inp[9]) ? 14'b00000001111111 : 14'b00000011111111;
											assign node1055 = (inp[3]) ? node1057 : 14'b00000001111111;
												assign node1057 = (inp[9]) ? 14'b00000000111111 : 14'b00000001111111;
									assign node1061 = (inp[2]) ? 14'b00000000011111 : node1062;
										assign node1062 = (inp[3]) ? 14'b00000000111111 : 14'b00000000011111;
							assign node1066 = (inp[4]) ? node1080 : node1067;
								assign node1067 = (inp[6]) ? node1073 : node1068;
									assign node1068 = (inp[13]) ? 14'b00000001111111 : node1069;
										assign node1069 = (inp[3]) ? 14'b00000000111111 : 14'b00000011111111;
									assign node1073 = (inp[9]) ? node1075 : 14'b00000000011111;
										assign node1075 = (inp[2]) ? node1077 : 14'b00000000111111;
											assign node1077 = (inp[13]) ? 14'b00000000111111 : 14'b00000001111111;
								assign node1080 = (inp[9]) ? node1094 : node1081;
									assign node1081 = (inp[10]) ? node1087 : node1082;
										assign node1082 = (inp[5]) ? 14'b00000000111111 : node1083;
											assign node1083 = (inp[3]) ? 14'b00000001111111 : 14'b00000011111111;
										assign node1087 = (inp[13]) ? 14'b00000000001111 : node1088;
											assign node1088 = (inp[6]) ? 14'b00000000111111 : node1089;
												assign node1089 = (inp[5]) ? 14'b00000000111111 : 14'b00000001111111;
									assign node1094 = (inp[6]) ? node1098 : node1095;
										assign node1095 = (inp[13]) ? 14'b00000000011111 : 14'b00000000111111;
										assign node1098 = (inp[10]) ? node1100 : 14'b00000000011111;
											assign node1100 = (inp[13]) ? node1102 : 14'b00000000001111;
												assign node1102 = (inp[5]) ? 14'b00000000001111 : 14'b00000000011111;
				assign node1105 = (inp[9]) ? node1245 : node1106;
					assign node1106 = (inp[5]) ? node1176 : node1107;
						assign node1107 = (inp[3]) ? node1145 : node1108;
							assign node1108 = (inp[2]) ? node1130 : node1109;
								assign node1109 = (inp[12]) ? node1119 : node1110;
									assign node1110 = (inp[10]) ? node1114 : node1111;
										assign node1111 = (inp[1]) ? 14'b00000111111111 : 14'b00001111111111;
										assign node1114 = (inp[11]) ? node1116 : 14'b00000111111111;
											assign node1116 = (inp[6]) ? 14'b00000011111111 : 14'b00000111111111;
									assign node1119 = (inp[13]) ? node1127 : node1120;
										assign node1120 = (inp[1]) ? node1122 : 14'b00000111111111;
											assign node1122 = (inp[11]) ? node1124 : 14'b00000111111111;
												assign node1124 = (inp[10]) ? 14'b00000011111111 : 14'b00000111111111;
										assign node1127 = (inp[10]) ? 14'b00000000111111 : 14'b00000011111111;
								assign node1130 = (inp[11]) ? node1138 : node1131;
									assign node1131 = (inp[13]) ? node1135 : node1132;
										assign node1132 = (inp[4]) ? 14'b00000111111111 : 14'b00001111111111;
										assign node1135 = (inp[12]) ? 14'b00000001111111 : 14'b00000011111111;
									assign node1138 = (inp[4]) ? node1142 : node1139;
										assign node1139 = (inp[6]) ? 14'b00000001111111 : 14'b00000011111111;
										assign node1142 = (inp[1]) ? 14'b00000000111111 : 14'b00000001111111;
							assign node1145 = (inp[10]) ? node1163 : node1146;
								assign node1146 = (inp[11]) ? node1156 : node1147;
									assign node1147 = (inp[6]) ? node1153 : node1148;
										assign node1148 = (inp[4]) ? node1150 : 14'b00000111111111;
											assign node1150 = (inp[1]) ? 14'b00000001111111 : 14'b00000111111111;
										assign node1153 = (inp[2]) ? 14'b00000001111111 : 14'b00000011111111;
									assign node1156 = (inp[1]) ? node1158 : 14'b00000011111111;
										assign node1158 = (inp[4]) ? node1160 : 14'b00000001111111;
											assign node1160 = (inp[6]) ? 14'b00000000111111 : 14'b00000001111111;
								assign node1163 = (inp[13]) ? node1171 : node1164;
									assign node1164 = (inp[1]) ? node1168 : node1165;
										assign node1165 = (inp[11]) ? 14'b00000111111111 : 14'b00000011111111;
										assign node1168 = (inp[4]) ? 14'b00000000011111 : 14'b00000000111111;
									assign node1171 = (inp[11]) ? 14'b00000000011111 : node1172;
										assign node1172 = (inp[12]) ? 14'b00000000011111 : 14'b00000000111111;
						assign node1176 = (inp[12]) ? node1214 : node1177;
							assign node1177 = (inp[4]) ? node1195 : node1178;
								assign node1178 = (inp[6]) ? node1190 : node1179;
									assign node1179 = (inp[10]) ? node1185 : node1180;
										assign node1180 = (inp[13]) ? 14'b00000011111111 : node1181;
											assign node1181 = (inp[1]) ? 14'b00000011111111 : 14'b00000111111111;
										assign node1185 = (inp[3]) ? node1187 : 14'b00000011111111;
											assign node1187 = (inp[11]) ? 14'b00000001111111 : 14'b00000011111111;
									assign node1190 = (inp[1]) ? 14'b00000000111111 : node1191;
										assign node1191 = (inp[11]) ? 14'b00000001111111 : 14'b00000011111111;
								assign node1195 = (inp[10]) ? node1203 : node1196;
									assign node1196 = (inp[3]) ? node1200 : node1197;
										assign node1197 = (inp[11]) ? 14'b00000001111111 : 14'b00000011111111;
										assign node1200 = (inp[6]) ? 14'b00000001111111 : 14'b00000000111111;
									assign node1203 = (inp[13]) ? node1211 : node1204;
										assign node1204 = (inp[6]) ? 14'b00000000111111 : node1205;
											assign node1205 = (inp[11]) ? node1207 : 14'b00000001111111;
												assign node1207 = (inp[1]) ? 14'b00000000111111 : 14'b00000001111111;
										assign node1211 = (inp[3]) ? 14'b00000000111111 : 14'b00000000011111;
							assign node1214 = (inp[10]) ? node1234 : node1215;
								assign node1215 = (inp[6]) ? node1227 : node1216;
									assign node1216 = (inp[1]) ? node1220 : node1217;
										assign node1217 = (inp[13]) ? 14'b00000001111111 : 14'b00000011111111;
										assign node1220 = (inp[4]) ? node1222 : 14'b00000001111111;
											assign node1222 = (inp[13]) ? 14'b00000000011111 : node1223;
												assign node1223 = (inp[2]) ? 14'b00000000111111 : 14'b00000001111111;
									assign node1227 = (inp[11]) ? node1231 : node1228;
										assign node1228 = (inp[13]) ? 14'b00000000111111 : 14'b00000111111111;
										assign node1231 = (inp[13]) ? 14'b00000000011111 : 14'b00000000111111;
								assign node1234 = (inp[4]) ? node1240 : node1235;
									assign node1235 = (inp[1]) ? node1237 : 14'b00000000111111;
										assign node1237 = (inp[13]) ? 14'b00000000111111 : 14'b00000001111111;
									assign node1240 = (inp[3]) ? node1242 : 14'b00000000111111;
										assign node1242 = (inp[1]) ? 14'b00000000001111 : 14'b00000000011111;
					assign node1245 = (inp[11]) ? node1325 : node1246;
						assign node1246 = (inp[12]) ? node1292 : node1247;
							assign node1247 = (inp[4]) ? node1263 : node1248;
								assign node1248 = (inp[10]) ? node1254 : node1249;
									assign node1249 = (inp[1]) ? 14'b00000011111111 : node1250;
										assign node1250 = (inp[2]) ? 14'b00000011111111 : 14'b00000111111111;
									assign node1254 = (inp[3]) ? node1260 : node1255;
										assign node1255 = (inp[13]) ? 14'b00000001111111 : node1256;
											assign node1256 = (inp[6]) ? 14'b00000011111111 : 14'b00000111111111;
										assign node1260 = (inp[5]) ? 14'b00000001111111 : 14'b00000000111111;
								assign node1263 = (inp[6]) ? node1281 : node1264;
									assign node1264 = (inp[2]) ? node1272 : node1265;
										assign node1265 = (inp[3]) ? node1269 : node1266;
											assign node1266 = (inp[5]) ? 14'b00000011111111 : 14'b00000111111111;
											assign node1269 = (inp[1]) ? 14'b00000001111111 : 14'b00000011111111;
										assign node1272 = (inp[10]) ? node1274 : 14'b00000001111111;
											assign node1274 = (inp[3]) ? node1276 : 14'b00000001111111;
												assign node1276 = (inp[5]) ? node1278 : 14'b00000000111111;
													assign node1278 = (inp[1]) ? 14'b00000000011111 : 14'b00000000111111;
									assign node1281 = (inp[5]) ? node1287 : node1282;
										assign node1282 = (inp[2]) ? 14'b00000000111111 : node1283;
											assign node1283 = (inp[13]) ? 14'b00000000011111 : 14'b00000000111111;
										assign node1287 = (inp[13]) ? node1289 : 14'b00000000011111;
											assign node1289 = (inp[2]) ? 14'b00000000001111 : 14'b00000000011111;
							assign node1292 = (inp[1]) ? node1302 : node1293;
								assign node1293 = (inp[3]) ? node1297 : node1294;
									assign node1294 = (inp[5]) ? 14'b00000001111111 : 14'b00000000111111;
									assign node1297 = (inp[5]) ? node1299 : 14'b00000001111111;
										assign node1299 = (inp[2]) ? 14'b00000000111111 : 14'b00000000011111;
								assign node1302 = (inp[5]) ? node1314 : node1303;
									assign node1303 = (inp[2]) ? node1307 : node1304;
										assign node1304 = (inp[3]) ? 14'b00000000111111 : 14'b00000001111111;
										assign node1307 = (inp[3]) ? 14'b00000000011111 : node1308;
											assign node1308 = (inp[4]) ? 14'b00000000111111 : node1309;
												assign node1309 = (inp[13]) ? 14'b00000000011111 : 14'b00000000111111;
									assign node1314 = (inp[13]) ? node1322 : node1315;
										assign node1315 = (inp[3]) ? node1319 : node1316;
											assign node1316 = (inp[6]) ? 14'b00000000011111 : 14'b00000000111111;
											assign node1319 = (inp[2]) ? 14'b00000000001111 : 14'b00000000011111;
										assign node1322 = (inp[10]) ? 14'b00000000001111 : 14'b00000000011111;
						assign node1325 = (inp[1]) ? node1373 : node1326;
							assign node1326 = (inp[6]) ? node1354 : node1327;
								assign node1327 = (inp[13]) ? node1339 : node1328;
									assign node1328 = (inp[10]) ? 14'b00000111111111 : node1329;
										assign node1329 = (inp[5]) ? 14'b00000001111111 : node1330;
											assign node1330 = (inp[2]) ? node1332 : 14'b00000011111111;
												assign node1332 = (inp[3]) ? 14'b00000001111111 : node1333;
													assign node1333 = (inp[4]) ? 14'b00000001111111 : 14'b00000011111111;
									assign node1339 = (inp[3]) ? node1347 : node1340;
										assign node1340 = (inp[2]) ? node1342 : 14'b00000000111111;
											assign node1342 = (inp[10]) ? 14'b00000001111111 : node1343;
												assign node1343 = (inp[4]) ? 14'b00000001111111 : 14'b00000011111111;
										assign node1347 = (inp[12]) ? 14'b00000000011111 : node1348;
											assign node1348 = (inp[2]) ? node1350 : 14'b00000001111111;
												assign node1350 = (inp[4]) ? 14'b00000000011111 : 14'b00000000111111;
								assign node1354 = (inp[13]) ? node1364 : node1355;
									assign node1355 = (inp[10]) ? node1361 : node1356;
										assign node1356 = (inp[2]) ? 14'b00000000111111 : node1357;
											assign node1357 = (inp[5]) ? 14'b00000000011111 : 14'b00000000111111;
										assign node1361 = (inp[5]) ? 14'b00000000001111 : 14'b00000000011111;
									assign node1364 = (inp[5]) ? node1368 : node1365;
										assign node1365 = (inp[10]) ? 14'b00000000011111 : 14'b00000000001111;
										assign node1368 = (inp[12]) ? 14'b00000000000111 : node1369;
											assign node1369 = (inp[3]) ? 14'b00000000000111 : 14'b00000000001111;
							assign node1373 = (inp[3]) ? node1401 : node1374;
								assign node1374 = (inp[6]) ? node1386 : node1375;
									assign node1375 = (inp[5]) ? node1377 : 14'b00000000111111;
										assign node1377 = (inp[2]) ? node1379 : 14'b00000000111111;
											assign node1379 = (inp[12]) ? 14'b00000000011111 : node1380;
												assign node1380 = (inp[10]) ? node1382 : 14'b00000000111111;
													assign node1382 = (inp[4]) ? 14'b00000000011111 : 14'b00000000111111;
									assign node1386 = (inp[4]) ? node1392 : node1387;
										assign node1387 = (inp[5]) ? node1389 : 14'b00000000111111;
											assign node1389 = (inp[12]) ? 14'b00000000011111 : 14'b00000000111111;
										assign node1392 = (inp[10]) ? node1396 : node1393;
											assign node1393 = (inp[13]) ? 14'b00000000001111 : 14'b00000000111111;
											assign node1396 = (inp[2]) ? node1398 : 14'b00000000001111;
												assign node1398 = (inp[13]) ? 14'b00000000000011 : 14'b00000000000111;
								assign node1401 = (inp[2]) ? node1411 : node1402;
									assign node1402 = (inp[5]) ? 14'b00000000001111 : node1403;
										assign node1403 = (inp[10]) ? node1407 : node1404;
											assign node1404 = (inp[12]) ? 14'b00000000011111 : 14'b00000000111111;
											assign node1407 = (inp[6]) ? 14'b00000000001111 : 14'b00000000011111;
									assign node1411 = (inp[4]) ? node1415 : node1412;
										assign node1412 = (inp[10]) ? 14'b00000000001111 : 14'b00000000011111;
										assign node1415 = (inp[13]) ? node1421 : node1416;
											assign node1416 = (inp[6]) ? node1418 : 14'b00000000001111;
												assign node1418 = (inp[12]) ? 14'b00000000000111 : 14'b00000000001111;
											assign node1421 = (inp[12]) ? 14'b00000000000111 : node1422;
												assign node1422 = (inp[10]) ? 14'b00000000000111 : 14'b00000000001111;
		assign node1426 = (inp[11]) ? node2138 : node1427;
			assign node1427 = (inp[6]) ? node1765 : node1428;
				assign node1428 = (inp[12]) ? node1610 : node1429;
					assign node1429 = (inp[3]) ? node1527 : node1430;
						assign node1430 = (inp[4]) ? node1478 : node1431;
							assign node1431 = (inp[2]) ? node1461 : node1432;
								assign node1432 = (inp[13]) ? node1450 : node1433;
									assign node1433 = (inp[9]) ? node1443 : node1434;
										assign node1434 = (inp[1]) ? node1438 : node1435;
											assign node1435 = (inp[5]) ? 14'b00011111111111 : 14'b00111111111111;
											assign node1438 = (inp[10]) ? 14'b00001111111111 : node1439;
												assign node1439 = (inp[7]) ? 14'b00001111111111 : 14'b00011111111111;
										assign node1443 = (inp[5]) ? node1447 : node1444;
											assign node1444 = (inp[0]) ? 14'b00001111111111 : 14'b00011111111111;
											assign node1447 = (inp[0]) ? 14'b00000011111111 : 14'b00000111111111;
									assign node1450 = (inp[1]) ? node1458 : node1451;
										assign node1451 = (inp[5]) ? 14'b00000111111111 : node1452;
											assign node1452 = (inp[7]) ? node1454 : 14'b00001111111111;
												assign node1454 = (inp[9]) ? 14'b00000111111111 : 14'b00001111111111;
										assign node1458 = (inp[0]) ? 14'b00000011111111 : 14'b00000111111111;
								assign node1461 = (inp[9]) ? node1469 : node1462;
									assign node1462 = (inp[13]) ? node1464 : 14'b00000011111111;
										assign node1464 = (inp[0]) ? 14'b00000111111111 : node1465;
											assign node1465 = (inp[7]) ? 14'b00000111111111 : 14'b00001111111111;
									assign node1469 = (inp[7]) ? 14'b00000011111111 : node1470;
										assign node1470 = (inp[13]) ? node1472 : 14'b00000111111111;
											assign node1472 = (inp[0]) ? 14'b00000011111111 : node1473;
												assign node1473 = (inp[10]) ? 14'b00000011111111 : 14'b00000111111111;
							assign node1478 = (inp[5]) ? node1498 : node1479;
								assign node1479 = (inp[13]) ? node1489 : node1480;
									assign node1480 = (inp[2]) ? node1486 : node1481;
										assign node1481 = (inp[9]) ? 14'b00000111111111 : node1482;
											assign node1482 = (inp[1]) ? 14'b00001111111111 : 14'b00011111111111;
										assign node1486 = (inp[7]) ? 14'b00000011111111 : 14'b00000111111111;
									assign node1489 = (inp[0]) ? node1493 : node1490;
										assign node1490 = (inp[1]) ? 14'b00000011111111 : 14'b00000111111111;
										assign node1493 = (inp[2]) ? node1495 : 14'b00000011111111;
											assign node1495 = (inp[1]) ? 14'b00000001111111 : 14'b00000011111111;
								assign node1498 = (inp[1]) ? node1514 : node1499;
									assign node1499 = (inp[10]) ? node1507 : node1500;
										assign node1500 = (inp[2]) ? node1502 : 14'b00000111111111;
											assign node1502 = (inp[0]) ? node1504 : 14'b00000111111111;
												assign node1504 = (inp[13]) ? 14'b00000011111111 : 14'b00000111111111;
										assign node1507 = (inp[13]) ? node1509 : 14'b00000011111111;
											assign node1509 = (inp[9]) ? 14'b00000001111111 : node1510;
												assign node1510 = (inp[0]) ? 14'b00000001111111 : 14'b00000011111111;
									assign node1514 = (inp[9]) ? node1522 : node1515;
										assign node1515 = (inp[2]) ? node1517 : 14'b00000011111111;
											assign node1517 = (inp[13]) ? node1519 : 14'b00000001111111;
												assign node1519 = (inp[0]) ? 14'b00000000111111 : 14'b00000001111111;
										assign node1522 = (inp[2]) ? 14'b00000000111111 : node1523;
											assign node1523 = (inp[7]) ? 14'b00000000111111 : 14'b00000001111111;
						assign node1527 = (inp[0]) ? node1577 : node1528;
							assign node1528 = (inp[4]) ? node1554 : node1529;
								assign node1529 = (inp[13]) ? node1541 : node1530;
									assign node1530 = (inp[7]) ? node1532 : 14'b00001111111111;
										assign node1532 = (inp[10]) ? node1536 : node1533;
											assign node1533 = (inp[2]) ? 14'b00000111111111 : 14'b00001111111111;
											assign node1536 = (inp[9]) ? 14'b00000011111111 : node1537;
												assign node1537 = (inp[2]) ? 14'b00000011111111 : 14'b00000111111111;
									assign node1541 = (inp[7]) ? node1549 : node1542;
										assign node1542 = (inp[5]) ? 14'b00000011111111 : node1543;
											assign node1543 = (inp[9]) ? 14'b00000111111111 : node1544;
												assign node1544 = (inp[2]) ? 14'b00000111111111 : 14'b00001111111111;
										assign node1549 = (inp[2]) ? 14'b00000001111111 : node1550;
											assign node1550 = (inp[1]) ? 14'b00000001111111 : 14'b00000011111111;
								assign node1554 = (inp[10]) ? node1568 : node1555;
									assign node1555 = (inp[1]) ? node1561 : node1556;
										assign node1556 = (inp[13]) ? node1558 : 14'b00000111111111;
											assign node1558 = (inp[7]) ? 14'b00000011111111 : 14'b00000111111111;
										assign node1561 = (inp[7]) ? node1565 : node1562;
											assign node1562 = (inp[9]) ? 14'b00000111111111 : 14'b00000011111111;
											assign node1565 = (inp[13]) ? 14'b00000000111111 : 14'b00000001111111;
									assign node1568 = (inp[7]) ? node1574 : node1569;
										assign node1569 = (inp[2]) ? 14'b00000000011111 : node1570;
											assign node1570 = (inp[5]) ? 14'b00000011111111 : 14'b00000001111111;
										assign node1574 = (inp[1]) ? 14'b00000000011111 : 14'b00000000111111;
							assign node1577 = (inp[9]) ? node1589 : node1578;
								assign node1578 = (inp[10]) ? node1584 : node1579;
									assign node1579 = (inp[4]) ? 14'b00000011111111 : node1580;
										assign node1580 = (inp[5]) ? 14'b00000001111111 : 14'b00000011111111;
									assign node1584 = (inp[7]) ? 14'b00000000111111 : node1585;
										assign node1585 = (inp[4]) ? 14'b00000001111111 : 14'b00000011111111;
								assign node1589 = (inp[2]) ? node1603 : node1590;
									assign node1590 = (inp[4]) ? node1598 : node1591;
										assign node1591 = (inp[10]) ? node1595 : node1592;
											assign node1592 = (inp[1]) ? 14'b00000001111111 : 14'b00000011111111;
											assign node1595 = (inp[7]) ? 14'b00000001111111 : 14'b00000000111111;
										assign node1598 = (inp[7]) ? 14'b00000000111111 : node1599;
											assign node1599 = (inp[10]) ? 14'b00000001111111 : 14'b00000000111111;
									assign node1603 = (inp[13]) ? node1607 : node1604;
										assign node1604 = (inp[4]) ? 14'b00000001111111 : 14'b00000000111111;
										assign node1607 = (inp[5]) ? 14'b00000000001111 : 14'b00000000011111;
					assign node1610 = (inp[2]) ? node1694 : node1611;
						assign node1611 = (inp[1]) ? node1661 : node1612;
							assign node1612 = (inp[10]) ? node1640 : node1613;
								assign node1613 = (inp[7]) ? node1629 : node1614;
									assign node1614 = (inp[13]) ? node1622 : node1615;
										assign node1615 = (inp[4]) ? node1619 : node1616;
											assign node1616 = (inp[9]) ? 14'b00001111111111 : 14'b00011111111111;
											assign node1619 = (inp[5]) ? 14'b00000011111111 : 14'b00000111111111;
										assign node1622 = (inp[3]) ? node1624 : 14'b00000111111111;
											assign node1624 = (inp[9]) ? 14'b00000011111111 : node1625;
												assign node1625 = (inp[0]) ? 14'b00000111111111 : 14'b00000011111111;
									assign node1629 = (inp[3]) ? node1633 : node1630;
										assign node1630 = (inp[13]) ? 14'b00000011111111 : 14'b00000111111111;
										assign node1633 = (inp[4]) ? node1635 : 14'b00000011111111;
											assign node1635 = (inp[13]) ? 14'b00000001111111 : node1636;
												assign node1636 = (inp[0]) ? 14'b00000001111111 : 14'b00000011111111;
								assign node1640 = (inp[0]) ? node1656 : node1641;
									assign node1641 = (inp[5]) ? node1649 : node1642;
										assign node1642 = (inp[3]) ? node1644 : 14'b00001111111111;
											assign node1644 = (inp[4]) ? 14'b00000011111111 : node1645;
												assign node1645 = (inp[7]) ? 14'b00000011111111 : 14'b00000111111111;
										assign node1649 = (inp[7]) ? 14'b00000000111111 : node1650;
											assign node1650 = (inp[9]) ? node1652 : 14'b00000011111111;
												assign node1652 = (inp[3]) ? 14'b00000001111111 : 14'b00000011111111;
									assign node1656 = (inp[4]) ? node1658 : 14'b00000001111111;
										assign node1658 = (inp[3]) ? 14'b00000000111111 : 14'b00000011111111;
							assign node1661 = (inp[3]) ? node1679 : node1662;
								assign node1662 = (inp[9]) ? node1670 : node1663;
									assign node1663 = (inp[0]) ? node1665 : 14'b00000011111111;
										assign node1665 = (inp[10]) ? node1667 : 14'b00000011111111;
											assign node1667 = (inp[4]) ? 14'b00000001111111 : 14'b00000011111111;
									assign node1670 = (inp[0]) ? node1676 : node1671;
										assign node1671 = (inp[7]) ? 14'b00000001111111 : node1672;
											assign node1672 = (inp[10]) ? 14'b00000001111111 : 14'b00000011111111;
										assign node1676 = (inp[5]) ? 14'b00000000111111 : 14'b00000001111111;
								assign node1679 = (inp[0]) ? node1691 : node1680;
									assign node1680 = (inp[4]) ? node1686 : node1681;
										assign node1681 = (inp[5]) ? 14'b00000001111111 : node1682;
											assign node1682 = (inp[7]) ? 14'b00000011111111 : 14'b00000111111111;
										assign node1686 = (inp[9]) ? node1688 : 14'b00000000111111;
											assign node1688 = (inp[13]) ? 14'b00000000011111 : 14'b00000000111111;
									assign node1691 = (inp[10]) ? 14'b00000000011111 : 14'b00000000111111;
						assign node1694 = (inp[9]) ? node1726 : node1695;
							assign node1695 = (inp[13]) ? node1713 : node1696;
								assign node1696 = (inp[5]) ? node1706 : node1697;
									assign node1697 = (inp[7]) ? 14'b00000011111111 : node1698;
										assign node1698 = (inp[1]) ? 14'b00000111111111 : node1699;
											assign node1699 = (inp[3]) ? 14'b00000111111111 : node1700;
												assign node1700 = (inp[4]) ? 14'b00000111111111 : 14'b00001111111111;
									assign node1706 = (inp[4]) ? 14'b00000001111111 : node1707;
										assign node1707 = (inp[3]) ? node1709 : 14'b00000111111111;
											assign node1709 = (inp[0]) ? 14'b00000001111111 : 14'b00000011111111;
								assign node1713 = (inp[0]) ? node1717 : node1714;
									assign node1714 = (inp[10]) ? 14'b00000001111111 : 14'b00000011111111;
									assign node1717 = (inp[5]) ? 14'b00000000111111 : node1718;
										assign node1718 = (inp[1]) ? node1720 : 14'b00000001111111;
											assign node1720 = (inp[3]) ? node1722 : 14'b00000000111111;
												assign node1722 = (inp[7]) ? 14'b00000000011111 : 14'b00000000111111;
							assign node1726 = (inp[10]) ? node1746 : node1727;
								assign node1727 = (inp[4]) ? node1735 : node1728;
									assign node1728 = (inp[1]) ? 14'b00000001111111 : node1729;
										assign node1729 = (inp[7]) ? 14'b00000001111111 : node1730;
											assign node1730 = (inp[3]) ? 14'b00000001111111 : 14'b00000011111111;
									assign node1735 = (inp[0]) ? node1743 : node1736;
										assign node1736 = (inp[5]) ? 14'b00000011111111 : node1737;
											assign node1737 = (inp[7]) ? node1739 : 14'b00000001111111;
												assign node1739 = (inp[3]) ? 14'b00000000111111 : 14'b00000001111111;
										assign node1743 = (inp[3]) ? 14'b00000000011111 : 14'b00000000111111;
								assign node1746 = (inp[0]) ? node1756 : node1747;
									assign node1747 = (inp[3]) ? node1751 : node1748;
										assign node1748 = (inp[1]) ? 14'b00000000111111 : 14'b00000001111111;
										assign node1751 = (inp[13]) ? 14'b00000000011111 : node1752;
											assign node1752 = (inp[1]) ? 14'b00000000001111 : 14'b00000000111111;
									assign node1756 = (inp[1]) ? node1762 : node1757;
										assign node1757 = (inp[7]) ? node1759 : 14'b00000000011111;
											assign node1759 = (inp[4]) ? 14'b00000000001111 : 14'b00000000011111;
										assign node1762 = (inp[3]) ? 14'b00000000011111 : 14'b00000000001111;
				assign node1765 = (inp[2]) ? node1941 : node1766;
					assign node1766 = (inp[10]) ? node1858 : node1767;
						assign node1767 = (inp[4]) ? node1817 : node1768;
							assign node1768 = (inp[5]) ? node1790 : node1769;
								assign node1769 = (inp[0]) ? node1781 : node1770;
									assign node1770 = (inp[9]) ? 14'b00000111111111 : node1771;
										assign node1771 = (inp[12]) ? 14'b00000111111111 : node1772;
											assign node1772 = (inp[7]) ? 14'b00001111111111 : node1773;
												assign node1773 = (inp[1]) ? node1775 : 14'b00011111111111;
													assign node1775 = (inp[13]) ? 14'b00001111111111 : 14'b00011111111111;
									assign node1781 = (inp[1]) ? node1787 : node1782;
										assign node1782 = (inp[13]) ? node1784 : 14'b00001111111111;
											assign node1784 = (inp[3]) ? 14'b00000011111111 : 14'b00000111111111;
										assign node1787 = (inp[7]) ? 14'b00000001111111 : 14'b00000011111111;
								assign node1790 = (inp[7]) ? node1808 : node1791;
									assign node1791 = (inp[12]) ? node1799 : node1792;
										assign node1792 = (inp[13]) ? 14'b00000001111111 : node1793;
											assign node1793 = (inp[9]) ? 14'b00000111111111 : node1794;
												assign node1794 = (inp[0]) ? 14'b00000111111111 : 14'b00001111111111;
										assign node1799 = (inp[0]) ? node1805 : node1800;
											assign node1800 = (inp[1]) ? node1802 : 14'b00000011111111;
												assign node1802 = (inp[9]) ? 14'b00000011111111 : 14'b00000111111111;
											assign node1805 = (inp[9]) ? 14'b00000001111111 : 14'b00000011111111;
									assign node1808 = (inp[3]) ? node1814 : node1809;
										assign node1809 = (inp[12]) ? 14'b00000001111111 : node1810;
											assign node1810 = (inp[9]) ? 14'b00000001111111 : 14'b00000011111111;
										assign node1814 = (inp[0]) ? 14'b00000001111111 : 14'b00000000111111;
							assign node1817 = (inp[3]) ? node1831 : node1818;
								assign node1818 = (inp[1]) ? node1826 : node1819;
									assign node1819 = (inp[0]) ? node1823 : node1820;
										assign node1820 = (inp[9]) ? 14'b00000011111111 : 14'b00001111111111;
										assign node1823 = (inp[9]) ? 14'b00000001111111 : 14'b00000011111111;
									assign node1826 = (inp[13]) ? 14'b00000001111111 : node1827;
										assign node1827 = (inp[5]) ? 14'b00000001111111 : 14'b00000011111111;
								assign node1831 = (inp[13]) ? node1849 : node1832;
									assign node1832 = (inp[7]) ? node1840 : node1833;
										assign node1833 = (inp[5]) ? 14'b00000001111111 : node1834;
											assign node1834 = (inp[12]) ? node1836 : 14'b00000011111111;
												assign node1836 = (inp[9]) ? 14'b00000001111111 : 14'b00000011111111;
										assign node1840 = (inp[9]) ? node1842 : 14'b00000001111111;
											assign node1842 = (inp[12]) ? 14'b00000000111111 : node1843;
												assign node1843 = (inp[5]) ? node1845 : 14'b00000001111111;
													assign node1845 = (inp[1]) ? 14'b00000000111111 : 14'b00000001111111;
									assign node1849 = (inp[7]) ? node1855 : node1850;
										assign node1850 = (inp[9]) ? node1852 : 14'b00000001111111;
											assign node1852 = (inp[5]) ? 14'b00000000111111 : 14'b00000001111111;
										assign node1855 = (inp[9]) ? 14'b00000000001111 : 14'b00000000011111;
						assign node1858 = (inp[9]) ? node1900 : node1859;
							assign node1859 = (inp[0]) ? node1879 : node1860;
								assign node1860 = (inp[12]) ? node1874 : node1861;
									assign node1861 = (inp[7]) ? node1869 : node1862;
										assign node1862 = (inp[3]) ? node1866 : node1863;
											assign node1863 = (inp[4]) ? 14'b00000111111111 : 14'b00001111111111;
											assign node1866 = (inp[1]) ? 14'b00000011111111 : 14'b00000111111111;
										assign node1869 = (inp[3]) ? 14'b00000001111111 : node1870;
											assign node1870 = (inp[13]) ? 14'b00000111111111 : 14'b00000011111111;
									assign node1874 = (inp[3]) ? 14'b00000001111111 : node1875;
										assign node1875 = (inp[1]) ? 14'b00000001111111 : 14'b00000011111111;
								assign node1879 = (inp[3]) ? node1893 : node1880;
									assign node1880 = (inp[4]) ? node1890 : node1881;
										assign node1881 = (inp[1]) ? node1885 : node1882;
											assign node1882 = (inp[5]) ? 14'b00000011111111 : 14'b00000111111111;
											assign node1885 = (inp[13]) ? 14'b00000001111111 : node1886;
												assign node1886 = (inp[12]) ? 14'b00000011111111 : 14'b00000001111111;
										assign node1890 = (inp[12]) ? 14'b00000000111111 : 14'b00000001111111;
									assign node1893 = (inp[4]) ? node1895 : 14'b00000000111111;
										assign node1895 = (inp[7]) ? 14'b00000000001111 : node1896;
											assign node1896 = (inp[13]) ? 14'b00000000011111 : 14'b00000000111111;
							assign node1900 = (inp[13]) ? node1918 : node1901;
								assign node1901 = (inp[0]) ? node1909 : node1902;
									assign node1902 = (inp[5]) ? 14'b00000011111111 : node1903;
										assign node1903 = (inp[7]) ? node1905 : 14'b00000001111111;
											assign node1905 = (inp[3]) ? 14'b00000001111111 : 14'b00000000111111;
									assign node1909 = (inp[4]) ? node1913 : node1910;
										assign node1910 = (inp[7]) ? 14'b00000000111111 : 14'b00000001111111;
										assign node1913 = (inp[5]) ? node1915 : 14'b00000000111111;
											assign node1915 = (inp[3]) ? 14'b00000000011111 : 14'b00000000111111;
								assign node1918 = (inp[1]) ? node1928 : node1919;
									assign node1919 = (inp[5]) ? node1921 : 14'b00000001111111;
										assign node1921 = (inp[3]) ? node1923 : 14'b00000000111111;
											assign node1923 = (inp[0]) ? 14'b00000000011111 : node1924;
												assign node1924 = (inp[4]) ? 14'b00000000011111 : 14'b00000000111111;
									assign node1928 = (inp[3]) ? node1934 : node1929;
										assign node1929 = (inp[12]) ? node1931 : 14'b00000000011111;
											assign node1931 = (inp[7]) ? 14'b00000000001111 : 14'b00000000011111;
										assign node1934 = (inp[4]) ? node1936 : 14'b00000000000111;
											assign node1936 = (inp[12]) ? node1938 : 14'b00000000001111;
												assign node1938 = (inp[7]) ? 14'b00000000000111 : 14'b00000000001111;
					assign node1941 = (inp[13]) ? node2025 : node1942;
						assign node1942 = (inp[9]) ? node1988 : node1943;
							assign node1943 = (inp[0]) ? node1965 : node1944;
								assign node1944 = (inp[10]) ? node1952 : node1945;
									assign node1945 = (inp[12]) ? 14'b00000011111111 : node1946;
										assign node1946 = (inp[5]) ? 14'b00000011111111 : node1947;
											assign node1947 = (inp[1]) ? 14'b00000111111111 : 14'b00001111111111;
									assign node1952 = (inp[4]) ? node1960 : node1953;
										assign node1953 = (inp[12]) ? node1957 : node1954;
											assign node1954 = (inp[3]) ? 14'b00000011111111 : 14'b00000111111111;
											assign node1957 = (inp[3]) ? 14'b00000001111111 : 14'b00000011111111;
										assign node1960 = (inp[5]) ? node1962 : 14'b00000001111111;
											assign node1962 = (inp[3]) ? 14'b00000000111111 : 14'b00000001111111;
								assign node1965 = (inp[4]) ? node1977 : node1966;
									assign node1966 = (inp[1]) ? node1974 : node1967;
										assign node1967 = (inp[7]) ? node1969 : 14'b00000011111111;
											assign node1969 = (inp[5]) ? 14'b00000001111111 : node1970;
												assign node1970 = (inp[12]) ? 14'b00000001111111 : 14'b00000111111111;
										assign node1974 = (inp[7]) ? 14'b00000000111111 : 14'b00000001111111;
									assign node1977 = (inp[3]) ? node1983 : node1978;
										assign node1978 = (inp[12]) ? 14'b00000000111111 : node1979;
											assign node1979 = (inp[1]) ? 14'b00000000111111 : 14'b00000001111111;
										assign node1983 = (inp[7]) ? node1985 : 14'b00000000111111;
											assign node1985 = (inp[12]) ? 14'b00000000001111 : 14'b00000000011111;
							assign node1988 = (inp[5]) ? node2010 : node1989;
								assign node1989 = (inp[10]) ? node1999 : node1990;
									assign node1990 = (inp[0]) ? node1996 : node1991;
										assign node1991 = (inp[12]) ? 14'b00000001111111 : node1992;
											assign node1992 = (inp[3]) ? 14'b00000001111111 : 14'b00000011111111;
										assign node1996 = (inp[7]) ? 14'b00000000011111 : 14'b00000001111111;
									assign node1999 = (inp[1]) ? node2005 : node2000;
										assign node2000 = (inp[12]) ? node2002 : 14'b00000001111111;
											assign node2002 = (inp[0]) ? 14'b00000000111111 : 14'b00000001111111;
										assign node2005 = (inp[4]) ? 14'b00000000011111 : node2006;
											assign node2006 = (inp[0]) ? 14'b00000000011111 : 14'b00000001111111;
								assign node2010 = (inp[1]) ? node2016 : node2011;
									assign node2011 = (inp[0]) ? 14'b00000000011111 : node2012;
										assign node2012 = (inp[3]) ? 14'b00000000111111 : 14'b00000001111111;
									assign node2016 = (inp[10]) ? node2020 : node2017;
										assign node2017 = (inp[0]) ? 14'b00000000011111 : 14'b00000000111111;
										assign node2020 = (inp[4]) ? 14'b00000000001111 : node2021;
											assign node2021 = (inp[0]) ? 14'b00000000001111 : 14'b00000000011111;
						assign node2025 = (inp[10]) ? node2083 : node2026;
							assign node2026 = (inp[0]) ? node2056 : node2027;
								assign node2027 = (inp[9]) ? node2045 : node2028;
									assign node2028 = (inp[7]) ? node2038 : node2029;
										assign node2029 = (inp[12]) ? 14'b00000001111111 : node2030;
											assign node2030 = (inp[5]) ? node2032 : 14'b00000011111111;
												assign node2032 = (inp[3]) ? 14'b00000001111111 : node2033;
													assign node2033 = (inp[4]) ? 14'b00000001111111 : 14'b00000011111111;
										assign node2038 = (inp[3]) ? node2040 : 14'b00000001111111;
											assign node2040 = (inp[5]) ? 14'b00000000111111 : node2041;
												assign node2041 = (inp[4]) ? 14'b00000001111111 : 14'b00000000111111;
									assign node2045 = (inp[5]) ? node2053 : node2046;
										assign node2046 = (inp[12]) ? 14'b00000000111111 : node2047;
											assign node2047 = (inp[4]) ? node2049 : 14'b00000011111111;
												assign node2049 = (inp[3]) ? 14'b00000000111111 : 14'b00000001111111;
										assign node2053 = (inp[12]) ? 14'b00000000011111 : 14'b00000000111111;
								assign node2056 = (inp[1]) ? node2072 : node2057;
									assign node2057 = (inp[9]) ? node2065 : node2058;
										assign node2058 = (inp[7]) ? node2060 : 14'b00000001111111;
											assign node2060 = (inp[5]) ? 14'b00000000111111 : node2061;
												assign node2061 = (inp[4]) ? 14'b00000000111111 : 14'b00000001111111;
										assign node2065 = (inp[7]) ? 14'b00000000000111 : node2066;
											assign node2066 = (inp[3]) ? node2068 : 14'b00000000111111;
												assign node2068 = (inp[5]) ? 14'b00000000001111 : 14'b00000000111111;
									assign node2072 = (inp[12]) ? node2076 : node2073;
										assign node2073 = (inp[5]) ? 14'b00000000011111 : 14'b00000000111111;
										assign node2076 = (inp[7]) ? node2080 : node2077;
											assign node2077 = (inp[3]) ? 14'b00000000001111 : 14'b00000000011111;
											assign node2080 = (inp[9]) ? 14'b00000000001111 : 14'b00000000000111;
							assign node2083 = (inp[4]) ? node2113 : node2084;
								assign node2084 = (inp[1]) ? node2100 : node2085;
									assign node2085 = (inp[3]) ? node2093 : node2086;
										assign node2086 = (inp[0]) ? 14'b00000000111111 : node2087;
											assign node2087 = (inp[5]) ? 14'b00000001111111 : node2088;
												assign node2088 = (inp[9]) ? 14'b00000001111111 : 14'b00000011111111;
										assign node2093 = (inp[0]) ? 14'b00000001111111 : node2094;
											assign node2094 = (inp[9]) ? node2096 : 14'b00000000111111;
												assign node2096 = (inp[7]) ? 14'b00000000001111 : 14'b00000000111111;
									assign node2100 = (inp[0]) ? node2110 : node2101;
										assign node2101 = (inp[9]) ? node2105 : node2102;
											assign node2102 = (inp[7]) ? 14'b00000000011111 : 14'b00000000111111;
											assign node2105 = (inp[5]) ? 14'b00000000011111 : node2106;
												assign node2106 = (inp[12]) ? 14'b00000000001111 : 14'b00000000011111;
										assign node2110 = (inp[5]) ? 14'b00000000000011 : 14'b00000000011111;
								assign node2113 = (inp[1]) ? node2127 : node2114;
									assign node2114 = (inp[7]) ? node2120 : node2115;
										assign node2115 = (inp[9]) ? node2117 : 14'b00000000011111;
											assign node2117 = (inp[12]) ? 14'b00000000011111 : 14'b00000000111111;
										assign node2120 = (inp[12]) ? 14'b00000000000111 : node2121;
											assign node2121 = (inp[5]) ? node2123 : 14'b00000000011111;
												assign node2123 = (inp[0]) ? 14'b00000000011111 : 14'b00000000001111;
									assign node2127 = (inp[0]) ? node2131 : node2128;
										assign node2128 = (inp[3]) ? 14'b00000000001111 : 14'b00000000011111;
										assign node2131 = (inp[3]) ? node2133 : 14'b00000000001111;
											assign node2133 = (inp[12]) ? 14'b00000000000111 : node2134;
												assign node2134 = (inp[9]) ? 14'b00000000000111 : 14'b00000000001111;
			assign node2138 = (inp[9]) ? node2490 : node2139;
				assign node2139 = (inp[13]) ? node2311 : node2140;
					assign node2140 = (inp[0]) ? node2222 : node2141;
						assign node2141 = (inp[5]) ? node2183 : node2142;
							assign node2142 = (inp[2]) ? node2162 : node2143;
								assign node2143 = (inp[7]) ? node2151 : node2144;
									assign node2144 = (inp[3]) ? node2148 : node2145;
										assign node2145 = (inp[10]) ? 14'b00001111111111 : 14'b00011111111111;
										assign node2148 = (inp[10]) ? 14'b00000011111111 : 14'b00000111111111;
									assign node2151 = (inp[10]) ? node2159 : node2152;
										assign node2152 = (inp[6]) ? node2154 : 14'b00000111111111;
											assign node2154 = (inp[1]) ? 14'b00000011111111 : node2155;
												assign node2155 = (inp[12]) ? 14'b00000011111111 : 14'b00000111111111;
										assign node2159 = (inp[3]) ? 14'b00000001111111 : 14'b00000011111111;
								assign node2162 = (inp[12]) ? node2168 : node2163;
									assign node2163 = (inp[4]) ? 14'b00000011111111 : node2164;
										assign node2164 = (inp[10]) ? 14'b00000011111111 : 14'b00000111111111;
									assign node2168 = (inp[6]) ? node2180 : node2169;
										assign node2169 = (inp[3]) ? node2175 : node2170;
											assign node2170 = (inp[7]) ? 14'b00000011111111 : node2171;
												assign node2171 = (inp[4]) ? 14'b00000011111111 : 14'b00000111111111;
											assign node2175 = (inp[10]) ? node2177 : 14'b00000011111111;
												assign node2177 = (inp[4]) ? 14'b00000000111111 : 14'b00000001111111;
										assign node2180 = (inp[10]) ? 14'b00000000111111 : 14'b00000001111111;
							assign node2183 = (inp[3]) ? node2205 : node2184;
								assign node2184 = (inp[4]) ? node2196 : node2185;
									assign node2185 = (inp[10]) ? node2189 : node2186;
										assign node2186 = (inp[6]) ? 14'b00000011111111 : 14'b00000111111111;
										assign node2189 = (inp[1]) ? 14'b00000001111111 : node2190;
											assign node2190 = (inp[2]) ? node2192 : 14'b00000011111111;
												assign node2192 = (inp[7]) ? 14'b00000001111111 : 14'b00000011111111;
									assign node2196 = (inp[1]) ? 14'b00000000111111 : node2197;
										assign node2197 = (inp[6]) ? node2199 : 14'b00000011111111;
											assign node2199 = (inp[2]) ? 14'b00000001111111 : node2200;
												assign node2200 = (inp[7]) ? 14'b00000001111111 : 14'b00000011111111;
								assign node2205 = (inp[10]) ? node2209 : node2206;
									assign node2206 = (inp[1]) ? 14'b00000001111111 : 14'b00000011111111;
									assign node2209 = (inp[6]) ? node2217 : node2210;
										assign node2210 = (inp[7]) ? node2214 : node2211;
											assign node2211 = (inp[2]) ? 14'b00000011111111 : 14'b00000001111111;
											assign node2214 = (inp[1]) ? 14'b00000001111111 : 14'b00000000111111;
										assign node2217 = (inp[1]) ? node2219 : 14'b00000000111111;
											assign node2219 = (inp[7]) ? 14'b00000000001111 : 14'b00000000011111;
						assign node2222 = (inp[6]) ? node2280 : node2223;
							assign node2223 = (inp[12]) ? node2245 : node2224;
								assign node2224 = (inp[3]) ? node2236 : node2225;
									assign node2225 = (inp[2]) ? node2231 : node2226;
										assign node2226 = (inp[4]) ? 14'b00000011111111 : node2227;
											assign node2227 = (inp[10]) ? 14'b00000111111111 : 14'b00001111111111;
										assign node2231 = (inp[4]) ? 14'b00000011111111 : node2232;
											assign node2232 = (inp[7]) ? 14'b00000001111111 : 14'b00000011111111;
									assign node2236 = (inp[7]) ? 14'b00000000111111 : node2237;
										assign node2237 = (inp[4]) ? 14'b00000001111111 : node2238;
											assign node2238 = (inp[1]) ? node2240 : 14'b00000111111111;
												assign node2240 = (inp[10]) ? 14'b00000001111111 : 14'b00000011111111;
								assign node2245 = (inp[2]) ? node2259 : node2246;
									assign node2246 = (inp[3]) ? node2256 : node2247;
										assign node2247 = (inp[7]) ? node2249 : 14'b00000011111111;
											assign node2249 = (inp[1]) ? 14'b00000001111111 : node2250;
												assign node2250 = (inp[5]) ? 14'b00000001111111 : node2251;
													assign node2251 = (inp[10]) ? 14'b00000001111111 : 14'b00000011111111;
										assign node2256 = (inp[4]) ? 14'b00000001111111 : 14'b00000000111111;
									assign node2259 = (inp[1]) ? node2271 : node2260;
										assign node2260 = (inp[4]) ? node2264 : node2261;
											assign node2261 = (inp[10]) ? 14'b00000011111111 : 14'b00000001111111;
											assign node2264 = (inp[5]) ? 14'b00000000111111 : node2265;
												assign node2265 = (inp[10]) ? node2267 : 14'b00000001111111;
													assign node2267 = (inp[3]) ? 14'b00000000111111 : 14'b00000001111111;
										assign node2271 = (inp[5]) ? node2277 : node2272;
											assign node2272 = (inp[10]) ? 14'b00000000111111 : node2273;
												assign node2273 = (inp[7]) ? 14'b00000000111111 : 14'b00000001111111;
											assign node2277 = (inp[7]) ? 14'b00000000011111 : 14'b00000000111111;
							assign node2280 = (inp[12]) ? node2296 : node2281;
								assign node2281 = (inp[10]) ? node2287 : node2282;
									assign node2282 = (inp[7]) ? node2284 : 14'b00000011111111;
										assign node2284 = (inp[5]) ? 14'b00000000111111 : 14'b00000001111111;
									assign node2287 = (inp[5]) ? node2291 : node2288;
										assign node2288 = (inp[7]) ? 14'b00000001111111 : 14'b00000000111111;
										assign node2291 = (inp[1]) ? node2293 : 14'b00000000111111;
											assign node2293 = (inp[4]) ? 14'b00000000011111 : 14'b00000000111111;
								assign node2296 = (inp[2]) ? node2304 : node2297;
									assign node2297 = (inp[4]) ? node2301 : node2298;
										assign node2298 = (inp[5]) ? 14'b00000000111111 : 14'b00000001111111;
										assign node2301 = (inp[1]) ? 14'b00000000011111 : 14'b00000000111111;
									assign node2304 = (inp[7]) ? node2308 : node2305;
										assign node2305 = (inp[4]) ? 14'b00000000011111 : 14'b00000000111111;
										assign node2308 = (inp[3]) ? 14'b00000000001111 : 14'b00000000011111;
					assign node2311 = (inp[0]) ? node2409 : node2312;
						assign node2312 = (inp[4]) ? node2360 : node2313;
							assign node2313 = (inp[1]) ? node2339 : node2314;
								assign node2314 = (inp[2]) ? node2326 : node2315;
									assign node2315 = (inp[3]) ? node2321 : node2316;
										assign node2316 = (inp[7]) ? 14'b00000011111111 : node2317;
											assign node2317 = (inp[6]) ? 14'b00000111111111 : 14'b00001111111111;
										assign node2321 = (inp[5]) ? 14'b00000001111111 : node2322;
											assign node2322 = (inp[10]) ? 14'b00000001111111 : 14'b00000011111111;
									assign node2326 = (inp[6]) ? node2334 : node2327;
										assign node2327 = (inp[7]) ? node2329 : 14'b00000011111111;
											assign node2329 = (inp[3]) ? 14'b00000001111111 : node2330;
												assign node2330 = (inp[12]) ? 14'b00000001111111 : 14'b00000011111111;
										assign node2334 = (inp[3]) ? 14'b00000000111111 : node2335;
											assign node2335 = (inp[7]) ? 14'b00000001111111 : 14'b00000000111111;
								assign node2339 = (inp[3]) ? node2353 : node2340;
									assign node2340 = (inp[6]) ? node2348 : node2341;
										assign node2341 = (inp[5]) ? node2343 : 14'b00000011111111;
											assign node2343 = (inp[10]) ? 14'b00000001111111 : node2344;
												assign node2344 = (inp[12]) ? 14'b00000001111111 : 14'b00000011111111;
										assign node2348 = (inp[12]) ? node2350 : 14'b00000011111111;
											assign node2350 = (inp[7]) ? 14'b00000000011111 : 14'b00000000111111;
									assign node2353 = (inp[2]) ? node2357 : node2354;
										assign node2354 = (inp[10]) ? 14'b00000000111111 : 14'b00000001111111;
										assign node2357 = (inp[7]) ? 14'b00000000011111 : 14'b00000000111111;
							assign node2360 = (inp[12]) ? node2382 : node2361;
								assign node2361 = (inp[6]) ? node2373 : node2362;
									assign node2362 = (inp[7]) ? node2370 : node2363;
										assign node2363 = (inp[5]) ? 14'b00000001111111 : node2364;
											assign node2364 = (inp[10]) ? node2366 : 14'b00000011111111;
												assign node2366 = (inp[1]) ? 14'b00000001111111 : 14'b00000011111111;
										assign node2370 = (inp[1]) ? 14'b00000000111111 : 14'b00000001111111;
									assign node2373 = (inp[2]) ? node2379 : node2374;
										assign node2374 = (inp[7]) ? node2376 : 14'b00000000111111;
											assign node2376 = (inp[5]) ? 14'b00000001111111 : 14'b00000011111111;
										assign node2379 = (inp[7]) ? 14'b00000000011111 : 14'b00000000111111;
								assign node2382 = (inp[3]) ? node2398 : node2383;
									assign node2383 = (inp[7]) ? node2389 : node2384;
										assign node2384 = (inp[5]) ? 14'b00000000111111 : node2385;
											assign node2385 = (inp[2]) ? 14'b00000000111111 : 14'b00000011111111;
										assign node2389 = (inp[1]) ? node2395 : node2390;
											assign node2390 = (inp[5]) ? node2392 : 14'b00000000111111;
												assign node2392 = (inp[2]) ? 14'b00000000011111 : 14'b00000000111111;
											assign node2395 = (inp[5]) ? 14'b00000000000111 : 14'b00000000011111;
									assign node2398 = (inp[6]) ? node2406 : node2399;
										assign node2399 = (inp[7]) ? node2401 : 14'b00000000111111;
											assign node2401 = (inp[5]) ? node2403 : 14'b00000000011111;
												assign node2403 = (inp[1]) ? 14'b00000000001111 : 14'b00000000011111;
										assign node2406 = (inp[5]) ? 14'b00000000000011 : 14'b00000000001111;
						assign node2409 = (inp[3]) ? node2449 : node2410;
							assign node2410 = (inp[4]) ? node2432 : node2411;
								assign node2411 = (inp[10]) ? node2421 : node2412;
									assign node2412 = (inp[1]) ? node2416 : node2413;
										assign node2413 = (inp[7]) ? 14'b00000001111111 : 14'b00000111111111;
										assign node2416 = (inp[12]) ? node2418 : 14'b00000001111111;
											assign node2418 = (inp[7]) ? 14'b00000000011111 : 14'b00000000111111;
									assign node2421 = (inp[6]) ? node2423 : 14'b00000000111111;
										assign node2423 = (inp[12]) ? node2425 : 14'b00000000111111;
											assign node2425 = (inp[7]) ? 14'b00000000011111 : node2426;
												assign node2426 = (inp[5]) ? node2428 : 14'b00000000111111;
													assign node2428 = (inp[2]) ? 14'b00000000011111 : 14'b00000000111111;
								assign node2432 = (inp[2]) ? node2440 : node2433;
									assign node2433 = (inp[6]) ? node2435 : 14'b00000000111111;
										assign node2435 = (inp[12]) ? 14'b00000000011111 : node2436;
											assign node2436 = (inp[7]) ? 14'b00000000011111 : 14'b00000000111111;
									assign node2440 = (inp[5]) ? node2444 : node2441;
										assign node2441 = (inp[12]) ? 14'b00000000011111 : 14'b00000000111111;
										assign node2444 = (inp[7]) ? 14'b00000000001111 : node2445;
											assign node2445 = (inp[12]) ? 14'b00000000001111 : 14'b00000000011111;
							assign node2449 = (inp[10]) ? node2467 : node2450;
								assign node2450 = (inp[12]) ? node2458 : node2451;
									assign node2451 = (inp[4]) ? node2453 : 14'b00000001111111;
										assign node2453 = (inp[7]) ? node2455 : 14'b00000000111111;
											assign node2455 = (inp[1]) ? 14'b00000000011111 : 14'b00000000111111;
									assign node2458 = (inp[2]) ? node2460 : 14'b00000001111111;
										assign node2460 = (inp[5]) ? node2462 : 14'b00000000011111;
											assign node2462 = (inp[1]) ? 14'b00000000000111 : node2463;
												assign node2463 = (inp[6]) ? 14'b00000000011111 : 14'b00000000001111;
								assign node2467 = (inp[1]) ? node2477 : node2468;
									assign node2468 = (inp[4]) ? node2472 : node2469;
										assign node2469 = (inp[12]) ? 14'b00000000011111 : 14'b00000000111111;
										assign node2472 = (inp[12]) ? node2474 : 14'b00000000011111;
											assign node2474 = (inp[6]) ? 14'b00000000001111 : 14'b00000000011111;
									assign node2477 = (inp[2]) ? node2483 : node2478;
										assign node2478 = (inp[4]) ? 14'b00000000001111 : node2479;
											assign node2479 = (inp[5]) ? 14'b00000000111111 : 14'b00000000011111;
										assign node2483 = (inp[5]) ? 14'b00000000000111 : node2484;
											assign node2484 = (inp[6]) ? 14'b00000000001111 : node2485;
												assign node2485 = (inp[12]) ? 14'b00000000001111 : 14'b00000000011111;
				assign node2490 = (inp[3]) ? node2690 : node2491;
					assign node2491 = (inp[1]) ? node2587 : node2492;
						assign node2492 = (inp[7]) ? node2540 : node2493;
							assign node2493 = (inp[4]) ? node2515 : node2494;
								assign node2494 = (inp[6]) ? node2508 : node2495;
									assign node2495 = (inp[0]) ? node2501 : node2496;
										assign node2496 = (inp[13]) ? 14'b00000011111111 : node2497;
											assign node2497 = (inp[2]) ? 14'b00000111111111 : 14'b00001111111111;
										assign node2501 = (inp[2]) ? 14'b00000001111111 : node2502;
											assign node2502 = (inp[5]) ? node2504 : 14'b00000011111111;
												assign node2504 = (inp[12]) ? 14'b00000001111111 : 14'b00000011111111;
									assign node2508 = (inp[0]) ? node2510 : 14'b00000001111111;
										assign node2510 = (inp[2]) ? 14'b00000001111111 : node2511;
											assign node2511 = (inp[10]) ? 14'b00000001111111 : 14'b00000011111111;
								assign node2515 = (inp[10]) ? node2531 : node2516;
									assign node2516 = (inp[5]) ? node2526 : node2517;
										assign node2517 = (inp[13]) ? node2521 : node2518;
											assign node2518 = (inp[6]) ? 14'b00000011111111 : 14'b00001111111111;
											assign node2521 = (inp[6]) ? node2523 : 14'b00000001111111;
												assign node2523 = (inp[12]) ? 14'b00000001111111 : 14'b00000011111111;
										assign node2526 = (inp[13]) ? node2528 : 14'b00000001111111;
											assign node2528 = (inp[12]) ? 14'b00000001111111 : 14'b00000000111111;
									assign node2531 = (inp[2]) ? node2535 : node2532;
										assign node2532 = (inp[5]) ? 14'b00000000111111 : 14'b00000001111111;
										assign node2535 = (inp[0]) ? 14'b00000000011111 : node2536;
											assign node2536 = (inp[12]) ? 14'b00000000011111 : 14'b00000001111111;
							assign node2540 = (inp[6]) ? node2560 : node2541;
								assign node2541 = (inp[12]) ? node2553 : node2542;
									assign node2542 = (inp[0]) ? node2550 : node2543;
										assign node2543 = (inp[13]) ? node2545 : 14'b00000011111111;
											assign node2545 = (inp[10]) ? 14'b00000001111111 : node2546;
												assign node2546 = (inp[2]) ? 14'b00000001111111 : 14'b00000011111111;
										assign node2550 = (inp[10]) ? 14'b00000000111111 : 14'b00000001111111;
									assign node2553 = (inp[10]) ? node2557 : node2554;
										assign node2554 = (inp[4]) ? 14'b00000000111111 : 14'b00000001111111;
										assign node2557 = (inp[0]) ? 14'b00000000011111 : 14'b00000000111111;
								assign node2560 = (inp[4]) ? node2568 : node2561;
									assign node2561 = (inp[5]) ? node2563 : 14'b00000001111111;
										assign node2563 = (inp[13]) ? 14'b00000000011111 : node2564;
											assign node2564 = (inp[2]) ? 14'b00000000011111 : 14'b00000001111111;
									assign node2568 = (inp[5]) ? node2580 : node2569;
										assign node2569 = (inp[12]) ? node2577 : node2570;
											assign node2570 = (inp[0]) ? node2574 : node2571;
												assign node2571 = (inp[2]) ? 14'b00000001111111 : 14'b00000000111111;
												assign node2574 = (inp[10]) ? 14'b00000000011111 : 14'b00000000111111;
											assign node2577 = (inp[0]) ? 14'b00000000001111 : 14'b00000000011111;
										assign node2580 = (inp[0]) ? node2584 : node2581;
											assign node2581 = (inp[2]) ? 14'b00000000001111 : 14'b00000000011111;
											assign node2584 = (inp[12]) ? 14'b00000000000011 : 14'b00000000000111;
						assign node2587 = (inp[2]) ? node2643 : node2588;
							assign node2588 = (inp[5]) ? node2612 : node2589;
								assign node2589 = (inp[7]) ? node2599 : node2590;
									assign node2590 = (inp[13]) ? node2592 : 14'b00000111111111;
										assign node2592 = (inp[10]) ? node2594 : 14'b00000001111111;
											assign node2594 = (inp[4]) ? 14'b00000000111111 : node2595;
												assign node2595 = (inp[0]) ? 14'b00000000111111 : 14'b00000001111111;
									assign node2599 = (inp[4]) ? node2607 : node2600;
										assign node2600 = (inp[0]) ? node2602 : 14'b00000001111111;
											assign node2602 = (inp[10]) ? node2604 : 14'b00000000111111;
												assign node2604 = (inp[12]) ? 14'b00000000011111 : 14'b00000000111111;
										assign node2607 = (inp[0]) ? 14'b00000000011111 : node2608;
											assign node2608 = (inp[13]) ? 14'b00000000011111 : 14'b00000000111111;
								assign node2612 = (inp[6]) ? node2632 : node2613;
									assign node2613 = (inp[10]) ? node2617 : node2614;
										assign node2614 = (inp[12]) ? 14'b00000000111111 : 14'b00000001111111;
										assign node2617 = (inp[12]) ? node2619 : 14'b00000000111111;
											assign node2619 = (inp[7]) ? 14'b00000000001111 : node2620;
												assign node2620 = (inp[4]) ? node2626 : node2621;
													assign node2621 = (inp[13]) ? node2623 : 14'b00000000111111;
														assign node2623 = (inp[0]) ? 14'b00000000011111 : 14'b00000000111111;
													assign node2626 = (inp[0]) ? 14'b00000000011111 : node2627;
														assign node2627 = (inp[13]) ? 14'b00000000011111 : 14'b00000000111111;
									assign node2632 = (inp[10]) ? node2636 : node2633;
										assign node2633 = (inp[12]) ? 14'b00000000011111 : 14'b00000000111111;
										assign node2636 = (inp[0]) ? node2638 : 14'b00000000011111;
											assign node2638 = (inp[7]) ? 14'b00000000001111 : node2639;
												assign node2639 = (inp[4]) ? 14'b00000000001111 : 14'b00000000011111;
							assign node2643 = (inp[10]) ? node2667 : node2644;
								assign node2644 = (inp[7]) ? node2656 : node2645;
									assign node2645 = (inp[5]) ? node2649 : node2646;
										assign node2646 = (inp[13]) ? 14'b00000001111111 : 14'b00000000111111;
										assign node2649 = (inp[6]) ? node2651 : 14'b00000000111111;
											assign node2651 = (inp[0]) ? 14'b00000000001111 : node2652;
												assign node2652 = (inp[4]) ? 14'b00000000011111 : 14'b00000000111111;
									assign node2656 = (inp[6]) ? 14'b00000000001111 : node2657;
										assign node2657 = (inp[4]) ? node2663 : node2658;
											assign node2658 = (inp[13]) ? node2660 : 14'b00000001111111;
												assign node2660 = (inp[5]) ? 14'b00000000011111 : 14'b00000000111111;
											assign node2663 = (inp[13]) ? 14'b00000000001111 : 14'b00000000011111;
								assign node2667 = (inp[12]) ? node2679 : node2668;
									assign node2668 = (inp[5]) ? node2674 : node2669;
										assign node2669 = (inp[6]) ? 14'b00000000011111 : node2670;
											assign node2670 = (inp[7]) ? 14'b00000000111111 : 14'b00000001111111;
										assign node2674 = (inp[13]) ? 14'b00000000000111 : node2675;
											assign node2675 = (inp[4]) ? 14'b00000000001111 : 14'b00000000011111;
									assign node2679 = (inp[7]) ? node2687 : node2680;
										assign node2680 = (inp[0]) ? node2682 : 14'b00000000001111;
											assign node2682 = (inp[4]) ? node2684 : 14'b00000000001111;
												assign node2684 = (inp[6]) ? 14'b00000000000011 : 14'b00000000001111;
										assign node2687 = (inp[0]) ? 14'b00000000000011 : 14'b00000000000111;
					assign node2690 = (inp[2]) ? node2782 : node2691;
						assign node2691 = (inp[6]) ? node2727 : node2692;
							assign node2692 = (inp[5]) ? node2720 : node2693;
								assign node2693 = (inp[12]) ? node2707 : node2694;
									assign node2694 = (inp[0]) ? node2702 : node2695;
										assign node2695 = (inp[7]) ? node2697 : 14'b00000011111111;
											assign node2697 = (inp[4]) ? 14'b00000001111111 : node2698;
												assign node2698 = (inp[13]) ? 14'b00000001111111 : 14'b00000011111111;
										assign node2702 = (inp[13]) ? 14'b00000000111111 : node2703;
											assign node2703 = (inp[1]) ? 14'b00000000111111 : 14'b00000001111111;
									assign node2707 = (inp[10]) ? node2715 : node2708;
										assign node2708 = (inp[13]) ? 14'b00000000011111 : node2709;
											assign node2709 = (inp[0]) ? 14'b00000000111111 : node2710;
												assign node2710 = (inp[7]) ? 14'b00000001111111 : 14'b00000011111111;
										assign node2715 = (inp[0]) ? 14'b00000000000111 : node2716;
											assign node2716 = (inp[1]) ? 14'b00000000011111 : 14'b00000000111111;
								assign node2720 = (inp[7]) ? 14'b00000000011111 : node2721;
									assign node2721 = (inp[13]) ? node2723 : 14'b00000000111111;
										assign node2723 = (inp[1]) ? 14'b00000000011111 : 14'b00000000111111;
							assign node2727 = (inp[10]) ? node2755 : node2728;
								assign node2728 = (inp[13]) ? node2742 : node2729;
									assign node2729 = (inp[12]) ? node2733 : node2730;
										assign node2730 = (inp[5]) ? 14'b00000000111111 : 14'b00000111111111;
										assign node2733 = (inp[4]) ? node2739 : node2734;
											assign node2734 = (inp[7]) ? 14'b00000000111111 : node2735;
												assign node2735 = (inp[5]) ? 14'b00000000111111 : 14'b00000001111111;
											assign node2739 = (inp[0]) ? 14'b00000000111111 : 14'b00000000011111;
									assign node2742 = (inp[4]) ? node2750 : node2743;
										assign node2743 = (inp[7]) ? 14'b00000000001111 : node2744;
											assign node2744 = (inp[0]) ? node2746 : 14'b00000000111111;
												assign node2746 = (inp[12]) ? 14'b00000000011111 : 14'b00000000111111;
										assign node2750 = (inp[0]) ? node2752 : 14'b00000000011111;
											assign node2752 = (inp[5]) ? 14'b00000000000111 : 14'b00000000011111;
								assign node2755 = (inp[1]) ? node2767 : node2756;
									assign node2756 = (inp[12]) ? node2760 : node2757;
										assign node2757 = (inp[13]) ? 14'b00000000011111 : 14'b00000000111111;
										assign node2760 = (inp[4]) ? node2762 : 14'b00000000011111;
											assign node2762 = (inp[5]) ? node2764 : 14'b00000000011111;
												assign node2764 = (inp[7]) ? 14'b00000000001111 : 14'b00000000011111;
									assign node2767 = (inp[4]) ? node2769 : 14'b00000000011111;
										assign node2769 = (inp[0]) ? node2773 : node2770;
											assign node2770 = (inp[12]) ? 14'b00000000000111 : 14'b00000000001111;
											assign node2773 = (inp[13]) ? node2775 : 14'b00000000001111;
												assign node2775 = (inp[5]) ? 14'b00000000000011 : node2776;
													assign node2776 = (inp[12]) ? node2778 : 14'b00000000000111;
														assign node2778 = (inp[7]) ? 14'b00000000000011 : 14'b00000000000111;
						assign node2782 = (inp[13]) ? node2820 : node2783;
							assign node2783 = (inp[1]) ? node2805 : node2784;
								assign node2784 = (inp[7]) ? node2790 : node2785;
									assign node2785 = (inp[10]) ? 14'b00000000111111 : node2786;
										assign node2786 = (inp[6]) ? 14'b00000000011111 : 14'b00000001111111;
									assign node2790 = (inp[4]) ? node2794 : node2791;
										assign node2791 = (inp[10]) ? 14'b00000000111111 : 14'b00000000011111;
										assign node2794 = (inp[0]) ? node2800 : node2795;
											assign node2795 = (inp[5]) ? node2797 : 14'b00000000011111;
												assign node2797 = (inp[6]) ? 14'b00000000001111 : 14'b00000000011111;
											assign node2800 = (inp[10]) ? 14'b00000000001111 : node2801;
												assign node2801 = (inp[6]) ? 14'b00000000001111 : 14'b00000000011111;
								assign node2805 = (inp[4]) ? node2813 : node2806;
									assign node2806 = (inp[6]) ? 14'b00000000001111 : node2807;
										assign node2807 = (inp[7]) ? node2809 : 14'b00000000111111;
											assign node2809 = (inp[0]) ? 14'b00000000001111 : 14'b00000000011111;
									assign node2813 = (inp[10]) ? node2817 : node2814;
										assign node2814 = (inp[0]) ? 14'b00000000001111 : 14'b00000000011111;
										assign node2817 = (inp[7]) ? 14'b00000000000001 : 14'b00000000001111;
							assign node2820 = (inp[4]) ? node2840 : node2821;
								assign node2821 = (inp[10]) ? node2823 : 14'b00000000011111;
									assign node2823 = (inp[0]) ? node2831 : node2824;
										assign node2824 = (inp[5]) ? 14'b00000000001111 : node2825;
											assign node2825 = (inp[12]) ? 14'b00000000011111 : node2826;
												assign node2826 = (inp[1]) ? 14'b00000000011111 : 14'b00000000111111;
										assign node2831 = (inp[1]) ? node2833 : 14'b00000000001111;
											assign node2833 = (inp[7]) ? 14'b00000000000111 : node2834;
												assign node2834 = (inp[5]) ? node2836 : 14'b00000000001111;
													assign node2836 = (inp[6]) ? 14'b00000000000111 : 14'b00000000001111;
								assign node2840 = (inp[10]) ? node2852 : node2841;
									assign node2841 = (inp[0]) ? node2847 : node2842;
										assign node2842 = (inp[12]) ? node2844 : 14'b00000000011111;
											assign node2844 = (inp[5]) ? 14'b00000000001111 : 14'b00000000011111;
										assign node2847 = (inp[5]) ? node2849 : 14'b00000000001111;
											assign node2849 = (inp[6]) ? 14'b00000000000111 : 14'b00000000001111;
									assign node2852 = (inp[5]) ? node2858 : node2853;
										assign node2853 = (inp[12]) ? 14'b00000000000111 : node2854;
											assign node2854 = (inp[6]) ? 14'b00000000000111 : 14'b00000000001111;
										assign node2858 = (inp[7]) ? 14'b00000000000111 : node2859;
											assign node2859 = (inp[1]) ? node2861 : 14'b00000000000011;
												assign node2861 = (inp[0]) ? 14'b00000000000001 : 14'b00000000000011;

endmodule