module dtc_split33_bm47 (
	input  wire [16-1:0] inp,
	output wire [1-1:0] outp
);

	wire [1-1:0] node1;
	wire [1-1:0] node2;
	wire [1-1:0] node3;
	wire [1-1:0] node4;
	wire [1-1:0] node5;
	wire [1-1:0] node6;
	wire [1-1:0] node8;
	wire [1-1:0] node9;
	wire [1-1:0] node11;
	wire [1-1:0] node14;
	wire [1-1:0] node15;
	wire [1-1:0] node17;
	wire [1-1:0] node20;
	wire [1-1:0] node21;
	wire [1-1:0] node26;
	wire [1-1:0] node27;
	wire [1-1:0] node28;
	wire [1-1:0] node29;
	wire [1-1:0] node30;
	wire [1-1:0] node31;
	wire [1-1:0] node35;
	wire [1-1:0] node36;
	wire [1-1:0] node40;
	wire [1-1:0] node41;
	wire [1-1:0] node45;
	wire [1-1:0] node47;
	wire [1-1:0] node48;
	wire [1-1:0] node50;
	wire [1-1:0] node53;
	wire [1-1:0] node54;
	wire [1-1:0] node55;
	wire [1-1:0] node59;
	wire [1-1:0] node61;
	wire [1-1:0] node64;
	wire [1-1:0] node65;
	wire [1-1:0] node67;
	wire [1-1:0] node68;
	wire [1-1:0] node69;
	wire [1-1:0] node71;
	wire [1-1:0] node74;
	wire [1-1:0] node75;
	wire [1-1:0] node79;
	wire [1-1:0] node80;
	wire [1-1:0] node85;
	wire [1-1:0] node86;
	wire [1-1:0] node87;
	wire [1-1:0] node88;
	wire [1-1:0] node89;
	wire [1-1:0] node90;
	wire [1-1:0] node92;
	wire [1-1:0] node93;
	wire [1-1:0] node94;
	wire [1-1:0] node95;
	wire [1-1:0] node99;
	wire [1-1:0] node103;
	wire [1-1:0] node104;
	wire [1-1:0] node105;
	wire [1-1:0] node106;
	wire [1-1:0] node108;
	wire [1-1:0] node109;
	wire [1-1:0] node114;
	wire [1-1:0] node116;
	wire [1-1:0] node117;
	wire [1-1:0] node121;
	wire [1-1:0] node122;
	wire [1-1:0] node124;
	wire [1-1:0] node126;
	wire [1-1:0] node130;
	wire [1-1:0] node131;
	wire [1-1:0] node133;
	wire [1-1:0] node135;
	wire [1-1:0] node138;
	wire [1-1:0] node139;
	wire [1-1:0] node140;
	wire [1-1:0] node141;
	wire [1-1:0] node143;
	wire [1-1:0] node145;
	wire [1-1:0] node148;
	wire [1-1:0] node150;
	wire [1-1:0] node154;
	wire [1-1:0] node155;
	wire [1-1:0] node156;
	wire [1-1:0] node158;
	wire [1-1:0] node161;
	wire [1-1:0] node164;
	wire [1-1:0] node166;
	wire [1-1:0] node168;
	wire [1-1:0] node169;
	wire [1-1:0] node172;
	wire [1-1:0] node175;
	wire [1-1:0] node176;
	wire [1-1:0] node177;
	wire [1-1:0] node179;
	wire [1-1:0] node181;
	wire [1-1:0] node182;
	wire [1-1:0] node183;
	wire [1-1:0] node185;
	wire [1-1:0] node188;
	wire [1-1:0] node190;
	wire [1-1:0] node193;
	wire [1-1:0] node197;
	wire [1-1:0] node198;
	wire [1-1:0] node199;
	wire [1-1:0] node200;
	wire [1-1:0] node201;
	wire [1-1:0] node202;
	wire [1-1:0] node204;
	wire [1-1:0] node205;
	wire [1-1:0] node208;
	wire [1-1:0] node214;
	wire [1-1:0] node215;
	wire [1-1:0] node216;
	wire [1-1:0] node220;
	wire [1-1:0] node221;
	wire [1-1:0] node222;
	wire [1-1:0] node223;
	wire [1-1:0] node228;
	wire [1-1:0] node231;
	wire [1-1:0] node232;
	wire [1-1:0] node234;
	wire [1-1:0] node235;
	wire [1-1:0] node236;
	wire [1-1:0] node237;
	wire [1-1:0] node242;
	wire [1-1:0] node243;
	wire [1-1:0] node248;
	wire [1-1:0] node249;
	wire [1-1:0] node250;
	wire [1-1:0] node251;
	wire [1-1:0] node252;
	wire [1-1:0] node254;
	wire [1-1:0] node255;
	wire [1-1:0] node260;
	wire [1-1:0] node261;
	wire [1-1:0] node262;
	wire [1-1:0] node263;
	wire [1-1:0] node267;
	wire [1-1:0] node269;
	wire [1-1:0] node271;
	wire [1-1:0] node273;
	wire [1-1:0] node276;
	wire [1-1:0] node278;
	wire [1-1:0] node279;
	wire [1-1:0] node280;
	wire [1-1:0] node285;
	wire [1-1:0] node286;
	wire [1-1:0] node287;
	wire [1-1:0] node288;
	wire [1-1:0] node289;
	wire [1-1:0] node293;
	wire [1-1:0] node294;
	wire [1-1:0] node296;
	wire [1-1:0] node299;
	wire [1-1:0] node300;
	wire [1-1:0] node302;
	wire [1-1:0] node306;
	wire [1-1:0] node307;
	wire [1-1:0] node309;
	wire [1-1:0] node311;
	wire [1-1:0] node312;
	wire [1-1:0] node314;
	wire [1-1:0] node317;
	wire [1-1:0] node321;
	wire [1-1:0] node322;
	wire [1-1:0] node323;
	wire [1-1:0] node325;
	wire [1-1:0] node327;
	wire [1-1:0] node331;
	wire [1-1:0] node332;
	wire [1-1:0] node334;
	wire [1-1:0] node335;
	wire [1-1:0] node339;
	wire [1-1:0] node340;
	wire [1-1:0] node341;
	wire [1-1:0] node343;
	wire [1-1:0] node346;
	wire [1-1:0] node350;
	wire [1-1:0] node351;
	wire [1-1:0] node352;
	wire [1-1:0] node354;
	wire [1-1:0] node355;
	wire [1-1:0] node356;
	wire [1-1:0] node357;
	wire [1-1:0] node358;
	wire [1-1:0] node362;
	wire [1-1:0] node364;
	wire [1-1:0] node369;
	wire [1-1:0] node370;
	wire [1-1:0] node371;
	wire [1-1:0] node373;
	wire [1-1:0] node375;
	wire [1-1:0] node378;
	wire [1-1:0] node381;
	wire [1-1:0] node382;
	wire [1-1:0] node383;
	wire [1-1:0] node387;
	wire [1-1:0] node388;
	wire [1-1:0] node391;
	wire [1-1:0] node394;
	wire [1-1:0] node395;
	wire [1-1:0] node397;
	wire [1-1:0] node398;
	wire [1-1:0] node400;
	wire [1-1:0] node403;
	wire [1-1:0] node404;
	wire [1-1:0] node405;
	wire [1-1:0] node411;
	wire [1-1:0] node412;
	wire [1-1:0] node413;
	wire [1-1:0] node414;
	wire [1-1:0] node416;
	wire [1-1:0] node417;
	wire [1-1:0] node418;
	wire [1-1:0] node419;
	wire [1-1:0] node420;
	wire [1-1:0] node423;
	wire [1-1:0] node427;
	wire [1-1:0] node428;
	wire [1-1:0] node433;
	wire [1-1:0] node434;
	wire [1-1:0] node435;
	wire [1-1:0] node436;
	wire [1-1:0] node437;
	wire [1-1:0] node441;
	wire [1-1:0] node442;
	wire [1-1:0] node443;
	wire [1-1:0] node447;
	wire [1-1:0] node448;
	wire [1-1:0] node451;
	wire [1-1:0] node454;
	wire [1-1:0] node456;
	wire [1-1:0] node457;
	wire [1-1:0] node458;
	wire [1-1:0] node461;
	wire [1-1:0] node462;
	wire [1-1:0] node463;
	wire [1-1:0] node467;
	wire [1-1:0] node468;
	wire [1-1:0] node472;
	wire [1-1:0] node474;
	wire [1-1:0] node477;
	wire [1-1:0] node479;
	wire [1-1:0] node480;
	wire [1-1:0] node482;
	wire [1-1:0] node483;
	wire [1-1:0] node486;
	wire [1-1:0] node490;
	wire [1-1:0] node491;
	wire [1-1:0] node493;
	wire [1-1:0] node494;
	wire [1-1:0] node495;
	wire [1-1:0] node496;
	wire [1-1:0] node500;
	wire [1-1:0] node501;
	wire [1-1:0] node503;
	wire [1-1:0] node506;
	wire [1-1:0] node510;
	wire [1-1:0] node511;
	wire [1-1:0] node512;
	wire [1-1:0] node513;
	wire [1-1:0] node515;
	wire [1-1:0] node518;
	wire [1-1:0] node519;
	wire [1-1:0] node521;
	wire [1-1:0] node524;
	wire [1-1:0] node526;
	wire [1-1:0] node527;
	wire [1-1:0] node531;
	wire [1-1:0] node533;
	wire [1-1:0] node534;
	wire [1-1:0] node535;
	wire [1-1:0] node537;
	wire [1-1:0] node540;
	wire [1-1:0] node542;
	wire [1-1:0] node543;
	wire [1-1:0] node546;
	wire [1-1:0] node550;
	wire [1-1:0] node552;
	wire [1-1:0] node553;
	wire [1-1:0] node555;
	wire [1-1:0] node556;
	wire [1-1:0] node561;
	wire [1-1:0] node562;
	wire [1-1:0] node563;
	wire [1-1:0] node564;
	wire [1-1:0] node566;
	wire [1-1:0] node567;
	wire [1-1:0] node569;
	wire [1-1:0] node572;
	wire [1-1:0] node574;
	wire [1-1:0] node576;
	wire [1-1:0] node577;
	wire [1-1:0] node582;
	wire [1-1:0] node583;
	wire [1-1:0] node584;
	wire [1-1:0] node585;
	wire [1-1:0] node587;
	wire [1-1:0] node590;
	wire [1-1:0] node591;
	wire [1-1:0] node593;
	wire [1-1:0] node596;
	wire [1-1:0] node600;
	wire [1-1:0] node601;
	wire [1-1:0] node603;
	wire [1-1:0] node606;
	wire [1-1:0] node607;
	wire [1-1:0] node608;
	wire [1-1:0] node612;
	wire [1-1:0] node614;
	wire [1-1:0] node617;
	wire [1-1:0] node618;
	wire [1-1:0] node620;
	wire [1-1:0] node621;
	wire [1-1:0] node622;
	wire [1-1:0] node626;
	wire [1-1:0] node627;
	wire [1-1:0] node628;
	wire [1-1:0] node630;
	wire [1-1:0] node633;
	wire [1-1:0] node634;
	wire [1-1:0] node635;
	wire [1-1:0] node640;
	wire [1-1:0] node641;
	wire [1-1:0] node643;
	wire [1-1:0] node645;
	wire [1-1:0] node648;
	wire [1-1:0] node652;
	wire [1-1:0] node653;
	wire [1-1:0] node654;
	wire [1-1:0] node655;
	wire [1-1:0] node657;
	wire [1-1:0] node658;
	wire [1-1:0] node659;
	wire [1-1:0] node663;
	wire [1-1:0] node664;
	wire [1-1:0] node665;
	wire [1-1:0] node669;
	wire [1-1:0] node670;
	wire [1-1:0] node675;
	wire [1-1:0] node676;
	wire [1-1:0] node677;
	wire [1-1:0] node678;
	wire [1-1:0] node680;
	wire [1-1:0] node683;
	wire [1-1:0] node684;
	wire [1-1:0] node685;
	wire [1-1:0] node689;
	wire [1-1:0] node690;
	wire [1-1:0] node695;
	wire [1-1:0] node696;
	wire [1-1:0] node698;
	wire [1-1:0] node701;
	wire [1-1:0] node702;
	wire [1-1:0] node704;
	wire [1-1:0] node707;
	wire [1-1:0] node708;
	wire [1-1:0] node712;
	wire [1-1:0] node713;
	wire [1-1:0] node715;
	wire [1-1:0] node716;
	wire [1-1:0] node717;
	wire [1-1:0] node718;
	wire [1-1:0] node722;
	wire [1-1:0] node723;
	wire [1-1:0] node727;
	wire [1-1:0] node728;
	wire [1-1:0] node733;
	wire [1-1:0] node734;
	wire [1-1:0] node735;
	wire [1-1:0] node736;
	wire [1-1:0] node737;
	wire [1-1:0] node738;
	wire [1-1:0] node739;
	wire [1-1:0] node740;
	wire [1-1:0] node741;
	wire [1-1:0] node743;
	wire [1-1:0] node744;
	wire [1-1:0] node745;
	wire [1-1:0] node751;
	wire [1-1:0] node752;
	wire [1-1:0] node753;
	wire [1-1:0] node756;
	wire [1-1:0] node757;
	wire [1-1:0] node759;
	wire [1-1:0] node763;
	wire [1-1:0] node765;
	wire [1-1:0] node766;
	wire [1-1:0] node768;
	wire [1-1:0] node769;
	wire [1-1:0] node774;
	wire [1-1:0] node775;
	wire [1-1:0] node776;
	wire [1-1:0] node777;
	wire [1-1:0] node779;
	wire [1-1:0] node783;
	wire [1-1:0] node784;
	wire [1-1:0] node785;
	wire [1-1:0] node786;
	wire [1-1:0] node791;
	wire [1-1:0] node792;
	wire [1-1:0] node794;
	wire [1-1:0] node798;
	wire [1-1:0] node799;
	wire [1-1:0] node800;
	wire [1-1:0] node801;
	wire [1-1:0] node804;
	wire [1-1:0] node805;
	wire [1-1:0] node807;
	wire [1-1:0] node812;
	wire [1-1:0] node813;
	wire [1-1:0] node814;
	wire [1-1:0] node816;
	wire [1-1:0] node821;
	wire [1-1:0] node822;
	wire [1-1:0] node823;
	wire [1-1:0] node824;
	wire [1-1:0] node826;
	wire [1-1:0] node828;
	wire [1-1:0] node829;
	wire [1-1:0] node830;
	wire [1-1:0] node836;
	wire [1-1:0] node837;
	wire [1-1:0] node838;
	wire [1-1:0] node839;
	wire [1-1:0] node841;
	wire [1-1:0] node845;
	wire [1-1:0] node846;
	wire [1-1:0] node850;
	wire [1-1:0] node851;
	wire [1-1:0] node853;
	wire [1-1:0] node854;
	wire [1-1:0] node858;
	wire [1-1:0] node859;
	wire [1-1:0] node860;
	wire [1-1:0] node865;
	wire [1-1:0] node866;
	wire [1-1:0] node868;
	wire [1-1:0] node869;
	wire [1-1:0] node870;
	wire [1-1:0] node871;
	wire [1-1:0] node878;
	wire [1-1:0] node879;
	wire [1-1:0] node880;
	wire [1-1:0] node881;
	wire [1-1:0] node882;
	wire [1-1:0] node884;
	wire [1-1:0] node885;
	wire [1-1:0] node886;
	wire [1-1:0] node889;
	wire [1-1:0] node890;
	wire [1-1:0] node894;
	wire [1-1:0] node896;
	wire [1-1:0] node900;
	wire [1-1:0] node901;
	wire [1-1:0] node902;
	wire [1-1:0] node903;
	wire [1-1:0] node905;
	wire [1-1:0] node909;
	wire [1-1:0] node910;
	wire [1-1:0] node911;
	wire [1-1:0] node914;
	wire [1-1:0] node917;
	wire [1-1:0] node920;
	wire [1-1:0] node921;
	wire [1-1:0] node923;
	wire [1-1:0] node926;
	wire [1-1:0] node928;
	wire [1-1:0] node929;
	wire [1-1:0] node933;
	wire [1-1:0] node935;
	wire [1-1:0] node936;
	wire [1-1:0] node937;
	wire [1-1:0] node938;
	wire [1-1:0] node940;
	wire [1-1:0] node944;
	wire [1-1:0] node946;
	wire [1-1:0] node950;
	wire [1-1:0] node951;
	wire [1-1:0] node952;
	wire [1-1:0] node953;
	wire [1-1:0] node954;
	wire [1-1:0] node955;
	wire [1-1:0] node959;
	wire [1-1:0] node961;
	wire [1-1:0] node962;
	wire [1-1:0] node964;
	wire [1-1:0] node968;
	wire [1-1:0] node970;
	wire [1-1:0] node971;
	wire [1-1:0] node973;
	wire [1-1:0] node977;
	wire [1-1:0] node979;
	wire [1-1:0] node980;
	wire [1-1:0] node981;
	wire [1-1:0] node983;
	wire [1-1:0] node987;
	wire [1-1:0] node988;
	wire [1-1:0] node992;
	wire [1-1:0] node993;
	wire [1-1:0] node994;
	wire [1-1:0] node996;
	wire [1-1:0] node997;
	wire [1-1:0] node998;
	wire [1-1:0] node1003;
	wire [1-1:0] node1004;
	wire [1-1:0] node1006;
	wire [1-1:0] node1009;
	wire [1-1:0] node1011;
	wire [1-1:0] node1012;
	wire [1-1:0] node1013;
	wire [1-1:0] node1018;
	wire [1-1:0] node1019;
	wire [1-1:0] node1020;
	wire [1-1:0] node1022;
	wire [1-1:0] node1026;
	wire [1-1:0] node1028;
	wire [1-1:0] node1029;
	wire [1-1:0] node1033;
	wire [1-1:0] node1034;
	wire [1-1:0] node1035;
	wire [1-1:0] node1036;
	wire [1-1:0] node1038;
	wire [1-1:0] node1039;
	wire [1-1:0] node1041;
	wire [1-1:0] node1044;
	wire [1-1:0] node1045;
	wire [1-1:0] node1047;
	wire [1-1:0] node1048;
	wire [1-1:0] node1050;
	wire [1-1:0] node1054;
	wire [1-1:0] node1056;
	wire [1-1:0] node1057;
	wire [1-1:0] node1062;
	wire [1-1:0] node1063;
	wire [1-1:0] node1064;
	wire [1-1:0] node1065;
	wire [1-1:0] node1066;
	wire [1-1:0] node1067;
	wire [1-1:0] node1071;
	wire [1-1:0] node1073;
	wire [1-1:0] node1076;
	wire [1-1:0] node1078;
	wire [1-1:0] node1079;
	wire [1-1:0] node1080;
	wire [1-1:0] node1085;
	wire [1-1:0] node1086;
	wire [1-1:0] node1087;
	wire [1-1:0] node1089;
	wire [1-1:0] node1093;
	wire [1-1:0] node1094;
	wire [1-1:0] node1098;
	wire [1-1:0] node1099;
	wire [1-1:0] node1101;
	wire [1-1:0] node1102;
	wire [1-1:0] node1104;
	wire [1-1:0] node1107;
	wire [1-1:0] node1108;
	wire [1-1:0] node1110;
	wire [1-1:0] node1111;
	wire [1-1:0] node1113;
	wire [1-1:0] node1116;
	wire [1-1:0] node1117;
	wire [1-1:0] node1123;
	wire [1-1:0] node1124;
	wire [1-1:0] node1125;
	wire [1-1:0] node1126;
	wire [1-1:0] node1127;
	wire [1-1:0] node1129;
	wire [1-1:0] node1130;
	wire [1-1:0] node1135;
	wire [1-1:0] node1136;
	wire [1-1:0] node1137;
	wire [1-1:0] node1138;
	wire [1-1:0] node1139;
	wire [1-1:0] node1141;
	wire [1-1:0] node1142;
	wire [1-1:0] node1145;
	wire [1-1:0] node1148;
	wire [1-1:0] node1151;
	wire [1-1:0] node1153;
	wire [1-1:0] node1157;
	wire [1-1:0] node1158;
	wire [1-1:0] node1159;
	wire [1-1:0] node1163;
	wire [1-1:0] node1164;
	wire [1-1:0] node1165;
	wire [1-1:0] node1169;
	wire [1-1:0] node1170;
	wire [1-1:0] node1172;
	wire [1-1:0] node1176;
	wire [1-1:0] node1177;
	wire [1-1:0] node1179;
	wire [1-1:0] node1180;
	wire [1-1:0] node1181;
	wire [1-1:0] node1184;
	wire [1-1:0] node1185;
	wire [1-1:0] node1188;
	wire [1-1:0] node1191;
	wire [1-1:0] node1193;
	wire [1-1:0] node1197;
	wire [1-1:0] node1198;
	wire [1-1:0] node1199;
	wire [1-1:0] node1201;
	wire [1-1:0] node1202;
	wire [1-1:0] node1203;
	wire [1-1:0] node1204;
	wire [1-1:0] node1205;
	wire [1-1:0] node1206;
	wire [1-1:0] node1214;
	wire [1-1:0] node1215;
	wire [1-1:0] node1216;
	wire [1-1:0] node1217;
	wire [1-1:0] node1219;
	wire [1-1:0] node1222;
	wire [1-1:0] node1224;
	wire [1-1:0] node1227;
	wire [1-1:0] node1228;
	wire [1-1:0] node1232;
	wire [1-1:0] node1234;
	wire [1-1:0] node1235;
	wire [1-1:0] node1236;
	wire [1-1:0] node1237;
	wire [1-1:0] node1241;
	wire [1-1:0] node1243;
	wire [1-1:0] node1246;
	wire [1-1:0] node1247;
	wire [1-1:0] node1251;
	wire [1-1:0] node1252;
	wire [1-1:0] node1254;
	wire [1-1:0] node1255;
	wire [1-1:0] node1256;
	wire [1-1:0] node1257;
	wire [1-1:0] node1261;
	wire [1-1:0] node1262;
	wire [1-1:0] node1264;
	wire [1-1:0] node1268;
	wire [1-1:0] node1270;
	wire [1-1:0] node1274;
	wire [1-1:0] node1275;
	wire [1-1:0] node1276;
	wire [1-1:0] node1278;
	wire [1-1:0] node1279;
	wire [1-1:0] node1281;
	wire [1-1:0] node1284;
	wire [1-1:0] node1285;
	wire [1-1:0] node1287;
	wire [1-1:0] node1290;
	wire [1-1:0] node1292;
	wire [1-1:0] node1296;
	wire [1-1:0] node1297;
	wire [1-1:0] node1298;
	wire [1-1:0] node1299;
	wire [1-1:0] node1300;
	wire [1-1:0] node1301;
	wire [1-1:0] node1305;
	wire [1-1:0] node1306;
	wire [1-1:0] node1307;
	wire [1-1:0] node1311;
	wire [1-1:0] node1312;
	wire [1-1:0] node1317;
	wire [1-1:0] node1318;
	wire [1-1:0] node1319;
	wire [1-1:0] node1321;
	wire [1-1:0] node1324;
	wire [1-1:0] node1326;
	wire [1-1:0] node1329;
	wire [1-1:0] node1331;
	wire [1-1:0] node1334;
	wire [1-1:0] node1335;
	wire [1-1:0] node1337;
	wire [1-1:0] node1338;
	wire [1-1:0] node1339;
	wire [1-1:0] node1341;
	wire [1-1:0] node1344;
	wire [1-1:0] node1345;
	wire [1-1:0] node1349;
	wire [1-1:0] node1351;
	wire [1-1:0] node1355;
	wire [1-1:0] node1356;
	wire [1-1:0] node1357;
	wire [1-1:0] node1358;
	wire [1-1:0] node1359;
	wire [1-1:0] node1360;
	wire [1-1:0] node1361;
	wire [1-1:0] node1362;
	wire [1-1:0] node1364;
	wire [1-1:0] node1366;
	wire [1-1:0] node1368;
	wire [1-1:0] node1371;
	wire [1-1:0] node1372;
	wire [1-1:0] node1374;
	wire [1-1:0] node1377;
	wire [1-1:0] node1380;
	wire [1-1:0] node1381;
	wire [1-1:0] node1383;
	wire [1-1:0] node1384;
	wire [1-1:0] node1385;
	wire [1-1:0] node1391;
	wire [1-1:0] node1392;
	wire [1-1:0] node1393;
	wire [1-1:0] node1394;
	wire [1-1:0] node1397;
	wire [1-1:0] node1398;
	wire [1-1:0] node1401;
	wire [1-1:0] node1405;
	wire [1-1:0] node1406;
	wire [1-1:0] node1407;
	wire [1-1:0] node1408;
	wire [1-1:0] node1409;
	wire [1-1:0] node1415;
	wire [1-1:0] node1416;
	wire [1-1:0] node1417;
	wire [1-1:0] node1421;
	wire [1-1:0] node1423;
	wire [1-1:0] node1426;
	wire [1-1:0] node1428;
	wire [1-1:0] node1429;
	wire [1-1:0] node1430;
	wire [1-1:0] node1431;
	wire [1-1:0] node1432;
	wire [1-1:0] node1436;
	wire [1-1:0] node1437;
	wire [1-1:0] node1441;
	wire [1-1:0] node1443;
	wire [1-1:0] node1447;
	wire [1-1:0] node1448;
	wire [1-1:0] node1449;
	wire [1-1:0] node1450;
	wire [1-1:0] node1451;
	wire [1-1:0] node1453;
	wire [1-1:0] node1454;
	wire [1-1:0] node1456;
	wire [1-1:0] node1459;
	wire [1-1:0] node1461;
	wire [1-1:0] node1465;
	wire [1-1:0] node1466;
	wire [1-1:0] node1467;
	wire [1-1:0] node1468;
	wire [1-1:0] node1472;
	wire [1-1:0] node1473;
	wire [1-1:0] node1474;
	wire [1-1:0] node1478;
	wire [1-1:0] node1481;
	wire [1-1:0] node1483;
	wire [1-1:0] node1484;
	wire [1-1:0] node1485;
	wire [1-1:0] node1489;
	wire [1-1:0] node1491;
	wire [1-1:0] node1493;
	wire [1-1:0] node1496;
	wire [1-1:0] node1497;
	wire [1-1:0] node1499;
	wire [1-1:0] node1500;
	wire [1-1:0] node1502;
	wire [1-1:0] node1504;
	wire [1-1:0] node1509;
	wire [1-1:0] node1510;
	wire [1-1:0] node1511;
	wire [1-1:0] node1512;
	wire [1-1:0] node1514;
	wire [1-1:0] node1517;
	wire [1-1:0] node1518;
	wire [1-1:0] node1519;
	wire [1-1:0] node1520;
	wire [1-1:0] node1525;
	wire [1-1:0] node1526;
	wire [1-1:0] node1528;
	wire [1-1:0] node1531;
	wire [1-1:0] node1533;
	wire [1-1:0] node1536;
	wire [1-1:0] node1537;
	wire [1-1:0] node1539;
	wire [1-1:0] node1540;
	wire [1-1:0] node1545;
	wire [1-1:0] node1546;
	wire [1-1:0] node1547;
	wire [1-1:0] node1549;
	wire [1-1:0] node1552;
	wire [1-1:0] node1553;
	wire [1-1:0] node1554;
	wire [1-1:0] node1558;
	wire [1-1:0] node1561;
	wire [1-1:0] node1563;
	wire [1-1:0] node1564;
	wire [1-1:0] node1565;
	wire [1-1:0] node1567;
	wire [1-1:0] node1571;
	wire [1-1:0] node1573;
	wire [1-1:0] node1575;
	wire [1-1:0] node1578;
	wire [1-1:0] node1579;
	wire [1-1:0] node1580;
	wire [1-1:0] node1582;
	wire [1-1:0] node1583;
	wire [1-1:0] node1584;
	wire [1-1:0] node1586;
	wire [1-1:0] node1587;
	wire [1-1:0] node1591;
	wire [1-1:0] node1593;
	wire [1-1:0] node1597;
	wire [1-1:0] node1598;
	wire [1-1:0] node1599;
	wire [1-1:0] node1600;
	wire [1-1:0] node1601;
	wire [1-1:0] node1602;
	wire [1-1:0] node1606;
	wire [1-1:0] node1608;
	wire [1-1:0] node1611;
	wire [1-1:0] node1613;
	wire [1-1:0] node1616;
	wire [1-1:0] node1618;
	wire [1-1:0] node1619;
	wire [1-1:0] node1620;
	wire [1-1:0] node1623;
	wire [1-1:0] node1624;
	wire [1-1:0] node1628;
	wire [1-1:0] node1629;
	wire [1-1:0] node1631;
	wire [1-1:0] node1633;
	wire [1-1:0] node1636;
	wire [1-1:0] node1637;
	wire [1-1:0] node1641;
	wire [1-1:0] node1643;
	wire [1-1:0] node1644;
	wire [1-1:0] node1645;
	wire [1-1:0] node1646;
	wire [1-1:0] node1647;
	wire [1-1:0] node1650;
	wire [1-1:0] node1653;
	wire [1-1:0] node1655;
	wire [1-1:0] node1658;
	wire [1-1:0] node1660;
	wire [1-1:0] node1664;
	wire [1-1:0] node1665;
	wire [1-1:0] node1666;
	wire [1-1:0] node1667;
	wire [1-1:0] node1669;
	wire [1-1:0] node1670;
	wire [1-1:0] node1671;
	wire [1-1:0] node1672;
	wire [1-1:0] node1674;
	wire [1-1:0] node1676;
	wire [1-1:0] node1682;
	wire [1-1:0] node1683;
	wire [1-1:0] node1684;
	wire [1-1:0] node1685;
	wire [1-1:0] node1687;
	wire [1-1:0] node1690;
	wire [1-1:0] node1691;
	wire [1-1:0] node1692;
	wire [1-1:0] node1695;
	wire [1-1:0] node1700;
	wire [1-1:0] node1701;
	wire [1-1:0] node1702;
	wire [1-1:0] node1706;
	wire [1-1:0] node1707;
	wire [1-1:0] node1709;
	wire [1-1:0] node1712;
	wire [1-1:0] node1714;
	wire [1-1:0] node1717;
	wire [1-1:0] node1718;
	wire [1-1:0] node1720;
	wire [1-1:0] node1721;
	wire [1-1:0] node1722;
	wire [1-1:0] node1726;
	wire [1-1:0] node1728;
	wire [1-1:0] node1732;
	wire [1-1:0] node1733;
	wire [1-1:0] node1734;
	wire [1-1:0] node1736;
	wire [1-1:0] node1737;
	wire [1-1:0] node1738;
	wire [1-1:0] node1739;
	wire [1-1:0] node1740;
	wire [1-1:0] node1747;
	wire [1-1:0] node1748;
	wire [1-1:0] node1749;
	wire [1-1:0] node1750;
	wire [1-1:0] node1751;
	wire [1-1:0] node1754;
	wire [1-1:0] node1755;
	wire [1-1:0] node1759;
	wire [1-1:0] node1761;
	wire [1-1:0] node1765;
	wire [1-1:0] node1766;
	wire [1-1:0] node1767;
	wire [1-1:0] node1769;
	wire [1-1:0] node1772;
	wire [1-1:0] node1773;
	wire [1-1:0] node1777;
	wire [1-1:0] node1779;
	wire [1-1:0] node1782;
	wire [1-1:0] node1783;
	wire [1-1:0] node1785;
	wire [1-1:0] node1786;
	wire [1-1:0] node1787;
	wire [1-1:0] node1788;
	wire [1-1:0] node1791;
	wire [1-1:0] node1794;
	wire [1-1:0] node1797;
	wire [1-1:0] node1799;
	wire [1-1:0] node1803;
	wire [1-1:0] node1804;
	wire [1-1:0] node1805;
	wire [1-1:0] node1806;
	wire [1-1:0] node1807;
	wire [1-1:0] node1809;
	wire [1-1:0] node1810;
	wire [1-1:0] node1811;
	wire [1-1:0] node1812;
	wire [1-1:0] node1815;
	wire [1-1:0] node1817;
	wire [1-1:0] node1820;
	wire [1-1:0] node1822;
	wire [1-1:0] node1826;
	wire [1-1:0] node1827;
	wire [1-1:0] node1828;
	wire [1-1:0] node1829;
	wire [1-1:0] node1830;
	wire [1-1:0] node1831;
	wire [1-1:0] node1832;
	wire [1-1:0] node1836;
	wire [1-1:0] node1839;
	wire [1-1:0] node1844;
	wire [1-1:0] node1845;
	wire [1-1:0] node1846;
	wire [1-1:0] node1848;
	wire [1-1:0] node1851;
	wire [1-1:0] node1853;
	wire [1-1:0] node1856;
	wire [1-1:0] node1858;
	wire [1-1:0] node1861;
	wire [1-1:0] node1863;
	wire [1-1:0] node1864;
	wire [1-1:0] node1865;
	wire [1-1:0] node1867;
	wire [1-1:0] node1870;
	wire [1-1:0] node1871;
	wire [1-1:0] node1872;
	wire [1-1:0] node1876;
	wire [1-1:0] node1880;
	wire [1-1:0] node1881;
	wire [1-1:0] node1882;
	wire [1-1:0] node1884;
	wire [1-1:0] node1885;
	wire [1-1:0] node1886;
	wire [1-1:0] node1890;
	wire [1-1:0] node1891;
	wire [1-1:0] node1892;
	wire [1-1:0] node1894;
	wire [1-1:0] node1898;
	wire [1-1:0] node1902;
	wire [1-1:0] node1903;
	wire [1-1:0] node1904;
	wire [1-1:0] node1905;
	wire [1-1:0] node1906;
	wire [1-1:0] node1910;
	wire [1-1:0] node1912;
	wire [1-1:0] node1914;
	wire [1-1:0] node1917;
	wire [1-1:0] node1918;
	wire [1-1:0] node1920;
	wire [1-1:0] node1921;
	wire [1-1:0] node1922;
	wire [1-1:0] node1927;
	wire [1-1:0] node1929;
	wire [1-1:0] node1931;
	wire [1-1:0] node1933;
	wire [1-1:0] node1936;
	wire [1-1:0] node1938;
	wire [1-1:0] node1939;
	wire [1-1:0] node1940;
	wire [1-1:0] node1941;
	wire [1-1:0] node1944;
	wire [1-1:0] node1946;
	wire [1-1:0] node1949;
	wire [1-1:0] node1950;
	wire [1-1:0] node1955;
	wire [1-1:0] node1956;
	wire [1-1:0] node1957;
	wire [1-1:0] node1958;
	wire [1-1:0] node1960;
	wire [1-1:0] node1961;
	wire [1-1:0] node1962;
	wire [1-1:0] node1964;
	wire [1-1:0] node1968;
	wire [1-1:0] node1969;
	wire [1-1:0] node1974;
	wire [1-1:0] node1975;
	wire [1-1:0] node1976;
	wire [1-1:0] node1977;
	wire [1-1:0] node1981;
	wire [1-1:0] node1982;
	wire [1-1:0] node1984;
	wire [1-1:0] node1987;
	wire [1-1:0] node1989;
	wire [1-1:0] node1992;
	wire [1-1:0] node1994;
	wire [1-1:0] node1995;
	wire [1-1:0] node1996;
	wire [1-1:0] node1998;
	wire [1-1:0] node2001;
	wire [1-1:0] node2002;
	wire [1-1:0] node2006;
	wire [1-1:0] node2008;
	wire [1-1:0] node2011;
	wire [1-1:0] node2013;
	wire [1-1:0] node2014;
	wire [1-1:0] node2015;
	wire [1-1:0] node2016;
	wire [1-1:0] node2018;
	wire [1-1:0] node2021;
	wire [1-1:0] node2023;
	wire [1-1:0] node2026;
	wire [1-1:0] node2028;
	wire [1-1:0] node2032;
	wire [1-1:0] node2033;
	wire [1-1:0] node2034;
	wire [1-1:0] node2035;
	wire [1-1:0] node2037;
	wire [1-1:0] node2038;
	wire [1-1:0] node2039;
	wire [1-1:0] node2040;
	wire [1-1:0] node2044;
	wire [1-1:0] node2045;
	wire [1-1:0] node2046;
	wire [1-1:0] node2050;
	wire [1-1:0] node2051;
	wire [1-1:0] node2056;
	wire [1-1:0] node2057;
	wire [1-1:0] node2058;
	wire [1-1:0] node2059;
	wire [1-1:0] node2063;
	wire [1-1:0] node2064;
	wire [1-1:0] node2065;
	wire [1-1:0] node2069;
	wire [1-1:0] node2070;
	wire [1-1:0] node2074;
	wire [1-1:0] node2076;
	wire [1-1:0] node2077;
	wire [1-1:0] node2078;
	wire [1-1:0] node2080;
	wire [1-1:0] node2083;
	wire [1-1:0] node2084;
	wire [1-1:0] node2088;
	wire [1-1:0] node2090;
	wire [1-1:0] node2093;
	wire [1-1:0] node2095;
	wire [1-1:0] node2096;
	wire [1-1:0] node2097;
	wire [1-1:0] node2099;
	wire [1-1:0] node2102;
	wire [1-1:0] node2103;
	wire [1-1:0] node2104;
	wire [1-1:0] node2108;
	wire [1-1:0] node2109;
	wire [1-1:0] node2114;
	wire [1-1:0] node2115;
	wire [1-1:0] node2116;
	wire [1-1:0] node2117;
	wire [1-1:0] node2118;
	wire [1-1:0] node2119;
	wire [1-1:0] node2120;
	wire [1-1:0] node2121;
	wire [1-1:0] node2122;
	wire [1-1:0] node2124;
	wire [1-1:0] node2126;
	wire [1-1:0] node2130;
	wire [1-1:0] node2131;
	wire [1-1:0] node2132;
	wire [1-1:0] node2133;
	wire [1-1:0] node2137;
	wire [1-1:0] node2139;
	wire [1-1:0] node2140;
	wire [1-1:0] node2144;
	wire [1-1:0] node2146;
	wire [1-1:0] node2147;
	wire [1-1:0] node2149;
	wire [1-1:0] node2152;
	wire [1-1:0] node2154;
	wire [1-1:0] node2155;
	wire [1-1:0] node2158;
	wire [1-1:0] node2161;
	wire [1-1:0] node2163;
	wire [1-1:0] node2164;
	wire [1-1:0] node2165;
	wire [1-1:0] node2167;
	wire [1-1:0] node2170;
	wire [1-1:0] node2172;
	wire [1-1:0] node2173;
	wire [1-1:0] node2178;
	wire [1-1:0] node2179;
	wire [1-1:0] node2181;
	wire [1-1:0] node2182;
	wire [1-1:0] node2183;
	wire [1-1:0] node2185;
	wire [1-1:0] node2188;
	wire [1-1:0] node2189;
	wire [1-1:0] node2191;
	wire [1-1:0] node2192;
	wire [1-1:0] node2196;
	wire [1-1:0] node2200;
	wire [1-1:0] node2201;
	wire [1-1:0] node2202;
	wire [1-1:0] node2203;
	wire [1-1:0] node2205;
	wire [1-1:0] node2206;
	wire [1-1:0] node2209;
	wire [1-1:0] node2213;
	wire [1-1:0] node2214;
	wire [1-1:0] node2215;
	wire [1-1:0] node2217;
	wire [1-1:0] node2220;
	wire [1-1:0] node2222;
	wire [1-1:0] node2225;
	wire [1-1:0] node2227;
	wire [1-1:0] node2230;
	wire [1-1:0] node2231;
	wire [1-1:0] node2233;
	wire [1-1:0] node2235;
	wire [1-1:0] node2237;
	wire [1-1:0] node2241;
	wire [1-1:0] node2242;
	wire [1-1:0] node2243;
	wire [1-1:0] node2245;
	wire [1-1:0] node2246;
	wire [1-1:0] node2247;
	wire [1-1:0] node2248;
	wire [1-1:0] node2249;
	wire [1-1:0] node2253;
	wire [1-1:0] node2256;
	wire [1-1:0] node2257;
	wire [1-1:0] node2262;
	wire [1-1:0] node2263;
	wire [1-1:0] node2264;
	wire [1-1:0] node2266;
	wire [1-1:0] node2269;
	wire [1-1:0] node2270;
	wire [1-1:0] node2271;
	wire [1-1:0] node2275;
	wire [1-1:0] node2276;
	wire [1-1:0] node2280;
	wire [1-1:0] node2282;
	wire [1-1:0] node2283;
	wire [1-1:0] node2284;
	wire [1-1:0] node2285;
	wire [1-1:0] node2290;
	wire [1-1:0] node2292;
	wire [1-1:0] node2295;
	wire [1-1:0] node2297;
	wire [1-1:0] node2298;
	wire [1-1:0] node2299;
	wire [1-1:0] node2301;
	wire [1-1:0] node2304;
	wire [1-1:0] node2305;
	wire [1-1:0] node2307;
	wire [1-1:0] node2309;
	wire [1-1:0] node2311;
	wire [1-1:0] node2314;
	wire [1-1:0] node2318;
	wire [1-1:0] node2319;
	wire [1-1:0] node2320;
	wire [1-1:0] node2321;
	wire [1-1:0] node2322;
	wire [1-1:0] node2323;
	wire [1-1:0] node2325;
	wire [1-1:0] node2327;
	wire [1-1:0] node2329;
	wire [1-1:0] node2333;
	wire [1-1:0] node2334;
	wire [1-1:0] node2335;
	wire [1-1:0] node2336;
	wire [1-1:0] node2338;
	wire [1-1:0] node2341;
	wire [1-1:0] node2343;
	wire [1-1:0] node2347;
	wire [1-1:0] node2348;
	wire [1-1:0] node2349;
	wire [1-1:0] node2353;
	wire [1-1:0] node2355;
	wire [1-1:0] node2358;
	wire [1-1:0] node2359;
	wire [1-1:0] node2361;
	wire [1-1:0] node2362;
	wire [1-1:0] node2363;
	wire [1-1:0] node2367;
	wire [1-1:0] node2369;
	wire [1-1:0] node2373;
	wire [1-1:0] node2374;
	wire [1-1:0] node2375;
	wire [1-1:0] node2376;
	wire [1-1:0] node2377;
	wire [1-1:0] node2381;
	wire [1-1:0] node2382;
	wire [1-1:0] node2383;
	wire [1-1:0] node2387;
	wire [1-1:0] node2389;
	wire [1-1:0] node2390;
	wire [1-1:0] node2393;
	wire [1-1:0] node2396;
	wire [1-1:0] node2397;
	wire [1-1:0] node2398;
	wire [1-1:0] node2400;
	wire [1-1:0] node2405;
	wire [1-1:0] node2406;
	wire [1-1:0] node2407;
	wire [1-1:0] node2408;
	wire [1-1:0] node2409;
	wire [1-1:0] node2413;
	wire [1-1:0] node2414;
	wire [1-1:0] node2418;
	wire [1-1:0] node2420;
	wire [1-1:0] node2423;
	wire [1-1:0] node2425;
	wire [1-1:0] node2426;
	wire [1-1:0] node2428;
	wire [1-1:0] node2431;
	wire [1-1:0] node2432;
	wire [1-1:0] node2433;
	wire [1-1:0] node2434;
	wire [1-1:0] node2435;
	wire [1-1:0] node2438;
	wire [1-1:0] node2441;
	wire [1-1:0] node2443;
	wire [1-1:0] node2446;
	wire [1-1:0] node2448;
	wire [1-1:0] node2452;
	wire [1-1:0] node2453;
	wire [1-1:0] node2454;
	wire [1-1:0] node2456;
	wire [1-1:0] node2457;
	wire [1-1:0] node2458;
	wire [1-1:0] node2460;
	wire [1-1:0] node2461;
	wire [1-1:0] node2465;
	wire [1-1:0] node2466;
	wire [1-1:0] node2471;
	wire [1-1:0] node2472;
	wire [1-1:0] node2473;
	wire [1-1:0] node2474;
	wire [1-1:0] node2478;
	wire [1-1:0] node2479;
	wire [1-1:0] node2481;
	wire [1-1:0] node2484;
	wire [1-1:0] node2485;
	wire [1-1:0] node2489;
	wire [1-1:0] node2491;
	wire [1-1:0] node2493;
	wire [1-1:0] node2494;
	wire [1-1:0] node2495;
	wire [1-1:0] node2499;
	wire [1-1:0] node2500;
	wire [1-1:0] node2504;
	wire [1-1:0] node2505;
	wire [1-1:0] node2507;
	wire [1-1:0] node2508;
	wire [1-1:0] node2509;
	wire [1-1:0] node2510;
	wire [1-1:0] node2513;
	wire [1-1:0] node2515;
	wire [1-1:0] node2516;
	wire [1-1:0] node2520;
	wire [1-1:0] node2523;
	wire [1-1:0] node2524;
	wire [1-1:0] node2525;
	wire [1-1:0] node2529;
	wire [1-1:0] node2530;
	wire [1-1:0] node2531;
	wire [1-1:0] node2535;
	wire [1-1:0] node2539;
	wire [1-1:0] node2540;
	wire [1-1:0] node2541;
	wire [1-1:0] node2542;
	wire [1-1:0] node2543;
	wire [1-1:0] node2544;
	wire [1-1:0] node2546;
	wire [1-1:0] node2547;
	wire [1-1:0] node2548;
	wire [1-1:0] node2550;
	wire [1-1:0] node2553;
	wire [1-1:0] node2555;
	wire [1-1:0] node2558;
	wire [1-1:0] node2560;
	wire [1-1:0] node2564;
	wire [1-1:0] node2565;
	wire [1-1:0] node2566;
	wire [1-1:0] node2567;
	wire [1-1:0] node2571;
	wire [1-1:0] node2572;
	wire [1-1:0] node2573;
	wire [1-1:0] node2577;
	wire [1-1:0] node2579;
	wire [1-1:0] node2582;
	wire [1-1:0] node2584;
	wire [1-1:0] node2585;
	wire [1-1:0] node2586;
	wire [1-1:0] node2590;
	wire [1-1:0] node2591;
	wire [1-1:0] node2592;
	wire [1-1:0] node2597;
	wire [1-1:0] node2599;
	wire [1-1:0] node2600;
	wire [1-1:0] node2601;
	wire [1-1:0] node2602;
	wire [1-1:0] node2603;
	wire [1-1:0] node2607;
	wire [1-1:0] node2608;
	wire [1-1:0] node2612;
	wire [1-1:0] node2614;
	wire [1-1:0] node2618;
	wire [1-1:0] node2619;
	wire [1-1:0] node2620;
	wire [1-1:0] node2622;
	wire [1-1:0] node2623;
	wire [1-1:0] node2624;
	wire [1-1:0] node2626;
	wire [1-1:0] node2629;
	wire [1-1:0] node2630;
	wire [1-1:0] node2634;
	wire [1-1:0] node2636;
	wire [1-1:0] node2640;
	wire [1-1:0] node2641;
	wire [1-1:0] node2642;
	wire [1-1:0] node2643;
	wire [1-1:0] node2644;
	wire [1-1:0] node2645;
	wire [1-1:0] node2649;
	wire [1-1:0] node2650;
	wire [1-1:0] node2652;
	wire [1-1:0] node2657;
	wire [1-1:0] node2658;
	wire [1-1:0] node2659;
	wire [1-1:0] node2660;
	wire [1-1:0] node2662;
	wire [1-1:0] node2666;
	wire [1-1:0] node2668;
	wire [1-1:0] node2671;
	wire [1-1:0] node2672;
	wire [1-1:0] node2676;
	wire [1-1:0] node2678;
	wire [1-1:0] node2679;
	wire [1-1:0] node2680;
	wire [1-1:0] node2682;
	wire [1-1:0] node2685;
	wire [1-1:0] node2686;
	wire [1-1:0] node2687;
	wire [1-1:0] node2691;
	wire [1-1:0] node2693;
	wire [1-1:0] node2697;
	wire [1-1:0] node2698;
	wire [1-1:0] node2700;
	wire [1-1:0] node2701;
	wire [1-1:0] node2702;
	wire [1-1:0] node2704;
	wire [1-1:0] node2707;
	wire [1-1:0] node2708;
	wire [1-1:0] node2711;
	wire [1-1:0] node2712;
	wire [1-1:0] node2715;
	wire [1-1:0] node2719;
	wire [1-1:0] node2720;
	wire [1-1:0] node2721;
	wire [1-1:0] node2722;
	wire [1-1:0] node2723;
	wire [1-1:0] node2724;
	wire [1-1:0] node2728;
	wire [1-1:0] node2729;
	wire [1-1:0] node2730;
	wire [1-1:0] node2734;
	wire [1-1:0] node2735;
	wire [1-1:0] node2740;
	wire [1-1:0] node2741;
	wire [1-1:0] node2742;
	wire [1-1:0] node2744;
	wire [1-1:0] node2747;
	wire [1-1:0] node2749;
	wire [1-1:0] node2752;
	wire [1-1:0] node2754;
	wire [1-1:0] node2757;
	wire [1-1:0] node2758;
	wire [1-1:0] node2760;
	wire [1-1:0] node2761;
	wire [1-1:0] node2762;
	wire [1-1:0] node2766;
	wire [1-1:0] node2767;
	wire [1-1:0] node2769;
	wire [1-1:0] node2772;
	wire [1-1:0] node2774;
	wire [1-1:0] node2778;
	wire [1-1:0] node2779;
	wire [1-1:0] node2780;
	wire [1-1:0] node2781;
	wire [1-1:0] node2783;
	wire [1-1:0] node2784;
	wire [1-1:0] node2786;
	wire [1-1:0] node2789;
	wire [1-1:0] node2790;
	wire [1-1:0] node2791;
	wire [1-1:0] node2795;
	wire [1-1:0] node2796;
	wire [1-1:0] node2801;
	wire [1-1:0] node2802;
	wire [1-1:0] node2803;
	wire [1-1:0] node2805;
	wire [1-1:0] node2808;
	wire [1-1:0] node2809;
	wire [1-1:0] node2811;
	wire [1-1:0] node2814;
	wire [1-1:0] node2816;
	wire [1-1:0] node2819;
	wire [1-1:0] node2821;
	wire [1-1:0] node2822;
	wire [1-1:0] node2823;
	wire [1-1:0] node2825;
	wire [1-1:0] node2828;
	wire [1-1:0] node2829;
	wire [1-1:0] node2833;
	wire [1-1:0] node2834;
	wire [1-1:0] node2838;
	wire [1-1:0] node2839;
	wire [1-1:0] node2841;
	wire [1-1:0] node2842;
	wire [1-1:0] node2844;
	wire [1-1:0] node2847;
	wire [1-1:0] node2848;
	wire [1-1:0] node2849;
	wire [1-1:0] node2853;
	wire [1-1:0] node2854;

	assign outp = (inp[4]) ? node2032 : node1;
		assign node1 = (inp[0]) ? node733 : node2;
			assign node2 = (inp[8]) ? node652 : node3;
				assign node3 = (inp[1]) ? node85 : node4;
					assign node4 = (inp[6]) ? node26 : node5;
						assign node5 = (inp[15]) ? 1'b1 : node6;
							assign node6 = (inp[12]) ? node8 : 1'b1;
								assign node8 = (inp[3]) ? node14 : node9;
									assign node9 = (inp[9]) ? node11 : 1'b0;
										assign node11 = (inp[10]) ? 1'b0 : 1'b1;
									assign node14 = (inp[7]) ? node20 : node15;
										assign node15 = (inp[9]) ? node17 : 1'b1;
											assign node17 = (inp[10]) ? 1'b1 : 1'b0;
										assign node20 = (inp[10]) ? 1'b0 : node21;
											assign node21 = (inp[9]) ? 1'b1 : 1'b0;
						assign node26 = (inp[5]) ? node64 : node27;
							assign node27 = (inp[12]) ? node45 : node28;
								assign node28 = (inp[7]) ? node40 : node29;
									assign node29 = (inp[3]) ? node35 : node30;
										assign node30 = (inp[10]) ? 1'b0 : node31;
											assign node31 = (inp[9]) ? 1'b1 : 1'b0;
										assign node35 = (inp[10]) ? 1'b1 : node36;
											assign node36 = (inp[9]) ? 1'b0 : 1'b1;
									assign node40 = (inp[10]) ? 1'b0 : node41;
										assign node41 = (inp[9]) ? 1'b1 : 1'b0;
								assign node45 = (inp[15]) ? node47 : 1'b1;
									assign node47 = (inp[9]) ? node53 : node48;
										assign node48 = (inp[3]) ? node50 : 1'b0;
											assign node50 = (inp[7]) ? 1'b0 : 1'b1;
										assign node53 = (inp[10]) ? node59 : node54;
											assign node54 = (inp[7]) ? 1'b1 : node55;
												assign node55 = (inp[3]) ? 1'b0 : 1'b1;
											assign node59 = (inp[3]) ? node61 : 1'b0;
												assign node61 = (inp[7]) ? 1'b0 : 1'b1;
							assign node64 = (inp[15]) ? 1'b1 : node65;
								assign node65 = (inp[12]) ? node67 : 1'b1;
									assign node67 = (inp[7]) ? node79 : node68;
										assign node68 = (inp[3]) ? node74 : node69;
											assign node69 = (inp[9]) ? node71 : 1'b0;
												assign node71 = (inp[10]) ? 1'b0 : 1'b1;
											assign node74 = (inp[10]) ? 1'b1 : node75;
												assign node75 = (inp[9]) ? 1'b0 : 1'b1;
										assign node79 = (inp[10]) ? 1'b0 : node80;
											assign node80 = (inp[9]) ? 1'b1 : 1'b0;
					assign node85 = (inp[11]) ? node411 : node86;
						assign node86 = (inp[13]) ? node248 : node87;
							assign node87 = (inp[2]) ? node175 : node88;
								assign node88 = (inp[14]) ? node130 : node89;
									assign node89 = (inp[6]) ? node103 : node90;
										assign node90 = (inp[12]) ? node92 : 1'b0;
											assign node92 = (inp[15]) ? 1'b0 : node93;
												assign node93 = (inp[3]) ? node99 : node94;
													assign node94 = (inp[10]) ? 1'b1 : node95;
														assign node95 = (inp[9]) ? 1'b0 : 1'b1;
													assign node99 = (inp[10]) ? 1'b0 : 1'b1;
										assign node103 = (inp[5]) ? node121 : node104;
											assign node104 = (inp[15]) ? node114 : node105;
												assign node105 = (inp[12]) ? 1'b0 : node106;
													assign node106 = (inp[7]) ? node108 : 1'b0;
														assign node108 = (inp[3]) ? 1'b1 : node109;
															assign node109 = (inp[9]) ? 1'b0 : 1'b1;
												assign node114 = (inp[3]) ? node116 : 1'b1;
													assign node116 = (inp[10]) ? 1'b1 : node117;
														assign node117 = (inp[7]) ? 1'b0 : 1'b1;
											assign node121 = (inp[15]) ? 1'b0 : node122;
												assign node122 = (inp[12]) ? node124 : 1'b0;
													assign node124 = (inp[9]) ? node126 : 1'b1;
														assign node126 = (inp[10]) ? 1'b1 : 1'b0;
									assign node130 = (inp[6]) ? node138 : node131;
										assign node131 = (inp[12]) ? node133 : 1'b1;
											assign node133 = (inp[7]) ? node135 : 1'b1;
												assign node135 = (inp[15]) ? 1'b1 : 1'b0;
										assign node138 = (inp[10]) ? node154 : node139;
											assign node139 = (inp[15]) ? 1'b1 : node140;
												assign node140 = (inp[9]) ? node148 : node141;
													assign node141 = (inp[7]) ? node143 : 1'b1;
														assign node143 = (inp[5]) ? node145 : 1'b0;
															assign node145 = (inp[3]) ? 1'b0 : 1'b1;
													assign node148 = (inp[5]) ? node150 : 1'b1;
														assign node150 = (inp[7]) ? 1'b1 : 1'b0;
											assign node154 = (inp[3]) ? node164 : node155;
												assign node155 = (inp[15]) ? node161 : node156;
													assign node156 = (inp[5]) ? node158 : 1'b1;
														assign node158 = (inp[12]) ? 1'b0 : 1'b1;
													assign node161 = (inp[5]) ? 1'b1 : 1'b0;
												assign node164 = (inp[7]) ? node166 : 1'b1;
													assign node166 = (inp[9]) ? node168 : 1'b0;
														assign node168 = (inp[5]) ? node172 : node169;
															assign node169 = (inp[12]) ? 1'b1 : 1'b0;
															assign node172 = (inp[12]) ? 1'b0 : 1'b1;
								assign node175 = (inp[12]) ? node197 : node176;
									assign node176 = (inp[5]) ? 1'b0 : node177;
										assign node177 = (inp[6]) ? node179 : 1'b0;
											assign node179 = (inp[15]) ? node181 : 1'b1;
												assign node181 = (inp[10]) ? node193 : node182;
													assign node182 = (inp[9]) ? node188 : node183;
														assign node183 = (inp[3]) ? node185 : 1'b1;
															assign node185 = (inp[14]) ? 1'b0 : 1'b1;
														assign node188 = (inp[3]) ? node190 : 1'b0;
															assign node190 = (inp[7]) ? 1'b0 : 1'b1;
													assign node193 = (inp[3]) ? 1'b0 : 1'b1;
									assign node197 = (inp[15]) ? node231 : node198;
										assign node198 = (inp[5]) ? node214 : node199;
											assign node199 = (inp[6]) ? 1'b0 : node200;
												assign node200 = (inp[7]) ? 1'b1 : node201;
													assign node201 = (inp[14]) ? 1'b0 : node202;
														assign node202 = (inp[9]) ? node204 : 1'b0;
															assign node204 = (inp[3]) ? node208 : node205;
																assign node205 = (inp[10]) ? 1'b1 : 1'b0;
																assign node208 = (inp[10]) ? 1'b0 : 1'b1;
											assign node214 = (inp[3]) ? node220 : node215;
												assign node215 = (inp[10]) ? 1'b1 : node216;
													assign node216 = (inp[9]) ? 1'b0 : 1'b1;
												assign node220 = (inp[10]) ? node228 : node221;
													assign node221 = (inp[14]) ? 1'b1 : node222;
														assign node222 = (inp[7]) ? 1'b0 : node223;
															assign node223 = (inp[9]) ? 1'b1 : 1'b0;
													assign node228 = (inp[7]) ? 1'b1 : 1'b0;
										assign node231 = (inp[5]) ? 1'b0 : node232;
											assign node232 = (inp[6]) ? node234 : 1'b0;
												assign node234 = (inp[14]) ? node242 : node235;
													assign node235 = (inp[10]) ? 1'b1 : node236;
														assign node236 = (inp[7]) ? 1'b1 : node237;
															assign node237 = (inp[3]) ? 1'b1 : 1'b0;
													assign node242 = (inp[3]) ? 1'b0 : node243;
														assign node243 = (inp[9]) ? 1'b0 : 1'b1;
							assign node248 = (inp[2]) ? node350 : node249;
								assign node249 = (inp[14]) ? node285 : node250;
									assign node250 = (inp[12]) ? node260 : node251;
										assign node251 = (inp[5]) ? 1'b1 : node252;
											assign node252 = (inp[6]) ? node254 : 1'b1;
												assign node254 = (inp[7]) ? 1'b0 : node255;
													assign node255 = (inp[9]) ? 1'b0 : 1'b1;
										assign node260 = (inp[15]) ? node276 : node261;
											assign node261 = (inp[10]) ? node267 : node262;
												assign node262 = (inp[9]) ? 1'b1 : node263;
													assign node263 = (inp[7]) ? 1'b0 : 1'b1;
												assign node267 = (inp[6]) ? node269 : 1'b0;
													assign node269 = (inp[5]) ? node271 : 1'b1;
														assign node271 = (inp[3]) ? node273 : 1'b0;
															assign node273 = (inp[7]) ? 1'b0 : 1'b1;
											assign node276 = (inp[6]) ? node278 : 1'b1;
												assign node278 = (inp[5]) ? 1'b1 : node279;
													assign node279 = (inp[7]) ? 1'b0 : node280;
														assign node280 = (inp[10]) ? 1'b0 : 1'b1;
									assign node285 = (inp[7]) ? node321 : node286;
										assign node286 = (inp[3]) ? node306 : node287;
											assign node287 = (inp[10]) ? node293 : node288;
												assign node288 = (inp[9]) ? 1'b0 : node289;
													assign node289 = (inp[12]) ? 1'b1 : 1'b0;
												assign node293 = (inp[9]) ? node299 : node294;
													assign node294 = (inp[6]) ? node296 : 1'b0;
														assign node296 = (inp[5]) ? 1'b0 : 1'b1;
													assign node299 = (inp[12]) ? 1'b1 : node300;
														assign node300 = (inp[15]) ? node302 : 1'b0;
															assign node302 = (inp[6]) ? 1'b1 : 1'b0;
											assign node306 = (inp[10]) ? 1'b0 : node307;
												assign node307 = (inp[9]) ? node309 : 1'b0;
													assign node309 = (inp[6]) ? node311 : 1'b0;
														assign node311 = (inp[15]) ? node317 : node312;
															assign node312 = (inp[5]) ? node314 : 1'b0;
																assign node314 = (inp[12]) ? 1'b1 : 1'b0;
															assign node317 = (inp[5]) ? 1'b0 : 1'b1;
										assign node321 = (inp[12]) ? node331 : node322;
											assign node322 = (inp[5]) ? 1'b0 : node323;
												assign node323 = (inp[6]) ? node325 : 1'b0;
													assign node325 = (inp[9]) ? node327 : 1'b1;
														assign node327 = (inp[10]) ? 1'b1 : 1'b0;
											assign node331 = (inp[3]) ? node339 : node332;
												assign node332 = (inp[15]) ? node334 : 1'b1;
													assign node334 = (inp[5]) ? 1'b0 : node335;
														assign node335 = (inp[6]) ? 1'b1 : 1'b0;
												assign node339 = (inp[9]) ? 1'b0 : node340;
													assign node340 = (inp[5]) ? node346 : node341;
														assign node341 = (inp[15]) ? node343 : 1'b0;
															assign node343 = (inp[6]) ? 1'b1 : 1'b0;
														assign node346 = (inp[15]) ? 1'b0 : 1'b1;
								assign node350 = (inp[15]) ? node394 : node351;
									assign node351 = (inp[12]) ? node369 : node352;
										assign node352 = (inp[6]) ? node354 : 1'b1;
											assign node354 = (inp[5]) ? 1'b1 : node355;
												assign node355 = (inp[10]) ? 1'b0 : node356;
													assign node356 = (inp[9]) ? node362 : node357;
														assign node357 = (inp[7]) ? 1'b0 : node358;
															assign node358 = (inp[3]) ? 1'b1 : 1'b0;
														assign node362 = (inp[14]) ? node364 : 1'b1;
															assign node364 = (inp[7]) ? 1'b1 : 1'b0;
										assign node369 = (inp[3]) ? node381 : node370;
											assign node370 = (inp[6]) ? node378 : node371;
												assign node371 = (inp[5]) ? node373 : 1'b0;
													assign node373 = (inp[9]) ? node375 : 1'b0;
														assign node375 = (inp[10]) ? 1'b0 : 1'b1;
												assign node378 = (inp[5]) ? 1'b0 : 1'b1;
											assign node381 = (inp[5]) ? node387 : node382;
												assign node382 = (inp[6]) ? 1'b1 : node383;
													assign node383 = (inp[9]) ? 1'b1 : 1'b0;
												assign node387 = (inp[10]) ? node391 : node388;
													assign node388 = (inp[7]) ? 1'b1 : 1'b0;
													assign node391 = (inp[7]) ? 1'b0 : 1'b1;
									assign node394 = (inp[5]) ? 1'b1 : node395;
										assign node395 = (inp[6]) ? node397 : 1'b1;
											assign node397 = (inp[9]) ? node403 : node398;
												assign node398 = (inp[3]) ? node400 : 1'b0;
													assign node400 = (inp[7]) ? 1'b0 : 1'b1;
												assign node403 = (inp[10]) ? 1'b0 : node404;
													assign node404 = (inp[7]) ? 1'b1 : node405;
														assign node405 = (inp[12]) ? 1'b0 : 1'b1;
						assign node411 = (inp[2]) ? node561 : node412;
							assign node412 = (inp[14]) ? node490 : node413;
								assign node413 = (inp[6]) ? node433 : node414;
									assign node414 = (inp[12]) ? node416 : 1'b0;
										assign node416 = (inp[15]) ? 1'b0 : node417;
											assign node417 = (inp[7]) ? node427 : node418;
												assign node418 = (inp[10]) ? 1'b0 : node419;
													assign node419 = (inp[9]) ? node423 : node420;
														assign node420 = (inp[3]) ? 1'b0 : 1'b1;
														assign node423 = (inp[3]) ? 1'b1 : 1'b0;
												assign node427 = (inp[10]) ? 1'b1 : node428;
													assign node428 = (inp[9]) ? 1'b0 : 1'b1;
									assign node433 = (inp[5]) ? node477 : node434;
										assign node434 = (inp[12]) ? node454 : node435;
											assign node435 = (inp[9]) ? node441 : node436;
												assign node436 = (inp[7]) ? 1'b1 : node437;
													assign node437 = (inp[3]) ? 1'b0 : 1'b1;
												assign node441 = (inp[15]) ? node447 : node442;
													assign node442 = (inp[10]) ? 1'b1 : node443;
														assign node443 = (inp[3]) ? 1'b1 : 1'b0;
													assign node447 = (inp[3]) ? node451 : node448;
														assign node448 = (inp[10]) ? 1'b1 : 1'b0;
														assign node451 = (inp[10]) ? 1'b0 : 1'b1;
											assign node454 = (inp[15]) ? node456 : 1'b0;
												assign node456 = (inp[7]) ? node472 : node457;
													assign node457 = (inp[9]) ? node461 : node458;
														assign node458 = (inp[3]) ? 1'b0 : 1'b1;
														assign node461 = (inp[13]) ? node467 : node462;
															assign node462 = (inp[10]) ? 1'b0 : node463;
																assign node463 = (inp[3]) ? 1'b1 : 1'b0;
															assign node467 = (inp[3]) ? 1'b1 : node468;
																assign node468 = (inp[10]) ? 1'b1 : 1'b0;
													assign node472 = (inp[9]) ? node474 : 1'b1;
														assign node474 = (inp[10]) ? 1'b1 : 1'b0;
										assign node477 = (inp[12]) ? node479 : 1'b0;
											assign node479 = (inp[15]) ? 1'b0 : node480;
												assign node480 = (inp[13]) ? node482 : 1'b1;
													assign node482 = (inp[3]) ? node486 : node483;
														assign node483 = (inp[7]) ? 1'b0 : 1'b1;
														assign node486 = (inp[7]) ? 1'b1 : 1'b0;
								assign node490 = (inp[6]) ? node510 : node491;
									assign node491 = (inp[12]) ? node493 : 1'b1;
										assign node493 = (inp[15]) ? 1'b1 : node494;
											assign node494 = (inp[3]) ? node500 : node495;
												assign node495 = (inp[7]) ? 1'b0 : node496;
													assign node496 = (inp[9]) ? 1'b1 : 1'b0;
												assign node500 = (inp[10]) ? node506 : node501;
													assign node501 = (inp[7]) ? node503 : 1'b0;
														assign node503 = (inp[9]) ? 1'b1 : 1'b0;
													assign node506 = (inp[7]) ? 1'b0 : 1'b1;
									assign node510 = (inp[5]) ? node550 : node511;
										assign node511 = (inp[12]) ? node531 : node512;
											assign node512 = (inp[3]) ? node518 : node513;
												assign node513 = (inp[9]) ? node515 : 1'b0;
													assign node515 = (inp[10]) ? 1'b0 : 1'b1;
												assign node518 = (inp[15]) ? node524 : node519;
													assign node519 = (inp[10]) ? node521 : 1'b0;
														assign node521 = (inp[13]) ? 1'b0 : 1'b1;
													assign node524 = (inp[9]) ? node526 : 1'b1;
														assign node526 = (inp[7]) ? 1'b1 : node527;
															assign node527 = (inp[10]) ? 1'b1 : 1'b0;
											assign node531 = (inp[15]) ? node533 : 1'b1;
												assign node533 = (inp[10]) ? 1'b0 : node534;
													assign node534 = (inp[13]) ? node540 : node535;
														assign node535 = (inp[3]) ? node537 : 1'b0;
															assign node537 = (inp[7]) ? 1'b0 : 1'b1;
														assign node540 = (inp[3]) ? node542 : 1'b1;
															assign node542 = (inp[9]) ? node546 : node543;
																assign node543 = (inp[7]) ? 1'b0 : 1'b1;
																assign node546 = (inp[7]) ? 1'b1 : 1'b0;
										assign node550 = (inp[12]) ? node552 : 1'b1;
											assign node552 = (inp[15]) ? 1'b1 : node553;
												assign node553 = (inp[7]) ? node555 : 1'b1;
													assign node555 = (inp[10]) ? 1'b0 : node556;
														assign node556 = (inp[3]) ? 1'b0 : 1'b1;
							assign node561 = (inp[5]) ? node617 : node562;
								assign node562 = (inp[6]) ? node582 : node563;
									assign node563 = (inp[15]) ? 1'b0 : node564;
										assign node564 = (inp[12]) ? node566 : 1'b0;
											assign node566 = (inp[3]) ? node572 : node567;
												assign node567 = (inp[9]) ? node569 : 1'b1;
													assign node569 = (inp[10]) ? 1'b1 : 1'b0;
												assign node572 = (inp[9]) ? node574 : 1'b0;
													assign node574 = (inp[14]) ? node576 : 1'b1;
														assign node576 = (inp[10]) ? 1'b0 : node577;
															assign node577 = (inp[7]) ? 1'b0 : 1'b1;
									assign node582 = (inp[15]) ? node600 : node583;
										assign node583 = (inp[12]) ? 1'b0 : node584;
											assign node584 = (inp[9]) ? node590 : node585;
												assign node585 = (inp[10]) ? node587 : 1'b1;
													assign node587 = (inp[14]) ? 1'b1 : 1'b0;
												assign node590 = (inp[10]) ? node596 : node591;
													assign node591 = (inp[3]) ? node593 : 1'b0;
														assign node593 = (inp[7]) ? 1'b0 : 1'b1;
													assign node596 = (inp[7]) ? 1'b1 : 1'b0;
										assign node600 = (inp[3]) ? node606 : node601;
											assign node601 = (inp[9]) ? node603 : 1'b1;
												assign node603 = (inp[10]) ? 1'b1 : 1'b0;
											assign node606 = (inp[7]) ? node612 : node607;
												assign node607 = (inp[10]) ? 1'b0 : node608;
													assign node608 = (inp[9]) ? 1'b1 : 1'b0;
												assign node612 = (inp[9]) ? node614 : 1'b1;
													assign node614 = (inp[10]) ? 1'b1 : 1'b0;
								assign node617 = (inp[15]) ? 1'b0 : node618;
									assign node618 = (inp[12]) ? node620 : 1'b0;
										assign node620 = (inp[9]) ? node626 : node621;
											assign node621 = (inp[7]) ? 1'b1 : node622;
												assign node622 = (inp[3]) ? 1'b0 : 1'b1;
											assign node626 = (inp[6]) ? node640 : node627;
												assign node627 = (inp[13]) ? node633 : node628;
													assign node628 = (inp[3]) ? node630 : 1'b1;
														assign node630 = (inp[14]) ? 1'b1 : 1'b0;
													assign node633 = (inp[14]) ? 1'b0 : node634;
														assign node634 = (inp[7]) ? 1'b1 : node635;
															assign node635 = (inp[10]) ? 1'b0 : 1'b1;
												assign node640 = (inp[10]) ? node648 : node641;
													assign node641 = (inp[13]) ? node643 : 1'b0;
														assign node643 = (inp[3]) ? node645 : 1'b0;
															assign node645 = (inp[7]) ? 1'b0 : 1'b1;
													assign node648 = (inp[3]) ? 1'b0 : 1'b1;
				assign node652 = (inp[15]) ? node712 : node653;
					assign node653 = (inp[12]) ? node675 : node654;
						assign node654 = (inp[5]) ? 1'b1 : node655;
							assign node655 = (inp[6]) ? node657 : 1'b1;
								assign node657 = (inp[9]) ? node663 : node658;
									assign node658 = (inp[7]) ? 1'b0 : node659;
										assign node659 = (inp[3]) ? 1'b1 : 1'b0;
									assign node663 = (inp[10]) ? node669 : node664;
										assign node664 = (inp[7]) ? 1'b1 : node665;
											assign node665 = (inp[3]) ? 1'b0 : 1'b1;
										assign node669 = (inp[7]) ? 1'b0 : node670;
											assign node670 = (inp[3]) ? 1'b1 : 1'b0;
						assign node675 = (inp[5]) ? node695 : node676;
							assign node676 = (inp[6]) ? 1'b1 : node677;
								assign node677 = (inp[3]) ? node683 : node678;
									assign node678 = (inp[9]) ? node680 : 1'b0;
										assign node680 = (inp[10]) ? 1'b0 : 1'b1;
									assign node683 = (inp[7]) ? node689 : node684;
										assign node684 = (inp[10]) ? 1'b1 : node685;
											assign node685 = (inp[9]) ? 1'b0 : 1'b1;
										assign node689 = (inp[10]) ? 1'b0 : node690;
											assign node690 = (inp[9]) ? 1'b1 : 1'b0;
							assign node695 = (inp[9]) ? node701 : node696;
								assign node696 = (inp[3]) ? node698 : 1'b0;
									assign node698 = (inp[7]) ? 1'b0 : 1'b1;
								assign node701 = (inp[10]) ? node707 : node702;
									assign node702 = (inp[3]) ? node704 : 1'b1;
										assign node704 = (inp[7]) ? 1'b1 : 1'b0;
									assign node707 = (inp[7]) ? 1'b0 : node708;
										assign node708 = (inp[3]) ? 1'b1 : 1'b0;
					assign node712 = (inp[5]) ? 1'b1 : node713;
						assign node713 = (inp[6]) ? node715 : 1'b1;
							assign node715 = (inp[10]) ? node727 : node716;
								assign node716 = (inp[9]) ? node722 : node717;
									assign node717 = (inp[7]) ? 1'b0 : node718;
										assign node718 = (inp[3]) ? 1'b1 : 1'b0;
									assign node722 = (inp[7]) ? 1'b1 : node723;
										assign node723 = (inp[3]) ? 1'b0 : 1'b1;
								assign node727 = (inp[7]) ? 1'b0 : node728;
									assign node728 = (inp[3]) ? 1'b1 : 1'b0;
			assign node733 = (inp[8]) ? node1355 : node734;
				assign node734 = (inp[1]) ? node1274 : node735;
					assign node735 = (inp[11]) ? node1033 : node736;
						assign node736 = (inp[13]) ? node878 : node737;
							assign node737 = (inp[2]) ? node821 : node738;
								assign node738 = (inp[14]) ? node774 : node739;
									assign node739 = (inp[12]) ? node751 : node740;
										assign node740 = (inp[5]) ? 1'b0 : node741;
											assign node741 = (inp[6]) ? node743 : 1'b0;
												assign node743 = (inp[10]) ? 1'b1 : node744;
													assign node744 = (inp[9]) ? 1'b0 : node745;
														assign node745 = (inp[3]) ? 1'b0 : 1'b1;
										assign node751 = (inp[15]) ? node763 : node752;
											assign node752 = (inp[5]) ? node756 : node753;
												assign node753 = (inp[6]) ? 1'b0 : 1'b1;
												assign node756 = (inp[10]) ? 1'b1 : node757;
													assign node757 = (inp[9]) ? node759 : 1'b1;
														assign node759 = (inp[7]) ? 1'b0 : 1'b1;
											assign node763 = (inp[10]) ? node765 : 1'b0;
												assign node765 = (inp[5]) ? 1'b0 : node766;
													assign node766 = (inp[6]) ? node768 : 1'b0;
														assign node768 = (inp[7]) ? 1'b1 : node769;
															assign node769 = (inp[9]) ? 1'b0 : 1'b1;
									assign node774 = (inp[3]) ? node798 : node775;
										assign node775 = (inp[6]) ? node783 : node776;
											assign node776 = (inp[15]) ? 1'b1 : node777;
												assign node777 = (inp[12]) ? node779 : 1'b1;
													assign node779 = (inp[10]) ? 1'b0 : 1'b1;
											assign node783 = (inp[5]) ? node791 : node784;
												assign node784 = (inp[15]) ? 1'b0 : node785;
													assign node785 = (inp[10]) ? 1'b1 : node786;
														assign node786 = (inp[7]) ? 1'b0 : 1'b1;
												assign node791 = (inp[15]) ? 1'b1 : node792;
													assign node792 = (inp[7]) ? node794 : 1'b1;
														assign node794 = (inp[9]) ? 1'b1 : 1'b0;
										assign node798 = (inp[5]) ? node812 : node799;
											assign node799 = (inp[10]) ? 1'b1 : node800;
												assign node800 = (inp[9]) ? node804 : node801;
													assign node801 = (inp[7]) ? 1'b0 : 1'b1;
													assign node804 = (inp[7]) ? 1'b1 : node805;
														assign node805 = (inp[15]) ? node807 : 1'b0;
															assign node807 = (inp[12]) ? 1'b1 : 1'b0;
											assign node812 = (inp[15]) ? 1'b1 : node813;
												assign node813 = (inp[9]) ? 1'b1 : node814;
													assign node814 = (inp[7]) ? node816 : 1'b1;
														assign node816 = (inp[12]) ? 1'b0 : 1'b1;
								assign node821 = (inp[5]) ? node865 : node822;
									assign node822 = (inp[6]) ? node836 : node823;
										assign node823 = (inp[15]) ? 1'b0 : node824;
											assign node824 = (inp[12]) ? node826 : 1'b0;
												assign node826 = (inp[14]) ? node828 : 1'b1;
													assign node828 = (inp[7]) ? 1'b1 : node829;
														assign node829 = (inp[3]) ? 1'b0 : node830;
															assign node830 = (inp[9]) ? 1'b0 : 1'b1;
										assign node836 = (inp[9]) ? node850 : node837;
											assign node837 = (inp[15]) ? node845 : node838;
												assign node838 = (inp[12]) ? 1'b0 : node839;
													assign node839 = (inp[3]) ? node841 : 1'b1;
														assign node841 = (inp[7]) ? 1'b1 : 1'b0;
												assign node845 = (inp[7]) ? 1'b1 : node846;
													assign node846 = (inp[3]) ? 1'b0 : 1'b1;
											assign node850 = (inp[10]) ? node858 : node851;
												assign node851 = (inp[3]) ? node853 : 1'b0;
													assign node853 = (inp[7]) ? 1'b0 : node854;
														assign node854 = (inp[15]) ? 1'b1 : 1'b0;
												assign node858 = (inp[15]) ? 1'b1 : node859;
													assign node859 = (inp[3]) ? 1'b0 : node860;
														assign node860 = (inp[12]) ? 1'b0 : 1'b1;
									assign node865 = (inp[15]) ? 1'b0 : node866;
										assign node866 = (inp[12]) ? node868 : 1'b0;
											assign node868 = (inp[7]) ? 1'b1 : node869;
												assign node869 = (inp[3]) ? 1'b0 : node870;
													assign node870 = (inp[6]) ? 1'b1 : node871;
														assign node871 = (inp[9]) ? 1'b0 : 1'b1;
							assign node878 = (inp[14]) ? node950 : node879;
								assign node879 = (inp[5]) ? node933 : node880;
									assign node880 = (inp[6]) ? node900 : node881;
										assign node881 = (inp[15]) ? 1'b1 : node882;
											assign node882 = (inp[12]) ? node884 : 1'b1;
												assign node884 = (inp[10]) ? node894 : node885;
													assign node885 = (inp[3]) ? node889 : node886;
														assign node886 = (inp[9]) ? 1'b1 : 1'b0;
														assign node889 = (inp[2]) ? 1'b0 : node890;
															assign node890 = (inp[7]) ? 1'b0 : 1'b1;
													assign node894 = (inp[3]) ? node896 : 1'b0;
														assign node896 = (inp[7]) ? 1'b0 : 1'b1;
										assign node900 = (inp[7]) ? node920 : node901;
											assign node901 = (inp[15]) ? node909 : node902;
												assign node902 = (inp[12]) ? 1'b1 : node903;
													assign node903 = (inp[3]) ? node905 : 1'b1;
														assign node905 = (inp[10]) ? 1'b1 : 1'b0;
												assign node909 = (inp[10]) ? node917 : node910;
													assign node910 = (inp[3]) ? node914 : node911;
														assign node911 = (inp[9]) ? 1'b1 : 1'b0;
														assign node914 = (inp[9]) ? 1'b0 : 1'b1;
													assign node917 = (inp[3]) ? 1'b1 : 1'b0;
											assign node920 = (inp[12]) ? node926 : node921;
												assign node921 = (inp[9]) ? node923 : 1'b0;
													assign node923 = (inp[10]) ? 1'b0 : 1'b1;
												assign node926 = (inp[15]) ? node928 : 1'b1;
													assign node928 = (inp[10]) ? 1'b0 : node929;
														assign node929 = (inp[2]) ? 1'b0 : 1'b1;
									assign node933 = (inp[12]) ? node935 : 1'b1;
										assign node935 = (inp[15]) ? 1'b1 : node936;
											assign node936 = (inp[10]) ? node944 : node937;
												assign node937 = (inp[9]) ? 1'b1 : node938;
													assign node938 = (inp[3]) ? node940 : 1'b0;
														assign node940 = (inp[7]) ? 1'b0 : 1'b1;
												assign node944 = (inp[3]) ? node946 : 1'b0;
													assign node946 = (inp[7]) ? 1'b0 : 1'b1;
								assign node950 = (inp[2]) ? node992 : node951;
									assign node951 = (inp[9]) ? node977 : node952;
										assign node952 = (inp[15]) ? node968 : node953;
											assign node953 = (inp[3]) ? node959 : node954;
												assign node954 = (inp[12]) ? 1'b1 : node955;
													assign node955 = (inp[5]) ? 1'b0 : 1'b1;
												assign node959 = (inp[7]) ? node961 : 1'b0;
													assign node961 = (inp[12]) ? 1'b1 : node962;
														assign node962 = (inp[6]) ? node964 : 1'b0;
															assign node964 = (inp[5]) ? 1'b0 : 1'b1;
											assign node968 = (inp[6]) ? node970 : 1'b0;
												assign node970 = (inp[5]) ? 1'b0 : node971;
													assign node971 = (inp[3]) ? node973 : 1'b1;
														assign node973 = (inp[7]) ? 1'b1 : 1'b0;
										assign node977 = (inp[12]) ? node979 : 1'b0;
											assign node979 = (inp[10]) ? node987 : node980;
												assign node980 = (inp[15]) ? 1'b0 : node981;
													assign node981 = (inp[6]) ? node983 : 1'b0;
														assign node983 = (inp[3]) ? 1'b1 : 1'b0;
												assign node987 = (inp[7]) ? 1'b1 : node988;
													assign node988 = (inp[6]) ? 1'b1 : 1'b0;
									assign node992 = (inp[3]) ? node1018 : node993;
										assign node993 = (inp[6]) ? node1003 : node994;
											assign node994 = (inp[12]) ? node996 : 1'b1;
												assign node996 = (inp[15]) ? 1'b1 : node997;
													assign node997 = (inp[10]) ? 1'b0 : node998;
														assign node998 = (inp[7]) ? 1'b0 : 1'b1;
											assign node1003 = (inp[9]) ? node1009 : node1004;
												assign node1004 = (inp[5]) ? node1006 : 1'b0;
													assign node1006 = (inp[15]) ? 1'b1 : 1'b0;
												assign node1009 = (inp[10]) ? node1011 : 1'b1;
													assign node1011 = (inp[5]) ? 1'b1 : node1012;
														assign node1012 = (inp[7]) ? 1'b0 : node1013;
															assign node1013 = (inp[12]) ? 1'b1 : 1'b0;
										assign node1018 = (inp[5]) ? node1026 : node1019;
											assign node1019 = (inp[9]) ? 1'b1 : node1020;
												assign node1020 = (inp[6]) ? node1022 : 1'b1;
													assign node1022 = (inp[7]) ? 1'b0 : 1'b1;
											assign node1026 = (inp[12]) ? node1028 : 1'b1;
												assign node1028 = (inp[15]) ? 1'b1 : node1029;
													assign node1029 = (inp[10]) ? 1'b1 : 1'b0;
						assign node1033 = (inp[14]) ? node1123 : node1034;
							assign node1034 = (inp[6]) ? node1062 : node1035;
								assign node1035 = (inp[15]) ? 1'b0 : node1036;
									assign node1036 = (inp[12]) ? node1038 : 1'b0;
										assign node1038 = (inp[3]) ? node1044 : node1039;
											assign node1039 = (inp[9]) ? node1041 : 1'b1;
												assign node1041 = (inp[10]) ? 1'b1 : 1'b0;
											assign node1044 = (inp[13]) ? node1054 : node1045;
												assign node1045 = (inp[2]) ? node1047 : 1'b1;
													assign node1047 = (inp[10]) ? 1'b0 : node1048;
														assign node1048 = (inp[7]) ? node1050 : 1'b1;
															assign node1050 = (inp[5]) ? 1'b0 : 1'b1;
												assign node1054 = (inp[7]) ? node1056 : 1'b0;
													assign node1056 = (inp[10]) ? 1'b1 : node1057;
														assign node1057 = (inp[9]) ? 1'b0 : 1'b1;
								assign node1062 = (inp[5]) ? node1098 : node1063;
									assign node1063 = (inp[10]) ? node1085 : node1064;
										assign node1064 = (inp[9]) ? node1076 : node1065;
											assign node1065 = (inp[7]) ? node1071 : node1066;
												assign node1066 = (inp[3]) ? 1'b0 : node1067;
													assign node1067 = (inp[15]) ? 1'b1 : 1'b0;
												assign node1071 = (inp[12]) ? node1073 : 1'b1;
													assign node1073 = (inp[15]) ? 1'b1 : 1'b0;
											assign node1076 = (inp[15]) ? node1078 : 1'b0;
												assign node1078 = (inp[13]) ? 1'b0 : node1079;
													assign node1079 = (inp[7]) ? 1'b0 : node1080;
														assign node1080 = (inp[3]) ? 1'b1 : 1'b0;
										assign node1085 = (inp[7]) ? node1093 : node1086;
											assign node1086 = (inp[3]) ? 1'b0 : node1087;
												assign node1087 = (inp[12]) ? node1089 : 1'b1;
													assign node1089 = (inp[15]) ? 1'b1 : 1'b0;
											assign node1093 = (inp[15]) ? 1'b1 : node1094;
												assign node1094 = (inp[12]) ? 1'b0 : 1'b1;
									assign node1098 = (inp[15]) ? 1'b0 : node1099;
										assign node1099 = (inp[12]) ? node1101 : 1'b0;
											assign node1101 = (inp[3]) ? node1107 : node1102;
												assign node1102 = (inp[9]) ? node1104 : 1'b1;
													assign node1104 = (inp[10]) ? 1'b1 : 1'b0;
												assign node1107 = (inp[13]) ? 1'b0 : node1108;
													assign node1108 = (inp[2]) ? node1110 : 1'b1;
														assign node1110 = (inp[7]) ? node1116 : node1111;
															assign node1111 = (inp[9]) ? node1113 : 1'b0;
																assign node1113 = (inp[10]) ? 1'b0 : 1'b1;
															assign node1116 = (inp[10]) ? 1'b1 : node1117;
																assign node1117 = (inp[9]) ? 1'b0 : 1'b1;
							assign node1123 = (inp[2]) ? node1197 : node1124;
								assign node1124 = (inp[15]) ? node1176 : node1125;
									assign node1125 = (inp[12]) ? node1135 : node1126;
										assign node1126 = (inp[5]) ? 1'b1 : node1127;
											assign node1127 = (inp[6]) ? node1129 : 1'b1;
												assign node1129 = (inp[7]) ? 1'b0 : node1130;
													assign node1130 = (inp[3]) ? 1'b1 : 1'b0;
										assign node1135 = (inp[5]) ? node1157 : node1136;
											assign node1136 = (inp[6]) ? 1'b1 : node1137;
												assign node1137 = (inp[7]) ? node1151 : node1138;
													assign node1138 = (inp[10]) ? node1148 : node1139;
														assign node1139 = (inp[13]) ? node1141 : 1'b1;
															assign node1141 = (inp[9]) ? node1145 : node1142;
																assign node1142 = (inp[3]) ? 1'b1 : 1'b0;
																assign node1145 = (inp[3]) ? 1'b0 : 1'b1;
														assign node1148 = (inp[9]) ? 1'b0 : 1'b1;
													assign node1151 = (inp[9]) ? node1153 : 1'b0;
														assign node1153 = (inp[10]) ? 1'b0 : 1'b1;
											assign node1157 = (inp[9]) ? node1163 : node1158;
												assign node1158 = (inp[7]) ? 1'b0 : node1159;
													assign node1159 = (inp[3]) ? 1'b1 : 1'b0;
												assign node1163 = (inp[10]) ? node1169 : node1164;
													assign node1164 = (inp[7]) ? 1'b1 : node1165;
														assign node1165 = (inp[3]) ? 1'b0 : 1'b1;
													assign node1169 = (inp[13]) ? 1'b0 : node1170;
														assign node1170 = (inp[3]) ? node1172 : 1'b0;
															assign node1172 = (inp[7]) ? 1'b0 : 1'b1;
									assign node1176 = (inp[5]) ? 1'b1 : node1177;
										assign node1177 = (inp[6]) ? node1179 : 1'b1;
											assign node1179 = (inp[7]) ? node1191 : node1180;
												assign node1180 = (inp[9]) ? node1184 : node1181;
													assign node1181 = (inp[3]) ? 1'b1 : 1'b0;
													assign node1184 = (inp[3]) ? node1188 : node1185;
														assign node1185 = (inp[10]) ? 1'b0 : 1'b1;
														assign node1188 = (inp[10]) ? 1'b1 : 1'b0;
												assign node1191 = (inp[9]) ? node1193 : 1'b0;
													assign node1193 = (inp[10]) ? 1'b0 : 1'b1;
								assign node1197 = (inp[15]) ? node1251 : node1198;
									assign node1198 = (inp[12]) ? node1214 : node1199;
										assign node1199 = (inp[6]) ? node1201 : 1'b0;
											assign node1201 = (inp[5]) ? 1'b0 : node1202;
												assign node1202 = (inp[10]) ? 1'b1 : node1203;
													assign node1203 = (inp[13]) ? 1'b0 : node1204;
														assign node1204 = (inp[7]) ? 1'b1 : node1205;
															assign node1205 = (inp[9]) ? 1'b1 : node1206;
																assign node1206 = (inp[3]) ? 1'b0 : 1'b1;
										assign node1214 = (inp[6]) ? node1232 : node1215;
											assign node1215 = (inp[7]) ? node1227 : node1216;
												assign node1216 = (inp[3]) ? node1222 : node1217;
													assign node1217 = (inp[9]) ? node1219 : 1'b1;
														assign node1219 = (inp[10]) ? 1'b1 : 1'b0;
													assign node1222 = (inp[9]) ? node1224 : 1'b0;
														assign node1224 = (inp[5]) ? 1'b1 : 1'b0;
												assign node1227 = (inp[10]) ? 1'b1 : node1228;
													assign node1228 = (inp[9]) ? 1'b0 : 1'b1;
											assign node1232 = (inp[5]) ? node1234 : 1'b0;
												assign node1234 = (inp[10]) ? node1246 : node1235;
													assign node1235 = (inp[13]) ? node1241 : node1236;
														assign node1236 = (inp[7]) ? 1'b0 : node1237;
															assign node1237 = (inp[9]) ? 1'b1 : 1'b0;
														assign node1241 = (inp[9]) ? node1243 : 1'b1;
															assign node1243 = (inp[7]) ? 1'b0 : 1'b1;
													assign node1246 = (inp[7]) ? 1'b1 : node1247;
														assign node1247 = (inp[9]) ? 1'b0 : 1'b1;
									assign node1251 = (inp[5]) ? 1'b0 : node1252;
										assign node1252 = (inp[6]) ? node1254 : 1'b0;
											assign node1254 = (inp[7]) ? node1268 : node1255;
												assign node1255 = (inp[12]) ? node1261 : node1256;
													assign node1256 = (inp[10]) ? 1'b0 : node1257;
														assign node1257 = (inp[9]) ? 1'b0 : 1'b1;
													assign node1261 = (inp[13]) ? 1'b1 : node1262;
														assign node1262 = (inp[9]) ? node1264 : 1'b0;
															assign node1264 = (inp[10]) ? 1'b1 : 1'b0;
												assign node1268 = (inp[9]) ? node1270 : 1'b1;
													assign node1270 = (inp[10]) ? 1'b1 : 1'b0;
					assign node1274 = (inp[12]) ? node1296 : node1275;
						assign node1275 = (inp[5]) ? 1'b1 : node1276;
							assign node1276 = (inp[6]) ? node1278 : 1'b1;
								assign node1278 = (inp[3]) ? node1284 : node1279;
									assign node1279 = (inp[9]) ? node1281 : 1'b0;
										assign node1281 = (inp[10]) ? 1'b0 : 1'b1;
									assign node1284 = (inp[7]) ? node1290 : node1285;
										assign node1285 = (inp[9]) ? node1287 : 1'b1;
											assign node1287 = (inp[10]) ? 1'b1 : 1'b0;
										assign node1290 = (inp[9]) ? node1292 : 1'b0;
											assign node1292 = (inp[10]) ? 1'b0 : 1'b1;
						assign node1296 = (inp[15]) ? node1334 : node1297;
							assign node1297 = (inp[5]) ? node1317 : node1298;
								assign node1298 = (inp[6]) ? 1'b1 : node1299;
									assign node1299 = (inp[3]) ? node1305 : node1300;
										assign node1300 = (inp[10]) ? 1'b0 : node1301;
											assign node1301 = (inp[9]) ? 1'b1 : 1'b0;
										assign node1305 = (inp[7]) ? node1311 : node1306;
											assign node1306 = (inp[10]) ? 1'b1 : node1307;
												assign node1307 = (inp[9]) ? 1'b0 : 1'b1;
											assign node1311 = (inp[10]) ? 1'b0 : node1312;
												assign node1312 = (inp[9]) ? 1'b1 : 1'b0;
								assign node1317 = (inp[7]) ? node1329 : node1318;
									assign node1318 = (inp[3]) ? node1324 : node1319;
										assign node1319 = (inp[9]) ? node1321 : 1'b0;
											assign node1321 = (inp[10]) ? 1'b0 : 1'b1;
										assign node1324 = (inp[9]) ? node1326 : 1'b1;
											assign node1326 = (inp[10]) ? 1'b1 : 1'b0;
									assign node1329 = (inp[9]) ? node1331 : 1'b0;
										assign node1331 = (inp[10]) ? 1'b0 : 1'b1;
							assign node1334 = (inp[5]) ? 1'b1 : node1335;
								assign node1335 = (inp[6]) ? node1337 : 1'b1;
									assign node1337 = (inp[10]) ? node1349 : node1338;
										assign node1338 = (inp[9]) ? node1344 : node1339;
											assign node1339 = (inp[3]) ? node1341 : 1'b0;
												assign node1341 = (inp[7]) ? 1'b0 : 1'b1;
											assign node1344 = (inp[7]) ? 1'b1 : node1345;
												assign node1345 = (inp[3]) ? 1'b0 : 1'b1;
										assign node1349 = (inp[3]) ? node1351 : 1'b0;
											assign node1351 = (inp[7]) ? 1'b0 : 1'b1;
				assign node1355 = (inp[11]) ? node1803 : node1356;
					assign node1356 = (inp[13]) ? node1578 : node1357;
						assign node1357 = (inp[14]) ? node1447 : node1358;
							assign node1358 = (inp[5]) ? node1426 : node1359;
								assign node1359 = (inp[10]) ? node1391 : node1360;
									assign node1360 = (inp[9]) ? node1380 : node1361;
										assign node1361 = (inp[6]) ? node1371 : node1362;
											assign node1362 = (inp[12]) ? node1364 : 1'b0;
												assign node1364 = (inp[2]) ? node1366 : 1'b0;
													assign node1366 = (inp[3]) ? node1368 : 1'b1;
														assign node1368 = (inp[7]) ? 1'b1 : 1'b0;
											assign node1371 = (inp[3]) ? node1377 : node1372;
												assign node1372 = (inp[12]) ? node1374 : 1'b1;
													assign node1374 = (inp[15]) ? 1'b1 : 1'b0;
												assign node1377 = (inp[2]) ? 1'b0 : 1'b1;
										assign node1380 = (inp[7]) ? 1'b0 : node1381;
											assign node1381 = (inp[3]) ? node1383 : 1'b0;
												assign node1383 = (inp[15]) ? 1'b1 : node1384;
													assign node1384 = (inp[6]) ? 1'b0 : node1385;
														assign node1385 = (inp[12]) ? 1'b1 : 1'b0;
									assign node1391 = (inp[7]) ? node1405 : node1392;
										assign node1392 = (inp[3]) ? 1'b0 : node1393;
											assign node1393 = (inp[12]) ? node1397 : node1394;
												assign node1394 = (inp[6]) ? 1'b1 : 1'b0;
												assign node1397 = (inp[6]) ? node1401 : node1398;
													assign node1398 = (inp[15]) ? 1'b0 : 1'b1;
													assign node1401 = (inp[15]) ? 1'b1 : 1'b0;
										assign node1405 = (inp[1]) ? node1415 : node1406;
											assign node1406 = (inp[9]) ? 1'b1 : node1407;
												assign node1407 = (inp[15]) ? 1'b0 : node1408;
													assign node1408 = (inp[3]) ? 1'b1 : node1409;
														assign node1409 = (inp[6]) ? 1'b0 : 1'b1;
											assign node1415 = (inp[6]) ? node1421 : node1416;
												assign node1416 = (inp[15]) ? 1'b0 : node1417;
													assign node1417 = (inp[12]) ? 1'b1 : 1'b0;
												assign node1421 = (inp[12]) ? node1423 : 1'b1;
													assign node1423 = (inp[15]) ? 1'b1 : 1'b0;
								assign node1426 = (inp[12]) ? node1428 : 1'b0;
									assign node1428 = (inp[15]) ? 1'b0 : node1429;
										assign node1429 = (inp[10]) ? node1441 : node1430;
											assign node1430 = (inp[9]) ? node1436 : node1431;
												assign node1431 = (inp[7]) ? 1'b1 : node1432;
													assign node1432 = (inp[3]) ? 1'b0 : 1'b1;
												assign node1436 = (inp[7]) ? 1'b0 : node1437;
													assign node1437 = (inp[3]) ? 1'b1 : 1'b0;
											assign node1441 = (inp[3]) ? node1443 : 1'b1;
												assign node1443 = (inp[7]) ? 1'b1 : 1'b0;
							assign node1447 = (inp[2]) ? node1509 : node1448;
								assign node1448 = (inp[15]) ? node1496 : node1449;
									assign node1449 = (inp[12]) ? node1465 : node1450;
										assign node1450 = (inp[5]) ? 1'b1 : node1451;
											assign node1451 = (inp[6]) ? node1453 : 1'b1;
												assign node1453 = (inp[3]) ? node1459 : node1454;
													assign node1454 = (inp[9]) ? node1456 : 1'b0;
														assign node1456 = (inp[10]) ? 1'b0 : 1'b1;
													assign node1459 = (inp[7]) ? node1461 : 1'b1;
														assign node1461 = (inp[10]) ? 1'b0 : 1'b1;
										assign node1465 = (inp[6]) ? node1481 : node1466;
											assign node1466 = (inp[9]) ? node1472 : node1467;
												assign node1467 = (inp[7]) ? 1'b0 : node1468;
													assign node1468 = (inp[3]) ? 1'b1 : 1'b0;
												assign node1472 = (inp[7]) ? node1478 : node1473;
													assign node1473 = (inp[10]) ? 1'b1 : node1474;
														assign node1474 = (inp[3]) ? 1'b0 : 1'b1;
													assign node1478 = (inp[10]) ? 1'b0 : 1'b1;
											assign node1481 = (inp[5]) ? node1483 : 1'b1;
												assign node1483 = (inp[3]) ? node1489 : node1484;
													assign node1484 = (inp[10]) ? 1'b0 : node1485;
														assign node1485 = (inp[9]) ? 1'b1 : 1'b0;
													assign node1489 = (inp[7]) ? node1491 : 1'b1;
														assign node1491 = (inp[9]) ? node1493 : 1'b0;
															assign node1493 = (inp[1]) ? 1'b0 : 1'b1;
									assign node1496 = (inp[5]) ? 1'b1 : node1497;
										assign node1497 = (inp[6]) ? node1499 : 1'b1;
											assign node1499 = (inp[10]) ? 1'b0 : node1500;
												assign node1500 = (inp[9]) ? node1502 : 1'b0;
													assign node1502 = (inp[3]) ? node1504 : 1'b1;
														assign node1504 = (inp[7]) ? 1'b1 : 1'b0;
								assign node1509 = (inp[10]) ? node1545 : node1510;
									assign node1510 = (inp[5]) ? node1536 : node1511;
										assign node1511 = (inp[6]) ? node1517 : node1512;
											assign node1512 = (inp[12]) ? node1514 : 1'b0;
												assign node1514 = (inp[15]) ? 1'b0 : 1'b1;
											assign node1517 = (inp[15]) ? node1525 : node1518;
												assign node1518 = (inp[12]) ? 1'b0 : node1519;
													assign node1519 = (inp[3]) ? 1'b0 : node1520;
														assign node1520 = (inp[9]) ? 1'b0 : 1'b1;
												assign node1525 = (inp[9]) ? node1531 : node1526;
													assign node1526 = (inp[3]) ? node1528 : 1'b1;
														assign node1528 = (inp[7]) ? 1'b1 : 1'b0;
													assign node1531 = (inp[3]) ? node1533 : 1'b0;
														assign node1533 = (inp[7]) ? 1'b0 : 1'b1;
										assign node1536 = (inp[15]) ? 1'b0 : node1537;
											assign node1537 = (inp[12]) ? node1539 : 1'b0;
												assign node1539 = (inp[3]) ? 1'b1 : node1540;
													assign node1540 = (inp[6]) ? 1'b0 : 1'b1;
									assign node1545 = (inp[3]) ? node1561 : node1546;
										assign node1546 = (inp[6]) ? node1552 : node1547;
											assign node1547 = (inp[12]) ? node1549 : 1'b0;
												assign node1549 = (inp[15]) ? 1'b0 : 1'b1;
											assign node1552 = (inp[5]) ? node1558 : node1553;
												assign node1553 = (inp[15]) ? 1'b1 : node1554;
													assign node1554 = (inp[12]) ? 1'b0 : 1'b1;
												assign node1558 = (inp[15]) ? 1'b0 : 1'b1;
										assign node1561 = (inp[7]) ? node1563 : 1'b0;
											assign node1563 = (inp[15]) ? node1571 : node1564;
												assign node1564 = (inp[12]) ? 1'b1 : node1565;
													assign node1565 = (inp[6]) ? node1567 : 1'b0;
														assign node1567 = (inp[5]) ? 1'b0 : 1'b1;
												assign node1571 = (inp[1]) ? node1573 : 1'b0;
													assign node1573 = (inp[6]) ? node1575 : 1'b0;
														assign node1575 = (inp[5]) ? 1'b0 : 1'b1;
						assign node1578 = (inp[14]) ? node1664 : node1579;
							assign node1579 = (inp[6]) ? node1597 : node1580;
								assign node1580 = (inp[12]) ? node1582 : 1'b1;
									assign node1582 = (inp[15]) ? 1'b1 : node1583;
										assign node1583 = (inp[7]) ? node1591 : node1584;
											assign node1584 = (inp[3]) ? node1586 : 1'b0;
												assign node1586 = (inp[10]) ? 1'b1 : node1587;
													assign node1587 = (inp[9]) ? 1'b0 : 1'b1;
											assign node1591 = (inp[9]) ? node1593 : 1'b0;
												assign node1593 = (inp[10]) ? 1'b0 : 1'b1;
								assign node1597 = (inp[5]) ? node1641 : node1598;
									assign node1598 = (inp[12]) ? node1616 : node1599;
										assign node1599 = (inp[7]) ? node1611 : node1600;
											assign node1600 = (inp[3]) ? node1606 : node1601;
												assign node1601 = (inp[2]) ? 1'b0 : node1602;
													assign node1602 = (inp[10]) ? 1'b0 : 1'b1;
												assign node1606 = (inp[9]) ? node1608 : 1'b1;
													assign node1608 = (inp[10]) ? 1'b1 : 1'b0;
											assign node1611 = (inp[9]) ? node1613 : 1'b0;
												assign node1613 = (inp[10]) ? 1'b0 : 1'b1;
										assign node1616 = (inp[15]) ? node1618 : 1'b1;
											assign node1618 = (inp[2]) ? node1628 : node1619;
												assign node1619 = (inp[9]) ? node1623 : node1620;
													assign node1620 = (inp[10]) ? 1'b1 : 1'b0;
													assign node1623 = (inp[3]) ? 1'b0 : node1624;
														assign node1624 = (inp[10]) ? 1'b0 : 1'b1;
												assign node1628 = (inp[10]) ? node1636 : node1629;
													assign node1629 = (inp[3]) ? node1631 : 1'b1;
														assign node1631 = (inp[9]) ? node1633 : 1'b1;
															assign node1633 = (inp[1]) ? 1'b1 : 1'b0;
													assign node1636 = (inp[7]) ? 1'b0 : node1637;
														assign node1637 = (inp[3]) ? 1'b1 : 1'b0;
									assign node1641 = (inp[12]) ? node1643 : 1'b1;
										assign node1643 = (inp[15]) ? 1'b1 : node1644;
											assign node1644 = (inp[7]) ? node1658 : node1645;
												assign node1645 = (inp[2]) ? node1653 : node1646;
													assign node1646 = (inp[10]) ? node1650 : node1647;
														assign node1647 = (inp[3]) ? 1'b0 : 1'b1;
														assign node1650 = (inp[3]) ? 1'b1 : 1'b0;
													assign node1653 = (inp[9]) ? node1655 : 1'b1;
														assign node1655 = (inp[3]) ? 1'b0 : 1'b1;
												assign node1658 = (inp[9]) ? node1660 : 1'b0;
													assign node1660 = (inp[10]) ? 1'b0 : 1'b1;
							assign node1664 = (inp[2]) ? node1732 : node1665;
								assign node1665 = (inp[5]) ? node1717 : node1666;
									assign node1666 = (inp[6]) ? node1682 : node1667;
										assign node1667 = (inp[12]) ? node1669 : 1'b0;
											assign node1669 = (inp[15]) ? 1'b0 : node1670;
												assign node1670 = (inp[7]) ? 1'b1 : node1671;
													assign node1671 = (inp[10]) ? 1'b0 : node1672;
														assign node1672 = (inp[1]) ? node1674 : 1'b1;
															assign node1674 = (inp[3]) ? node1676 : 1'b0;
																assign node1676 = (inp[9]) ? 1'b1 : 1'b0;
										assign node1682 = (inp[15]) ? node1700 : node1683;
											assign node1683 = (inp[12]) ? 1'b0 : node1684;
												assign node1684 = (inp[9]) ? node1690 : node1685;
													assign node1685 = (inp[3]) ? node1687 : 1'b1;
														assign node1687 = (inp[7]) ? 1'b1 : 1'b0;
													assign node1690 = (inp[7]) ? 1'b0 : node1691;
														assign node1691 = (inp[10]) ? node1695 : node1692;
															assign node1692 = (inp[1]) ? 1'b1 : 1'b0;
															assign node1695 = (inp[3]) ? 1'b0 : 1'b1;
											assign node1700 = (inp[3]) ? node1706 : node1701;
												assign node1701 = (inp[10]) ? 1'b1 : node1702;
													assign node1702 = (inp[9]) ? 1'b0 : 1'b1;
												assign node1706 = (inp[7]) ? node1712 : node1707;
													assign node1707 = (inp[9]) ? node1709 : 1'b0;
														assign node1709 = (inp[10]) ? 1'b0 : 1'b1;
													assign node1712 = (inp[9]) ? node1714 : 1'b1;
														assign node1714 = (inp[10]) ? 1'b1 : 1'b0;
									assign node1717 = (inp[15]) ? 1'b0 : node1718;
										assign node1718 = (inp[12]) ? node1720 : 1'b0;
											assign node1720 = (inp[3]) ? node1726 : node1721;
												assign node1721 = (inp[10]) ? 1'b1 : node1722;
													assign node1722 = (inp[9]) ? 1'b0 : 1'b1;
												assign node1726 = (inp[7]) ? node1728 : 1'b0;
													assign node1728 = (inp[6]) ? 1'b0 : 1'b1;
								assign node1732 = (inp[15]) ? node1782 : node1733;
									assign node1733 = (inp[12]) ? node1747 : node1734;
										assign node1734 = (inp[6]) ? node1736 : 1'b1;
											assign node1736 = (inp[5]) ? 1'b1 : node1737;
												assign node1737 = (inp[10]) ? 1'b0 : node1738;
													assign node1738 = (inp[1]) ? 1'b0 : node1739;
														assign node1739 = (inp[7]) ? 1'b1 : node1740;
															assign node1740 = (inp[3]) ? 1'b0 : 1'b1;
										assign node1747 = (inp[5]) ? node1765 : node1748;
											assign node1748 = (inp[6]) ? 1'b1 : node1749;
												assign node1749 = (inp[10]) ? node1759 : node1750;
													assign node1750 = (inp[9]) ? node1754 : node1751;
														assign node1751 = (inp[7]) ? 1'b0 : 1'b1;
														assign node1754 = (inp[7]) ? 1'b1 : node1755;
															assign node1755 = (inp[3]) ? 1'b0 : 1'b1;
													assign node1759 = (inp[3]) ? node1761 : 1'b0;
														assign node1761 = (inp[7]) ? 1'b0 : 1'b1;
											assign node1765 = (inp[10]) ? node1777 : node1766;
												assign node1766 = (inp[6]) ? node1772 : node1767;
													assign node1767 = (inp[9]) ? node1769 : 1'b0;
														assign node1769 = (inp[3]) ? 1'b0 : 1'b1;
													assign node1772 = (inp[3]) ? 1'b1 : node1773;
														assign node1773 = (inp[7]) ? 1'b1 : 1'b0;
												assign node1777 = (inp[3]) ? node1779 : 1'b0;
													assign node1779 = (inp[7]) ? 1'b0 : 1'b1;
									assign node1782 = (inp[5]) ? 1'b1 : node1783;
										assign node1783 = (inp[6]) ? node1785 : 1'b1;
											assign node1785 = (inp[10]) ? node1797 : node1786;
												assign node1786 = (inp[7]) ? node1794 : node1787;
													assign node1787 = (inp[9]) ? node1791 : node1788;
														assign node1788 = (inp[3]) ? 1'b1 : 1'b0;
														assign node1791 = (inp[3]) ? 1'b0 : 1'b1;
													assign node1794 = (inp[9]) ? 1'b1 : 1'b0;
												assign node1797 = (inp[3]) ? node1799 : 1'b0;
													assign node1799 = (inp[1]) ? 1'b1 : 1'b0;
					assign node1803 = (inp[2]) ? node1955 : node1804;
						assign node1804 = (inp[14]) ? node1880 : node1805;
							assign node1805 = (inp[5]) ? node1861 : node1806;
								assign node1806 = (inp[6]) ? node1826 : node1807;
									assign node1807 = (inp[12]) ? node1809 : 1'b0;
										assign node1809 = (inp[15]) ? 1'b0 : node1810;
											assign node1810 = (inp[10]) ? node1820 : node1811;
												assign node1811 = (inp[3]) ? node1815 : node1812;
													assign node1812 = (inp[9]) ? 1'b0 : 1'b1;
													assign node1815 = (inp[9]) ? node1817 : 1'b0;
														assign node1817 = (inp[1]) ? 1'b0 : 1'b1;
												assign node1820 = (inp[3]) ? node1822 : 1'b1;
													assign node1822 = (inp[7]) ? 1'b1 : 1'b0;
									assign node1826 = (inp[15]) ? node1844 : node1827;
										assign node1827 = (inp[12]) ? 1'b0 : node1828;
											assign node1828 = (inp[7]) ? 1'b1 : node1829;
												assign node1829 = (inp[10]) ? node1839 : node1830;
													assign node1830 = (inp[1]) ? node1836 : node1831;
														assign node1831 = (inp[9]) ? 1'b1 : node1832;
															assign node1832 = (inp[3]) ? 1'b0 : 1'b1;
														assign node1836 = (inp[13]) ? 1'b0 : 1'b1;
													assign node1839 = (inp[3]) ? 1'b0 : 1'b1;
										assign node1844 = (inp[7]) ? node1856 : node1845;
											assign node1845 = (inp[3]) ? node1851 : node1846;
												assign node1846 = (inp[9]) ? node1848 : 1'b1;
													assign node1848 = (inp[10]) ? 1'b1 : 1'b0;
												assign node1851 = (inp[9]) ? node1853 : 1'b0;
													assign node1853 = (inp[10]) ? 1'b0 : 1'b1;
											assign node1856 = (inp[9]) ? node1858 : 1'b1;
												assign node1858 = (inp[10]) ? 1'b1 : 1'b0;
								assign node1861 = (inp[12]) ? node1863 : 1'b0;
									assign node1863 = (inp[15]) ? 1'b0 : node1864;
										assign node1864 = (inp[3]) ? node1870 : node1865;
											assign node1865 = (inp[9]) ? node1867 : 1'b1;
												assign node1867 = (inp[10]) ? 1'b1 : 1'b0;
											assign node1870 = (inp[7]) ? node1876 : node1871;
												assign node1871 = (inp[10]) ? 1'b0 : node1872;
													assign node1872 = (inp[9]) ? 1'b1 : 1'b0;
												assign node1876 = (inp[10]) ? 1'b1 : 1'b0;
							assign node1880 = (inp[6]) ? node1902 : node1881;
								assign node1881 = (inp[15]) ? 1'b1 : node1882;
									assign node1882 = (inp[12]) ? node1884 : 1'b1;
										assign node1884 = (inp[3]) ? node1890 : node1885;
											assign node1885 = (inp[10]) ? 1'b0 : node1886;
												assign node1886 = (inp[9]) ? 1'b1 : 1'b0;
											assign node1890 = (inp[7]) ? node1898 : node1891;
												assign node1891 = (inp[1]) ? 1'b1 : node1892;
													assign node1892 = (inp[9]) ? node1894 : 1'b1;
														assign node1894 = (inp[10]) ? 1'b1 : 1'b0;
												assign node1898 = (inp[9]) ? 1'b1 : 1'b0;
								assign node1902 = (inp[5]) ? node1936 : node1903;
									assign node1903 = (inp[3]) ? node1917 : node1904;
										assign node1904 = (inp[9]) ? node1910 : node1905;
											assign node1905 = (inp[15]) ? 1'b0 : node1906;
												assign node1906 = (inp[12]) ? 1'b1 : 1'b0;
											assign node1910 = (inp[10]) ? node1912 : 1'b1;
												assign node1912 = (inp[12]) ? node1914 : 1'b0;
													assign node1914 = (inp[15]) ? 1'b0 : 1'b1;
										assign node1917 = (inp[7]) ? node1927 : node1918;
											assign node1918 = (inp[9]) ? node1920 : 1'b1;
												assign node1920 = (inp[10]) ? 1'b1 : node1921;
													assign node1921 = (inp[1]) ? 1'b0 : node1922;
														assign node1922 = (inp[12]) ? 1'b1 : 1'b0;
											assign node1927 = (inp[13]) ? node1929 : 1'b0;
												assign node1929 = (inp[1]) ? node1931 : 1'b1;
													assign node1931 = (inp[15]) ? node1933 : 1'b0;
														assign node1933 = (inp[10]) ? 1'b0 : 1'b1;
									assign node1936 = (inp[12]) ? node1938 : 1'b1;
										assign node1938 = (inp[15]) ? 1'b1 : node1939;
											assign node1939 = (inp[10]) ? node1949 : node1940;
												assign node1940 = (inp[9]) ? node1944 : node1941;
													assign node1941 = (inp[7]) ? 1'b0 : 1'b1;
													assign node1944 = (inp[3]) ? node1946 : 1'b1;
														assign node1946 = (inp[7]) ? 1'b1 : 1'b0;
												assign node1949 = (inp[7]) ? 1'b0 : node1950;
													assign node1950 = (inp[3]) ? 1'b1 : 1'b0;
						assign node1955 = (inp[15]) ? node2011 : node1956;
							assign node1956 = (inp[12]) ? node1974 : node1957;
								assign node1957 = (inp[5]) ? 1'b0 : node1958;
									assign node1958 = (inp[6]) ? node1960 : 1'b0;
										assign node1960 = (inp[7]) ? node1968 : node1961;
											assign node1961 = (inp[3]) ? 1'b0 : node1962;
												assign node1962 = (inp[9]) ? node1964 : 1'b1;
													assign node1964 = (inp[10]) ? 1'b1 : 1'b0;
											assign node1968 = (inp[10]) ? 1'b1 : node1969;
												assign node1969 = (inp[9]) ? 1'b0 : 1'b1;
								assign node1974 = (inp[6]) ? node1992 : node1975;
									assign node1975 = (inp[3]) ? node1981 : node1976;
										assign node1976 = (inp[10]) ? 1'b1 : node1977;
											assign node1977 = (inp[9]) ? 1'b0 : 1'b1;
										assign node1981 = (inp[7]) ? node1987 : node1982;
											assign node1982 = (inp[9]) ? node1984 : 1'b0;
												assign node1984 = (inp[10]) ? 1'b0 : 1'b1;
											assign node1987 = (inp[9]) ? node1989 : 1'b1;
												assign node1989 = (inp[10]) ? 1'b1 : 1'b0;
									assign node1992 = (inp[5]) ? node1994 : 1'b0;
										assign node1994 = (inp[10]) ? node2006 : node1995;
											assign node1995 = (inp[9]) ? node2001 : node1996;
												assign node1996 = (inp[3]) ? node1998 : 1'b1;
													assign node1998 = (inp[7]) ? 1'b1 : 1'b0;
												assign node2001 = (inp[7]) ? 1'b0 : node2002;
													assign node2002 = (inp[3]) ? 1'b1 : 1'b0;
											assign node2006 = (inp[3]) ? node2008 : 1'b1;
												assign node2008 = (inp[7]) ? 1'b1 : 1'b0;
							assign node2011 = (inp[6]) ? node2013 : 1'b0;
								assign node2013 = (inp[5]) ? 1'b0 : node2014;
									assign node2014 = (inp[7]) ? node2026 : node2015;
										assign node2015 = (inp[3]) ? node2021 : node2016;
											assign node2016 = (inp[9]) ? node2018 : 1'b1;
												assign node2018 = (inp[10]) ? 1'b1 : 1'b0;
											assign node2021 = (inp[9]) ? node2023 : 1'b0;
												assign node2023 = (inp[10]) ? 1'b0 : 1'b1;
										assign node2026 = (inp[9]) ? node2028 : 1'b1;
											assign node2028 = (inp[10]) ? 1'b1 : 1'b0;
		assign node2032 = (inp[1]) ? node2114 : node2033;
			assign node2033 = (inp[15]) ? node2093 : node2034;
				assign node2034 = (inp[12]) ? node2056 : node2035;
					assign node2035 = (inp[6]) ? node2037 : 1'b1;
						assign node2037 = (inp[5]) ? 1'b1 : node2038;
							assign node2038 = (inp[9]) ? node2044 : node2039;
								assign node2039 = (inp[7]) ? 1'b0 : node2040;
									assign node2040 = (inp[3]) ? 1'b1 : 1'b0;
								assign node2044 = (inp[10]) ? node2050 : node2045;
									assign node2045 = (inp[7]) ? 1'b1 : node2046;
										assign node2046 = (inp[3]) ? 1'b0 : 1'b1;
									assign node2050 = (inp[7]) ? 1'b0 : node2051;
										assign node2051 = (inp[3]) ? 1'b1 : 1'b0;
					assign node2056 = (inp[6]) ? node2074 : node2057;
						assign node2057 = (inp[3]) ? node2063 : node2058;
							assign node2058 = (inp[10]) ? 1'b0 : node2059;
								assign node2059 = (inp[9]) ? 1'b1 : 1'b0;
							assign node2063 = (inp[7]) ? node2069 : node2064;
								assign node2064 = (inp[10]) ? 1'b1 : node2065;
									assign node2065 = (inp[9]) ? 1'b0 : 1'b1;
								assign node2069 = (inp[10]) ? 1'b0 : node2070;
									assign node2070 = (inp[9]) ? 1'b1 : 1'b0;
						assign node2074 = (inp[5]) ? node2076 : 1'b1;
							assign node2076 = (inp[7]) ? node2088 : node2077;
								assign node2077 = (inp[3]) ? node2083 : node2078;
									assign node2078 = (inp[9]) ? node2080 : 1'b0;
										assign node2080 = (inp[10]) ? 1'b0 : 1'b1;
									assign node2083 = (inp[10]) ? 1'b1 : node2084;
										assign node2084 = (inp[9]) ? 1'b0 : 1'b1;
								assign node2088 = (inp[9]) ? node2090 : 1'b0;
									assign node2090 = (inp[10]) ? 1'b0 : 1'b1;
				assign node2093 = (inp[6]) ? node2095 : 1'b1;
					assign node2095 = (inp[5]) ? 1'b1 : node2096;
						assign node2096 = (inp[9]) ? node2102 : node2097;
							assign node2097 = (inp[3]) ? node2099 : 1'b0;
								assign node2099 = (inp[7]) ? 1'b0 : 1'b1;
							assign node2102 = (inp[10]) ? node2108 : node2103;
								assign node2103 = (inp[7]) ? 1'b1 : node2104;
									assign node2104 = (inp[3]) ? 1'b0 : 1'b1;
								assign node2108 = (inp[7]) ? 1'b0 : node2109;
									assign node2109 = (inp[3]) ? 1'b1 : 1'b0;
			assign node2114 = (inp[8]) ? node2778 : node2115;
				assign node2115 = (inp[2]) ? node2539 : node2116;
					assign node2116 = (inp[14]) ? node2318 : node2117;
						assign node2117 = (inp[11]) ? node2241 : node2118;
							assign node2118 = (inp[13]) ? node2178 : node2119;
								assign node2119 = (inp[5]) ? node2161 : node2120;
									assign node2120 = (inp[6]) ? node2130 : node2121;
										assign node2121 = (inp[15]) ? 1'b0 : node2122;
											assign node2122 = (inp[12]) ? node2124 : 1'b0;
												assign node2124 = (inp[0]) ? node2126 : 1'b1;
													assign node2126 = (inp[10]) ? 1'b1 : 1'b0;
										assign node2130 = (inp[12]) ? node2144 : node2131;
											assign node2131 = (inp[9]) ? node2137 : node2132;
												assign node2132 = (inp[7]) ? 1'b1 : node2133;
													assign node2133 = (inp[3]) ? 1'b0 : 1'b1;
												assign node2137 = (inp[10]) ? node2139 : 1'b0;
													assign node2139 = (inp[7]) ? 1'b1 : node2140;
														assign node2140 = (inp[3]) ? 1'b0 : 1'b1;
											assign node2144 = (inp[15]) ? node2146 : 1'b0;
												assign node2146 = (inp[9]) ? node2152 : node2147;
													assign node2147 = (inp[3]) ? node2149 : 1'b1;
														assign node2149 = (inp[7]) ? 1'b1 : 1'b0;
													assign node2152 = (inp[3]) ? node2154 : 1'b0;
														assign node2154 = (inp[0]) ? node2158 : node2155;
															assign node2155 = (inp[10]) ? 1'b1 : 1'b0;
															assign node2158 = (inp[10]) ? 1'b0 : 1'b1;
									assign node2161 = (inp[12]) ? node2163 : 1'b0;
										assign node2163 = (inp[15]) ? 1'b0 : node2164;
											assign node2164 = (inp[9]) ? node2170 : node2165;
												assign node2165 = (inp[3]) ? node2167 : 1'b1;
													assign node2167 = (inp[7]) ? 1'b1 : 1'b0;
												assign node2170 = (inp[10]) ? node2172 : 1'b0;
													assign node2172 = (inp[7]) ? 1'b1 : node2173;
														assign node2173 = (inp[3]) ? 1'b0 : 1'b1;
								assign node2178 = (inp[12]) ? node2200 : node2179;
									assign node2179 = (inp[6]) ? node2181 : 1'b1;
										assign node2181 = (inp[5]) ? 1'b1 : node2182;
											assign node2182 = (inp[3]) ? node2188 : node2183;
												assign node2183 = (inp[15]) ? node2185 : 1'b0;
													assign node2185 = (inp[9]) ? 1'b1 : 1'b0;
												assign node2188 = (inp[10]) ? node2196 : node2189;
													assign node2189 = (inp[0]) ? node2191 : 1'b0;
														assign node2191 = (inp[9]) ? 1'b1 : node2192;
															assign node2192 = (inp[7]) ? 1'b0 : 1'b1;
													assign node2196 = (inp[7]) ? 1'b0 : 1'b1;
									assign node2200 = (inp[15]) ? node2230 : node2201;
										assign node2201 = (inp[5]) ? node2213 : node2202;
											assign node2202 = (inp[6]) ? 1'b1 : node2203;
												assign node2203 = (inp[9]) ? node2205 : 1'b0;
													assign node2205 = (inp[7]) ? node2209 : node2206;
														assign node2206 = (inp[10]) ? 1'b1 : 1'b0;
														assign node2209 = (inp[10]) ? 1'b0 : 1'b1;
											assign node2213 = (inp[10]) ? node2225 : node2214;
												assign node2214 = (inp[9]) ? node2220 : node2215;
													assign node2215 = (inp[3]) ? node2217 : 1'b0;
														assign node2217 = (inp[7]) ? 1'b0 : 1'b1;
													assign node2220 = (inp[3]) ? node2222 : 1'b1;
														assign node2222 = (inp[7]) ? 1'b1 : 1'b0;
												assign node2225 = (inp[3]) ? node2227 : 1'b0;
													assign node2227 = (inp[7]) ? 1'b0 : 1'b1;
										assign node2230 = (inp[5]) ? 1'b1 : node2231;
											assign node2231 = (inp[6]) ? node2233 : 1'b1;
												assign node2233 = (inp[3]) ? node2235 : 1'b0;
													assign node2235 = (inp[7]) ? node2237 : 1'b1;
														assign node2237 = (inp[10]) ? 1'b0 : 1'b1;
							assign node2241 = (inp[5]) ? node2295 : node2242;
								assign node2242 = (inp[6]) ? node2262 : node2243;
									assign node2243 = (inp[12]) ? node2245 : 1'b0;
										assign node2245 = (inp[15]) ? 1'b0 : node2246;
											assign node2246 = (inp[10]) ? node2256 : node2247;
												assign node2247 = (inp[9]) ? node2253 : node2248;
													assign node2248 = (inp[7]) ? 1'b1 : node2249;
														assign node2249 = (inp[13]) ? 1'b0 : 1'b1;
													assign node2253 = (inp[13]) ? 1'b1 : 1'b0;
												assign node2256 = (inp[7]) ? 1'b1 : node2257;
													assign node2257 = (inp[3]) ? 1'b0 : 1'b1;
									assign node2262 = (inp[12]) ? node2280 : node2263;
										assign node2263 = (inp[9]) ? node2269 : node2264;
											assign node2264 = (inp[3]) ? node2266 : 1'b1;
												assign node2266 = (inp[7]) ? 1'b1 : 1'b0;
											assign node2269 = (inp[10]) ? node2275 : node2270;
												assign node2270 = (inp[7]) ? 1'b0 : node2271;
													assign node2271 = (inp[3]) ? 1'b1 : 1'b0;
												assign node2275 = (inp[7]) ? 1'b1 : node2276;
													assign node2276 = (inp[3]) ? 1'b0 : 1'b1;
										assign node2280 = (inp[15]) ? node2282 : 1'b0;
											assign node2282 = (inp[7]) ? node2290 : node2283;
												assign node2283 = (inp[3]) ? 1'b0 : node2284;
													assign node2284 = (inp[10]) ? 1'b1 : node2285;
														assign node2285 = (inp[9]) ? 1'b0 : 1'b1;
												assign node2290 = (inp[9]) ? node2292 : 1'b1;
													assign node2292 = (inp[10]) ? 1'b1 : 1'b0;
								assign node2295 = (inp[12]) ? node2297 : 1'b0;
									assign node2297 = (inp[15]) ? 1'b0 : node2298;
										assign node2298 = (inp[9]) ? node2304 : node2299;
											assign node2299 = (inp[3]) ? node2301 : 1'b1;
												assign node2301 = (inp[7]) ? 1'b1 : 1'b0;
											assign node2304 = (inp[7]) ? node2314 : node2305;
												assign node2305 = (inp[0]) ? node2307 : 1'b1;
													assign node2307 = (inp[6]) ? node2309 : 1'b0;
														assign node2309 = (inp[3]) ? node2311 : 1'b1;
															assign node2311 = (inp[13]) ? 1'b0 : 1'b1;
												assign node2314 = (inp[10]) ? 1'b1 : 1'b0;
						assign node2318 = (inp[11]) ? node2452 : node2319;
							assign node2319 = (inp[13]) ? node2373 : node2320;
								assign node2320 = (inp[5]) ? node2358 : node2321;
									assign node2321 = (inp[6]) ? node2333 : node2322;
										assign node2322 = (inp[15]) ? 1'b1 : node2323;
											assign node2323 = (inp[12]) ? node2325 : 1'b1;
												assign node2325 = (inp[3]) ? node2327 : 1'b0;
													assign node2327 = (inp[10]) ? node2329 : 1'b1;
														assign node2329 = (inp[7]) ? 1'b0 : 1'b1;
										assign node2333 = (inp[7]) ? node2347 : node2334;
											assign node2334 = (inp[12]) ? 1'b1 : node2335;
												assign node2335 = (inp[3]) ? node2341 : node2336;
													assign node2336 = (inp[9]) ? node2338 : 1'b0;
														assign node2338 = (inp[15]) ? 1'b0 : 1'b1;
													assign node2341 = (inp[9]) ? node2343 : 1'b1;
														assign node2343 = (inp[15]) ? 1'b0 : 1'b1;
											assign node2347 = (inp[10]) ? node2353 : node2348;
												assign node2348 = (inp[9]) ? 1'b1 : node2349;
													assign node2349 = (inp[15]) ? 1'b0 : 1'b1;
												assign node2353 = (inp[12]) ? node2355 : 1'b0;
													assign node2355 = (inp[15]) ? 1'b0 : 1'b1;
									assign node2358 = (inp[15]) ? 1'b1 : node2359;
										assign node2359 = (inp[12]) ? node2361 : 1'b1;
											assign node2361 = (inp[7]) ? node2367 : node2362;
												assign node2362 = (inp[3]) ? 1'b1 : node2363;
													assign node2363 = (inp[10]) ? 1'b0 : 1'b1;
												assign node2367 = (inp[9]) ? node2369 : 1'b0;
													assign node2369 = (inp[10]) ? 1'b0 : 1'b1;
								assign node2373 = (inp[10]) ? node2405 : node2374;
									assign node2374 = (inp[9]) ? node2396 : node2375;
										assign node2375 = (inp[7]) ? node2381 : node2376;
											assign node2376 = (inp[3]) ? 1'b0 : node2377;
												assign node2377 = (inp[0]) ? 1'b0 : 1'b1;
											assign node2381 = (inp[6]) ? node2387 : node2382;
												assign node2382 = (inp[15]) ? 1'b0 : node2383;
													assign node2383 = (inp[12]) ? 1'b1 : 1'b0;
												assign node2387 = (inp[0]) ? node2389 : 1'b1;
													assign node2389 = (inp[5]) ? node2393 : node2390;
														assign node2390 = (inp[15]) ? 1'b1 : 1'b0;
														assign node2393 = (inp[15]) ? 1'b0 : 1'b1;
										assign node2396 = (inp[6]) ? 1'b0 : node2397;
											assign node2397 = (inp[15]) ? 1'b0 : node2398;
												assign node2398 = (inp[3]) ? node2400 : 1'b0;
													assign node2400 = (inp[7]) ? 1'b0 : 1'b1;
									assign node2405 = (inp[3]) ? node2423 : node2406;
										assign node2406 = (inp[5]) ? node2418 : node2407;
											assign node2407 = (inp[6]) ? node2413 : node2408;
												assign node2408 = (inp[15]) ? 1'b0 : node2409;
													assign node2409 = (inp[12]) ? 1'b1 : 1'b0;
												assign node2413 = (inp[15]) ? 1'b1 : node2414;
													assign node2414 = (inp[12]) ? 1'b0 : 1'b1;
											assign node2418 = (inp[12]) ? node2420 : 1'b0;
												assign node2420 = (inp[15]) ? 1'b0 : 1'b1;
										assign node2423 = (inp[7]) ? node2425 : 1'b0;
											assign node2425 = (inp[12]) ? node2431 : node2426;
												assign node2426 = (inp[6]) ? node2428 : 1'b0;
													assign node2428 = (inp[5]) ? 1'b0 : 1'b1;
												assign node2431 = (inp[5]) ? 1'b1 : node2432;
													assign node2432 = (inp[0]) ? node2446 : node2433;
														assign node2433 = (inp[9]) ? node2441 : node2434;
															assign node2434 = (inp[6]) ? node2438 : node2435;
																assign node2435 = (inp[15]) ? 1'b0 : 1'b1;
																assign node2438 = (inp[15]) ? 1'b1 : 1'b0;
															assign node2441 = (inp[15]) ? node2443 : 1'b1;
																assign node2443 = (inp[6]) ? 1'b1 : 1'b0;
														assign node2446 = (inp[6]) ? node2448 : 1'b0;
															assign node2448 = (inp[15]) ? 1'b1 : 1'b0;
							assign node2452 = (inp[5]) ? node2504 : node2453;
								assign node2453 = (inp[6]) ? node2471 : node2454;
									assign node2454 = (inp[12]) ? node2456 : 1'b1;
										assign node2456 = (inp[15]) ? 1'b1 : node2457;
											assign node2457 = (inp[10]) ? node2465 : node2458;
												assign node2458 = (inp[3]) ? node2460 : 1'b1;
													assign node2460 = (inp[7]) ? 1'b0 : node2461;
														assign node2461 = (inp[9]) ? 1'b0 : 1'b1;
												assign node2465 = (inp[7]) ? 1'b0 : node2466;
													assign node2466 = (inp[3]) ? 1'b1 : 1'b0;
									assign node2471 = (inp[12]) ? node2489 : node2472;
										assign node2472 = (inp[9]) ? node2478 : node2473;
											assign node2473 = (inp[7]) ? 1'b0 : node2474;
												assign node2474 = (inp[3]) ? 1'b1 : 1'b0;
											assign node2478 = (inp[10]) ? node2484 : node2479;
												assign node2479 = (inp[3]) ? node2481 : 1'b1;
													assign node2481 = (inp[7]) ? 1'b1 : 1'b0;
												assign node2484 = (inp[7]) ? 1'b0 : node2485;
													assign node2485 = (inp[3]) ? 1'b1 : 1'b0;
										assign node2489 = (inp[15]) ? node2491 : 1'b1;
											assign node2491 = (inp[3]) ? node2493 : 1'b0;
												assign node2493 = (inp[7]) ? node2499 : node2494;
													assign node2494 = (inp[10]) ? 1'b1 : node2495;
														assign node2495 = (inp[9]) ? 1'b0 : 1'b1;
													assign node2499 = (inp[10]) ? 1'b0 : node2500;
														assign node2500 = (inp[9]) ? 1'b1 : 1'b0;
								assign node2504 = (inp[15]) ? 1'b1 : node2505;
									assign node2505 = (inp[12]) ? node2507 : 1'b1;
										assign node2507 = (inp[0]) ? node2523 : node2508;
											assign node2508 = (inp[10]) ? node2520 : node2509;
												assign node2509 = (inp[3]) ? node2513 : node2510;
													assign node2510 = (inp[9]) ? 1'b1 : 1'b0;
													assign node2513 = (inp[6]) ? node2515 : 1'b1;
														assign node2515 = (inp[7]) ? 1'b1 : node2516;
															assign node2516 = (inp[9]) ? 1'b0 : 1'b1;
												assign node2520 = (inp[3]) ? 1'b1 : 1'b0;
											assign node2523 = (inp[9]) ? node2529 : node2524;
												assign node2524 = (inp[7]) ? 1'b0 : node2525;
													assign node2525 = (inp[3]) ? 1'b1 : 1'b0;
												assign node2529 = (inp[10]) ? node2535 : node2530;
													assign node2530 = (inp[7]) ? 1'b1 : node2531;
														assign node2531 = (inp[13]) ? 1'b0 : 1'b1;
													assign node2535 = (inp[3]) ? 1'b1 : 1'b0;
					assign node2539 = (inp[11]) ? node2697 : node2540;
						assign node2540 = (inp[13]) ? node2618 : node2541;
							assign node2541 = (inp[15]) ? node2597 : node2542;
								assign node2542 = (inp[12]) ? node2564 : node2543;
									assign node2543 = (inp[5]) ? 1'b0 : node2544;
										assign node2544 = (inp[6]) ? node2546 : 1'b0;
											assign node2546 = (inp[10]) ? node2558 : node2547;
												assign node2547 = (inp[9]) ? node2553 : node2548;
													assign node2548 = (inp[3]) ? node2550 : 1'b1;
														assign node2550 = (inp[0]) ? 1'b1 : 1'b0;
													assign node2553 = (inp[3]) ? node2555 : 1'b0;
														assign node2555 = (inp[7]) ? 1'b0 : 1'b1;
												assign node2558 = (inp[3]) ? node2560 : 1'b1;
													assign node2560 = (inp[7]) ? 1'b1 : 1'b0;
									assign node2564 = (inp[6]) ? node2582 : node2565;
										assign node2565 = (inp[9]) ? node2571 : node2566;
											assign node2566 = (inp[7]) ? 1'b1 : node2567;
												assign node2567 = (inp[3]) ? 1'b0 : 1'b1;
											assign node2571 = (inp[10]) ? node2577 : node2572;
												assign node2572 = (inp[7]) ? 1'b0 : node2573;
													assign node2573 = (inp[3]) ? 1'b1 : 1'b0;
												assign node2577 = (inp[3]) ? node2579 : 1'b1;
													assign node2579 = (inp[7]) ? 1'b1 : 1'b0;
										assign node2582 = (inp[5]) ? node2584 : 1'b0;
											assign node2584 = (inp[10]) ? node2590 : node2585;
												assign node2585 = (inp[9]) ? 1'b0 : node2586;
													assign node2586 = (inp[7]) ? 1'b1 : 1'b0;
												assign node2590 = (inp[0]) ? 1'b1 : node2591;
													assign node2591 = (inp[14]) ? 1'b1 : node2592;
														assign node2592 = (inp[7]) ? 1'b1 : 1'b0;
								assign node2597 = (inp[6]) ? node2599 : 1'b0;
									assign node2599 = (inp[5]) ? 1'b0 : node2600;
										assign node2600 = (inp[10]) ? node2612 : node2601;
											assign node2601 = (inp[12]) ? node2607 : node2602;
												assign node2602 = (inp[9]) ? 1'b0 : node2603;
													assign node2603 = (inp[3]) ? 1'b0 : 1'b1;
												assign node2607 = (inp[7]) ? 1'b0 : node2608;
													assign node2608 = (inp[9]) ? 1'b1 : 1'b0;
											assign node2612 = (inp[3]) ? node2614 : 1'b1;
												assign node2614 = (inp[7]) ? 1'b1 : 1'b0;
							assign node2618 = (inp[12]) ? node2640 : node2619;
								assign node2619 = (inp[5]) ? 1'b1 : node2620;
									assign node2620 = (inp[6]) ? node2622 : 1'b1;
										assign node2622 = (inp[7]) ? node2634 : node2623;
											assign node2623 = (inp[3]) ? node2629 : node2624;
												assign node2624 = (inp[9]) ? node2626 : 1'b0;
													assign node2626 = (inp[10]) ? 1'b0 : 1'b1;
												assign node2629 = (inp[10]) ? 1'b1 : node2630;
													assign node2630 = (inp[9]) ? 1'b0 : 1'b1;
											assign node2634 = (inp[9]) ? node2636 : 1'b0;
												assign node2636 = (inp[10]) ? 1'b0 : 1'b1;
								assign node2640 = (inp[15]) ? node2676 : node2641;
									assign node2641 = (inp[5]) ? node2657 : node2642;
										assign node2642 = (inp[6]) ? 1'b1 : node2643;
											assign node2643 = (inp[9]) ? node2649 : node2644;
												assign node2644 = (inp[7]) ? 1'b0 : node2645;
													assign node2645 = (inp[3]) ? 1'b1 : 1'b0;
												assign node2649 = (inp[10]) ? 1'b0 : node2650;
													assign node2650 = (inp[3]) ? node2652 : 1'b1;
														assign node2652 = (inp[7]) ? 1'b1 : 1'b0;
										assign node2657 = (inp[7]) ? node2671 : node2658;
											assign node2658 = (inp[3]) ? node2666 : node2659;
												assign node2659 = (inp[6]) ? 1'b0 : node2660;
													assign node2660 = (inp[9]) ? node2662 : 1'b0;
														assign node2662 = (inp[10]) ? 1'b0 : 1'b1;
												assign node2666 = (inp[9]) ? node2668 : 1'b1;
													assign node2668 = (inp[10]) ? 1'b1 : 1'b0;
											assign node2671 = (inp[10]) ? 1'b0 : node2672;
												assign node2672 = (inp[9]) ? 1'b1 : 1'b0;
									assign node2676 = (inp[6]) ? node2678 : 1'b1;
										assign node2678 = (inp[5]) ? 1'b1 : node2679;
											assign node2679 = (inp[3]) ? node2685 : node2680;
												assign node2680 = (inp[9]) ? node2682 : 1'b0;
													assign node2682 = (inp[10]) ? 1'b0 : 1'b1;
												assign node2685 = (inp[7]) ? node2691 : node2686;
													assign node2686 = (inp[10]) ? 1'b1 : node2687;
														assign node2687 = (inp[9]) ? 1'b0 : 1'b1;
													assign node2691 = (inp[9]) ? node2693 : 1'b0;
														assign node2693 = (inp[10]) ? 1'b0 : 1'b1;
						assign node2697 = (inp[12]) ? node2719 : node2698;
							assign node2698 = (inp[6]) ? node2700 : 1'b0;
								assign node2700 = (inp[5]) ? 1'b0 : node2701;
									assign node2701 = (inp[3]) ? node2707 : node2702;
										assign node2702 = (inp[9]) ? node2704 : 1'b1;
											assign node2704 = (inp[10]) ? 1'b1 : 1'b0;
										assign node2707 = (inp[9]) ? node2711 : node2708;
											assign node2708 = (inp[7]) ? 1'b1 : 1'b0;
											assign node2711 = (inp[7]) ? node2715 : node2712;
												assign node2712 = (inp[10]) ? 1'b0 : 1'b1;
												assign node2715 = (inp[10]) ? 1'b1 : 1'b0;
							assign node2719 = (inp[15]) ? node2757 : node2720;
								assign node2720 = (inp[5]) ? node2740 : node2721;
									assign node2721 = (inp[6]) ? 1'b0 : node2722;
										assign node2722 = (inp[9]) ? node2728 : node2723;
											assign node2723 = (inp[7]) ? 1'b1 : node2724;
												assign node2724 = (inp[3]) ? 1'b0 : 1'b1;
											assign node2728 = (inp[10]) ? node2734 : node2729;
												assign node2729 = (inp[7]) ? 1'b0 : node2730;
													assign node2730 = (inp[3]) ? 1'b1 : 1'b0;
												assign node2734 = (inp[7]) ? 1'b1 : node2735;
													assign node2735 = (inp[3]) ? 1'b0 : 1'b1;
									assign node2740 = (inp[7]) ? node2752 : node2741;
										assign node2741 = (inp[3]) ? node2747 : node2742;
											assign node2742 = (inp[9]) ? node2744 : 1'b1;
												assign node2744 = (inp[10]) ? 1'b1 : 1'b0;
											assign node2747 = (inp[9]) ? node2749 : 1'b0;
												assign node2749 = (inp[10]) ? 1'b0 : 1'b1;
										assign node2752 = (inp[9]) ? node2754 : 1'b1;
											assign node2754 = (inp[10]) ? 1'b1 : 1'b0;
								assign node2757 = (inp[5]) ? 1'b0 : node2758;
									assign node2758 = (inp[6]) ? node2760 : 1'b0;
										assign node2760 = (inp[9]) ? node2766 : node2761;
											assign node2761 = (inp[7]) ? 1'b1 : node2762;
												assign node2762 = (inp[3]) ? 1'b0 : 1'b1;
											assign node2766 = (inp[10]) ? node2772 : node2767;
												assign node2767 = (inp[3]) ? node2769 : 1'b0;
													assign node2769 = (inp[7]) ? 1'b0 : 1'b1;
												assign node2772 = (inp[3]) ? node2774 : 1'b1;
													assign node2774 = (inp[7]) ? 1'b1 : 1'b0;
				assign node2778 = (inp[5]) ? node2838 : node2779;
					assign node2779 = (inp[6]) ? node2801 : node2780;
						assign node2780 = (inp[15]) ? 1'b1 : node2781;
							assign node2781 = (inp[12]) ? node2783 : 1'b1;
								assign node2783 = (inp[9]) ? node2789 : node2784;
									assign node2784 = (inp[3]) ? node2786 : 1'b0;
										assign node2786 = (inp[7]) ? 1'b0 : 1'b1;
									assign node2789 = (inp[10]) ? node2795 : node2790;
										assign node2790 = (inp[7]) ? 1'b1 : node2791;
											assign node2791 = (inp[3]) ? 1'b0 : 1'b1;
										assign node2795 = (inp[7]) ? 1'b0 : node2796;
											assign node2796 = (inp[3]) ? 1'b1 : 1'b0;
						assign node2801 = (inp[12]) ? node2819 : node2802;
							assign node2802 = (inp[3]) ? node2808 : node2803;
								assign node2803 = (inp[9]) ? node2805 : 1'b0;
									assign node2805 = (inp[10]) ? 1'b0 : 1'b1;
								assign node2808 = (inp[7]) ? node2814 : node2809;
									assign node2809 = (inp[9]) ? node2811 : 1'b1;
										assign node2811 = (inp[10]) ? 1'b1 : 1'b0;
									assign node2814 = (inp[9]) ? node2816 : 1'b0;
										assign node2816 = (inp[10]) ? 1'b0 : 1'b1;
							assign node2819 = (inp[15]) ? node2821 : 1'b1;
								assign node2821 = (inp[7]) ? node2833 : node2822;
									assign node2822 = (inp[3]) ? node2828 : node2823;
										assign node2823 = (inp[9]) ? node2825 : 1'b0;
											assign node2825 = (inp[10]) ? 1'b0 : 1'b1;
										assign node2828 = (inp[10]) ? 1'b1 : node2829;
											assign node2829 = (inp[9]) ? 1'b0 : 1'b1;
									assign node2833 = (inp[10]) ? 1'b0 : node2834;
										assign node2834 = (inp[9]) ? 1'b1 : 1'b0;
					assign node2838 = (inp[15]) ? 1'b1 : node2839;
						assign node2839 = (inp[12]) ? node2841 : 1'b1;
							assign node2841 = (inp[3]) ? node2847 : node2842;
								assign node2842 = (inp[9]) ? node2844 : 1'b0;
									assign node2844 = (inp[10]) ? 1'b0 : 1'b1;
								assign node2847 = (inp[7]) ? node2853 : node2848;
									assign node2848 = (inp[10]) ? 1'b1 : node2849;
										assign node2849 = (inp[9]) ? 1'b0 : 1'b1;
									assign node2853 = (inp[10]) ? 1'b0 : node2854;
										assign node2854 = (inp[9]) ? 1'b1 : 1'b0;

endmodule