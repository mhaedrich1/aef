module dtc_split875_bm83 (
	input  wire [12-1:0] inp,
	output wire [3-1:0] outp
);

	wire [3-1:0] node1;
	wire [3-1:0] node2;
	wire [3-1:0] node3;
	wire [3-1:0] node4;
	wire [3-1:0] node5;
	wire [3-1:0] node6;
	wire [3-1:0] node7;
	wire [3-1:0] node8;
	wire [3-1:0] node9;
	wire [3-1:0] node12;
	wire [3-1:0] node15;
	wire [3-1:0] node16;
	wire [3-1:0] node19;
	wire [3-1:0] node22;
	wire [3-1:0] node23;
	wire [3-1:0] node24;
	wire [3-1:0] node28;
	wire [3-1:0] node29;
	wire [3-1:0] node32;
	wire [3-1:0] node35;
	wire [3-1:0] node36;
	wire [3-1:0] node37;
	wire [3-1:0] node38;
	wire [3-1:0] node41;
	wire [3-1:0] node44;
	wire [3-1:0] node45;
	wire [3-1:0] node48;
	wire [3-1:0] node51;
	wire [3-1:0] node52;
	wire [3-1:0] node53;
	wire [3-1:0] node56;
	wire [3-1:0] node59;
	wire [3-1:0] node60;
	wire [3-1:0] node63;
	wire [3-1:0] node66;
	wire [3-1:0] node67;
	wire [3-1:0] node68;
	wire [3-1:0] node69;
	wire [3-1:0] node72;
	wire [3-1:0] node74;
	wire [3-1:0] node77;
	wire [3-1:0] node78;
	wire [3-1:0] node79;
	wire [3-1:0] node82;
	wire [3-1:0] node85;
	wire [3-1:0] node86;
	wire [3-1:0] node90;
	wire [3-1:0] node91;
	wire [3-1:0] node92;
	wire [3-1:0] node93;
	wire [3-1:0] node96;
	wire [3-1:0] node99;
	wire [3-1:0] node100;
	wire [3-1:0] node103;
	wire [3-1:0] node107;
	wire [3-1:0] node108;
	wire [3-1:0] node109;
	wire [3-1:0] node110;
	wire [3-1:0] node112;
	wire [3-1:0] node114;
	wire [3-1:0] node118;
	wire [3-1:0] node119;
	wire [3-1:0] node120;
	wire [3-1:0] node122;
	wire [3-1:0] node125;
	wire [3-1:0] node126;
	wire [3-1:0] node131;
	wire [3-1:0] node132;
	wire [3-1:0] node133;
	wire [3-1:0] node134;
	wire [3-1:0] node135;
	wire [3-1:0] node139;
	wire [3-1:0] node140;
	wire [3-1:0] node143;
	wire [3-1:0] node146;
	wire [3-1:0] node148;
	wire [3-1:0] node149;
	wire [3-1:0] node153;
	wire [3-1:0] node155;
	wire [3-1:0] node156;
	wire [3-1:0] node157;
	wire [3-1:0] node160;
	wire [3-1:0] node164;
	wire [3-1:0] node165;
	wire [3-1:0] node166;
	wire [3-1:0] node167;
	wire [3-1:0] node168;
	wire [3-1:0] node169;
	wire [3-1:0] node170;
	wire [3-1:0] node173;
	wire [3-1:0] node176;
	wire [3-1:0] node177;
	wire [3-1:0] node181;
	wire [3-1:0] node182;
	wire [3-1:0] node183;
	wire [3-1:0] node186;
	wire [3-1:0] node189;
	wire [3-1:0] node190;
	wire [3-1:0] node193;
	wire [3-1:0] node196;
	wire [3-1:0] node197;
	wire [3-1:0] node198;
	wire [3-1:0] node199;
	wire [3-1:0] node202;
	wire [3-1:0] node205;
	wire [3-1:0] node206;
	wire [3-1:0] node209;
	wire [3-1:0] node212;
	wire [3-1:0] node213;
	wire [3-1:0] node214;
	wire [3-1:0] node218;
	wire [3-1:0] node219;
	wire [3-1:0] node222;
	wire [3-1:0] node225;
	wire [3-1:0] node226;
	wire [3-1:0] node227;
	wire [3-1:0] node228;
	wire [3-1:0] node229;
	wire [3-1:0] node232;
	wire [3-1:0] node235;
	wire [3-1:0] node236;
	wire [3-1:0] node239;
	wire [3-1:0] node242;
	wire [3-1:0] node243;
	wire [3-1:0] node244;
	wire [3-1:0] node247;
	wire [3-1:0] node250;
	wire [3-1:0] node251;
	wire [3-1:0] node254;
	wire [3-1:0] node257;
	wire [3-1:0] node258;
	wire [3-1:0] node259;
	wire [3-1:0] node260;
	wire [3-1:0] node263;
	wire [3-1:0] node266;
	wire [3-1:0] node267;
	wire [3-1:0] node270;
	wire [3-1:0] node273;
	wire [3-1:0] node274;
	wire [3-1:0] node275;
	wire [3-1:0] node278;
	wire [3-1:0] node281;
	wire [3-1:0] node282;
	wire [3-1:0] node285;
	wire [3-1:0] node288;
	wire [3-1:0] node289;
	wire [3-1:0] node290;
	wire [3-1:0] node291;
	wire [3-1:0] node292;
	wire [3-1:0] node294;
	wire [3-1:0] node297;
	wire [3-1:0] node298;
	wire [3-1:0] node301;
	wire [3-1:0] node304;
	wire [3-1:0] node305;
	wire [3-1:0] node307;
	wire [3-1:0] node310;
	wire [3-1:0] node311;
	wire [3-1:0] node314;
	wire [3-1:0] node317;
	wire [3-1:0] node318;
	wire [3-1:0] node319;
	wire [3-1:0] node320;
	wire [3-1:0] node323;
	wire [3-1:0] node326;
	wire [3-1:0] node327;
	wire [3-1:0] node330;
	wire [3-1:0] node333;
	wire [3-1:0] node334;
	wire [3-1:0] node335;
	wire [3-1:0] node338;
	wire [3-1:0] node341;
	wire [3-1:0] node342;
	wire [3-1:0] node345;
	wire [3-1:0] node348;
	wire [3-1:0] node349;
	wire [3-1:0] node350;
	wire [3-1:0] node351;
	wire [3-1:0] node352;
	wire [3-1:0] node355;
	wire [3-1:0] node358;
	wire [3-1:0] node359;
	wire [3-1:0] node362;
	wire [3-1:0] node365;
	wire [3-1:0] node366;
	wire [3-1:0] node368;
	wire [3-1:0] node371;
	wire [3-1:0] node372;
	wire [3-1:0] node375;
	wire [3-1:0] node378;
	wire [3-1:0] node379;
	wire [3-1:0] node381;
	wire [3-1:0] node382;
	wire [3-1:0] node386;
	wire [3-1:0] node387;
	wire [3-1:0] node388;
	wire [3-1:0] node392;
	wire [3-1:0] node393;
	wire [3-1:0] node396;
	wire [3-1:0] node399;
	wire [3-1:0] node400;
	wire [3-1:0] node401;
	wire [3-1:0] node402;
	wire [3-1:0] node403;
	wire [3-1:0] node404;
	wire [3-1:0] node405;
	wire [3-1:0] node406;
	wire [3-1:0] node409;
	wire [3-1:0] node412;
	wire [3-1:0] node413;
	wire [3-1:0] node416;
	wire [3-1:0] node419;
	wire [3-1:0] node420;
	wire [3-1:0] node421;
	wire [3-1:0] node424;
	wire [3-1:0] node427;
	wire [3-1:0] node428;
	wire [3-1:0] node431;
	wire [3-1:0] node434;
	wire [3-1:0] node435;
	wire [3-1:0] node436;
	wire [3-1:0] node437;
	wire [3-1:0] node440;
	wire [3-1:0] node443;
	wire [3-1:0] node444;
	wire [3-1:0] node447;
	wire [3-1:0] node450;
	wire [3-1:0] node451;
	wire [3-1:0] node452;
	wire [3-1:0] node455;
	wire [3-1:0] node458;
	wire [3-1:0] node459;
	wire [3-1:0] node462;
	wire [3-1:0] node465;
	wire [3-1:0] node466;
	wire [3-1:0] node467;
	wire [3-1:0] node468;
	wire [3-1:0] node469;
	wire [3-1:0] node472;
	wire [3-1:0] node475;
	wire [3-1:0] node476;
	wire [3-1:0] node479;
	wire [3-1:0] node482;
	wire [3-1:0] node483;
	wire [3-1:0] node484;
	wire [3-1:0] node487;
	wire [3-1:0] node490;
	wire [3-1:0] node491;
	wire [3-1:0] node494;
	wire [3-1:0] node497;
	wire [3-1:0] node498;
	wire [3-1:0] node499;
	wire [3-1:0] node500;
	wire [3-1:0] node503;
	wire [3-1:0] node506;
	wire [3-1:0] node507;
	wire [3-1:0] node510;
	wire [3-1:0] node513;
	wire [3-1:0] node514;
	wire [3-1:0] node515;
	wire [3-1:0] node518;
	wire [3-1:0] node521;
	wire [3-1:0] node522;
	wire [3-1:0] node525;
	wire [3-1:0] node528;
	wire [3-1:0] node529;
	wire [3-1:0] node530;
	wire [3-1:0] node531;
	wire [3-1:0] node532;
	wire [3-1:0] node533;
	wire [3-1:0] node536;
	wire [3-1:0] node539;
	wire [3-1:0] node540;
	wire [3-1:0] node543;
	wire [3-1:0] node546;
	wire [3-1:0] node547;
	wire [3-1:0] node549;
	wire [3-1:0] node552;
	wire [3-1:0] node553;
	wire [3-1:0] node556;
	wire [3-1:0] node559;
	wire [3-1:0] node560;
	wire [3-1:0] node561;
	wire [3-1:0] node562;
	wire [3-1:0] node565;
	wire [3-1:0] node568;
	wire [3-1:0] node569;
	wire [3-1:0] node572;
	wire [3-1:0] node575;
	wire [3-1:0] node577;
	wire [3-1:0] node578;
	wire [3-1:0] node581;
	wire [3-1:0] node584;
	wire [3-1:0] node585;
	wire [3-1:0] node586;
	wire [3-1:0] node587;
	wire [3-1:0] node588;
	wire [3-1:0] node591;
	wire [3-1:0] node594;
	wire [3-1:0] node595;
	wire [3-1:0] node598;
	wire [3-1:0] node601;
	wire [3-1:0] node602;
	wire [3-1:0] node603;
	wire [3-1:0] node606;
	wire [3-1:0] node609;
	wire [3-1:0] node610;
	wire [3-1:0] node613;
	wire [3-1:0] node616;
	wire [3-1:0] node617;
	wire [3-1:0] node618;
	wire [3-1:0] node619;
	wire [3-1:0] node622;
	wire [3-1:0] node625;
	wire [3-1:0] node626;
	wire [3-1:0] node629;
	wire [3-1:0] node632;
	wire [3-1:0] node633;
	wire [3-1:0] node634;
	wire [3-1:0] node637;
	wire [3-1:0] node640;
	wire [3-1:0] node641;
	wire [3-1:0] node644;
	wire [3-1:0] node647;
	wire [3-1:0] node648;
	wire [3-1:0] node649;
	wire [3-1:0] node650;
	wire [3-1:0] node651;
	wire [3-1:0] node652;
	wire [3-1:0] node653;
	wire [3-1:0] node656;
	wire [3-1:0] node659;
	wire [3-1:0] node660;
	wire [3-1:0] node663;
	wire [3-1:0] node666;
	wire [3-1:0] node667;
	wire [3-1:0] node668;
	wire [3-1:0] node671;
	wire [3-1:0] node674;
	wire [3-1:0] node675;
	wire [3-1:0] node678;
	wire [3-1:0] node681;
	wire [3-1:0] node682;
	wire [3-1:0] node683;
	wire [3-1:0] node684;
	wire [3-1:0] node687;
	wire [3-1:0] node690;
	wire [3-1:0] node691;
	wire [3-1:0] node694;
	wire [3-1:0] node697;
	wire [3-1:0] node698;
	wire [3-1:0] node699;
	wire [3-1:0] node702;
	wire [3-1:0] node705;
	wire [3-1:0] node707;
	wire [3-1:0] node710;
	wire [3-1:0] node711;
	wire [3-1:0] node712;
	wire [3-1:0] node713;
	wire [3-1:0] node714;
	wire [3-1:0] node717;
	wire [3-1:0] node720;
	wire [3-1:0] node721;
	wire [3-1:0] node724;
	wire [3-1:0] node727;
	wire [3-1:0] node728;
	wire [3-1:0] node729;
	wire [3-1:0] node732;
	wire [3-1:0] node735;
	wire [3-1:0] node736;
	wire [3-1:0] node739;
	wire [3-1:0] node742;
	wire [3-1:0] node743;
	wire [3-1:0] node744;
	wire [3-1:0] node745;
	wire [3-1:0] node748;
	wire [3-1:0] node751;
	wire [3-1:0] node752;
	wire [3-1:0] node755;
	wire [3-1:0] node758;
	wire [3-1:0] node759;
	wire [3-1:0] node760;
	wire [3-1:0] node763;
	wire [3-1:0] node766;
	wire [3-1:0] node767;
	wire [3-1:0] node770;
	wire [3-1:0] node773;
	wire [3-1:0] node774;
	wire [3-1:0] node775;
	wire [3-1:0] node776;
	wire [3-1:0] node777;
	wire [3-1:0] node778;
	wire [3-1:0] node781;
	wire [3-1:0] node784;
	wire [3-1:0] node785;
	wire [3-1:0] node788;
	wire [3-1:0] node791;
	wire [3-1:0] node792;
	wire [3-1:0] node793;
	wire [3-1:0] node796;
	wire [3-1:0] node799;
	wire [3-1:0] node800;
	wire [3-1:0] node803;
	wire [3-1:0] node806;
	wire [3-1:0] node807;
	wire [3-1:0] node808;
	wire [3-1:0] node809;
	wire [3-1:0] node812;
	wire [3-1:0] node815;
	wire [3-1:0] node816;
	wire [3-1:0] node819;
	wire [3-1:0] node822;
	wire [3-1:0] node823;
	wire [3-1:0] node824;
	wire [3-1:0] node827;
	wire [3-1:0] node830;
	wire [3-1:0] node831;
	wire [3-1:0] node834;
	wire [3-1:0] node837;
	wire [3-1:0] node838;
	wire [3-1:0] node839;
	wire [3-1:0] node840;
	wire [3-1:0] node841;
	wire [3-1:0] node844;
	wire [3-1:0] node847;
	wire [3-1:0] node848;
	wire [3-1:0] node851;
	wire [3-1:0] node854;
	wire [3-1:0] node855;
	wire [3-1:0] node856;
	wire [3-1:0] node859;
	wire [3-1:0] node862;
	wire [3-1:0] node863;
	wire [3-1:0] node866;
	wire [3-1:0] node869;
	wire [3-1:0] node870;
	wire [3-1:0] node871;
	wire [3-1:0] node872;
	wire [3-1:0] node875;
	wire [3-1:0] node878;
	wire [3-1:0] node879;
	wire [3-1:0] node882;
	wire [3-1:0] node885;
	wire [3-1:0] node886;
	wire [3-1:0] node887;
	wire [3-1:0] node890;
	wire [3-1:0] node893;
	wire [3-1:0] node894;
	wire [3-1:0] node897;
	wire [3-1:0] node900;
	wire [3-1:0] node901;
	wire [3-1:0] node902;
	wire [3-1:0] node903;
	wire [3-1:0] node904;
	wire [3-1:0] node905;
	wire [3-1:0] node906;
	wire [3-1:0] node907;
	wire [3-1:0] node908;
	wire [3-1:0] node911;
	wire [3-1:0] node914;
	wire [3-1:0] node915;
	wire [3-1:0] node919;
	wire [3-1:0] node920;
	wire [3-1:0] node921;
	wire [3-1:0] node924;
	wire [3-1:0] node928;
	wire [3-1:0] node929;
	wire [3-1:0] node930;
	wire [3-1:0] node933;
	wire [3-1:0] node934;
	wire [3-1:0] node937;
	wire [3-1:0] node940;
	wire [3-1:0] node941;
	wire [3-1:0] node942;
	wire [3-1:0] node946;
	wire [3-1:0] node947;
	wire [3-1:0] node950;
	wire [3-1:0] node953;
	wire [3-1:0] node954;
	wire [3-1:0] node955;
	wire [3-1:0] node956;
	wire [3-1:0] node957;
	wire [3-1:0] node960;
	wire [3-1:0] node963;
	wire [3-1:0] node964;
	wire [3-1:0] node967;
	wire [3-1:0] node970;
	wire [3-1:0] node972;
	wire [3-1:0] node973;
	wire [3-1:0] node976;
	wire [3-1:0] node979;
	wire [3-1:0] node980;
	wire [3-1:0] node981;
	wire [3-1:0] node982;
	wire [3-1:0] node985;
	wire [3-1:0] node988;
	wire [3-1:0] node989;
	wire [3-1:0] node992;
	wire [3-1:0] node995;
	wire [3-1:0] node996;
	wire [3-1:0] node997;
	wire [3-1:0] node1000;
	wire [3-1:0] node1003;
	wire [3-1:0] node1004;
	wire [3-1:0] node1007;
	wire [3-1:0] node1010;
	wire [3-1:0] node1011;
	wire [3-1:0] node1012;
	wire [3-1:0] node1013;
	wire [3-1:0] node1014;
	wire [3-1:0] node1015;
	wire [3-1:0] node1018;
	wire [3-1:0] node1021;
	wire [3-1:0] node1022;
	wire [3-1:0] node1025;
	wire [3-1:0] node1028;
	wire [3-1:0] node1029;
	wire [3-1:0] node1030;
	wire [3-1:0] node1033;
	wire [3-1:0] node1036;
	wire [3-1:0] node1037;
	wire [3-1:0] node1040;
	wire [3-1:0] node1043;
	wire [3-1:0] node1044;
	wire [3-1:0] node1045;
	wire [3-1:0] node1046;
	wire [3-1:0] node1049;
	wire [3-1:0] node1052;
	wire [3-1:0] node1053;
	wire [3-1:0] node1056;
	wire [3-1:0] node1059;
	wire [3-1:0] node1060;
	wire [3-1:0] node1061;
	wire [3-1:0] node1064;
	wire [3-1:0] node1067;
	wire [3-1:0] node1068;
	wire [3-1:0] node1071;
	wire [3-1:0] node1074;
	wire [3-1:0] node1075;
	wire [3-1:0] node1076;
	wire [3-1:0] node1077;
	wire [3-1:0] node1078;
	wire [3-1:0] node1081;
	wire [3-1:0] node1084;
	wire [3-1:0] node1085;
	wire [3-1:0] node1088;
	wire [3-1:0] node1091;
	wire [3-1:0] node1092;
	wire [3-1:0] node1093;
	wire [3-1:0] node1096;
	wire [3-1:0] node1099;
	wire [3-1:0] node1100;
	wire [3-1:0] node1103;
	wire [3-1:0] node1106;
	wire [3-1:0] node1107;
	wire [3-1:0] node1108;
	wire [3-1:0] node1109;
	wire [3-1:0] node1112;
	wire [3-1:0] node1115;
	wire [3-1:0] node1116;
	wire [3-1:0] node1119;
	wire [3-1:0] node1122;
	wire [3-1:0] node1123;
	wire [3-1:0] node1124;
	wire [3-1:0] node1127;
	wire [3-1:0] node1130;
	wire [3-1:0] node1131;
	wire [3-1:0] node1134;
	wire [3-1:0] node1137;
	wire [3-1:0] node1138;
	wire [3-1:0] node1139;
	wire [3-1:0] node1141;
	wire [3-1:0] node1142;
	wire [3-1:0] node1143;
	wire [3-1:0] node1144;
	wire [3-1:0] node1148;
	wire [3-1:0] node1149;
	wire [3-1:0] node1152;
	wire [3-1:0] node1155;
	wire [3-1:0] node1156;
	wire [3-1:0] node1158;
	wire [3-1:0] node1162;
	wire [3-1:0] node1163;
	wire [3-1:0] node1164;
	wire [3-1:0] node1165;
	wire [3-1:0] node1166;
	wire [3-1:0] node1169;
	wire [3-1:0] node1172;
	wire [3-1:0] node1173;
	wire [3-1:0] node1176;
	wire [3-1:0] node1179;
	wire [3-1:0] node1180;
	wire [3-1:0] node1182;
	wire [3-1:0] node1185;
	wire [3-1:0] node1186;
	wire [3-1:0] node1189;
	wire [3-1:0] node1192;
	wire [3-1:0] node1193;
	wire [3-1:0] node1194;
	wire [3-1:0] node1196;
	wire [3-1:0] node1199;
	wire [3-1:0] node1200;
	wire [3-1:0] node1203;
	wire [3-1:0] node1206;
	wire [3-1:0] node1207;
	wire [3-1:0] node1209;
	wire [3-1:0] node1213;
	wire [3-1:0] node1214;
	wire [3-1:0] node1215;
	wire [3-1:0] node1216;
	wire [3-1:0] node1217;
	wire [3-1:0] node1218;
	wire [3-1:0] node1221;
	wire [3-1:0] node1224;
	wire [3-1:0] node1225;
	wire [3-1:0] node1228;
	wire [3-1:0] node1231;
	wire [3-1:0] node1232;
	wire [3-1:0] node1233;
	wire [3-1:0] node1236;
	wire [3-1:0] node1239;
	wire [3-1:0] node1240;
	wire [3-1:0] node1243;
	wire [3-1:0] node1246;
	wire [3-1:0] node1247;
	wire [3-1:0] node1248;
	wire [3-1:0] node1250;
	wire [3-1:0] node1253;
	wire [3-1:0] node1254;
	wire [3-1:0] node1257;
	wire [3-1:0] node1260;
	wire [3-1:0] node1262;
	wire [3-1:0] node1264;
	wire [3-1:0] node1267;
	wire [3-1:0] node1268;
	wire [3-1:0] node1269;
	wire [3-1:0] node1270;
	wire [3-1:0] node1271;
	wire [3-1:0] node1274;
	wire [3-1:0] node1277;
	wire [3-1:0] node1278;
	wire [3-1:0] node1281;
	wire [3-1:0] node1284;
	wire [3-1:0] node1285;
	wire [3-1:0] node1286;
	wire [3-1:0] node1289;
	wire [3-1:0] node1292;
	wire [3-1:0] node1293;
	wire [3-1:0] node1296;
	wire [3-1:0] node1299;
	wire [3-1:0] node1300;
	wire [3-1:0] node1301;
	wire [3-1:0] node1302;
	wire [3-1:0] node1305;
	wire [3-1:0] node1308;
	wire [3-1:0] node1309;
	wire [3-1:0] node1312;
	wire [3-1:0] node1315;
	wire [3-1:0] node1316;
	wire [3-1:0] node1317;
	wire [3-1:0] node1320;
	wire [3-1:0] node1323;
	wire [3-1:0] node1324;
	wire [3-1:0] node1327;
	wire [3-1:0] node1330;
	wire [3-1:0] node1331;
	wire [3-1:0] node1332;
	wire [3-1:0] node1333;
	wire [3-1:0] node1335;
	wire [3-1:0] node1337;
	wire [3-1:0] node1338;
	wire [3-1:0] node1339;
	wire [3-1:0] node1342;
	wire [3-1:0] node1345;
	wire [3-1:0] node1346;
	wire [3-1:0] node1350;
	wire [3-1:0] node1351;
	wire [3-1:0] node1353;
	wire [3-1:0] node1354;
	wire [3-1:0] node1355;
	wire [3-1:0] node1358;
	wire [3-1:0] node1361;
	wire [3-1:0] node1362;
	wire [3-1:0] node1366;
	wire [3-1:0] node1367;
	wire [3-1:0] node1368;
	wire [3-1:0] node1369;
	wire [3-1:0] node1372;
	wire [3-1:0] node1375;
	wire [3-1:0] node1376;
	wire [3-1:0] node1380;
	wire [3-1:0] node1381;
	wire [3-1:0] node1382;
	wire [3-1:0] node1385;
	wire [3-1:0] node1388;
	wire [3-1:0] node1389;
	wire [3-1:0] node1392;
	wire [3-1:0] node1395;
	wire [3-1:0] node1396;
	wire [3-1:0] node1397;
	wire [3-1:0] node1398;
	wire [3-1:0] node1399;
	wire [3-1:0] node1401;
	wire [3-1:0] node1404;
	wire [3-1:0] node1405;
	wire [3-1:0] node1408;
	wire [3-1:0] node1411;
	wire [3-1:0] node1412;
	wire [3-1:0] node1413;
	wire [3-1:0] node1416;
	wire [3-1:0] node1419;
	wire [3-1:0] node1420;
	wire [3-1:0] node1424;
	wire [3-1:0] node1425;
	wire [3-1:0] node1426;
	wire [3-1:0] node1427;
	wire [3-1:0] node1432;
	wire [3-1:0] node1433;
	wire [3-1:0] node1434;
	wire [3-1:0] node1438;
	wire [3-1:0] node1440;
	wire [3-1:0] node1443;
	wire [3-1:0] node1444;
	wire [3-1:0] node1445;
	wire [3-1:0] node1446;
	wire [3-1:0] node1447;
	wire [3-1:0] node1450;
	wire [3-1:0] node1453;
	wire [3-1:0] node1454;
	wire [3-1:0] node1457;
	wire [3-1:0] node1460;
	wire [3-1:0] node1461;
	wire [3-1:0] node1462;
	wire [3-1:0] node1465;
	wire [3-1:0] node1468;
	wire [3-1:0] node1469;
	wire [3-1:0] node1472;
	wire [3-1:0] node1475;
	wire [3-1:0] node1476;
	wire [3-1:0] node1477;
	wire [3-1:0] node1478;
	wire [3-1:0] node1481;
	wire [3-1:0] node1484;
	wire [3-1:0] node1485;
	wire [3-1:0] node1488;
	wire [3-1:0] node1491;
	wire [3-1:0] node1492;
	wire [3-1:0] node1493;
	wire [3-1:0] node1496;
	wire [3-1:0] node1499;
	wire [3-1:0] node1500;
	wire [3-1:0] node1503;
	wire [3-1:0] node1506;
	wire [3-1:0] node1507;
	wire [3-1:0] node1509;
	wire [3-1:0] node1510;
	wire [3-1:0] node1511;
	wire [3-1:0] node1513;
	wire [3-1:0] node1514;
	wire [3-1:0] node1518;
	wire [3-1:0] node1519;
	wire [3-1:0] node1520;
	wire [3-1:0] node1526;
	wire [3-1:0] node1527;
	wire [3-1:0] node1529;
	wire [3-1:0] node1531;
	wire [3-1:0] node1532;
	wire [3-1:0] node1533;
	wire [3-1:0] node1536;
	wire [3-1:0] node1539;
	wire [3-1:0] node1541;
	wire [3-1:0] node1544;
	wire [3-1:0] node1545;
	wire [3-1:0] node1546;
	wire [3-1:0] node1547;
	wire [3-1:0] node1550;
	wire [3-1:0] node1551;
	wire [3-1:0] node1554;
	wire [3-1:0] node1557;
	wire [3-1:0] node1559;
	wire [3-1:0] node1560;
	wire [3-1:0] node1563;
	wire [3-1:0] node1566;
	wire [3-1:0] node1568;
	wire [3-1:0] node1569;
	wire [3-1:0] node1570;
	wire [3-1:0] node1574;
	wire [3-1:0] node1575;
	wire [3-1:0] node1578;

	assign outp = (inp[3]) ? node900 : node1;
		assign node1 = (inp[4]) ? node399 : node2;
			assign node2 = (inp[9]) ? node164 : node3;
				assign node3 = (inp[7]) ? node107 : node4;
					assign node4 = (inp[0]) ? node66 : node5;
						assign node5 = (inp[6]) ? node35 : node6;
							assign node6 = (inp[1]) ? node22 : node7;
								assign node7 = (inp[10]) ? node15 : node8;
									assign node8 = (inp[2]) ? node12 : node9;
										assign node9 = (inp[5]) ? 3'b001 : 3'b001;
										assign node12 = (inp[8]) ? 3'b001 : 3'b101;
									assign node15 = (inp[11]) ? node19 : node16;
										assign node16 = (inp[5]) ? 3'b001 : 3'b101;
										assign node19 = (inp[5]) ? 3'b110 : 3'b001;
								assign node22 = (inp[8]) ? node28 : node23;
									assign node23 = (inp[5]) ? 3'b001 : node24;
										assign node24 = (inp[11]) ? 3'b111 : 3'b001;
									assign node28 = (inp[2]) ? node32 : node29;
										assign node29 = (inp[10]) ? 3'b101 : 3'b001;
										assign node32 = (inp[5]) ? 3'b001 : 3'b111;
							assign node35 = (inp[10]) ? node51 : node36;
								assign node36 = (inp[5]) ? node44 : node37;
									assign node37 = (inp[11]) ? node41 : node38;
										assign node38 = (inp[8]) ? 3'b001 : 3'b001;
										assign node41 = (inp[1]) ? 3'b101 : 3'b011;
									assign node44 = (inp[11]) ? node48 : node45;
										assign node45 = (inp[8]) ? 3'b111 : 3'b011;
										assign node48 = (inp[1]) ? 3'b011 : 3'b011;
								assign node51 = (inp[5]) ? node59 : node52;
									assign node52 = (inp[11]) ? node56 : node53;
										assign node53 = (inp[1]) ? 3'b011 : 3'b111;
										assign node56 = (inp[1]) ? 3'b111 : 3'b011;
									assign node59 = (inp[1]) ? node63 : node60;
										assign node60 = (inp[11]) ? 3'b101 : 3'b011;
										assign node63 = (inp[11]) ? 3'b011 : 3'b111;
						assign node66 = (inp[1]) ? node90 : node67;
							assign node67 = (inp[5]) ? node77 : node68;
								assign node68 = (inp[2]) ? node72 : node69;
									assign node69 = (inp[8]) ? 3'b111 : 3'b011;
									assign node72 = (inp[8]) ? node74 : 3'b111;
										assign node74 = (inp[11]) ? 3'b111 : 3'b011;
								assign node77 = (inp[11]) ? node85 : node78;
									assign node78 = (inp[6]) ? node82 : node79;
										assign node79 = (inp[2]) ? 3'b001 : 3'b001;
										assign node82 = (inp[10]) ? 3'b001 : 3'b001;
									assign node85 = (inp[2]) ? 3'b101 : node86;
										assign node86 = (inp[8]) ? 3'b101 : 3'b001;
							assign node90 = (inp[6]) ? 3'b111 : node91;
								assign node91 = (inp[5]) ? node99 : node92;
									assign node92 = (inp[8]) ? node96 : node93;
										assign node93 = (inp[2]) ? 3'b111 : 3'b011;
										assign node96 = (inp[11]) ? 3'b111 : 3'b011;
									assign node99 = (inp[2]) ? node103 : node100;
										assign node100 = (inp[8]) ? 3'b011 : 3'b011;
										assign node103 = (inp[8]) ? 3'b111 : 3'b011;
					assign node107 = (inp[5]) ? node131 : node108;
						assign node108 = (inp[2]) ? node118 : node109;
							assign node109 = (inp[8]) ? 3'b111 : node110;
								assign node110 = (inp[1]) ? node112 : 3'b111;
									assign node112 = (inp[11]) ? node114 : 3'b111;
										assign node114 = (inp[6]) ? 3'b111 : 3'b011;
							assign node118 = (inp[11]) ? 3'b111 : node119;
								assign node119 = (inp[0]) ? node125 : node120;
									assign node120 = (inp[8]) ? node122 : 3'b111;
										assign node122 = (inp[6]) ? 3'b101 : 3'b001;
									assign node125 = (inp[6]) ? 3'b111 : node126;
										assign node126 = (inp[1]) ? 3'b011 : 3'b111;
						assign node131 = (inp[0]) ? node153 : node132;
							assign node132 = (inp[6]) ? node146 : node133;
								assign node133 = (inp[1]) ? node139 : node134;
									assign node134 = (inp[8]) ? 3'b111 : node135;
										assign node135 = (inp[2]) ? 3'b111 : 3'b101;
									assign node139 = (inp[11]) ? node143 : node140;
										assign node140 = (inp[8]) ? 3'b011 : 3'b011;
										assign node143 = (inp[2]) ? 3'b011 : 3'b101;
								assign node146 = (inp[11]) ? node148 : 3'b111;
									assign node148 = (inp[2]) ? 3'b111 : node149;
										assign node149 = (inp[8]) ? 3'b111 : 3'b101;
							assign node153 = (inp[1]) ? node155 : 3'b011;
								assign node155 = (inp[6]) ? 3'b111 : node156;
									assign node156 = (inp[11]) ? node160 : node157;
										assign node157 = (inp[2]) ? 3'b011 : 3'b011;
										assign node160 = (inp[2]) ? 3'b011 : 3'b111;
				assign node164 = (inp[6]) ? node288 : node165;
					assign node165 = (inp[0]) ? node225 : node166;
						assign node166 = (inp[5]) ? node196 : node167;
							assign node167 = (inp[10]) ? node181 : node168;
								assign node168 = (inp[1]) ? node176 : node169;
									assign node169 = (inp[7]) ? node173 : node170;
										assign node170 = (inp[8]) ? 3'b001 : 3'b110;
										assign node173 = (inp[11]) ? 3'b001 : 3'b101;
									assign node176 = (inp[2]) ? 3'b101 : node177;
										assign node177 = (inp[7]) ? 3'b101 : 3'b001;
								assign node181 = (inp[7]) ? node189 : node182;
									assign node182 = (inp[11]) ? node186 : node183;
										assign node183 = (inp[1]) ? 3'b001 : 3'b110;
										assign node186 = (inp[1]) ? 3'b110 : 3'b010;
									assign node189 = (inp[1]) ? node193 : node190;
										assign node190 = (inp[11]) ? 3'b110 : 3'b001;
										assign node193 = (inp[8]) ? 3'b001 : 3'b001;
							assign node196 = (inp[10]) ? node212 : node197;
								assign node197 = (inp[11]) ? node205 : node198;
									assign node198 = (inp[1]) ? node202 : node199;
										assign node199 = (inp[7]) ? 3'b001 : 3'b110;
										assign node202 = (inp[2]) ? 3'b001 : 3'b001;
									assign node205 = (inp[7]) ? node209 : node206;
										assign node206 = (inp[1]) ? 3'b110 : 3'b010;
										assign node209 = (inp[8]) ? 3'b001 : 3'b110;
								assign node212 = (inp[7]) ? node218 : node213;
									assign node213 = (inp[1]) ? 3'b010 : node214;
										assign node214 = (inp[2]) ? 3'b010 : 3'b100;
									assign node218 = (inp[1]) ? node222 : node219;
										assign node219 = (inp[11]) ? 3'b010 : 3'b110;
										assign node222 = (inp[2]) ? 3'b110 : 3'b110;
						assign node225 = (inp[10]) ? node257 : node226;
							assign node226 = (inp[7]) ? node242 : node227;
								assign node227 = (inp[1]) ? node235 : node228;
									assign node228 = (inp[5]) ? node232 : node229;
										assign node229 = (inp[11]) ? 3'b101 : 3'b101;
										assign node232 = (inp[2]) ? 3'b001 : 3'b001;
									assign node235 = (inp[5]) ? node239 : node236;
										assign node236 = (inp[8]) ? 3'b011 : 3'b001;
										assign node239 = (inp[2]) ? 3'b101 : 3'b101;
								assign node242 = (inp[5]) ? node250 : node243;
									assign node243 = (inp[1]) ? node247 : node244;
										assign node244 = (inp[2]) ? 3'b011 : 3'b001;
										assign node247 = (inp[11]) ? 3'b011 : 3'b111;
									assign node250 = (inp[8]) ? node254 : node251;
										assign node251 = (inp[2]) ? 3'b101 : 3'b101;
										assign node254 = (inp[1]) ? 3'b011 : 3'b101;
							assign node257 = (inp[5]) ? node273 : node258;
								assign node258 = (inp[2]) ? node266 : node259;
									assign node259 = (inp[1]) ? node263 : node260;
										assign node260 = (inp[7]) ? 3'b101 : 3'b001;
										assign node263 = (inp[8]) ? 3'b101 : 3'b101;
									assign node266 = (inp[7]) ? node270 : node267;
										assign node267 = (inp[11]) ? 3'b001 : 3'b101;
										assign node270 = (inp[11]) ? 3'b101 : 3'b011;
								assign node273 = (inp[7]) ? node281 : node274;
									assign node274 = (inp[1]) ? node278 : node275;
										assign node275 = (inp[8]) ? 3'b110 : 3'b110;
										assign node278 = (inp[11]) ? 3'b110 : 3'b001;
									assign node281 = (inp[8]) ? node285 : node282;
										assign node282 = (inp[1]) ? 3'b001 : 3'b110;
										assign node285 = (inp[1]) ? 3'b101 : 3'b001;
					assign node288 = (inp[0]) ? node348 : node289;
						assign node289 = (inp[7]) ? node317 : node290;
							assign node290 = (inp[5]) ? node304 : node291;
								assign node291 = (inp[1]) ? node297 : node292;
									assign node292 = (inp[10]) ? node294 : 3'b101;
										assign node294 = (inp[8]) ? 3'b001 : 3'b001;
									assign node297 = (inp[10]) ? node301 : node298;
										assign node298 = (inp[8]) ? 3'b011 : 3'b011;
										assign node301 = (inp[2]) ? 3'b101 : 3'b101;
								assign node304 = (inp[1]) ? node310 : node305;
									assign node305 = (inp[10]) ? node307 : 3'b001;
										assign node307 = (inp[11]) ? 3'b110 : 3'b110;
									assign node310 = (inp[10]) ? node314 : node311;
										assign node311 = (inp[8]) ? 3'b001 : 3'b101;
										assign node314 = (inp[2]) ? 3'b001 : 3'b001;
							assign node317 = (inp[5]) ? node333 : node318;
								assign node318 = (inp[10]) ? node326 : node319;
									assign node319 = (inp[1]) ? node323 : node320;
										assign node320 = (inp[2]) ? 3'b011 : 3'b011;
										assign node323 = (inp[2]) ? 3'b001 : 3'b111;
									assign node326 = (inp[8]) ? node330 : node327;
										assign node327 = (inp[11]) ? 3'b101 : 3'b001;
										assign node330 = (inp[1]) ? 3'b011 : 3'b001;
								assign node333 = (inp[10]) ? node341 : node334;
									assign node334 = (inp[1]) ? node338 : node335;
										assign node335 = (inp[8]) ? 3'b101 : 3'b101;
										assign node338 = (inp[11]) ? 3'b011 : 3'b011;
									assign node341 = (inp[11]) ? node345 : node342;
										assign node342 = (inp[1]) ? 3'b101 : 3'b001;
										assign node345 = (inp[2]) ? 3'b001 : 3'b001;
						assign node348 = (inp[7]) ? node378 : node349;
							assign node349 = (inp[1]) ? node365 : node350;
								assign node350 = (inp[10]) ? node358 : node351;
									assign node351 = (inp[11]) ? node355 : node352;
										assign node352 = (inp[5]) ? 3'b011 : 3'b011;
										assign node355 = (inp[5]) ? 3'b101 : 3'b011;
									assign node358 = (inp[5]) ? node362 : node359;
										assign node359 = (inp[2]) ? 3'b011 : 3'b101;
										assign node362 = (inp[11]) ? 3'b001 : 3'b101;
								assign node365 = (inp[11]) ? node371 : node366;
									assign node366 = (inp[10]) ? node368 : 3'b111;
										assign node368 = (inp[5]) ? 3'b011 : 3'b111;
									assign node371 = (inp[5]) ? node375 : node372;
										assign node372 = (inp[8]) ? 3'b011 : 3'b011;
										assign node375 = (inp[10]) ? 3'b101 : 3'b011;
							assign node378 = (inp[10]) ? node386 : node379;
								assign node379 = (inp[5]) ? node381 : 3'b111;
									assign node381 = (inp[1]) ? 3'b111 : node382;
										assign node382 = (inp[2]) ? 3'b111 : 3'b011;
								assign node386 = (inp[5]) ? node392 : node387;
									assign node387 = (inp[1]) ? 3'b111 : node388;
										assign node388 = (inp[2]) ? 3'b111 : 3'b011;
									assign node392 = (inp[1]) ? node396 : node393;
										assign node393 = (inp[11]) ? 3'b101 : 3'b011;
										assign node396 = (inp[8]) ? 3'b011 : 3'b011;
			assign node399 = (inp[0]) ? node647 : node400;
				assign node400 = (inp[9]) ? node528 : node401;
					assign node401 = (inp[11]) ? node465 : node402;
						assign node402 = (inp[5]) ? node434 : node403;
							assign node403 = (inp[2]) ? node419 : node404;
								assign node404 = (inp[1]) ? node412 : node405;
									assign node405 = (inp[10]) ? node409 : node406;
										assign node406 = (inp[7]) ? 3'b001 : 3'b001;
										assign node409 = (inp[6]) ? 3'b101 : 3'b101;
									assign node412 = (inp[10]) ? node416 : node413;
										assign node413 = (inp[8]) ? 3'b101 : 3'b001;
										assign node416 = (inp[6]) ? 3'b001 : 3'b001;
								assign node419 = (inp[10]) ? node427 : node420;
									assign node420 = (inp[1]) ? node424 : node421;
										assign node421 = (inp[7]) ? 3'b101 : 3'b000;
										assign node424 = (inp[7]) ? 3'b110 : 3'b101;
									assign node427 = (inp[1]) ? node431 : node428;
										assign node428 = (inp[7]) ? 3'b001 : 3'b110;
										assign node431 = (inp[7]) ? 3'b011 : 3'b001;
							assign node434 = (inp[7]) ? node450 : node435;
								assign node435 = (inp[1]) ? node443 : node436;
									assign node436 = (inp[6]) ? node440 : node437;
										assign node437 = (inp[10]) ? 3'b010 : 3'b110;
										assign node440 = (inp[10]) ? 3'b000 : 3'b101;
									assign node443 = (inp[10]) ? node447 : node444;
										assign node444 = (inp[2]) ? 3'b010 : 3'b010;
										assign node447 = (inp[2]) ? 3'b110 : 3'b010;
								assign node450 = (inp[1]) ? node458 : node451;
									assign node451 = (inp[10]) ? node455 : node452;
										assign node452 = (inp[8]) ? 3'b001 : 3'b101;
										assign node455 = (inp[6]) ? 3'b001 : 3'b101;
									assign node458 = (inp[10]) ? node462 : node459;
										assign node459 = (inp[2]) ? 3'b011 : 3'b001;
										assign node462 = (inp[6]) ? 3'b101 : 3'b110;
						assign node465 = (inp[6]) ? node497 : node466;
							assign node466 = (inp[1]) ? node482 : node467;
								assign node467 = (inp[5]) ? node475 : node468;
									assign node468 = (inp[7]) ? node472 : node469;
										assign node469 = (inp[10]) ? 3'b010 : 3'b110;
										assign node472 = (inp[10]) ? 3'b110 : 3'b010;
									assign node475 = (inp[7]) ? node479 : node476;
										assign node476 = (inp[10]) ? 3'b100 : 3'b010;
										assign node479 = (inp[8]) ? 3'b110 : 3'b110;
								assign node482 = (inp[7]) ? node490 : node483;
									assign node483 = (inp[5]) ? node487 : node484;
										assign node484 = (inp[10]) ? 3'b110 : 3'b010;
										assign node487 = (inp[10]) ? 3'b010 : 3'b110;
									assign node490 = (inp[10]) ? node494 : node491;
										assign node491 = (inp[5]) ? 3'b000 : 3'b101;
										assign node494 = (inp[5]) ? 3'b110 : 3'b000;
							assign node497 = (inp[8]) ? node513 : node498;
								assign node498 = (inp[7]) ? node506 : node499;
									assign node499 = (inp[1]) ? node503 : node500;
										assign node500 = (inp[5]) ? 3'b000 : 3'b001;
										assign node503 = (inp[5]) ? 3'b010 : 3'b010;
									assign node506 = (inp[1]) ? node510 : node507;
										assign node507 = (inp[10]) ? 3'b010 : 3'b010;
										assign node510 = (inp[2]) ? 3'b001 : 3'b000;
								assign node513 = (inp[2]) ? node521 : node514;
									assign node514 = (inp[7]) ? node518 : node515;
										assign node515 = (inp[1]) ? 3'b010 : 3'b001;
										assign node518 = (inp[1]) ? 3'b001 : 3'b010;
									assign node521 = (inp[5]) ? node525 : node522;
										assign node522 = (inp[1]) ? 3'b110 : 3'b111;
										assign node525 = (inp[10]) ? 3'b010 : 3'b110;
					assign node528 = (inp[6]) ? node584 : node529;
						assign node529 = (inp[10]) ? node559 : node530;
							assign node530 = (inp[1]) ? node546 : node531;
								assign node531 = (inp[8]) ? node539 : node532;
									assign node532 = (inp[5]) ? node536 : node533;
										assign node533 = (inp[11]) ? 3'b100 : 3'b100;
										assign node536 = (inp[7]) ? 3'b100 : 3'b000;
									assign node539 = (inp[7]) ? node543 : node540;
										assign node540 = (inp[5]) ? 3'b100 : 3'b010;
										assign node543 = (inp[11]) ? 3'b000 : 3'b010;
								assign node546 = (inp[5]) ? node552 : node547;
									assign node547 = (inp[7]) ? node549 : 3'b010;
										assign node549 = (inp[11]) ? 3'b110 : 3'b010;
									assign node552 = (inp[7]) ? node556 : node553;
										assign node553 = (inp[11]) ? 3'b100 : 3'b100;
										assign node556 = (inp[8]) ? 3'b010 : 3'b010;
							assign node559 = (inp[5]) ? node575 : node560;
								assign node560 = (inp[7]) ? node568 : node561;
									assign node561 = (inp[11]) ? node565 : node562;
										assign node562 = (inp[1]) ? 3'b100 : 3'b100;
										assign node565 = (inp[1]) ? 3'b100 : 3'b000;
									assign node568 = (inp[1]) ? node572 : node569;
										assign node569 = (inp[8]) ? 3'b100 : 3'b100;
										assign node572 = (inp[11]) ? 3'b010 : 3'b010;
								assign node575 = (inp[1]) ? node577 : 3'b000;
									assign node577 = (inp[7]) ? node581 : node578;
										assign node578 = (inp[2]) ? 3'b000 : 3'b000;
										assign node581 = (inp[11]) ? 3'b100 : 3'b100;
						assign node584 = (inp[5]) ? node616 : node585;
							assign node585 = (inp[10]) ? node601 : node586;
								assign node586 = (inp[8]) ? node594 : node587;
									assign node587 = (inp[7]) ? node591 : node588;
										assign node588 = (inp[1]) ? 3'b111 : 3'b110;
										assign node591 = (inp[2]) ? 3'b001 : 3'b010;
									assign node594 = (inp[1]) ? node598 : node595;
										assign node595 = (inp[7]) ? 3'b001 : 3'b110;
										assign node598 = (inp[7]) ? 3'b101 : 3'b001;
								assign node601 = (inp[7]) ? node609 : node602;
									assign node602 = (inp[1]) ? node606 : node603;
										assign node603 = (inp[11]) ? 3'b010 : 3'b010;
										assign node606 = (inp[2]) ? 3'b110 : 3'b110;
									assign node609 = (inp[1]) ? node613 : node610;
										assign node610 = (inp[2]) ? 3'b110 : 3'b110;
										assign node613 = (inp[11]) ? 3'b110 : 3'b001;
							assign node616 = (inp[7]) ? node632 : node617;
								assign node617 = (inp[10]) ? node625 : node618;
									assign node618 = (inp[8]) ? node622 : node619;
										assign node619 = (inp[1]) ? 3'b110 : 3'b010;
										assign node622 = (inp[1]) ? 3'b000 : 3'b010;
									assign node625 = (inp[1]) ? node629 : node626;
										assign node626 = (inp[8]) ? 3'b100 : 3'b100;
										assign node629 = (inp[11]) ? 3'b100 : 3'b010;
								assign node632 = (inp[10]) ? node640 : node633;
									assign node633 = (inp[2]) ? node637 : node634;
										assign node634 = (inp[1]) ? 3'b110 : 3'b110;
										assign node637 = (inp[1]) ? 3'b001 : 3'b110;
									assign node640 = (inp[2]) ? node644 : node641;
										assign node641 = (inp[1]) ? 3'b010 : 3'b010;
										assign node644 = (inp[11]) ? 3'b010 : 3'b110;
				assign node647 = (inp[9]) ? node773 : node648;
					assign node648 = (inp[7]) ? node710 : node649;
						assign node649 = (inp[6]) ? node681 : node650;
							assign node650 = (inp[5]) ? node666 : node651;
								assign node651 = (inp[1]) ? node659 : node652;
									assign node652 = (inp[10]) ? node656 : node653;
										assign node653 = (inp[8]) ? 3'b101 : 3'b001;
										assign node656 = (inp[8]) ? 3'b001 : 3'b001;
									assign node659 = (inp[8]) ? node663 : node660;
										assign node660 = (inp[11]) ? 3'b001 : 3'b101;
										assign node663 = (inp[11]) ? 3'b101 : 3'b011;
								assign node666 = (inp[10]) ? node674 : node667;
									assign node667 = (inp[1]) ? node671 : node668;
										assign node668 = (inp[8]) ? 3'b011 : 3'b011;
										assign node671 = (inp[11]) ? 3'b100 : 3'b001;
									assign node674 = (inp[1]) ? node678 : node675;
										assign node675 = (inp[2]) ? 3'b000 : 3'b110;
										assign node678 = (inp[11]) ? 3'b110 : 3'b001;
							assign node681 = (inp[5]) ? node697 : node682;
								assign node682 = (inp[1]) ? node690 : node683;
									assign node683 = (inp[11]) ? node687 : node684;
										assign node684 = (inp[8]) ? 3'b000 : 3'b000;
										assign node687 = (inp[2]) ? 3'b100 : 3'b101;
									assign node690 = (inp[11]) ? node694 : node691;
										assign node691 = (inp[8]) ? 3'b001 : 3'b101;
										assign node694 = (inp[2]) ? 3'b011 : 3'b011;
								assign node697 = (inp[1]) ? node705 : node698;
									assign node698 = (inp[2]) ? node702 : node699;
										assign node699 = (inp[11]) ? 3'b101 : 3'b011;
										assign node702 = (inp[8]) ? 3'b001 : 3'b011;
									assign node705 = (inp[2]) ? node707 : 3'b101;
										assign node707 = (inp[8]) ? 3'b011 : 3'b101;
						assign node710 = (inp[5]) ? node742 : node711;
							assign node711 = (inp[1]) ? node727 : node712;
								assign node712 = (inp[10]) ? node720 : node713;
									assign node713 = (inp[6]) ? node717 : node714;
										assign node714 = (inp[11]) ? 3'b011 : 3'b011;
										assign node717 = (inp[11]) ? 3'b111 : 3'b011;
									assign node720 = (inp[11]) ? node724 : node721;
										assign node721 = (inp[2]) ? 3'b111 : 3'b111;
										assign node724 = (inp[8]) ? 3'b111 : 3'b000;
								assign node727 = (inp[10]) ? node735 : node728;
									assign node728 = (inp[11]) ? node732 : node729;
										assign node729 = (inp[6]) ? 3'b101 : 3'b111;
										assign node732 = (inp[6]) ? 3'b001 : 3'b011;
									assign node735 = (inp[11]) ? node739 : node736;
										assign node736 = (inp[6]) ? 3'b011 : 3'b011;
										assign node739 = (inp[6]) ? 3'b111 : 3'b101;
							assign node742 = (inp[1]) ? node758 : node743;
								assign node743 = (inp[10]) ? node751 : node744;
									assign node744 = (inp[11]) ? node748 : node745;
										assign node745 = (inp[2]) ? 3'b101 : 3'b101;
										assign node748 = (inp[2]) ? 3'b101 : 3'b010;
									assign node751 = (inp[11]) ? node755 : node752;
										assign node752 = (inp[8]) ? 3'b001 : 3'b001;
										assign node755 = (inp[8]) ? 3'b001 : 3'b100;
								assign node758 = (inp[10]) ? node766 : node759;
									assign node759 = (inp[11]) ? node763 : node760;
										assign node760 = (inp[8]) ? 3'b011 : 3'b011;
										assign node763 = (inp[8]) ? 3'b111 : 3'b111;
									assign node766 = (inp[6]) ? node770 : node767;
										assign node767 = (inp[2]) ? 3'b101 : 3'b001;
										assign node770 = (inp[11]) ? 3'b011 : 3'b111;
					assign node773 = (inp[6]) ? node837 : node774;
						assign node774 = (inp[10]) ? node806 : node775;
							assign node775 = (inp[7]) ? node791 : node776;
								assign node776 = (inp[5]) ? node784 : node777;
									assign node777 = (inp[11]) ? node781 : node778;
										assign node778 = (inp[1]) ? 3'b001 : 3'b110;
										assign node781 = (inp[2]) ? 3'b110 : 3'b110;
									assign node784 = (inp[11]) ? node788 : node785;
										assign node785 = (inp[1]) ? 3'b110 : 3'b010;
										assign node788 = (inp[2]) ? 3'b010 : 3'b010;
								assign node791 = (inp[1]) ? node799 : node792;
									assign node792 = (inp[5]) ? node796 : node793;
										assign node793 = (inp[11]) ? 3'b001 : 3'b001;
										assign node796 = (inp[2]) ? 3'b110 : 3'b110;
									assign node799 = (inp[2]) ? node803 : node800;
										assign node800 = (inp[8]) ? 3'b001 : 3'b000;
										assign node803 = (inp[5]) ? 3'b001 : 3'b101;
							assign node806 = (inp[5]) ? node822 : node807;
								assign node807 = (inp[1]) ? node815 : node808;
									assign node808 = (inp[11]) ? node812 : node809;
										assign node809 = (inp[7]) ? 3'b110 : 3'b010;
										assign node812 = (inp[7]) ? 3'b010 : 3'b100;
									assign node815 = (inp[7]) ? node819 : node816;
										assign node816 = (inp[11]) ? 3'b010 : 3'b110;
										assign node819 = (inp[8]) ? 3'b001 : 3'b110;
								assign node822 = (inp[1]) ? node830 : node823;
									assign node823 = (inp[7]) ? node827 : node824;
										assign node824 = (inp[2]) ? 3'b100 : 3'b100;
										assign node827 = (inp[8]) ? 3'b010 : 3'b100;
									assign node830 = (inp[7]) ? node834 : node831;
										assign node831 = (inp[8]) ? 3'b010 : 3'b100;
										assign node834 = (inp[8]) ? 3'b110 : 3'b010;
						assign node837 = (inp[7]) ? node869 : node838;
							assign node838 = (inp[1]) ? node854 : node839;
								assign node839 = (inp[5]) ? node847 : node840;
									assign node840 = (inp[8]) ? node844 : node841;
										assign node841 = (inp[10]) ? 3'b110 : 3'b011;
										assign node844 = (inp[10]) ? 3'b001 : 3'b101;
									assign node847 = (inp[10]) ? node851 : node848;
										assign node848 = (inp[11]) ? 3'b111 : 3'b011;
										assign node851 = (inp[2]) ? 3'b110 : 3'b010;
								assign node854 = (inp[10]) ? node862 : node855;
									assign node855 = (inp[5]) ? node859 : node856;
										assign node856 = (inp[11]) ? 3'b101 : 3'b011;
										assign node859 = (inp[8]) ? 3'b001 : 3'b001;
									assign node862 = (inp[5]) ? node866 : node863;
										assign node863 = (inp[11]) ? 3'b001 : 3'b100;
										assign node866 = (inp[11]) ? 3'b110 : 3'b001;
							assign node869 = (inp[10]) ? node885 : node870;
								assign node870 = (inp[5]) ? node878 : node871;
									assign node871 = (inp[1]) ? node875 : node872;
										assign node872 = (inp[8]) ? 3'b011 : 3'b101;
										assign node875 = (inp[8]) ? 3'b011 : 3'b011;
									assign node878 = (inp[8]) ? node882 : node879;
										assign node879 = (inp[11]) ? 3'b001 : 3'b101;
										assign node882 = (inp[1]) ? 3'b101 : 3'b101;
								assign node885 = (inp[5]) ? node893 : node886;
									assign node886 = (inp[1]) ? node890 : node887;
										assign node887 = (inp[11]) ? 3'b001 : 3'b101;
										assign node890 = (inp[2]) ? 3'b101 : 3'b101;
									assign node893 = (inp[1]) ? node897 : node894;
										assign node894 = (inp[11]) ? 3'b110 : 3'b000;
										assign node897 = (inp[8]) ? 3'b001 : 3'b001;
		assign node900 = (inp[4]) ? node1330 : node901;
			assign node901 = (inp[9]) ? node1137 : node902;
				assign node902 = (inp[6]) ? node1010 : node903;
					assign node903 = (inp[0]) ? node953 : node904;
						assign node904 = (inp[7]) ? node928 : node905;
							assign node905 = (inp[5]) ? node919 : node906;
								assign node906 = (inp[10]) ? node914 : node907;
									assign node907 = (inp[1]) ? node911 : node908;
										assign node908 = (inp[8]) ? 3'b000 : 3'b100;
										assign node911 = (inp[11]) ? 3'b010 : 3'b100;
									assign node914 = (inp[1]) ? 3'b100 : node915;
										assign node915 = (inp[11]) ? 3'b000 : 3'b100;
								assign node919 = (inp[10]) ? 3'b000 : node920;
									assign node920 = (inp[1]) ? node924 : node921;
										assign node921 = (inp[11]) ? 3'b000 : 3'b100;
										assign node924 = (inp[11]) ? 3'b100 : 3'b010;
							assign node928 = (inp[11]) ? node940 : node929;
								assign node929 = (inp[8]) ? node933 : node930;
									assign node930 = (inp[1]) ? 3'b110 : 3'b100;
									assign node933 = (inp[1]) ? node937 : node934;
										assign node934 = (inp[2]) ? 3'b000 : 3'b010;
										assign node937 = (inp[5]) ? 3'b110 : 3'b010;
								assign node940 = (inp[1]) ? node946 : node941;
									assign node941 = (inp[5]) ? 3'b100 : node942;
										assign node942 = (inp[10]) ? 3'b100 : 3'b110;
									assign node946 = (inp[5]) ? node950 : node947;
										assign node947 = (inp[8]) ? 3'b000 : 3'b100;
										assign node950 = (inp[2]) ? 3'b000 : 3'b000;
						assign node953 = (inp[7]) ? node979 : node954;
							assign node954 = (inp[1]) ? node970 : node955;
								assign node955 = (inp[10]) ? node963 : node956;
									assign node956 = (inp[5]) ? node960 : node957;
										assign node957 = (inp[8]) ? 3'b110 : 3'b010;
										assign node960 = (inp[2]) ? 3'b010 : 3'b010;
									assign node963 = (inp[5]) ? node967 : node964;
										assign node964 = (inp[2]) ? 3'b010 : 3'b010;
										assign node967 = (inp[2]) ? 3'b100 : 3'b100;
								assign node970 = (inp[10]) ? node972 : 3'b110;
									assign node972 = (inp[5]) ? node976 : node973;
										assign node973 = (inp[8]) ? 3'b110 : 3'b010;
										assign node976 = (inp[11]) ? 3'b100 : 3'b010;
							assign node979 = (inp[1]) ? node995 : node980;
								assign node980 = (inp[2]) ? node988 : node981;
									assign node981 = (inp[8]) ? node985 : node982;
										assign node982 = (inp[5]) ? 3'b000 : 3'b010;
										assign node985 = (inp[11]) ? 3'b100 : 3'b110;
									assign node988 = (inp[8]) ? node992 : node989;
										assign node989 = (inp[11]) ? 3'b100 : 3'b110;
										assign node992 = (inp[11]) ? 3'b110 : 3'b010;
								assign node995 = (inp[5]) ? node1003 : node996;
									assign node996 = (inp[8]) ? node1000 : node997;
										assign node997 = (inp[10]) ? 3'b100 : 3'b101;
										assign node1000 = (inp[10]) ? 3'b001 : 3'b011;
									assign node1003 = (inp[10]) ? node1007 : node1004;
										assign node1004 = (inp[11]) ? 3'b110 : 3'b001;
										assign node1007 = (inp[11]) ? 3'b010 : 3'b110;
					assign node1010 = (inp[0]) ? node1074 : node1011;
						assign node1011 = (inp[7]) ? node1043 : node1012;
							assign node1012 = (inp[1]) ? node1028 : node1013;
								assign node1013 = (inp[8]) ? node1021 : node1014;
									assign node1014 = (inp[5]) ? node1018 : node1015;
										assign node1015 = (inp[10]) ? 3'b000 : 3'b100;
										assign node1018 = (inp[10]) ? 3'b100 : 3'b000;
									assign node1021 = (inp[2]) ? node1025 : node1022;
										assign node1022 = (inp[5]) ? 3'b000 : 3'b000;
										assign node1025 = (inp[5]) ? 3'b000 : 3'b000;
								assign node1028 = (inp[10]) ? node1036 : node1029;
									assign node1029 = (inp[5]) ? node1033 : node1030;
										assign node1030 = (inp[8]) ? 3'b000 : 3'b000;
										assign node1033 = (inp[8]) ? 3'b110 : 3'b110;
									assign node1036 = (inp[5]) ? node1040 : node1037;
										assign node1037 = (inp[2]) ? 3'b110 : 3'b110;
										assign node1040 = (inp[2]) ? 3'b010 : 3'b010;
							assign node1043 = (inp[10]) ? node1059 : node1044;
								assign node1044 = (inp[1]) ? node1052 : node1045;
									assign node1045 = (inp[5]) ? node1049 : node1046;
										assign node1046 = (inp[8]) ? 3'b001 : 3'b100;
										assign node1049 = (inp[11]) ? 3'b110 : 3'b110;
									assign node1052 = (inp[8]) ? node1056 : node1053;
										assign node1053 = (inp[11]) ? 3'b000 : 3'b101;
										assign node1056 = (inp[11]) ? 3'b001 : 3'b011;
								assign node1059 = (inp[8]) ? node1067 : node1060;
									assign node1060 = (inp[1]) ? node1064 : node1061;
										assign node1061 = (inp[11]) ? 3'b110 : 3'b110;
										assign node1064 = (inp[11]) ? 3'b010 : 3'b110;
									assign node1067 = (inp[5]) ? node1071 : node1068;
										assign node1068 = (inp[11]) ? 3'b110 : 3'b011;
										assign node1071 = (inp[2]) ? 3'b110 : 3'b010;
						assign node1074 = (inp[1]) ? node1106 : node1075;
							assign node1075 = (inp[7]) ? node1091 : node1076;
								assign node1076 = (inp[11]) ? node1084 : node1077;
									assign node1077 = (inp[5]) ? node1081 : node1078;
										assign node1078 = (inp[10]) ? 3'b001 : 3'b000;
										assign node1081 = (inp[10]) ? 3'b110 : 3'b001;
									assign node1084 = (inp[2]) ? node1088 : node1085;
										assign node1085 = (inp[10]) ? 3'b110 : 3'b110;
										assign node1088 = (inp[8]) ? 3'b001 : 3'b010;
								assign node1091 = (inp[10]) ? node1099 : node1092;
									assign node1092 = (inp[5]) ? node1096 : node1093;
										assign node1093 = (inp[8]) ? 3'b010 : 3'b101;
										assign node1096 = (inp[2]) ? 3'b101 : 3'b001;
									assign node1099 = (inp[5]) ? node1103 : node1100;
										assign node1100 = (inp[11]) ? 3'b001 : 3'b101;
										assign node1103 = (inp[11]) ? 3'b110 : 3'b001;
							assign node1106 = (inp[7]) ? node1122 : node1107;
								assign node1107 = (inp[10]) ? node1115 : node1108;
									assign node1108 = (inp[5]) ? node1112 : node1109;
										assign node1109 = (inp[8]) ? 3'b011 : 3'b101;
										assign node1112 = (inp[8]) ? 3'b101 : 3'b001;
									assign node1115 = (inp[8]) ? node1119 : node1116;
										assign node1116 = (inp[11]) ? 3'b001 : 3'b000;
										assign node1119 = (inp[5]) ? 3'b001 : 3'b100;
								assign node1122 = (inp[5]) ? node1130 : node1123;
									assign node1123 = (inp[11]) ? node1127 : node1124;
										assign node1124 = (inp[10]) ? 3'b011 : 3'b111;
										assign node1127 = (inp[10]) ? 3'b101 : 3'b011;
									assign node1130 = (inp[10]) ? node1134 : node1131;
										assign node1131 = (inp[11]) ? 3'b101 : 3'b011;
										assign node1134 = (inp[11]) ? 3'b001 : 3'b001;
				assign node1137 = (inp[6]) ? node1213 : node1138;
					assign node1138 = (inp[0]) ? node1162 : node1139;
						assign node1139 = (inp[1]) ? node1141 : 3'b000;
							assign node1141 = (inp[10]) ? node1155 : node1142;
								assign node1142 = (inp[7]) ? node1148 : node1143;
									assign node1143 = (inp[11]) ? 3'b000 : node1144;
										assign node1144 = (inp[2]) ? 3'b000 : 3'b000;
									assign node1148 = (inp[5]) ? node1152 : node1149;
										assign node1149 = (inp[8]) ? 3'b100 : 3'b100;
										assign node1152 = (inp[8]) ? 3'b000 : 3'b000;
								assign node1155 = (inp[5]) ? 3'b000 : node1156;
									assign node1156 = (inp[8]) ? node1158 : 3'b000;
										assign node1158 = (inp[11]) ? 3'b000 : 3'b000;
						assign node1162 = (inp[5]) ? node1192 : node1163;
							assign node1163 = (inp[10]) ? node1179 : node1164;
								assign node1164 = (inp[7]) ? node1172 : node1165;
									assign node1165 = (inp[11]) ? node1169 : node1166;
										assign node1166 = (inp[2]) ? 3'b010 : 3'b100;
										assign node1169 = (inp[2]) ? 3'b100 : 3'b100;
									assign node1172 = (inp[1]) ? node1176 : node1173;
										assign node1173 = (inp[11]) ? 3'b100 : 3'b010;
										assign node1176 = (inp[11]) ? 3'b010 : 3'b110;
								assign node1179 = (inp[1]) ? node1185 : node1180;
									assign node1180 = (inp[7]) ? node1182 : 3'b000;
										assign node1182 = (inp[8]) ? 3'b100 : 3'b000;
									assign node1185 = (inp[11]) ? node1189 : node1186;
										assign node1186 = (inp[7]) ? 3'b010 : 3'b100;
										assign node1189 = (inp[7]) ? 3'b100 : 3'b000;
							assign node1192 = (inp[10]) ? node1206 : node1193;
								assign node1193 = (inp[2]) ? node1199 : node1194;
									assign node1194 = (inp[7]) ? node1196 : 3'b000;
										assign node1196 = (inp[1]) ? 3'b100 : 3'b000;
									assign node1199 = (inp[11]) ? node1203 : node1200;
										assign node1200 = (inp[7]) ? 3'b100 : 3'b100;
										assign node1203 = (inp[8]) ? 3'b000 : 3'b000;
								assign node1206 = (inp[11]) ? 3'b000 : node1207;
									assign node1207 = (inp[1]) ? node1209 : 3'b000;
										assign node1209 = (inp[7]) ? 3'b100 : 3'b000;
					assign node1213 = (inp[0]) ? node1267 : node1214;
						assign node1214 = (inp[10]) ? node1246 : node1215;
							assign node1215 = (inp[7]) ? node1231 : node1216;
								assign node1216 = (inp[5]) ? node1224 : node1217;
									assign node1217 = (inp[1]) ? node1221 : node1218;
										assign node1218 = (inp[11]) ? 3'b100 : 3'b100;
										assign node1221 = (inp[8]) ? 3'b110 : 3'b010;
									assign node1224 = (inp[1]) ? node1228 : node1225;
										assign node1225 = (inp[11]) ? 3'b000 : 3'b000;
										assign node1228 = (inp[8]) ? 3'b100 : 3'b000;
								assign node1231 = (inp[8]) ? node1239 : node1232;
									assign node1232 = (inp[11]) ? node1236 : node1233;
										assign node1233 = (inp[2]) ? 3'b000 : 3'b010;
										assign node1236 = (inp[5]) ? 3'b100 : 3'b000;
									assign node1239 = (inp[1]) ? node1243 : node1240;
										assign node1240 = (inp[5]) ? 3'b000 : 3'b010;
										assign node1243 = (inp[5]) ? 3'b010 : 3'b100;
							assign node1246 = (inp[5]) ? node1260 : node1247;
								assign node1247 = (inp[7]) ? node1253 : node1248;
									assign node1248 = (inp[1]) ? node1250 : 3'b000;
										assign node1250 = (inp[11]) ? 3'b000 : 3'b100;
									assign node1253 = (inp[1]) ? node1257 : node1254;
										assign node1254 = (inp[11]) ? 3'b000 : 3'b100;
										assign node1257 = (inp[11]) ? 3'b100 : 3'b010;
								assign node1260 = (inp[7]) ? node1262 : 3'b000;
									assign node1262 = (inp[1]) ? node1264 : 3'b000;
										assign node1264 = (inp[2]) ? 3'b100 : 3'b000;
						assign node1267 = (inp[10]) ? node1299 : node1268;
							assign node1268 = (inp[5]) ? node1284 : node1269;
								assign node1269 = (inp[11]) ? node1277 : node1270;
									assign node1270 = (inp[1]) ? node1274 : node1271;
										assign node1271 = (inp[7]) ? 3'b001 : 3'b110;
										assign node1274 = (inp[7]) ? 3'b001 : 3'b001;
									assign node1277 = (inp[7]) ? node1281 : node1278;
										assign node1278 = (inp[1]) ? 3'b110 : 3'b010;
										assign node1281 = (inp[2]) ? 3'b001 : 3'b110;
								assign node1284 = (inp[7]) ? node1292 : node1285;
									assign node1285 = (inp[2]) ? node1289 : node1286;
										assign node1286 = (inp[1]) ? 3'b010 : 3'b110;
										assign node1289 = (inp[1]) ? 3'b010 : 3'b010;
									assign node1292 = (inp[1]) ? node1296 : node1293;
										assign node1293 = (inp[8]) ? 3'b110 : 3'b010;
										assign node1296 = (inp[8]) ? 3'b110 : 3'b110;
							assign node1299 = (inp[5]) ? node1315 : node1300;
								assign node1300 = (inp[7]) ? node1308 : node1301;
									assign node1301 = (inp[1]) ? node1305 : node1302;
										assign node1302 = (inp[11]) ? 3'b100 : 3'b010;
										assign node1305 = (inp[11]) ? 3'b010 : 3'b010;
									assign node1308 = (inp[11]) ? node1312 : node1309;
										assign node1309 = (inp[8]) ? 3'b110 : 3'b110;
										assign node1312 = (inp[1]) ? 3'b110 : 3'b010;
								assign node1315 = (inp[7]) ? node1323 : node1316;
									assign node1316 = (inp[1]) ? node1320 : node1317;
										assign node1317 = (inp[8]) ? 3'b100 : 3'b000;
										assign node1320 = (inp[8]) ? 3'b100 : 3'b100;
									assign node1323 = (inp[11]) ? node1327 : node1324;
										assign node1324 = (inp[1]) ? 3'b010 : 3'b010;
										assign node1327 = (inp[1]) ? 3'b010 : 3'b100;
			assign node1330 = (inp[9]) ? node1506 : node1331;
				assign node1331 = (inp[6]) ? node1395 : node1332;
					assign node1332 = (inp[0]) ? node1350 : node1333;
						assign node1333 = (inp[1]) ? node1335 : 3'b000;
							assign node1335 = (inp[7]) ? node1337 : 3'b000;
								assign node1337 = (inp[5]) ? node1345 : node1338;
									assign node1338 = (inp[8]) ? node1342 : node1339;
										assign node1339 = (inp[10]) ? 3'b000 : 3'b000;
										assign node1342 = (inp[11]) ? 3'b000 : 3'b100;
									assign node1345 = (inp[10]) ? 3'b000 : node1346;
										assign node1346 = (inp[2]) ? 3'b000 : 3'b000;
						assign node1350 = (inp[7]) ? node1366 : node1351;
							assign node1351 = (inp[1]) ? node1353 : 3'b000;
								assign node1353 = (inp[5]) ? node1361 : node1354;
									assign node1354 = (inp[10]) ? node1358 : node1355;
										assign node1355 = (inp[11]) ? 3'b100 : 3'b001;
										assign node1358 = (inp[8]) ? 3'b100 : 3'b000;
									assign node1361 = (inp[10]) ? 3'b000 : node1362;
										assign node1362 = (inp[11]) ? 3'b000 : 3'b100;
							assign node1366 = (inp[1]) ? node1380 : node1367;
								assign node1367 = (inp[5]) ? node1375 : node1368;
									assign node1368 = (inp[10]) ? node1372 : node1369;
										assign node1369 = (inp[11]) ? 3'b100 : 3'b001;
										assign node1372 = (inp[11]) ? 3'b000 : 3'b100;
									assign node1375 = (inp[10]) ? 3'b000 : node1376;
										assign node1376 = (inp[11]) ? 3'b000 : 3'b100;
								assign node1380 = (inp[8]) ? node1388 : node1381;
									assign node1381 = (inp[5]) ? node1385 : node1382;
										assign node1382 = (inp[10]) ? 3'b100 : 3'b110;
										assign node1385 = (inp[10]) ? 3'b000 : 3'b100;
									assign node1388 = (inp[2]) ? node1392 : node1389;
										assign node1389 = (inp[10]) ? 3'b000 : 3'b000;
										assign node1392 = (inp[5]) ? 3'b010 : 3'b010;
					assign node1395 = (inp[0]) ? node1443 : node1396;
						assign node1396 = (inp[10]) ? node1424 : node1397;
							assign node1397 = (inp[7]) ? node1411 : node1398;
								assign node1398 = (inp[8]) ? node1404 : node1399;
									assign node1399 = (inp[2]) ? node1401 : 3'b000;
										assign node1401 = (inp[11]) ? 3'b000 : 3'b000;
									assign node1404 = (inp[5]) ? node1408 : node1405;
										assign node1405 = (inp[1]) ? 3'b000 : 3'b000;
										assign node1408 = (inp[1]) ? 3'b100 : 3'b000;
								assign node1411 = (inp[5]) ? node1419 : node1412;
									assign node1412 = (inp[1]) ? node1416 : node1413;
										assign node1413 = (inp[11]) ? 3'b110 : 3'b000;
										assign node1416 = (inp[8]) ? 3'b110 : 3'b010;
									assign node1419 = (inp[11]) ? 3'b100 : node1420;
										assign node1420 = (inp[1]) ? 3'b010 : 3'b000;
							assign node1424 = (inp[7]) ? node1432 : node1425;
								assign node1425 = (inp[1]) ? 3'b000 : node1426;
									assign node1426 = (inp[5]) ? 3'b000 : node1427;
										assign node1427 = (inp[8]) ? 3'b100 : 3'b000;
								assign node1432 = (inp[5]) ? node1438 : node1433;
									assign node1433 = (inp[11]) ? 3'b000 : node1434;
										assign node1434 = (inp[1]) ? 3'b010 : 3'b000;
									assign node1438 = (inp[1]) ? node1440 : 3'b000;
										assign node1440 = (inp[8]) ? 3'b100 : 3'b000;
						assign node1443 = (inp[5]) ? node1475 : node1444;
							assign node1444 = (inp[10]) ? node1460 : node1445;
								assign node1445 = (inp[11]) ? node1453 : node1446;
									assign node1446 = (inp[1]) ? node1450 : node1447;
										assign node1447 = (inp[8]) ? 3'b000 : 3'b000;
										assign node1450 = (inp[8]) ? 3'b101 : 3'b001;
									assign node1453 = (inp[1]) ? node1457 : node1454;
										assign node1454 = (inp[2]) ? 3'b000 : 3'b110;
										assign node1457 = (inp[7]) ? 3'b001 : 3'b010;
								assign node1460 = (inp[11]) ? node1468 : node1461;
									assign node1461 = (inp[8]) ? node1465 : node1462;
										assign node1462 = (inp[2]) ? 3'b110 : 3'b110;
										assign node1465 = (inp[2]) ? 3'b010 : 3'b110;
									assign node1468 = (inp[1]) ? node1472 : node1469;
										assign node1469 = (inp[8]) ? 3'b010 : 3'b100;
										assign node1472 = (inp[7]) ? 3'b110 : 3'b010;
							assign node1475 = (inp[10]) ? node1491 : node1476;
								assign node1476 = (inp[1]) ? node1484 : node1477;
									assign node1477 = (inp[7]) ? node1481 : node1478;
										assign node1478 = (inp[8]) ? 3'b010 : 3'b100;
										assign node1481 = (inp[11]) ? 3'b010 : 3'b110;
									assign node1484 = (inp[11]) ? node1488 : node1485;
										assign node1485 = (inp[8]) ? 3'b110 : 3'b110;
										assign node1488 = (inp[7]) ? 3'b110 : 3'b010;
								assign node1491 = (inp[7]) ? node1499 : node1492;
									assign node1492 = (inp[1]) ? node1496 : node1493;
										assign node1493 = (inp[2]) ? 3'b100 : 3'b000;
										assign node1496 = (inp[11]) ? 3'b100 : 3'b000;
									assign node1499 = (inp[1]) ? node1503 : node1500;
										assign node1500 = (inp[11]) ? 3'b100 : 3'b010;
										assign node1503 = (inp[11]) ? 3'b010 : 3'b010;
				assign node1506 = (inp[6]) ? node1526 : node1507;
					assign node1507 = (inp[7]) ? node1509 : 3'b000;
						assign node1509 = (inp[11]) ? 3'b000 : node1510;
							assign node1510 = (inp[1]) ? node1518 : node1511;
								assign node1511 = (inp[0]) ? node1513 : 3'b000;
									assign node1513 = (inp[5]) ? 3'b000 : node1514;
										assign node1514 = (inp[10]) ? 3'b000 : 3'b010;
								assign node1518 = (inp[5]) ? 3'b000 : node1519;
									assign node1519 = (inp[10]) ? 3'b000 : node1520;
										assign node1520 = (inp[0]) ? 3'b100 : 3'b000;
					assign node1526 = (inp[7]) ? node1544 : node1527;
						assign node1527 = (inp[1]) ? node1529 : 3'b000;
							assign node1529 = (inp[0]) ? node1531 : 3'b000;
								assign node1531 = (inp[5]) ? node1539 : node1532;
									assign node1532 = (inp[10]) ? node1536 : node1533;
										assign node1533 = (inp[2]) ? 3'b100 : 3'b000;
										assign node1536 = (inp[8]) ? 3'b000 : 3'b000;
									assign node1539 = (inp[8]) ? node1541 : 3'b000;
										assign node1541 = (inp[11]) ? 3'b000 : 3'b000;
						assign node1544 = (inp[10]) ? node1566 : node1545;
							assign node1545 = (inp[5]) ? node1557 : node1546;
								assign node1546 = (inp[0]) ? node1550 : node1547;
									assign node1547 = (inp[1]) ? 3'b100 : 3'b000;
									assign node1550 = (inp[11]) ? node1554 : node1551;
										assign node1551 = (inp[1]) ? 3'b010 : 3'b010;
										assign node1554 = (inp[1]) ? 3'b010 : 3'b100;
								assign node1557 = (inp[0]) ? node1559 : 3'b000;
									assign node1559 = (inp[11]) ? node1563 : node1560;
										assign node1560 = (inp[1]) ? 3'b100 : 3'b000;
										assign node1563 = (inp[1]) ? 3'b000 : 3'b000;
							assign node1566 = (inp[0]) ? node1568 : 3'b000;
								assign node1568 = (inp[1]) ? node1574 : node1569;
									assign node1569 = (inp[5]) ? 3'b000 : node1570;
										assign node1570 = (inp[11]) ? 3'b000 : 3'b000;
									assign node1574 = (inp[5]) ? node1578 : node1575;
										assign node1575 = (inp[8]) ? 3'b100 : 3'b000;
										assign node1578 = (inp[2]) ? 3'b000 : 3'b000;

endmodule