module dtc_split66_bm13 (
	input  wire [11-1:0] inp,
	output wire [1-1:0] outp
);

	wire [1-1:0] node1;
	wire [1-1:0] node2;
	wire [1-1:0] node3;
	wire [1-1:0] node4;
	wire [1-1:0] node6;
	wire [1-1:0] node8;
	wire [1-1:0] node10;
	wire [1-1:0] node12;
	wire [1-1:0] node15;
	wire [1-1:0] node16;
	wire [1-1:0] node18;
	wire [1-1:0] node20;
	wire [1-1:0] node22;
	wire [1-1:0] node25;
	wire [1-1:0] node26;
	wire [1-1:0] node28;
	wire [1-1:0] node30;
	wire [1-1:0] node33;
	wire [1-1:0] node34;
	wire [1-1:0] node36;
	wire [1-1:0] node39;
	wire [1-1:0] node40;
	wire [1-1:0] node44;
	wire [1-1:0] node45;
	wire [1-1:0] node46;
	wire [1-1:0] node48;
	wire [1-1:0] node50;
	wire [1-1:0] node52;
	wire [1-1:0] node55;
	wire [1-1:0] node56;
	wire [1-1:0] node58;
	wire [1-1:0] node60;
	wire [1-1:0] node63;
	wire [1-1:0] node64;
	wire [1-1:0] node66;
	wire [1-1:0] node69;
	wire [1-1:0] node70;
	wire [1-1:0] node74;
	wire [1-1:0] node75;
	wire [1-1:0] node76;
	wire [1-1:0] node78;
	wire [1-1:0] node79;
	wire [1-1:0] node82;
	wire [1-1:0] node85;
	wire [1-1:0] node86;
	wire [1-1:0] node89;
	wire [1-1:0] node90;
	wire [1-1:0] node94;
	wire [1-1:0] node95;
	wire [1-1:0] node96;
	wire [1-1:0] node98;
	wire [1-1:0] node101;
	wire [1-1:0] node102;
	wire [1-1:0] node106;
	wire [1-1:0] node107;
	wire [1-1:0] node108;
	wire [1-1:0] node113;
	wire [1-1:0] node114;
	wire [1-1:0] node115;
	wire [1-1:0] node116;
	wire [1-1:0] node118;
	wire [1-1:0] node120;
	wire [1-1:0] node122;
	wire [1-1:0] node125;
	wire [1-1:0] node126;
	wire [1-1:0] node128;
	wire [1-1:0] node130;
	wire [1-1:0] node133;
	wire [1-1:0] node134;
	wire [1-1:0] node136;
	wire [1-1:0] node139;
	wire [1-1:0] node140;
	wire [1-1:0] node144;
	wire [1-1:0] node145;
	wire [1-1:0] node146;
	wire [1-1:0] node148;
	wire [1-1:0] node150;
	wire [1-1:0] node153;
	wire [1-1:0] node154;
	wire [1-1:0] node156;
	wire [1-1:0] node159;
	wire [1-1:0] node160;
	wire [1-1:0] node164;
	wire [1-1:0] node165;
	wire [1-1:0] node166;
	wire [1-1:0] node168;
	wire [1-1:0] node171;
	wire [1-1:0] node172;
	wire [1-1:0] node176;
	wire [1-1:0] node177;
	wire [1-1:0] node178;
	wire [1-1:0] node183;
	wire [1-1:0] node184;
	wire [1-1:0] node185;
	wire [1-1:0] node186;
	wire [1-1:0] node188;
	wire [1-1:0] node190;
	wire [1-1:0] node193;
	wire [1-1:0] node194;
	wire [1-1:0] node196;
	wire [1-1:0] node199;
	wire [1-1:0] node200;
	wire [1-1:0] node204;
	wire [1-1:0] node205;
	wire [1-1:0] node206;
	wire [1-1:0] node208;
	wire [1-1:0] node211;
	wire [1-1:0] node212;
	wire [1-1:0] node216;
	wire [1-1:0] node217;
	wire [1-1:0] node218;
	wire [1-1:0] node223;
	wire [1-1:0] node224;
	wire [1-1:0] node225;
	wire [1-1:0] node226;
	wire [1-1:0] node228;
	wire [1-1:0] node231;
	wire [1-1:0] node232;
	wire [1-1:0] node236;
	wire [1-1:0] node237;
	wire [1-1:0] node238;
	wire [1-1:0] node243;
	wire [1-1:0] node244;
	wire [1-1:0] node245;
	wire [1-1:0] node246;
	wire [1-1:0] node252;
	wire [1-1:0] node253;
	wire [1-1:0] node254;
	wire [1-1:0] node255;
	wire [1-1:0] node256;
	wire [1-1:0] node258;
	wire [1-1:0] node260;
	wire [1-1:0] node262;
	wire [1-1:0] node265;
	wire [1-1:0] node266;
	wire [1-1:0] node268;
	wire [1-1:0] node270;
	wire [1-1:0] node273;
	wire [1-1:0] node274;
	wire [1-1:0] node276;
	wire [1-1:0] node279;
	wire [1-1:0] node280;
	wire [1-1:0] node284;
	wire [1-1:0] node285;
	wire [1-1:0] node286;
	wire [1-1:0] node288;
	wire [1-1:0] node290;
	wire [1-1:0] node293;
	wire [1-1:0] node294;
	wire [1-1:0] node296;
	wire [1-1:0] node299;
	wire [1-1:0] node300;
	wire [1-1:0] node303;
	wire [1-1:0] node306;
	wire [1-1:0] node307;
	wire [1-1:0] node308;
	wire [1-1:0] node310;
	wire [1-1:0] node313;
	wire [1-1:0] node314;
	wire [1-1:0] node318;
	wire [1-1:0] node319;
	wire [1-1:0] node320;
	wire [1-1:0] node325;
	wire [1-1:0] node326;
	wire [1-1:0] node327;
	wire [1-1:0] node328;
	wire [1-1:0] node330;
	wire [1-1:0] node332;
	wire [1-1:0] node335;
	wire [1-1:0] node336;
	wire [1-1:0] node338;
	wire [1-1:0] node341;
	wire [1-1:0] node342;
	wire [1-1:0] node345;
	wire [1-1:0] node348;
	wire [1-1:0] node349;
	wire [1-1:0] node350;
	wire [1-1:0] node352;
	wire [1-1:0] node355;
	wire [1-1:0] node356;
	wire [1-1:0] node360;
	wire [1-1:0] node361;
	wire [1-1:0] node362;
	wire [1-1:0] node367;
	wire [1-1:0] node368;
	wire [1-1:0] node369;
	wire [1-1:0] node370;
	wire [1-1:0] node372;
	wire [1-1:0] node375;
	wire [1-1:0] node376;
	wire [1-1:0] node380;
	wire [1-1:0] node381;
	wire [1-1:0] node382;
	wire [1-1:0] node387;
	wire [1-1:0] node388;
	wire [1-1:0] node389;
	wire [1-1:0] node390;
	wire [1-1:0] node396;
	wire [1-1:0] node397;
	wire [1-1:0] node398;
	wire [1-1:0] node399;
	wire [1-1:0] node400;
	wire [1-1:0] node402;
	wire [1-1:0] node404;
	wire [1-1:0] node407;
	wire [1-1:0] node408;
	wire [1-1:0] node410;
	wire [1-1:0] node413;
	wire [1-1:0] node414;
	wire [1-1:0] node418;
	wire [1-1:0] node419;
	wire [1-1:0] node420;
	wire [1-1:0] node422;
	wire [1-1:0] node425;
	wire [1-1:0] node426;
	wire [1-1:0] node430;
	wire [1-1:0] node431;
	wire [1-1:0] node432;
	wire [1-1:0] node437;
	wire [1-1:0] node438;
	wire [1-1:0] node439;
	wire [1-1:0] node440;
	wire [1-1:0] node442;
	wire [1-1:0] node445;
	wire [1-1:0] node446;
	wire [1-1:0] node450;
	wire [1-1:0] node451;
	wire [1-1:0] node452;
	wire [1-1:0] node457;
	wire [1-1:0] node458;
	wire [1-1:0] node459;
	wire [1-1:0] node460;
	wire [1-1:0] node466;
	wire [1-1:0] node467;
	wire [1-1:0] node468;
	wire [1-1:0] node469;
	wire [1-1:0] node470;
	wire [1-1:0] node472;
	wire [1-1:0] node475;
	wire [1-1:0] node476;
	wire [1-1:0] node480;
	wire [1-1:0] node481;
	wire [1-1:0] node482;
	wire [1-1:0] node487;
	wire [1-1:0] node488;
	wire [1-1:0] node489;
	wire [1-1:0] node490;
	wire [1-1:0] node496;
	wire [1-1:0] node497;
	wire [1-1:0] node498;
	wire [1-1:0] node499;
	wire [1-1:0] node500;

	assign outp = (inp[9]) ? node252 : node1;
		assign node1 = (inp[7]) ? node113 : node2;
			assign node2 = (inp[8]) ? node44 : node3;
				assign node3 = (inp[5]) ? node15 : node4;
					assign node4 = (inp[3]) ? node6 : 1'b1;
						assign node6 = (inp[6]) ? node8 : 1'b1;
							assign node8 = (inp[0]) ? node10 : 1'b1;
								assign node10 = (inp[2]) ? node12 : 1'b1;
									assign node12 = (inp[10]) ? 1'b0 : 1'b1;
					assign node15 = (inp[4]) ? node25 : node16;
						assign node16 = (inp[2]) ? node18 : 1'b1;
							assign node18 = (inp[6]) ? node20 : 1'b1;
								assign node20 = (inp[10]) ? node22 : 1'b1;
									assign node22 = (inp[3]) ? 1'b0 : 1'b1;
						assign node25 = (inp[10]) ? node33 : node26;
							assign node26 = (inp[6]) ? node28 : 1'b1;
								assign node28 = (inp[1]) ? node30 : 1'b1;
									assign node30 = (inp[2]) ? 1'b0 : 1'b1;
							assign node33 = (inp[1]) ? node39 : node34;
								assign node34 = (inp[2]) ? node36 : 1'b1;
									assign node36 = (inp[6]) ? 1'b0 : 1'b1;
								assign node39 = (inp[0]) ? 1'b0 : node40;
									assign node40 = (inp[2]) ? 1'b0 : 1'b1;
				assign node44 = (inp[0]) ? node74 : node45;
					assign node45 = (inp[4]) ? node55 : node46;
						assign node46 = (inp[2]) ? node48 : 1'b1;
							assign node48 = (inp[3]) ? node50 : 1'b1;
								assign node50 = (inp[1]) ? node52 : 1'b1;
									assign node52 = (inp[6]) ? 1'b0 : 1'b1;
						assign node55 = (inp[5]) ? node63 : node56;
							assign node56 = (inp[1]) ? node58 : 1'b1;
								assign node58 = (inp[3]) ? node60 : 1'b1;
									assign node60 = (inp[10]) ? 1'b0 : 1'b1;
							assign node63 = (inp[2]) ? node69 : node64;
								assign node64 = (inp[3]) ? node66 : 1'b1;
									assign node66 = (inp[1]) ? 1'b0 : 1'b1;
								assign node69 = (inp[6]) ? 1'b0 : node70;
									assign node70 = (inp[10]) ? 1'b0 : 1'b1;
					assign node74 = (inp[4]) ? node94 : node75;
						assign node75 = (inp[1]) ? node85 : node76;
							assign node76 = (inp[5]) ? node78 : 1'b1;
								assign node78 = (inp[3]) ? node82 : node79;
									assign node79 = (inp[2]) ? 1'b1 : 1'b1;
									assign node82 = (inp[10]) ? 1'b0 : 1'b0;
							assign node85 = (inp[6]) ? node89 : node86;
								assign node86 = (inp[2]) ? 1'b0 : 1'b1;
								assign node89 = (inp[10]) ? 1'b0 : node90;
									assign node90 = (inp[3]) ? 1'b0 : 1'b1;
						assign node94 = (inp[6]) ? node106 : node95;
							assign node95 = (inp[3]) ? node101 : node96;
								assign node96 = (inp[2]) ? node98 : 1'b1;
									assign node98 = (inp[10]) ? 1'b0 : 1'b1;
								assign node101 = (inp[5]) ? 1'b0 : node102;
									assign node102 = (inp[1]) ? 1'b0 : 1'b1;
							assign node106 = (inp[2]) ? 1'b0 : node107;
								assign node107 = (inp[5]) ? 1'b0 : node108;
									assign node108 = (inp[10]) ? 1'b0 : 1'b1;
			assign node113 = (inp[6]) ? node183 : node114;
				assign node114 = (inp[4]) ? node144 : node115;
					assign node115 = (inp[5]) ? node125 : node116;
						assign node116 = (inp[8]) ? node118 : 1'b1;
							assign node118 = (inp[0]) ? node120 : 1'b1;
								assign node120 = (inp[3]) ? node122 : 1'b1;
									assign node122 = (inp[2]) ? 1'b0 : 1'b1;
						assign node125 = (inp[10]) ? node133 : node126;
							assign node126 = (inp[2]) ? node128 : 1'b1;
								assign node128 = (inp[0]) ? node130 : 1'b1;
									assign node130 = (inp[8]) ? 1'b0 : 1'b1;
							assign node133 = (inp[8]) ? node139 : node134;
								assign node134 = (inp[0]) ? node136 : 1'b1;
									assign node136 = (inp[1]) ? 1'b0 : 1'b1;
								assign node139 = (inp[3]) ? 1'b0 : node140;
									assign node140 = (inp[2]) ? 1'b0 : 1'b1;
					assign node144 = (inp[2]) ? node164 : node145;
						assign node145 = (inp[1]) ? node153 : node146;
							assign node146 = (inp[0]) ? node148 : 1'b1;
								assign node148 = (inp[5]) ? node150 : 1'b1;
									assign node150 = (inp[10]) ? 1'b1 : 1'b0;
							assign node153 = (inp[5]) ? node159 : node154;
								assign node154 = (inp[8]) ? node156 : 1'b1;
									assign node156 = (inp[3]) ? 1'b0 : 1'b1;
								assign node159 = (inp[0]) ? 1'b0 : node160;
									assign node160 = (inp[10]) ? 1'b0 : 1'b1;
						assign node164 = (inp[0]) ? node176 : node165;
							assign node165 = (inp[3]) ? node171 : node166;
								assign node166 = (inp[10]) ? node168 : 1'b1;
									assign node168 = (inp[1]) ? 1'b0 : 1'b1;
								assign node171 = (inp[1]) ? 1'b0 : node172;
									assign node172 = (inp[5]) ? 1'b0 : 1'b1;
							assign node176 = (inp[10]) ? 1'b0 : node177;
								assign node177 = (inp[5]) ? 1'b0 : node178;
									assign node178 = (inp[8]) ? 1'b0 : 1'b1;
				assign node183 = (inp[10]) ? node223 : node184;
					assign node184 = (inp[0]) ? node204 : node185;
						assign node185 = (inp[4]) ? node193 : node186;
							assign node186 = (inp[2]) ? node188 : 1'b1;
								assign node188 = (inp[5]) ? node190 : 1'b1;
									assign node190 = (inp[8]) ? 1'b0 : 1'b1;
							assign node193 = (inp[1]) ? node199 : node194;
								assign node194 = (inp[5]) ? node196 : 1'b1;
									assign node196 = (inp[2]) ? 1'b0 : 1'b1;
								assign node199 = (inp[2]) ? 1'b0 : node200;
									assign node200 = (inp[3]) ? 1'b0 : 1'b1;
						assign node204 = (inp[2]) ? node216 : node205;
							assign node205 = (inp[8]) ? node211 : node206;
								assign node206 = (inp[1]) ? node208 : 1'b1;
									assign node208 = (inp[4]) ? 1'b0 : 1'b1;
								assign node211 = (inp[4]) ? 1'b0 : node212;
									assign node212 = (inp[3]) ? 1'b0 : 1'b1;
							assign node216 = (inp[1]) ? 1'b0 : node217;
								assign node217 = (inp[3]) ? 1'b0 : node218;
									assign node218 = (inp[8]) ? 1'b0 : 1'b1;
					assign node223 = (inp[4]) ? node243 : node224;
						assign node224 = (inp[2]) ? node236 : node225;
							assign node225 = (inp[0]) ? node231 : node226;
								assign node226 = (inp[5]) ? node228 : 1'b1;
									assign node228 = (inp[8]) ? 1'b0 : 1'b1;
								assign node231 = (inp[1]) ? 1'b0 : node232;
									assign node232 = (inp[3]) ? 1'b0 : 1'b1;
							assign node236 = (inp[8]) ? 1'b0 : node237;
								assign node237 = (inp[1]) ? 1'b0 : node238;
									assign node238 = (inp[0]) ? 1'b0 : 1'b1;
						assign node243 = (inp[8]) ? 1'b0 : node244;
							assign node244 = (inp[3]) ? 1'b0 : node245;
								assign node245 = (inp[0]) ? 1'b0 : node246;
									assign node246 = (inp[5]) ? 1'b0 : 1'b1;
		assign node252 = (inp[10]) ? node396 : node253;
			assign node253 = (inp[5]) ? node325 : node254;
				assign node254 = (inp[2]) ? node284 : node255;
					assign node255 = (inp[6]) ? node265 : node256;
						assign node256 = (inp[4]) ? node258 : 1'b1;
							assign node258 = (inp[7]) ? node260 : 1'b1;
								assign node260 = (inp[1]) ? node262 : 1'b1;
									assign node262 = (inp[8]) ? 1'b0 : 1'b1;
						assign node265 = (inp[8]) ? node273 : node266;
							assign node266 = (inp[0]) ? node268 : 1'b1;
								assign node268 = (inp[1]) ? node270 : 1'b1;
									assign node270 = (inp[7]) ? 1'b0 : 1'b1;
							assign node273 = (inp[4]) ? node279 : node274;
								assign node274 = (inp[0]) ? node276 : 1'b1;
									assign node276 = (inp[7]) ? 1'b0 : 1'b1;
								assign node279 = (inp[7]) ? 1'b0 : node280;
									assign node280 = (inp[0]) ? 1'b0 : 1'b1;
					assign node284 = (inp[3]) ? node306 : node285;
						assign node285 = (inp[0]) ? node293 : node286;
							assign node286 = (inp[8]) ? node288 : 1'b1;
								assign node288 = (inp[1]) ? node290 : 1'b1;
									assign node290 = (inp[4]) ? 1'b0 : 1'b1;
							assign node293 = (inp[4]) ? node299 : node294;
								assign node294 = (inp[8]) ? node296 : 1'b1;
									assign node296 = (inp[6]) ? 1'b0 : 1'b1;
								assign node299 = (inp[6]) ? node303 : node300;
									assign node300 = (inp[1]) ? 1'b0 : 1'b1;
									assign node303 = (inp[7]) ? 1'b0 : 1'b0;
						assign node306 = (inp[8]) ? node318 : node307;
							assign node307 = (inp[1]) ? node313 : node308;
								assign node308 = (inp[7]) ? node310 : 1'b1;
									assign node310 = (inp[6]) ? 1'b0 : 1'b1;
								assign node313 = (inp[4]) ? 1'b0 : node314;
									assign node314 = (inp[6]) ? 1'b0 : 1'b1;
							assign node318 = (inp[6]) ? 1'b0 : node319;
								assign node319 = (inp[4]) ? 1'b0 : node320;
									assign node320 = (inp[1]) ? 1'b0 : 1'b1;
				assign node325 = (inp[3]) ? node367 : node326;
					assign node326 = (inp[7]) ? node348 : node327;
						assign node327 = (inp[6]) ? node335 : node328;
							assign node328 = (inp[4]) ? node330 : 1'b1;
								assign node330 = (inp[0]) ? node332 : 1'b1;
									assign node332 = (inp[2]) ? 1'b0 : 1'b1;
							assign node335 = (inp[8]) ? node341 : node336;
								assign node336 = (inp[4]) ? node338 : 1'b1;
									assign node338 = (inp[2]) ? 1'b0 : 1'b1;
								assign node341 = (inp[1]) ? node345 : node342;
									assign node342 = (inp[0]) ? 1'b0 : 1'b1;
									assign node345 = (inp[2]) ? 1'b0 : 1'b0;
						assign node348 = (inp[1]) ? node360 : node349;
							assign node349 = (inp[6]) ? node355 : node350;
								assign node350 = (inp[8]) ? node352 : 1'b1;
									assign node352 = (inp[2]) ? 1'b0 : 1'b1;
								assign node355 = (inp[0]) ? 1'b0 : node356;
									assign node356 = (inp[4]) ? 1'b0 : 1'b1;
							assign node360 = (inp[8]) ? 1'b0 : node361;
								assign node361 = (inp[6]) ? 1'b0 : node362;
									assign node362 = (inp[2]) ? 1'b0 : 1'b1;
					assign node367 = (inp[0]) ? node387 : node368;
						assign node368 = (inp[4]) ? node380 : node369;
							assign node369 = (inp[2]) ? node375 : node370;
								assign node370 = (inp[1]) ? node372 : 1'b1;
									assign node372 = (inp[7]) ? 1'b0 : 1'b1;
								assign node375 = (inp[1]) ? 1'b0 : node376;
									assign node376 = (inp[8]) ? 1'b0 : 1'b1;
							assign node380 = (inp[6]) ? 1'b0 : node381;
								assign node381 = (inp[8]) ? 1'b0 : node382;
									assign node382 = (inp[7]) ? 1'b0 : 1'b1;
						assign node387 = (inp[7]) ? 1'b0 : node388;
							assign node388 = (inp[4]) ? 1'b0 : node389;
								assign node389 = (inp[1]) ? 1'b0 : node390;
									assign node390 = (inp[6]) ? 1'b0 : 1'b1;
			assign node396 = (inp[8]) ? node466 : node397;
				assign node397 = (inp[6]) ? node437 : node398;
					assign node398 = (inp[0]) ? node418 : node399;
						assign node399 = (inp[4]) ? node407 : node400;
							assign node400 = (inp[3]) ? node402 : 1'b1;
								assign node402 = (inp[1]) ? node404 : 1'b1;
									assign node404 = (inp[7]) ? 1'b0 : 1'b1;
							assign node407 = (inp[7]) ? node413 : node408;
								assign node408 = (inp[5]) ? node410 : 1'b1;
									assign node410 = (inp[2]) ? 1'b0 : 1'b1;
								assign node413 = (inp[1]) ? 1'b0 : node414;
									assign node414 = (inp[2]) ? 1'b0 : 1'b1;
						assign node418 = (inp[2]) ? node430 : node419;
							assign node419 = (inp[7]) ? node425 : node420;
								assign node420 = (inp[5]) ? node422 : 1'b1;
									assign node422 = (inp[3]) ? 1'b0 : 1'b1;
								assign node425 = (inp[1]) ? 1'b0 : node426;
									assign node426 = (inp[5]) ? 1'b0 : 1'b1;
							assign node430 = (inp[1]) ? 1'b0 : node431;
								assign node431 = (inp[3]) ? 1'b0 : node432;
									assign node432 = (inp[4]) ? 1'b0 : 1'b1;
					assign node437 = (inp[7]) ? node457 : node438;
						assign node438 = (inp[2]) ? node450 : node439;
							assign node439 = (inp[3]) ? node445 : node440;
								assign node440 = (inp[1]) ? node442 : 1'b1;
									assign node442 = (inp[4]) ? 1'b0 : 1'b1;
								assign node445 = (inp[4]) ? 1'b0 : node446;
									assign node446 = (inp[1]) ? 1'b0 : 1'b1;
							assign node450 = (inp[3]) ? 1'b0 : node451;
								assign node451 = (inp[1]) ? 1'b0 : node452;
									assign node452 = (inp[0]) ? 1'b0 : 1'b1;
						assign node457 = (inp[4]) ? 1'b0 : node458;
							assign node458 = (inp[5]) ? 1'b0 : node459;
								assign node459 = (inp[1]) ? 1'b0 : node460;
									assign node460 = (inp[3]) ? 1'b0 : 1'b1;
				assign node466 = (inp[1]) ? node496 : node467;
					assign node467 = (inp[0]) ? node487 : node468;
						assign node468 = (inp[6]) ? node480 : node469;
							assign node469 = (inp[5]) ? node475 : node470;
								assign node470 = (inp[2]) ? node472 : 1'b1;
									assign node472 = (inp[7]) ? 1'b0 : 1'b1;
								assign node475 = (inp[3]) ? 1'b0 : node476;
									assign node476 = (inp[7]) ? 1'b0 : 1'b1;
							assign node480 = (inp[3]) ? 1'b0 : node481;
								assign node481 = (inp[5]) ? 1'b0 : node482;
									assign node482 = (inp[2]) ? 1'b0 : 1'b1;
						assign node487 = (inp[5]) ? 1'b0 : node488;
							assign node488 = (inp[3]) ? 1'b0 : node489;
								assign node489 = (inp[7]) ? 1'b0 : node490;
									assign node490 = (inp[4]) ? 1'b0 : 1'b1;
					assign node496 = (inp[3]) ? 1'b0 : node497;
						assign node497 = (inp[6]) ? 1'b0 : node498;
							assign node498 = (inp[5]) ? 1'b0 : node499;
								assign node499 = (inp[4]) ? 1'b0 : node500;
									assign node500 = (inp[0]) ? 1'b0 : 1'b1;

endmodule