module dtc_split125_bm84 (
	input  wire [12-1:0] inp,
	output wire [3-1:0] outp
);

	wire [3-1:0] node1;
	wire [3-1:0] node2;
	wire [3-1:0] node3;
	wire [3-1:0] node4;
	wire [3-1:0] node6;
	wire [3-1:0] node8;
	wire [3-1:0] node11;
	wire [3-1:0] node12;
	wire [3-1:0] node13;
	wire [3-1:0] node15;
	wire [3-1:0] node18;
	wire [3-1:0] node19;
	wire [3-1:0] node22;
	wire [3-1:0] node25;
	wire [3-1:0] node26;
	wire [3-1:0] node27;
	wire [3-1:0] node31;
	wire [3-1:0] node34;
	wire [3-1:0] node35;
	wire [3-1:0] node36;
	wire [3-1:0] node37;
	wire [3-1:0] node40;
	wire [3-1:0] node42;
	wire [3-1:0] node45;
	wire [3-1:0] node46;
	wire [3-1:0] node47;
	wire [3-1:0] node51;
	wire [3-1:0] node52;
	wire [3-1:0] node56;
	wire [3-1:0] node57;
	wire [3-1:0] node59;
	wire [3-1:0] node62;
	wire [3-1:0] node64;
	wire [3-1:0] node65;
	wire [3-1:0] node69;
	wire [3-1:0] node70;
	wire [3-1:0] node71;
	wire [3-1:0] node72;
	wire [3-1:0] node73;
	wire [3-1:0] node75;
	wire [3-1:0] node78;
	wire [3-1:0] node79;
	wire [3-1:0] node82;
	wire [3-1:0] node85;
	wire [3-1:0] node86;
	wire [3-1:0] node88;
	wire [3-1:0] node92;
	wire [3-1:0] node93;
	wire [3-1:0] node96;
	wire [3-1:0] node99;
	wire [3-1:0] node100;
	wire [3-1:0] node101;
	wire [3-1:0] node104;
	wire [3-1:0] node107;
	wire [3-1:0] node108;
	wire [3-1:0] node110;
	wire [3-1:0] node112;
	wire [3-1:0] node116;
	wire [3-1:0] node117;
	wire [3-1:0] node118;
	wire [3-1:0] node119;
	wire [3-1:0] node120;
	wire [3-1:0] node121;
	wire [3-1:0] node122;
	wire [3-1:0] node126;
	wire [3-1:0] node128;
	wire [3-1:0] node131;
	wire [3-1:0] node133;
	wire [3-1:0] node136;
	wire [3-1:0] node137;
	wire [3-1:0] node139;
	wire [3-1:0] node142;
	wire [3-1:0] node144;
	wire [3-1:0] node147;
	wire [3-1:0] node148;
	wire [3-1:0] node149;
	wire [3-1:0] node150;
	wire [3-1:0] node153;
	wire [3-1:0] node156;
	wire [3-1:0] node160;
	wire [3-1:0] node161;
	wire [3-1:0] node162;
	wire [3-1:0] node163;

	assign outp = (inp[9]) ? node116 : node1;
		assign node1 = (inp[6]) ? node69 : node2;
			assign node2 = (inp[10]) ? node34 : node3;
				assign node3 = (inp[7]) ? node11 : node4;
					assign node4 = (inp[11]) ? node6 : 3'b111;
						assign node6 = (inp[8]) ? node8 : 3'b111;
							assign node8 = (inp[3]) ? 3'b011 : 3'b111;
					assign node11 = (inp[8]) ? node25 : node12;
						assign node12 = (inp[0]) ? node18 : node13;
							assign node13 = (inp[3]) ? node15 : 3'b011;
								assign node15 = (inp[11]) ? 3'b011 : 3'b111;
							assign node18 = (inp[11]) ? node22 : node19;
								assign node19 = (inp[2]) ? 3'b111 : 3'b111;
								assign node22 = (inp[5]) ? 3'b101 : 3'b111;
						assign node25 = (inp[11]) ? node31 : node26;
							assign node26 = (inp[3]) ? 3'b011 : node27;
								assign node27 = (inp[4]) ? 3'b111 : 3'b011;
							assign node31 = (inp[3]) ? 3'b101 : 3'b011;
				assign node34 = (inp[11]) ? node56 : node35;
					assign node35 = (inp[7]) ? node45 : node36;
						assign node36 = (inp[8]) ? node40 : node37;
							assign node37 = (inp[3]) ? 3'b011 : 3'b111;
							assign node40 = (inp[3]) ? node42 : 3'b011;
								assign node42 = (inp[4]) ? 3'b101 : 3'b001;
						assign node45 = (inp[4]) ? node51 : node46;
							assign node46 = (inp[8]) ? 3'b001 : node47;
								assign node47 = (inp[3]) ? 3'b111 : 3'b011;
							assign node51 = (inp[3]) ? 3'b001 : node52;
								assign node52 = (inp[8]) ? 3'b001 : 3'b101;
					assign node56 = (inp[7]) ? node62 : node57;
						assign node57 = (inp[4]) ? node59 : 3'b101;
							assign node59 = (inp[3]) ? 3'b001 : 3'b101;
						assign node62 = (inp[8]) ? node64 : 3'b101;
							assign node64 = (inp[3]) ? 3'b110 : node65;
								assign node65 = (inp[0]) ? 3'b101 : 3'b110;
			assign node69 = (inp[10]) ? node99 : node70;
				assign node70 = (inp[11]) ? node92 : node71;
					assign node71 = (inp[7]) ? node85 : node72;
						assign node72 = (inp[8]) ? node78 : node73;
							assign node73 = (inp[3]) ? node75 : 3'b011;
								assign node75 = (inp[4]) ? 3'b101 : 3'b011;
							assign node78 = (inp[5]) ? node82 : node79;
								assign node79 = (inp[4]) ? 3'b001 : 3'b011;
								assign node82 = (inp[0]) ? 3'b001 : 3'b001;
						assign node85 = (inp[8]) ? 3'b110 : node86;
							assign node86 = (inp[4]) ? node88 : 3'b001;
								assign node88 = (inp[3]) ? 3'b110 : 3'b001;
					assign node92 = (inp[8]) ? node96 : node93;
						assign node93 = (inp[7]) ? 3'b110 : 3'b001;
						assign node96 = (inp[7]) ? 3'b010 : 3'b110;
				assign node99 = (inp[7]) ? node107 : node100;
					assign node100 = (inp[11]) ? node104 : node101;
						assign node101 = (inp[8]) ? 3'b010 : 3'b110;
						assign node104 = (inp[8]) ? 3'b100 : 3'b010;
					assign node107 = (inp[11]) ? 3'b000 : node108;
						assign node108 = (inp[4]) ? node110 : 3'b100;
							assign node110 = (inp[0]) ? node112 : 3'b100;
								assign node112 = (inp[2]) ? 3'b100 : 3'b000;
		assign node116 = (inp[6]) ? node160 : node117;
			assign node117 = (inp[10]) ? node147 : node118;
				assign node118 = (inp[7]) ? node136 : node119;
					assign node119 = (inp[8]) ? node131 : node120;
						assign node120 = (inp[4]) ? node126 : node121;
							assign node121 = (inp[3]) ? 3'b001 : node122;
								assign node122 = (inp[11]) ? 3'b001 : 3'b101;
							assign node126 = (inp[3]) ? node128 : 3'b101;
								assign node128 = (inp[2]) ? 3'b110 : 3'b101;
						assign node131 = (inp[11]) ? node133 : 3'b000;
							assign node133 = (inp[3]) ? 3'b010 : 3'b110;
					assign node136 = (inp[11]) ? node142 : node137;
						assign node137 = (inp[8]) ? node139 : 3'b010;
							assign node139 = (inp[3]) ? 3'b100 : 3'b010;
						assign node142 = (inp[4]) ? node144 : 3'b100;
							assign node144 = (inp[8]) ? 3'b000 : 3'b100;
				assign node147 = (inp[7]) ? 3'b000 : node148;
					assign node148 = (inp[0]) ? node156 : node149;
						assign node149 = (inp[11]) ? node153 : node150;
							assign node150 = (inp[8]) ? 3'b100 : 3'b010;
							assign node153 = (inp[8]) ? 3'b000 : 3'b100;
						assign node156 = (inp[11]) ? 3'b000 : 3'b010;
			assign node160 = (inp[10]) ? 3'b000 : node161;
				assign node161 = (inp[7]) ? 3'b000 : node162;
					assign node162 = (inp[8]) ? 3'b000 : node163;
						assign node163 = (inp[11]) ? 3'b000 : 3'b100;

endmodule