module dtc_split75_bm64 (
	input  wire [16-1:0] inp,
	output wire [4-1:0] outp
);

	wire [4-1:0] node2;
	wire [4-1:0] node3;
	wire [4-1:0] node4;
	wire [4-1:0] node5;
	wire [4-1:0] node6;
	wire [4-1:0] node7;
	wire [4-1:0] node8;
	wire [4-1:0] node9;
	wire [4-1:0] node10;
	wire [4-1:0] node11;
	wire [4-1:0] node12;
	wire [4-1:0] node13;
	wire [4-1:0] node14;
	wire [4-1:0] node18;
	wire [4-1:0] node20;
	wire [4-1:0] node21;
	wire [4-1:0] node26;
	wire [4-1:0] node28;
	wire [4-1:0] node29;
	wire [4-1:0] node31;
	wire [4-1:0] node32;
	wire [4-1:0] node36;
	wire [4-1:0] node38;
	wire [4-1:0] node42;
	wire [4-1:0] node44;
	wire [4-1:0] node45;
	wire [4-1:0] node46;
	wire [4-1:0] node47;
	wire [4-1:0] node49;
	wire [4-1:0] node50;
	wire [4-1:0] node54;
	wire [4-1:0] node56;
	wire [4-1:0] node60;
	wire [4-1:0] node62;
	wire [4-1:0] node63;
	wire [4-1:0] node65;
	wire [4-1:0] node66;
	wire [4-1:0] node70;
	wire [4-1:0] node72;
	wire [4-1:0] node74;
	wire [4-1:0] node78;
	wire [4-1:0] node80;
	wire [4-1:0] node81;
	wire [4-1:0] node82;
	wire [4-1:0] node83;
	wire [4-1:0] node84;
	wire [4-1:0] node85;
	wire [4-1:0] node86;
	wire [4-1:0] node88;
	wire [4-1:0] node92;
	wire [4-1:0] node94;
	wire [4-1:0] node95;
	wire [4-1:0] node100;
	wire [4-1:0] node102;
	wire [4-1:0] node103;
	wire [4-1:0] node104;
	wire [4-1:0] node106;
	wire [4-1:0] node110;
	wire [4-1:0] node112;
	wire [4-1:0] node114;
	wire [4-1:0] node118;
	wire [4-1:0] node120;
	wire [4-1:0] node121;
	wire [4-1:0] node122;
	wire [4-1:0] node123;
	wire [4-1:0] node125;
	wire [4-1:0] node126;
	wire [4-1:0] node130;
	wire [4-1:0] node132;
	wire [4-1:0] node133;
	wire [4-1:0] node138;
	wire [4-1:0] node140;
	wire [4-1:0] node141;
	wire [4-1:0] node142;
	wire [4-1:0] node146;
	wire [4-1:0] node147;
	wire [4-1:0] node149;
	wire [4-1:0] node154;
	wire [4-1:0] node155;
	wire [4-1:0] node156;
	wire [4-1:0] node157;
	wire [4-1:0] node158;
	wire [4-1:0] node159;
	wire [4-1:0] node160;
	wire [4-1:0] node161;
	wire [4-1:0] node162;
	wire [4-1:0] node164;
	wire [4-1:0] node168;
	wire [4-1:0] node170;
	wire [4-1:0] node171;
	wire [4-1:0] node176;
	wire [4-1:0] node178;
	wire [4-1:0] node179;
	wire [4-1:0] node180;
	wire [4-1:0] node182;
	wire [4-1:0] node186;
	wire [4-1:0] node188;
	wire [4-1:0] node190;
	wire [4-1:0] node194;
	wire [4-1:0] node196;
	wire [4-1:0] node197;
	wire [4-1:0] node198;
	wire [4-1:0] node199;
	wire [4-1:0] node201;
	wire [4-1:0] node202;
	wire [4-1:0] node206;
	wire [4-1:0] node208;
	wire [4-1:0] node210;
	wire [4-1:0] node214;
	wire [4-1:0] node216;
	wire [4-1:0] node217;
	wire [4-1:0] node219;
	wire [4-1:0] node220;
	wire [4-1:0] node224;
	wire [4-1:0] node226;
	wire [4-1:0] node228;
	wire [4-1:0] node232;
	wire [4-1:0] node233;
	wire [4-1:0] node234;
	wire [4-1:0] node235;
	wire [4-1:0] node237;
	wire [4-1:0] node238;
	wire [4-1:0] node239;
	wire [4-1:0] node241;
	wire [4-1:0] node242;
	wire [4-1:0] node246;
	wire [4-1:0] node248;
	wire [4-1:0] node249;
	wire [4-1:0] node250;
	wire [4-1:0] node257;
	wire [4-1:0] node258;
	wire [4-1:0] node259;
	wire [4-1:0] node261;
	wire [4-1:0] node262;
	wire [4-1:0] node263;
	wire [4-1:0] node265;
	wire [4-1:0] node266;
	wire [4-1:0] node270;
	wire [4-1:0] node272;
	wire [4-1:0] node277;
	wire [4-1:0] node278;
	wire [4-1:0] node279;
	wire [4-1:0] node280;
	wire [4-1:0] node282;
	wire [4-1:0] node283;
	wire [4-1:0] node284;
	wire [4-1:0] node291;
	wire [4-1:0] node292;
	wire [4-1:0] node294;
	wire [4-1:0] node295;
	wire [4-1:0] node296;
	wire [4-1:0] node298;
	wire [4-1:0] node303;
	wire [4-1:0] node304;
	wire [4-1:0] node305;
	wire [4-1:0] node306;
	wire [4-1:0] node307;
	wire [4-1:0] node313;
	wire [4-1:0] node314;
	wire [4-1:0] node316;
	wire [4-1:0] node317;
	wire [4-1:0] node322;
	wire [4-1:0] node323;
	wire [4-1:0] node324;
	wire [4-1:0] node325;
	wire [4-1:0] node326;
	wire [4-1:0] node327;
	wire [4-1:0] node328;
	wire [4-1:0] node330;
	wire [4-1:0] node334;
	wire [4-1:0] node335;
	wire [4-1:0] node337;
	wire [4-1:0] node342;
	wire [4-1:0] node344;
	wire [4-1:0] node345;
	wire [4-1:0] node346;
	wire [4-1:0] node348;
	wire [4-1:0] node352;
	wire [4-1:0] node353;
	wire [4-1:0] node355;
	wire [4-1:0] node360;
	wire [4-1:0] node362;
	wire [4-1:0] node363;
	wire [4-1:0] node364;
	wire [4-1:0] node365;
	wire [4-1:0] node366;
	wire [4-1:0] node368;
	wire [4-1:0] node372;
	wire [4-1:0] node374;
	wire [4-1:0] node375;
	wire [4-1:0] node380;
	wire [4-1:0] node382;
	wire [4-1:0] node383;
	wire [4-1:0] node384;
	wire [4-1:0] node386;
	wire [4-1:0] node390;
	wire [4-1:0] node392;
	wire [4-1:0] node393;
	wire [4-1:0] node397;
	wire [4-1:0] node398;
	wire [4-1:0] node400;
	wire [4-1:0] node401;
	wire [4-1:0] node402;
	wire [4-1:0] node403;
	wire [4-1:0] node404;
	wire [4-1:0] node405;
	wire [4-1:0] node406;
	wire [4-1:0] node407;
	wire [4-1:0] node408;
	wire [4-1:0] node410;
	wire [4-1:0] node414;
	wire [4-1:0] node415;
	wire [4-1:0] node417;
	wire [4-1:0] node422;
	wire [4-1:0] node424;
	wire [4-1:0] node425;
	wire [4-1:0] node426;
	wire [4-1:0] node428;
	wire [4-1:0] node432;
	wire [4-1:0] node434;
	wire [4-1:0] node435;
	wire [4-1:0] node440;
	wire [4-1:0] node442;
	wire [4-1:0] node443;
	wire [4-1:0] node444;
	wire [4-1:0] node445;
	wire [4-1:0] node446;
	wire [4-1:0] node447;
	wire [4-1:0] node448;
	wire [4-1:0] node454;
	wire [4-1:0] node456;
	wire [4-1:0] node457;
	wire [4-1:0] node462;
	wire [4-1:0] node464;
	wire [4-1:0] node465;
	wire [4-1:0] node466;
	wire [4-1:0] node470;
	wire [4-1:0] node472;
	wire [4-1:0] node474;
	wire [4-1:0] node478;
	wire [4-1:0] node480;
	wire [4-1:0] node481;
	wire [4-1:0] node482;
	wire [4-1:0] node483;
	wire [4-1:0] node484;
	wire [4-1:0] node485;
	wire [4-1:0] node487;
	wire [4-1:0] node488;
	wire [4-1:0] node489;
	wire [4-1:0] node494;
	wire [4-1:0] node496;
	wire [4-1:0] node498;
	wire [4-1:0] node502;
	wire [4-1:0] node504;
	wire [4-1:0] node506;
	wire [4-1:0] node508;
	wire [4-1:0] node510;
	wire [4-1:0] node514;
	wire [4-1:0] node516;
	wire [4-1:0] node517;
	wire [4-1:0] node518;
	wire [4-1:0] node519;
	wire [4-1:0] node520;
	wire [4-1:0] node521;
	wire [4-1:0] node526;
	wire [4-1:0] node527;
	wire [4-1:0] node529;
	wire [4-1:0] node534;
	wire [4-1:0] node536;
	wire [4-1:0] node538;
	wire [4-1:0] node540;
	wire [4-1:0] node542;
	wire [4-1:0] node545;
	wire [4-1:0] node546;
	wire [4-1:0] node547;
	wire [4-1:0] node548;
	wire [4-1:0] node549;
	wire [4-1:0] node550;
	wire [4-1:0] node551;
	wire [4-1:0] node553;
	wire [4-1:0] node554;
	wire [4-1:0] node558;
	wire [4-1:0] node560;
	wire [4-1:0] node562;
	wire [4-1:0] node565;
	wire [4-1:0] node567;
	wire [4-1:0] node568;
	wire [4-1:0] node569;
	wire [4-1:0] node570;
	wire [4-1:0] node572;
	wire [4-1:0] node578;
	wire [4-1:0] node580;
	wire [4-1:0] node581;
	wire [4-1:0] node582;
	wire [4-1:0] node583;
	wire [4-1:0] node588;
	wire [4-1:0] node590;
	wire [4-1:0] node592;
	wire [4-1:0] node595;
	wire [4-1:0] node596;
	wire [4-1:0] node597;
	wire [4-1:0] node598;
	wire [4-1:0] node599;
	wire [4-1:0] node600;
	wire [4-1:0] node601;
	wire [4-1:0] node605;
	wire [4-1:0] node606;
	wire [4-1:0] node611;
	wire [4-1:0] node613;
	wire [4-1:0] node614;
	wire [4-1:0] node615;
	wire [4-1:0] node616;
	wire [4-1:0] node622;
	wire [4-1:0] node623;
	wire [4-1:0] node625;
	wire [4-1:0] node627;
	wire [4-1:0] node629;
	wire [4-1:0] node631;
	wire [4-1:0] node635;
	wire [4-1:0] node636;
	wire [4-1:0] node638;
	wire [4-1:0] node639;
	wire [4-1:0] node641;
	wire [4-1:0] node643;
	wire [4-1:0] node646;
	wire [4-1:0] node648;
	wire [4-1:0] node649;
	wire [4-1:0] node650;
	wire [4-1:0] node656;
	wire [4-1:0] node657;
	wire [4-1:0] node658;
	wire [4-1:0] node659;
	wire [4-1:0] node660;
	wire [4-1:0] node661;
	wire [4-1:0] node662;
	wire [4-1:0] node665;
	wire [4-1:0] node666;
	wire [4-1:0] node670;
	wire [4-1:0] node671;
	wire [4-1:0] node673;
	wire [4-1:0] node675;
	wire [4-1:0] node678;
	wire [4-1:0] node681;
	wire [4-1:0] node682;
	wire [4-1:0] node683;
	wire [4-1:0] node686;
	wire [4-1:0] node689;
	wire [4-1:0] node690;
	wire [4-1:0] node691;
	wire [4-1:0] node695;
	wire [4-1:0] node696;
	wire [4-1:0] node698;
	wire [4-1:0] node702;
	wire [4-1:0] node703;
	wire [4-1:0] node704;
	wire [4-1:0] node705;
	wire [4-1:0] node709;
	wire [4-1:0] node710;
	wire [4-1:0] node713;
	wire [4-1:0] node716;
	wire [4-1:0] node717;
	wire [4-1:0] node718;
	wire [4-1:0] node719;
	wire [4-1:0] node723;
	wire [4-1:0] node724;
	wire [4-1:0] node728;
	wire [4-1:0] node729;
	wire [4-1:0] node732;
	wire [4-1:0] node735;
	wire [4-1:0] node736;
	wire [4-1:0] node737;
	wire [4-1:0] node738;
	wire [4-1:0] node739;
	wire [4-1:0] node743;
	wire [4-1:0] node744;
	wire [4-1:0] node745;
	wire [4-1:0] node749;
	wire [4-1:0] node751;
	wire [4-1:0] node754;
	wire [4-1:0] node755;
	wire [4-1:0] node756;
	wire [4-1:0] node760;
	wire [4-1:0] node761;
	wire [4-1:0] node764;
	wire [4-1:0] node767;
	wire [4-1:0] node768;
	wire [4-1:0] node769;
	wire [4-1:0] node770;
	wire [4-1:0] node772;
	wire [4-1:0] node774;
	wire [4-1:0] node777;
	wire [4-1:0] node780;
	wire [4-1:0] node781;
	wire [4-1:0] node782;
	wire [4-1:0] node784;
	wire [4-1:0] node789;
	wire [4-1:0] node790;
	wire [4-1:0] node792;
	wire [4-1:0] node795;
	wire [4-1:0] node797;
	wire [4-1:0] node798;
	wire [4-1:0] node799;
	wire [4-1:0] node804;
	wire [4-1:0] node805;
	wire [4-1:0] node806;
	wire [4-1:0] node807;
	wire [4-1:0] node808;
	wire [4-1:0] node809;
	wire [4-1:0] node811;
	wire [4-1:0] node815;
	wire [4-1:0] node816;
	wire [4-1:0] node820;
	wire [4-1:0] node821;
	wire [4-1:0] node823;
	wire [4-1:0] node826;
	wire [4-1:0] node828;
	wire [4-1:0] node829;
	wire [4-1:0] node833;
	wire [4-1:0] node834;
	wire [4-1:0] node835;
	wire [4-1:0] node837;
	wire [4-1:0] node839;
	wire [4-1:0] node842;
	wire [4-1:0] node843;
	wire [4-1:0] node847;
	wire [4-1:0] node848;
	wire [4-1:0] node849;
	wire [4-1:0] node850;
	wire [4-1:0] node851;
	wire [4-1:0] node857;
	wire [4-1:0] node858;
	wire [4-1:0] node860;
	wire [4-1:0] node862;
	wire [4-1:0] node865;
	wire [4-1:0] node868;
	wire [4-1:0] node869;
	wire [4-1:0] node870;
	wire [4-1:0] node871;
	wire [4-1:0] node873;
	wire [4-1:0] node875;
	wire [4-1:0] node878;
	wire [4-1:0] node881;
	wire [4-1:0] node882;
	wire [4-1:0] node883;
	wire [4-1:0] node884;
	wire [4-1:0] node886;
	wire [4-1:0] node891;
	wire [4-1:0] node892;
	wire [4-1:0] node893;
	wire [4-1:0] node895;
	wire [4-1:0] node898;
	wire [4-1:0] node900;
	wire [4-1:0] node901;
	wire [4-1:0] node905;
	wire [4-1:0] node906;
	wire [4-1:0] node908;
	wire [4-1:0] node911;
	wire [4-1:0] node912;
	wire [4-1:0] node916;
	wire [4-1:0] node917;
	wire [4-1:0] node918;
	wire [4-1:0] node920;
	wire [4-1:0] node921;
	wire [4-1:0] node926;
	wire [4-1:0] node927;
	wire [4-1:0] node928;
	wire [4-1:0] node930;
	wire [4-1:0] node932;
	wire [4-1:0] node937;
	wire [4-1:0] node938;
	wire [4-1:0] node939;
	wire [4-1:0] node940;
	wire [4-1:0] node941;
	wire [4-1:0] node942;
	wire [4-1:0] node944;
	wire [4-1:0] node945;
	wire [4-1:0] node946;
	wire [4-1:0] node951;
	wire [4-1:0] node952;
	wire [4-1:0] node954;
	wire [4-1:0] node955;
	wire [4-1:0] node956;
	wire [4-1:0] node962;
	wire [4-1:0] node963;
	wire [4-1:0] node964;
	wire [4-1:0] node966;
	wire [4-1:0] node968;
	wire [4-1:0] node971;
	wire [4-1:0] node972;
	wire [4-1:0] node973;
	wire [4-1:0] node978;
	wire [4-1:0] node979;
	wire [4-1:0] node981;
	wire [4-1:0] node982;
	wire [4-1:0] node983;
	wire [4-1:0] node989;
	wire [4-1:0] node990;
	wire [4-1:0] node991;
	wire [4-1:0] node992;
	wire [4-1:0] node993;
	wire [4-1:0] node995;
	wire [4-1:0] node1000;
	wire [4-1:0] node1001;
	wire [4-1:0] node1003;
	wire [4-1:0] node1005;
	wire [4-1:0] node1006;
	wire [4-1:0] node1010;
	wire [4-1:0] node1012;
	wire [4-1:0] node1015;
	wire [4-1:0] node1016;
	wire [4-1:0] node1018;
	wire [4-1:0] node1019;
	wire [4-1:0] node1023;
	wire [4-1:0] node1024;
	wire [4-1:0] node1026;
	wire [4-1:0] node1027;
	wire [4-1:0] node1032;
	wire [4-1:0] node1033;
	wire [4-1:0] node1034;
	wire [4-1:0] node1035;
	wire [4-1:0] node1036;
	wire [4-1:0] node1037;
	wire [4-1:0] node1042;
	wire [4-1:0] node1044;
	wire [4-1:0] node1046;
	wire [4-1:0] node1049;
	wire [4-1:0] node1051;
	wire [4-1:0] node1052;
	wire [4-1:0] node1053;
	wire [4-1:0] node1055;
	wire [4-1:0] node1058;
	wire [4-1:0] node1059;
	wire [4-1:0] node1064;
	wire [4-1:0] node1065;
	wire [4-1:0] node1066;
	wire [4-1:0] node1067;
	wire [4-1:0] node1068;
	wire [4-1:0] node1069;
	wire [4-1:0] node1070;
	wire [4-1:0] node1075;
	wire [4-1:0] node1077;
	wire [4-1:0] node1081;
	wire [4-1:0] node1083;
	wire [4-1:0] node1084;
	wire [4-1:0] node1085;
	wire [4-1:0] node1086;
	wire [4-1:0] node1088;
	wire [4-1:0] node1094;
	wire [4-1:0] node1095;
	wire [4-1:0] node1096;
	wire [4-1:0] node1097;
	wire [4-1:0] node1102;
	wire [4-1:0] node1104;
	wire [4-1:0] node1105;
	wire [4-1:0] node1109;
	wire [4-1:0] node1110;
	wire [4-1:0] node1111;
	wire [4-1:0] node1112;
	wire [4-1:0] node1113;
	wire [4-1:0] node1114;
	wire [4-1:0] node1115;
	wire [4-1:0] node1116;
	wire [4-1:0] node1120;
	wire [4-1:0] node1121;
	wire [4-1:0] node1125;
	wire [4-1:0] node1126;
	wire [4-1:0] node1127;
	wire [4-1:0] node1131;
	wire [4-1:0] node1133;
	wire [4-1:0] node1136;
	wire [4-1:0] node1137;
	wire [4-1:0] node1138;
	wire [4-1:0] node1140;
	wire [4-1:0] node1142;
	wire [4-1:0] node1145;
	wire [4-1:0] node1147;
	wire [4-1:0] node1150;
	wire [4-1:0] node1151;
	wire [4-1:0] node1152;
	wire [4-1:0] node1156;
	wire [4-1:0] node1159;
	wire [4-1:0] node1160;
	wire [4-1:0] node1161;
	wire [4-1:0] node1162;
	wire [4-1:0] node1163;
	wire [4-1:0] node1165;
	wire [4-1:0] node1169;
	wire [4-1:0] node1170;
	wire [4-1:0] node1174;
	wire [4-1:0] node1177;
	wire [4-1:0] node1178;
	wire [4-1:0] node1179;
	wire [4-1:0] node1181;
	wire [4-1:0] node1182;
	wire [4-1:0] node1187;
	wire [4-1:0] node1188;
	wire [4-1:0] node1189;
	wire [4-1:0] node1191;
	wire [4-1:0] node1196;
	wire [4-1:0] node1197;
	wire [4-1:0] node1198;
	wire [4-1:0] node1199;
	wire [4-1:0] node1200;
	wire [4-1:0] node1203;
	wire [4-1:0] node1204;
	wire [4-1:0] node1205;
	wire [4-1:0] node1210;
	wire [4-1:0] node1211;
	wire [4-1:0] node1212;
	wire [4-1:0] node1215;
	wire [4-1:0] node1217;
	wire [4-1:0] node1220;
	wire [4-1:0] node1221;
	wire [4-1:0] node1224;
	wire [4-1:0] node1227;
	wire [4-1:0] node1228;
	wire [4-1:0] node1229;
	wire [4-1:0] node1230;
	wire [4-1:0] node1232;
	wire [4-1:0] node1236;
	wire [4-1:0] node1237;
	wire [4-1:0] node1241;
	wire [4-1:0] node1242;
	wire [4-1:0] node1243;
	wire [4-1:0] node1246;
	wire [4-1:0] node1249;
	wire [4-1:0] node1250;
	wire [4-1:0] node1251;
	wire [4-1:0] node1255;
	wire [4-1:0] node1257;
	wire [4-1:0] node1260;
	wire [4-1:0] node1261;
	wire [4-1:0] node1262;
	wire [4-1:0] node1263;
	wire [4-1:0] node1264;
	wire [4-1:0] node1266;
	wire [4-1:0] node1269;
	wire [4-1:0] node1271;
	wire [4-1:0] node1274;
	wire [4-1:0] node1275;
	wire [4-1:0] node1276;
	wire [4-1:0] node1280;
	wire [4-1:0] node1281;
	wire [4-1:0] node1285;
	wire [4-1:0] node1288;
	wire [4-1:0] node1289;
	wire [4-1:0] node1290;
	wire [4-1:0] node1291;
	wire [4-1:0] node1292;
	wire [4-1:0] node1296;
	wire [4-1:0] node1298;
	wire [4-1:0] node1301;
	wire [4-1:0] node1302;
	wire [4-1:0] node1304;
	wire [4-1:0] node1307;
	wire [4-1:0] node1309;
	wire [4-1:0] node1312;
	wire [4-1:0] node1315;
	wire [4-1:0] node1316;
	wire [4-1:0] node1317;
	wire [4-1:0] node1318;
	wire [4-1:0] node1319;
	wire [4-1:0] node1320;
	wire [4-1:0] node1321;
	wire [4-1:0] node1322;
	wire [4-1:0] node1325;
	wire [4-1:0] node1328;
	wire [4-1:0] node1329;
	wire [4-1:0] node1333;
	wire [4-1:0] node1334;
	wire [4-1:0] node1337;
	wire [4-1:0] node1338;
	wire [4-1:0] node1341;
	wire [4-1:0] node1344;
	wire [4-1:0] node1345;
	wire [4-1:0] node1346;
	wire [4-1:0] node1347;
	wire [4-1:0] node1351;
	wire [4-1:0] node1353;
	wire [4-1:0] node1356;
	wire [4-1:0] node1357;
	wire [4-1:0] node1358;
	wire [4-1:0] node1361;
	wire [4-1:0] node1364;
	wire [4-1:0] node1366;
	wire [4-1:0] node1369;
	wire [4-1:0] node1370;
	wire [4-1:0] node1371;
	wire [4-1:0] node1373;
	wire [4-1:0] node1376;
	wire [4-1:0] node1377;
	wire [4-1:0] node1378;
	wire [4-1:0] node1382;
	wire [4-1:0] node1385;
	wire [4-1:0] node1386;
	wire [4-1:0] node1387;
	wire [4-1:0] node1390;
	wire [4-1:0] node1391;
	wire [4-1:0] node1395;
	wire [4-1:0] node1396;
	wire [4-1:0] node1398;
	wire [4-1:0] node1401;
	wire [4-1:0] node1402;
	wire [4-1:0] node1405;
	wire [4-1:0] node1408;
	wire [4-1:0] node1409;
	wire [4-1:0] node1410;
	wire [4-1:0] node1413;
	wire [4-1:0] node1416;
	wire [4-1:0] node1417;
	wire [4-1:0] node1420;
	wire [4-1:0] node1423;
	wire [4-1:0] node1424;
	wire [4-1:0] node1425;
	wire [4-1:0] node1426;
	wire [4-1:0] node1429;
	wire [4-1:0] node1432;
	wire [4-1:0] node1433;
	wire [4-1:0] node1436;
	wire [4-1:0] node1440;
	wire [4-1:0] node1442;
	wire [4-1:0] node1443;
	wire [4-1:0] node1444;
	wire [4-1:0] node1445;
	wire [4-1:0] node1446;
	wire [4-1:0] node1447;
	wire [4-1:0] node1448;
	wire [4-1:0] node1449;
	wire [4-1:0] node1450;
	wire [4-1:0] node1451;
	wire [4-1:0] node1452;
	wire [4-1:0] node1454;
	wire [4-1:0] node1458;
	wire [4-1:0] node1459;
	wire [4-1:0] node1461;
	wire [4-1:0] node1466;
	wire [4-1:0] node1468;
	wire [4-1:0] node1469;
	wire [4-1:0] node1470;
	wire [4-1:0] node1474;
	wire [4-1:0] node1476;
	wire [4-1:0] node1480;
	wire [4-1:0] node1482;
	wire [4-1:0] node1483;
	wire [4-1:0] node1484;
	wire [4-1:0] node1485;
	wire [4-1:0] node1486;
	wire [4-1:0] node1488;
	wire [4-1:0] node1492;
	wire [4-1:0] node1494;
	wire [4-1:0] node1496;
	wire [4-1:0] node1500;
	wire [4-1:0] node1502;
	wire [4-1:0] node1503;
	wire [4-1:0] node1504;
	wire [4-1:0] node1505;
	wire [4-1:0] node1510;
	wire [4-1:0] node1511;
	wire [4-1:0] node1513;
	wire [4-1:0] node1518;
	wire [4-1:0] node1519;
	wire [4-1:0] node1520;
	wire [4-1:0] node1521;
	wire [4-1:0] node1522;
	wire [4-1:0] node1523;
	wire [4-1:0] node1524;
	wire [4-1:0] node1526;
	wire [4-1:0] node1530;
	wire [4-1:0] node1532;
	wire [4-1:0] node1533;
	wire [4-1:0] node1538;
	wire [4-1:0] node1540;
	wire [4-1:0] node1541;
	wire [4-1:0] node1542;
	wire [4-1:0] node1544;
	wire [4-1:0] node1548;
	wire [4-1:0] node1550;
	wire [4-1:0] node1551;
	wire [4-1:0] node1556;
	wire [4-1:0] node1557;
	wire [4-1:0] node1558;
	wire [4-1:0] node1559;
	wire [4-1:0] node1561;
	wire [4-1:0] node1562;
	wire [4-1:0] node1563;
	wire [4-1:0] node1564;
	wire [4-1:0] node1570;
	wire [4-1:0] node1572;
	wire [4-1:0] node1574;
	wire [4-1:0] node1576;
	wire [4-1:0] node1577;
	wire [4-1:0] node1581;
	wire [4-1:0] node1582;
	wire [4-1:0] node1583;
	wire [4-1:0] node1584;
	wire [4-1:0] node1586;
	wire [4-1:0] node1590;
	wire [4-1:0] node1592;
	wire [4-1:0] node1594;
	wire [4-1:0] node1598;
	wire [4-1:0] node1599;
	wire [4-1:0] node1601;
	wire [4-1:0] node1602;
	wire [4-1:0] node1603;
	wire [4-1:0] node1605;
	wire [4-1:0] node1606;
	wire [4-1:0] node1611;
	wire [4-1:0] node1613;
	wire [4-1:0] node1614;
	wire [4-1:0] node1615;
	wire [4-1:0] node1620;
	wire [4-1:0] node1622;
	wire [4-1:0] node1623;
	wire [4-1:0] node1625;
	wire [4-1:0] node1626;
	wire [4-1:0] node1630;
	wire [4-1:0] node1632;
	wire [4-1:0] node1634;
	wire [4-1:0] node1637;
	wire [4-1:0] node1638;
	wire [4-1:0] node1640;
	wire [4-1:0] node1641;
	wire [4-1:0] node1642;
	wire [4-1:0] node1643;
	wire [4-1:0] node1644;
	wire [4-1:0] node1645;
	wire [4-1:0] node1647;
	wire [4-1:0] node1650;
	wire [4-1:0] node1652;
	wire [4-1:0] node1656;
	wire [4-1:0] node1658;
	wire [4-1:0] node1659;
	wire [4-1:0] node1660;
	wire [4-1:0] node1662;
	wire [4-1:0] node1666;
	wire [4-1:0] node1668;
	wire [4-1:0] node1670;
	wire [4-1:0] node1674;
	wire [4-1:0] node1676;
	wire [4-1:0] node1677;
	wire [4-1:0] node1678;
	wire [4-1:0] node1679;
	wire [4-1:0] node1681;
	wire [4-1:0] node1684;
	wire [4-1:0] node1686;
	wire [4-1:0] node1687;
	wire [4-1:0] node1692;
	wire [4-1:0] node1694;
	wire [4-1:0] node1695;
	wire [4-1:0] node1696;
	wire [4-1:0] node1700;
	wire [4-1:0] node1701;
	wire [4-1:0] node1705;
	wire [4-1:0] node1706;
	wire [4-1:0] node1707;
	wire [4-1:0] node1708;
	wire [4-1:0] node1709;
	wire [4-1:0] node1710;
	wire [4-1:0] node1711;
	wire [4-1:0] node1715;
	wire [4-1:0] node1716;
	wire [4-1:0] node1717;
	wire [4-1:0] node1718;
	wire [4-1:0] node1723;
	wire [4-1:0] node1726;
	wire [4-1:0] node1728;
	wire [4-1:0] node1729;
	wire [4-1:0] node1731;
	wire [4-1:0] node1733;
	wire [4-1:0] node1736;
	wire [4-1:0] node1737;
	wire [4-1:0] node1741;
	wire [4-1:0] node1742;
	wire [4-1:0] node1743;
	wire [4-1:0] node1745;
	wire [4-1:0] node1747;
	wire [4-1:0] node1748;
	wire [4-1:0] node1752;
	wire [4-1:0] node1753;
	wire [4-1:0] node1756;
	wire [4-1:0] node1757;
	wire [4-1:0] node1761;
	wire [4-1:0] node1762;
	wire [4-1:0] node1764;
	wire [4-1:0] node1768;
	wire [4-1:0] node1769;
	wire [4-1:0] node1770;
	wire [4-1:0] node1772;
	wire [4-1:0] node1773;
	wire [4-1:0] node1775;
	wire [4-1:0] node1779;
	wire [4-1:0] node1781;
	wire [4-1:0] node1782;
	wire [4-1:0] node1783;
	wire [4-1:0] node1784;
	wire [4-1:0] node1790;
	wire [4-1:0] node1791;
	wire [4-1:0] node1792;
	wire [4-1:0] node1793;
	wire [4-1:0] node1794;
	wire [4-1:0] node1796;
	wire [4-1:0] node1799;
	wire [4-1:0] node1801;
	wire [4-1:0] node1804;
	wire [4-1:0] node1806;
	wire [4-1:0] node1809;
	wire [4-1:0] node1810;
	wire [4-1:0] node1812;
	wire [4-1:0] node1813;
	wire [4-1:0] node1815;
	wire [4-1:0] node1818;
	wire [4-1:0] node1819;
	wire [4-1:0] node1823;
	wire [4-1:0] node1824;
	wire [4-1:0] node1826;
	wire [4-1:0] node1829;
	wire [4-1:0] node1832;
	wire [4-1:0] node1833;
	wire [4-1:0] node1834;
	wire [4-1:0] node1836;
	wire [4-1:0] node1838;
	wire [4-1:0] node1841;
	wire [4-1:0] node1844;
	wire [4-1:0] node1846;
	wire [4-1:0] node1849;
	wire [4-1:0] node1850;
	wire [4-1:0] node1851;
	wire [4-1:0] node1852;
	wire [4-1:0] node1853;
	wire [4-1:0] node1854;
	wire [4-1:0] node1855;
	wire [4-1:0] node1858;
	wire [4-1:0] node1860;
	wire [4-1:0] node1863;
	wire [4-1:0] node1864;
	wire [4-1:0] node1865;
	wire [4-1:0] node1868;
	wire [4-1:0] node1871;
	wire [4-1:0] node1872;
	wire [4-1:0] node1873;
	wire [4-1:0] node1877;
	wire [4-1:0] node1878;
	wire [4-1:0] node1881;
	wire [4-1:0] node1884;
	wire [4-1:0] node1886;
	wire [4-1:0] node1889;
	wire [4-1:0] node1890;
	wire [4-1:0] node1891;
	wire [4-1:0] node1892;
	wire [4-1:0] node1893;
	wire [4-1:0] node1895;
	wire [4-1:0] node1898;
	wire [4-1:0] node1901;
	wire [4-1:0] node1903;
	wire [4-1:0] node1906;
	wire [4-1:0] node1907;
	wire [4-1:0] node1909;
	wire [4-1:0] node1912;
	wire [4-1:0] node1913;
	wire [4-1:0] node1914;
	wire [4-1:0] node1919;
	wire [4-1:0] node1920;
	wire [4-1:0] node1922;
	wire [4-1:0] node1923;
	wire [4-1:0] node1927;
	wire [4-1:0] node1928;
	wire [4-1:0] node1930;
	wire [4-1:0] node1934;
	wire [4-1:0] node1935;
	wire [4-1:0] node1936;
	wire [4-1:0] node1937;
	wire [4-1:0] node1941;
	wire [4-1:0] node1942;
	wire [4-1:0] node1943;
	wire [4-1:0] node1945;
	wire [4-1:0] node1950;
	wire [4-1:0] node1951;
	wire [4-1:0] node1953;
	wire [4-1:0] node1955;
	wire [4-1:0] node1958;
	wire [4-1:0] node1959;
	wire [4-1:0] node1963;
	wire [4-1:0] node1964;
	wire [4-1:0] node1965;
	wire [4-1:0] node1966;
	wire [4-1:0] node1967;
	wire [4-1:0] node1968;
	wire [4-1:0] node1969;
	wire [4-1:0] node1973;
	wire [4-1:0] node1975;
	wire [4-1:0] node1978;
	wire [4-1:0] node1979;
	wire [4-1:0] node1982;
	wire [4-1:0] node1983;
	wire [4-1:0] node1987;
	wire [4-1:0] node1990;
	wire [4-1:0] node1991;
	wire [4-1:0] node1992;
	wire [4-1:0] node1993;
	wire [4-1:0] node1995;
	wire [4-1:0] node1999;
	wire [4-1:0] node2000;
	wire [4-1:0] node2004;
	wire [4-1:0] node2005;
	wire [4-1:0] node2006;
	wire [4-1:0] node2007;
	wire [4-1:0] node2011;
	wire [4-1:0] node2013;
	wire [4-1:0] node2016;
	wire [4-1:0] node2019;
	wire [4-1:0] node2020;
	wire [4-1:0] node2021;
	wire [4-1:0] node2022;
	wire [4-1:0] node2025;
	wire [4-1:0] node2028;
	wire [4-1:0] node2029;
	wire [4-1:0] node2032;
	wire [4-1:0] node2036;
	wire [4-1:0] node2038;
	wire [4-1:0] node2039;
	wire [4-1:0] node2040;
	wire [4-1:0] node2041;
	wire [4-1:0] node2042;
	wire [4-1:0] node2043;
	wire [4-1:0] node2044;
	wire [4-1:0] node2045;
	wire [4-1:0] node2046;
	wire [4-1:0] node2047;
	wire [4-1:0] node2052;
	wire [4-1:0] node2054;
	wire [4-1:0] node2056;
	wire [4-1:0] node2060;
	wire [4-1:0] node2062;
	wire [4-1:0] node2063;
	wire [4-1:0] node2064;
	wire [4-1:0] node2066;
	wire [4-1:0] node2070;
	wire [4-1:0] node2072;
	wire [4-1:0] node2073;
	wire [4-1:0] node2078;
	wire [4-1:0] node2079;
	wire [4-1:0] node2080;
	wire [4-1:0] node2081;
	wire [4-1:0] node2082;
	wire [4-1:0] node2084;
	wire [4-1:0] node2088;
	wire [4-1:0] node2089;
	wire [4-1:0] node2091;
	wire [4-1:0] node2096;
	wire [4-1:0] node2097;
	wire [4-1:0] node2098;
	wire [4-1:0] node2100;
	wire [4-1:0] node2102;
	wire [4-1:0] node2103;
	wire [4-1:0] node2107;
	wire [4-1:0] node2108;
	wire [4-1:0] node2109;
	wire [4-1:0] node2113;
	wire [4-1:0] node2114;
	wire [4-1:0] node2118;
	wire [4-1:0] node2119;
	wire [4-1:0] node2120;
	wire [4-1:0] node2121;
	wire [4-1:0] node2126;
	wire [4-1:0] node2127;
	wire [4-1:0] node2131;
	wire [4-1:0] node2132;
	wire [4-1:0] node2134;
	wire [4-1:0] node2135;
	wire [4-1:0] node2136;
	wire [4-1:0] node2137;
	wire [4-1:0] node2138;
	wire [4-1:0] node2139;
	wire [4-1:0] node2144;
	wire [4-1:0] node2145;
	wire [4-1:0] node2147;
	wire [4-1:0] node2152;
	wire [4-1:0] node2154;
	wire [4-1:0] node2155;
	wire [4-1:0] node2156;
	wire [4-1:0] node2157;
	wire [4-1:0] node2162;
	wire [4-1:0] node2164;
	wire [4-1:0] node2166;
	wire [4-1:0] node2169;
	wire [4-1:0] node2170;
	wire [4-1:0] node2171;
	wire [4-1:0] node2172;
	wire [4-1:0] node2173;
	wire [4-1:0] node2176;
	wire [4-1:0] node2177;
	wire [4-1:0] node2181;
	wire [4-1:0] node2182;
	wire [4-1:0] node2184;
	wire [4-1:0] node2186;
	wire [4-1:0] node2189;
	wire [4-1:0] node2190;
	wire [4-1:0] node2194;
	wire [4-1:0] node2195;
	wire [4-1:0] node2196;
	wire [4-1:0] node2198;
	wire [4-1:0] node2202;
	wire [4-1:0] node2203;
	wire [4-1:0] node2204;
	wire [4-1:0] node2206;
	wire [4-1:0] node2211;
	wire [4-1:0] node2212;
	wire [4-1:0] node2213;
	wire [4-1:0] node2214;
	wire [4-1:0] node2215;
	wire [4-1:0] node2216;
	wire [4-1:0] node2220;
	wire [4-1:0] node2223;
	wire [4-1:0] node2226;
	wire [4-1:0] node2227;
	wire [4-1:0] node2228;
	wire [4-1:0] node2231;
	wire [4-1:0] node2232;
	wire [4-1:0] node2236;
	wire [4-1:0] node2239;
	wire [4-1:0] node2240;
	wire [4-1:0] node2241;
	wire [4-1:0] node2244;
	wire [4-1:0] node2248;
	wire [4-1:0] node2250;
	wire [4-1:0] node2251;
	wire [4-1:0] node2252;
	wire [4-1:0] node2253;
	wire [4-1:0] node2254;
	wire [4-1:0] node2255;
	wire [4-1:0] node2256;
	wire [4-1:0] node2258;
	wire [4-1:0] node2262;
	wire [4-1:0] node2264;
	wire [4-1:0] node2268;
	wire [4-1:0] node2269;
	wire [4-1:0] node2270;
	wire [4-1:0] node2272;
	wire [4-1:0] node2275;
	wire [4-1:0] node2276;
	wire [4-1:0] node2277;
	wire [4-1:0] node2282;
	wire [4-1:0] node2284;
	wire [4-1:0] node2285;
	wire [4-1:0] node2289;
	wire [4-1:0] node2290;
	wire [4-1:0] node2292;
	wire [4-1:0] node2293;
	wire [4-1:0] node2294;
	wire [4-1:0] node2296;
	wire [4-1:0] node2300;
	wire [4-1:0] node2302;
	wire [4-1:0] node2304;
	wire [4-1:0] node2307;
	wire [4-1:0] node2308;
	wire [4-1:0] node2309;
	wire [4-1:0] node2310;
	wire [4-1:0] node2312;
	wire [4-1:0] node2316;
	wire [4-1:0] node2317;
	wire [4-1:0] node2321;
	wire [4-1:0] node2322;
	wire [4-1:0] node2324;
	wire [4-1:0] node2325;
	wire [4-1:0] node2329;
	wire [4-1:0] node2330;
	wire [4-1:0] node2334;
	wire [4-1:0] node2336;
	wire [4-1:0] node2337;
	wire [4-1:0] node2338;
	wire [4-1:0] node2339;
	wire [4-1:0] node2340;
	wire [4-1:0] node2341;
	wire [4-1:0] node2346;
	wire [4-1:0] node2347;
	wire [4-1:0] node2349;
	wire [4-1:0] node2353;
	wire [4-1:0] node2354;
	wire [4-1:0] node2355;
	wire [4-1:0] node2356;
	wire [4-1:0] node2359;
	wire [4-1:0] node2362;
	wire [4-1:0] node2364;
	wire [4-1:0] node2367;
	wire [4-1:0] node2368;
	wire [4-1:0] node2372;
	wire [4-1:0] node2374;
	wire [4-1:0] node2375;
	wire [4-1:0] node2376;
	wire [4-1:0] node2377;
	wire [4-1:0] node2381;
	wire [4-1:0] node2382;
	wire [4-1:0] node2386;
	wire [4-1:0] node2388;
	wire [4-1:0] node2389;

	assign outp = (inp[14]) ? node2 : 4'b0000;
		assign node2 = (inp[12]) ? node1440 : node3;
			assign node3 = (inp[3]) ? node397 : node4;
				assign node4 = (inp[0]) ? node154 : node5;
					assign node5 = (inp[4]) ? 4'b0000 : node6;
						assign node6 = (inp[11]) ? node78 : node7;
							assign node7 = (inp[7]) ? 4'b0010 : node8;
								assign node8 = (inp[9]) ? node42 : node9;
									assign node9 = (inp[5]) ? 4'b0000 : node10;
										assign node10 = (inp[13]) ? node26 : node11;
											assign node11 = (inp[15]) ? 4'b0000 : node12;
												assign node12 = (inp[1]) ? node18 : node13;
													assign node13 = (inp[8]) ? 4'b0000 : node14;
														assign node14 = (inp[10]) ? 4'b0000 : 4'b0010;
													assign node18 = (inp[8]) ? node20 : 4'b0010;
														assign node20 = (inp[6]) ? 4'b0010 : node21;
															assign node21 = (inp[10]) ? 4'b0000 : 4'b0010;
											assign node26 = (inp[15]) ? node28 : 4'b0010;
												assign node28 = (inp[8]) ? node36 : node29;
													assign node29 = (inp[10]) ? node31 : 4'b0010;
														assign node31 = (inp[6]) ? 4'b0010 : node32;
															assign node32 = (inp[1]) ? 4'b0010 : 4'b0000;
													assign node36 = (inp[1]) ? node38 : 4'b0000;
														assign node38 = (inp[6]) ? 4'b0010 : 4'b0000;
									assign node42 = (inp[5]) ? node44 : 4'b0010;
										assign node44 = (inp[13]) ? node60 : node45;
											assign node45 = (inp[15]) ? 4'b0000 : node46;
												assign node46 = (inp[8]) ? node54 : node47;
													assign node47 = (inp[10]) ? node49 : 4'b0010;
														assign node49 = (inp[6]) ? 4'b0010 : node50;
															assign node50 = (inp[1]) ? 4'b0010 : 4'b0000;
													assign node54 = (inp[1]) ? node56 : 4'b0000;
														assign node56 = (inp[10]) ? 4'b0000 : 4'b0010;
											assign node60 = (inp[15]) ? node62 : 4'b0010;
												assign node62 = (inp[8]) ? node70 : node63;
													assign node63 = (inp[10]) ? node65 : 4'b0010;
														assign node65 = (inp[1]) ? 4'b0010 : node66;
															assign node66 = (inp[6]) ? 4'b0010 : 4'b0000;
													assign node70 = (inp[1]) ? node72 : 4'b0000;
														assign node72 = (inp[10]) ? node74 : 4'b0010;
															assign node74 = (inp[6]) ? 4'b0010 : 4'b0000;
							assign node78 = (inp[7]) ? node80 : 4'b0000;
								assign node80 = (inp[5]) ? node118 : node81;
									assign node81 = (inp[9]) ? 4'b0010 : node82;
										assign node82 = (inp[13]) ? node100 : node83;
											assign node83 = (inp[15]) ? 4'b0000 : node84;
												assign node84 = (inp[8]) ? node92 : node85;
													assign node85 = (inp[6]) ? 4'b0010 : node86;
														assign node86 = (inp[10]) ? node88 : 4'b0010;
															assign node88 = (inp[1]) ? 4'b0010 : 4'b0000;
													assign node92 = (inp[1]) ? node94 : 4'b0000;
														assign node94 = (inp[6]) ? 4'b0010 : node95;
															assign node95 = (inp[10]) ? 4'b0000 : 4'b0010;
											assign node100 = (inp[15]) ? node102 : 4'b0010;
												assign node102 = (inp[1]) ? node110 : node103;
													assign node103 = (inp[8]) ? 4'b0000 : node104;
														assign node104 = (inp[10]) ? node106 : 4'b0010;
															assign node106 = (inp[6]) ? 4'b0010 : 4'b0000;
													assign node110 = (inp[10]) ? node112 : 4'b0010;
														assign node112 = (inp[8]) ? node114 : 4'b0010;
															assign node114 = (inp[6]) ? 4'b0010 : 4'b0000;
									assign node118 = (inp[9]) ? node120 : 4'b0000;
										assign node120 = (inp[15]) ? node138 : node121;
											assign node121 = (inp[13]) ? 4'b0010 : node122;
												assign node122 = (inp[8]) ? node130 : node123;
													assign node123 = (inp[10]) ? node125 : 4'b0010;
														assign node125 = (inp[6]) ? 4'b0010 : node126;
															assign node126 = (inp[1]) ? 4'b0010 : 4'b0000;
													assign node130 = (inp[1]) ? node132 : 4'b0000;
														assign node132 = (inp[6]) ? 4'b0010 : node133;
															assign node133 = (inp[10]) ? 4'b0000 : 4'b0010;
											assign node138 = (inp[13]) ? node140 : 4'b0000;
												assign node140 = (inp[1]) ? node146 : node141;
													assign node141 = (inp[8]) ? 4'b0000 : node142;
														assign node142 = (inp[10]) ? 4'b0000 : 4'b0010;
													assign node146 = (inp[6]) ? 4'b0010 : node147;
														assign node147 = (inp[10]) ? node149 : 4'b0010;
															assign node149 = (inp[8]) ? 4'b0000 : 4'b0010;
					assign node154 = (inp[7]) ? node232 : node155;
						assign node155 = (inp[4]) ? 4'b0010 : node156;
							assign node156 = (inp[9]) ? node194 : node157;
								assign node157 = (inp[11]) ? 4'b0010 : node158;
									assign node158 = (inp[5]) ? node176 : node159;
										assign node159 = (inp[13]) ? 4'b0000 : node160;
											assign node160 = (inp[15]) ? node168 : node161;
												assign node161 = (inp[1]) ? 4'b0000 : node162;
													assign node162 = (inp[8]) ? node164 : 4'b0000;
														assign node164 = (inp[6]) ? 4'b0000 : 4'b0010;
												assign node168 = (inp[1]) ? node170 : 4'b0010;
													assign node170 = (inp[6]) ? 4'b0000 : node171;
														assign node171 = (inp[8]) ? 4'b0010 : 4'b0000;
										assign node176 = (inp[13]) ? node178 : 4'b0010;
											assign node178 = (inp[1]) ? node186 : node179;
												assign node179 = (inp[15]) ? 4'b0010 : node180;
													assign node180 = (inp[8]) ? node182 : 4'b0000;
														assign node182 = (inp[6]) ? 4'b0000 : 4'b0010;
												assign node186 = (inp[15]) ? node188 : 4'b0000;
													assign node188 = (inp[8]) ? node190 : 4'b0000;
														assign node190 = (inp[6]) ? 4'b0000 : 4'b0010;
								assign node194 = (inp[11]) ? node196 : 4'b0000;
									assign node196 = (inp[5]) ? node214 : node197;
										assign node197 = (inp[13]) ? 4'b0000 : node198;
											assign node198 = (inp[15]) ? node206 : node199;
												assign node199 = (inp[8]) ? node201 : 4'b0000;
													assign node201 = (inp[1]) ? 4'b0000 : node202;
														assign node202 = (inp[6]) ? 4'b0000 : 4'b0010;
												assign node206 = (inp[1]) ? node208 : 4'b0010;
													assign node208 = (inp[8]) ? node210 : 4'b0000;
														assign node210 = (inp[6]) ? 4'b0000 : 4'b0010;
										assign node214 = (inp[13]) ? node216 : 4'b0010;
											assign node216 = (inp[15]) ? node224 : node217;
												assign node217 = (inp[8]) ? node219 : 4'b0000;
													assign node219 = (inp[1]) ? 4'b0000 : node220;
														assign node220 = (inp[6]) ? 4'b0000 : 4'b0010;
												assign node224 = (inp[1]) ? node226 : 4'b0010;
													assign node226 = (inp[8]) ? node228 : 4'b0000;
														assign node228 = (inp[6]) ? 4'b0000 : 4'b0010;
						assign node232 = (inp[4]) ? node322 : node233;
							assign node233 = (inp[9]) ? node257 : node234;
								assign node234 = (inp[5]) ? 4'b0000 : node235;
									assign node235 = (inp[13]) ? node237 : 4'b0000;
										assign node237 = (inp[11]) ? 4'b0000 : node238;
											assign node238 = (inp[1]) ? node246 : node239;
												assign node239 = (inp[6]) ? node241 : 4'b0000;
													assign node241 = (inp[15]) ? 4'b0000 : node242;
														assign node242 = (inp[8]) ? 4'b0000 : 4'b0010;
												assign node246 = (inp[15]) ? node248 : 4'b0010;
													assign node248 = (inp[6]) ? 4'b0010 : node249;
														assign node249 = (inp[10]) ? 4'b0000 : node250;
															assign node250 = (inp[8]) ? 4'b0000 : 4'b0010;
								assign node257 = (inp[11]) ? node277 : node258;
									assign node258 = (inp[1]) ? 4'b0010 : node259;
										assign node259 = (inp[5]) ? node261 : 4'b0010;
											assign node261 = (inp[13]) ? 4'b0010 : node262;
												assign node262 = (inp[15]) ? node270 : node263;
													assign node263 = (inp[10]) ? node265 : 4'b0010;
														assign node265 = (inp[6]) ? 4'b0010 : node266;
															assign node266 = (inp[8]) ? 4'b0000 : 4'b0010;
													assign node270 = (inp[6]) ? node272 : 4'b0000;
														assign node272 = (inp[8]) ? 4'b0000 : 4'b0010;
									assign node277 = (inp[13]) ? node291 : node278;
										assign node278 = (inp[15]) ? 4'b0000 : node279;
											assign node279 = (inp[5]) ? 4'b0000 : node280;
												assign node280 = (inp[1]) ? node282 : 4'b0000;
													assign node282 = (inp[6]) ? 4'b0010 : node283;
														assign node283 = (inp[8]) ? 4'b0000 : node284;
															assign node284 = (inp[10]) ? 4'b0000 : 4'b0010;
										assign node291 = (inp[5]) ? node303 : node292;
											assign node292 = (inp[15]) ? node294 : 4'b0010;
												assign node294 = (inp[1]) ? 4'b0010 : node295;
													assign node295 = (inp[6]) ? 4'b0010 : node296;
														assign node296 = (inp[8]) ? node298 : 4'b0010;
															assign node298 = (inp[10]) ? 4'b0000 : 4'b0010;
											assign node303 = (inp[1]) ? node313 : node304;
												assign node304 = (inp[15]) ? 4'b0000 : node305;
													assign node305 = (inp[10]) ? 4'b0000 : node306;
														assign node306 = (inp[8]) ? 4'b0000 : node307;
															assign node307 = (inp[6]) ? 4'b0010 : 4'b0000;
												assign node313 = (inp[6]) ? 4'b0010 : node314;
													assign node314 = (inp[15]) ? node316 : 4'b0010;
														assign node316 = (inp[8]) ? 4'b0000 : node317;
															assign node317 = (inp[10]) ? 4'b0000 : 4'b0010;
							assign node322 = (inp[11]) ? node360 : node323;
								assign node323 = (inp[9]) ? 4'b0000 : node324;
									assign node324 = (inp[13]) ? node342 : node325;
										assign node325 = (inp[5]) ? 4'b0010 : node326;
											assign node326 = (inp[1]) ? node334 : node327;
												assign node327 = (inp[15]) ? 4'b0010 : node328;
													assign node328 = (inp[8]) ? node330 : 4'b0000;
														assign node330 = (inp[6]) ? 4'b0000 : 4'b0010;
												assign node334 = (inp[6]) ? 4'b0000 : node335;
													assign node335 = (inp[8]) ? node337 : 4'b0000;
														assign node337 = (inp[15]) ? 4'b0010 : 4'b0000;
										assign node342 = (inp[5]) ? node344 : 4'b0000;
											assign node344 = (inp[1]) ? node352 : node345;
												assign node345 = (inp[15]) ? 4'b0010 : node346;
													assign node346 = (inp[8]) ? node348 : 4'b0000;
														assign node348 = (inp[6]) ? 4'b0000 : 4'b0010;
												assign node352 = (inp[6]) ? 4'b0000 : node353;
													assign node353 = (inp[8]) ? node355 : 4'b0000;
														assign node355 = (inp[15]) ? 4'b0010 : 4'b0000;
								assign node360 = (inp[9]) ? node362 : 4'b0010;
									assign node362 = (inp[5]) ? node380 : node363;
										assign node363 = (inp[13]) ? 4'b0000 : node364;
											assign node364 = (inp[15]) ? node372 : node365;
												assign node365 = (inp[6]) ? 4'b0000 : node366;
													assign node366 = (inp[8]) ? node368 : 4'b0000;
														assign node368 = (inp[1]) ? 4'b0000 : 4'b0010;
												assign node372 = (inp[1]) ? node374 : 4'b0010;
													assign node374 = (inp[6]) ? 4'b0000 : node375;
														assign node375 = (inp[8]) ? 4'b0010 : 4'b0000;
										assign node380 = (inp[13]) ? node382 : 4'b0010;
											assign node382 = (inp[1]) ? node390 : node383;
												assign node383 = (inp[15]) ? 4'b0010 : node384;
													assign node384 = (inp[8]) ? node386 : 4'b0000;
														assign node386 = (inp[6]) ? 4'b0000 : 4'b0010;
												assign node390 = (inp[8]) ? node392 : 4'b0000;
													assign node392 = (inp[6]) ? 4'b0000 : node393;
														assign node393 = (inp[15]) ? 4'b0010 : 4'b0000;
				assign node397 = (inp[0]) ? node545 : node398;
					assign node398 = (inp[4]) ? node400 : 4'b0010;
						assign node400 = (inp[7]) ? node478 : node401;
							assign node401 = (inp[11]) ? 4'b0000 : node402;
								assign node402 = (inp[9]) ? node440 : node403;
									assign node403 = (inp[5]) ? 4'b0000 : node404;
										assign node404 = (inp[13]) ? node422 : node405;
											assign node405 = (inp[15]) ? 4'b0000 : node406;
												assign node406 = (inp[1]) ? node414 : node407;
													assign node407 = (inp[8]) ? 4'b0000 : node408;
														assign node408 = (inp[10]) ? node410 : 4'b0010;
															assign node410 = (inp[6]) ? 4'b0010 : 4'b0000;
													assign node414 = (inp[6]) ? 4'b0010 : node415;
														assign node415 = (inp[8]) ? node417 : 4'b0010;
															assign node417 = (inp[10]) ? 4'b0000 : 4'b0010;
											assign node422 = (inp[15]) ? node424 : 4'b0010;
												assign node424 = (inp[1]) ? node432 : node425;
													assign node425 = (inp[8]) ? 4'b0000 : node426;
														assign node426 = (inp[2]) ? node428 : 4'b0010;
															assign node428 = (inp[6]) ? 4'b0010 : 4'b0000;
													assign node432 = (inp[10]) ? node434 : 4'b0010;
														assign node434 = (inp[6]) ? 4'b0010 : node435;
															assign node435 = (inp[8]) ? 4'b0000 : 4'b0010;
									assign node440 = (inp[5]) ? node442 : 4'b0010;
										assign node442 = (inp[13]) ? node462 : node443;
											assign node443 = (inp[15]) ? 4'b0000 : node444;
												assign node444 = (inp[8]) ? node454 : node445;
													assign node445 = (inp[1]) ? 4'b0010 : node446;
														assign node446 = (inp[2]) ? 4'b0010 : node447;
															assign node447 = (inp[6]) ? 4'b0010 : node448;
																assign node448 = (inp[10]) ? 4'b0000 : 4'b0010;
													assign node454 = (inp[1]) ? node456 : 4'b0000;
														assign node456 = (inp[6]) ? 4'b0010 : node457;
															assign node457 = (inp[10]) ? 4'b0000 : 4'b0010;
											assign node462 = (inp[15]) ? node464 : 4'b0010;
												assign node464 = (inp[1]) ? node470 : node465;
													assign node465 = (inp[8]) ? 4'b0000 : node466;
														assign node466 = (inp[10]) ? 4'b0000 : 4'b0010;
													assign node470 = (inp[10]) ? node472 : 4'b0010;
														assign node472 = (inp[8]) ? node474 : 4'b0010;
															assign node474 = (inp[6]) ? 4'b0010 : 4'b0000;
							assign node478 = (inp[11]) ? node480 : 4'b0010;
								assign node480 = (inp[9]) ? node514 : node481;
									assign node481 = (inp[5]) ? 4'b0000 : node482;
										assign node482 = (inp[15]) ? node502 : node483;
											assign node483 = (inp[13]) ? 4'b0010 : node484;
												assign node484 = (inp[8]) ? node494 : node485;
													assign node485 = (inp[2]) ? node487 : 4'b0010;
														assign node487 = (inp[6]) ? 4'b0010 : node488;
															assign node488 = (inp[1]) ? 4'b0010 : node489;
																assign node489 = (inp[10]) ? 4'b0000 : 4'b0010;
													assign node494 = (inp[1]) ? node496 : 4'b0000;
														assign node496 = (inp[10]) ? node498 : 4'b0010;
															assign node498 = (inp[6]) ? 4'b0010 : 4'b0000;
											assign node502 = (inp[13]) ? node504 : 4'b0000;
												assign node504 = (inp[8]) ? node506 : 4'b0010;
													assign node506 = (inp[1]) ? node508 : 4'b0000;
														assign node508 = (inp[10]) ? node510 : 4'b0010;
															assign node510 = (inp[6]) ? 4'b0010 : 4'b0000;
									assign node514 = (inp[5]) ? node516 : 4'b0010;
										assign node516 = (inp[13]) ? node534 : node517;
											assign node517 = (inp[15]) ? 4'b0000 : node518;
												assign node518 = (inp[1]) ? node526 : node519;
													assign node519 = (inp[8]) ? 4'b0000 : node520;
														assign node520 = (inp[6]) ? 4'b0010 : node521;
															assign node521 = (inp[10]) ? 4'b0000 : 4'b0010;
													assign node526 = (inp[6]) ? 4'b0010 : node527;
														assign node527 = (inp[10]) ? node529 : 4'b0010;
															assign node529 = (inp[8]) ? 4'b0000 : 4'b0010;
											assign node534 = (inp[15]) ? node536 : 4'b0010;
												assign node536 = (inp[8]) ? node538 : 4'b0010;
													assign node538 = (inp[1]) ? node540 : 4'b0000;
														assign node540 = (inp[10]) ? node542 : 4'b0010;
															assign node542 = (inp[6]) ? 4'b0010 : 4'b0000;
					assign node545 = (inp[9]) ? node937 : node546;
						assign node546 = (inp[7]) ? node656 : node547;
							assign node547 = (inp[4]) ? node595 : node548;
								assign node548 = (inp[11]) ? node578 : node549;
									assign node549 = (inp[13]) ? node565 : node550;
										assign node550 = (inp[5]) ? node558 : node551;
											assign node551 = (inp[15]) ? node553 : 4'b1000;
												assign node553 = (inp[6]) ? 4'b1000 : node554;
													assign node554 = (inp[1]) ? 4'b1000 : 4'b0010;
											assign node558 = (inp[1]) ? node560 : 4'b0010;
												assign node560 = (inp[15]) ? node562 : 4'b1000;
													assign node562 = (inp[6]) ? 4'b1000 : 4'b0010;
										assign node565 = (inp[1]) ? node567 : 4'b1000;
											assign node567 = (inp[5]) ? 4'b1000 : node568;
												assign node568 = (inp[6]) ? 4'b1010 : node569;
													assign node569 = (inp[15]) ? 4'b1000 : node570;
														assign node570 = (inp[10]) ? node572 : 4'b1010;
															assign node572 = (inp[8]) ? 4'b1000 : 4'b1010;
									assign node578 = (inp[13]) ? node580 : 4'b0010;
										assign node580 = (inp[1]) ? node588 : node581;
											assign node581 = (inp[5]) ? 4'b0010 : node582;
												assign node582 = (inp[6]) ? 4'b1000 : node583;
													assign node583 = (inp[15]) ? 4'b0010 : 4'b1000;
											assign node588 = (inp[15]) ? node590 : 4'b1000;
												assign node590 = (inp[5]) ? node592 : 4'b1000;
													assign node592 = (inp[6]) ? 4'b1000 : 4'b0010;
								assign node595 = (inp[11]) ? node635 : node596;
									assign node596 = (inp[13]) ? node622 : node597;
										assign node597 = (inp[5]) ? node611 : node598;
											assign node598 = (inp[1]) ? 4'b0010 : node599;
												assign node599 = (inp[15]) ? node605 : node600;
													assign node600 = (inp[6]) ? 4'b0010 : node601;
														assign node601 = (inp[10]) ? 4'b0000 : 4'b0010;
													assign node605 = (inp[8]) ? 4'b0000 : node606;
														assign node606 = (inp[6]) ? 4'b0010 : 4'b0000;
											assign node611 = (inp[1]) ? node613 : 4'b0000;
												assign node613 = (inp[15]) ? 4'b0000 : node614;
													assign node614 = (inp[6]) ? 4'b0010 : node615;
														assign node615 = (inp[10]) ? 4'b0000 : node616;
															assign node616 = (inp[8]) ? 4'b0000 : 4'b0010;
										assign node622 = (inp[1]) ? 4'b0010 : node623;
											assign node623 = (inp[5]) ? node625 : 4'b0010;
												assign node625 = (inp[15]) ? node627 : 4'b0010;
													assign node627 = (inp[8]) ? node629 : 4'b0010;
														assign node629 = (inp[10]) ? node631 : 4'b0010;
															assign node631 = (inp[6]) ? 4'b0010 : 4'b0000;
									assign node635 = (inp[5]) ? 4'b0000 : node636;
										assign node636 = (inp[13]) ? node638 : 4'b0000;
											assign node638 = (inp[1]) ? node646 : node639;
												assign node639 = (inp[6]) ? node641 : 4'b0000;
													assign node641 = (inp[10]) ? node643 : 4'b0000;
														assign node643 = (inp[15]) ? 4'b0000 : 4'b0010;
												assign node646 = (inp[15]) ? node648 : 4'b0010;
													assign node648 = (inp[6]) ? 4'b0010 : node649;
														assign node649 = (inp[10]) ? 4'b0000 : node650;
															assign node650 = (inp[8]) ? 4'b0000 : 4'b0010;
							assign node656 = (inp[4]) ? node804 : node657;
								assign node657 = (inp[15]) ? node735 : node658;
									assign node658 = (inp[11]) ? node702 : node659;
										assign node659 = (inp[13]) ? node681 : node660;
											assign node660 = (inp[1]) ? node670 : node661;
												assign node661 = (inp[6]) ? node665 : node662;
													assign node662 = (inp[5]) ? 4'b1010 : 4'b0000;
													assign node665 = (inp[5]) ? 4'b0000 : node666;
														assign node666 = (inp[8]) ? 4'b0000 : 4'b0010;
												assign node670 = (inp[6]) ? node678 : node671;
													assign node671 = (inp[8]) ? node673 : 4'b0010;
														assign node673 = (inp[5]) ? node675 : 4'b0010;
															assign node675 = (inp[10]) ? 4'b0000 : 4'b0010;
													assign node678 = (inp[5]) ? 4'b0010 : 4'b0000;
											assign node681 = (inp[1]) ? node689 : node682;
												assign node682 = (inp[5]) ? node686 : node683;
													assign node683 = (inp[6]) ? 4'b1000 : 4'b0010;
													assign node686 = (inp[6]) ? 4'b0010 : 4'b0000;
												assign node689 = (inp[5]) ? node695 : node690;
													assign node690 = (inp[6]) ? 4'b1010 : node691;
														assign node691 = (inp[8]) ? 4'b1010 : 4'b1000;
													assign node695 = (inp[6]) ? 4'b1000 : node696;
														assign node696 = (inp[10]) ? node698 : 4'b1010;
															assign node698 = (inp[8]) ? 4'b1000 : 4'b1010;
										assign node702 = (inp[13]) ? node716 : node703;
											assign node703 = (inp[1]) ? node709 : node704;
												assign node704 = (inp[6]) ? 4'b1010 : node705;
													assign node705 = (inp[5]) ? 4'b1000 : 4'b1010;
												assign node709 = (inp[6]) ? node713 : node710;
													assign node710 = (inp[5]) ? 4'b1010 : 4'b0000;
													assign node713 = (inp[5]) ? 4'b0000 : 4'b0010;
											assign node716 = (inp[1]) ? node728 : node717;
												assign node717 = (inp[6]) ? node723 : node718;
													assign node718 = (inp[5]) ? 4'b0010 : node719;
														assign node719 = (inp[8]) ? 4'b0010 : 4'b0000;
													assign node723 = (inp[5]) ? 4'b0000 : node724;
														assign node724 = (inp[8]) ? 4'b0000 : 4'b0010;
												assign node728 = (inp[5]) ? node732 : node729;
													assign node729 = (inp[6]) ? 4'b1010 : 4'b1000;
													assign node732 = (inp[6]) ? 4'b1000 : 4'b0010;
									assign node735 = (inp[13]) ? node767 : node736;
										assign node736 = (inp[1]) ? node754 : node737;
											assign node737 = (inp[11]) ? node743 : node738;
												assign node738 = (inp[6]) ? 4'b0000 : node739;
													assign node739 = (inp[5]) ? 4'b1010 : 4'b0000;
												assign node743 = (inp[5]) ? node749 : node744;
													assign node744 = (inp[6]) ? 4'b1010 : node745;
														assign node745 = (inp[10]) ? 4'b1000 : 4'b1010;
													assign node749 = (inp[6]) ? node751 : 4'b1000;
														assign node751 = (inp[8]) ? 4'b1000 : 4'b1010;
											assign node754 = (inp[5]) ? node760 : node755;
												assign node755 = (inp[11]) ? 4'b0000 : node756;
													assign node756 = (inp[6]) ? 4'b0000 : 4'b0010;
												assign node760 = (inp[6]) ? node764 : node761;
													assign node761 = (inp[11]) ? 4'b1010 : 4'b0000;
													assign node764 = (inp[11]) ? 4'b0000 : 4'b0010;
										assign node767 = (inp[1]) ? node789 : node768;
											assign node768 = (inp[5]) ? node780 : node769;
												assign node769 = (inp[6]) ? node777 : node770;
													assign node770 = (inp[10]) ? node772 : 4'b0010;
														assign node772 = (inp[8]) ? node774 : 4'b0010;
															assign node774 = (inp[11]) ? 4'b0010 : 4'b0000;
													assign node777 = (inp[11]) ? 4'b0000 : 4'b1000;
												assign node780 = (inp[6]) ? 4'b0010 : node781;
													assign node781 = (inp[10]) ? 4'b0000 : node782;
														assign node782 = (inp[11]) ? node784 : 4'b0000;
															assign node784 = (inp[8]) ? 4'b0000 : 4'b0010;
											assign node789 = (inp[5]) ? node795 : node790;
												assign node790 = (inp[11]) ? node792 : 4'b1010;
													assign node792 = (inp[6]) ? 4'b1010 : 4'b0010;
												assign node795 = (inp[11]) ? node797 : 4'b1000;
													assign node797 = (inp[6]) ? 4'b1000 : node798;
														assign node798 = (inp[8]) ? 4'b0000 : node799;
															assign node799 = (inp[10]) ? 4'b0000 : 4'b0010;
								assign node804 = (inp[13]) ? node868 : node805;
									assign node805 = (inp[1]) ? node833 : node806;
										assign node806 = (inp[6]) ? node820 : node807;
											assign node807 = (inp[11]) ? node815 : node808;
												assign node808 = (inp[5]) ? 4'b1010 : node809;
													assign node809 = (inp[8]) ? node811 : 4'b1000;
														assign node811 = (inp[15]) ? 4'b1010 : 4'b1000;
												assign node815 = (inp[5]) ? 4'b1000 : node816;
													assign node816 = (inp[15]) ? 4'b1000 : 4'b1010;
											assign node820 = (inp[11]) ? node826 : node821;
												assign node821 = (inp[5]) ? node823 : 4'b1000;
													assign node823 = (inp[15]) ? 4'b1010 : 4'b1000;
												assign node826 = (inp[5]) ? node828 : 4'b1010;
													assign node828 = (inp[15]) ? 4'b1000 : node829;
														assign node829 = (inp[8]) ? 4'b1000 : 4'b1010;
										assign node833 = (inp[15]) ? node847 : node834;
											assign node834 = (inp[5]) ? node842 : node835;
												assign node835 = (inp[11]) ? node837 : 4'b1010;
													assign node837 = (inp[8]) ? node839 : 4'b1000;
														assign node839 = (inp[6]) ? 4'b1000 : 4'b1010;
												assign node842 = (inp[11]) ? 4'b1010 : node843;
													assign node843 = (inp[6]) ? 4'b1010 : 4'b1000;
											assign node847 = (inp[11]) ? node857 : node848;
												assign node848 = (inp[5]) ? 4'b1000 : node849;
													assign node849 = (inp[6]) ? 4'b1010 : node850;
														assign node850 = (inp[8]) ? 4'b1000 : node851;
															assign node851 = (inp[10]) ? 4'b1000 : 4'b1010;
												assign node857 = (inp[6]) ? node865 : node858;
													assign node858 = (inp[8]) ? node860 : 4'b1010;
														assign node860 = (inp[10]) ? node862 : 4'b1010;
															assign node862 = (inp[5]) ? 4'b1000 : 4'b1010;
													assign node865 = (inp[5]) ? 4'b1010 : 4'b1000;
									assign node868 = (inp[1]) ? node916 : node869;
										assign node869 = (inp[11]) ? node881 : node870;
											assign node870 = (inp[5]) ? node878 : node871;
												assign node871 = (inp[6]) ? node873 : 4'b0000;
													assign node873 = (inp[15]) ? node875 : 4'b0010;
														assign node875 = (inp[8]) ? 4'b0000 : 4'b0010;
												assign node878 = (inp[6]) ? 4'b0000 : 4'b1010;
											assign node881 = (inp[5]) ? node891 : node882;
												assign node882 = (inp[6]) ? 4'b1010 : node883;
													assign node883 = (inp[15]) ? 4'b1000 : node884;
														assign node884 = (inp[8]) ? node886 : 4'b1010;
															assign node886 = (inp[10]) ? 4'b1000 : 4'b1010;
												assign node891 = (inp[2]) ? node905 : node892;
													assign node892 = (inp[10]) ? node898 : node893;
														assign node893 = (inp[8]) ? node895 : 4'b1000;
															assign node895 = (inp[15]) ? 4'b1010 : 4'b1000;
														assign node898 = (inp[6]) ? node900 : 4'b1000;
															assign node900 = (inp[15]) ? 4'b1000 : node901;
																assign node901 = (inp[8]) ? 4'b1000 : 4'b1010;
													assign node905 = (inp[6]) ? node911 : node906;
														assign node906 = (inp[15]) ? node908 : 4'b1000;
															assign node908 = (inp[8]) ? 4'b1010 : 4'b1000;
														assign node911 = (inp[8]) ? 4'b1000 : node912;
															assign node912 = (inp[15]) ? 4'b1000 : 4'b1010;
										assign node916 = (inp[5]) ? node926 : node917;
											assign node917 = (inp[6]) ? 4'b0010 : node918;
												assign node918 = (inp[15]) ? node920 : 4'b0000;
													assign node920 = (inp[11]) ? 4'b0000 : node921;
														assign node921 = (inp[8]) ? 4'b0010 : 4'b0000;
											assign node926 = (inp[6]) ? 4'b0000 : node927;
												assign node927 = (inp[11]) ? 4'b1010 : node928;
													assign node928 = (inp[15]) ? node930 : 4'b0010;
														assign node930 = (inp[8]) ? node932 : 4'b0010;
															assign node932 = (inp[10]) ? 4'b0000 : 4'b0010;
						assign node937 = (inp[7]) ? node1109 : node938;
							assign node938 = (inp[4]) ? node1032 : node939;
								assign node939 = (inp[11]) ? node989 : node940;
									assign node940 = (inp[13]) ? node962 : node941;
										assign node941 = (inp[5]) ? node951 : node942;
											assign node942 = (inp[1]) ? node944 : 4'b1010;
												assign node944 = (inp[6]) ? 4'b1000 : node945;
													assign node945 = (inp[8]) ? 4'b1010 : node946;
														assign node946 = (inp[15]) ? 4'b1010 : 4'b1000;
											assign node951 = (inp[6]) ? 4'b1010 : node952;
												assign node952 = (inp[15]) ? node954 : 4'b1010;
													assign node954 = (inp[1]) ? 4'b1010 : node955;
														assign node955 = (inp[8]) ? 4'b1000 : node956;
															assign node956 = (inp[10]) ? 4'b1000 : 4'b1010;
										assign node962 = (inp[1]) ? node978 : node963;
											assign node963 = (inp[6]) ? node971 : node964;
												assign node964 = (inp[15]) ? node966 : 4'b1000;
													assign node966 = (inp[8]) ? node968 : 4'b1000;
														assign node968 = (inp[5]) ? 4'b1010 : 4'b1000;
												assign node971 = (inp[5]) ? 4'b1000 : node972;
													assign node972 = (inp[8]) ? 4'b1000 : node973;
														assign node973 = (inp[15]) ? 4'b1000 : 4'b1010;
											assign node978 = (inp[6]) ? 4'b1010 : node979;
												assign node979 = (inp[5]) ? node981 : 4'b1010;
													assign node981 = (inp[15]) ? 4'b1000 : node982;
														assign node982 = (inp[8]) ? 4'b1000 : node983;
															assign node983 = (inp[10]) ? 4'b1000 : 4'b1010;
									assign node989 = (inp[13]) ? node1015 : node990;
										assign node990 = (inp[1]) ? node1000 : node991;
											assign node991 = (inp[5]) ? 4'b1000 : node992;
												assign node992 = (inp[8]) ? 4'b1000 : node993;
													assign node993 = (inp[6]) ? node995 : 4'b1000;
														assign node995 = (inp[15]) ? 4'b1000 : 4'b1010;
											assign node1000 = (inp[5]) ? node1010 : node1001;
												assign node1001 = (inp[10]) ? node1003 : 4'b1010;
													assign node1003 = (inp[15]) ? node1005 : 4'b1010;
														assign node1005 = (inp[6]) ? 4'b1010 : node1006;
															assign node1006 = (inp[8]) ? 4'b1000 : 4'b1010;
												assign node1010 = (inp[6]) ? node1012 : 4'b1000;
													assign node1012 = (inp[15]) ? 4'b1000 : 4'b1010;
										assign node1015 = (inp[1]) ? node1023 : node1016;
											assign node1016 = (inp[6]) ? node1018 : 4'b1010;
												assign node1018 = (inp[15]) ? 4'b1010 : node1019;
													assign node1019 = (inp[5]) ? 4'b1010 : 4'b1000;
											assign node1023 = (inp[6]) ? 4'b1000 : node1024;
												assign node1024 = (inp[5]) ? node1026 : 4'b1000;
													assign node1026 = (inp[15]) ? 4'b1010 : node1027;
														assign node1027 = (inp[8]) ? 4'b1010 : 4'b1000;
								assign node1032 = (inp[13]) ? node1064 : node1033;
									assign node1033 = (inp[11]) ? node1049 : node1034;
										assign node1034 = (inp[5]) ? node1042 : node1035;
											assign node1035 = (inp[6]) ? 4'b1000 : node1036;
												assign node1036 = (inp[1]) ? 4'b1000 : node1037;
													assign node1037 = (inp[15]) ? 4'b0010 : 4'b1000;
											assign node1042 = (inp[1]) ? node1044 : 4'b0010;
												assign node1044 = (inp[15]) ? node1046 : 4'b1000;
													assign node1046 = (inp[6]) ? 4'b1000 : 4'b0010;
										assign node1049 = (inp[5]) ? node1051 : 4'b0010;
											assign node1051 = (inp[1]) ? 4'b0010 : node1052;
												assign node1052 = (inp[15]) ? node1058 : node1053;
													assign node1053 = (inp[10]) ? node1055 : 4'b0010;
														assign node1055 = (inp[6]) ? 4'b0010 : 4'b0000;
													assign node1058 = (inp[8]) ? 4'b0000 : node1059;
														assign node1059 = (inp[6]) ? 4'b0010 : 4'b0000;
									assign node1064 = (inp[11]) ? node1094 : node1065;
										assign node1065 = (inp[1]) ? node1081 : node1066;
											assign node1066 = (inp[5]) ? 4'b1000 : node1067;
												assign node1067 = (inp[6]) ? node1075 : node1068;
													assign node1068 = (inp[15]) ? 4'b1000 : node1069;
														assign node1069 = (inp[10]) ? 4'b1000 : node1070;
															assign node1070 = (inp[8]) ? 4'b1000 : 4'b1010;
													assign node1075 = (inp[8]) ? node1077 : 4'b1010;
														assign node1077 = (inp[15]) ? 4'b1000 : 4'b1010;
											assign node1081 = (inp[5]) ? node1083 : 4'b1010;
												assign node1083 = (inp[6]) ? 4'b1010 : node1084;
													assign node1084 = (inp[15]) ? 4'b1000 : node1085;
														assign node1085 = (inp[2]) ? 4'b1010 : node1086;
															assign node1086 = (inp[8]) ? node1088 : 4'b1010;
																assign node1088 = (inp[10]) ? 4'b1000 : 4'b1010;
										assign node1094 = (inp[1]) ? node1102 : node1095;
											assign node1095 = (inp[5]) ? 4'b0010 : node1096;
												assign node1096 = (inp[6]) ? 4'b1000 : node1097;
													assign node1097 = (inp[15]) ? 4'b0010 : 4'b1000;
											assign node1102 = (inp[5]) ? node1104 : 4'b1000;
												assign node1104 = (inp[6]) ? 4'b1000 : node1105;
													assign node1105 = (inp[15]) ? 4'b0010 : 4'b1000;
							assign node1109 = (inp[13]) ? node1315 : node1110;
								assign node1110 = (inp[4]) ? node1196 : node1111;
									assign node1111 = (inp[1]) ? node1159 : node1112;
										assign node1112 = (inp[11]) ? node1136 : node1113;
											assign node1113 = (inp[6]) ? node1125 : node1114;
												assign node1114 = (inp[5]) ? node1120 : node1115;
													assign node1115 = (inp[15]) ? 4'b0011 : node1116;
														assign node1116 = (inp[8]) ? 4'b0011 : 4'b0001;
													assign node1120 = (inp[8]) ? 4'b0001 : node1121;
														assign node1121 = (inp[15]) ? 4'b0001 : 4'b0011;
												assign node1125 = (inp[5]) ? node1131 : node1126;
													assign node1126 = (inp[8]) ? 4'b1001 : node1127;
														assign node1127 = (inp[15]) ? 4'b1001 : 4'b1011;
													assign node1131 = (inp[8]) ? node1133 : 4'b0011;
														assign node1133 = (inp[15]) ? 4'b0001 : 4'b0011;
											assign node1136 = (inp[6]) ? node1150 : node1137;
												assign node1137 = (inp[5]) ? node1145 : node1138;
													assign node1138 = (inp[15]) ? node1140 : 4'b1010;
														assign node1140 = (inp[10]) ? node1142 : 4'b1010;
															assign node1142 = (inp[8]) ? 4'b1000 : 4'b1010;
													assign node1145 = (inp[15]) ? node1147 : 4'b1000;
														assign node1147 = (inp[8]) ? 4'b1010 : 4'b1000;
												assign node1150 = (inp[15]) ? node1156 : node1151;
													assign node1151 = (inp[8]) ? 4'b0001 : node1152;
														assign node1152 = (inp[5]) ? 4'b0011 : 4'b0001;
													assign node1156 = (inp[5]) ? 4'b0001 : 4'b0011;
										assign node1159 = (inp[15]) ? node1177 : node1160;
											assign node1160 = (inp[6]) ? node1174 : node1161;
												assign node1161 = (inp[11]) ? node1169 : node1162;
													assign node1162 = (inp[5]) ? 4'b1011 : node1163;
														assign node1163 = (inp[8]) ? node1165 : 4'b0011;
															assign node1165 = (inp[10]) ? 4'b0001 : 4'b0011;
													assign node1169 = (inp[5]) ? 4'b1001 : node1170;
														assign node1170 = (inp[8]) ? 4'b1011 : 4'b1001;
												assign node1174 = (inp[11]) ? 4'b0011 : 4'b1011;
											assign node1177 = (inp[11]) ? node1187 : node1178;
												assign node1178 = (inp[6]) ? 4'b1001 : node1179;
													assign node1179 = (inp[5]) ? node1181 : 4'b0001;
														assign node1181 = (inp[2]) ? 4'b1001 : node1182;
															assign node1182 = (inp[10]) ? 4'b1001 : 4'b1011;
												assign node1187 = (inp[6]) ? 4'b0001 : node1188;
													assign node1188 = (inp[5]) ? 4'b0011 : node1189;
														assign node1189 = (inp[8]) ? node1191 : 4'b1011;
															assign node1191 = (inp[10]) ? 4'b1001 : 4'b1011;
									assign node1196 = (inp[1]) ? node1260 : node1197;
										assign node1197 = (inp[11]) ? node1227 : node1198;
											assign node1198 = (inp[8]) ? node1210 : node1199;
												assign node1199 = (inp[15]) ? node1203 : node1200;
													assign node1200 = (inp[5]) ? 4'b1000 : 4'b1010;
													assign node1203 = (inp[6]) ? 4'b1010 : node1204;
														assign node1204 = (inp[5]) ? 4'b0010 : node1205;
															assign node1205 = (inp[10]) ? 4'b1000 : 4'b1010;
												assign node1210 = (inp[2]) ? node1220 : node1211;
													assign node1211 = (inp[15]) ? node1215 : node1212;
														assign node1212 = (inp[5]) ? 4'b1000 : 4'b1010;
														assign node1215 = (inp[5]) ? node1217 : 4'b1000;
															assign node1217 = (inp[6]) ? 4'b1010 : 4'b0010;
													assign node1220 = (inp[15]) ? node1224 : node1221;
														assign node1221 = (inp[5]) ? 4'b1000 : 4'b1010;
														assign node1224 = (inp[5]) ? 4'b1010 : 4'b1000;
											assign node1227 = (inp[5]) ? node1241 : node1228;
												assign node1228 = (inp[6]) ? node1236 : node1229;
													assign node1229 = (inp[15]) ? 4'b0000 : node1230;
														assign node1230 = (inp[8]) ? node1232 : 4'b0010;
															assign node1232 = (inp[2]) ? 4'b0000 : 4'b0010;
													assign node1236 = (inp[8]) ? 4'b1000 : node1237;
														assign node1237 = (inp[15]) ? 4'b1000 : 4'b1010;
												assign node1241 = (inp[10]) ? node1249 : node1242;
													assign node1242 = (inp[15]) ? node1246 : node1243;
														assign node1243 = (inp[8]) ? 4'b0010 : 4'b0000;
														assign node1246 = (inp[8]) ? 4'b0000 : 4'b0010;
													assign node1249 = (inp[6]) ? node1255 : node1250;
														assign node1250 = (inp[8]) ? 4'b0010 : node1251;
															assign node1251 = (inp[15]) ? 4'b0010 : 4'b0000;
														assign node1255 = (inp[15]) ? node1257 : 4'b0010;
															assign node1257 = (inp[8]) ? 4'b0000 : 4'b0010;
										assign node1260 = (inp[11]) ? node1288 : node1261;
											assign node1261 = (inp[6]) ? node1285 : node1262;
												assign node1262 = (inp[10]) ? node1274 : node1263;
													assign node1263 = (inp[15]) ? node1269 : node1264;
														assign node1264 = (inp[8]) ? node1266 : 4'b0011;
															assign node1266 = (inp[5]) ? 4'b0011 : 4'b0001;
														assign node1269 = (inp[8]) ? node1271 : 4'b0001;
															assign node1271 = (inp[5]) ? 4'b0001 : 4'b0011;
													assign node1274 = (inp[15]) ? node1280 : node1275;
														assign node1275 = (inp[8]) ? 4'b0001 : node1276;
															assign node1276 = (inp[5]) ? 4'b0011 : 4'b0001;
														assign node1280 = (inp[5]) ? 4'b0001 : node1281;
															assign node1281 = (inp[8]) ? 4'b0011 : 4'b0001;
												assign node1285 = (inp[15]) ? 4'b1001 : 4'b1011;
											assign node1288 = (inp[6]) ? node1312 : node1289;
												assign node1289 = (inp[10]) ? node1301 : node1290;
													assign node1290 = (inp[15]) ? node1296 : node1291;
														assign node1291 = (inp[8]) ? 4'b1010 : node1292;
															assign node1292 = (inp[5]) ? 4'b1000 : 4'b1010;
														assign node1296 = (inp[8]) ? node1298 : 4'b1010;
															assign node1298 = (inp[5]) ? 4'b1010 : 4'b1000;
													assign node1301 = (inp[15]) ? node1307 : node1302;
														assign node1302 = (inp[5]) ? node1304 : 4'b1010;
															assign node1304 = (inp[8]) ? 4'b1010 : 4'b1000;
														assign node1307 = (inp[5]) ? node1309 : 4'b1000;
															assign node1309 = (inp[8]) ? 4'b1000 : 4'b1010;
												assign node1312 = (inp[15]) ? 4'b0001 : 4'b0011;
								assign node1315 = (inp[6]) ? node1423 : node1316;
									assign node1316 = (inp[1]) ? node1408 : node1317;
										assign node1317 = (inp[4]) ? node1369 : node1318;
											assign node1318 = (inp[10]) ? node1344 : node1319;
												assign node1319 = (inp[5]) ? node1333 : node1320;
													assign node1320 = (inp[15]) ? node1328 : node1321;
														assign node1321 = (inp[11]) ? node1325 : node1322;
															assign node1322 = (inp[8]) ? 4'b0010 : 4'b0000;
															assign node1325 = (inp[8]) ? 4'b1000 : 4'b1010;
														assign node1328 = (inp[11]) ? 4'b0010 : node1329;
															assign node1329 = (inp[8]) ? 4'b0000 : 4'b0010;
													assign node1333 = (inp[11]) ? node1337 : node1334;
														assign node1334 = (inp[8]) ? 4'b1010 : 4'b1000;
														assign node1337 = (inp[8]) ? node1341 : node1338;
															assign node1338 = (inp[15]) ? 4'b0010 : 4'b0000;
															assign node1341 = (inp[15]) ? 4'b0000 : 4'b0010;
												assign node1344 = (inp[5]) ? node1356 : node1345;
													assign node1345 = (inp[11]) ? node1351 : node1346;
														assign node1346 = (inp[15]) ? 4'b0000 : node1347;
															assign node1347 = (inp[8]) ? 4'b0010 : 4'b0000;
														assign node1351 = (inp[15]) ? node1353 : 4'b1000;
															assign node1353 = (inp[8]) ? 4'b0000 : 4'b0010;
													assign node1356 = (inp[11]) ? node1364 : node1357;
														assign node1357 = (inp[15]) ? node1361 : node1358;
															assign node1358 = (inp[8]) ? 4'b1000 : 4'b1010;
															assign node1361 = (inp[8]) ? 4'b1010 : 4'b1000;
														assign node1364 = (inp[2]) ? node1366 : 4'b0000;
															assign node1366 = (inp[15]) ? 4'b0000 : 4'b0010;
											assign node1369 = (inp[11]) ? node1385 : node1370;
												assign node1370 = (inp[5]) ? node1376 : node1371;
													assign node1371 = (inp[15]) ? node1373 : 4'b1011;
														assign node1373 = (inp[8]) ? 4'b1011 : 4'b1001;
													assign node1376 = (inp[15]) ? node1382 : node1377;
														assign node1377 = (inp[10]) ? 4'b1001 : node1378;
															assign node1378 = (inp[2]) ? 4'b1011 : 4'b1001;
														assign node1382 = (inp[10]) ? 4'b0001 : 4'b0011;
												assign node1385 = (inp[5]) ? node1395 : node1386;
													assign node1386 = (inp[15]) ? node1390 : node1387;
														assign node1387 = (inp[8]) ? 4'b0011 : 4'b0001;
														assign node1390 = (inp[8]) ? 4'b0001 : node1391;
															assign node1391 = (inp[10]) ? 4'b0001 : 4'b0011;
													assign node1395 = (inp[10]) ? node1401 : node1396;
														assign node1396 = (inp[15]) ? node1398 : 4'b1011;
															assign node1398 = (inp[8]) ? 4'b1011 : 4'b1001;
														assign node1401 = (inp[8]) ? node1405 : node1402;
															assign node1402 = (inp[15]) ? 4'b1001 : 4'b1011;
															assign node1405 = (inp[15]) ? 4'b1011 : 4'b1001;
										assign node1408 = (inp[11]) ? node1416 : node1409;
											assign node1409 = (inp[10]) ? node1413 : node1410;
												assign node1410 = (inp[15]) ? 4'b0111 : 4'b1111;
												assign node1413 = (inp[15]) ? 4'b0101 : 4'b1101;
											assign node1416 = (inp[15]) ? node1420 : node1417;
												assign node1417 = (inp[10]) ? 4'b1100 : 4'b1110;
												assign node1420 = (inp[10]) ? 4'b0100 : 4'b0110;
									assign node1423 = (inp[1]) ? 4'b0000 : node1424;
										assign node1424 = (inp[4]) ? node1432 : node1425;
											assign node1425 = (inp[5]) ? node1429 : node1426;
												assign node1426 = (inp[8]) ? 4'b1001 : 4'b1011;
												assign node1429 = (inp[8]) ? 4'b0001 : 4'b0011;
											assign node1432 = (inp[5]) ? node1436 : node1433;
												assign node1433 = (inp[8]) ? 4'b1000 : 4'b1010;
												assign node1436 = (inp[8]) ? 4'b0000 : 4'b0010;
			assign node1440 = (inp[0]) ? node1442 : 4'b0000;
				assign node1442 = (inp[4]) ? node2036 : node1443;
					assign node1443 = (inp[7]) ? node1637 : node1444;
						assign node1444 = (inp[3]) ? node1518 : node1445;
							assign node1445 = (inp[11]) ? 4'b0000 : node1446;
								assign node1446 = (inp[9]) ? node1480 : node1447;
									assign node1447 = (inp[5]) ? 4'b0000 : node1448;
										assign node1448 = (inp[15]) ? node1466 : node1449;
											assign node1449 = (inp[13]) ? 4'b0010 : node1450;
												assign node1450 = (inp[1]) ? node1458 : node1451;
													assign node1451 = (inp[8]) ? 4'b0000 : node1452;
														assign node1452 = (inp[10]) ? node1454 : 4'b0010;
															assign node1454 = (inp[6]) ? 4'b0010 : 4'b0000;
													assign node1458 = (inp[6]) ? 4'b0010 : node1459;
														assign node1459 = (inp[8]) ? node1461 : 4'b0010;
															assign node1461 = (inp[10]) ? 4'b0000 : 4'b0010;
											assign node1466 = (inp[13]) ? node1468 : 4'b0000;
												assign node1468 = (inp[8]) ? node1474 : node1469;
													assign node1469 = (inp[6]) ? 4'b0010 : node1470;
														assign node1470 = (inp[2]) ? 4'b0010 : 4'b0000;
													assign node1474 = (inp[1]) ? node1476 : 4'b0000;
														assign node1476 = (inp[10]) ? 4'b0000 : 4'b0010;
									assign node1480 = (inp[5]) ? node1482 : 4'b0010;
										assign node1482 = (inp[15]) ? node1500 : node1483;
											assign node1483 = (inp[13]) ? 4'b0010 : node1484;
												assign node1484 = (inp[1]) ? node1492 : node1485;
													assign node1485 = (inp[8]) ? 4'b0000 : node1486;
														assign node1486 = (inp[10]) ? node1488 : 4'b0010;
															assign node1488 = (inp[6]) ? 4'b0010 : 4'b0000;
													assign node1492 = (inp[8]) ? node1494 : 4'b0010;
														assign node1494 = (inp[10]) ? node1496 : 4'b0010;
															assign node1496 = (inp[6]) ? 4'b0010 : 4'b0000;
											assign node1500 = (inp[13]) ? node1502 : 4'b0000;
												assign node1502 = (inp[1]) ? node1510 : node1503;
													assign node1503 = (inp[8]) ? 4'b0000 : node1504;
														assign node1504 = (inp[6]) ? 4'b0010 : node1505;
															assign node1505 = (inp[10]) ? 4'b0000 : 4'b0010;
													assign node1510 = (inp[6]) ? 4'b0010 : node1511;
														assign node1511 = (inp[8]) ? node1513 : 4'b0010;
															assign node1513 = (inp[10]) ? 4'b0000 : 4'b0010;
							assign node1518 = (inp[9]) ? node1556 : node1519;
								assign node1519 = (inp[11]) ? 4'b0010 : node1520;
									assign node1520 = (inp[13]) ? node1538 : node1521;
										assign node1521 = (inp[5]) ? 4'b0010 : node1522;
											assign node1522 = (inp[15]) ? node1530 : node1523;
												assign node1523 = (inp[6]) ? 4'b0000 : node1524;
													assign node1524 = (inp[8]) ? node1526 : 4'b0000;
														assign node1526 = (inp[1]) ? 4'b0000 : 4'b0010;
												assign node1530 = (inp[1]) ? node1532 : 4'b0010;
													assign node1532 = (inp[6]) ? 4'b0000 : node1533;
														assign node1533 = (inp[8]) ? 4'b0010 : 4'b0000;
										assign node1538 = (inp[5]) ? node1540 : 4'b0000;
											assign node1540 = (inp[1]) ? node1548 : node1541;
												assign node1541 = (inp[15]) ? 4'b0010 : node1542;
													assign node1542 = (inp[8]) ? node1544 : 4'b0000;
														assign node1544 = (inp[6]) ? 4'b0000 : 4'b0010;
												assign node1548 = (inp[15]) ? node1550 : 4'b0000;
													assign node1550 = (inp[6]) ? 4'b0000 : node1551;
														assign node1551 = (inp[8]) ? 4'b0010 : 4'b0000;
								assign node1556 = (inp[5]) ? node1598 : node1557;
									assign node1557 = (inp[11]) ? node1581 : node1558;
										assign node1558 = (inp[13]) ? node1570 : node1559;
											assign node1559 = (inp[1]) ? node1561 : 4'b0000;
												assign node1561 = (inp[15]) ? 4'b0000 : node1562;
													assign node1562 = (inp[6]) ? 4'b0010 : node1563;
														assign node1563 = (inp[8]) ? 4'b0000 : node1564;
															assign node1564 = (inp[10]) ? 4'b0000 : 4'b0010;
											assign node1570 = (inp[15]) ? node1572 : 4'b0010;
												assign node1572 = (inp[10]) ? node1574 : 4'b0010;
													assign node1574 = (inp[8]) ? node1576 : 4'b0010;
														assign node1576 = (inp[6]) ? 4'b0010 : node1577;
															assign node1577 = (inp[1]) ? 4'b0010 : 4'b0000;
										assign node1581 = (inp[13]) ? 4'b0000 : node1582;
											assign node1582 = (inp[1]) ? node1590 : node1583;
												assign node1583 = (inp[15]) ? 4'b0010 : node1584;
													assign node1584 = (inp[8]) ? node1586 : 4'b0000;
														assign node1586 = (inp[6]) ? 4'b0000 : 4'b0010;
												assign node1590 = (inp[15]) ? node1592 : 4'b0000;
													assign node1592 = (inp[8]) ? node1594 : 4'b0000;
														assign node1594 = (inp[6]) ? 4'b0000 : 4'b0010;
									assign node1598 = (inp[11]) ? node1620 : node1599;
										assign node1599 = (inp[13]) ? node1601 : 4'b0000;
											assign node1601 = (inp[1]) ? node1611 : node1602;
												assign node1602 = (inp[15]) ? 4'b0000 : node1603;
													assign node1603 = (inp[10]) ? node1605 : 4'b0000;
														assign node1605 = (inp[8]) ? 4'b0000 : node1606;
															assign node1606 = (inp[6]) ? 4'b0010 : 4'b0000;
												assign node1611 = (inp[15]) ? node1613 : 4'b0010;
													assign node1613 = (inp[6]) ? 4'b0010 : node1614;
														assign node1614 = (inp[10]) ? 4'b0000 : node1615;
															assign node1615 = (inp[8]) ? 4'b0000 : 4'b0010;
										assign node1620 = (inp[13]) ? node1622 : 4'b0010;
											assign node1622 = (inp[15]) ? node1630 : node1623;
												assign node1623 = (inp[8]) ? node1625 : 4'b0000;
													assign node1625 = (inp[1]) ? 4'b0000 : node1626;
														assign node1626 = (inp[6]) ? 4'b0000 : 4'b0010;
												assign node1630 = (inp[1]) ? node1632 : 4'b0010;
													assign node1632 = (inp[8]) ? node1634 : 4'b0000;
														assign node1634 = (inp[6]) ? 4'b0000 : 4'b0010;
						assign node1637 = (inp[3]) ? node1705 : node1638;
							assign node1638 = (inp[11]) ? node1640 : 4'b0010;
								assign node1640 = (inp[5]) ? node1674 : node1641;
									assign node1641 = (inp[9]) ? 4'b0010 : node1642;
										assign node1642 = (inp[13]) ? node1656 : node1643;
											assign node1643 = (inp[15]) ? 4'b0000 : node1644;
												assign node1644 = (inp[8]) ? node1650 : node1645;
													assign node1645 = (inp[10]) ? node1647 : 4'b0010;
														assign node1647 = (inp[6]) ? 4'b0010 : 4'b0000;
													assign node1650 = (inp[1]) ? node1652 : 4'b0000;
														assign node1652 = (inp[10]) ? 4'b0000 : 4'b0010;
											assign node1656 = (inp[15]) ? node1658 : 4'b0010;
												assign node1658 = (inp[1]) ? node1666 : node1659;
													assign node1659 = (inp[8]) ? 4'b0000 : node1660;
														assign node1660 = (inp[10]) ? node1662 : 4'b0010;
															assign node1662 = (inp[6]) ? 4'b0010 : 4'b0000;
													assign node1666 = (inp[8]) ? node1668 : 4'b0010;
														assign node1668 = (inp[10]) ? node1670 : 4'b0010;
															assign node1670 = (inp[6]) ? 4'b0010 : 4'b0000;
									assign node1674 = (inp[9]) ? node1676 : 4'b0000;
										assign node1676 = (inp[13]) ? node1692 : node1677;
											assign node1677 = (inp[15]) ? 4'b0000 : node1678;
												assign node1678 = (inp[10]) ? node1684 : node1679;
													assign node1679 = (inp[8]) ? node1681 : 4'b0010;
														assign node1681 = (inp[1]) ? 4'b0010 : 4'b0000;
													assign node1684 = (inp[6]) ? node1686 : 4'b0000;
														assign node1686 = (inp[1]) ? 4'b0010 : node1687;
															assign node1687 = (inp[8]) ? 4'b0000 : 4'b0010;
											assign node1692 = (inp[15]) ? node1694 : 4'b0010;
												assign node1694 = (inp[1]) ? node1700 : node1695;
													assign node1695 = (inp[8]) ? 4'b0000 : node1696;
														assign node1696 = (inp[6]) ? 4'b0010 : 4'b0000;
													assign node1700 = (inp[6]) ? 4'b0010 : node1701;
														assign node1701 = (inp[10]) ? 4'b0000 : 4'b0010;
							assign node1705 = (inp[13]) ? node1849 : node1706;
								assign node1706 = (inp[11]) ? node1768 : node1707;
									assign node1707 = (inp[1]) ? node1741 : node1708;
										assign node1708 = (inp[5]) ? node1726 : node1709;
											assign node1709 = (inp[9]) ? node1715 : node1710;
												assign node1710 = (inp[6]) ? 4'b1000 : node1711;
													assign node1711 = (inp[15]) ? 4'b0010 : 4'b1000;
												assign node1715 = (inp[6]) ? node1723 : node1716;
													assign node1716 = (inp[15]) ? 4'b0000 : node1717;
														assign node1717 = (inp[10]) ? 4'b0000 : node1718;
															assign node1718 = (inp[8]) ? 4'b0000 : 4'b0010;
													assign node1723 = (inp[15]) ? 4'b0010 : 4'b0000;
											assign node1726 = (inp[9]) ? node1728 : 4'b0010;
												assign node1728 = (inp[6]) ? node1736 : node1729;
													assign node1729 = (inp[15]) ? node1731 : 4'b1010;
														assign node1731 = (inp[10]) ? node1733 : 4'b1010;
															assign node1733 = (inp[8]) ? 4'b1000 : 4'b1010;
													assign node1736 = (inp[15]) ? 4'b0000 : node1737;
														assign node1737 = (inp[8]) ? 4'b0000 : 4'b0010;
										assign node1741 = (inp[6]) ? node1761 : node1742;
											assign node1742 = (inp[15]) ? node1752 : node1743;
												assign node1743 = (inp[9]) ? node1745 : 4'b1000;
													assign node1745 = (inp[5]) ? node1747 : 4'b1000;
														assign node1747 = (inp[8]) ? 4'b0000 : node1748;
															assign node1748 = (inp[10]) ? 4'b0000 : 4'b0010;
												assign node1752 = (inp[5]) ? node1756 : node1753;
													assign node1753 = (inp[9]) ? 4'b0010 : 4'b1000;
													assign node1756 = (inp[8]) ? 4'b0010 : node1757;
														assign node1757 = (inp[9]) ? 4'b0000 : 4'b0010;
											assign node1761 = (inp[15]) ? 4'b1000 : node1762;
												assign node1762 = (inp[5]) ? node1764 : 4'b1010;
													assign node1764 = (inp[9]) ? 4'b1010 : 4'b1000;
									assign node1768 = (inp[9]) ? node1790 : node1769;
										assign node1769 = (inp[5]) ? node1779 : node1770;
											assign node1770 = (inp[15]) ? node1772 : 4'b0010;
												assign node1772 = (inp[1]) ? 4'b0010 : node1773;
													assign node1773 = (inp[6]) ? node1775 : 4'b0000;
														assign node1775 = (inp[8]) ? 4'b0000 : 4'b0010;
											assign node1779 = (inp[1]) ? node1781 : 4'b0000;
												assign node1781 = (inp[15]) ? 4'b0000 : node1782;
													assign node1782 = (inp[6]) ? 4'b0010 : node1783;
														assign node1783 = (inp[10]) ? 4'b0000 : node1784;
															assign node1784 = (inp[8]) ? 4'b0000 : 4'b0010;
										assign node1790 = (inp[1]) ? node1832 : node1791;
											assign node1791 = (inp[10]) ? node1809 : node1792;
												assign node1792 = (inp[6]) ? node1804 : node1793;
													assign node1793 = (inp[5]) ? node1799 : node1794;
														assign node1794 = (inp[15]) ? node1796 : 4'b1000;
															assign node1796 = (inp[2]) ? 4'b1010 : 4'b1000;
														assign node1799 = (inp[15]) ? node1801 : 4'b1010;
															assign node1801 = (inp[8]) ? 4'b1000 : 4'b1010;
													assign node1804 = (inp[5]) ? node1806 : 4'b1010;
														assign node1806 = (inp[15]) ? 4'b1010 : 4'b1000;
												assign node1809 = (inp[6]) ? node1823 : node1810;
													assign node1810 = (inp[2]) ? node1812 : 4'b1000;
														assign node1812 = (inp[8]) ? node1818 : node1813;
															assign node1813 = (inp[5]) ? node1815 : 4'b1000;
																assign node1815 = (inp[15]) ? 4'b1000 : 4'b1010;
															assign node1818 = (inp[5]) ? 4'b1000 : node1819;
																assign node1819 = (inp[15]) ? 4'b1010 : 4'b1000;
													assign node1823 = (inp[5]) ? node1829 : node1824;
														assign node1824 = (inp[15]) ? node1826 : 4'b1010;
															assign node1826 = (inp[8]) ? 4'b1000 : 4'b1010;
														assign node1829 = (inp[15]) ? 4'b1010 : 4'b1000;
											assign node1832 = (inp[15]) ? node1844 : node1833;
												assign node1833 = (inp[5]) ? node1841 : node1834;
													assign node1834 = (inp[10]) ? node1836 : 4'b0010;
														assign node1836 = (inp[8]) ? node1838 : 4'b0010;
															assign node1838 = (inp[6]) ? 4'b0010 : 4'b0000;
													assign node1841 = (inp[6]) ? 4'b0010 : 4'b1010;
												assign node1844 = (inp[5]) ? node1846 : 4'b0000;
													assign node1846 = (inp[6]) ? 4'b0000 : 4'b1000;
								assign node1849 = (inp[9]) ? node1963 : node1850;
									assign node1850 = (inp[11]) ? node1934 : node1851;
										assign node1851 = (inp[5]) ? node1889 : node1852;
											assign node1852 = (inp[15]) ? node1884 : node1853;
												assign node1853 = (inp[10]) ? node1863 : node1854;
													assign node1854 = (inp[1]) ? node1858 : node1855;
														assign node1855 = (inp[6]) ? 4'b1000 : 4'b1010;
														assign node1858 = (inp[8]) ? node1860 : 4'b1010;
															assign node1860 = (inp[6]) ? 4'b1010 : 4'b1000;
													assign node1863 = (inp[2]) ? node1871 : node1864;
														assign node1864 = (inp[1]) ? node1868 : node1865;
															assign node1865 = (inp[6]) ? 4'b1000 : 4'b1010;
															assign node1868 = (inp[6]) ? 4'b1010 : 4'b1000;
														assign node1871 = (inp[8]) ? node1877 : node1872;
															assign node1872 = (inp[6]) ? 4'b1010 : node1873;
																assign node1873 = (inp[1]) ? 4'b1000 : 4'b1010;
															assign node1877 = (inp[1]) ? node1881 : node1878;
																assign node1878 = (inp[6]) ? 4'b1000 : 4'b1010;
																assign node1881 = (inp[6]) ? 4'b1010 : 4'b1000;
												assign node1884 = (inp[1]) ? node1886 : 4'b1010;
													assign node1886 = (inp[6]) ? 4'b1010 : 4'b1000;
											assign node1889 = (inp[10]) ? node1919 : node1890;
												assign node1890 = (inp[2]) ? node1906 : node1891;
													assign node1891 = (inp[8]) ? node1901 : node1892;
														assign node1892 = (inp[6]) ? node1898 : node1893;
															assign node1893 = (inp[15]) ? node1895 : 4'b1000;
																assign node1895 = (inp[1]) ? 4'b1010 : 4'b1000;
															assign node1898 = (inp[1]) ? 4'b1000 : 4'b1010;
														assign node1901 = (inp[1]) ? node1903 : 4'b1000;
															assign node1903 = (inp[6]) ? 4'b1000 : 4'b1010;
													assign node1906 = (inp[8]) ? node1912 : node1907;
														assign node1907 = (inp[1]) ? node1909 : 4'b1010;
															assign node1909 = (inp[6]) ? 4'b1000 : 4'b1010;
														assign node1912 = (inp[1]) ? 4'b1010 : node1913;
															assign node1913 = (inp[15]) ? 4'b1000 : node1914;
																assign node1914 = (inp[6]) ? 4'b1010 : 4'b1000;
												assign node1919 = (inp[6]) ? node1927 : node1920;
													assign node1920 = (inp[1]) ? node1922 : 4'b1000;
														assign node1922 = (inp[15]) ? 4'b1010 : node1923;
															assign node1923 = (inp[8]) ? 4'b1010 : 4'b1000;
													assign node1927 = (inp[1]) ? 4'b1000 : node1928;
														assign node1928 = (inp[8]) ? node1930 : 4'b1010;
															assign node1930 = (inp[2]) ? 4'b1010 : 4'b1000;
										assign node1934 = (inp[5]) ? node1950 : node1935;
											assign node1935 = (inp[1]) ? node1941 : node1936;
												assign node1936 = (inp[6]) ? 4'b1000 : node1937;
													assign node1937 = (inp[15]) ? 4'b0010 : 4'b1000;
												assign node1941 = (inp[6]) ? 4'b1010 : node1942;
													assign node1942 = (inp[15]) ? 4'b1000 : node1943;
														assign node1943 = (inp[8]) ? node1945 : 4'b1010;
															assign node1945 = (inp[10]) ? 4'b1000 : 4'b1010;
											assign node1950 = (inp[1]) ? node1958 : node1951;
												assign node1951 = (inp[8]) ? node1953 : 4'b0010;
													assign node1953 = (inp[10]) ? node1955 : 4'b0010;
														assign node1955 = (inp[6]) ? 4'b0010 : 4'b0000;
												assign node1958 = (inp[6]) ? 4'b1000 : node1959;
													assign node1959 = (inp[15]) ? 4'b0010 : 4'b1000;
									assign node1963 = (inp[1]) ? node2019 : node1964;
										assign node1964 = (inp[5]) ? node1990 : node1965;
											assign node1965 = (inp[6]) ? node1987 : node1966;
												assign node1966 = (inp[11]) ? node1978 : node1967;
													assign node1967 = (inp[15]) ? node1973 : node1968;
														assign node1968 = (inp[8]) ? 4'b1001 : node1969;
															assign node1969 = (inp[10]) ? 4'b1001 : 4'b1011;
														assign node1973 = (inp[8]) ? node1975 : 4'b0011;
															assign node1975 = (inp[10]) ? 4'b0001 : 4'b0011;
													assign node1978 = (inp[8]) ? node1982 : node1979;
														assign node1979 = (inp[15]) ? 4'b1000 : 4'b1010;
														assign node1982 = (inp[15]) ? 4'b1010 : node1983;
															assign node1983 = (inp[10]) ? 4'b1000 : 4'b1010;
												assign node1987 = (inp[8]) ? 4'b1001 : 4'b1011;
											assign node1990 = (inp[11]) ? node2004 : node1991;
												assign node1991 = (inp[8]) ? node1999 : node1992;
													assign node1992 = (inp[6]) ? 4'b0011 : node1993;
														assign node1993 = (inp[15]) ? node1995 : 4'b0001;
															assign node1995 = (inp[10]) ? 4'b0001 : 4'b0011;
													assign node1999 = (inp[15]) ? 4'b0001 : node2000;
														assign node2000 = (inp[6]) ? 4'b0001 : 4'b0011;
												assign node2004 = (inp[6]) ? node2016 : node2005;
													assign node2005 = (inp[15]) ? node2011 : node2006;
														assign node2006 = (inp[10]) ? 4'b1000 : node2007;
															assign node2007 = (inp[8]) ? 4'b1000 : 4'b1010;
														assign node2011 = (inp[8]) ? node2013 : 4'b0010;
															assign node2013 = (inp[10]) ? 4'b0000 : 4'b0010;
													assign node2016 = (inp[8]) ? 4'b0001 : 4'b0011;
										assign node2019 = (inp[6]) ? 4'b0000 : node2020;
											assign node2020 = (inp[10]) ? node2028 : node2021;
												assign node2021 = (inp[11]) ? node2025 : node2022;
													assign node2022 = (inp[15]) ? 4'b0011 : 4'b1011;
													assign node2025 = (inp[15]) ? 4'b0010 : 4'b1010;
												assign node2028 = (inp[15]) ? node2032 : node2029;
													assign node2029 = (inp[11]) ? 4'b1000 : 4'b1001;
													assign node2032 = (inp[11]) ? 4'b0000 : 4'b0001;
					assign node2036 = (inp[3]) ? node2038 : 4'b0000;
						assign node2038 = (inp[11]) ? node2248 : node2039;
							assign node2039 = (inp[9]) ? node2131 : node2040;
								assign node2040 = (inp[7]) ? node2078 : node2041;
									assign node2041 = (inp[5]) ? 4'b0000 : node2042;
										assign node2042 = (inp[13]) ? node2060 : node2043;
											assign node2043 = (inp[15]) ? 4'b0000 : node2044;
												assign node2044 = (inp[1]) ? node2052 : node2045;
													assign node2045 = (inp[8]) ? 4'b0000 : node2046;
														assign node2046 = (inp[6]) ? 4'b0010 : node2047;
															assign node2047 = (inp[10]) ? 4'b0000 : 4'b0010;
													assign node2052 = (inp[10]) ? node2054 : 4'b0010;
														assign node2054 = (inp[8]) ? node2056 : 4'b0010;
															assign node2056 = (inp[6]) ? 4'b0010 : 4'b0000;
											assign node2060 = (inp[15]) ? node2062 : 4'b0010;
												assign node2062 = (inp[8]) ? node2070 : node2063;
													assign node2063 = (inp[6]) ? 4'b0010 : node2064;
														assign node2064 = (inp[10]) ? node2066 : 4'b0010;
															assign node2066 = (inp[1]) ? 4'b0010 : 4'b0000;
													assign node2070 = (inp[1]) ? node2072 : 4'b0000;
														assign node2072 = (inp[6]) ? 4'b0010 : node2073;
															assign node2073 = (inp[10]) ? 4'b0000 : 4'b0010;
									assign node2078 = (inp[13]) ? node2096 : node2079;
										assign node2079 = (inp[5]) ? 4'b0010 : node2080;
											assign node2080 = (inp[1]) ? node2088 : node2081;
												assign node2081 = (inp[15]) ? 4'b0010 : node2082;
													assign node2082 = (inp[8]) ? node2084 : 4'b0000;
														assign node2084 = (inp[6]) ? 4'b0000 : 4'b0010;
												assign node2088 = (inp[6]) ? 4'b0000 : node2089;
													assign node2089 = (inp[15]) ? node2091 : 4'b0000;
														assign node2091 = (inp[8]) ? 4'b0010 : 4'b0000;
										assign node2096 = (inp[6]) ? node2118 : node2097;
											assign node2097 = (inp[5]) ? node2107 : node2098;
												assign node2098 = (inp[1]) ? node2100 : 4'b0000;
													assign node2100 = (inp[15]) ? node2102 : 4'b0010;
														assign node2102 = (inp[8]) ? 4'b0000 : node2103;
															assign node2103 = (inp[10]) ? 4'b0000 : 4'b0010;
												assign node2107 = (inp[15]) ? node2113 : node2108;
													assign node2108 = (inp[1]) ? 4'b0000 : node2109;
														assign node2109 = (inp[8]) ? 4'b0010 : 4'b0000;
													assign node2113 = (inp[8]) ? 4'b0010 : node2114;
														assign node2114 = (inp[1]) ? 4'b0000 : 4'b0010;
											assign node2118 = (inp[5]) ? node2126 : node2119;
												assign node2119 = (inp[1]) ? 4'b0010 : node2120;
													assign node2120 = (inp[8]) ? 4'b0000 : node2121;
														assign node2121 = (inp[15]) ? 4'b0000 : 4'b0010;
												assign node2126 = (inp[1]) ? 4'b0000 : node2127;
													assign node2127 = (inp[15]) ? 4'b0010 : 4'b0000;
								assign node2131 = (inp[7]) ? node2169 : node2132;
									assign node2132 = (inp[5]) ? node2134 : 4'b0010;
										assign node2134 = (inp[15]) ? node2152 : node2135;
											assign node2135 = (inp[13]) ? 4'b0010 : node2136;
												assign node2136 = (inp[1]) ? node2144 : node2137;
													assign node2137 = (inp[8]) ? 4'b0000 : node2138;
														assign node2138 = (inp[6]) ? 4'b0010 : node2139;
															assign node2139 = (inp[10]) ? 4'b0000 : 4'b0010;
													assign node2144 = (inp[6]) ? 4'b0010 : node2145;
														assign node2145 = (inp[10]) ? node2147 : 4'b0010;
															assign node2147 = (inp[8]) ? 4'b0000 : 4'b0010;
											assign node2152 = (inp[13]) ? node2154 : 4'b0000;
												assign node2154 = (inp[8]) ? node2162 : node2155;
													assign node2155 = (inp[2]) ? 4'b0010 : node2156;
														assign node2156 = (inp[6]) ? 4'b0010 : node2157;
															assign node2157 = (inp[10]) ? 4'b0000 : 4'b0010;
													assign node2162 = (inp[1]) ? node2164 : 4'b0000;
														assign node2164 = (inp[10]) ? node2166 : 4'b0010;
															assign node2166 = (inp[6]) ? 4'b0010 : 4'b0000;
									assign node2169 = (inp[13]) ? node2211 : node2170;
										assign node2170 = (inp[1]) ? node2194 : node2171;
											assign node2171 = (inp[5]) ? node2181 : node2172;
												assign node2172 = (inp[6]) ? node2176 : node2173;
													assign node2173 = (inp[15]) ? 4'b0010 : 4'b1000;
													assign node2176 = (inp[15]) ? 4'b1000 : node2177;
														assign node2177 = (inp[8]) ? 4'b1000 : 4'b1010;
												assign node2181 = (inp[15]) ? node2189 : node2182;
													assign node2182 = (inp[10]) ? node2184 : 4'b0010;
														assign node2184 = (inp[8]) ? node2186 : 4'b0010;
															assign node2186 = (inp[6]) ? 4'b0010 : 4'b0000;
													assign node2189 = (inp[8]) ? 4'b0000 : node2190;
														assign node2190 = (inp[6]) ? 4'b0010 : 4'b0000;
											assign node2194 = (inp[15]) ? node2202 : node2195;
												assign node2195 = (inp[6]) ? 4'b1010 : node2196;
													assign node2196 = (inp[8]) ? node2198 : 4'b1000;
														assign node2198 = (inp[5]) ? 4'b1000 : 4'b1010;
												assign node2202 = (inp[6]) ? 4'b1000 : node2203;
													assign node2203 = (inp[5]) ? 4'b0010 : node2204;
														assign node2204 = (inp[8]) ? node2206 : 4'b1010;
															assign node2206 = (inp[10]) ? 4'b1000 : 4'b1010;
										assign node2211 = (inp[1]) ? node2239 : node2212;
											assign node2212 = (inp[8]) ? node2226 : node2213;
												assign node2213 = (inp[6]) ? node2223 : node2214;
													assign node2214 = (inp[5]) ? node2220 : node2215;
														assign node2215 = (inp[10]) ? 4'b0000 : node2216;
															assign node2216 = (inp[15]) ? 4'b0010 : 4'b0000;
														assign node2220 = (inp[15]) ? 4'b1000 : 4'b1010;
													assign node2223 = (inp[5]) ? 4'b0010 : 4'b1010;
												assign node2226 = (inp[6]) ? node2236 : node2227;
													assign node2227 = (inp[5]) ? node2231 : node2228;
														assign node2228 = (inp[15]) ? 4'b0000 : 4'b0010;
														assign node2231 = (inp[15]) ? 4'b1010 : node2232;
															assign node2232 = (inp[10]) ? 4'b1000 : 4'b1010;
													assign node2236 = (inp[5]) ? 4'b0000 : 4'b1000;
											assign node2239 = (inp[6]) ? 4'b0000 : node2240;
												assign node2240 = (inp[15]) ? node2244 : node2241;
													assign node2241 = (inp[10]) ? 4'b1001 : 4'b1011;
													assign node2244 = (inp[10]) ? 4'b0001 : 4'b0011;
							assign node2248 = (inp[7]) ? node2250 : 4'b0000;
								assign node2250 = (inp[5]) ? node2334 : node2251;
									assign node2251 = (inp[13]) ? node2289 : node2252;
										assign node2252 = (inp[9]) ? node2268 : node2253;
											assign node2253 = (inp[15]) ? 4'b0000 : node2254;
												assign node2254 = (inp[1]) ? node2262 : node2255;
													assign node2255 = (inp[8]) ? 4'b0000 : node2256;
														assign node2256 = (inp[10]) ? node2258 : 4'b0010;
															assign node2258 = (inp[6]) ? 4'b0010 : 4'b0000;
													assign node2262 = (inp[10]) ? node2264 : 4'b0010;
														assign node2264 = (inp[6]) ? 4'b0010 : 4'b0000;
											assign node2268 = (inp[15]) ? node2282 : node2269;
												assign node2269 = (inp[1]) ? node2275 : node2270;
													assign node2270 = (inp[8]) ? node2272 : 4'b0000;
														assign node2272 = (inp[6]) ? 4'b0000 : 4'b0010;
													assign node2275 = (inp[6]) ? 4'b0010 : node2276;
														assign node2276 = (inp[10]) ? 4'b0000 : node2277;
															assign node2277 = (inp[8]) ? 4'b0000 : 4'b0010;
												assign node2282 = (inp[1]) ? node2284 : 4'b0010;
													assign node2284 = (inp[6]) ? 4'b0000 : node2285;
														assign node2285 = (inp[8]) ? 4'b0010 : 4'b0000;
										assign node2289 = (inp[9]) ? node2307 : node2290;
											assign node2290 = (inp[15]) ? node2292 : 4'b0010;
												assign node2292 = (inp[1]) ? node2300 : node2293;
													assign node2293 = (inp[8]) ? 4'b0000 : node2294;
														assign node2294 = (inp[10]) ? node2296 : 4'b0010;
															assign node2296 = (inp[6]) ? 4'b0010 : 4'b0000;
													assign node2300 = (inp[8]) ? node2302 : 4'b0010;
														assign node2302 = (inp[10]) ? node2304 : 4'b0010;
															assign node2304 = (inp[6]) ? 4'b0010 : 4'b0000;
											assign node2307 = (inp[15]) ? node2321 : node2308;
												assign node2308 = (inp[1]) ? node2316 : node2309;
													assign node2309 = (inp[8]) ? 4'b1000 : node2310;
														assign node2310 = (inp[10]) ? node2312 : 4'b1010;
															assign node2312 = (inp[6]) ? 4'b1010 : 4'b1000;
													assign node2316 = (inp[6]) ? 4'b0000 : node2317;
														assign node2317 = (inp[10]) ? 4'b1000 : 4'b1010;
												assign node2321 = (inp[6]) ? node2329 : node2322;
													assign node2322 = (inp[10]) ? node2324 : 4'b0010;
														assign node2324 = (inp[8]) ? 4'b0000 : node2325;
															assign node2325 = (inp[1]) ? 4'b0000 : 4'b0010;
													assign node2329 = (inp[1]) ? 4'b0000 : node2330;
														assign node2330 = (inp[8]) ? 4'b1000 : 4'b1010;
									assign node2334 = (inp[9]) ? node2336 : 4'b0000;
										assign node2336 = (inp[15]) ? node2372 : node2337;
											assign node2337 = (inp[13]) ? node2353 : node2338;
												assign node2338 = (inp[1]) ? node2346 : node2339;
													assign node2339 = (inp[8]) ? 4'b0000 : node2340;
														assign node2340 = (inp[6]) ? 4'b0010 : node2341;
															assign node2341 = (inp[10]) ? 4'b0000 : 4'b0010;
													assign node2346 = (inp[6]) ? 4'b0010 : node2347;
														assign node2347 = (inp[10]) ? node2349 : 4'b0010;
															assign node2349 = (inp[8]) ? 4'b0000 : 4'b0010;
												assign node2353 = (inp[1]) ? node2367 : node2354;
													assign node2354 = (inp[10]) ? node2362 : node2355;
														assign node2355 = (inp[8]) ? node2359 : node2356;
															assign node2356 = (inp[6]) ? 4'b0010 : 4'b0000;
															assign node2359 = (inp[6]) ? 4'b0000 : 4'b0010;
														assign node2362 = (inp[8]) ? node2364 : 4'b0000;
															assign node2364 = (inp[6]) ? 4'b0000 : 4'b0010;
													assign node2367 = (inp[6]) ? 4'b0000 : node2368;
														assign node2368 = (inp[10]) ? 4'b1000 : 4'b1010;
											assign node2372 = (inp[13]) ? node2374 : 4'b0000;
												assign node2374 = (inp[10]) ? node2386 : node2375;
													assign node2375 = (inp[6]) ? node2381 : node2376;
														assign node2376 = (inp[1]) ? 4'b0010 : node2377;
															assign node2377 = (inp[8]) ? 4'b0000 : 4'b0010;
														assign node2381 = (inp[1]) ? 4'b0000 : node2382;
															assign node2382 = (inp[8]) ? 4'b0000 : 4'b0010;
													assign node2386 = (inp[6]) ? node2388 : 4'b0000;
														assign node2388 = (inp[1]) ? 4'b0000 : node2389;
															assign node2389 = (inp[8]) ? 4'b0000 : 4'b0010;

endmodule