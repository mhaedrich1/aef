module dtc_split125_bm56 (
	input  wire [12-1:0] inp,
	output wire [3-1:0] outp
);

	wire [3-1:0] node1;
	wire [3-1:0] node2;
	wire [3-1:0] node3;
	wire [3-1:0] node4;
	wire [3-1:0] node5;
	wire [3-1:0] node6;
	wire [3-1:0] node8;
	wire [3-1:0] node9;
	wire [3-1:0] node13;
	wire [3-1:0] node14;
	wire [3-1:0] node15;
	wire [3-1:0] node19;
	wire [3-1:0] node20;
	wire [3-1:0] node22;
	wire [3-1:0] node26;
	wire [3-1:0] node27;
	wire [3-1:0] node28;
	wire [3-1:0] node31;
	wire [3-1:0] node32;
	wire [3-1:0] node34;
	wire [3-1:0] node35;
	wire [3-1:0] node40;
	wire [3-1:0] node41;
	wire [3-1:0] node43;
	wire [3-1:0] node46;
	wire [3-1:0] node49;
	wire [3-1:0] node50;
	wire [3-1:0] node51;
	wire [3-1:0] node52;
	wire [3-1:0] node55;
	wire [3-1:0] node56;
	wire [3-1:0] node59;
	wire [3-1:0] node62;
	wire [3-1:0] node64;
	wire [3-1:0] node66;
	wire [3-1:0] node67;
	wire [3-1:0] node71;
	wire [3-1:0] node72;
	wire [3-1:0] node73;
	wire [3-1:0] node74;
	wire [3-1:0] node76;
	wire [3-1:0] node79;
	wire [3-1:0] node82;
	wire [3-1:0] node83;
	wire [3-1:0] node84;
	wire [3-1:0] node85;
	wire [3-1:0] node90;
	wire [3-1:0] node93;
	wire [3-1:0] node94;
	wire [3-1:0] node97;
	wire [3-1:0] node98;
	wire [3-1:0] node102;
	wire [3-1:0] node103;
	wire [3-1:0] node104;
	wire [3-1:0] node105;
	wire [3-1:0] node106;
	wire [3-1:0] node107;
	wire [3-1:0] node110;
	wire [3-1:0] node113;
	wire [3-1:0] node115;
	wire [3-1:0] node118;
	wire [3-1:0] node119;
	wire [3-1:0] node120;
	wire [3-1:0] node124;
	wire [3-1:0] node126;
	wire [3-1:0] node129;
	wire [3-1:0] node130;
	wire [3-1:0] node132;
	wire [3-1:0] node133;
	wire [3-1:0] node136;
	wire [3-1:0] node137;
	wire [3-1:0] node139;
	wire [3-1:0] node143;
	wire [3-1:0] node144;
	wire [3-1:0] node147;
	wire [3-1:0] node148;
	wire [3-1:0] node151;
	wire [3-1:0] node153;
	wire [3-1:0] node156;
	wire [3-1:0] node157;
	wire [3-1:0] node158;
	wire [3-1:0] node159;
	wire [3-1:0] node160;
	wire [3-1:0] node163;
	wire [3-1:0] node165;
	wire [3-1:0] node166;
	wire [3-1:0] node171;
	wire [3-1:0] node172;
	wire [3-1:0] node176;
	wire [3-1:0] node177;
	wire [3-1:0] node178;
	wire [3-1:0] node179;
	wire [3-1:0] node181;
	wire [3-1:0] node185;
	wire [3-1:0] node187;
	wire [3-1:0] node190;
	wire [3-1:0] node191;
	wire [3-1:0] node192;
	wire [3-1:0] node193;
	wire [3-1:0] node194;
	wire [3-1:0] node199;
	wire [3-1:0] node200;
	wire [3-1:0] node204;
	wire [3-1:0] node207;
	wire [3-1:0] node208;
	wire [3-1:0] node209;
	wire [3-1:0] node210;
	wire [3-1:0] node211;
	wire [3-1:0] node212;
	wire [3-1:0] node213;
	wire [3-1:0] node214;
	wire [3-1:0] node220;
	wire [3-1:0] node221;
	wire [3-1:0] node223;
	wire [3-1:0] node227;
	wire [3-1:0] node228;
	wire [3-1:0] node230;
	wire [3-1:0] node232;
	wire [3-1:0] node235;
	wire [3-1:0] node236;
	wire [3-1:0] node238;
	wire [3-1:0] node239;
	wire [3-1:0] node243;
	wire [3-1:0] node245;
	wire [3-1:0] node246;
	wire [3-1:0] node249;
	wire [3-1:0] node252;
	wire [3-1:0] node253;
	wire [3-1:0] node254;
	wire [3-1:0] node255;
	wire [3-1:0] node256;
	wire [3-1:0] node257;
	wire [3-1:0] node260;
	wire [3-1:0] node263;
	wire [3-1:0] node265;
	wire [3-1:0] node268;
	wire [3-1:0] node269;
	wire [3-1:0] node272;
	wire [3-1:0] node275;
	wire [3-1:0] node276;
	wire [3-1:0] node279;
	wire [3-1:0] node280;
	wire [3-1:0] node282;
	wire [3-1:0] node286;
	wire [3-1:0] node287;
	wire [3-1:0] node289;
	wire [3-1:0] node290;
	wire [3-1:0] node294;
	wire [3-1:0] node295;
	wire [3-1:0] node296;
	wire [3-1:0] node298;
	wire [3-1:0] node301;
	wire [3-1:0] node304;
	wire [3-1:0] node307;
	wire [3-1:0] node308;
	wire [3-1:0] node309;
	wire [3-1:0] node310;
	wire [3-1:0] node311;
	wire [3-1:0] node312;
	wire [3-1:0] node315;
	wire [3-1:0] node318;
	wire [3-1:0] node320;
	wire [3-1:0] node323;
	wire [3-1:0] node324;
	wire [3-1:0] node326;
	wire [3-1:0] node329;
	wire [3-1:0] node332;
	wire [3-1:0] node333;
	wire [3-1:0] node334;
	wire [3-1:0] node337;
	wire [3-1:0] node340;
	wire [3-1:0] node341;
	wire [3-1:0] node343;
	wire [3-1:0] node346;
	wire [3-1:0] node348;
	wire [3-1:0] node351;
	wire [3-1:0] node352;
	wire [3-1:0] node353;
	wire [3-1:0] node354;
	wire [3-1:0] node355;
	wire [3-1:0] node358;
	wire [3-1:0] node361;
	wire [3-1:0] node365;
	wire [3-1:0] node366;
	wire [3-1:0] node367;
	wire [3-1:0] node369;
	wire [3-1:0] node373;
	wire [3-1:0] node374;
	wire [3-1:0] node377;
	wire [3-1:0] node379;
	wire [3-1:0] node381;
	wire [3-1:0] node384;
	wire [3-1:0] node385;
	wire [3-1:0] node386;
	wire [3-1:0] node387;
	wire [3-1:0] node388;
	wire [3-1:0] node389;
	wire [3-1:0] node390;
	wire [3-1:0] node392;
	wire [3-1:0] node393;
	wire [3-1:0] node398;
	wire [3-1:0] node399;
	wire [3-1:0] node400;
	wire [3-1:0] node405;
	wire [3-1:0] node406;
	wire [3-1:0] node407;
	wire [3-1:0] node409;
	wire [3-1:0] node412;
	wire [3-1:0] node414;
	wire [3-1:0] node417;
	wire [3-1:0] node419;
	wire [3-1:0] node421;
	wire [3-1:0] node422;
	wire [3-1:0] node425;
	wire [3-1:0] node426;
	wire [3-1:0] node430;
	wire [3-1:0] node431;
	wire [3-1:0] node432;
	wire [3-1:0] node433;
	wire [3-1:0] node434;
	wire [3-1:0] node436;
	wire [3-1:0] node440;
	wire [3-1:0] node443;
	wire [3-1:0] node445;
	wire [3-1:0] node446;
	wire [3-1:0] node447;
	wire [3-1:0] node452;
	wire [3-1:0] node453;
	wire [3-1:0] node454;
	wire [3-1:0] node455;
	wire [3-1:0] node457;
	wire [3-1:0] node461;
	wire [3-1:0] node463;
	wire [3-1:0] node464;
	wire [3-1:0] node468;
	wire [3-1:0] node469;
	wire [3-1:0] node471;
	wire [3-1:0] node473;
	wire [3-1:0] node476;
	wire [3-1:0] node479;
	wire [3-1:0] node480;
	wire [3-1:0] node481;
	wire [3-1:0] node482;
	wire [3-1:0] node483;
	wire [3-1:0] node485;
	wire [3-1:0] node488;
	wire [3-1:0] node489;
	wire [3-1:0] node491;
	wire [3-1:0] node494;
	wire [3-1:0] node497;
	wire [3-1:0] node498;
	wire [3-1:0] node499;
	wire [3-1:0] node503;
	wire [3-1:0] node506;
	wire [3-1:0] node507;
	wire [3-1:0] node508;
	wire [3-1:0] node509;
	wire [3-1:0] node513;
	wire [3-1:0] node514;
	wire [3-1:0] node517;
	wire [3-1:0] node520;
	wire [3-1:0] node521;
	wire [3-1:0] node523;
	wire [3-1:0] node526;
	wire [3-1:0] node527;
	wire [3-1:0] node530;
	wire [3-1:0] node533;
	wire [3-1:0] node534;
	wire [3-1:0] node535;
	wire [3-1:0] node536;
	wire [3-1:0] node540;
	wire [3-1:0] node543;
	wire [3-1:0] node544;
	wire [3-1:0] node546;
	wire [3-1:0] node547;
	wire [3-1:0] node551;
	wire [3-1:0] node552;
	wire [3-1:0] node556;
	wire [3-1:0] node557;
	wire [3-1:0] node558;
	wire [3-1:0] node559;
	wire [3-1:0] node560;
	wire [3-1:0] node561;
	wire [3-1:0] node563;
	wire [3-1:0] node567;
	wire [3-1:0] node568;
	wire [3-1:0] node572;
	wire [3-1:0] node573;
	wire [3-1:0] node575;
	wire [3-1:0] node577;
	wire [3-1:0] node578;
	wire [3-1:0] node582;
	wire [3-1:0] node583;
	wire [3-1:0] node584;
	wire [3-1:0] node588;
	wire [3-1:0] node589;
	wire [3-1:0] node592;
	wire [3-1:0] node594;
	wire [3-1:0] node597;
	wire [3-1:0] node598;
	wire [3-1:0] node599;
	wire [3-1:0] node600;
	wire [3-1:0] node601;
	wire [3-1:0] node603;
	wire [3-1:0] node607;
	wire [3-1:0] node608;
	wire [3-1:0] node610;
	wire [3-1:0] node613;
	wire [3-1:0] node616;
	wire [3-1:0] node617;
	wire [3-1:0] node619;
	wire [3-1:0] node622;
	wire [3-1:0] node625;
	wire [3-1:0] node626;
	wire [3-1:0] node627;
	wire [3-1:0] node628;
	wire [3-1:0] node629;
	wire [3-1:0] node634;
	wire [3-1:0] node637;
	wire [3-1:0] node638;
	wire [3-1:0] node640;
	wire [3-1:0] node643;
	wire [3-1:0] node645;
	wire [3-1:0] node648;
	wire [3-1:0] node649;
	wire [3-1:0] node650;
	wire [3-1:0] node651;
	wire [3-1:0] node654;
	wire [3-1:0] node655;
	wire [3-1:0] node658;
	wire [3-1:0] node661;
	wire [3-1:0] node662;
	wire [3-1:0] node665;
	wire [3-1:0] node666;
	wire [3-1:0] node667;
	wire [3-1:0] node671;
	wire [3-1:0] node672;
	wire [3-1:0] node675;
	wire [3-1:0] node678;
	wire [3-1:0] node679;
	wire [3-1:0] node680;
	wire [3-1:0] node681;
	wire [3-1:0] node682;
	wire [3-1:0] node687;
	wire [3-1:0] node688;
	wire [3-1:0] node691;
	wire [3-1:0] node692;
	wire [3-1:0] node696;
	wire [3-1:0] node697;
	wire [3-1:0] node698;
	wire [3-1:0] node701;
	wire [3-1:0] node704;
	wire [3-1:0] node705;
	wire [3-1:0] node706;
	wire [3-1:0] node709;

	assign outp = (inp[9]) ? node384 : node1;
		assign node1 = (inp[7]) ? node207 : node2;
			assign node2 = (inp[2]) ? node102 : node3;
				assign node3 = (inp[0]) ? node49 : node4;
					assign node4 = (inp[8]) ? node26 : node5;
						assign node5 = (inp[3]) ? node13 : node6;
							assign node6 = (inp[4]) ? node8 : 3'b011;
								assign node8 = (inp[10]) ? 3'b111 : node9;
									assign node9 = (inp[11]) ? 3'b001 : 3'b101;
							assign node13 = (inp[4]) ? node19 : node14;
								assign node14 = (inp[10]) ? 3'b101 : node15;
									assign node15 = (inp[1]) ? 3'b101 : 3'b111;
								assign node19 = (inp[5]) ? 3'b111 : node20;
									assign node20 = (inp[10]) ? node22 : 3'b001;
										assign node22 = (inp[1]) ? 3'b111 : 3'b001;
						assign node26 = (inp[3]) ? node40 : node27;
							assign node27 = (inp[6]) ? node31 : node28;
								assign node28 = (inp[11]) ? 3'b011 : 3'b001;
								assign node31 = (inp[10]) ? 3'b001 : node32;
									assign node32 = (inp[1]) ? node34 : 3'b001;
										assign node34 = (inp[11]) ? 3'b111 : node35;
											assign node35 = (inp[4]) ? 3'b101 : 3'b101;
							assign node40 = (inp[11]) ? node46 : node41;
								assign node41 = (inp[4]) ? node43 : 3'b011;
									assign node43 = (inp[6]) ? 3'b001 : 3'b011;
								assign node46 = (inp[5]) ? 3'b111 : 3'b011;
					assign node49 = (inp[8]) ? node71 : node50;
						assign node50 = (inp[3]) ? node62 : node51;
							assign node51 = (inp[1]) ? node55 : node52;
								assign node52 = (inp[4]) ? 3'b001 : 3'b101;
								assign node55 = (inp[5]) ? node59 : node56;
									assign node56 = (inp[4]) ? 3'b101 : 3'b011;
									assign node59 = (inp[4]) ? 3'b110 : 3'b101;
							assign node62 = (inp[4]) ? node64 : 3'b101;
								assign node64 = (inp[11]) ? node66 : 3'b010;
									assign node66 = (inp[1]) ? 3'b110 : node67;
										assign node67 = (inp[6]) ? 3'b010 : 3'b110;
						assign node71 = (inp[1]) ? node93 : node72;
							assign node72 = (inp[4]) ? node82 : node73;
								assign node73 = (inp[10]) ? node79 : node74;
									assign node74 = (inp[11]) ? node76 : 3'b001;
										assign node76 = (inp[6]) ? 3'b110 : 3'b001;
									assign node79 = (inp[5]) ? 3'b010 : 3'b110;
								assign node82 = (inp[3]) ? node90 : node83;
									assign node83 = (inp[5]) ? 3'b010 : node84;
										assign node84 = (inp[11]) ? 3'b010 : node85;
											assign node85 = (inp[10]) ? 3'b110 : 3'b010;
									assign node90 = (inp[10]) ? 3'b100 : 3'b010;
							assign node93 = (inp[6]) ? node97 : node94;
								assign node94 = (inp[10]) ? 3'b100 : 3'b000;
								assign node97 = (inp[10]) ? 3'b010 : node98;
									assign node98 = (inp[4]) ? 3'b100 : 3'b110;
				assign node102 = (inp[0]) ? node156 : node103;
					assign node103 = (inp[8]) ? node129 : node104;
						assign node104 = (inp[4]) ? node118 : node105;
							assign node105 = (inp[3]) ? node113 : node106;
								assign node106 = (inp[11]) ? node110 : node107;
									assign node107 = (inp[1]) ? 3'b011 : 3'b111;
									assign node110 = (inp[6]) ? 3'b001 : 3'b101;
								assign node113 = (inp[11]) ? node115 : 3'b101;
									assign node115 = (inp[10]) ? 3'b001 : 3'b101;
							assign node118 = (inp[5]) ? node124 : node119;
								assign node119 = (inp[1]) ? 3'b110 : node120;
									assign node120 = (inp[10]) ? 3'b101 : 3'b001;
								assign node124 = (inp[10]) ? node126 : 3'b110;
									assign node126 = (inp[6]) ? 3'b010 : 3'b110;
						assign node129 = (inp[4]) ? node143 : node130;
							assign node130 = (inp[10]) ? node132 : 3'b110;
								assign node132 = (inp[5]) ? node136 : node133;
									assign node133 = (inp[11]) ? 3'b110 : 3'b001;
									assign node136 = (inp[11]) ? 3'b010 : node137;
										assign node137 = (inp[3]) ? node139 : 3'b110;
											assign node139 = (inp[6]) ? 3'b010 : 3'b110;
							assign node143 = (inp[5]) ? node147 : node144;
								assign node144 = (inp[1]) ? 3'b100 : 3'b110;
								assign node147 = (inp[11]) ? node151 : node148;
									assign node148 = (inp[1]) ? 3'b100 : 3'b010;
									assign node151 = (inp[6]) ? node153 : 3'b000;
										assign node153 = (inp[10]) ? 3'b000 : 3'b100;
					assign node156 = (inp[6]) ? node176 : node157;
						assign node157 = (inp[10]) ? node171 : node158;
							assign node158 = (inp[5]) ? 3'b010 : node159;
								assign node159 = (inp[11]) ? node163 : node160;
									assign node160 = (inp[1]) ? 3'b010 : 3'b110;
									assign node163 = (inp[3]) ? node165 : 3'b000;
										assign node165 = (inp[4]) ? 3'b010 : node166;
											assign node166 = (inp[8]) ? 3'b000 : 3'b010;
							assign node171 = (inp[1]) ? 3'b110 : node172;
								assign node172 = (inp[11]) ? 3'b110 : 3'b000;
						assign node176 = (inp[11]) ? node190 : node177;
							assign node177 = (inp[3]) ? node185 : node178;
								assign node178 = (inp[5]) ? 3'b000 : node179;
									assign node179 = (inp[1]) ? node181 : 3'b010;
										assign node181 = (inp[8]) ? 3'b010 : 3'b000;
								assign node185 = (inp[10]) ? node187 : 3'b010;
									assign node187 = (inp[8]) ? 3'b010 : 3'b100;
							assign node190 = (inp[10]) ? node204 : node191;
								assign node191 = (inp[4]) ? node199 : node192;
									assign node192 = (inp[8]) ? 3'b110 : node193;
										assign node193 = (inp[5]) ? 3'b100 : node194;
											assign node194 = (inp[3]) ? 3'b100 : 3'b110;
									assign node199 = (inp[8]) ? 3'b100 : node200;
										assign node200 = (inp[3]) ? 3'b110 : 3'b100;
								assign node204 = (inp[3]) ? 3'b010 : 3'b000;
			assign node207 = (inp[0]) ? node307 : node208;
				assign node208 = (inp[2]) ? node252 : node209;
					assign node209 = (inp[11]) ? node227 : node210;
						assign node210 = (inp[3]) ? node220 : node211;
							assign node211 = (inp[5]) ? 3'b010 : node212;
								assign node212 = (inp[10]) ? 3'b100 : node213;
									assign node213 = (inp[1]) ? 3'b000 : node214;
										assign node214 = (inp[4]) ? 3'b000 : 3'b010;
							assign node220 = (inp[1]) ? 3'b110 : node221;
								assign node221 = (inp[5]) ? node223 : 3'b110;
									assign node223 = (inp[10]) ? 3'b010 : 3'b000;
						assign node227 = (inp[10]) ? node235 : node228;
							assign node228 = (inp[6]) ? node230 : 3'b010;
								assign node230 = (inp[8]) ? node232 : 3'b110;
									assign node232 = (inp[4]) ? 3'b100 : 3'b110;
							assign node235 = (inp[6]) ? node243 : node236;
								assign node236 = (inp[5]) ? node238 : 3'b100;
									assign node238 = (inp[8]) ? 3'b110 : node239;
										assign node239 = (inp[4]) ? 3'b110 : 3'b100;
								assign node243 = (inp[3]) ? node245 : 3'b000;
									assign node245 = (inp[4]) ? node249 : node246;
										assign node246 = (inp[8]) ? 3'b010 : 3'b000;
										assign node249 = (inp[8]) ? 3'b000 : 3'b010;
					assign node252 = (inp[8]) ? node286 : node253;
						assign node253 = (inp[3]) ? node275 : node254;
							assign node254 = (inp[4]) ? node268 : node255;
								assign node255 = (inp[5]) ? node263 : node256;
									assign node256 = (inp[6]) ? node260 : node257;
										assign node257 = (inp[10]) ? 3'b110 : 3'b010;
										assign node260 = (inp[10]) ? 3'b010 : 3'b110;
									assign node263 = (inp[11]) ? node265 : 3'b010;
										assign node265 = (inp[10]) ? 3'b100 : 3'b010;
								assign node268 = (inp[6]) ? node272 : node269;
									assign node269 = (inp[1]) ? 3'b000 : 3'b100;
									assign node272 = (inp[10]) ? 3'b011 : 3'b111;
							assign node275 = (inp[6]) ? node279 : node276;
								assign node276 = (inp[11]) ? 3'b010 : 3'b000;
								assign node279 = (inp[4]) ? 3'b111 : node280;
									assign node280 = (inp[10]) ? node282 : 3'b100;
										assign node282 = (inp[1]) ? 3'b000 : 3'b100;
						assign node286 = (inp[4]) ? node294 : node287;
							assign node287 = (inp[5]) ? node289 : 3'b000;
								assign node289 = (inp[3]) ? 3'b011 : node290;
									assign node290 = (inp[11]) ? 3'b111 : 3'b011;
							assign node294 = (inp[3]) ? node304 : node295;
								assign node295 = (inp[1]) ? node301 : node296;
									assign node296 = (inp[11]) ? node298 : 3'b011;
										assign node298 = (inp[6]) ? 3'b101 : 3'b011;
									assign node301 = (inp[5]) ? 3'b101 : 3'b111;
								assign node304 = (inp[10]) ? 3'b001 : 3'b101;
				assign node307 = (inp[2]) ? node351 : node308;
					assign node308 = (inp[4]) ? node332 : node309;
						assign node309 = (inp[3]) ? node323 : node310;
							assign node310 = (inp[11]) ? node318 : node311;
								assign node311 = (inp[1]) ? node315 : node312;
									assign node312 = (inp[6]) ? 3'b000 : 3'b100;
									assign node315 = (inp[8]) ? 3'b111 : 3'b100;
								assign node318 = (inp[10]) ? node320 : 3'b000;
									assign node320 = (inp[6]) ? 3'b000 : 3'b100;
							assign node323 = (inp[8]) ? node329 : node324;
								assign node324 = (inp[6]) ? node326 : 3'b010;
									assign node326 = (inp[1]) ? 3'b000 : 3'b100;
								assign node329 = (inp[5]) ? 3'b011 : 3'b111;
						assign node332 = (inp[8]) ? node340 : node333;
							assign node333 = (inp[11]) ? node337 : node334;
								assign node334 = (inp[1]) ? 3'b111 : 3'b100;
								assign node337 = (inp[1]) ? 3'b111 : 3'b011;
							assign node340 = (inp[6]) ? node346 : node341;
								assign node341 = (inp[5]) ? node343 : 3'b011;
									assign node343 = (inp[10]) ? 3'b101 : 3'b001;
								assign node346 = (inp[1]) ? node348 : 3'b101;
									assign node348 = (inp[3]) ? 3'b101 : 3'b001;
					assign node351 = (inp[10]) ? node365 : node352;
						assign node352 = (inp[4]) ? 3'b101 : node353;
							assign node353 = (inp[11]) ? node361 : node354;
								assign node354 = (inp[3]) ? node358 : node355;
									assign node355 = (inp[5]) ? 3'b001 : 3'b011;
									assign node358 = (inp[5]) ? 3'b011 : 3'b101;
								assign node361 = (inp[8]) ? 3'b111 : 3'b101;
						assign node365 = (inp[6]) ? node373 : node366;
							assign node366 = (inp[11]) ? 3'b111 : node367;
								assign node367 = (inp[1]) ? node369 : 3'b011;
									assign node369 = (inp[4]) ? 3'b111 : 3'b101;
							assign node373 = (inp[11]) ? node377 : node374;
								assign node374 = (inp[4]) ? 3'b001 : 3'b011;
								assign node377 = (inp[5]) ? node379 : 3'b011;
									assign node379 = (inp[1]) ? node381 : 3'b011;
										assign node381 = (inp[3]) ? 3'b011 : 3'b001;
		assign node384 = (inp[6]) ? node556 : node385;
			assign node385 = (inp[10]) ? node479 : node386;
				assign node386 = (inp[11]) ? node430 : node387;
					assign node387 = (inp[1]) ? node405 : node388;
						assign node388 = (inp[5]) ? node398 : node389;
							assign node389 = (inp[3]) ? 3'b101 : node390;
								assign node390 = (inp[2]) ? node392 : 3'b100;
									assign node392 = (inp[7]) ? 3'b110 : node393;
										assign node393 = (inp[8]) ? 3'b100 : 3'b110;
							assign node398 = (inp[8]) ? 3'b111 : node399;
								assign node399 = (inp[3]) ? 3'b101 : node400;
									assign node400 = (inp[4]) ? 3'b101 : 3'b111;
						assign node405 = (inp[4]) ? node417 : node406;
							assign node406 = (inp[5]) ? node412 : node407;
								assign node407 = (inp[0]) ? node409 : 3'b010;
									assign node409 = (inp[8]) ? 3'b001 : 3'b011;
								assign node412 = (inp[2]) ? node414 : 3'b011;
									assign node414 = (inp[8]) ? 3'b000 : 3'b001;
							assign node417 = (inp[7]) ? node419 : 3'b010;
								assign node419 = (inp[0]) ? node421 : 3'b001;
									assign node421 = (inp[3]) ? node425 : node422;
										assign node422 = (inp[2]) ? 3'b000 : 3'b001;
										assign node425 = (inp[8]) ? 3'b000 : node426;
											assign node426 = (inp[5]) ? 3'b010 : 3'b000;
					assign node430 = (inp[1]) ? node452 : node431;
						assign node431 = (inp[7]) ? node443 : node432;
							assign node432 = (inp[0]) ? node440 : node433;
								assign node433 = (inp[2]) ? 3'b010 : node434;
									assign node434 = (inp[4]) ? node436 : 3'b000;
										assign node436 = (inp[5]) ? 3'b000 : 3'b010;
								assign node440 = (inp[2]) ? 3'b011 : 3'b010;
							assign node443 = (inp[4]) ? node445 : 3'b001;
								assign node445 = (inp[0]) ? 3'b000 : node446;
									assign node446 = (inp[8]) ? 3'b010 : node447;
										assign node447 = (inp[2]) ? 3'b001 : 3'b011;
						assign node452 = (inp[2]) ? node468 : node453;
							assign node453 = (inp[4]) ? node461 : node454;
								assign node454 = (inp[0]) ? 3'b010 : node455;
									assign node455 = (inp[8]) ? node457 : 3'b011;
										assign node457 = (inp[3]) ? 3'b011 : 3'b001;
								assign node461 = (inp[8]) ? node463 : 3'b000;
									assign node463 = (inp[3]) ? 3'b010 : node464;
										assign node464 = (inp[0]) ? 3'b011 : 3'b010;
							assign node468 = (inp[3]) ? node476 : node469;
								assign node469 = (inp[5]) ? node471 : 3'b011;
									assign node471 = (inp[8]) ? node473 : 3'b010;
										assign node473 = (inp[4]) ? 3'b010 : 3'b000;
								assign node476 = (inp[8]) ? 3'b000 : 3'b001;
				assign node479 = (inp[11]) ? node533 : node480;
					assign node480 = (inp[1]) ? node506 : node481;
						assign node481 = (inp[5]) ? node497 : node482;
							assign node482 = (inp[3]) ? node488 : node483;
								assign node483 = (inp[2]) ? node485 : 3'b010;
									assign node485 = (inp[0]) ? 3'b010 : 3'b011;
								assign node488 = (inp[4]) ? node494 : node489;
									assign node489 = (inp[7]) ? node491 : 3'b000;
										assign node491 = (inp[8]) ? 3'b001 : 3'b011;
									assign node494 = (inp[7]) ? 3'b010 : 3'b011;
							assign node497 = (inp[4]) ? node503 : node498;
								assign node498 = (inp[7]) ? 3'b000 : node499;
									assign node499 = (inp[3]) ? 3'b000 : 3'b010;
								assign node503 = (inp[8]) ? 3'b011 : 3'b000;
						assign node506 = (inp[4]) ? node520 : node507;
							assign node507 = (inp[3]) ? node513 : node508;
								assign node508 = (inp[0]) ? 3'b100 : node509;
									assign node509 = (inp[8]) ? 3'b101 : 3'b111;
								assign node513 = (inp[0]) ? node517 : node514;
									assign node514 = (inp[7]) ? 3'b111 : 3'b110;
									assign node517 = (inp[7]) ? 3'b110 : 3'b111;
							assign node520 = (inp[8]) ? node526 : node521;
								assign node521 = (inp[5]) ? node523 : 3'b101;
									assign node523 = (inp[7]) ? 3'b110 : 3'b111;
								assign node526 = (inp[7]) ? node530 : node527;
									assign node527 = (inp[3]) ? 3'b100 : 3'b110;
									assign node530 = (inp[5]) ? 3'b100 : 3'b101;
					assign node533 = (inp[7]) ? node543 : node534;
						assign node534 = (inp[8]) ? node540 : node535;
							assign node535 = (inp[3]) ? 3'b111 : node536;
								assign node536 = (inp[0]) ? 3'b100 : 3'b110;
							assign node540 = (inp[4]) ? 3'b101 : 3'b111;
						assign node543 = (inp[0]) ? node551 : node544;
							assign node544 = (inp[5]) ? node546 : 3'b101;
								assign node546 = (inp[4]) ? 3'b110 : node547;
									assign node547 = (inp[8]) ? 3'b111 : 3'b101;
							assign node551 = (inp[4]) ? 3'b100 : node552;
								assign node552 = (inp[8]) ? 3'b101 : 3'b100;
			assign node556 = (inp[10]) ? node648 : node557;
				assign node557 = (inp[1]) ? node597 : node558;
					assign node558 = (inp[11]) ? node572 : node559;
						assign node559 = (inp[3]) ? node567 : node560;
							assign node560 = (inp[8]) ? 3'b011 : node561;
								assign node561 = (inp[5]) ? node563 : 3'b011;
									assign node563 = (inp[2]) ? 3'b011 : 3'b010;
							assign node567 = (inp[8]) ? 3'b010 : node568;
								assign node568 = (inp[2]) ? 3'b010 : 3'b001;
						assign node572 = (inp[4]) ? node582 : node573;
							assign node573 = (inp[2]) ? node575 : 3'b100;
								assign node575 = (inp[5]) ? node577 : 3'b100;
									assign node577 = (inp[3]) ? 3'b101 : node578;
										assign node578 = (inp[0]) ? 3'b101 : 3'b100;
							assign node582 = (inp[8]) ? node588 : node583;
								assign node583 = (inp[2]) ? 3'b110 : node584;
									assign node584 = (inp[0]) ? 3'b110 : 3'b111;
								assign node588 = (inp[3]) ? node592 : node589;
									assign node589 = (inp[5]) ? 3'b101 : 3'b111;
									assign node592 = (inp[7]) ? node594 : 3'b101;
										assign node594 = (inp[2]) ? 3'b100 : 3'b101;
					assign node597 = (inp[0]) ? node625 : node598;
						assign node598 = (inp[7]) ? node616 : node599;
							assign node599 = (inp[3]) ? node607 : node600;
								assign node600 = (inp[4]) ? 3'b100 : node601;
									assign node601 = (inp[2]) ? node603 : 3'b100;
										assign node603 = (inp[5]) ? 3'b100 : 3'b110;
								assign node607 = (inp[2]) ? node613 : node608;
									assign node608 = (inp[5]) ? node610 : 3'b110;
										assign node610 = (inp[4]) ? 3'b110 : 3'b100;
									assign node613 = (inp[5]) ? 3'b101 : 3'b100;
							assign node616 = (inp[2]) ? node622 : node617;
								assign node617 = (inp[8]) ? node619 : 3'b101;
									assign node619 = (inp[4]) ? 3'b101 : 3'b111;
								assign node622 = (inp[4]) ? 3'b100 : 3'b101;
						assign node625 = (inp[7]) ? node637 : node626;
							assign node626 = (inp[2]) ? node634 : node627;
								assign node627 = (inp[5]) ? 3'b111 : node628;
									assign node628 = (inp[8]) ? 3'b100 : node629;
										assign node629 = (inp[4]) ? 3'b100 : 3'b110;
								assign node634 = (inp[8]) ? 3'b101 : 3'b111;
							assign node637 = (inp[2]) ? node643 : node638;
								assign node638 = (inp[5]) ? node640 : 3'b101;
									assign node640 = (inp[4]) ? 3'b100 : 3'b110;
								assign node643 = (inp[8]) ? node645 : 3'b110;
									assign node645 = (inp[4]) ? 3'b110 : 3'b100;
				assign node648 = (inp[11]) ? node678 : node649;
					assign node649 = (inp[1]) ? node661 : node650;
						assign node650 = (inp[2]) ? node654 : node651;
							assign node651 = (inp[8]) ? 3'b110 : 3'b111;
							assign node654 = (inp[7]) ? node658 : node655;
								assign node655 = (inp[3]) ? 3'b111 : 3'b101;
								assign node658 = (inp[0]) ? 3'b100 : 3'b101;
						assign node661 = (inp[0]) ? node665 : node662;
							assign node662 = (inp[8]) ? 3'b010 : 3'b000;
							assign node665 = (inp[5]) ? node671 : node666;
								assign node666 = (inp[4]) ? 3'b010 : node667;
									assign node667 = (inp[3]) ? 3'b010 : 3'b001;
								assign node671 = (inp[8]) ? node675 : node672;
									assign node672 = (inp[7]) ? 3'b001 : 3'b011;
									assign node675 = (inp[7]) ? 3'b000 : 3'b001;
					assign node678 = (inp[0]) ? node696 : node679;
						assign node679 = (inp[3]) ? node687 : node680;
							assign node680 = (inp[5]) ? 3'b011 : node681;
								assign node681 = (inp[1]) ? 3'b000 : node682;
									assign node682 = (inp[8]) ? 3'b001 : 3'b011;
							assign node687 = (inp[2]) ? node691 : node688;
								assign node688 = (inp[7]) ? 3'b001 : 3'b000;
								assign node691 = (inp[5]) ? 3'b001 : node692;
									assign node692 = (inp[8]) ? 3'b010 : 3'b001;
						assign node696 = (inp[7]) ? node704 : node697;
							assign node697 = (inp[5]) ? node701 : node698;
								assign node698 = (inp[2]) ? 3'b001 : 3'b000;
								assign node701 = (inp[8]) ? 3'b001 : 3'b011;
							assign node704 = (inp[4]) ? 3'b000 : node705;
								assign node705 = (inp[8]) ? node709 : node706;
									assign node706 = (inp[2]) ? 3'b000 : 3'b001;
									assign node709 = (inp[3]) ? 3'b010 : 3'b000;

endmodule