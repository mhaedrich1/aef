module dtc_split33_bm90 (
	input  wire [12-1:0] inp,
	output wire [3-1:0] outp
);

	wire [3-1:0] node1;
	wire [3-1:0] node2;
	wire [3-1:0] node3;
	wire [3-1:0] node5;
	wire [3-1:0] node7;
	wire [3-1:0] node9;
	wire [3-1:0] node11;
	wire [3-1:0] node14;
	wire [3-1:0] node15;
	wire [3-1:0] node16;
	wire [3-1:0] node18;
	wire [3-1:0] node19;
	wire [3-1:0] node21;
	wire [3-1:0] node25;
	wire [3-1:0] node27;
	wire [3-1:0] node28;
	wire [3-1:0] node30;
	wire [3-1:0] node33;
	wire [3-1:0] node35;
	wire [3-1:0] node39;
	wire [3-1:0] node40;
	wire [3-1:0] node41;
	wire [3-1:0] node42;
	wire [3-1:0] node43;
	wire [3-1:0] node44;
	wire [3-1:0] node45;
	wire [3-1:0] node48;
	wire [3-1:0] node51;
	wire [3-1:0] node52;
	wire [3-1:0] node55;
	wire [3-1:0] node58;
	wire [3-1:0] node59;
	wire [3-1:0] node60;
	wire [3-1:0] node64;
	wire [3-1:0] node65;
	wire [3-1:0] node68;
	wire [3-1:0] node71;
	wire [3-1:0] node72;
	wire [3-1:0] node73;
	wire [3-1:0] node74;
	wire [3-1:0] node78;
	wire [3-1:0] node79;
	wire [3-1:0] node82;
	wire [3-1:0] node85;
	wire [3-1:0] node86;
	wire [3-1:0] node87;
	wire [3-1:0] node91;
	wire [3-1:0] node92;
	wire [3-1:0] node95;
	wire [3-1:0] node98;
	wire [3-1:0] node99;
	wire [3-1:0] node100;
	wire [3-1:0] node101;
	wire [3-1:0] node102;
	wire [3-1:0] node106;
	wire [3-1:0] node107;
	wire [3-1:0] node110;
	wire [3-1:0] node113;
	wire [3-1:0] node114;
	wire [3-1:0] node115;
	wire [3-1:0] node118;
	wire [3-1:0] node122;
	wire [3-1:0] node123;
	wire [3-1:0] node124;
	wire [3-1:0] node125;
	wire [3-1:0] node128;
	wire [3-1:0] node131;
	wire [3-1:0] node132;
	wire [3-1:0] node135;
	wire [3-1:0] node138;
	wire [3-1:0] node139;
	wire [3-1:0] node140;
	wire [3-1:0] node143;
	wire [3-1:0] node146;
	wire [3-1:0] node147;
	wire [3-1:0] node150;
	wire [3-1:0] node153;
	wire [3-1:0] node154;
	wire [3-1:0] node155;
	wire [3-1:0] node156;
	wire [3-1:0] node157;
	wire [3-1:0] node158;
	wire [3-1:0] node161;
	wire [3-1:0] node165;
	wire [3-1:0] node166;
	wire [3-1:0] node167;
	wire [3-1:0] node170;
	wire [3-1:0] node173;
	wire [3-1:0] node174;
	wire [3-1:0] node177;
	wire [3-1:0] node180;
	wire [3-1:0] node181;
	wire [3-1:0] node182;
	wire [3-1:0] node183;
	wire [3-1:0] node186;
	wire [3-1:0] node189;
	wire [3-1:0] node190;
	wire [3-1:0] node194;
	wire [3-1:0] node195;
	wire [3-1:0] node196;
	wire [3-1:0] node199;
	wire [3-1:0] node202;
	wire [3-1:0] node203;
	wire [3-1:0] node206;
	wire [3-1:0] node209;
	wire [3-1:0] node210;
	wire [3-1:0] node211;
	wire [3-1:0] node212;
	wire [3-1:0] node213;
	wire [3-1:0] node216;
	wire [3-1:0] node219;
	wire [3-1:0] node221;
	wire [3-1:0] node224;
	wire [3-1:0] node225;
	wire [3-1:0] node226;
	wire [3-1:0] node230;
	wire [3-1:0] node231;
	wire [3-1:0] node234;
	wire [3-1:0] node237;
	wire [3-1:0] node238;
	wire [3-1:0] node239;
	wire [3-1:0] node240;
	wire [3-1:0] node243;
	wire [3-1:0] node246;
	wire [3-1:0] node247;
	wire [3-1:0] node250;
	wire [3-1:0] node253;
	wire [3-1:0] node254;
	wire [3-1:0] node255;
	wire [3-1:0] node258;
	wire [3-1:0] node261;
	wire [3-1:0] node262;
	wire [3-1:0] node265;
	wire [3-1:0] node268;
	wire [3-1:0] node269;
	wire [3-1:0] node270;
	wire [3-1:0] node271;
	wire [3-1:0] node272;
	wire [3-1:0] node273;
	wire [3-1:0] node274;
	wire [3-1:0] node275;
	wire [3-1:0] node278;
	wire [3-1:0] node281;
	wire [3-1:0] node282;
	wire [3-1:0] node285;
	wire [3-1:0] node288;
	wire [3-1:0] node289;
	wire [3-1:0] node290;
	wire [3-1:0] node293;
	wire [3-1:0] node296;
	wire [3-1:0] node298;
	wire [3-1:0] node301;
	wire [3-1:0] node302;
	wire [3-1:0] node304;
	wire [3-1:0] node306;
	wire [3-1:0] node309;
	wire [3-1:0] node310;
	wire [3-1:0] node311;
	wire [3-1:0] node314;
	wire [3-1:0] node317;
	wire [3-1:0] node318;
	wire [3-1:0] node321;
	wire [3-1:0] node324;
	wire [3-1:0] node325;
	wire [3-1:0] node326;
	wire [3-1:0] node327;
	wire [3-1:0] node329;
	wire [3-1:0] node332;
	wire [3-1:0] node334;
	wire [3-1:0] node337;
	wire [3-1:0] node338;
	wire [3-1:0] node339;
	wire [3-1:0] node342;
	wire [3-1:0] node345;
	wire [3-1:0] node346;
	wire [3-1:0] node349;
	wire [3-1:0] node352;
	wire [3-1:0] node353;
	wire [3-1:0] node354;
	wire [3-1:0] node355;
	wire [3-1:0] node359;
	wire [3-1:0] node360;
	wire [3-1:0] node363;
	wire [3-1:0] node366;
	wire [3-1:0] node367;
	wire [3-1:0] node368;
	wire [3-1:0] node371;
	wire [3-1:0] node374;
	wire [3-1:0] node375;
	wire [3-1:0] node379;
	wire [3-1:0] node380;
	wire [3-1:0] node381;
	wire [3-1:0] node382;
	wire [3-1:0] node383;
	wire [3-1:0] node384;
	wire [3-1:0] node387;
	wire [3-1:0] node391;
	wire [3-1:0] node392;
	wire [3-1:0] node393;
	wire [3-1:0] node397;
	wire [3-1:0] node398;
	wire [3-1:0] node401;
	wire [3-1:0] node404;
	wire [3-1:0] node405;
	wire [3-1:0] node406;
	wire [3-1:0] node407;
	wire [3-1:0] node410;
	wire [3-1:0] node413;
	wire [3-1:0] node414;
	wire [3-1:0] node417;
	wire [3-1:0] node420;
	wire [3-1:0] node421;
	wire [3-1:0] node422;
	wire [3-1:0] node425;
	wire [3-1:0] node428;
	wire [3-1:0] node429;
	wire [3-1:0] node432;
	wire [3-1:0] node435;
	wire [3-1:0] node436;
	wire [3-1:0] node437;
	wire [3-1:0] node438;
	wire [3-1:0] node439;
	wire [3-1:0] node442;
	wire [3-1:0] node445;
	wire [3-1:0] node446;
	wire [3-1:0] node449;
	wire [3-1:0] node452;
	wire [3-1:0] node453;
	wire [3-1:0] node455;
	wire [3-1:0] node459;
	wire [3-1:0] node460;
	wire [3-1:0] node461;
	wire [3-1:0] node462;
	wire [3-1:0] node465;
	wire [3-1:0] node468;
	wire [3-1:0] node469;
	wire [3-1:0] node472;
	wire [3-1:0] node475;
	wire [3-1:0] node476;
	wire [3-1:0] node477;
	wire [3-1:0] node480;
	wire [3-1:0] node483;
	wire [3-1:0] node484;
	wire [3-1:0] node488;
	wire [3-1:0] node489;
	wire [3-1:0] node490;
	wire [3-1:0] node491;
	wire [3-1:0] node492;
	wire [3-1:0] node493;
	wire [3-1:0] node494;
	wire [3-1:0] node497;
	wire [3-1:0] node500;
	wire [3-1:0] node502;
	wire [3-1:0] node505;
	wire [3-1:0] node506;
	wire [3-1:0] node508;
	wire [3-1:0] node511;
	wire [3-1:0] node512;
	wire [3-1:0] node515;
	wire [3-1:0] node518;
	wire [3-1:0] node519;
	wire [3-1:0] node520;
	wire [3-1:0] node521;
	wire [3-1:0] node524;
	wire [3-1:0] node527;
	wire [3-1:0] node528;
	wire [3-1:0] node531;
	wire [3-1:0] node534;
	wire [3-1:0] node535;
	wire [3-1:0] node537;
	wire [3-1:0] node540;
	wire [3-1:0] node541;
	wire [3-1:0] node545;
	wire [3-1:0] node546;
	wire [3-1:0] node547;
	wire [3-1:0] node549;
	wire [3-1:0] node551;
	wire [3-1:0] node554;
	wire [3-1:0] node555;
	wire [3-1:0] node556;
	wire [3-1:0] node560;
	wire [3-1:0] node561;
	wire [3-1:0] node565;
	wire [3-1:0] node566;
	wire [3-1:0] node567;
	wire [3-1:0] node569;
	wire [3-1:0] node572;
	wire [3-1:0] node573;
	wire [3-1:0] node576;
	wire [3-1:0] node579;
	wire [3-1:0] node580;
	wire [3-1:0] node581;
	wire [3-1:0] node584;
	wire [3-1:0] node587;
	wire [3-1:0] node588;
	wire [3-1:0] node591;
	wire [3-1:0] node594;
	wire [3-1:0] node595;
	wire [3-1:0] node596;
	wire [3-1:0] node597;
	wire [3-1:0] node599;
	wire [3-1:0] node600;
	wire [3-1:0] node605;
	wire [3-1:0] node607;
	wire [3-1:0] node608;
	wire [3-1:0] node609;
	wire [3-1:0] node612;
	wire [3-1:0] node615;
	wire [3-1:0] node617;
	wire [3-1:0] node620;
	wire [3-1:0] node621;
	wire [3-1:0] node622;
	wire [3-1:0] node623;
	wire [3-1:0] node625;
	wire [3-1:0] node629;
	wire [3-1:0] node630;
	wire [3-1:0] node631;
	wire [3-1:0] node634;
	wire [3-1:0] node637;
	wire [3-1:0] node639;
	wire [3-1:0] node642;
	wire [3-1:0] node643;
	wire [3-1:0] node644;
	wire [3-1:0] node645;
	wire [3-1:0] node648;
	wire [3-1:0] node651;
	wire [3-1:0] node652;
	wire [3-1:0] node656;
	wire [3-1:0] node657;
	wire [3-1:0] node658;
	wire [3-1:0] node661;
	wire [3-1:0] node664;
	wire [3-1:0] node665;
	wire [3-1:0] node668;

	assign outp = (inp[0]) ? node268 : node1;
		assign node1 = (inp[6]) ? node39 : node2;
			assign node2 = (inp[3]) ? node14 : node3;
				assign node3 = (inp[4]) ? node5 : 3'b011;
					assign node5 = (inp[7]) ? node7 : 3'b011;
						assign node7 = (inp[8]) ? node9 : 3'b111;
							assign node9 = (inp[2]) ? node11 : 3'b111;
								assign node11 = (inp[1]) ? 3'b011 : 3'b111;
				assign node14 = (inp[9]) ? 3'b111 : node15;
					assign node15 = (inp[1]) ? node25 : node16;
						assign node16 = (inp[2]) ? node18 : 3'b111;
							assign node18 = (inp[4]) ? 3'b111 : node19;
								assign node19 = (inp[5]) ? node21 : 3'b111;
									assign node21 = (inp[8]) ? 3'b011 : 3'b111;
						assign node25 = (inp[7]) ? node27 : 3'b111;
							assign node27 = (inp[4]) ? node33 : node28;
								assign node28 = (inp[8]) ? node30 : 3'b001;
									assign node30 = (inp[10]) ? 3'b101 : 3'b001;
								assign node33 = (inp[10]) ? node35 : 3'b011;
									assign node35 = (inp[8]) ? 3'b011 : 3'b111;
			assign node39 = (inp[7]) ? node153 : node40;
				assign node40 = (inp[3]) ? node98 : node41;
					assign node41 = (inp[4]) ? node71 : node42;
						assign node42 = (inp[8]) ? node58 : node43;
							assign node43 = (inp[9]) ? node51 : node44;
								assign node44 = (inp[5]) ? node48 : node45;
									assign node45 = (inp[11]) ? 3'b001 : 3'b101;
									assign node48 = (inp[1]) ? 3'b101 : 3'b101;
								assign node51 = (inp[2]) ? node55 : node52;
									assign node52 = (inp[1]) ? 3'b001 : 3'b001;
									assign node55 = (inp[1]) ? 3'b001 : 3'b001;
							assign node58 = (inp[2]) ? node64 : node59;
								assign node59 = (inp[5]) ? 3'b001 : node60;
									assign node60 = (inp[9]) ? 3'b001 : 3'b101;
								assign node64 = (inp[1]) ? node68 : node65;
									assign node65 = (inp[11]) ? 3'b001 : 3'b001;
									assign node68 = (inp[5]) ? 3'b010 : 3'b110;
						assign node71 = (inp[9]) ? node85 : node72;
							assign node72 = (inp[2]) ? node78 : node73;
								assign node73 = (inp[8]) ? 3'b011 : node74;
									assign node74 = (inp[11]) ? 3'b001 : 3'b111;
								assign node78 = (inp[8]) ? node82 : node79;
									assign node79 = (inp[10]) ? 3'b001 : 3'b101;
									assign node82 = (inp[5]) ? 3'b101 : 3'b101;
							assign node85 = (inp[1]) ? node91 : node86;
								assign node86 = (inp[10]) ? 3'b111 : node87;
									assign node87 = (inp[2]) ? 3'b011 : 3'b111;
								assign node91 = (inp[10]) ? node95 : node92;
									assign node92 = (inp[11]) ? 3'b001 : 3'b101;
									assign node95 = (inp[11]) ? 3'b101 : 3'b001;
					assign node98 = (inp[1]) ? node122 : node99;
						assign node99 = (inp[5]) ? node113 : node100;
							assign node100 = (inp[8]) ? node106 : node101;
								assign node101 = (inp[10]) ? 3'b111 : node102;
									assign node102 = (inp[4]) ? 3'b111 : 3'b101;
								assign node106 = (inp[4]) ? node110 : node107;
									assign node107 = (inp[2]) ? 3'b101 : 3'b111;
									assign node110 = (inp[10]) ? 3'b101 : 3'b101;
							assign node113 = (inp[9]) ? 3'b111 : node114;
								assign node114 = (inp[2]) ? node118 : node115;
									assign node115 = (inp[4]) ? 3'b111 : 3'b111;
									assign node118 = (inp[4]) ? 3'b111 : 3'b011;
						assign node122 = (inp[9]) ? node138 : node123;
							assign node123 = (inp[4]) ? node131 : node124;
								assign node124 = (inp[11]) ? node128 : node125;
									assign node125 = (inp[10]) ? 3'b010 : 3'b001;
									assign node128 = (inp[5]) ? 3'b101 : 3'b100;
								assign node131 = (inp[5]) ? node135 : node132;
									assign node132 = (inp[11]) ? 3'b001 : 3'b001;
									assign node135 = (inp[8]) ? 3'b101 : 3'b111;
							assign node138 = (inp[4]) ? node146 : node139;
								assign node139 = (inp[2]) ? node143 : node140;
									assign node140 = (inp[5]) ? 3'b111 : 3'b001;
									assign node143 = (inp[8]) ? 3'b011 : 3'b001;
								assign node146 = (inp[11]) ? node150 : node147;
									assign node147 = (inp[5]) ? 3'b011 : 3'b011;
									assign node150 = (inp[10]) ? 3'b001 : 3'b111;
				assign node153 = (inp[3]) ? node209 : node154;
					assign node154 = (inp[4]) ? node180 : node155;
						assign node155 = (inp[9]) ? node165 : node156;
							assign node156 = (inp[1]) ? 3'b000 : node157;
								assign node157 = (inp[10]) ? node161 : node158;
									assign node158 = (inp[2]) ? 3'b000 : 3'b000;
									assign node161 = (inp[8]) ? 3'b100 : 3'b000;
							assign node165 = (inp[2]) ? node173 : node166;
								assign node166 = (inp[5]) ? node170 : node167;
									assign node167 = (inp[8]) ? 3'b000 : 3'b110;
									assign node170 = (inp[8]) ? 3'b110 : 3'b001;
								assign node173 = (inp[5]) ? node177 : node174;
									assign node174 = (inp[1]) ? 3'b000 : 3'b010;
									assign node177 = (inp[1]) ? 3'b110 : 3'b100;
						assign node180 = (inp[1]) ? node194 : node181;
							assign node181 = (inp[9]) ? node189 : node182;
								assign node182 = (inp[2]) ? node186 : node183;
									assign node183 = (inp[10]) ? 3'b001 : 3'b011;
									assign node186 = (inp[10]) ? 3'b000 : 3'b010;
								assign node189 = (inp[8]) ? 3'b001 : node190;
									assign node190 = (inp[2]) ? 3'b111 : 3'b011;
							assign node194 = (inp[9]) ? node202 : node195;
								assign node195 = (inp[10]) ? node199 : node196;
									assign node196 = (inp[2]) ? 3'b000 : 3'b000;
									assign node199 = (inp[11]) ? 3'b000 : 3'b100;
								assign node202 = (inp[8]) ? node206 : node203;
									assign node203 = (inp[10]) ? 3'b001 : 3'b010;
									assign node206 = (inp[11]) ? 3'b110 : 3'b000;
					assign node209 = (inp[1]) ? node237 : node210;
						assign node210 = (inp[9]) ? node224 : node211;
							assign node211 = (inp[11]) ? node219 : node212;
								assign node212 = (inp[4]) ? node216 : node213;
									assign node213 = (inp[5]) ? 3'b001 : 3'b000;
									assign node216 = (inp[2]) ? 3'b001 : 3'b101;
								assign node219 = (inp[4]) ? node221 : 3'b101;
									assign node221 = (inp[5]) ? 3'b111 : 3'b011;
							assign node224 = (inp[2]) ? node230 : node225;
								assign node225 = (inp[10]) ? 3'b111 : node226;
									assign node226 = (inp[5]) ? 3'b101 : 3'b011;
								assign node230 = (inp[11]) ? node234 : node231;
									assign node231 = (inp[4]) ? 3'b011 : 3'b101;
									assign node234 = (inp[10]) ? 3'b011 : 3'b011;
						assign node237 = (inp[9]) ? node253 : node238;
							assign node238 = (inp[2]) ? node246 : node239;
								assign node239 = (inp[10]) ? node243 : node240;
									assign node240 = (inp[5]) ? 3'b010 : 3'b100;
									assign node243 = (inp[8]) ? 3'b001 : 3'b001;
								assign node246 = (inp[8]) ? node250 : node247;
									assign node247 = (inp[5]) ? 3'b110 : 3'b100;
									assign node250 = (inp[10]) ? 3'b010 : 3'b010;
							assign node253 = (inp[8]) ? node261 : node254;
								assign node254 = (inp[4]) ? node258 : node255;
									assign node255 = (inp[10]) ? 3'b111 : 3'b100;
									assign node258 = (inp[5]) ? 3'b011 : 3'b011;
								assign node261 = (inp[2]) ? node265 : node262;
									assign node262 = (inp[4]) ? 3'b011 : 3'b001;
									assign node265 = (inp[4]) ? 3'b101 : 3'b110;
		assign node268 = (inp[6]) ? node488 : node269;
			assign node269 = (inp[4]) ? node379 : node270;
				assign node270 = (inp[3]) ? node324 : node271;
					assign node271 = (inp[9]) ? node301 : node272;
						assign node272 = (inp[8]) ? node288 : node273;
							assign node273 = (inp[5]) ? node281 : node274;
								assign node274 = (inp[11]) ? node278 : node275;
									assign node275 = (inp[10]) ? 3'b000 : 3'b000;
									assign node278 = (inp[7]) ? 3'b000 : 3'b010;
								assign node281 = (inp[7]) ? node285 : node282;
									assign node282 = (inp[10]) ? 3'b010 : 3'b100;
									assign node285 = (inp[2]) ? 3'b010 : 3'b100;
							assign node288 = (inp[2]) ? node296 : node289;
								assign node289 = (inp[11]) ? node293 : node290;
									assign node290 = (inp[10]) ? 3'b000 : 3'b000;
									assign node293 = (inp[5]) ? 3'b110 : 3'b000;
								assign node296 = (inp[5]) ? node298 : 3'b100;
									assign node298 = (inp[1]) ? 3'b100 : 3'b000;
						assign node301 = (inp[1]) ? node309 : node302;
							assign node302 = (inp[7]) ? node304 : 3'b110;
								assign node304 = (inp[2]) ? node306 : 3'b110;
									assign node306 = (inp[10]) ? 3'b110 : 3'b010;
							assign node309 = (inp[2]) ? node317 : node310;
								assign node310 = (inp[8]) ? node314 : node311;
									assign node311 = (inp[5]) ? 3'b110 : 3'b010;
									assign node314 = (inp[5]) ? 3'b010 : 3'b010;
								assign node317 = (inp[7]) ? node321 : node318;
									assign node318 = (inp[10]) ? 3'b110 : 3'b000;
									assign node321 = (inp[10]) ? 3'b100 : 3'b110;
					assign node324 = (inp[9]) ? node352 : node325;
						assign node325 = (inp[1]) ? node337 : node326;
							assign node326 = (inp[7]) ? node332 : node327;
								assign node327 = (inp[5]) ? node329 : 3'b111;
									assign node329 = (inp[2]) ? 3'b011 : 3'b111;
								assign node332 = (inp[10]) ? node334 : 3'b110;
									assign node334 = (inp[5]) ? 3'b100 : 3'b000;
							assign node337 = (inp[8]) ? node345 : node338;
								assign node338 = (inp[5]) ? node342 : node339;
									assign node339 = (inp[7]) ? 3'b000 : 3'b010;
									assign node342 = (inp[11]) ? 3'b010 : 3'b110;
								assign node345 = (inp[5]) ? node349 : node346;
									assign node346 = (inp[10]) ? 3'b100 : 3'b000;
									assign node349 = (inp[7]) ? 3'b100 : 3'b010;
						assign node352 = (inp[7]) ? node366 : node353;
							assign node353 = (inp[1]) ? node359 : node354;
								assign node354 = (inp[10]) ? 3'b111 : node355;
									assign node355 = (inp[2]) ? 3'b011 : 3'b111;
								assign node359 = (inp[2]) ? node363 : node360;
									assign node360 = (inp[5]) ? 3'b011 : 3'b011;
									assign node363 = (inp[8]) ? 3'b001 : 3'b001;
							assign node366 = (inp[1]) ? node374 : node367;
								assign node367 = (inp[10]) ? node371 : node368;
									assign node368 = (inp[11]) ? 3'b101 : 3'b001;
									assign node371 = (inp[2]) ? 3'b011 : 3'b011;
								assign node374 = (inp[8]) ? 3'b010 : node375;
									assign node375 = (inp[10]) ? 3'b001 : 3'b000;
				assign node379 = (inp[3]) ? node435 : node380;
					assign node380 = (inp[11]) ? node404 : node381;
						assign node381 = (inp[7]) ? node391 : node382;
							assign node382 = (inp[2]) ? 3'b001 : node383;
								assign node383 = (inp[9]) ? node387 : node384;
									assign node384 = (inp[1]) ? 3'b001 : 3'b001;
									assign node387 = (inp[8]) ? 3'b001 : 3'b000;
							assign node391 = (inp[1]) ? node397 : node392;
								assign node392 = (inp[2]) ? 3'b001 : node393;
									assign node393 = (inp[10]) ? 3'b101 : 3'b001;
								assign node397 = (inp[9]) ? node401 : node398;
									assign node398 = (inp[10]) ? 3'b000 : 3'b000;
									assign node401 = (inp[8]) ? 3'b100 : 3'b010;
						assign node404 = (inp[1]) ? node420 : node405;
							assign node405 = (inp[7]) ? node413 : node406;
								assign node406 = (inp[2]) ? node410 : node407;
									assign node407 = (inp[10]) ? 3'b110 : 3'b001;
									assign node410 = (inp[5]) ? 3'b001 : 3'b000;
								assign node413 = (inp[5]) ? node417 : node414;
									assign node414 = (inp[10]) ? 3'b001 : 3'b001;
									assign node417 = (inp[8]) ? 3'b001 : 3'b011;
							assign node420 = (inp[9]) ? node428 : node421;
								assign node421 = (inp[7]) ? node425 : node422;
									assign node422 = (inp[10]) ? 3'b000 : 3'b001;
									assign node425 = (inp[2]) ? 3'b000 : 3'b000;
								assign node428 = (inp[10]) ? node432 : node429;
									assign node429 = (inp[7]) ? 3'b010 : 3'b110;
									assign node432 = (inp[5]) ? 3'b001 : 3'b100;
					assign node435 = (inp[1]) ? node459 : node436;
						assign node436 = (inp[9]) ? node452 : node437;
							assign node437 = (inp[7]) ? node445 : node438;
								assign node438 = (inp[5]) ? node442 : node439;
									assign node439 = (inp[2]) ? 3'b101 : 3'b011;
									assign node442 = (inp[8]) ? 3'b011 : 3'b111;
								assign node445 = (inp[8]) ? node449 : node446;
									assign node446 = (inp[2]) ? 3'b101 : 3'b101;
									assign node449 = (inp[2]) ? 3'b101 : 3'b001;
							assign node452 = (inp[10]) ? 3'b111 : node453;
								assign node453 = (inp[7]) ? node455 : 3'b111;
									assign node455 = (inp[2]) ? 3'b011 : 3'b111;
						assign node459 = (inp[9]) ? node475 : node460;
							assign node460 = (inp[5]) ? node468 : node461;
								assign node461 = (inp[2]) ? node465 : node462;
									assign node462 = (inp[7]) ? 3'b010 : 3'b001;
									assign node465 = (inp[8]) ? 3'b100 : 3'b010;
								assign node468 = (inp[10]) ? node472 : node469;
									assign node469 = (inp[11]) ? 3'b101 : 3'b110;
									assign node472 = (inp[11]) ? 3'b001 : 3'b011;
							assign node475 = (inp[7]) ? node483 : node476;
								assign node476 = (inp[11]) ? node480 : node477;
									assign node477 = (inp[2]) ? 3'b011 : 3'b111;
									assign node480 = (inp[8]) ? 3'b001 : 3'b011;
								assign node483 = (inp[10]) ? 3'b001 : node484;
									assign node484 = (inp[5]) ? 3'b110 : 3'b001;
			assign node488 = (inp[1]) ? node594 : node489;
				assign node489 = (inp[7]) ? node545 : node490;
					assign node490 = (inp[4]) ? node518 : node491;
						assign node491 = (inp[2]) ? node505 : node492;
							assign node492 = (inp[5]) ? node500 : node493;
								assign node493 = (inp[10]) ? node497 : node494;
									assign node494 = (inp[3]) ? 3'b100 : 3'b110;
									assign node497 = (inp[11]) ? 3'b010 : 3'b000;
								assign node500 = (inp[9]) ? node502 : 3'b010;
									assign node502 = (inp[8]) ? 3'b110 : 3'b010;
							assign node505 = (inp[10]) ? node511 : node506;
								assign node506 = (inp[8]) ? node508 : 3'b100;
									assign node508 = (inp[5]) ? 3'b000 : 3'b010;
								assign node511 = (inp[11]) ? node515 : node512;
									assign node512 = (inp[3]) ? 3'b100 : 3'b000;
									assign node515 = (inp[5]) ? 3'b100 : 3'b100;
						assign node518 = (inp[2]) ? node534 : node519;
							assign node519 = (inp[3]) ? node527 : node520;
								assign node520 = (inp[9]) ? node524 : node521;
									assign node521 = (inp[11]) ? 3'b101 : 3'b100;
									assign node524 = (inp[10]) ? 3'b110 : 3'b000;
								assign node527 = (inp[9]) ? node531 : node528;
									assign node528 = (inp[8]) ? 3'b010 : 3'b110;
									assign node531 = (inp[10]) ? 3'b111 : 3'b101;
							assign node534 = (inp[3]) ? node540 : node535;
								assign node535 = (inp[9]) ? node537 : 3'b110;
									assign node537 = (inp[8]) ? 3'b010 : 3'b110;
								assign node540 = (inp[9]) ? 3'b101 : node541;
									assign node541 = (inp[8]) ? 3'b110 : 3'b110;
					assign node545 = (inp[3]) ? node565 : node546;
						assign node546 = (inp[9]) ? node554 : node547;
							assign node547 = (inp[10]) ? node549 : 3'b000;
								assign node549 = (inp[11]) ? node551 : 3'b000;
									assign node551 = (inp[5]) ? 3'b100 : 3'b000;
							assign node554 = (inp[5]) ? node560 : node555;
								assign node555 = (inp[8]) ? 3'b000 : node556;
									assign node556 = (inp[10]) ? 3'b010 : 3'b100;
								assign node560 = (inp[2]) ? 3'b010 : node561;
									assign node561 = (inp[10]) ? 3'b000 : 3'b100;
						assign node565 = (inp[9]) ? node579 : node566;
							assign node566 = (inp[4]) ? node572 : node567;
								assign node567 = (inp[10]) ? node569 : 3'b000;
									assign node569 = (inp[2]) ? 3'b000 : 3'b100;
								assign node572 = (inp[2]) ? node576 : node573;
									assign node573 = (inp[11]) ? 3'b110 : 3'b010;
									assign node576 = (inp[10]) ? 3'b100 : 3'b000;
							assign node579 = (inp[4]) ? node587 : node580;
								assign node580 = (inp[8]) ? node584 : node581;
									assign node581 = (inp[2]) ? 3'b010 : 3'b011;
									assign node584 = (inp[2]) ? 3'b100 : 3'b110;
								assign node587 = (inp[10]) ? node591 : node588;
									assign node588 = (inp[2]) ? 3'b010 : 3'b001;
									assign node591 = (inp[2]) ? 3'b001 : 3'b001;
				assign node594 = (inp[3]) ? node620 : node595;
					assign node595 = (inp[9]) ? node605 : node596;
						assign node596 = (inp[5]) ? 3'b000 : node597;
							assign node597 = (inp[11]) ? node599 : 3'b000;
								assign node599 = (inp[2]) ? 3'b000 : node600;
									assign node600 = (inp[8]) ? 3'b000 : 3'b000;
						assign node605 = (inp[4]) ? node607 : 3'b000;
							assign node607 = (inp[8]) ? node615 : node608;
								assign node608 = (inp[5]) ? node612 : node609;
									assign node609 = (inp[7]) ? 3'b000 : 3'b000;
									assign node612 = (inp[2]) ? 3'b000 : 3'b100;
								assign node615 = (inp[10]) ? node617 : 3'b000;
									assign node617 = (inp[2]) ? 3'b000 : 3'b100;
					assign node620 = (inp[9]) ? node642 : node621;
						assign node621 = (inp[5]) ? node629 : node622;
							assign node622 = (inp[7]) ? 3'b000 : node623;
								assign node623 = (inp[4]) ? node625 : 3'b000;
									assign node625 = (inp[2]) ? 3'b000 : 3'b000;
							assign node629 = (inp[2]) ? node637 : node630;
								assign node630 = (inp[4]) ? node634 : node631;
									assign node631 = (inp[7]) ? 3'b010 : 3'b000;
									assign node634 = (inp[7]) ? 3'b000 : 3'b010;
								assign node637 = (inp[10]) ? node639 : 3'b000;
									assign node639 = (inp[7]) ? 3'b000 : 3'b100;
						assign node642 = (inp[4]) ? node656 : node643;
							assign node643 = (inp[2]) ? node651 : node644;
								assign node644 = (inp[10]) ? node648 : node645;
									assign node645 = (inp[7]) ? 3'b000 : 3'b001;
									assign node648 = (inp[11]) ? 3'b010 : 3'b010;
								assign node651 = (inp[7]) ? 3'b000 : node652;
									assign node652 = (inp[11]) ? 3'b100 : 3'b000;
							assign node656 = (inp[7]) ? node664 : node657;
								assign node657 = (inp[2]) ? node661 : node658;
									assign node658 = (inp[11]) ? 3'b001 : 3'b001;
									assign node661 = (inp[5]) ? 3'b010 : 3'b100;
								assign node664 = (inp[10]) ? node668 : node665;
									assign node665 = (inp[8]) ? 3'b000 : 3'b100;
									assign node668 = (inp[8]) ? 3'b100 : 3'b110;

endmodule