module dtc_split875_bm93 (
	input  wire [12-1:0] inp,
	output wire [3-1:0] outp
);

	wire [3-1:0] node1;
	wire [3-1:0] node2;
	wire [3-1:0] node4;
	wire [3-1:0] node5;
	wire [3-1:0] node6;
	wire [3-1:0] node7;
	wire [3-1:0] node11;
	wire [3-1:0] node12;
	wire [3-1:0] node14;
	wire [3-1:0] node17;
	wire [3-1:0] node18;
	wire [3-1:0] node24;
	wire [3-1:0] node25;
	wire [3-1:0] node26;
	wire [3-1:0] node27;
	wire [3-1:0] node29;
	wire [3-1:0] node30;
	wire [3-1:0] node34;
	wire [3-1:0] node35;
	wire [3-1:0] node36;
	wire [3-1:0] node37;
	wire [3-1:0] node38;
	wire [3-1:0] node39;
	wire [3-1:0] node43;
	wire [3-1:0] node44;
	wire [3-1:0] node46;
	wire [3-1:0] node50;
	wire [3-1:0] node51;
	wire [3-1:0] node55;
	wire [3-1:0] node56;
	wire [3-1:0] node61;
	wire [3-1:0] node62;
	wire [3-1:0] node63;
	wire [3-1:0] node64;
	wire [3-1:0] node69;
	wire [3-1:0] node70;
	wire [3-1:0] node71;
	wire [3-1:0] node72;
	wire [3-1:0] node73;
	wire [3-1:0] node74;
	wire [3-1:0] node75;
	wire [3-1:0] node84;
	wire [3-1:0] node86;
	wire [3-1:0] node87;
	wire [3-1:0] node88;
	wire [3-1:0] node90;
	wire [3-1:0] node92;
	wire [3-1:0] node93;
	wire [3-1:0] node94;
	wire [3-1:0] node95;
	wire [3-1:0] node100;
	wire [3-1:0] node103;
	wire [3-1:0] node104;
	wire [3-1:0] node106;
	wire [3-1:0] node108;
	wire [3-1:0] node109;
	wire [3-1:0] node111;
	wire [3-1:0] node115;
	wire [3-1:0] node116;
	wire [3-1:0] node118;
	wire [3-1:0] node122;
	wire [3-1:0] node124;
	wire [3-1:0] node126;
	wire [3-1:0] node128;
	wire [3-1:0] node130;
	wire [3-1:0] node131;

	assign outp = (inp[0]) ? node24 : node1;
		assign node1 = (inp[6]) ? 3'b000 : node2;
			assign node2 = (inp[3]) ? node4 : 3'b000;
				assign node4 = (inp[7]) ? 3'b000 : node5;
					assign node5 = (inp[5]) ? node11 : node6;
						assign node6 = (inp[8]) ? 3'b000 : node7;
							assign node7 = (inp[4]) ? 3'b100 : 3'b000;
						assign node11 = (inp[8]) ? node17 : node12;
							assign node12 = (inp[4]) ? node14 : 3'b010;
								assign node14 = (inp[10]) ? 3'b010 : 3'b100;
							assign node17 = (inp[10]) ? 3'b100 : node18;
								assign node18 = (inp[4]) ? 3'b000 : 3'b100;
		assign node24 = (inp[7]) ? node84 : node25;
			assign node25 = (inp[3]) ? node61 : node26;
				assign node26 = (inp[5]) ? node34 : node27;
					assign node27 = (inp[4]) ? node29 : 3'b000;
						assign node29 = (inp[6]) ? 3'b000 : node30;
							assign node30 = (inp[8]) ? 3'b000 : 3'b110;
					assign node34 = (inp[6]) ? 3'b100 : node35;
						assign node35 = (inp[8]) ? node55 : node36;
							assign node36 = (inp[10]) ? node50 : node37;
								assign node37 = (inp[4]) ? node43 : node38;
									assign node38 = (inp[2]) ? 3'b100 : node39;
										assign node39 = (inp[1]) ? 3'b100 : 3'b000;
									assign node43 = (inp[1]) ? 3'b110 : node44;
										assign node44 = (inp[11]) ? node46 : 3'b110;
											assign node46 = (inp[2]) ? 3'b110 : 3'b010;
								assign node50 = (inp[1]) ? 3'b100 : node51;
									assign node51 = (inp[2]) ? 3'b100 : 3'b000;
							assign node55 = (inp[10]) ? 3'b110 : node56;
								assign node56 = (inp[4]) ? 3'b100 : 3'b110;
				assign node61 = (inp[5]) ? node69 : node62;
					assign node62 = (inp[6]) ? 3'b011 : node63;
						assign node63 = (inp[8]) ? 3'b011 : node64;
							assign node64 = (inp[4]) ? 3'b111 : 3'b011;
					assign node69 = (inp[6]) ? 3'b110 : node70;
						assign node70 = (inp[2]) ? 3'b111 : node71;
							assign node71 = (inp[8]) ? 3'b111 : node72;
								assign node72 = (inp[1]) ? 3'b111 : node73;
									assign node73 = (inp[10]) ? 3'b011 : node74;
										assign node74 = (inp[11]) ? 3'b011 : node75;
											assign node75 = (inp[4]) ? 3'b101 : 3'b011;
			assign node84 = (inp[5]) ? node86 : 3'b000;
				assign node86 = (inp[6]) ? node122 : node87;
					assign node87 = (inp[3]) ? node103 : node88;
						assign node88 = (inp[2]) ? node90 : 3'b000;
							assign node90 = (inp[1]) ? node92 : 3'b000;
								assign node92 = (inp[8]) ? node100 : node93;
									assign node93 = (inp[11]) ? 3'b100 : node94;
										assign node94 = (inp[10]) ? 3'b100 : node95;
											assign node95 = (inp[4]) ? 3'b000 : 3'b100;
									assign node100 = (inp[11]) ? 3'b000 : 3'b100;
						assign node103 = (inp[8]) ? node115 : node104;
							assign node104 = (inp[2]) ? node106 : 3'b011;
								assign node106 = (inp[1]) ? node108 : 3'b011;
									assign node108 = (inp[11]) ? 3'b111 : node109;
										assign node109 = (inp[4]) ? node111 : 3'b111;
											assign node111 = (inp[10]) ? 3'b111 : 3'b011;
							assign node115 = (inp[11]) ? 3'b011 : node116;
								assign node116 = (inp[2]) ? node118 : 3'b001;
									assign node118 = (inp[1]) ? 3'b101 : 3'b001;
					assign node122 = (inp[4]) ? node124 : 3'b000;
						assign node124 = (inp[9]) ? node126 : 3'b000;
							assign node126 = (inp[1]) ? node128 : 3'b000;
								assign node128 = (inp[2]) ? node130 : 3'b000;
									assign node130 = (inp[10]) ? 3'b000 : node131;
										assign node131 = (inp[8]) ? 3'b100 : 3'b000;

endmodule