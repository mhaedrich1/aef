module dtc_split5_bm71 (
	input  wire [12-1:0] inp,
	output wire [3-1:0] outp
);

	wire [3-1:0] node1;
	wire [3-1:0] node2;
	wire [3-1:0] node3;
	wire [3-1:0] node4;
	wire [3-1:0] node5;
	wire [3-1:0] node6;
	wire [3-1:0] node7;
	wire [3-1:0] node8;
	wire [3-1:0] node10;
	wire [3-1:0] node13;
	wire [3-1:0] node14;
	wire [3-1:0] node15;
	wire [3-1:0] node19;
	wire [3-1:0] node22;
	wire [3-1:0] node23;
	wire [3-1:0] node25;
	wire [3-1:0] node28;
	wire [3-1:0] node29;
	wire [3-1:0] node30;
	wire [3-1:0] node35;
	wire [3-1:0] node36;
	wire [3-1:0] node37;
	wire [3-1:0] node38;
	wire [3-1:0] node40;
	wire [3-1:0] node44;
	wire [3-1:0] node46;
	wire [3-1:0] node49;
	wire [3-1:0] node50;
	wire [3-1:0] node51;
	wire [3-1:0] node55;
	wire [3-1:0] node57;
	wire [3-1:0] node60;
	wire [3-1:0] node61;
	wire [3-1:0] node62;
	wire [3-1:0] node63;
	wire [3-1:0] node64;
	wire [3-1:0] node65;
	wire [3-1:0] node71;
	wire [3-1:0] node72;
	wire [3-1:0] node74;
	wire [3-1:0] node76;
	wire [3-1:0] node81;
	wire [3-1:0] node82;
	wire [3-1:0] node83;
	wire [3-1:0] node84;
	wire [3-1:0] node85;
	wire [3-1:0] node87;
	wire [3-1:0] node89;
	wire [3-1:0] node92;
	wire [3-1:0] node93;
	wire [3-1:0] node96;
	wire [3-1:0] node99;
	wire [3-1:0] node100;
	wire [3-1:0] node101;
	wire [3-1:0] node103;
	wire [3-1:0] node106;
	wire [3-1:0] node108;
	wire [3-1:0] node111;
	wire [3-1:0] node112;
	wire [3-1:0] node115;
	wire [3-1:0] node117;
	wire [3-1:0] node120;
	wire [3-1:0] node121;
	wire [3-1:0] node122;
	wire [3-1:0] node124;
	wire [3-1:0] node125;
	wire [3-1:0] node129;
	wire [3-1:0] node131;
	wire [3-1:0] node134;
	wire [3-1:0] node135;
	wire [3-1:0] node137;
	wire [3-1:0] node140;
	wire [3-1:0] node142;
	wire [3-1:0] node145;
	wire [3-1:0] node146;
	wire [3-1:0] node147;
	wire [3-1:0] node148;
	wire [3-1:0] node149;
	wire [3-1:0] node150;
	wire [3-1:0] node154;
	wire [3-1:0] node157;
	wire [3-1:0] node159;
	wire [3-1:0] node161;
	wire [3-1:0] node164;
	wire [3-1:0] node165;
	wire [3-1:0] node166;
	wire [3-1:0] node170;
	wire [3-1:0] node173;
	wire [3-1:0] node174;
	wire [3-1:0] node175;
	wire [3-1:0] node177;
	wire [3-1:0] node181;
	wire [3-1:0] node182;
	wire [3-1:0] node183;
	wire [3-1:0] node184;
	wire [3-1:0] node188;
	wire [3-1:0] node191;
	wire [3-1:0] node193;
	wire [3-1:0] node195;
	wire [3-1:0] node198;
	wire [3-1:0] node199;
	wire [3-1:0] node200;
	wire [3-1:0] node202;
	wire [3-1:0] node203;
	wire [3-1:0] node204;
	wire [3-1:0] node210;
	wire [3-1:0] node211;
	wire [3-1:0] node212;
	wire [3-1:0] node213;
	wire [3-1:0] node214;
	wire [3-1:0] node215;
	wire [3-1:0] node217;
	wire [3-1:0] node221;
	wire [3-1:0] node223;
	wire [3-1:0] node224;
	wire [3-1:0] node228;
	wire [3-1:0] node229;
	wire [3-1:0] node231;
	wire [3-1:0] node234;
	wire [3-1:0] node236;
	wire [3-1:0] node239;
	wire [3-1:0] node240;
	wire [3-1:0] node241;
	wire [3-1:0] node242;
	wire [3-1:0] node246;
	wire [3-1:0] node247;
	wire [3-1:0] node251;
	wire [3-1:0] node252;
	wire [3-1:0] node253;
	wire [3-1:0] node258;
	wire [3-1:0] node259;
	wire [3-1:0] node261;
	wire [3-1:0] node262;
	wire [3-1:0] node264;
	wire [3-1:0] node265;
	wire [3-1:0] node271;
	wire [3-1:0] node273;
	wire [3-1:0] node274;
	wire [3-1:0] node275;
	wire [3-1:0] node276;
	wire [3-1:0] node277;
	wire [3-1:0] node278;
	wire [3-1:0] node282;
	wire [3-1:0] node283;
	wire [3-1:0] node284;
	wire [3-1:0] node288;
	wire [3-1:0] node289;
	wire [3-1:0] node293;
	wire [3-1:0] node294;
	wire [3-1:0] node295;
	wire [3-1:0] node302;
	wire [3-1:0] node303;
	wire [3-1:0] node304;
	wire [3-1:0] node305;
	wire [3-1:0] node306;
	wire [3-1:0] node307;
	wire [3-1:0] node308;
	wire [3-1:0] node309;
	wire [3-1:0] node310;
	wire [3-1:0] node314;
	wire [3-1:0] node317;
	wire [3-1:0] node319;
	wire [3-1:0] node320;
	wire [3-1:0] node324;
	wire [3-1:0] node325;
	wire [3-1:0] node326;
	wire [3-1:0] node327;
	wire [3-1:0] node328;
	wire [3-1:0] node331;
	wire [3-1:0] node335;
	wire [3-1:0] node336;
	wire [3-1:0] node338;
	wire [3-1:0] node341;
	wire [3-1:0] node344;
	wire [3-1:0] node346;
	wire [3-1:0] node347;
	wire [3-1:0] node350;
	wire [3-1:0] node352;
	wire [3-1:0] node355;
	wire [3-1:0] node356;
	wire [3-1:0] node357;
	wire [3-1:0] node358;
	wire [3-1:0] node359;
	wire [3-1:0] node363;
	wire [3-1:0] node366;
	wire [3-1:0] node367;
	wire [3-1:0] node368;
	wire [3-1:0] node372;
	wire [3-1:0] node374;
	wire [3-1:0] node375;
	wire [3-1:0] node379;
	wire [3-1:0] node380;
	wire [3-1:0] node381;
	wire [3-1:0] node382;
	wire [3-1:0] node384;
	wire [3-1:0] node387;
	wire [3-1:0] node389;
	wire [3-1:0] node392;
	wire [3-1:0] node393;
	wire [3-1:0] node397;
	wire [3-1:0] node398;
	wire [3-1:0] node401;
	wire [3-1:0] node402;
	wire [3-1:0] node404;
	wire [3-1:0] node408;
	wire [3-1:0] node409;
	wire [3-1:0] node410;
	wire [3-1:0] node412;
	wire [3-1:0] node416;
	wire [3-1:0] node417;
	wire [3-1:0] node418;
	wire [3-1:0] node420;
	wire [3-1:0] node423;
	wire [3-1:0] node424;
	wire [3-1:0] node427;
	wire [3-1:0] node428;
	wire [3-1:0] node429;
	wire [3-1:0] node434;
	wire [3-1:0] node435;
	wire [3-1:0] node436;
	wire [3-1:0] node437;
	wire [3-1:0] node441;
	wire [3-1:0] node442;
	wire [3-1:0] node446;
	wire [3-1:0] node447;
	wire [3-1:0] node448;
	wire [3-1:0] node452;
	wire [3-1:0] node455;
	wire [3-1:0] node456;
	wire [3-1:0] node457;
	wire [3-1:0] node458;
	wire [3-1:0] node459;
	wire [3-1:0] node460;
	wire [3-1:0] node463;
	wire [3-1:0] node466;
	wire [3-1:0] node467;
	wire [3-1:0] node469;
	wire [3-1:0] node471;
	wire [3-1:0] node474;
	wire [3-1:0] node475;
	wire [3-1:0] node477;
	wire [3-1:0] node481;
	wire [3-1:0] node482;
	wire [3-1:0] node483;
	wire [3-1:0] node484;
	wire [3-1:0] node485;
	wire [3-1:0] node489;
	wire [3-1:0] node490;
	wire [3-1:0] node494;
	wire [3-1:0] node497;
	wire [3-1:0] node498;
	wire [3-1:0] node499;
	wire [3-1:0] node502;
	wire [3-1:0] node506;
	wire [3-1:0] node507;
	wire [3-1:0] node508;
	wire [3-1:0] node509;
	wire [3-1:0] node511;
	wire [3-1:0] node515;
	wire [3-1:0] node516;
	wire [3-1:0] node518;
	wire [3-1:0] node521;
	wire [3-1:0] node522;
	wire [3-1:0] node524;
	wire [3-1:0] node528;
	wire [3-1:0] node529;
	wire [3-1:0] node530;
	wire [3-1:0] node531;
	wire [3-1:0] node533;
	wire [3-1:0] node538;
	wire [3-1:0] node539;
	wire [3-1:0] node541;
	wire [3-1:0] node542;
	wire [3-1:0] node546;
	wire [3-1:0] node549;
	wire [3-1:0] node550;
	wire [3-1:0] node551;
	wire [3-1:0] node552;
	wire [3-1:0] node553;
	wire [3-1:0] node554;
	wire [3-1:0] node557;
	wire [3-1:0] node560;
	wire [3-1:0] node562;
	wire [3-1:0] node565;
	wire [3-1:0] node566;
	wire [3-1:0] node568;
	wire [3-1:0] node570;
	wire [3-1:0] node573;
	wire [3-1:0] node575;
	wire [3-1:0] node577;
	wire [3-1:0] node580;
	wire [3-1:0] node581;
	wire [3-1:0] node582;
	wire [3-1:0] node584;
	wire [3-1:0] node585;
	wire [3-1:0] node589;
	wire [3-1:0] node591;
	wire [3-1:0] node594;
	wire [3-1:0] node595;
	wire [3-1:0] node598;
	wire [3-1:0] node600;
	wire [3-1:0] node602;
	wire [3-1:0] node605;
	wire [3-1:0] node606;
	wire [3-1:0] node607;
	wire [3-1:0] node608;
	wire [3-1:0] node610;
	wire [3-1:0] node611;
	wire [3-1:0] node615;
	wire [3-1:0] node617;
	wire [3-1:0] node620;
	wire [3-1:0] node621;
	wire [3-1:0] node622;
	wire [3-1:0] node624;
	wire [3-1:0] node627;
	wire [3-1:0] node629;
	wire [3-1:0] node632;
	wire [3-1:0] node633;
	wire [3-1:0] node636;
	wire [3-1:0] node639;
	wire [3-1:0] node640;
	wire [3-1:0] node641;
	wire [3-1:0] node644;
	wire [3-1:0] node647;
	wire [3-1:0] node648;
	wire [3-1:0] node650;
	wire [3-1:0] node653;
	wire [3-1:0] node655;
	wire [3-1:0] node658;
	wire [3-1:0] node659;
	wire [3-1:0] node660;
	wire [3-1:0] node661;
	wire [3-1:0] node662;
	wire [3-1:0] node663;
	wire [3-1:0] node664;
	wire [3-1:0] node665;
	wire [3-1:0] node667;
	wire [3-1:0] node671;
	wire [3-1:0] node672;
	wire [3-1:0] node674;
	wire [3-1:0] node678;
	wire [3-1:0] node679;
	wire [3-1:0] node680;
	wire [3-1:0] node682;
	wire [3-1:0] node686;
	wire [3-1:0] node689;
	wire [3-1:0] node690;
	wire [3-1:0] node691;
	wire [3-1:0] node692;
	wire [3-1:0] node695;
	wire [3-1:0] node698;
	wire [3-1:0] node699;
	wire [3-1:0] node702;
	wire [3-1:0] node705;
	wire [3-1:0] node706;
	wire [3-1:0] node709;
	wire [3-1:0] node712;
	wire [3-1:0] node713;
	wire [3-1:0] node714;
	wire [3-1:0] node715;
	wire [3-1:0] node716;
	wire [3-1:0] node718;
	wire [3-1:0] node724;
	wire [3-1:0] node725;
	wire [3-1:0] node726;
	wire [3-1:0] node727;
	wire [3-1:0] node729;
	wire [3-1:0] node733;
	wire [3-1:0] node736;
	wire [3-1:0] node737;
	wire [3-1:0] node741;
	wire [3-1:0] node742;
	wire [3-1:0] node743;
	wire [3-1:0] node744;
	wire [3-1:0] node746;
	wire [3-1:0] node749;
	wire [3-1:0] node750;
	wire [3-1:0] node753;
	wire [3-1:0] node756;
	wire [3-1:0] node757;
	wire [3-1:0] node758;
	wire [3-1:0] node759;
	wire [3-1:0] node761;
	wire [3-1:0] node764;
	wire [3-1:0] node767;
	wire [3-1:0] node770;
	wire [3-1:0] node771;
	wire [3-1:0] node772;
	wire [3-1:0] node776;
	wire [3-1:0] node779;
	wire [3-1:0] node780;
	wire [3-1:0] node781;
	wire [3-1:0] node782;
	wire [3-1:0] node784;
	wire [3-1:0] node785;
	wire [3-1:0] node789;
	wire [3-1:0] node791;
	wire [3-1:0] node792;
	wire [3-1:0] node796;
	wire [3-1:0] node797;
	wire [3-1:0] node799;
	wire [3-1:0] node802;
	wire [3-1:0] node805;
	wire [3-1:0] node806;
	wire [3-1:0] node807;
	wire [3-1:0] node809;
	wire [3-1:0] node810;
	wire [3-1:0] node813;
	wire [3-1:0] node816;
	wire [3-1:0] node819;
	wire [3-1:0] node820;
	wire [3-1:0] node821;
	wire [3-1:0] node823;
	wire [3-1:0] node827;
	wire [3-1:0] node830;
	wire [3-1:0] node831;
	wire [3-1:0] node832;
	wire [3-1:0] node833;
	wire [3-1:0] node835;
	wire [3-1:0] node836;
	wire [3-1:0] node837;
	wire [3-1:0] node839;
	wire [3-1:0] node843;
	wire [3-1:0] node844;
	wire [3-1:0] node850;
	wire [3-1:0] node851;
	wire [3-1:0] node852;
	wire [3-1:0] node853;
	wire [3-1:0] node854;
	wire [3-1:0] node855;
	wire [3-1:0] node856;
	wire [3-1:0] node860;
	wire [3-1:0] node863;
	wire [3-1:0] node864;
	wire [3-1:0] node866;
	wire [3-1:0] node870;
	wire [3-1:0] node871;
	wire [3-1:0] node872;
	wire [3-1:0] node876;
	wire [3-1:0] node877;
	wire [3-1:0] node881;
	wire [3-1:0] node882;
	wire [3-1:0] node883;
	wire [3-1:0] node885;
	wire [3-1:0] node886;
	wire [3-1:0] node891;
	wire [3-1:0] node892;
	wire [3-1:0] node895;
	wire [3-1:0] node896;
	wire [3-1:0] node898;
	wire [3-1:0] node901;
	wire [3-1:0] node903;
	wire [3-1:0] node906;
	wire [3-1:0] node907;
	wire [3-1:0] node908;
	wire [3-1:0] node909;
	wire [3-1:0] node910;
	wire [3-1:0] node914;
	wire [3-1:0] node916;
	wire [3-1:0] node919;
	wire [3-1:0] node920;
	wire [3-1:0] node922;

	assign outp = (inp[6]) ? node302 : node1;
		assign node1 = (inp[9]) ? node271 : node2;
			assign node2 = (inp[0]) ? node198 : node3;
				assign node3 = (inp[7]) ? node81 : node4;
					assign node4 = (inp[10]) ? node60 : node5;
						assign node5 = (inp[1]) ? node35 : node6;
							assign node6 = (inp[8]) ? node22 : node7;
								assign node7 = (inp[11]) ? node13 : node8;
									assign node8 = (inp[5]) ? node10 : 3'b010;
										assign node10 = (inp[3]) ? 3'b100 : 3'b010;
									assign node13 = (inp[3]) ? node19 : node14;
										assign node14 = (inp[4]) ? 3'b100 : node15;
											assign node15 = (inp[5]) ? 3'b100 : 3'b000;
										assign node19 = (inp[2]) ? 3'b000 : 3'b100;
								assign node22 = (inp[11]) ? node28 : node23;
									assign node23 = (inp[3]) ? node25 : 3'b110;
										assign node25 = (inp[2]) ? 3'b010 : 3'b110;
									assign node28 = (inp[3]) ? 3'b010 : node29;
										assign node29 = (inp[4]) ? 3'b010 : node30;
											assign node30 = (inp[5]) ? 3'b010 : 3'b110;
							assign node35 = (inp[3]) ? node49 : node36;
								assign node36 = (inp[8]) ? node44 : node37;
									assign node37 = (inp[11]) ? 3'b000 : node38;
										assign node38 = (inp[2]) ? node40 : 3'b100;
											assign node40 = (inp[4]) ? 3'b000 : 3'b100;
									assign node44 = (inp[11]) ? node46 : 3'b010;
										assign node46 = (inp[4]) ? 3'b000 : 3'b100;
								assign node49 = (inp[8]) ? node55 : node50;
									assign node50 = (inp[2]) ? 3'b000 : node51;
										assign node51 = (inp[11]) ? 3'b000 : 3'b100;
									assign node55 = (inp[2]) ? node57 : 3'b100;
										assign node57 = (inp[11]) ? 3'b000 : 3'b100;
						assign node60 = (inp[1]) ? 3'b000 : node61;
							assign node61 = (inp[8]) ? node71 : node62;
								assign node62 = (inp[3]) ? 3'b000 : node63;
									assign node63 = (inp[2]) ? 3'b000 : node64;
										assign node64 = (inp[5]) ? 3'b000 : node65;
											assign node65 = (inp[11]) ? 3'b000 : 3'b100;
								assign node71 = (inp[11]) ? 3'b000 : node72;
									assign node72 = (inp[4]) ? node74 : 3'b100;
										assign node74 = (inp[5]) ? node76 : 3'b100;
											assign node76 = (inp[3]) ? 3'b000 : 3'b100;
					assign node81 = (inp[10]) ? node145 : node82;
						assign node82 = (inp[1]) ? node120 : node83;
							assign node83 = (inp[8]) ? node99 : node84;
								assign node84 = (inp[11]) ? node92 : node85;
									assign node85 = (inp[3]) ? node87 : 3'b001;
										assign node87 = (inp[5]) ? node89 : 3'b001;
											assign node89 = (inp[2]) ? 3'b110 : 3'b001;
									assign node92 = (inp[2]) ? node96 : node93;
										assign node93 = (inp[3]) ? 3'b110 : 3'b001;
										assign node96 = (inp[4]) ? 3'b010 : 3'b110;
								assign node99 = (inp[11]) ? node111 : node100;
									assign node100 = (inp[2]) ? node106 : node101;
										assign node101 = (inp[4]) ? node103 : 3'b011;
											assign node103 = (inp[5]) ? 3'b101 : 3'b001;
										assign node106 = (inp[3]) ? node108 : 3'b101;
											assign node108 = (inp[4]) ? 3'b001 : 3'b101;
									assign node111 = (inp[2]) ? node115 : node112;
										assign node112 = (inp[3]) ? 3'b001 : 3'b101;
										assign node115 = (inp[3]) ? node117 : 3'b001;
											assign node117 = (inp[5]) ? 3'b110 : 3'b001;
							assign node120 = (inp[8]) ? node134 : node121;
								assign node121 = (inp[11]) ? node129 : node122;
									assign node122 = (inp[2]) ? node124 : 3'b110;
										assign node124 = (inp[3]) ? 3'b010 : node125;
											assign node125 = (inp[4]) ? 3'b010 : 3'b110;
									assign node129 = (inp[2]) ? node131 : 3'b010;
										assign node131 = (inp[3]) ? 3'b100 : 3'b010;
								assign node134 = (inp[3]) ? node140 : node135;
									assign node135 = (inp[11]) ? node137 : 3'b001;
										assign node137 = (inp[5]) ? 3'b110 : 3'b001;
									assign node140 = (inp[11]) ? node142 : 3'b110;
										assign node142 = (inp[2]) ? 3'b010 : 3'b110;
						assign node145 = (inp[1]) ? node173 : node146;
							assign node146 = (inp[8]) ? node164 : node147;
								assign node147 = (inp[11]) ? node157 : node148;
									assign node148 = (inp[4]) ? node154 : node149;
										assign node149 = (inp[2]) ? 3'b010 : node150;
											assign node150 = (inp[3]) ? 3'b010 : 3'b110;
										assign node154 = (inp[5]) ? 3'b100 : 3'b010;
									assign node157 = (inp[5]) ? node159 : 3'b100;
										assign node159 = (inp[4]) ? node161 : 3'b010;
											assign node161 = (inp[2]) ? 3'b100 : 3'b000;
								assign node164 = (inp[2]) ? node170 : node165;
									assign node165 = (inp[3]) ? 3'b110 : node166;
										assign node166 = (inp[11]) ? 3'b110 : 3'b001;
									assign node170 = (inp[11]) ? 3'b010 : 3'b110;
							assign node173 = (inp[8]) ? node181 : node174;
								assign node174 = (inp[11]) ? 3'b000 : node175;
									assign node175 = (inp[2]) ? node177 : 3'b100;
										assign node177 = (inp[3]) ? 3'b000 : 3'b100;
								assign node181 = (inp[11]) ? node191 : node182;
									assign node182 = (inp[2]) ? node188 : node183;
										assign node183 = (inp[3]) ? 3'b010 : node184;
											assign node184 = (inp[4]) ? 3'b010 : 3'b010;
										assign node188 = (inp[3]) ? 3'b100 : 3'b010;
									assign node191 = (inp[4]) ? node193 : 3'b010;
										assign node193 = (inp[2]) ? node195 : 3'b100;
											assign node195 = (inp[3]) ? 3'b000 : 3'b100;
				assign node198 = (inp[7]) ? node210 : node199;
					assign node199 = (inp[2]) ? 3'b000 : node200;
						assign node200 = (inp[8]) ? node202 : 3'b000;
							assign node202 = (inp[4]) ? 3'b000 : node203;
								assign node203 = (inp[1]) ? 3'b000 : node204;
									assign node204 = (inp[3]) ? 3'b000 : 3'b100;
					assign node210 = (inp[10]) ? node258 : node211;
						assign node211 = (inp[1]) ? node239 : node212;
							assign node212 = (inp[8]) ? node228 : node213;
								assign node213 = (inp[2]) ? node221 : node214;
									assign node214 = (inp[11]) ? 3'b100 : node215;
										assign node215 = (inp[4]) ? node217 : 3'b010;
											assign node217 = (inp[3]) ? 3'b100 : 3'b010;
									assign node221 = (inp[11]) ? node223 : 3'b100;
										assign node223 = (inp[5]) ? 3'b000 : node224;
											assign node224 = (inp[4]) ? 3'b000 : 3'b000;
								assign node228 = (inp[11]) ? node234 : node229;
									assign node229 = (inp[4]) ? node231 : 3'b110;
										assign node231 = (inp[2]) ? 3'b010 : 3'b110;
									assign node234 = (inp[4]) ? node236 : 3'b010;
										assign node236 = (inp[5]) ? 3'b010 : 3'b100;
							assign node239 = (inp[11]) ? node251 : node240;
								assign node240 = (inp[8]) ? node246 : node241;
									assign node241 = (inp[2]) ? 3'b000 : node242;
										assign node242 = (inp[3]) ? 3'b000 : 3'b100;
									assign node246 = (inp[2]) ? 3'b100 : node247;
										assign node247 = (inp[4]) ? 3'b100 : 3'b010;
								assign node251 = (inp[2]) ? 3'b000 : node252;
									assign node252 = (inp[3]) ? 3'b000 : node253;
										assign node253 = (inp[8]) ? 3'b100 : 3'b000;
						assign node258 = (inp[11]) ? 3'b000 : node259;
							assign node259 = (inp[8]) ? node261 : 3'b000;
								assign node261 = (inp[1]) ? 3'b000 : node262;
									assign node262 = (inp[2]) ? node264 : 3'b100;
										assign node264 = (inp[3]) ? 3'b000 : node265;
											assign node265 = (inp[5]) ? 3'b000 : 3'b100;
			assign node271 = (inp[7]) ? node273 : 3'b000;
				assign node273 = (inp[0]) ? 3'b000 : node274;
					assign node274 = (inp[10]) ? 3'b000 : node275;
						assign node275 = (inp[1]) ? node293 : node276;
							assign node276 = (inp[8]) ? node282 : node277;
								assign node277 = (inp[3]) ? 3'b000 : node278;
									assign node278 = (inp[11]) ? 3'b000 : 3'b100;
								assign node282 = (inp[11]) ? node288 : node283;
									assign node283 = (inp[2]) ? 3'b100 : node284;
										assign node284 = (inp[5]) ? 3'b100 : 3'b010;
									assign node288 = (inp[3]) ? 3'b000 : node289;
										assign node289 = (inp[2]) ? 3'b000 : 3'b100;
							assign node293 = (inp[11]) ? 3'b000 : node294;
								assign node294 = (inp[3]) ? 3'b000 : node295;
									assign node295 = (inp[4]) ? 3'b000 : 3'b100;
		assign node302 = (inp[9]) ? node658 : node303;
			assign node303 = (inp[0]) ? node455 : node304;
				assign node304 = (inp[7]) ? node408 : node305;
					assign node305 = (inp[10]) ? node355 : node306;
						assign node306 = (inp[1]) ? node324 : node307;
							assign node307 = (inp[8]) ? node317 : node308;
								assign node308 = (inp[11]) ? node314 : node309;
									assign node309 = (inp[2]) ? 3'b011 : node310;
										assign node310 = (inp[3]) ? 3'b011 : 3'b111;
									assign node314 = (inp[3]) ? 3'b101 : 3'b011;
								assign node317 = (inp[11]) ? node319 : 3'b111;
									assign node319 = (inp[2]) ? 3'b011 : node320;
										assign node320 = (inp[3]) ? 3'b011 : 3'b111;
							assign node324 = (inp[8]) ? node344 : node325;
								assign node325 = (inp[11]) ? node335 : node326;
									assign node326 = (inp[5]) ? 3'b101 : node327;
										assign node327 = (inp[4]) ? node331 : node328;
											assign node328 = (inp[2]) ? 3'b101 : 3'b011;
											assign node331 = (inp[3]) ? 3'b001 : 3'b101;
									assign node335 = (inp[3]) ? node341 : node336;
										assign node336 = (inp[5]) ? node338 : 3'b001;
											assign node338 = (inp[4]) ? 3'b001 : 3'b101;
										assign node341 = (inp[4]) ? 3'b110 : 3'b001;
								assign node344 = (inp[11]) ? node346 : 3'b011;
									assign node346 = (inp[2]) ? node350 : node347;
										assign node347 = (inp[3]) ? 3'b101 : 3'b011;
										assign node350 = (inp[3]) ? node352 : 3'b101;
											assign node352 = (inp[4]) ? 3'b001 : 3'b101;
						assign node355 = (inp[8]) ? node379 : node356;
							assign node356 = (inp[1]) ? node366 : node357;
								assign node357 = (inp[11]) ? node363 : node358;
									assign node358 = (inp[2]) ? 3'b001 : node359;
										assign node359 = (inp[3]) ? 3'b001 : 3'b101;
									assign node363 = (inp[2]) ? 3'b110 : 3'b001;
								assign node366 = (inp[11]) ? node372 : node367;
									assign node367 = (inp[4]) ? 3'b110 : node368;
										assign node368 = (inp[3]) ? 3'b110 : 3'b001;
									assign node372 = (inp[4]) ? node374 : 3'b010;
										assign node374 = (inp[3]) ? 3'b100 : node375;
											assign node375 = (inp[5]) ? 3'b010 : 3'b110;
							assign node379 = (inp[2]) ? node397 : node380;
								assign node380 = (inp[1]) ? node392 : node381;
									assign node381 = (inp[11]) ? node387 : node382;
										assign node382 = (inp[4]) ? node384 : 3'b011;
											assign node384 = (inp[3]) ? 3'b101 : 3'b011;
										assign node387 = (inp[4]) ? node389 : 3'b101;
											assign node389 = (inp[3]) ? 3'b001 : 3'b101;
									assign node392 = (inp[3]) ? 3'b001 : node393;
										assign node393 = (inp[11]) ? 3'b001 : 3'b101;
								assign node397 = (inp[1]) ? node401 : node398;
									assign node398 = (inp[11]) ? 3'b001 : 3'b101;
									assign node401 = (inp[11]) ? 3'b110 : node402;
										assign node402 = (inp[5]) ? node404 : 3'b001;
											assign node404 = (inp[3]) ? 3'b000 : 3'b001;
					assign node408 = (inp[10]) ? node416 : node409;
						assign node409 = (inp[8]) ? 3'b111 : node410;
							assign node410 = (inp[1]) ? node412 : 3'b111;
								assign node412 = (inp[11]) ? 3'b011 : 3'b111;
						assign node416 = (inp[1]) ? node434 : node417;
							assign node417 = (inp[2]) ? node423 : node418;
								assign node418 = (inp[11]) ? node420 : 3'b111;
									assign node420 = (inp[8]) ? 3'b111 : 3'b011;
								assign node423 = (inp[11]) ? node427 : node424;
									assign node424 = (inp[8]) ? 3'b111 : 3'b011;
									assign node427 = (inp[8]) ? 3'b011 : node428;
										assign node428 = (inp[4]) ? 3'b101 : node429;
											assign node429 = (inp[3]) ? 3'b101 : 3'b011;
							assign node434 = (inp[8]) ? node446 : node435;
								assign node435 = (inp[11]) ? node441 : node436;
									assign node436 = (inp[2]) ? 3'b101 : node437;
										assign node437 = (inp[3]) ? 3'b101 : 3'b011;
									assign node441 = (inp[2]) ? 3'b001 : node442;
										assign node442 = (inp[3]) ? 3'b001 : 3'b101;
								assign node446 = (inp[11]) ? node452 : node447;
									assign node447 = (inp[2]) ? 3'b011 : node448;
										assign node448 = (inp[3]) ? 3'b011 : 3'b111;
									assign node452 = (inp[2]) ? 3'b101 : 3'b011;
				assign node455 = (inp[7]) ? node549 : node456;
					assign node456 = (inp[10]) ? node506 : node457;
						assign node457 = (inp[2]) ? node481 : node458;
							assign node458 = (inp[1]) ? node466 : node459;
								assign node459 = (inp[11]) ? node463 : node460;
									assign node460 = (inp[8]) ? 3'b101 : 3'b001;
									assign node463 = (inp[8]) ? 3'b001 : 3'b110;
								assign node466 = (inp[8]) ? node474 : node467;
									assign node467 = (inp[3]) ? node469 : 3'b110;
										assign node469 = (inp[5]) ? node471 : 3'b010;
											assign node471 = (inp[4]) ? 3'b000 : 3'b010;
									assign node474 = (inp[11]) ? 3'b110 : node475;
										assign node475 = (inp[4]) ? node477 : 3'b001;
											assign node477 = (inp[5]) ? 3'b110 : 3'b001;
							assign node481 = (inp[8]) ? node497 : node482;
								assign node482 = (inp[1]) ? node494 : node483;
									assign node483 = (inp[11]) ? node489 : node484;
										assign node484 = (inp[5]) ? 3'b110 : node485;
											assign node485 = (inp[4]) ? 3'b110 : 3'b001;
										assign node489 = (inp[5]) ? 3'b010 : node490;
											assign node490 = (inp[4]) ? 3'b110 : 3'b010;
									assign node494 = (inp[11]) ? 3'b100 : 3'b010;
								assign node497 = (inp[4]) ? 3'b110 : node498;
									assign node498 = (inp[5]) ? node502 : node499;
										assign node499 = (inp[11]) ? 3'b110 : 3'b001;
										assign node502 = (inp[11]) ? 3'b010 : 3'b110;
						assign node506 = (inp[1]) ? node528 : node507;
							assign node507 = (inp[11]) ? node515 : node508;
								assign node508 = (inp[8]) ? 3'b110 : node509;
									assign node509 = (inp[5]) ? node511 : 3'b010;
										assign node511 = (inp[2]) ? 3'b100 : 3'b010;
								assign node515 = (inp[8]) ? node521 : node516;
									assign node516 = (inp[3]) ? node518 : 3'b100;
										assign node518 = (inp[2]) ? 3'b000 : 3'b100;
									assign node521 = (inp[4]) ? 3'b010 : node522;
										assign node522 = (inp[2]) ? node524 : 3'b010;
											assign node524 = (inp[3]) ? 3'b100 : 3'b010;
							assign node528 = (inp[8]) ? node538 : node529;
								assign node529 = (inp[11]) ? 3'b000 : node530;
									assign node530 = (inp[2]) ? 3'b000 : node531;
										assign node531 = (inp[5]) ? node533 : 3'b100;
											assign node533 = (inp[4]) ? 3'b000 : 3'b100;
								assign node538 = (inp[11]) ? node546 : node539;
									assign node539 = (inp[2]) ? node541 : 3'b010;
										assign node541 = (inp[3]) ? 3'b100 : node542;
											assign node542 = (inp[5]) ? 3'b100 : 3'b010;
									assign node546 = (inp[2]) ? 3'b000 : 3'b100;
					assign node549 = (inp[10]) ? node605 : node550;
						assign node550 = (inp[1]) ? node580 : node551;
							assign node551 = (inp[8]) ? node565 : node552;
								assign node552 = (inp[11]) ? node560 : node553;
									assign node553 = (inp[3]) ? node557 : node554;
										assign node554 = (inp[2]) ? 3'b011 : 3'b111;
										assign node557 = (inp[2]) ? 3'b101 : 3'b011;
									assign node560 = (inp[3]) ? node562 : 3'b101;
										assign node562 = (inp[2]) ? 3'b001 : 3'b101;
								assign node565 = (inp[11]) ? node573 : node566;
									assign node566 = (inp[3]) ? node568 : 3'b111;
										assign node568 = (inp[5]) ? node570 : 3'b111;
											assign node570 = (inp[2]) ? 3'b011 : 3'b111;
									assign node573 = (inp[5]) ? node575 : 3'b011;
										assign node575 = (inp[4]) ? node577 : 3'b111;
											assign node577 = (inp[2]) ? 3'b001 : 3'b011;
							assign node580 = (inp[11]) ? node594 : node581;
								assign node581 = (inp[8]) ? node589 : node582;
									assign node582 = (inp[2]) ? node584 : 3'b101;
										assign node584 = (inp[3]) ? 3'b001 : node585;
											assign node585 = (inp[4]) ? 3'b001 : 3'b101;
									assign node589 = (inp[2]) ? node591 : 3'b011;
										assign node591 = (inp[4]) ? 3'b101 : 3'b011;
								assign node594 = (inp[8]) ? node598 : node595;
									assign node595 = (inp[2]) ? 3'b110 : 3'b001;
									assign node598 = (inp[4]) ? node600 : 3'b101;
										assign node600 = (inp[2]) ? node602 : 3'b101;
											assign node602 = (inp[3]) ? 3'b001 : 3'b101;
						assign node605 = (inp[1]) ? node639 : node606;
							assign node606 = (inp[2]) ? node620 : node607;
								assign node607 = (inp[11]) ? node615 : node608;
									assign node608 = (inp[8]) ? node610 : 3'b001;
										assign node610 = (inp[3]) ? 3'b101 : node611;
											assign node611 = (inp[4]) ? 3'b101 : 3'b011;
									assign node615 = (inp[8]) ? node617 : 3'b110;
										assign node617 = (inp[4]) ? 3'b001 : 3'b101;
								assign node620 = (inp[8]) ? node632 : node621;
									assign node621 = (inp[11]) ? node627 : node622;
										assign node622 = (inp[3]) ? node624 : 3'b001;
											assign node624 = (inp[5]) ? 3'b110 : 3'b001;
										assign node627 = (inp[3]) ? node629 : 3'b110;
											assign node629 = (inp[5]) ? 3'b010 : 3'b010;
									assign node632 = (inp[3]) ? node636 : node633;
										assign node633 = (inp[11]) ? 3'b001 : 3'b101;
										assign node636 = (inp[4]) ? 3'b110 : 3'b001;
							assign node639 = (inp[2]) ? node647 : node640;
								assign node640 = (inp[11]) ? node644 : node641;
									assign node641 = (inp[8]) ? 3'b001 : 3'b110;
									assign node644 = (inp[8]) ? 3'b110 : 3'b010;
								assign node647 = (inp[11]) ? node653 : node648;
									assign node648 = (inp[8]) ? node650 : 3'b010;
										assign node650 = (inp[3]) ? 3'b110 : 3'b001;
									assign node653 = (inp[8]) ? node655 : 3'b100;
										assign node655 = (inp[3]) ? 3'b010 : 3'b110;
			assign node658 = (inp[0]) ? node830 : node659;
				assign node659 = (inp[7]) ? node741 : node660;
					assign node660 = (inp[10]) ? node712 : node661;
						assign node661 = (inp[1]) ? node689 : node662;
							assign node662 = (inp[11]) ? node678 : node663;
								assign node663 = (inp[8]) ? node671 : node664;
									assign node664 = (inp[2]) ? 3'b010 : node665;
										assign node665 = (inp[4]) ? node667 : 3'b110;
											assign node667 = (inp[3]) ? 3'b010 : 3'b110;
									assign node671 = (inp[2]) ? 3'b110 : node672;
										assign node672 = (inp[3]) ? node674 : 3'b001;
											assign node674 = (inp[5]) ? 3'b000 : 3'b001;
								assign node678 = (inp[2]) ? node686 : node679;
									assign node679 = (inp[8]) ? 3'b110 : node680;
										assign node680 = (inp[3]) ? node682 : 3'b010;
											assign node682 = (inp[4]) ? 3'b100 : 3'b010;
									assign node686 = (inp[8]) ? 3'b010 : 3'b100;
							assign node689 = (inp[3]) ? node705 : node690;
								assign node690 = (inp[8]) ? node698 : node691;
									assign node691 = (inp[2]) ? node695 : node692;
										assign node692 = (inp[11]) ? 3'b100 : 3'b010;
										assign node695 = (inp[11]) ? 3'b000 : 3'b100;
									assign node698 = (inp[11]) ? node702 : node699;
										assign node699 = (inp[2]) ? 3'b010 : 3'b110;
										assign node702 = (inp[2]) ? 3'b100 : 3'b010;
								assign node705 = (inp[11]) ? node709 : node706;
									assign node706 = (inp[8]) ? 3'b010 : 3'b100;
									assign node709 = (inp[8]) ? 3'b100 : 3'b000;
						assign node712 = (inp[8]) ? node724 : node713;
							assign node713 = (inp[11]) ? 3'b000 : node714;
								assign node714 = (inp[1]) ? 3'b000 : node715;
									assign node715 = (inp[2]) ? 3'b000 : node716;
										assign node716 = (inp[3]) ? node718 : 3'b100;
											assign node718 = (inp[5]) ? 3'b000 : 3'b100;
							assign node724 = (inp[1]) ? node736 : node725;
								assign node725 = (inp[2]) ? node733 : node726;
									assign node726 = (inp[11]) ? 3'b100 : node727;
										assign node727 = (inp[4]) ? node729 : 3'b010;
											assign node729 = (inp[5]) ? 3'b100 : 3'b010;
									assign node733 = (inp[11]) ? 3'b000 : 3'b100;
								assign node736 = (inp[2]) ? 3'b000 : node737;
									assign node737 = (inp[11]) ? 3'b000 : 3'b100;
					assign node741 = (inp[10]) ? node779 : node742;
						assign node742 = (inp[1]) ? node756 : node743;
							assign node743 = (inp[8]) ? node749 : node744;
								assign node744 = (inp[11]) ? node746 : 3'b001;
									assign node746 = (inp[2]) ? 3'b110 : 3'b001;
								assign node749 = (inp[11]) ? node753 : node750;
									assign node750 = (inp[2]) ? 3'b101 : 3'b011;
									assign node753 = (inp[2]) ? 3'b001 : 3'b101;
							assign node756 = (inp[8]) ? node770 : node757;
								assign node757 = (inp[2]) ? node767 : node758;
									assign node758 = (inp[11]) ? node764 : node759;
										assign node759 = (inp[5]) ? node761 : 3'b001;
											assign node761 = (inp[3]) ? 3'b110 : 3'b001;
										assign node764 = (inp[3]) ? 3'b010 : 3'b110;
									assign node767 = (inp[11]) ? 3'b010 : 3'b110;
								assign node770 = (inp[2]) ? node776 : node771;
									assign node771 = (inp[11]) ? 3'b001 : node772;
										assign node772 = (inp[3]) ? 3'b001 : 3'b101;
									assign node776 = (inp[11]) ? 3'b110 : 3'b001;
						assign node779 = (inp[1]) ? node805 : node780;
							assign node780 = (inp[8]) ? node796 : node781;
								assign node781 = (inp[11]) ? node789 : node782;
									assign node782 = (inp[2]) ? node784 : 3'b110;
										assign node784 = (inp[4]) ? 3'b010 : node785;
											assign node785 = (inp[3]) ? 3'b010 : 3'b110;
									assign node789 = (inp[2]) ? node791 : 3'b010;
										assign node791 = (inp[4]) ? 3'b100 : node792;
											assign node792 = (inp[3]) ? 3'b100 : 3'b010;
								assign node796 = (inp[11]) ? node802 : node797;
									assign node797 = (inp[2]) ? node799 : 3'b001;
										assign node799 = (inp[3]) ? 3'b110 : 3'b001;
									assign node802 = (inp[3]) ? 3'b010 : 3'b110;
							assign node805 = (inp[8]) ? node819 : node806;
								assign node806 = (inp[2]) ? node816 : node807;
									assign node807 = (inp[3]) ? node809 : 3'b100;
										assign node809 = (inp[4]) ? node813 : node810;
											assign node810 = (inp[11]) ? 3'b100 : 3'b010;
											assign node813 = (inp[11]) ? 3'b000 : 3'b100;
									assign node816 = (inp[11]) ? 3'b000 : 3'b100;
								assign node819 = (inp[11]) ? node827 : node820;
									assign node820 = (inp[2]) ? 3'b010 : node821;
										assign node821 = (inp[4]) ? node823 : 3'b110;
											assign node823 = (inp[3]) ? 3'b010 : 3'b110;
									assign node827 = (inp[2]) ? 3'b100 : 3'b010;
				assign node830 = (inp[7]) ? node850 : node831;
					assign node831 = (inp[10]) ? 3'b000 : node832;
						assign node832 = (inp[1]) ? 3'b000 : node833;
							assign node833 = (inp[8]) ? node835 : 3'b000;
								assign node835 = (inp[11]) ? node843 : node836;
									assign node836 = (inp[5]) ? 3'b100 : node837;
										assign node837 = (inp[3]) ? node839 : 3'b010;
											assign node839 = (inp[4]) ? 3'b000 : 3'b100;
									assign node843 = (inp[2]) ? 3'b000 : node844;
										assign node844 = (inp[4]) ? 3'b000 : 3'b100;
					assign node850 = (inp[10]) ? node906 : node851;
						assign node851 = (inp[1]) ? node881 : node852;
							assign node852 = (inp[8]) ? node870 : node853;
								assign node853 = (inp[11]) ? node863 : node854;
									assign node854 = (inp[2]) ? node860 : node855;
										assign node855 = (inp[4]) ? 3'b010 : node856;
											assign node856 = (inp[3]) ? 3'b010 : 3'b110;
										assign node860 = (inp[4]) ? 3'b100 : 3'b010;
									assign node863 = (inp[5]) ? 3'b100 : node864;
										assign node864 = (inp[3]) ? node866 : 3'b010;
											assign node866 = (inp[2]) ? 3'b000 : 3'b100;
								assign node870 = (inp[11]) ? node876 : node871;
									assign node871 = (inp[2]) ? 3'b110 : node872;
										assign node872 = (inp[3]) ? 3'b110 : 3'b001;
									assign node876 = (inp[3]) ? 3'b010 : node877;
										assign node877 = (inp[2]) ? 3'b010 : 3'b110;
							assign node881 = (inp[8]) ? node891 : node882;
								assign node882 = (inp[11]) ? 3'b000 : node883;
									assign node883 = (inp[2]) ? node885 : 3'b100;
										assign node885 = (inp[3]) ? 3'b000 : node886;
											assign node886 = (inp[5]) ? 3'b000 : 3'b100;
								assign node891 = (inp[11]) ? node895 : node892;
									assign node892 = (inp[3]) ? 3'b100 : 3'b010;
									assign node895 = (inp[4]) ? node901 : node896;
										assign node896 = (inp[5]) ? node898 : 3'b010;
											assign node898 = (inp[2]) ? 3'b000 : 3'b100;
										assign node901 = (inp[3]) ? node903 : 3'b100;
											assign node903 = (inp[2]) ? 3'b000 : 3'b100;
						assign node906 = (inp[1]) ? 3'b000 : node907;
							assign node907 = (inp[11]) ? node919 : node908;
								assign node908 = (inp[8]) ? node914 : node909;
									assign node909 = (inp[5]) ? 3'b000 : node910;
										assign node910 = (inp[2]) ? 3'b000 : 3'b100;
									assign node914 = (inp[4]) ? node916 : 3'b100;
										assign node916 = (inp[2]) ? 3'b100 : 3'b010;
								assign node919 = (inp[2]) ? 3'b000 : node920;
									assign node920 = (inp[5]) ? node922 : 3'b000;
										assign node922 = (inp[8]) ? 3'b100 : 3'b000;

endmodule