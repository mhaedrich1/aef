module dtc_split875_bm53 (
	input  wire [8-1:0] inp,
	output wire [2-1:0] outp
);

	wire [2-1:0] node1;
	wire [2-1:0] node2;
	wire [2-1:0] node3;
	wire [2-1:0] node4;
	wire [2-1:0] node5;
	wire [2-1:0] node7;
	wire [2-1:0] node10;
	wire [2-1:0] node12;
	wire [2-1:0] node15;
	wire [2-1:0] node17;
	wire [2-1:0] node18;
	wire [2-1:0] node21;
	wire [2-1:0] node25;
	wire [2-1:0] node26;
	wire [2-1:0] node27;
	wire [2-1:0] node28;
	wire [2-1:0] node30;
	wire [2-1:0] node33;
	wire [2-1:0] node34;
	wire [2-1:0] node38;
	wire [2-1:0] node39;
	wire [2-1:0] node40;
	wire [2-1:0] node43;
	wire [2-1:0] node47;
	wire [2-1:0] node48;
	wire [2-1:0] node49;
	wire [2-1:0] node50;
	wire [2-1:0] node56;
	wire [2-1:0] node57;
	wire [2-1:0] node58;
	wire [2-1:0] node59;
	wire [2-1:0] node61;
	wire [2-1:0] node62;
	wire [2-1:0] node66;
	wire [2-1:0] node67;
	wire [2-1:0] node68;
	wire [2-1:0] node71;
	wire [2-1:0] node74;
	wire [2-1:0] node76;
	wire [2-1:0] node79;
	wire [2-1:0] node80;
	wire [2-1:0] node81;
	wire [2-1:0] node82;
	wire [2-1:0] node86;
	wire [2-1:0] node88;
	wire [2-1:0] node91;
	wire [2-1:0] node93;
	wire [2-1:0] node94;

	assign outp = (inp[6]) ? node56 : node1;
		assign node1 = (inp[7]) ? node25 : node2;
			assign node2 = (inp[3]) ? 2'b01 : node3;
				assign node3 = (inp[0]) ? node15 : node4;
					assign node4 = (inp[2]) ? node10 : node5;
						assign node5 = (inp[4]) ? node7 : 2'b00;
							assign node7 = (inp[5]) ? 2'b00 : 2'b01;
						assign node10 = (inp[4]) ? node12 : 2'b01;
							assign node12 = (inp[5]) ? 2'b01 : 2'b00;
					assign node15 = (inp[1]) ? node17 : 2'b11;
						assign node17 = (inp[2]) ? node21 : node18;
							assign node18 = (inp[4]) ? 2'b00 : 2'b00;
							assign node21 = (inp[4]) ? 2'b00 : 2'b01;
			assign node25 = (inp[1]) ? node47 : node26;
				assign node26 = (inp[3]) ? node38 : node27;
					assign node27 = (inp[5]) ? node33 : node28;
						assign node28 = (inp[4]) ? node30 : 2'b00;
							assign node30 = (inp[2]) ? 2'b00 : 2'b00;
						assign node33 = (inp[2]) ? 2'b01 : node34;
							assign node34 = (inp[0]) ? 2'b00 : 2'b01;
					assign node38 = (inp[0]) ? 2'b01 : node39;
						assign node39 = (inp[2]) ? node43 : node40;
							assign node40 = (inp[5]) ? 2'b00 : 2'b00;
							assign node43 = (inp[5]) ? 2'b01 : 2'b00;
				assign node47 = (inp[5]) ? 2'b00 : node48;
					assign node48 = (inp[2]) ? 2'b00 : node49;
						assign node49 = (inp[3]) ? 2'b00 : node50;
							assign node50 = (inp[4]) ? 2'b00 : 2'b00;
		assign node56 = (inp[3]) ? 2'b00 : node57;
			assign node57 = (inp[7]) ? node79 : node58;
				assign node58 = (inp[1]) ? node66 : node59;
					assign node59 = (inp[2]) ? node61 : 2'b10;
						assign node61 = (inp[0]) ? 2'b10 : node62;
							assign node62 = (inp[4]) ? 2'b00 : 2'b00;
					assign node66 = (inp[0]) ? node74 : node67;
						assign node67 = (inp[2]) ? node71 : node68;
							assign node68 = (inp[5]) ? 2'b01 : 2'b00;
							assign node71 = (inp[5]) ? 2'b00 : 2'b00;
						assign node74 = (inp[2]) ? node76 : 2'b10;
							assign node76 = (inp[4]) ? 2'b10 : 2'b00;
				assign node79 = (inp[1]) ? node91 : node80;
					assign node80 = (inp[5]) ? node86 : node81;
						assign node81 = (inp[2]) ? 2'b01 : node82;
							assign node82 = (inp[4]) ? 2'b00 : 2'b01;
						assign node86 = (inp[0]) ? node88 : 2'b00;
							assign node88 = (inp[2]) ? 2'b00 : 2'b01;
					assign node91 = (inp[4]) ? node93 : 2'b00;
						assign node93 = (inp[5]) ? 2'b00 : node94;
							assign node94 = (inp[0]) ? 2'b01 : 2'b00;

endmodule