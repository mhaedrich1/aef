module dtc_split875_bm32 (
	input  wire [15-1:0] inp,
	output wire [9-1:0] outp
);

	wire [9-1:0] node1;
	wire [9-1:0] node2;
	wire [9-1:0] node5;
	wire [9-1:0] node6;
	wire [9-1:0] node7;
	wire [9-1:0] node9;
	wire [9-1:0] node11;
	wire [9-1:0] node12;
	wire [9-1:0] node14;
	wire [9-1:0] node18;
	wire [9-1:0] node21;
	wire [9-1:0] node22;
	wire [9-1:0] node24;
	wire [9-1:0] node26;
	wire [9-1:0] node29;
	wire [9-1:0] node30;
	wire [9-1:0] node31;
	wire [9-1:0] node34;
	wire [9-1:0] node35;
	wire [9-1:0] node37;
	wire [9-1:0] node41;
	wire [9-1:0] node43;
	wire [9-1:0] node45;
	wire [9-1:0] node48;
	wire [9-1:0] node49;
	wire [9-1:0] node50;
	wire [9-1:0] node51;
	wire [9-1:0] node52;
	wire [9-1:0] node53;
	wire [9-1:0] node54;
	wire [9-1:0] node55;
	wire [9-1:0] node60;
	wire [9-1:0] node61;
	wire [9-1:0] node62;
	wire [9-1:0] node63;
	wire [9-1:0] node68;
	wire [9-1:0] node71;
	wire [9-1:0] node72;
	wire [9-1:0] node73;
	wire [9-1:0] node74;
	wire [9-1:0] node79;
	wire [9-1:0] node80;
	wire [9-1:0] node81;
	wire [9-1:0] node82;
	wire [9-1:0] node87;
	wire [9-1:0] node90;
	wire [9-1:0] node91;
	wire [9-1:0] node92;
	wire [9-1:0] node93;
	wire [9-1:0] node94;
	wire [9-1:0] node99;
	wire [9-1:0] node100;
	wire [9-1:0] node101;
	wire [9-1:0] node102;
	wire [9-1:0] node107;
	wire [9-1:0] node110;
	wire [9-1:0] node111;
	wire [9-1:0] node112;
	wire [9-1:0] node113;
	wire [9-1:0] node114;
	wire [9-1:0] node115;
	wire [9-1:0] node119;
	wire [9-1:0] node120;
	wire [9-1:0] node121;
	wire [9-1:0] node126;
	wire [9-1:0] node127;
	wire [9-1:0] node129;
	wire [9-1:0] node131;
	wire [9-1:0] node134;
	wire [9-1:0] node136;
	wire [9-1:0] node139;
	wire [9-1:0] node140;
	wire [9-1:0] node143;
	wire [9-1:0] node146;
	wire [9-1:0] node147;
	wire [9-1:0] node148;
	wire [9-1:0] node149;
	wire [9-1:0] node150;
	wire [9-1:0] node154;
	wire [9-1:0] node155;
	wire [9-1:0] node156;
	wire [9-1:0] node161;
	wire [9-1:0] node162;
	wire [9-1:0] node164;
	wire [9-1:0] node166;
	wire [9-1:0] node169;
	wire [9-1:0] node171;
	wire [9-1:0] node174;
	wire [9-1:0] node176;
	wire [9-1:0] node179;
	wire [9-1:0] node180;
	wire [9-1:0] node181;
	wire [9-1:0] node182;
	wire [9-1:0] node183;
	wire [9-1:0] node184;
	wire [9-1:0] node189;
	wire [9-1:0] node190;
	wire [9-1:0] node191;
	wire [9-1:0] node192;
	wire [9-1:0] node197;
	wire [9-1:0] node200;
	wire [9-1:0] node201;
	wire [9-1:0] node202;
	wire [9-1:0] node203;
	wire [9-1:0] node208;
	wire [9-1:0] node209;
	wire [9-1:0] node210;
	wire [9-1:0] node211;
	wire [9-1:0] node216;
	wire [9-1:0] node219;
	wire [9-1:0] node220;
	wire [9-1:0] node221;
	wire [9-1:0] node222;
	wire [9-1:0] node223;
	wire [9-1:0] node228;
	wire [9-1:0] node229;
	wire [9-1:0] node230;
	wire [9-1:0] node231;
	wire [9-1:0] node236;
	wire [9-1:0] node239;
	wire [9-1:0] node240;
	wire [9-1:0] node241;
	wire [9-1:0] node242;
	wire [9-1:0] node243;
	wire [9-1:0] node244;
	wire [9-1:0] node246;
	wire [9-1:0] node248;
	wire [9-1:0] node251;
	wire [9-1:0] node253;
	wire [9-1:0] node256;
	wire [9-1:0] node257;
	wire [9-1:0] node259;
	wire [9-1:0] node261;
	wire [9-1:0] node264;
	wire [9-1:0] node266;
	wire [9-1:0] node269;
	wire [9-1:0] node271;
	wire [9-1:0] node274;
	wire [9-1:0] node275;
	wire [9-1:0] node276;
	wire [9-1:0] node277;
	wire [9-1:0] node278;
	wire [9-1:0] node282;
	wire [9-1:0] node283;
	wire [9-1:0] node284;
	wire [9-1:0] node289;
	wire [9-1:0] node290;
	wire [9-1:0] node291;
	wire [9-1:0] node295;
	wire [9-1:0] node296;
	wire [9-1:0] node297;
	wire [9-1:0] node302;
	wire [9-1:0] node303;
	wire [9-1:0] node306;
	wire [9-1:0] node309;
	wire [9-1:0] node310;
	wire [9-1:0] node311;
	wire [9-1:0] node312;
	wire [9-1:0] node313;
	wire [9-1:0] node314;
	wire [9-1:0] node318;
	wire [9-1:0] node319;
	wire [9-1:0] node320;
	wire [9-1:0] node325;
	wire [9-1:0] node326;
	wire [9-1:0] node327;
	wire [9-1:0] node331;
	wire [9-1:0] node332;
	wire [9-1:0] node333;
	wire [9-1:0] node338;
	wire [9-1:0] node340;
	wire [9-1:0] node343;
	wire [9-1:0] node344;
	wire [9-1:0] node345;
	wire [9-1:0] node346;
	wire [9-1:0] node347;
	wire [9-1:0] node351;
	wire [9-1:0] node352;
	wire [9-1:0] node353;
	wire [9-1:0] node358;
	wire [9-1:0] node359;
	wire [9-1:0] node360;
	wire [9-1:0] node364;
	wire [9-1:0] node365;
	wire [9-1:0] node366;
	wire [9-1:0] node371;
	wire [9-1:0] node372;
	wire [9-1:0] node375;
	wire [9-1:0] node378;
	wire [9-1:0] node379;
	wire [9-1:0] node380;
	wire [9-1:0] node381;
	wire [9-1:0] node383;
	wire [9-1:0] node386;
	wire [9-1:0] node387;
	wire [9-1:0] node390;
	wire [9-1:0] node391;
	wire [9-1:0] node394;
	wire [9-1:0] node395;
	wire [9-1:0] node398;
	wire [9-1:0] node401;
	wire [9-1:0] node402;
	wire [9-1:0] node404;
	wire [9-1:0] node407;
	wire [9-1:0] node408;
	wire [9-1:0] node411;
	wire [9-1:0] node412;
	wire [9-1:0] node415;
	wire [9-1:0] node416;
	wire [9-1:0] node419;
	wire [9-1:0] node422;
	wire [9-1:0] node423;
	wire [9-1:0] node424;
	wire [9-1:0] node425;
	wire [9-1:0] node428;
	wire [9-1:0] node430;
	wire [9-1:0] node433;
	wire [9-1:0] node434;
	wire [9-1:0] node437;
	wire [9-1:0] node439;
	wire [9-1:0] node440;
	wire [9-1:0] node443;
	wire [9-1:0] node446;
	wire [9-1:0] node447;
	wire [9-1:0] node448;
	wire [9-1:0] node451;
	wire [9-1:0] node454;
	wire [9-1:0] node455;
	wire [9-1:0] node458;
	wire [9-1:0] node459;
	wire [9-1:0] node460;
	wire [9-1:0] node463;
	wire [9-1:0] node464;
	wire [9-1:0] node467;
	wire [9-1:0] node470;
	wire [9-1:0] node471;
	wire [9-1:0] node474;
	wire [9-1:0] node475;
	wire [9-1:0] node478;

	assign outp = (inp[12]) ? node48 : node1;
		assign node1 = (inp[13]) ? node5 : node2;
			assign node2 = (inp[11]) ? 9'b101010101 : 9'b101010000;
			assign node5 = (inp[14]) ? node21 : node6;
				assign node6 = (inp[0]) ? node18 : node7;
					assign node7 = (inp[3]) ? node9 : 9'b101010001;
						assign node9 = (inp[8]) ? node11 : 9'b100010001;
							assign node11 = (inp[4]) ? 9'b100010001 : node12;
								assign node12 = (inp[9]) ? node14 : 9'b100010001;
									assign node14 = (inp[6]) ? 9'b001010001 : 9'b101010001;
					assign node18 = (inp[3]) ? 9'b000010101 : 9'b101010101;
				assign node21 = (inp[3]) ? node29 : node22;
					assign node22 = (inp[8]) ? node24 : 9'b111010101;
						assign node24 = (inp[9]) ? node26 : 9'b101010101;
							assign node26 = (inp[4]) ? 9'b111010101 : 9'b101010101;
					assign node29 = (inp[0]) ? node41 : node30;
						assign node30 = (inp[9]) ? node34 : node31;
							assign node31 = (inp[8]) ? 9'b101010111 : 9'b111010111;
							assign node34 = (inp[4]) ? 9'b111010111 : node35;
								assign node35 = (inp[8]) ? node37 : 9'b111010111;
									assign node37 = (inp[6]) ? 9'b011010101 : 9'b111010101;
						assign node41 = (inp[8]) ? node43 : 9'b011010111;
							assign node43 = (inp[9]) ? node45 : 9'b001010111;
								assign node45 = (inp[4]) ? 9'b001010101 : 9'b000010111;
		assign node48 = (inp[8]) ? node378 : node49;
			assign node49 = (inp[6]) ? node179 : node50;
				assign node50 = (inp[13]) ? node90 : node51;
					assign node51 = (inp[11]) ? node71 : node52;
						assign node52 = (inp[7]) ? node60 : node53;
							assign node53 = (inp[1]) ? 9'b111011000 : node54;
								assign node54 = (inp[9]) ? 9'b111011000 : node55;
									assign node55 = (inp[2]) ? 9'b111111000 : 9'b111110000;
							assign node60 = (inp[4]) ? node68 : node61;
								assign node61 = (inp[1]) ? 9'b111111000 : node62;
									assign node62 = (inp[9]) ? 9'b111111000 : node63;
										assign node63 = (inp[2]) ? 9'b111111000 : 9'b111110000;
								assign node68 = (inp[9]) ? 9'b111010000 : 9'b111110000;
						assign node71 = (inp[7]) ? node79 : node72;
							assign node72 = (inp[1]) ? 9'b111011100 : node73;
								assign node73 = (inp[9]) ? 9'b111011100 : node74;
									assign node74 = (inp[2]) ? 9'b111111100 : 9'b111110100;
							assign node79 = (inp[4]) ? node87 : node80;
								assign node80 = (inp[2]) ? 9'b111111100 : node81;
									assign node81 = (inp[9]) ? 9'b111111100 : node82;
										assign node82 = (inp[1]) ? 9'b111111100 : 9'b111110100;
								assign node87 = (inp[9]) ? 9'b111010100 : 9'b111110100;
					assign node90 = (inp[3]) ? node110 : node91;
						assign node91 = (inp[7]) ? node99 : node92;
							assign node92 = (inp[9]) ? 9'b111011100 : node93;
								assign node93 = (inp[1]) ? 9'b111011100 : node94;
									assign node94 = (inp[2]) ? 9'b111111100 : 9'b111110100;
							assign node99 = (inp[4]) ? node107 : node100;
								assign node100 = (inp[9]) ? 9'b111111100 : node101;
									assign node101 = (inp[1]) ? 9'b111111100 : node102;
										assign node102 = (inp[2]) ? 9'b111111100 : 9'b111110100;
								assign node107 = (inp[9]) ? 9'b111010100 : 9'b111110100;
						assign node110 = (inp[14]) ? node146 : node111;
							assign node111 = (inp[9]) ? node139 : node112;
								assign node112 = (inp[10]) ? node126 : node113;
									assign node113 = (inp[7]) ? node119 : node114;
										assign node114 = (inp[1]) ? 9'b110011100 : node115;
											assign node115 = (inp[2]) ? 9'b110111100 : 9'b110110100;
										assign node119 = (inp[4]) ? 9'b110110100 : node120;
											assign node120 = (inp[2]) ? 9'b110111100 : node121;
												assign node121 = (inp[1]) ? 9'b110111100 : 9'b110110100;
									assign node126 = (inp[1]) ? node134 : node127;
										assign node127 = (inp[2]) ? node129 : 9'b110110110;
											assign node129 = (inp[7]) ? node131 : 9'b110111110;
												assign node131 = (inp[4]) ? 9'b110110110 : 9'b110111110;
										assign node134 = (inp[7]) ? node136 : 9'b110011110;
											assign node136 = (inp[4]) ? 9'b110110110 : 9'b110111110;
								assign node139 = (inp[4]) ? node143 : node140;
									assign node140 = (inp[7]) ? 9'b110111110 : 9'b110011110;
									assign node143 = (inp[7]) ? 9'b110010110 : 9'b110011110;
							assign node146 = (inp[9]) ? node174 : node147;
								assign node147 = (inp[10]) ? node161 : node148;
									assign node148 = (inp[7]) ? node154 : node149;
										assign node149 = (inp[1]) ? 9'b111011100 : node150;
											assign node150 = (inp[2]) ? 9'b111111100 : 9'b111110100;
										assign node154 = (inp[4]) ? 9'b111110100 : node155;
											assign node155 = (inp[1]) ? 9'b111111100 : node156;
												assign node156 = (inp[2]) ? 9'b111111100 : 9'b111110100;
									assign node161 = (inp[1]) ? node169 : node162;
										assign node162 = (inp[2]) ? node164 : 9'b111110110;
											assign node164 = (inp[4]) ? node166 : 9'b111111110;
												assign node166 = (inp[7]) ? 9'b111110110 : 9'b111111110;
										assign node169 = (inp[7]) ? node171 : 9'b111011110;
											assign node171 = (inp[4]) ? 9'b111110110 : 9'b111111110;
								assign node174 = (inp[7]) ? node176 : 9'b111011110;
									assign node176 = (inp[4]) ? 9'b111010110 : 9'b111111110;
				assign node179 = (inp[13]) ? node219 : node180;
					assign node180 = (inp[11]) ? node200 : node181;
						assign node181 = (inp[7]) ? node189 : node182;
							assign node182 = (inp[9]) ? 9'b111011000 : node183;
								assign node183 = (inp[1]) ? 9'b111011000 : node184;
									assign node184 = (inp[2]) ? 9'b111111000 : 9'b111110000;
							assign node189 = (inp[4]) ? node197 : node190;
								assign node190 = (inp[9]) ? 9'b111111000 : node191;
									assign node191 = (inp[1]) ? 9'b111111000 : node192;
										assign node192 = (inp[2]) ? 9'b111111000 : 9'b111110000;
								assign node197 = (inp[9]) ? 9'b111010000 : 9'b111110000;
						assign node200 = (inp[7]) ? node208 : node201;
							assign node201 = (inp[1]) ? 9'b111011101 : node202;
								assign node202 = (inp[9]) ? 9'b111011101 : node203;
									assign node203 = (inp[2]) ? 9'b111111101 : 9'b111110101;
							assign node208 = (inp[4]) ? node216 : node209;
								assign node209 = (inp[9]) ? 9'b111111101 : node210;
									assign node210 = (inp[1]) ? 9'b111111101 : node211;
										assign node211 = (inp[2]) ? 9'b111111101 : 9'b111110101;
								assign node216 = (inp[9]) ? 9'b111010101 : 9'b111110101;
					assign node219 = (inp[3]) ? node239 : node220;
						assign node220 = (inp[7]) ? node228 : node221;
							assign node221 = (inp[1]) ? 9'b111011101 : node222;
								assign node222 = (inp[9]) ? 9'b111011101 : node223;
									assign node223 = (inp[2]) ? 9'b111111101 : 9'b111110101;
							assign node228 = (inp[4]) ? node236 : node229;
								assign node229 = (inp[2]) ? 9'b111111101 : node230;
									assign node230 = (inp[9]) ? 9'b111111101 : node231;
										assign node231 = (inp[1]) ? 9'b111111101 : 9'b111110101;
								assign node236 = (inp[9]) ? 9'b111010101 : 9'b111110101;
						assign node239 = (inp[5]) ? node309 : node240;
							assign node240 = (inp[14]) ? node274 : node241;
								assign node241 = (inp[9]) ? node269 : node242;
									assign node242 = (inp[10]) ? node256 : node243;
										assign node243 = (inp[1]) ? node251 : node244;
											assign node244 = (inp[2]) ? node246 : 9'b110100101;
												assign node246 = (inp[4]) ? node248 : 9'b110101101;
													assign node248 = (inp[7]) ? 9'b110100101 : 9'b110101101;
											assign node251 = (inp[7]) ? node253 : 9'b110001101;
												assign node253 = (inp[4]) ? 9'b110100101 : 9'b110101101;
										assign node256 = (inp[1]) ? node264 : node257;
											assign node257 = (inp[2]) ? node259 : 9'b110100111;
												assign node259 = (inp[7]) ? node261 : 9'b110101111;
													assign node261 = (inp[4]) ? 9'b110100111 : 9'b110101111;
											assign node264 = (inp[7]) ? node266 : 9'b110001111;
												assign node266 = (inp[4]) ? 9'b110100111 : 9'b110101111;
									assign node269 = (inp[7]) ? node271 : 9'b110001111;
										assign node271 = (inp[4]) ? 9'b110000111 : 9'b110101111;
								assign node274 = (inp[9]) ? node302 : node275;
									assign node275 = (inp[10]) ? node289 : node276;
										assign node276 = (inp[7]) ? node282 : node277;
											assign node277 = (inp[1]) ? 9'b111001101 : node278;
												assign node278 = (inp[2]) ? 9'b111101101 : 9'b111100101;
											assign node282 = (inp[4]) ? 9'b111100101 : node283;
												assign node283 = (inp[1]) ? 9'b111101101 : node284;
													assign node284 = (inp[2]) ? 9'b111101101 : 9'b111100101;
										assign node289 = (inp[7]) ? node295 : node290;
											assign node290 = (inp[1]) ? 9'b111001111 : node291;
												assign node291 = (inp[2]) ? 9'b111101111 : 9'b111100111;
											assign node295 = (inp[4]) ? 9'b111100111 : node296;
												assign node296 = (inp[1]) ? 9'b111101111 : node297;
													assign node297 = (inp[2]) ? 9'b111101111 : 9'b111100111;
									assign node302 = (inp[4]) ? node306 : node303;
										assign node303 = (inp[7]) ? 9'b111101111 : 9'b111001111;
										assign node306 = (inp[7]) ? 9'b111000111 : 9'b111001111;
							assign node309 = (inp[14]) ? node343 : node310;
								assign node310 = (inp[9]) ? node338 : node311;
									assign node311 = (inp[10]) ? node325 : node312;
										assign node312 = (inp[7]) ? node318 : node313;
											assign node313 = (inp[1]) ? 9'b110011101 : node314;
												assign node314 = (inp[2]) ? 9'b110111101 : 9'b110110101;
											assign node318 = (inp[4]) ? 9'b110110101 : node319;
												assign node319 = (inp[2]) ? 9'b110111101 : node320;
													assign node320 = (inp[1]) ? 9'b110111101 : 9'b110110101;
										assign node325 = (inp[7]) ? node331 : node326;
											assign node326 = (inp[1]) ? 9'b110011111 : node327;
												assign node327 = (inp[2]) ? 9'b110111111 : 9'b110110111;
											assign node331 = (inp[4]) ? 9'b110110111 : node332;
												assign node332 = (inp[2]) ? 9'b110111111 : node333;
													assign node333 = (inp[1]) ? 9'b110111111 : 9'b110110111;
									assign node338 = (inp[7]) ? node340 : 9'b110011111;
										assign node340 = (inp[4]) ? 9'b110010111 : 9'b110111111;
								assign node343 = (inp[9]) ? node371 : node344;
									assign node344 = (inp[10]) ? node358 : node345;
										assign node345 = (inp[7]) ? node351 : node346;
											assign node346 = (inp[1]) ? 9'b111011101 : node347;
												assign node347 = (inp[2]) ? 9'b111111101 : 9'b111110101;
											assign node351 = (inp[4]) ? 9'b111110101 : node352;
												assign node352 = (inp[1]) ? 9'b111111101 : node353;
													assign node353 = (inp[2]) ? 9'b111111101 : 9'b111110101;
										assign node358 = (inp[7]) ? node364 : node359;
											assign node359 = (inp[1]) ? 9'b111011111 : node360;
												assign node360 = (inp[2]) ? 9'b111111111 : 9'b111110111;
											assign node364 = (inp[4]) ? 9'b111110111 : node365;
												assign node365 = (inp[1]) ? 9'b111111111 : node366;
													assign node366 = (inp[2]) ? 9'b111111111 : 9'b111110111;
									assign node371 = (inp[4]) ? node375 : node372;
										assign node372 = (inp[7]) ? 9'b111111111 : 9'b111011111;
										assign node375 = (inp[7]) ? 9'b111010111 : 9'b111011111;
			assign node378 = (inp[9]) ? node422 : node379;
				assign node379 = (inp[4]) ? node401 : node380;
					assign node380 = (inp[13]) ? node386 : node381;
						assign node381 = (inp[11]) ? node383 : 9'b101111000;
							assign node383 = (inp[6]) ? 9'b101111101 : 9'b101111100;
						assign node386 = (inp[3]) ? node390 : node387;
							assign node387 = (inp[6]) ? 9'b101111101 : 9'b101111100;
							assign node390 = (inp[6]) ? node394 : node391;
								assign node391 = (inp[14]) ? 9'b101111110 : 9'b100111110;
								assign node394 = (inp[14]) ? node398 : node395;
									assign node395 = (inp[5]) ? 9'b100111111 : 9'b100101111;
									assign node398 = (inp[5]) ? 9'b101111111 : 9'b101101111;
					assign node401 = (inp[13]) ? node407 : node402;
						assign node402 = (inp[11]) ? node404 : 9'b101010000;
							assign node404 = (inp[6]) ? 9'b101010101 : 9'b101010100;
						assign node407 = (inp[3]) ? node411 : node408;
							assign node408 = (inp[6]) ? 9'b101010101 : 9'b101010100;
							assign node411 = (inp[6]) ? node415 : node412;
								assign node412 = (inp[14]) ? 9'b101010110 : 9'b100010110;
								assign node415 = (inp[14]) ? node419 : node416;
									assign node416 = (inp[5]) ? 9'b100010111 : 9'b100000111;
									assign node419 = (inp[5]) ? 9'b101010111 : 9'b101000111;
				assign node422 = (inp[6]) ? node446 : node423;
					assign node423 = (inp[4]) ? node433 : node424;
						assign node424 = (inp[13]) ? node428 : node425;
							assign node425 = (inp[11]) ? 9'b101010100 : 9'b101010000;
							assign node428 = (inp[3]) ? node430 : 9'b101010100;
								assign node430 = (inp[0]) ? 9'b100010110 : 9'b111010100;
						assign node433 = (inp[13]) ? node437 : node434;
							assign node434 = (inp[11]) ? 9'b111010100 : 9'b111010000;
							assign node437 = (inp[3]) ? node439 : 9'b111010100;
								assign node439 = (inp[0]) ? node443 : node440;
									assign node440 = (inp[14]) ? 9'b111010110 : 9'b110010110;
									assign node443 = (inp[14]) ? 9'b101010100 : 9'b100010100;
					assign node446 = (inp[13]) ? node454 : node447;
						assign node447 = (inp[11]) ? node451 : node448;
							assign node448 = (inp[4]) ? 9'b111010000 : 9'b101010000;
							assign node451 = (inp[4]) ? 9'b111010101 : 9'b101010101;
						assign node454 = (inp[3]) ? node458 : node455;
							assign node455 = (inp[4]) ? 9'b111010101 : 9'b101010101;
							assign node458 = (inp[0]) ? node470 : node459;
								assign node459 = (inp[4]) ? node463 : node460;
									assign node460 = (inp[5]) ? 9'b011010101 : 9'b011000101;
									assign node463 = (inp[5]) ? node467 : node464;
										assign node464 = (inp[14]) ? 9'b111000111 : 9'b110000111;
										assign node467 = (inp[14]) ? 9'b111010111 : 9'b110010111;
								assign node470 = (inp[4]) ? node474 : node471;
									assign node471 = (inp[5]) ? 9'b100010111 : 9'b100000111;
									assign node474 = (inp[5]) ? node478 : node475;
										assign node475 = (inp[14]) ? 9'b101000101 : 9'b100000101;
										assign node478 = (inp[14]) ? 9'b101010101 : 9'b100010101;

endmodule