module dtc_split66_bm39 (
	input  wire [14-1:0] inp,
	output wire [14-1:0] outp
);

	wire [14-1:0] node1;
	wire [14-1:0] node3;
	wire [14-1:0] node4;
	wire [14-1:0] node5;
	wire [14-1:0] node6;
	wire [14-1:0] node7;
	wire [14-1:0] node8;
	wire [14-1:0] node9;
	wire [14-1:0] node10;
	wire [14-1:0] node11;
	wire [14-1:0] node12;
	wire [14-1:0] node13;
	wire [14-1:0] node17;
	wire [14-1:0] node18;
	wire [14-1:0] node21;
	wire [14-1:0] node24;
	wire [14-1:0] node25;
	wire [14-1:0] node26;
	wire [14-1:0] node29;
	wire [14-1:0] node32;
	wire [14-1:0] node33;
	wire [14-1:0] node36;
	wire [14-1:0] node39;
	wire [14-1:0] node40;
	wire [14-1:0] node41;
	wire [14-1:0] node42;
	wire [14-1:0] node45;
	wire [14-1:0] node48;
	wire [14-1:0] node49;
	wire [14-1:0] node52;
	wire [14-1:0] node55;
	wire [14-1:0] node56;
	wire [14-1:0] node57;
	wire [14-1:0] node61;
	wire [14-1:0] node62;
	wire [14-1:0] node65;
	wire [14-1:0] node68;
	wire [14-1:0] node69;
	wire [14-1:0] node70;
	wire [14-1:0] node72;
	wire [14-1:0] node73;
	wire [14-1:0] node76;
	wire [14-1:0] node79;
	wire [14-1:0] node80;
	wire [14-1:0] node81;
	wire [14-1:0] node85;
	wire [14-1:0] node86;
	wire [14-1:0] node90;
	wire [14-1:0] node91;
	wire [14-1:0] node92;
	wire [14-1:0] node93;
	wire [14-1:0] node96;
	wire [14-1:0] node99;
	wire [14-1:0] node100;
	wire [14-1:0] node103;
	wire [14-1:0] node106;
	wire [14-1:0] node107;
	wire [14-1:0] node108;
	wire [14-1:0] node111;
	wire [14-1:0] node114;
	wire [14-1:0] node115;
	wire [14-1:0] node118;
	wire [14-1:0] node121;
	wire [14-1:0] node122;
	wire [14-1:0] node123;
	wire [14-1:0] node124;
	wire [14-1:0] node125;
	wire [14-1:0] node126;
	wire [14-1:0] node129;
	wire [14-1:0] node132;
	wire [14-1:0] node133;
	wire [14-1:0] node136;
	wire [14-1:0] node139;
	wire [14-1:0] node140;
	wire [14-1:0] node141;
	wire [14-1:0] node144;
	wire [14-1:0] node147;
	wire [14-1:0] node148;
	wire [14-1:0] node151;
	wire [14-1:0] node154;
	wire [14-1:0] node155;
	wire [14-1:0] node156;
	wire [14-1:0] node157;
	wire [14-1:0] node161;
	wire [14-1:0] node162;
	wire [14-1:0] node165;
	wire [14-1:0] node169;
	wire [14-1:0] node170;
	wire [14-1:0] node172;
	wire [14-1:0] node173;
	wire [14-1:0] node175;
	wire [14-1:0] node178;
	wire [14-1:0] node179;
	wire [14-1:0] node183;
	wire [14-1:0] node184;
	wire [14-1:0] node185;
	wire [14-1:0] node186;
	wire [14-1:0] node189;
	wire [14-1:0] node192;
	wire [14-1:0] node193;
	wire [14-1:0] node196;
	wire [14-1:0] node200;
	wire [14-1:0] node201;
	wire [14-1:0] node202;
	wire [14-1:0] node203;
	wire [14-1:0] node204;
	wire [14-1:0] node205;
	wire [14-1:0] node207;
	wire [14-1:0] node210;
	wire [14-1:0] node211;
	wire [14-1:0] node214;
	wire [14-1:0] node217;
	wire [14-1:0] node218;
	wire [14-1:0] node220;
	wire [14-1:0] node223;
	wire [14-1:0] node224;
	wire [14-1:0] node227;
	wire [14-1:0] node230;
	wire [14-1:0] node231;
	wire [14-1:0] node232;
	wire [14-1:0] node234;
	wire [14-1:0] node237;
	wire [14-1:0] node238;
	wire [14-1:0] node241;
	wire [14-1:0] node244;
	wire [14-1:0] node245;
	wire [14-1:0] node246;
	wire [14-1:0] node249;
	wire [14-1:0] node252;
	wire [14-1:0] node253;
	wire [14-1:0] node256;
	wire [14-1:0] node259;
	wire [14-1:0] node260;
	wire [14-1:0] node261;
	wire [14-1:0] node262;
	wire [14-1:0] node263;
	wire [14-1:0] node266;
	wire [14-1:0] node269;
	wire [14-1:0] node270;
	wire [14-1:0] node273;
	wire [14-1:0] node277;
	wire [14-1:0] node278;
	wire [14-1:0] node279;
	wire [14-1:0] node280;
	wire [14-1:0] node283;
	wire [14-1:0] node286;
	wire [14-1:0] node287;
	wire [14-1:0] node290;
	wire [14-1:0] node293;
	wire [14-1:0] node294;
	wire [14-1:0] node295;
	wire [14-1:0] node298;
	wire [14-1:0] node301;
	wire [14-1:0] node302;
	wire [14-1:0] node305;
	wire [14-1:0] node308;
	wire [14-1:0] node309;
	wire [14-1:0] node310;
	wire [14-1:0] node311;
	wire [14-1:0] node312;
	wire [14-1:0] node313;
	wire [14-1:0] node317;
	wire [14-1:0] node318;
	wire [14-1:0] node322;
	wire [14-1:0] node323;
	wire [14-1:0] node324;
	wire [14-1:0] node327;
	wire [14-1:0] node330;
	wire [14-1:0] node332;
	wire [14-1:0] node335;
	wire [14-1:0] node337;
	wire [14-1:0] node338;
	wire [14-1:0] node339;
	wire [14-1:0] node342;
	wire [14-1:0] node345;
	wire [14-1:0] node346;
	wire [14-1:0] node351;
	wire [14-1:0] node352;
	wire [14-1:0] node353;
	wire [14-1:0] node354;
	wire [14-1:0] node355;
	wire [14-1:0] node356;
	wire [14-1:0] node357;
	wire [14-1:0] node358;
	wire [14-1:0] node361;
	wire [14-1:0] node364;
	wire [14-1:0] node365;
	wire [14-1:0] node368;
	wire [14-1:0] node371;
	wire [14-1:0] node372;
	wire [14-1:0] node374;
	wire [14-1:0] node377;
	wire [14-1:0] node378;
	wire [14-1:0] node381;
	wire [14-1:0] node384;
	wire [14-1:0] node385;
	wire [14-1:0] node386;
	wire [14-1:0] node387;
	wire [14-1:0] node390;
	wire [14-1:0] node393;
	wire [14-1:0] node394;
	wire [14-1:0] node398;
	wire [14-1:0] node399;
	wire [14-1:0] node401;
	wire [14-1:0] node404;
	wire [14-1:0] node407;
	wire [14-1:0] node408;
	wire [14-1:0] node409;
	wire [14-1:0] node410;
	wire [14-1:0] node411;
	wire [14-1:0] node414;
	wire [14-1:0] node417;
	wire [14-1:0] node418;
	wire [14-1:0] node422;
	wire [14-1:0] node423;
	wire [14-1:0] node424;
	wire [14-1:0] node427;
	wire [14-1:0] node430;
	wire [14-1:0] node432;
	wire [14-1:0] node435;
	wire [14-1:0] node436;
	wire [14-1:0] node437;
	wire [14-1:0] node439;
	wire [14-1:0] node442;
	wire [14-1:0] node443;
	wire [14-1:0] node446;
	wire [14-1:0] node450;
	wire [14-1:0] node451;
	wire [14-1:0] node453;
	wire [14-1:0] node454;
	wire [14-1:0] node455;
	wire [14-1:0] node456;
	wire [14-1:0] node459;
	wire [14-1:0] node462;
	wire [14-1:0] node463;
	wire [14-1:0] node467;
	wire [14-1:0] node468;
	wire [14-1:0] node469;
	wire [14-1:0] node472;
	wire [14-1:0] node475;
	wire [14-1:0] node476;
	wire [14-1:0] node479;
	wire [14-1:0] node483;
	wire [14-1:0] node484;
	wire [14-1:0] node486;
	wire [14-1:0] node487;
	wire [14-1:0] node488;
	wire [14-1:0] node489;
	wire [14-1:0] node490;
	wire [14-1:0] node493;
	wire [14-1:0] node496;
	wire [14-1:0] node497;
	wire [14-1:0] node501;
	wire [14-1:0] node502;
	wire [14-1:0] node503;
	wire [14-1:0] node506;
	wire [14-1:0] node509;
	wire [14-1:0] node510;
	wire [14-1:0] node513;
	wire [14-1:0] node516;
	wire [14-1:0] node517;
	wire [14-1:0] node518;
	wire [14-1:0] node519;
	wire [14-1:0] node522;
	wire [14-1:0] node525;
	wire [14-1:0] node526;
	wire [14-1:0] node529;
	wire [14-1:0] node532;
	wire [14-1:0] node533;
	wire [14-1:0] node535;
	wire [14-1:0] node540;
	wire [14-1:0] node541;
	wire [14-1:0] node542;
	wire [14-1:0] node543;
	wire [14-1:0] node544;
	wire [14-1:0] node545;
	wire [14-1:0] node546;
	wire [14-1:0] node548;
	wire [14-1:0] node549;
	wire [14-1:0] node552;
	wire [14-1:0] node555;
	wire [14-1:0] node556;
	wire [14-1:0] node557;
	wire [14-1:0] node561;
	wire [14-1:0] node563;
	wire [14-1:0] node566;
	wire [14-1:0] node567;
	wire [14-1:0] node568;
	wire [14-1:0] node569;
	wire [14-1:0] node572;
	wire [14-1:0] node575;
	wire [14-1:0] node576;
	wire [14-1:0] node579;
	wire [14-1:0] node582;
	wire [14-1:0] node583;
	wire [14-1:0] node584;
	wire [14-1:0] node587;
	wire [14-1:0] node590;
	wire [14-1:0] node591;
	wire [14-1:0] node594;
	wire [14-1:0] node597;
	wire [14-1:0] node598;
	wire [14-1:0] node599;
	wire [14-1:0] node600;
	wire [14-1:0] node601;
	wire [14-1:0] node604;
	wire [14-1:0] node607;
	wire [14-1:0] node608;
	wire [14-1:0] node611;
	wire [14-1:0] node614;
	wire [14-1:0] node615;
	wire [14-1:0] node616;
	wire [14-1:0] node619;
	wire [14-1:0] node622;
	wire [14-1:0] node623;
	wire [14-1:0] node626;
	wire [14-1:0] node629;
	wire [14-1:0] node630;
	wire [14-1:0] node631;
	wire [14-1:0] node632;
	wire [14-1:0] node635;
	wire [14-1:0] node638;
	wire [14-1:0] node639;
	wire [14-1:0] node642;
	wire [14-1:0] node645;
	wire [14-1:0] node646;
	wire [14-1:0] node648;
	wire [14-1:0] node651;
	wire [14-1:0] node652;
	wire [14-1:0] node655;
	wire [14-1:0] node658;
	wire [14-1:0] node659;
	wire [14-1:0] node660;
	wire [14-1:0] node661;
	wire [14-1:0] node662;
	wire [14-1:0] node663;
	wire [14-1:0] node666;
	wire [14-1:0] node669;
	wire [14-1:0] node670;
	wire [14-1:0] node673;
	wire [14-1:0] node676;
	wire [14-1:0] node677;
	wire [14-1:0] node678;
	wire [14-1:0] node681;
	wire [14-1:0] node684;
	wire [14-1:0] node685;
	wire [14-1:0] node688;
	wire [14-1:0] node691;
	wire [14-1:0] node692;
	wire [14-1:0] node694;
	wire [14-1:0] node695;
	wire [14-1:0] node698;
	wire [14-1:0] node702;
	wire [14-1:0] node704;
	wire [14-1:0] node705;
	wire [14-1:0] node706;
	wire [14-1:0] node707;
	wire [14-1:0] node710;
	wire [14-1:0] node713;
	wire [14-1:0] node714;
	wire [14-1:0] node717;
	wire [14-1:0] node721;
	wire [14-1:0] node722;
	wire [14-1:0] node723;
	wire [14-1:0] node725;
	wire [14-1:0] node726;
	wire [14-1:0] node727;
	wire [14-1:0] node728;
	wire [14-1:0] node734;
	wire [14-1:0] node735;
	wire [14-1:0] node736;
	wire [14-1:0] node737;
	wire [14-1:0] node738;
	wire [14-1:0] node741;
	wire [14-1:0] node744;
	wire [14-1:0] node745;
	wire [14-1:0] node749;
	wire [14-1:0] node750;
	wire [14-1:0] node751;
	wire [14-1:0] node754;
	wire [14-1:0] node757;
	wire [14-1:0] node758;
	wire [14-1:0] node761;
	wire [14-1:0] node764;
	wire [14-1:0] node765;
	wire [14-1:0] node766;
	wire [14-1:0] node767;
	wire [14-1:0] node770;
	wire [14-1:0] node773;
	wire [14-1:0] node774;
	wire [14-1:0] node777;
	wire [14-1:0] node780;
	wire [14-1:0] node782;
	wire [14-1:0] node783;
	wire [14-1:0] node789;
	wire [14-1:0] node790;
	wire [14-1:0] node791;
	wire [14-1:0] node792;
	wire [14-1:0] node793;
	wire [14-1:0] node794;
	wire [14-1:0] node795;
	wire [14-1:0] node796;
	wire [14-1:0] node797;
	wire [14-1:0] node799;
	wire [14-1:0] node802;
	wire [14-1:0] node803;
	wire [14-1:0] node806;
	wire [14-1:0] node809;
	wire [14-1:0] node810;
	wire [14-1:0] node811;
	wire [14-1:0] node814;
	wire [14-1:0] node817;
	wire [14-1:0] node818;
	wire [14-1:0] node821;
	wire [14-1:0] node824;
	wire [14-1:0] node825;
	wire [14-1:0] node826;
	wire [14-1:0] node827;
	wire [14-1:0] node830;
	wire [14-1:0] node833;
	wire [14-1:0] node834;
	wire [14-1:0] node837;
	wire [14-1:0] node840;
	wire [14-1:0] node841;
	wire [14-1:0] node842;
	wire [14-1:0] node845;
	wire [14-1:0] node848;
	wire [14-1:0] node850;
	wire [14-1:0] node853;
	wire [14-1:0] node854;
	wire [14-1:0] node855;
	wire [14-1:0] node856;
	wire [14-1:0] node857;
	wire [14-1:0] node860;
	wire [14-1:0] node863;
	wire [14-1:0] node864;
	wire [14-1:0] node867;
	wire [14-1:0] node870;
	wire [14-1:0] node871;
	wire [14-1:0] node873;
	wire [14-1:0] node877;
	wire [14-1:0] node879;
	wire [14-1:0] node880;
	wire [14-1:0] node881;
	wire [14-1:0] node886;
	wire [14-1:0] node887;
	wire [14-1:0] node888;
	wire [14-1:0] node889;
	wire [14-1:0] node890;
	wire [14-1:0] node891;
	wire [14-1:0] node894;
	wire [14-1:0] node897;
	wire [14-1:0] node898;
	wire [14-1:0] node902;
	wire [14-1:0] node903;
	wire [14-1:0] node904;
	wire [14-1:0] node907;
	wire [14-1:0] node910;
	wire [14-1:0] node911;
	wire [14-1:0] node914;
	wire [14-1:0] node917;
	wire [14-1:0] node918;
	wire [14-1:0] node919;
	wire [14-1:0] node921;
	wire [14-1:0] node924;
	wire [14-1:0] node925;
	wire [14-1:0] node928;
	wire [14-1:0] node931;
	wire [14-1:0] node932;
	wire [14-1:0] node933;
	wire [14-1:0] node939;
	wire [14-1:0] node940;
	wire [14-1:0] node941;
	wire [14-1:0] node942;
	wire [14-1:0] node943;
	wire [14-1:0] node944;
	wire [14-1:0] node946;
	wire [14-1:0] node949;
	wire [14-1:0] node950;
	wire [14-1:0] node953;
	wire [14-1:0] node956;
	wire [14-1:0] node957;
	wire [14-1:0] node958;
	wire [14-1:0] node961;
	wire [14-1:0] node964;
	wire [14-1:0] node965;
	wire [14-1:0] node968;
	wire [14-1:0] node971;
	wire [14-1:0] node972;
	wire [14-1:0] node973;
	wire [14-1:0] node974;
	wire [14-1:0] node977;
	wire [14-1:0] node980;
	wire [14-1:0] node982;
	wire [14-1:0] node985;
	wire [14-1:0] node987;
	wire [14-1:0] node990;
	wire [14-1:0] node992;
	wire [14-1:0] node993;
	wire [14-1:0] node994;
	wire [14-1:0] node995;
	wire [14-1:0] node998;
	wire [14-1:0] node1001;
	wire [14-1:0] node1002;
	wire [14-1:0] node1005;
	wire [14-1:0] node1008;
	wire [14-1:0] node1009;
	wire [14-1:0] node1010;
	wire [14-1:0] node1015;
	wire [14-1:0] node1017;
	wire [14-1:0] node1018;
	wire [14-1:0] node1019;
	wire [14-1:0] node1020;
	wire [14-1:0] node1021;
	wire [14-1:0] node1024;
	wire [14-1:0] node1027;
	wire [14-1:0] node1028;
	wire [14-1:0] node1031;
	wire [14-1:0] node1034;
	wire [14-1:0] node1035;
	wire [14-1:0] node1038;
	wire [14-1:0] node1039;
	wire [14-1:0] node1042;
	wire [14-1:0] node1046;
	wire [14-1:0] node1047;
	wire [14-1:0] node1048;
	wire [14-1:0] node1049;
	wire [14-1:0] node1050;
	wire [14-1:0] node1051;
	wire [14-1:0] node1052;
	wire [14-1:0] node1053;
	wire [14-1:0] node1056;
	wire [14-1:0] node1059;
	wire [14-1:0] node1060;
	wire [14-1:0] node1063;
	wire [14-1:0] node1066;
	wire [14-1:0] node1067;
	wire [14-1:0] node1068;
	wire [14-1:0] node1071;
	wire [14-1:0] node1075;
	wire [14-1:0] node1076;
	wire [14-1:0] node1077;
	wire [14-1:0] node1078;
	wire [14-1:0] node1081;
	wire [14-1:0] node1084;
	wire [14-1:0] node1086;
	wire [14-1:0] node1089;
	wire [14-1:0] node1090;
	wire [14-1:0] node1092;
	wire [14-1:0] node1096;
	wire [14-1:0] node1097;
	wire [14-1:0] node1098;
	wire [14-1:0] node1099;
	wire [14-1:0] node1101;
	wire [14-1:0] node1104;
	wire [14-1:0] node1106;
	wire [14-1:0] node1109;
	wire [14-1:0] node1110;
	wire [14-1:0] node1112;
	wire [14-1:0] node1117;
	wire [14-1:0] node1118;
	wire [14-1:0] node1119;
	wire [14-1:0] node1120;
	wire [14-1:0] node1121;
	wire [14-1:0] node1123;
	wire [14-1:0] node1126;
	wire [14-1:0] node1127;
	wire [14-1:0] node1132;
	wire [14-1:0] node1133;
	wire [14-1:0] node1134;
	wire [14-1:0] node1135;
	wire [14-1:0] node1138;
	wire [14-1:0] node1141;
	wire [14-1:0] node1142;
	wire [14-1:0] node1146;
	wire [14-1:0] node1147;
	wire [14-1:0] node1148;
	wire [14-1:0] node1151;
	wire [14-1:0] node1154;
	wire [14-1:0] node1156;
	wire [14-1:0] node1159;
	wire [14-1:0] node1161;
	wire [14-1:0] node1162;
	wire [14-1:0] node1163;
	wire [14-1:0] node1164;
	wire [14-1:0] node1167;
	wire [14-1:0] node1170;
	wire [14-1:0] node1171;
	wire [14-1:0] node1174;
	wire [14-1:0] node1180;
	wire [14-1:0] node1181;
	wire [14-1:0] node1182;
	wire [14-1:0] node1183;
	wire [14-1:0] node1184;
	wire [14-1:0] node1185;
	wire [14-1:0] node1186;
	wire [14-1:0] node1187;
	wire [14-1:0] node1188;
	wire [14-1:0] node1189;
	wire [14-1:0] node1190;
	wire [14-1:0] node1191;
	wire [14-1:0] node1198;
	wire [14-1:0] node1199;
	wire [14-1:0] node1200;
	wire [14-1:0] node1201;
	wire [14-1:0] node1203;
	wire [14-1:0] node1206;
	wire [14-1:0] node1207;
	wire [14-1:0] node1211;
	wire [14-1:0] node1212;
	wire [14-1:0] node1213;
	wire [14-1:0] node1216;
	wire [14-1:0] node1219;
	wire [14-1:0] node1222;
	wire [14-1:0] node1223;
	wire [14-1:0] node1224;
	wire [14-1:0] node1225;
	wire [14-1:0] node1228;
	wire [14-1:0] node1231;
	wire [14-1:0] node1234;
	wire [14-1:0] node1235;
	wire [14-1:0] node1236;
	wire [14-1:0] node1239;
	wire [14-1:0] node1242;
	wire [14-1:0] node1245;
	wire [14-1:0] node1246;
	wire [14-1:0] node1247;
	wire [14-1:0] node1248;
	wire [14-1:0] node1249;
	wire [14-1:0] node1251;
	wire [14-1:0] node1255;
	wire [14-1:0] node1256;
	wire [14-1:0] node1257;
	wire [14-1:0] node1260;
	wire [14-1:0] node1263;
	wire [14-1:0] node1266;
	wire [14-1:0] node1267;
	wire [14-1:0] node1268;
	wire [14-1:0] node1271;
	wire [14-1:0] node1274;
	wire [14-1:0] node1275;
	wire [14-1:0] node1276;
	wire [14-1:0] node1279;
	wire [14-1:0] node1282;
	wire [14-1:0] node1285;
	wire [14-1:0] node1286;
	wire [14-1:0] node1287;
	wire [14-1:0] node1288;
	wire [14-1:0] node1290;
	wire [14-1:0] node1293;
	wire [14-1:0] node1296;
	wire [14-1:0] node1297;
	wire [14-1:0] node1298;
	wire [14-1:0] node1301;
	wire [14-1:0] node1304;
	wire [14-1:0] node1307;
	wire [14-1:0] node1308;
	wire [14-1:0] node1309;
	wire [14-1:0] node1310;
	wire [14-1:0] node1313;
	wire [14-1:0] node1316;
	wire [14-1:0] node1319;
	wire [14-1:0] node1320;
	wire [14-1:0] node1321;
	wire [14-1:0] node1324;
	wire [14-1:0] node1327;
	wire [14-1:0] node1330;
	wire [14-1:0] node1331;
	wire [14-1:0] node1332;
	wire [14-1:0] node1333;
	wire [14-1:0] node1334;
	wire [14-1:0] node1336;
	wire [14-1:0] node1337;
	wire [14-1:0] node1341;
	wire [14-1:0] node1342;
	wire [14-1:0] node1343;
	wire [14-1:0] node1346;
	wire [14-1:0] node1349;
	wire [14-1:0] node1352;
	wire [14-1:0] node1353;
	wire [14-1:0] node1354;
	wire [14-1:0] node1355;
	wire [14-1:0] node1358;
	wire [14-1:0] node1361;
	wire [14-1:0] node1364;
	wire [14-1:0] node1365;
	wire [14-1:0] node1366;
	wire [14-1:0] node1369;
	wire [14-1:0] node1372;
	wire [14-1:0] node1375;
	wire [14-1:0] node1376;
	wire [14-1:0] node1377;
	wire [14-1:0] node1378;
	wire [14-1:0] node1381;
	wire [14-1:0] node1384;
	wire [14-1:0] node1386;
	wire [14-1:0] node1389;
	wire [14-1:0] node1390;
	wire [14-1:0] node1391;
	wire [14-1:0] node1392;
	wire [14-1:0] node1395;
	wire [14-1:0] node1398;
	wire [14-1:0] node1401;
	wire [14-1:0] node1402;
	wire [14-1:0] node1403;
	wire [14-1:0] node1406;
	wire [14-1:0] node1409;
	wire [14-1:0] node1412;
	wire [14-1:0] node1413;
	wire [14-1:0] node1414;
	wire [14-1:0] node1415;
	wire [14-1:0] node1416;
	wire [14-1:0] node1419;
	wire [14-1:0] node1422;
	wire [14-1:0] node1423;
	wire [14-1:0] node1424;
	wire [14-1:0] node1427;
	wire [14-1:0] node1430;
	wire [14-1:0] node1433;
	wire [14-1:0] node1434;
	wire [14-1:0] node1435;
	wire [14-1:0] node1436;
	wire [14-1:0] node1439;
	wire [14-1:0] node1442;
	wire [14-1:0] node1445;
	wire [14-1:0] node1446;
	wire [14-1:0] node1447;
	wire [14-1:0] node1450;
	wire [14-1:0] node1453;
	wire [14-1:0] node1456;
	wire [14-1:0] node1457;
	wire [14-1:0] node1458;
	wire [14-1:0] node1459;
	wire [14-1:0] node1460;
	wire [14-1:0] node1464;
	wire [14-1:0] node1467;
	wire [14-1:0] node1468;
	wire [14-1:0] node1469;
	wire [14-1:0] node1472;
	wire [14-1:0] node1475;
	wire [14-1:0] node1476;
	wire [14-1:0] node1479;
	wire [14-1:0] node1482;
	wire [14-1:0] node1483;
	wire [14-1:0] node1484;
	wire [14-1:0] node1487;
	wire [14-1:0] node1490;
	wire [14-1:0] node1491;
	wire [14-1:0] node1494;
	wire [14-1:0] node1497;
	wire [14-1:0] node1498;
	wire [14-1:0] node1499;
	wire [14-1:0] node1500;
	wire [14-1:0] node1501;
	wire [14-1:0] node1502;
	wire [14-1:0] node1503;
	wire [14-1:0] node1506;
	wire [14-1:0] node1507;
	wire [14-1:0] node1510;
	wire [14-1:0] node1513;
	wire [14-1:0] node1514;
	wire [14-1:0] node1515;
	wire [14-1:0] node1518;
	wire [14-1:0] node1521;
	wire [14-1:0] node1522;
	wire [14-1:0] node1525;
	wire [14-1:0] node1528;
	wire [14-1:0] node1529;
	wire [14-1:0] node1530;
	wire [14-1:0] node1531;
	wire [14-1:0] node1534;
	wire [14-1:0] node1537;
	wire [14-1:0] node1539;
	wire [14-1:0] node1542;
	wire [14-1:0] node1543;
	wire [14-1:0] node1544;
	wire [14-1:0] node1548;
	wire [14-1:0] node1549;
	wire [14-1:0] node1552;
	wire [14-1:0] node1555;
	wire [14-1:0] node1556;
	wire [14-1:0] node1557;
	wire [14-1:0] node1559;
	wire [14-1:0] node1560;
	wire [14-1:0] node1563;
	wire [14-1:0] node1566;
	wire [14-1:0] node1567;
	wire [14-1:0] node1568;
	wire [14-1:0] node1571;
	wire [14-1:0] node1574;
	wire [14-1:0] node1575;
	wire [14-1:0] node1578;
	wire [14-1:0] node1581;
	wire [14-1:0] node1582;
	wire [14-1:0] node1583;
	wire [14-1:0] node1584;
	wire [14-1:0] node1587;
	wire [14-1:0] node1590;
	wire [14-1:0] node1591;
	wire [14-1:0] node1594;
	wire [14-1:0] node1597;
	wire [14-1:0] node1598;
	wire [14-1:0] node1600;
	wire [14-1:0] node1603;
	wire [14-1:0] node1604;
	wire [14-1:0] node1607;
	wire [14-1:0] node1610;
	wire [14-1:0] node1612;
	wire [14-1:0] node1613;
	wire [14-1:0] node1614;
	wire [14-1:0] node1616;
	wire [14-1:0] node1619;
	wire [14-1:0] node1620;
	wire [14-1:0] node1621;
	wire [14-1:0] node1624;
	wire [14-1:0] node1627;
	wire [14-1:0] node1628;
	wire [14-1:0] node1631;
	wire [14-1:0] node1634;
	wire [14-1:0] node1635;
	wire [14-1:0] node1636;
	wire [14-1:0] node1637;
	wire [14-1:0] node1640;
	wire [14-1:0] node1643;
	wire [14-1:0] node1644;
	wire [14-1:0] node1647;
	wire [14-1:0] node1650;
	wire [14-1:0] node1651;
	wire [14-1:0] node1653;
	wire [14-1:0] node1656;
	wire [14-1:0] node1657;
	wire [14-1:0] node1661;
	wire [14-1:0] node1662;
	wire [14-1:0] node1663;
	wire [14-1:0] node1664;
	wire [14-1:0] node1666;
	wire [14-1:0] node1667;
	wire [14-1:0] node1668;
	wire [14-1:0] node1671;
	wire [14-1:0] node1674;
	wire [14-1:0] node1675;
	wire [14-1:0] node1678;
	wire [14-1:0] node1681;
	wire [14-1:0] node1682;
	wire [14-1:0] node1683;
	wire [14-1:0] node1684;
	wire [14-1:0] node1687;
	wire [14-1:0] node1690;
	wire [14-1:0] node1691;
	wire [14-1:0] node1694;
	wire [14-1:0] node1697;
	wire [14-1:0] node1698;
	wire [14-1:0] node1700;
	wire [14-1:0] node1703;
	wire [14-1:0] node1704;
	wire [14-1:0] node1707;
	wire [14-1:0] node1712;
	wire [14-1:0] node1713;
	wire [14-1:0] node1714;
	wire [14-1:0] node1715;
	wire [14-1:0] node1716;
	wire [14-1:0] node1717;
	wire [14-1:0] node1718;
	wire [14-1:0] node1720;
	wire [14-1:0] node1724;
	wire [14-1:0] node1725;
	wire [14-1:0] node1726;
	wire [14-1:0] node1727;
	wire [14-1:0] node1730;
	wire [14-1:0] node1733;
	wire [14-1:0] node1734;
	wire [14-1:0] node1737;
	wire [14-1:0] node1740;
	wire [14-1:0] node1741;
	wire [14-1:0] node1744;
	wire [14-1:0] node1747;
	wire [14-1:0] node1748;
	wire [14-1:0] node1749;
	wire [14-1:0] node1750;
	wire [14-1:0] node1751;
	wire [14-1:0] node1754;
	wire [14-1:0] node1757;
	wire [14-1:0] node1758;
	wire [14-1:0] node1761;
	wire [14-1:0] node1764;
	wire [14-1:0] node1765;
	wire [14-1:0] node1766;
	wire [14-1:0] node1769;
	wire [14-1:0] node1772;
	wire [14-1:0] node1773;
	wire [14-1:0] node1776;
	wire [14-1:0] node1779;
	wire [14-1:0] node1780;
	wire [14-1:0] node1782;
	wire [14-1:0] node1785;
	wire [14-1:0] node1786;
	wire [14-1:0] node1789;
	wire [14-1:0] node1792;
	wire [14-1:0] node1793;
	wire [14-1:0] node1794;
	wire [14-1:0] node1795;
	wire [14-1:0] node1796;
	wire [14-1:0] node1797;
	wire [14-1:0] node1800;
	wire [14-1:0] node1803;
	wire [14-1:0] node1804;
	wire [14-1:0] node1808;
	wire [14-1:0] node1809;
	wire [14-1:0] node1812;
	wire [14-1:0] node1815;
	wire [14-1:0] node1816;
	wire [14-1:0] node1817;
	wire [14-1:0] node1818;
	wire [14-1:0] node1821;
	wire [14-1:0] node1824;
	wire [14-1:0] node1827;
	wire [14-1:0] node1828;
	wire [14-1:0] node1830;
	wire [14-1:0] node1833;
	wire [14-1:0] node1836;
	wire [14-1:0] node1837;
	wire [14-1:0] node1838;
	wire [14-1:0] node1839;
	wire [14-1:0] node1840;
	wire [14-1:0] node1843;
	wire [14-1:0] node1846;
	wire [14-1:0] node1849;
	wire [14-1:0] node1850;
	wire [14-1:0] node1851;
	wire [14-1:0] node1854;
	wire [14-1:0] node1857;
	wire [14-1:0] node1860;
	wire [14-1:0] node1861;
	wire [14-1:0] node1862;
	wire [14-1:0] node1863;
	wire [14-1:0] node1866;
	wire [14-1:0] node1869;
	wire [14-1:0] node1872;
	wire [14-1:0] node1873;
	wire [14-1:0] node1874;
	wire [14-1:0] node1877;
	wire [14-1:0] node1880;
	wire [14-1:0] node1883;
	wire [14-1:0] node1884;
	wire [14-1:0] node1885;
	wire [14-1:0] node1886;
	wire [14-1:0] node1887;
	wire [14-1:0] node1888;
	wire [14-1:0] node1890;
	wire [14-1:0] node1893;
	wire [14-1:0] node1894;
	wire [14-1:0] node1898;
	wire [14-1:0] node1899;
	wire [14-1:0] node1900;
	wire [14-1:0] node1903;
	wire [14-1:0] node1906;
	wire [14-1:0] node1907;
	wire [14-1:0] node1910;
	wire [14-1:0] node1913;
	wire [14-1:0] node1914;
	wire [14-1:0] node1915;
	wire [14-1:0] node1916;
	wire [14-1:0] node1919;
	wire [14-1:0] node1922;
	wire [14-1:0] node1923;
	wire [14-1:0] node1926;
	wire [14-1:0] node1929;
	wire [14-1:0] node1930;
	wire [14-1:0] node1931;
	wire [14-1:0] node1934;
	wire [14-1:0] node1937;
	wire [14-1:0] node1938;
	wire [14-1:0] node1941;
	wire [14-1:0] node1944;
	wire [14-1:0] node1946;
	wire [14-1:0] node1947;
	wire [14-1:0] node1948;
	wire [14-1:0] node1949;
	wire [14-1:0] node1952;
	wire [14-1:0] node1955;
	wire [14-1:0] node1956;
	wire [14-1:0] node1959;
	wire [14-1:0] node1962;
	wire [14-1:0] node1963;
	wire [14-1:0] node1964;
	wire [14-1:0] node1967;
	wire [14-1:0] node1970;
	wire [14-1:0] node1971;
	wire [14-1:0] node1974;
	wire [14-1:0] node1977;
	wire [14-1:0] node1978;
	wire [14-1:0] node1979;
	wire [14-1:0] node1980;
	wire [14-1:0] node1982;
	wire [14-1:0] node1985;
	wire [14-1:0] node1986;
	wire [14-1:0] node1987;
	wire [14-1:0] node1990;
	wire [14-1:0] node1993;
	wire [14-1:0] node1994;
	wire [14-1:0] node1997;
	wire [14-1:0] node2002;
	wire [14-1:0] node2004;
	wire [14-1:0] node2005;
	wire [14-1:0] node2006;
	wire [14-1:0] node2007;
	wire [14-1:0] node2008;
	wire [14-1:0] node2010;
	wire [14-1:0] node2011;
	wire [14-1:0] node2016;
	wire [14-1:0] node2017;
	wire [14-1:0] node2018;
	wire [14-1:0] node2020;
	wire [14-1:0] node2024;
	wire [14-1:0] node2026;
	wire [14-1:0] node2027;
	wire [14-1:0] node2033;
	wire [14-1:0] node2034;
	wire [14-1:0] node2035;
	wire [14-1:0] node2036;
	wire [14-1:0] node2037;
	wire [14-1:0] node2038;
	wire [14-1:0] node2039;
	wire [14-1:0] node2040;
	wire [14-1:0] node2041;
	wire [14-1:0] node2043;
	wire [14-1:0] node2046;
	wire [14-1:0] node2048;
	wire [14-1:0] node2051;
	wire [14-1:0] node2052;
	wire [14-1:0] node2053;
	wire [14-1:0] node2057;
	wire [14-1:0] node2058;
	wire [14-1:0] node2062;
	wire [14-1:0] node2063;
	wire [14-1:0] node2064;
	wire [14-1:0] node2067;
	wire [14-1:0] node2070;
	wire [14-1:0] node2071;
	wire [14-1:0] node2072;
	wire [14-1:0] node2076;
	wire [14-1:0] node2078;
	wire [14-1:0] node2081;
	wire [14-1:0] node2082;
	wire [14-1:0] node2083;
	wire [14-1:0] node2084;
	wire [14-1:0] node2085;
	wire [14-1:0] node2088;
	wire [14-1:0] node2091;
	wire [14-1:0] node2092;
	wire [14-1:0] node2095;
	wire [14-1:0] node2098;
	wire [14-1:0] node2099;
	wire [14-1:0] node2100;
	wire [14-1:0] node2103;
	wire [14-1:0] node2106;
	wire [14-1:0] node2108;
	wire [14-1:0] node2113;
	wire [14-1:0] node2114;
	wire [14-1:0] node2115;
	wire [14-1:0] node2116;
	wire [14-1:0] node2118;
	wire [14-1:0] node2119;
	wire [14-1:0] node2122;
	wire [14-1:0] node2125;
	wire [14-1:0] node2126;
	wire [14-1:0] node2127;
	wire [14-1:0] node2130;
	wire [14-1:0] node2133;
	wire [14-1:0] node2134;
	wire [14-1:0] node2137;
	wire [14-1:0] node2140;
	wire [14-1:0] node2141;
	wire [14-1:0] node2142;
	wire [14-1:0] node2143;
	wire [14-1:0] node2146;
	wire [14-1:0] node2149;
	wire [14-1:0] node2150;
	wire [14-1:0] node2153;
	wire [14-1:0] node2156;
	wire [14-1:0] node2157;
	wire [14-1:0] node2158;
	wire [14-1:0] node2161;
	wire [14-1:0] node2164;
	wire [14-1:0] node2165;
	wire [14-1:0] node2168;
	wire [14-1:0] node2171;
	wire [14-1:0] node2172;
	wire [14-1:0] node2173;
	wire [14-1:0] node2174;
	wire [14-1:0] node2175;
	wire [14-1:0] node2178;
	wire [14-1:0] node2181;
	wire [14-1:0] node2182;
	wire [14-1:0] node2185;
	wire [14-1:0] node2188;
	wire [14-1:0] node2189;
	wire [14-1:0] node2190;
	wire [14-1:0] node2193;
	wire [14-1:0] node2196;
	wire [14-1:0] node2197;
	wire [14-1:0] node2200;
	wire [14-1:0] node2204;
	wire [14-1:0] node2205;
	wire [14-1:0] node2206;
	wire [14-1:0] node2207;
	wire [14-1:0] node2208;
	wire [14-1:0] node2209;
	wire [14-1:0] node2210;
	wire [14-1:0] node2213;
	wire [14-1:0] node2214;
	wire [14-1:0] node2217;
	wire [14-1:0] node2220;
	wire [14-1:0] node2221;
	wire [14-1:0] node2223;
	wire [14-1:0] node2228;
	wire [14-1:0] node2230;
	wire [14-1:0] node2232;
	wire [14-1:0] node2233;
	wire [14-1:0] node2237;
	wire [14-1:0] node2238;
	wire [14-1:0] node2239;
	wire [14-1:0] node2240;
	wire [14-1:0] node2241;
	wire [14-1:0] node2242;
	wire [14-1:0] node2245;
	wire [14-1:0] node2248;
	wire [14-1:0] node2249;
	wire [14-1:0] node2253;
	wire [14-1:0] node2254;
	wire [14-1:0] node2255;
	wire [14-1:0] node2258;
	wire [14-1:0] node2263;
	wire [14-1:0] node2264;
	wire [14-1:0] node2265;
	wire [14-1:0] node2266;
	wire [14-1:0] node2269;
	wire [14-1:0] node2272;
	wire [14-1:0] node2273;
	wire [14-1:0] node2276;
	wire [14-1:0] node2279;
	wire [14-1:0] node2280;
	wire [14-1:0] node2281;
	wire [14-1:0] node2284;
	wire [14-1:0] node2289;
	wire [14-1:0] node2290;
	wire [14-1:0] node2291;
	wire [14-1:0] node2292;
	wire [14-1:0] node2293;
	wire [14-1:0] node2294;
	wire [14-1:0] node2295;
	wire [14-1:0] node2296;
	wire [14-1:0] node2298;
	wire [14-1:0] node2301;
	wire [14-1:0] node2302;
	wire [14-1:0] node2306;
	wire [14-1:0] node2307;
	wire [14-1:0] node2308;
	wire [14-1:0] node2311;
	wire [14-1:0] node2314;
	wire [14-1:0] node2315;
	wire [14-1:0] node2318;
	wire [14-1:0] node2321;
	wire [14-1:0] node2322;
	wire [14-1:0] node2323;
	wire [14-1:0] node2324;
	wire [14-1:0] node2328;
	wire [14-1:0] node2329;
	wire [14-1:0] node2332;
	wire [14-1:0] node2336;
	wire [14-1:0] node2338;
	wire [14-1:0] node2339;
	wire [14-1:0] node2340;
	wire [14-1:0] node2341;
	wire [14-1:0] node2344;
	wire [14-1:0] node2347;
	wire [14-1:0] node2350;
	wire [14-1:0] node2351;
	wire [14-1:0] node2352;
	wire [14-1:0] node2355;
	wire [14-1:0] node2359;
	wire [14-1:0] node2360;
	wire [14-1:0] node2362;
	wire [14-1:0] node2363;
	wire [14-1:0] node2364;
	wire [14-1:0] node2365;
	wire [14-1:0] node2368;
	wire [14-1:0] node2371;
	wire [14-1:0] node2372;
	wire [14-1:0] node2375;
	wire [14-1:0] node2378;
	wire [14-1:0] node2379;
	wire [14-1:0] node2381;
	wire [14-1:0] node2386;
	wire [14-1:0] node2387;
	wire [14-1:0] node2388;
	wire [14-1:0] node2389;
	wire [14-1:0] node2390;
	wire [14-1:0] node2392;
	wire [14-1:0] node2394;
	wire [14-1:0] node2398;
	wire [14-1:0] node2400;
	wire [14-1:0] node2401;
	wire [14-1:0] node2407;
	wire [14-1:0] node2408;
	wire [14-1:0] node2409;
	wire [14-1:0] node2411;
	wire [14-1:0] node2412;
	wire [14-1:0] node2414;
	wire [14-1:0] node2416;
	wire [14-1:0] node2417;
	wire [14-1:0] node2421;
	wire [14-1:0] node2422;
	wire [14-1:0] node2423;
	wire [14-1:0] node2425;
	wire [14-1:0] node2432;
	wire [14-1:0] node2433;
	wire [14-1:0] node2434;
	wire [14-1:0] node2435;
	wire [14-1:0] node2436;
	wire [14-1:0] node2437;
	wire [14-1:0] node2438;
	wire [14-1:0] node2439;
	wire [14-1:0] node2440;
	wire [14-1:0] node2442;
	wire [14-1:0] node2444;
	wire [14-1:0] node2447;
	wire [14-1:0] node2448;
	wire [14-1:0] node2449;
	wire [14-1:0] node2452;
	wire [14-1:0] node2455;
	wire [14-1:0] node2456;
	wire [14-1:0] node2459;
	wire [14-1:0] node2462;
	wire [14-1:0] node2464;
	wire [14-1:0] node2465;
	wire [14-1:0] node2468;
	wire [14-1:0] node2471;
	wire [14-1:0] node2472;
	wire [14-1:0] node2473;
	wire [14-1:0] node2474;
	wire [14-1:0] node2476;
	wire [14-1:0] node2479;
	wire [14-1:0] node2482;
	wire [14-1:0] node2483;
	wire [14-1:0] node2484;
	wire [14-1:0] node2487;
	wire [14-1:0] node2490;
	wire [14-1:0] node2493;
	wire [14-1:0] node2494;
	wire [14-1:0] node2495;
	wire [14-1:0] node2496;
	wire [14-1:0] node2499;
	wire [14-1:0] node2502;
	wire [14-1:0] node2505;
	wire [14-1:0] node2506;
	wire [14-1:0] node2509;
	wire [14-1:0] node2512;
	wire [14-1:0] node2513;
	wire [14-1:0] node2514;
	wire [14-1:0] node2515;
	wire [14-1:0] node2516;
	wire [14-1:0] node2517;
	wire [14-1:0] node2520;
	wire [14-1:0] node2523;
	wire [14-1:0] node2525;
	wire [14-1:0] node2528;
	wire [14-1:0] node2529;
	wire [14-1:0] node2532;
	wire [14-1:0] node2535;
	wire [14-1:0] node2536;
	wire [14-1:0] node2537;
	wire [14-1:0] node2538;
	wire [14-1:0] node2541;
	wire [14-1:0] node2544;
	wire [14-1:0] node2547;
	wire [14-1:0] node2548;
	wire [14-1:0] node2549;
	wire [14-1:0] node2552;
	wire [14-1:0] node2555;
	wire [14-1:0] node2558;
	wire [14-1:0] node2559;
	wire [14-1:0] node2560;
	wire [14-1:0] node2561;
	wire [14-1:0] node2563;
	wire [14-1:0] node2566;
	wire [14-1:0] node2569;
	wire [14-1:0] node2570;
	wire [14-1:0] node2572;
	wire [14-1:0] node2575;
	wire [14-1:0] node2578;
	wire [14-1:0] node2579;
	wire [14-1:0] node2580;
	wire [14-1:0] node2581;
	wire [14-1:0] node2585;
	wire [14-1:0] node2588;
	wire [14-1:0] node2589;
	wire [14-1:0] node2590;
	wire [14-1:0] node2593;
	wire [14-1:0] node2596;
	wire [14-1:0] node2599;
	wire [14-1:0] node2600;
	wire [14-1:0] node2601;
	wire [14-1:0] node2602;
	wire [14-1:0] node2603;
	wire [14-1:0] node2604;
	wire [14-1:0] node2605;
	wire [14-1:0] node2608;
	wire [14-1:0] node2611;
	wire [14-1:0] node2612;
	wire [14-1:0] node2615;
	wire [14-1:0] node2618;
	wire [14-1:0] node2619;
	wire [14-1:0] node2620;
	wire [14-1:0] node2623;
	wire [14-1:0] node2626;
	wire [14-1:0] node2627;
	wire [14-1:0] node2630;
	wire [14-1:0] node2633;
	wire [14-1:0] node2634;
	wire [14-1:0] node2635;
	wire [14-1:0] node2636;
	wire [14-1:0] node2639;
	wire [14-1:0] node2642;
	wire [14-1:0] node2643;
	wire [14-1:0] node2646;
	wire [14-1:0] node2649;
	wire [14-1:0] node2650;
	wire [14-1:0] node2651;
	wire [14-1:0] node2654;
	wire [14-1:0] node2657;
	wire [14-1:0] node2659;
	wire [14-1:0] node2662;
	wire [14-1:0] node2664;
	wire [14-1:0] node2665;
	wire [14-1:0] node2666;
	wire [14-1:0] node2667;
	wire [14-1:0] node2671;
	wire [14-1:0] node2672;
	wire [14-1:0] node2675;
	wire [14-1:0] node2678;
	wire [14-1:0] node2679;
	wire [14-1:0] node2680;
	wire [14-1:0] node2683;
	wire [14-1:0] node2686;
	wire [14-1:0] node2687;
	wire [14-1:0] node2691;
	wire [14-1:0] node2692;
	wire [14-1:0] node2693;
	wire [14-1:0] node2694;
	wire [14-1:0] node2696;
	wire [14-1:0] node2697;
	wire [14-1:0] node2700;
	wire [14-1:0] node2703;
	wire [14-1:0] node2704;
	wire [14-1:0] node2705;
	wire [14-1:0] node2708;
	wire [14-1:0] node2711;
	wire [14-1:0] node2712;
	wire [14-1:0] node2715;
	wire [14-1:0] node2720;
	wire [14-1:0] node2721;
	wire [14-1:0] node2722;
	wire [14-1:0] node2723;
	wire [14-1:0] node2724;
	wire [14-1:0] node2725;
	wire [14-1:0] node2726;
	wire [14-1:0] node2727;
	wire [14-1:0] node2730;
	wire [14-1:0] node2733;
	wire [14-1:0] node2734;
	wire [14-1:0] node2738;
	wire [14-1:0] node2739;
	wire [14-1:0] node2740;
	wire [14-1:0] node2744;
	wire [14-1:0] node2745;
	wire [14-1:0] node2748;
	wire [14-1:0] node2752;
	wire [14-1:0] node2753;
	wire [14-1:0] node2754;
	wire [14-1:0] node2755;
	wire [14-1:0] node2758;
	wire [14-1:0] node2761;
	wire [14-1:0] node2762;
	wire [14-1:0] node2765;
	wire [14-1:0] node2768;
	wire [14-1:0] node2769;
	wire [14-1:0] node2770;
	wire [14-1:0] node2773;
	wire [14-1:0] node2776;
	wire [14-1:0] node2777;
	wire [14-1:0] node2780;
	wire [14-1:0] node2783;
	wire [14-1:0] node2784;
	wire [14-1:0] node2785;
	wire [14-1:0] node2786;
	wire [14-1:0] node2787;
	wire [14-1:0] node2788;
	wire [14-1:0] node2791;
	wire [14-1:0] node2794;
	wire [14-1:0] node2796;
	wire [14-1:0] node2799;
	wire [14-1:0] node2801;
	wire [14-1:0] node2803;
	wire [14-1:0] node2806;
	wire [14-1:0] node2808;
	wire [14-1:0] node2810;
	wire [14-1:0] node2812;
	wire [14-1:0] node2816;
	wire [14-1:0] node2817;
	wire [14-1:0] node2818;
	wire [14-1:0] node2819;
	wire [14-1:0] node2820;
	wire [14-1:0] node2821;
	wire [14-1:0] node2822;
	wire [14-1:0] node2825;
	wire [14-1:0] node2828;
	wire [14-1:0] node2829;
	wire [14-1:0] node2832;
	wire [14-1:0] node2835;
	wire [14-1:0] node2837;
	wire [14-1:0] node2838;
	wire [14-1:0] node2842;
	wire [14-1:0] node2844;
	wire [14-1:0] node2845;
	wire [14-1:0] node2846;
	wire [14-1:0] node2849;
	wire [14-1:0] node2855;
	wire [14-1:0] node2856;
	wire [14-1:0] node2857;
	wire [14-1:0] node2858;
	wire [14-1:0] node2859;
	wire [14-1:0] node2861;
	wire [14-1:0] node2862;
	wire [14-1:0] node2863;
	wire [14-1:0] node2865;
	wire [14-1:0] node2868;
	wire [14-1:0] node2869;
	wire [14-1:0] node2877;
	wire [14-1:0] node2878;
	wire [14-1:0] node2879;
	wire [14-1:0] node2880;
	wire [14-1:0] node2881;
	wire [14-1:0] node2882;
	wire [14-1:0] node2883;
	wire [14-1:0] node2884;
	wire [14-1:0] node2887;
	wire [14-1:0] node2890;
	wire [14-1:0] node2893;
	wire [14-1:0] node2894;
	wire [14-1:0] node2895;
	wire [14-1:0] node2899;
	wire [14-1:0] node2901;
	wire [14-1:0] node2904;
	wire [14-1:0] node2905;
	wire [14-1:0] node2906;
	wire [14-1:0] node2907;
	wire [14-1:0] node2910;
	wire [14-1:0] node2913;
	wire [14-1:0] node2916;
	wire [14-1:0] node2917;
	wire [14-1:0] node2918;
	wire [14-1:0] node2922;
	wire [14-1:0] node2924;
	wire [14-1:0] node2927;
	wire [14-1:0] node2928;
	wire [14-1:0] node2929;
	wire [14-1:0] node2930;
	wire [14-1:0] node2931;
	wire [14-1:0] node2934;
	wire [14-1:0] node2938;
	wire [14-1:0] node2939;
	wire [14-1:0] node2942;
	wire [14-1:0] node2945;
	wire [14-1:0] node2946;
	wire [14-1:0] node2947;
	wire [14-1:0] node2948;
	wire [14-1:0] node2954;
	wire [14-1:0] node2955;
	wire [14-1:0] node2956;
	wire [14-1:0] node2957;
	wire [14-1:0] node2958;
	wire [14-1:0] node2959;
	wire [14-1:0] node2962;
	wire [14-1:0] node2965;
	wire [14-1:0] node2967;
	wire [14-1:0] node2970;
	wire [14-1:0] node2971;
	wire [14-1:0] node2972;
	wire [14-1:0] node2975;
	wire [14-1:0] node2979;
	wire [14-1:0] node2981;
	wire [14-1:0] node2982;
	wire [14-1:0] node2984;
	wire [14-1:0] node2988;
	wire [14-1:0] node2989;
	wire [14-1:0] node2990;
	wire [14-1:0] node2991;
	wire [14-1:0] node2993;
	wire [14-1:0] node2996;
	wire [14-1:0] node3002;
	wire [14-1:0] node3003;
	wire [14-1:0] node3004;
	wire [14-1:0] node3005;
	wire [14-1:0] node3006;
	wire [14-1:0] node3007;
	wire [14-1:0] node3008;
	wire [14-1:0] node3010;
	wire [14-1:0] node3011;
	wire [14-1:0] node3012;
	wire [14-1:0] node3015;
	wire [14-1:0] node3019;
	wire [14-1:0] node3020;
	wire [14-1:0] node3021;
	wire [14-1:0] node3023;
	wire [14-1:0] node3032;
	wire [14-1:0] node3033;
	wire [14-1:0] node3034;
	wire [14-1:0] node3035;
	wire [14-1:0] node3036;
	wire [14-1:0] node3037;
	wire [14-1:0] node3039;
	wire [14-1:0] node3040;
	wire [14-1:0] node3044;
	wire [14-1:0] node3046;
	wire [14-1:0] node3047;
	wire [14-1:0] node3054;
	wire [14-1:0] node3055;
	wire [14-1:0] node3056;
	wire [14-1:0] node3057;
	wire [14-1:0] node3058;
	wire [14-1:0] node3059;
	wire [14-1:0] node3061;
	wire [14-1:0] node3068;
	wire [14-1:0] node3069;
	wire [14-1:0] node3070;
	wire [14-1:0] node3071;
	wire [14-1:0] node3072;
	wire [14-1:0] node3073;
	wire [14-1:0] node3080;
	wire [14-1:0] node3082;
	wire [14-1:0] node3084;
	wire [14-1:0] node3086;
	wire [14-1:0] node3087;
	wire [14-1:0] node3090;

	assign outp = (inp[13]) ? node1180 : node1;
		assign node1 = (inp[8]) ? node3 : 14'b00000000000000;
			assign node3 = (inp[0]) ? node789 : node4;
				assign node4 = (inp[11]) ? node540 : node5;
					assign node5 = (inp[3]) ? node351 : node6;
						assign node6 = (inp[2]) ? node200 : node7;
							assign node7 = (inp[12]) ? node121 : node8;
								assign node8 = (inp[1]) ? node68 : node9;
									assign node9 = (inp[6]) ? node39 : node10;
										assign node10 = (inp[7]) ? node24 : node11;
											assign node11 = (inp[9]) ? node17 : node12;
												assign node12 = (inp[4]) ? 14'b00000000000001 : node13;
													assign node13 = (inp[10]) ? 14'b00000000000001 : 14'b10000000001000;
												assign node17 = (inp[5]) ? node21 : node18;
													assign node18 = (inp[4]) ? 14'b01101100000000 : 14'b01101100000010;
													assign node21 = (inp[4]) ? 14'b01100100000000 : 14'b00100100000010;
											assign node24 = (inp[10]) ? node32 : node25;
												assign node25 = (inp[4]) ? node29 : node26;
													assign node26 = (inp[5]) ? 14'b00100110010010 : 14'b00000000000001;
													assign node29 = (inp[9]) ? 14'b01100110010110 : 14'b01100110110110;
												assign node32 = (inp[9]) ? node36 : node33;
													assign node33 = (inp[5]) ? 14'b01100110110000 : 14'b01101110110000;
													assign node36 = (inp[5]) ? 14'b01100110010000 : 14'b01101110010000;
										assign node39 = (inp[9]) ? node55 : node40;
											assign node40 = (inp[5]) ? node48 : node41;
												assign node41 = (inp[10]) ? node45 : node42;
													assign node42 = (inp[7]) ? 14'b01101100110110 : 14'b01111100110110;
													assign node45 = (inp[4]) ? 14'b01101100110000 : 14'b01101100110010;
												assign node48 = (inp[7]) ? node52 : node49;
													assign node49 = (inp[10]) ? 14'b01110100110000 : 14'b00110100110010;
													assign node52 = (inp[4]) ? 14'b01100100110000 : 14'b00100100110010;
											assign node55 = (inp[7]) ? node61 : node56;
												assign node56 = (inp[5]) ? 14'b01110100010010 : node57;
													assign node57 = (inp[10]) ? 14'b01111100010000 : 14'b01111100010110;
												assign node61 = (inp[4]) ? node65 : node62;
													assign node62 = (inp[10]) ? 14'b01101100010010 : 14'b00000000000001;
													assign node65 = (inp[10]) ? 14'b01100100010000 : 14'b01100100010110;
									assign node68 = (inp[4]) ? node90 : node69;
										assign node69 = (inp[10]) ? node79 : node70;
											assign node70 = (inp[5]) ? node72 : 14'b00000000000001;
												assign node72 = (inp[6]) ? node76 : node73;
													assign node73 = (inp[9]) ? 14'b00100010010010 : 14'b00110010000010;
													assign node76 = (inp[7]) ? 14'b00100000010010 : 14'b00110000010010;
											assign node79 = (inp[6]) ? node85 : node80;
												assign node80 = (inp[7]) ? 14'b01101010110010 : node81;
													assign node81 = (inp[9]) ? 14'b01101000000010 : 14'b01111010000010;
												assign node85 = (inp[5]) ? 14'b01110000110010 : node86;
													assign node86 = (inp[7]) ? 14'b01101000110010 : 14'b01111000110010;
										assign node90 = (inp[10]) ? node106 : node91;
											assign node91 = (inp[7]) ? node99 : node92;
												assign node92 = (inp[9]) ? node96 : node93;
													assign node93 = (inp[5]) ? 14'b01110010000110 : 14'b01111010000110;
													assign node96 = (inp[6]) ? 14'b01110000010110 : 14'b01100000000110;
												assign node99 = (inp[5]) ? node103 : node100;
													assign node100 = (inp[6]) ? 14'b01101000010110 : 14'b01101010010110;
													assign node103 = (inp[6]) ? 14'b01100000110110 : 14'b01100010010110;
											assign node106 = (inp[7]) ? node114 : node107;
												assign node107 = (inp[6]) ? node111 : node108;
													assign node108 = (inp[9]) ? 14'b01100000000000 : 14'b01110010000000;
													assign node111 = (inp[5]) ? 14'b01110000010000 : 14'b01111000010000;
												assign node114 = (inp[5]) ? node118 : node115;
													assign node115 = (inp[9]) ? 14'b01101000010000 : 14'b01101010110000;
													assign node118 = (inp[6]) ? 14'b01100000110000 : 14'b01100010110000;
								assign node121 = (inp[4]) ? node169 : node122;
									assign node122 = (inp[10]) ? node154 : node123;
										assign node123 = (inp[6]) ? node139 : node124;
											assign node124 = (inp[7]) ? node132 : node125;
												assign node125 = (inp[9]) ? node129 : node126;
													assign node126 = (inp[1]) ? 14'b01011010000110 : 14'b00000000000001;
													assign node129 = (inp[1]) ? 14'b01000000000110 : 14'b01000100000110;
												assign node132 = (inp[5]) ? node136 : node133;
													assign node133 = (inp[1]) ? 14'b01001010010110 : 14'b01001110010110;
													assign node136 = (inp[9]) ? 14'b01000010010110 : 14'b01000010110110;
											assign node139 = (inp[5]) ? node147 : node140;
												assign node140 = (inp[7]) ? node144 : node141;
													assign node141 = (inp[9]) ? 14'b01011100010110 : 14'b01011000110110;
													assign node144 = (inp[9]) ? 14'b01001000010110 : 14'b01001100110110;
												assign node147 = (inp[1]) ? node151 : node148;
													assign node148 = (inp[9]) ? 14'b01000100010110 : 14'b01010100110110;
													assign node151 = (inp[9]) ? 14'b01010000010110 : 14'b01010000110110;
										assign node154 = (inp[5]) ? 14'b00000000000001 : node155;
											assign node155 = (inp[6]) ? node161 : node156;
												assign node156 = (inp[7]) ? 14'b01001110010010 : node157;
													assign node157 = (inp[1]) ? 14'b01001000000010 : 14'b00000000000001;
												assign node161 = (inp[1]) ? node165 : node162;
													assign node162 = (inp[7]) ? 14'b01001100010010 : 14'b01011100010010;
													assign node165 = (inp[9]) ? 14'b01011000010010 : 14'b01011000110010;
									assign node169 = (inp[5]) ? node183 : node170;
										assign node170 = (inp[10]) ? node172 : 14'b00000000000001;
											assign node172 = (inp[9]) ? node178 : node173;
												assign node173 = (inp[1]) ? node175 : 14'b00000000000001;
													assign node175 = (inp[7]) ? 14'b00101010110000 : 14'b00111000000000;
												assign node178 = (inp[1]) ? 14'b00101000010000 : node179;
													assign node179 = (inp[6]) ? 14'b00101100010000 : 14'b00101100000000;
										assign node183 = (inp[10]) ? 14'b00000000000001 : node184;
											assign node184 = (inp[7]) ? node192 : node185;
												assign node185 = (inp[6]) ? node189 : node186;
													assign node186 = (inp[1]) ? 14'b01000000000010 : 14'b00000000000000;
													assign node189 = (inp[9]) ? 14'b01010100010010 : 14'b01010100110010;
												assign node192 = (inp[1]) ? node196 : node193;
													assign node193 = (inp[9]) ? 14'b01000100010010 : 14'b01000100110010;
													assign node196 = (inp[6]) ? 14'b01000000110010 : 14'b01000010110010;
							assign node200 = (inp[4]) ? node308 : node201;
								assign node201 = (inp[5]) ? node259 : node202;
									assign node202 = (inp[7]) ? node230 : node203;
										assign node203 = (inp[6]) ? node217 : node204;
											assign node204 = (inp[1]) ? node210 : node205;
												assign node205 = (inp[9]) ? node207 : 14'b00000000000001;
													assign node207 = (inp[10]) ? 14'b00001100000010 : 14'b00001100000110;
												assign node210 = (inp[9]) ? node214 : node211;
													assign node211 = (inp[12]) ? 14'b00011010000010 : 14'b00011010000000;
													assign node214 = (inp[10]) ? 14'b00001000000010 : 14'b00001000000110;
											assign node217 = (inp[10]) ? node223 : node218;
												assign node218 = (inp[9]) ? node220 : 14'b00011000110000;
													assign node220 = (inp[1]) ? 14'b00011000010000 : 14'b00011100010000;
												assign node223 = (inp[9]) ? node227 : node224;
													assign node224 = (inp[1]) ? 14'b00111000110010 : 14'b00111100110010;
													assign node227 = (inp[1]) ? 14'b00011000010010 : 14'b00011100010010;
										assign node230 = (inp[6]) ? node244 : node231;
											assign node231 = (inp[1]) ? node237 : node232;
												assign node232 = (inp[12]) ? node234 : 14'b00001110110000;
													assign node234 = (inp[9]) ? 14'b00001110010110 : 14'b00001110110010;
												assign node237 = (inp[9]) ? node241 : node238;
													assign node238 = (inp[10]) ? 14'b00001010110010 : 14'b00001010110000;
													assign node241 = (inp[12]) ? 14'b00001010010010 : 14'b00001010010000;
											assign node244 = (inp[1]) ? node252 : node245;
												assign node245 = (inp[9]) ? node249 : node246;
													assign node246 = (inp[10]) ? 14'b00001100110010 : 14'b00001100110000;
													assign node249 = (inp[10]) ? 14'b00001100010010 : 14'b00001100010000;
												assign node252 = (inp[9]) ? node256 : node253;
													assign node253 = (inp[10]) ? 14'b00001000110010 : 14'b00001000110110;
													assign node256 = (inp[12]) ? 14'b00001000010010 : 14'b00001000010000;
									assign node259 = (inp[12]) ? node277 : node260;
										assign node260 = (inp[10]) ? 14'b00000000000001 : node261;
											assign node261 = (inp[7]) ? node269 : node262;
												assign node262 = (inp[6]) ? node266 : node263;
													assign node263 = (inp[9]) ? 14'b00000000000000 : 14'b00000000000001;
													assign node266 = (inp[1]) ? 14'b00010000010000 : 14'b00010100010000;
												assign node269 = (inp[9]) ? node273 : node270;
													assign node270 = (inp[1]) ? 14'b00000010110000 : 14'b00000100110000;
													assign node273 = (inp[6]) ? 14'b00000000010000 : 14'b00000010010000;
										assign node277 = (inp[7]) ? node293 : node278;
											assign node278 = (inp[6]) ? node286 : node279;
												assign node279 = (inp[9]) ? node283 : node280;
													assign node280 = (inp[1]) ? 14'b00010010000110 : 14'b00000000000001;
													assign node283 = (inp[1]) ? 14'b00000000000010 : 14'b00000100000010;
												assign node286 = (inp[10]) ? node290 : node287;
													assign node287 = (inp[9]) ? 14'b00010000010110 : 14'b00010100110110;
													assign node290 = (inp[9]) ? 14'b00010000010010 : 14'b00010000110010;
											assign node293 = (inp[6]) ? node301 : node294;
												assign node294 = (inp[9]) ? node298 : node295;
													assign node295 = (inp[1]) ? 14'b00000010110010 : 14'b00000110110010;
													assign node298 = (inp[10]) ? 14'b00000010010010 : 14'b00000110010110;
												assign node301 = (inp[1]) ? node305 : node302;
													assign node302 = (inp[10]) ? 14'b00000100110010 : 14'b00000100010110;
													assign node305 = (inp[9]) ? 14'b00000000010010 : 14'b00000000110110;
								assign node308 = (inp[12]) ? 14'b00000000000001 : node309;
									assign node309 = (inp[10]) ? node335 : node310;
										assign node310 = (inp[9]) ? node322 : node311;
											assign node311 = (inp[7]) ? node317 : node312;
												assign node312 = (inp[1]) ? 14'b00111000110110 : node313;
													assign node313 = (inp[5]) ? 14'b00110100110110 : 14'b00111100110110;
												assign node317 = (inp[6]) ? 14'b00100100110110 : node318;
													assign node318 = (inp[5]) ? 14'b00100110110110 : 14'b00101110110110;
											assign node322 = (inp[5]) ? node330 : node323;
												assign node323 = (inp[1]) ? node327 : node324;
													assign node324 = (inp[7]) ? 14'b00101100010110 : 14'b00101100000110;
													assign node327 = (inp[6]) ? 14'b00101000010110 : 14'b00101000000110;
												assign node330 = (inp[1]) ? node332 : 14'b00100110010110;
													assign node332 = (inp[6]) ? 14'b00100000010110 : 14'b00100010010110;
										assign node335 = (inp[5]) ? node337 : 14'b00000000000001;
											assign node337 = (inp[1]) ? node345 : node338;
												assign node338 = (inp[9]) ? node342 : node339;
													assign node339 = (inp[6]) ? 14'b00100100110000 : 14'b00100110110000;
													assign node342 = (inp[6]) ? 14'b00100100010000 : 14'b00100100000000;
												assign node345 = (inp[9]) ? 14'b00100010010000 : node346;
													assign node346 = (inp[6]) ? 14'b00100000110000 : 14'b00100010110000;
						assign node351 = (inp[7]) ? node483 : node352;
							assign node352 = (inp[6]) ? node450 : node353;
								assign node353 = (inp[12]) ? node407 : node354;
									assign node354 = (inp[2]) ? node384 : node355;
										assign node355 = (inp[9]) ? node371 : node356;
											assign node356 = (inp[1]) ? node364 : node357;
												assign node357 = (inp[5]) ? node361 : node358;
													assign node358 = (inp[10]) ? 14'b01111110110000 : 14'b01111110110110;
													assign node361 = (inp[10]) ? 14'b01110110110000 : 14'b00110110110010;
												assign node364 = (inp[5]) ? node368 : node365;
													assign node365 = (inp[4]) ? 14'b01111010110110 : 14'b01111010110010;
													assign node368 = (inp[4]) ? 14'b01110010110110 : 14'b00110010110010;
											assign node371 = (inp[4]) ? node377 : node372;
												assign node372 = (inp[5]) ? node374 : 14'b00000000000001;
													assign node374 = (inp[10]) ? 14'b01110010010010 : 14'b00110010010010;
												assign node377 = (inp[10]) ? node381 : node378;
													assign node378 = (inp[5]) ? 14'b01110110010110 : 14'b01111010010110;
													assign node381 = (inp[1]) ? 14'b01110010010000 : 14'b01110110010000;
										assign node384 = (inp[10]) ? node398 : node385;
											assign node385 = (inp[4]) ? node393 : node386;
												assign node386 = (inp[1]) ? node390 : node387;
													assign node387 = (inp[9]) ? 14'b00010110010000 : 14'b00010110110000;
													assign node390 = (inp[5]) ? 14'b00010010110000 : 14'b00011010110000;
												assign node393 = (inp[5]) ? 14'b00110010010110 : node394;
													assign node394 = (inp[1]) ? 14'b00111010110110 : 14'b00111110010110;
											assign node398 = (inp[9]) ? node404 : node399;
												assign node399 = (inp[1]) ? node401 : 14'b00000000000001;
													assign node401 = (inp[4]) ? 14'b00000000000001 : 14'b00111010110010;
												assign node404 = (inp[4]) ? 14'b00110010010000 : 14'b00111110010010;
									assign node407 = (inp[4]) ? node435 : node408;
										assign node408 = (inp[5]) ? node422 : node409;
											assign node409 = (inp[2]) ? node417 : node410;
												assign node410 = (inp[9]) ? node414 : node411;
													assign node411 = (inp[1]) ? 14'b01011010110010 : 14'b01011110110010;
													assign node414 = (inp[10]) ? 14'b01011010010010 : 14'b01011010010110;
												assign node417 = (inp[10]) ? 14'b00011110010010 : node418;
													assign node418 = (inp[1]) ? 14'b00011010010110 : 14'b00011110010110;
											assign node422 = (inp[10]) ? node430 : node423;
												assign node423 = (inp[2]) ? node427 : node424;
													assign node424 = (inp[1]) ? 14'b01010010010110 : 14'b01010110010110;
													assign node427 = (inp[1]) ? 14'b00010010010110 : 14'b00010110110110;
												assign node430 = (inp[2]) ? node432 : 14'b00000000000001;
													assign node432 = (inp[9]) ? 14'b00010110010010 : 14'b00010110110010;
										assign node435 = (inp[2]) ? 14'b00000000000001 : node436;
											assign node436 = (inp[9]) ? node442 : node437;
												assign node437 = (inp[10]) ? node439 : 14'b01010010110010;
													assign node439 = (inp[1]) ? 14'b00111010110000 : 14'b00111110110000;
												assign node442 = (inp[5]) ? node446 : node443;
													assign node443 = (inp[10]) ? 14'b00111010010000 : 14'b00000000000001;
													assign node446 = (inp[10]) ? 14'b00000000000001 : 14'b01010110010010;
								assign node450 = (inp[9]) ? 14'b00000000000001 : node451;
									assign node451 = (inp[1]) ? node453 : 14'b00000000000001;
										assign node453 = (inp[5]) ? node467 : node454;
											assign node454 = (inp[4]) ? node462 : node455;
												assign node455 = (inp[10]) ? node459 : node456;
													assign node456 = (inp[12]) ? 14'b00011000100110 : 14'b00000000000000;
													assign node459 = (inp[2]) ? 14'b00011000100010 : 14'b01011000100010;
												assign node462 = (inp[2]) ? 14'b00000000000001 : node463;
													assign node463 = (inp[12]) ? 14'b00000000000000 : 14'b01111000100110;
											assign node467 = (inp[10]) ? node475 : node468;
												assign node468 = (inp[4]) ? node472 : node469;
													assign node469 = (inp[2]) ? 14'b00010000100000 : 14'b00110000100010;
													assign node472 = (inp[12]) ? 14'b01010000100010 : 14'b00110000100110;
												assign node475 = (inp[12]) ? node479 : node476;
													assign node476 = (inp[2]) ? 14'b00000000000000 : 14'b01110000100000;
													assign node479 = (inp[2]) ? 14'b00010000100010 : 14'b00000000000001;
							assign node483 = (inp[9]) ? 14'b00000000000001 : node484;
								assign node484 = (inp[6]) ? node486 : 14'b00000000000001;
									assign node486 = (inp[12]) ? node516 : node487;
										assign node487 = (inp[4]) ? node501 : node488;
											assign node488 = (inp[10]) ? node496 : node489;
												assign node489 = (inp[2]) ? node493 : node490;
													assign node490 = (inp[5]) ? 14'b00100100100010 : 14'b00000000000001;
													assign node493 = (inp[5]) ? 14'b00000000100000 : 14'b00001000100000;
												assign node496 = (inp[5]) ? 14'b00000000000001 : node497;
													assign node497 = (inp[2]) ? 14'b00101000100010 : 14'b01101000100010;
											assign node501 = (inp[10]) ? node509 : node502;
												assign node502 = (inp[2]) ? node506 : node503;
													assign node503 = (inp[1]) ? 14'b01100000100110 : 14'b01100100100110;
													assign node506 = (inp[1]) ? 14'b00100000100110 : 14'b00101100100110;
												assign node509 = (inp[1]) ? node513 : node510;
													assign node510 = (inp[5]) ? 14'b01100100100000 : 14'b01101100100000;
													assign node513 = (inp[5]) ? 14'b00100000100000 : 14'b01101000100000;
										assign node516 = (inp[4]) ? node532 : node517;
											assign node517 = (inp[5]) ? node525 : node518;
												assign node518 = (inp[2]) ? node522 : node519;
													assign node519 = (inp[10]) ? 14'b01001000100010 : 14'b01001000100110;
													assign node522 = (inp[10]) ? 14'b00001000100010 : 14'b00001000100110;
												assign node525 = (inp[10]) ? node529 : node526;
													assign node526 = (inp[2]) ? 14'b00000000100110 : 14'b01000000100110;
													assign node529 = (inp[2]) ? 14'b00000100100010 : 14'b00000000000001;
											assign node532 = (inp[2]) ? 14'b00000000000001 : node533;
												assign node533 = (inp[1]) ? node535 : 14'b01000100100010;
													assign node535 = (inp[10]) ? 14'b00000000000000 : 14'b00000000000000;
					assign node540 = (inp[10]) ? 14'b00000000000001 : node541;
						assign node541 = (inp[4]) ? node721 : node542;
							assign node542 = (inp[3]) ? node658 : node543;
								assign node543 = (inp[6]) ? node597 : node544;
									assign node544 = (inp[7]) ? node566 : node545;
										assign node545 = (inp[9]) ? node555 : node546;
											assign node546 = (inp[1]) ? node548 : 14'b00000000000001;
												assign node548 = (inp[12]) ? node552 : node549;
													assign node549 = (inp[5]) ? 14'b00110010000100 : 14'b01111010000100;
													assign node552 = (inp[5]) ? 14'b00010010000100 : 14'b00011010000100;
											assign node555 = (inp[1]) ? node561 : node556;
												assign node556 = (inp[5]) ? 14'b00100100000100 : node557;
													assign node557 = (inp[2]) ? 14'b00101100000100 : 14'b01101100000100;
												assign node561 = (inp[2]) ? node563 : 14'b01000000000100;
													assign node563 = (inp[12]) ? 14'b00001000000100 : 14'b00100000000100;
										assign node566 = (inp[1]) ? node582 : node567;
											assign node567 = (inp[5]) ? node575 : node568;
												assign node568 = (inp[12]) ? node572 : node569;
													assign node569 = (inp[9]) ? 14'b00101110010100 : 14'b00101110110100;
													assign node572 = (inp[9]) ? 14'b00001110010100 : 14'b01001110110100;
												assign node575 = (inp[12]) ? node579 : node576;
													assign node576 = (inp[2]) ? 14'b00100110010100 : 14'b01100110010100;
													assign node579 = (inp[9]) ? 14'b00000110010100 : 14'b00000110110100;
											assign node582 = (inp[2]) ? node590 : node583;
												assign node583 = (inp[5]) ? node587 : node584;
													assign node584 = (inp[12]) ? 14'b01001010110100 : 14'b01101010110100;
													assign node587 = (inp[9]) ? 14'b01000010010100 : 14'b01100010110100;
												assign node590 = (inp[5]) ? node594 : node591;
													assign node591 = (inp[12]) ? 14'b00001010010100 : 14'b00101010010100;
													assign node594 = (inp[12]) ? 14'b00000010110100 : 14'b00100010010100;
									assign node597 = (inp[9]) ? node629 : node598;
										assign node598 = (inp[2]) ? node614 : node599;
											assign node599 = (inp[5]) ? node607 : node600;
												assign node600 = (inp[7]) ? node604 : node601;
													assign node601 = (inp[1]) ? 14'b01011000110100 : 14'b01011100110100;
													assign node604 = (inp[1]) ? 14'b01001000110100 : 14'b01001100110100;
												assign node607 = (inp[1]) ? node611 : node608;
													assign node608 = (inp[7]) ? 14'b01000100110100 : 14'b01010100110100;
													assign node611 = (inp[7]) ? 14'b01000000110100 : 14'b01010000110100;
											assign node614 = (inp[5]) ? node622 : node615;
												assign node615 = (inp[12]) ? node619 : node616;
													assign node616 = (inp[7]) ? 14'b00101100110100 : 14'b00111000110100;
													assign node619 = (inp[7]) ? 14'b00001000110100 : 14'b00011000110100;
												assign node622 = (inp[7]) ? node626 : node623;
													assign node623 = (inp[1]) ? 14'b00110000110100 : 14'b00010100110100;
													assign node626 = (inp[12]) ? 14'b00000100110100 : 14'b00100100110100;
										assign node629 = (inp[1]) ? node645 : node630;
											assign node630 = (inp[7]) ? node638 : node631;
												assign node631 = (inp[2]) ? node635 : node632;
													assign node632 = (inp[12]) ? 14'b01010100010100 : 14'b01110100010100;
													assign node635 = (inp[5]) ? 14'b00010100010100 : 14'b00011100010100;
												assign node638 = (inp[5]) ? node642 : node639;
													assign node639 = (inp[2]) ? 14'b00001100010100 : 14'b01001100010100;
													assign node642 = (inp[12]) ? 14'b00000100010100 : 14'b00100100010100;
											assign node645 = (inp[12]) ? node651 : node646;
												assign node646 = (inp[5]) ? node648 : 14'b01111000010100;
													assign node648 = (inp[2]) ? 14'b00110000010100 : 14'b01100000010100;
												assign node651 = (inp[5]) ? node655 : node652;
													assign node652 = (inp[7]) ? 14'b01001000010100 : 14'b01011000010100;
													assign node655 = (inp[2]) ? 14'b00000000010100 : 14'b01000000010100;
								assign node658 = (inp[7]) ? node702 : node659;
									assign node659 = (inp[6]) ? node691 : node660;
										assign node660 = (inp[5]) ? node676 : node661;
											assign node661 = (inp[1]) ? node669 : node662;
												assign node662 = (inp[12]) ? node666 : node663;
													assign node663 = (inp[9]) ? 14'b00111110010100 : 14'b00111110110100;
													assign node666 = (inp[9]) ? 14'b00011110010100 : 14'b00011110110100;
												assign node669 = (inp[9]) ? node673 : node670;
													assign node670 = (inp[2]) ? 14'b00011010110100 : 14'b01111010110100;
													assign node673 = (inp[12]) ? 14'b01011010010100 : 14'b00111010010100;
											assign node676 = (inp[1]) ? node684 : node677;
												assign node677 = (inp[12]) ? node681 : node678;
													assign node678 = (inp[9]) ? 14'b01110110010100 : 14'b01110110110100;
													assign node681 = (inp[2]) ? 14'b00010110010100 : 14'b01010110010100;
												assign node684 = (inp[9]) ? node688 : node685;
													assign node685 = (inp[2]) ? 14'b00010010110100 : 14'b01010010110100;
													assign node688 = (inp[2]) ? 14'b00010010010100 : 14'b01010010010100;
										assign node691 = (inp[9]) ? 14'b00000000000001 : node692;
											assign node692 = (inp[1]) ? node694 : 14'b00000000000001;
												assign node694 = (inp[12]) ? node698 : node695;
													assign node695 = (inp[2]) ? 14'b00110000100100 : 14'b01111000100100;
													assign node698 = (inp[5]) ? 14'b00010000100100 : 14'b00011000100100;
									assign node702 = (inp[6]) ? node704 : 14'b00000000000001;
										assign node704 = (inp[9]) ? 14'b00000000000001 : node705;
											assign node705 = (inp[2]) ? node713 : node706;
												assign node706 = (inp[1]) ? node710 : node707;
													assign node707 = (inp[12]) ? 14'b01000100100100 : 14'b01100100100100;
													assign node710 = (inp[12]) ? 14'b01001000100100 : 14'b01101000100100;
												assign node713 = (inp[5]) ? node717 : node714;
													assign node714 = (inp[1]) ? 14'b00101000100100 : 14'b00101100100100;
													assign node717 = (inp[12]) ? 14'b00000000100100 : 14'b00100000100100;
							assign node721 = (inp[2]) ? 14'b00000000000001 : node722;
								assign node722 = (inp[12]) ? node734 : node723;
									assign node723 = (inp[3]) ? node725 : 14'b00000000000001;
										assign node725 = (inp[1]) ? 14'b00000000000001 : node726;
											assign node726 = (inp[9]) ? 14'b00000000000001 : node727;
												assign node727 = (inp[5]) ? 14'b00000000000001 : node728;
													assign node728 = (inp[6]) ? 14'b10000001001000 : 14'b00000000000000;
									assign node734 = (inp[7]) ? node764 : node735;
										assign node735 = (inp[1]) ? node749 : node736;
											assign node736 = (inp[3]) ? node744 : node737;
												assign node737 = (inp[6]) ? node741 : node738;
													assign node738 = (inp[9]) ? 14'b01000100000000 : 14'b00000000000001;
													assign node741 = (inp[5]) ? 14'b01010100010000 : 14'b01011100010000;
												assign node744 = (inp[6]) ? 14'b00000000000001 : node745;
													assign node745 = (inp[9]) ? 14'b01010110010000 : 14'b01010110110000;
											assign node749 = (inp[6]) ? node757 : node750;
												assign node750 = (inp[3]) ? node754 : node751;
													assign node751 = (inp[9]) ? 14'b01000000000000 : 14'b01010010000000;
													assign node754 = (inp[5]) ? 14'b01010010010000 : 14'b01011010010000;
												assign node757 = (inp[9]) ? node761 : node758;
													assign node758 = (inp[5]) ? 14'b01010000100000 : 14'b01011000100000;
													assign node761 = (inp[3]) ? 14'b00000000000001 : 14'b01010000010000;
										assign node764 = (inp[3]) ? node780 : node765;
											assign node765 = (inp[9]) ? node773 : node766;
												assign node766 = (inp[6]) ? node770 : node767;
													assign node767 = (inp[5]) ? 14'b01000010110000 : 14'b01001010110000;
													assign node770 = (inp[5]) ? 14'b01000000110000 : 14'b01001000110000;
												assign node773 = (inp[1]) ? node777 : node774;
													assign node774 = (inp[6]) ? 14'b01000100010000 : 14'b01001110010000;
													assign node777 = (inp[5]) ? 14'b01000000010000 : 14'b01001000010000;
											assign node780 = (inp[6]) ? node782 : 14'b00000000000001;
												assign node782 = (inp[9]) ? 14'b00000000000001 : node783;
													assign node783 = (inp[1]) ? 14'b01001000100000 : 14'b01000100100000;
				assign node789 = (inp[7]) ? 14'b00000000000001 : node790;
					assign node790 = (inp[10]) ? node1046 : node791;
						assign node791 = (inp[1]) ? node939 : node792;
							assign node792 = (inp[3]) ? node886 : node793;
								assign node793 = (inp[4]) ? node853 : node794;
									assign node794 = (inp[12]) ? node824 : node795;
										assign node795 = (inp[11]) ? node809 : node796;
											assign node796 = (inp[5]) ? node802 : node797;
												assign node797 = (inp[2]) ? node799 : 14'b00000000000001;
													assign node799 = (inp[9]) ? 14'b00011110000000 : 14'b00011100100000;
												assign node802 = (inp[2]) ? node806 : node803;
													assign node803 = (inp[6]) ? 14'b00110100000010 : 14'b00110110000010;
													assign node806 = (inp[9]) ? 14'b00010110000000 : 14'b00010110100000;
											assign node809 = (inp[6]) ? node817 : node810;
												assign node810 = (inp[5]) ? node814 : node811;
													assign node811 = (inp[9]) ? 14'b01111110000100 : 14'b00111110100100;
													assign node814 = (inp[2]) ? 14'b00110110000100 : 14'b01110110000100;
												assign node817 = (inp[2]) ? node821 : node818;
													assign node818 = (inp[5]) ? 14'b01110100100100 : 14'b01111100100100;
													assign node821 = (inp[5]) ? 14'b00110100000100 : 14'b00111100000100;
										assign node824 = (inp[2]) ? node840 : node825;
											assign node825 = (inp[6]) ? node833 : node826;
												assign node826 = (inp[9]) ? node830 : node827;
													assign node827 = (inp[5]) ? 14'b01010110100110 : 14'b01011110100110;
													assign node830 = (inp[5]) ? 14'b01010110000100 : 14'b01011110000110;
												assign node833 = (inp[5]) ? node837 : node834;
													assign node834 = (inp[11]) ? 14'b01011100000100 : 14'b01011100000110;
													assign node837 = (inp[9]) ? 14'b01010100000110 : 14'b01010100100100;
											assign node840 = (inp[5]) ? node848 : node841;
												assign node841 = (inp[6]) ? node845 : node842;
													assign node842 = (inp[11]) ? 14'b00011110100100 : 14'b00011110100110;
													assign node845 = (inp[9]) ? 14'b00011100000100 : 14'b00011100100100;
												assign node848 = (inp[11]) ? node850 : 14'b00010110000110;
													assign node850 = (inp[6]) ? 14'b00010100000100 : 14'b00010110000100;
									assign node853 = (inp[11]) ? node877 : node854;
										assign node854 = (inp[12]) ? node870 : node855;
											assign node855 = (inp[9]) ? node863 : node856;
												assign node856 = (inp[6]) ? node860 : node857;
													assign node857 = (inp[5]) ? 14'b01110110100110 : 14'b01111110100110;
													assign node860 = (inp[5]) ? 14'b00110100100110 : 14'b00111100100110;
												assign node863 = (inp[2]) ? node867 : node864;
													assign node864 = (inp[6]) ? 14'b01111100000110 : 14'b01111110000110;
													assign node867 = (inp[5]) ? 14'b00110110000110 : 14'b00111110000110;
											assign node870 = (inp[2]) ? 14'b00000000000001 : node871;
												assign node871 = (inp[5]) ? node873 : 14'b00000000000001;
													assign node873 = (inp[6]) ? 14'b01010100000010 : 14'b01010110000010;
										assign node877 = (inp[12]) ? node879 : 14'b00000000000001;
											assign node879 = (inp[2]) ? 14'b00000000000001 : node880;
												assign node880 = (inp[5]) ? 14'b01010100100000 : node881;
													assign node881 = (inp[9]) ? 14'b01011100000000 : 14'b01011110100000;
								assign node886 = (inp[9]) ? 14'b00000000000001 : node887;
									assign node887 = (inp[4]) ? node917 : node888;
										assign node888 = (inp[12]) ? node902 : node889;
											assign node889 = (inp[11]) ? node897 : node890;
												assign node890 = (inp[5]) ? node894 : node891;
													assign node891 = (inp[2]) ? 14'b00001110000000 : 14'b00000000000001;
													assign node894 = (inp[2]) ? 14'b00000110100000 : 14'b00100110000010;
												assign node897 = (inp[5]) ? 14'b01100110100100 : node898;
													assign node898 = (inp[6]) ? 14'b01101110000100 : 14'b00101110100100;
											assign node902 = (inp[11]) ? node910 : node903;
												assign node903 = (inp[5]) ? node907 : node904;
													assign node904 = (inp[2]) ? 14'b00001110000110 : 14'b01001110100110;
													assign node907 = (inp[2]) ? 14'b00000110000110 : 14'b01000110000110;
												assign node910 = (inp[6]) ? node914 : node911;
													assign node911 = (inp[2]) ? 14'b00000110100100 : 14'b01000110100100;
													assign node914 = (inp[5]) ? 14'b00000110000100 : 14'b01001110000100;
										assign node917 = (inp[2]) ? node931 : node918;
											assign node918 = (inp[5]) ? node924 : node919;
												assign node919 = (inp[11]) ? node921 : 14'b00000000000001;
													assign node921 = (inp[12]) ? 14'b01001110000000 : 14'b00000000000001;
												assign node924 = (inp[11]) ? node928 : node925;
													assign node925 = (inp[12]) ? 14'b01000110000010 : 14'b01100110000110;
													assign node928 = (inp[12]) ? 14'b01000110000000 : 14'b00000000000001;
											assign node931 = (inp[12]) ? 14'b00000000000001 : node932;
												assign node932 = (inp[11]) ? 14'b00000000000001 : node933;
													assign node933 = (inp[6]) ? 14'b00101110000110 : 14'b00101110100110;
							assign node939 = (inp[6]) ? node1015 : node940;
								assign node940 = (inp[9]) ? node990 : node941;
									assign node941 = (inp[4]) ? node971 : node942;
										assign node942 = (inp[11]) ? node956 : node943;
											assign node943 = (inp[12]) ? node949 : node944;
												assign node944 = (inp[2]) ? node946 : 14'b00000000000001;
													assign node946 = (inp[3]) ? 14'b00000010100000 : 14'b00011010100000;
												assign node949 = (inp[3]) ? node953 : node950;
													assign node950 = (inp[2]) ? 14'b00010010100110 : 14'b01010010100110;
													assign node953 = (inp[2]) ? 14'b00000010100110 : 14'b01000010100110;
											assign node956 = (inp[12]) ? node964 : node957;
												assign node957 = (inp[2]) ? node961 : node958;
													assign node958 = (inp[5]) ? 14'b01100010100100 : 14'b01101010100100;
													assign node961 = (inp[5]) ? 14'b00100010100100 : 14'b00101010100100;
												assign node964 = (inp[2]) ? node968 : node965;
													assign node965 = (inp[5]) ? 14'b01010010100100 : 14'b01001010100100;
													assign node968 = (inp[5]) ? 14'b00000010100100 : 14'b00011010100100;
										assign node971 = (inp[11]) ? node985 : node972;
											assign node972 = (inp[12]) ? node980 : node973;
												assign node973 = (inp[2]) ? node977 : node974;
													assign node974 = (inp[3]) ? 14'b01101010100110 : 14'b01110010100110;
													assign node977 = (inp[3]) ? 14'b00100010100110 : 14'b00111010100110;
												assign node980 = (inp[5]) ? node982 : 14'b00000000000001;
													assign node982 = (inp[2]) ? 14'b00000000000001 : 14'b01000010100010;
											assign node985 = (inp[12]) ? node987 : 14'b00000000000001;
												assign node987 = (inp[2]) ? 14'b00000000000001 : 14'b01010010100000;
									assign node990 = (inp[3]) ? node992 : 14'b00000000000001;
										assign node992 = (inp[4]) ? node1008 : node993;
											assign node993 = (inp[12]) ? node1001 : node994;
												assign node994 = (inp[11]) ? node998 : node995;
													assign node995 = (inp[5]) ? 14'b00000010000000 : 14'b00000000000001;
													assign node998 = (inp[2]) ? 14'b00101010000100 : 14'b01100010000100;
												assign node1001 = (inp[5]) ? node1005 : node1002;
													assign node1002 = (inp[2]) ? 14'b00001010000110 : 14'b01001010000110;
													assign node1005 = (inp[11]) ? 14'b00000010000100 : 14'b00000010000110;
											assign node1008 = (inp[11]) ? 14'b00000000000001 : node1009;
												assign node1009 = (inp[12]) ? 14'b00000000000001 : node1010;
													assign node1010 = (inp[5]) ? 14'b00100010000110 : 14'b00101010000110;
								assign node1015 = (inp[9]) ? node1017 : 14'b00000000000001;
									assign node1017 = (inp[3]) ? 14'b00000000000001 : node1018;
										assign node1018 = (inp[2]) ? node1034 : node1019;
											assign node1019 = (inp[5]) ? node1027 : node1020;
												assign node1020 = (inp[11]) ? node1024 : node1021;
													assign node1021 = (inp[4]) ? 14'b00000000000000 : 14'b00000000000001;
													assign node1024 = (inp[12]) ? 14'b01011000000000 : 14'b00000000000001;
												assign node1027 = (inp[11]) ? node1031 : node1028;
													assign node1028 = (inp[4]) ? 14'b01110000000110 : 14'b01010000000110;
													assign node1031 = (inp[4]) ? 14'b00000000000000 : 14'b01110000000100;
											assign node1034 = (inp[5]) ? node1038 : node1035;
												assign node1035 = (inp[4]) ? 14'b00111000000110 : 14'b00011000000000;
												assign node1038 = (inp[4]) ? node1042 : node1039;
													assign node1039 = (inp[11]) ? 14'b00010000000100 : 14'b00010000000000;
													assign node1042 = (inp[12]) ? 14'b00000000000001 : 14'b00000000000000;
						assign node1046 = (inp[11]) ? 14'b00000000000001 : node1047;
							assign node1047 = (inp[2]) ? node1117 : node1048;
								assign node1048 = (inp[12]) ? node1096 : node1049;
									assign node1049 = (inp[1]) ? node1075 : node1050;
										assign node1050 = (inp[3]) ? node1066 : node1051;
											assign node1051 = (inp[9]) ? node1059 : node1052;
												assign node1052 = (inp[5]) ? node1056 : node1053;
													assign node1053 = (inp[4]) ? 14'b01111100100000 : 14'b01111100100010;
													assign node1056 = (inp[4]) ? 14'b01110100100000 : 14'b01110100100010;
												assign node1059 = (inp[4]) ? node1063 : node1060;
													assign node1060 = (inp[5]) ? 14'b01110100000010 : 14'b01111100000010;
													assign node1063 = (inp[6]) ? 14'b01110100000000 : 14'b01110110000000;
											assign node1066 = (inp[9]) ? 14'b00000000000001 : node1067;
												assign node1067 = (inp[6]) ? node1071 : node1068;
													assign node1068 = (inp[4]) ? 14'b01100110100000 : 14'b01100110100010;
													assign node1071 = (inp[4]) ? 14'b01101110000000 : 14'b01101110000010;
										assign node1075 = (inp[6]) ? node1089 : node1076;
											assign node1076 = (inp[9]) ? node1084 : node1077;
												assign node1077 = (inp[5]) ? node1081 : node1078;
													assign node1078 = (inp[3]) ? 14'b01101010100000 : 14'b01111010100000;
													assign node1081 = (inp[3]) ? 14'b01100010100010 : 14'b01110010100000;
												assign node1084 = (inp[3]) ? node1086 : 14'b00000000000001;
													assign node1086 = (inp[5]) ? 14'b01100010000000 : 14'b01101010000000;
											assign node1089 = (inp[3]) ? 14'b00000000000001 : node1090;
												assign node1090 = (inp[9]) ? node1092 : 14'b00000000000001;
													assign node1092 = (inp[5]) ? 14'b01110000000000 : 14'b01111000000010;
									assign node1096 = (inp[5]) ? 14'b00000000000001 : node1097;
										assign node1097 = (inp[6]) ? node1109 : node1098;
											assign node1098 = (inp[9]) ? node1104 : node1099;
												assign node1099 = (inp[4]) ? node1101 : 14'b01011010100010;
													assign node1101 = (inp[1]) ? 14'b00111010100000 : 14'b00101110100000;
												assign node1104 = (inp[4]) ? node1106 : 14'b00000000000001;
													assign node1106 = (inp[1]) ? 14'b00000000000000 : 14'b00000000000000;
											assign node1109 = (inp[3]) ? 14'b00000000000001 : node1110;
												assign node1110 = (inp[1]) ? node1112 : 14'b01011100100010;
													assign node1112 = (inp[9]) ? 14'b00111000000000 : 14'b00000000000001;
								assign node1117 = (inp[4]) ? node1159 : node1118;
									assign node1118 = (inp[12]) ? node1132 : node1119;
										assign node1119 = (inp[5]) ? 14'b00000000000001 : node1120;
											assign node1120 = (inp[6]) ? node1126 : node1121;
												assign node1121 = (inp[3]) ? node1123 : 14'b00000000000001;
													assign node1123 = (inp[9]) ? 14'b00101010000010 : 14'b00101010100010;
												assign node1126 = (inp[3]) ? 14'b00000000000001 : node1127;
													assign node1127 = (inp[9]) ? 14'b00111000000010 : 14'b00000000000001;
										assign node1132 = (inp[9]) ? node1146 : node1133;
											assign node1133 = (inp[1]) ? node1141 : node1134;
												assign node1134 = (inp[3]) ? node1138 : node1135;
													assign node1135 = (inp[5]) ? 14'b00010100100010 : 14'b00011100100010;
													assign node1138 = (inp[6]) ? 14'b00000110000010 : 14'b00001110100010;
												assign node1141 = (inp[6]) ? 14'b00000000000001 : node1142;
													assign node1142 = (inp[5]) ? 14'b00000010100010 : 14'b00001010100010;
											assign node1146 = (inp[3]) ? node1154 : node1147;
												assign node1147 = (inp[1]) ? node1151 : node1148;
													assign node1148 = (inp[6]) ? 14'b00010100000010 : 14'b00011110000010;
													assign node1151 = (inp[6]) ? 14'b00011000000010 : 14'b00000000000001;
												assign node1154 = (inp[1]) ? node1156 : 14'b00000000000001;
													assign node1156 = (inp[6]) ? 14'b00000000000001 : 14'b00000010000010;
									assign node1159 = (inp[5]) ? node1161 : 14'b00000000000001;
										assign node1161 = (inp[12]) ? 14'b00000000000001 : node1162;
											assign node1162 = (inp[3]) ? node1170 : node1163;
												assign node1163 = (inp[6]) ? node1167 : node1164;
													assign node1164 = (inp[1]) ? 14'b00110010100000 : 14'b00110110000000;
													assign node1167 = (inp[9]) ? 14'b00110000000000 : 14'b00000000000001;
												assign node1170 = (inp[9]) ? node1174 : node1171;
													assign node1171 = (inp[1]) ? 14'b00100010100000 : 14'b00100110000000;
													assign node1174 = (inp[1]) ? 14'b00000000000000 : 14'b00000000000001;
		assign node1180 = (inp[0]) ? node2432 : node1181;
			assign node1181 = (inp[5]) ? node2033 : node1182;
				assign node1182 = (inp[6]) ? node1712 : node1183;
					assign node1183 = (inp[2]) ? node1497 : node1184;
						assign node1184 = (inp[3]) ? node1330 : node1185;
							assign node1185 = (inp[1]) ? node1245 : node1186;
								assign node1186 = (inp[9]) ? node1198 : node1187;
									assign node1187 = (inp[4]) ? 14'b00000000000001 : node1188;
										assign node1188 = (inp[12]) ? 14'b00000000000001 : node1189;
											assign node1189 = (inp[8]) ? 14'b10000000001000 : node1190;
												assign node1190 = (inp[10]) ? 14'b00000000000001 : node1191;
													assign node1191 = (inp[7]) ? 14'b00000000000001 : 14'b10000000001000;
									assign node1198 = (inp[4]) ? node1222 : node1199;
										assign node1199 = (inp[12]) ? node1211 : node1200;
											assign node1200 = (inp[10]) ? node1206 : node1201;
												assign node1201 = (inp[7]) ? node1203 : 14'b00000000000001;
													assign node1203 = (inp[8]) ? 14'b00000000000000 : 14'b00000000000010;
												assign node1206 = (inp[8]) ? 14'b00000000000001 : node1207;
													assign node1207 = (inp[7]) ? 14'b01100000000010 : 14'b01100100000010;
											assign node1211 = (inp[8]) ? node1219 : node1212;
												assign node1212 = (inp[10]) ? node1216 : node1213;
													assign node1213 = (inp[7]) ? 14'b00000000000000 : 14'b01000000000100;
													assign node1216 = (inp[7]) ? 14'b01100000000000 : 14'b01100100000000;
												assign node1219 = (inp[7]) ? 14'b01000000000100 : 14'b01000100000100;
										assign node1222 = (inp[7]) ? node1234 : node1223;
											assign node1223 = (inp[8]) ? node1231 : node1224;
												assign node1224 = (inp[12]) ? node1228 : node1225;
													assign node1225 = (inp[10]) ? 14'b00100100000010 : 14'b00100100000110;
													assign node1228 = (inp[10]) ? 14'b00100100000000 : 14'b00100100000100;
												assign node1231 = (inp[12]) ? 14'b00000100000100 : 14'b00100100000100;
											assign node1234 = (inp[8]) ? node1242 : node1235;
												assign node1235 = (inp[10]) ? node1239 : node1236;
													assign node1236 = (inp[12]) ? 14'b00100000000100 : 14'b00100000000110;
													assign node1239 = (inp[12]) ? 14'b00100000000000 : 14'b00100000000010;
												assign node1242 = (inp[12]) ? 14'b00000000000100 : 14'b00100000000100;
								assign node1245 = (inp[4]) ? node1285 : node1246;
									assign node1246 = (inp[12]) ? node1266 : node1247;
										assign node1247 = (inp[7]) ? node1255 : node1248;
											assign node1248 = (inp[8]) ? 14'b00000000000001 : node1249;
												assign node1249 = (inp[10]) ? node1251 : 14'b00000000000001;
													assign node1251 = (inp[9]) ? 14'b01110110000010 : 14'b01110110100010;
											assign node1255 = (inp[8]) ? node1263 : node1256;
												assign node1256 = (inp[10]) ? node1260 : node1257;
													assign node1257 = (inp[9]) ? 14'b00010010000010 : 14'b00010010100010;
													assign node1260 = (inp[9]) ? 14'b01110010000010 : 14'b01110010100010;
												assign node1263 = (inp[9]) ? 14'b00010010000000 : 14'b00010010100000;
										assign node1266 = (inp[9]) ? node1274 : node1267;
											assign node1267 = (inp[8]) ? node1271 : node1268;
												assign node1268 = (inp[7]) ? 14'b00010010100000 : 14'b01010010100100;
												assign node1271 = (inp[7]) ? 14'b01010010100100 : 14'b01010110100100;
											assign node1274 = (inp[8]) ? node1282 : node1275;
												assign node1275 = (inp[10]) ? node1279 : node1276;
													assign node1276 = (inp[7]) ? 14'b00010010000000 : 14'b01010010000100;
													assign node1279 = (inp[7]) ? 14'b01110010000000 : 14'b01110110000000;
												assign node1282 = (inp[7]) ? 14'b01010010000100 : 14'b01010110000100;
									assign node1285 = (inp[9]) ? node1307 : node1286;
										assign node1286 = (inp[7]) ? node1296 : node1287;
											assign node1287 = (inp[8]) ? node1293 : node1288;
												assign node1288 = (inp[12]) ? node1290 : 14'b00110110100110;
													assign node1290 = (inp[11]) ? 14'b00110110100100 : 14'b00110110100000;
												assign node1293 = (inp[12]) ? 14'b00010110100100 : 14'b00110110100100;
											assign node1296 = (inp[8]) ? node1304 : node1297;
												assign node1297 = (inp[10]) ? node1301 : node1298;
													assign node1298 = (inp[12]) ? 14'b00110010100100 : 14'b00110010100110;
													assign node1301 = (inp[12]) ? 14'b00110010100000 : 14'b00110010100010;
												assign node1304 = (inp[12]) ? 14'b00010010100100 : 14'b00110010100100;
										assign node1307 = (inp[7]) ? node1319 : node1308;
											assign node1308 = (inp[8]) ? node1316 : node1309;
												assign node1309 = (inp[10]) ? node1313 : node1310;
													assign node1310 = (inp[12]) ? 14'b00110110000100 : 14'b00110110000110;
													assign node1313 = (inp[12]) ? 14'b00110110000000 : 14'b00110110000010;
												assign node1316 = (inp[12]) ? 14'b00010110000100 : 14'b00110110000100;
											assign node1319 = (inp[8]) ? node1327 : node1320;
												assign node1320 = (inp[12]) ? node1324 : node1321;
													assign node1321 = (inp[10]) ? 14'b00110010000010 : 14'b00110010000110;
													assign node1324 = (inp[10]) ? 14'b00110010000000 : 14'b00110010000100;
												assign node1327 = (inp[12]) ? 14'b00010010000100 : 14'b00110010000100;
							assign node1330 = (inp[1]) ? node1412 : node1331;
								assign node1331 = (inp[4]) ? node1375 : node1332;
									assign node1332 = (inp[12]) ? node1352 : node1333;
										assign node1333 = (inp[7]) ? node1341 : node1334;
											assign node1334 = (inp[10]) ? node1336 : 14'b00000000000001;
												assign node1336 = (inp[8]) ? 14'b00000000000001 : node1337;
													assign node1337 = (inp[9]) ? 14'b01110110010010 : 14'b01110110110010;
											assign node1341 = (inp[8]) ? node1349 : node1342;
												assign node1342 = (inp[10]) ? node1346 : node1343;
													assign node1343 = (inp[9]) ? 14'b00010010010010 : 14'b00010010110010;
													assign node1346 = (inp[9]) ? 14'b01110010010010 : 14'b01110010110010;
												assign node1349 = (inp[9]) ? 14'b00010010010000 : 14'b00010010110000;
										assign node1352 = (inp[9]) ? node1364 : node1353;
											assign node1353 = (inp[8]) ? node1361 : node1354;
												assign node1354 = (inp[10]) ? node1358 : node1355;
													assign node1355 = (inp[7]) ? 14'b00010010110000 : 14'b01010010110100;
													assign node1358 = (inp[11]) ? 14'b01110010110000 : 14'b01110110110000;
												assign node1361 = (inp[7]) ? 14'b01010010110100 : 14'b01010110110100;
											assign node1364 = (inp[8]) ? node1372 : node1365;
												assign node1365 = (inp[10]) ? node1369 : node1366;
													assign node1366 = (inp[11]) ? 14'b01010010010100 : 14'b00010010010000;
													assign node1369 = (inp[7]) ? 14'b01110010010000 : 14'b01110110010000;
												assign node1372 = (inp[7]) ? 14'b01010010010100 : 14'b01010110010100;
									assign node1375 = (inp[7]) ? node1389 : node1376;
										assign node1376 = (inp[8]) ? node1384 : node1377;
											assign node1377 = (inp[10]) ? node1381 : node1378;
												assign node1378 = (inp[9]) ? 14'b00110110010100 : 14'b00110110110100;
												assign node1381 = (inp[12]) ? 14'b00110110110000 : 14'b00110110110010;
											assign node1384 = (inp[12]) ? node1386 : 14'b00110110110100;
												assign node1386 = (inp[9]) ? 14'b00010110010100 : 14'b00010110110100;
										assign node1389 = (inp[9]) ? node1401 : node1390;
											assign node1390 = (inp[8]) ? node1398 : node1391;
												assign node1391 = (inp[12]) ? node1395 : node1392;
													assign node1392 = (inp[10]) ? 14'b00110010110010 : 14'b00110010110110;
													assign node1395 = (inp[10]) ? 14'b00110010110000 : 14'b00110010110100;
												assign node1398 = (inp[12]) ? 14'b00010010110100 : 14'b00110010110100;
											assign node1401 = (inp[8]) ? node1409 : node1402;
												assign node1402 = (inp[10]) ? node1406 : node1403;
													assign node1403 = (inp[12]) ? 14'b00110010010100 : 14'b00110010010110;
													assign node1406 = (inp[12]) ? 14'b00110010010000 : 14'b00110010010010;
												assign node1409 = (inp[12]) ? 14'b00010010010100 : 14'b00110010010100;
								assign node1412 = (inp[9]) ? node1456 : node1413;
									assign node1413 = (inp[4]) ? node1433 : node1414;
										assign node1414 = (inp[12]) ? node1422 : node1415;
											assign node1415 = (inp[8]) ? node1419 : node1416;
												assign node1416 = (inp[7]) ? 14'b00000010100010 : 14'b01100110100010;
												assign node1419 = (inp[7]) ? 14'b00000010100000 : 14'b00000000000001;
											assign node1422 = (inp[8]) ? node1430 : node1423;
												assign node1423 = (inp[10]) ? node1427 : node1424;
													assign node1424 = (inp[7]) ? 14'b00000010100000 : 14'b01000010100100;
													assign node1427 = (inp[7]) ? 14'b01100010100000 : 14'b01100110100000;
												assign node1430 = (inp[7]) ? 14'b01000010100100 : 14'b01000110100100;
										assign node1433 = (inp[7]) ? node1445 : node1434;
											assign node1434 = (inp[8]) ? node1442 : node1435;
												assign node1435 = (inp[10]) ? node1439 : node1436;
													assign node1436 = (inp[12]) ? 14'b00100110100100 : 14'b00100110100110;
													assign node1439 = (inp[12]) ? 14'b00100110100000 : 14'b00100110100010;
												assign node1442 = (inp[12]) ? 14'b00000110100100 : 14'b00100110100100;
											assign node1445 = (inp[8]) ? node1453 : node1446;
												assign node1446 = (inp[12]) ? node1450 : node1447;
													assign node1447 = (inp[10]) ? 14'b00100010100010 : 14'b00100010100110;
													assign node1450 = (inp[10]) ? 14'b00100010100000 : 14'b00100010100100;
												assign node1453 = (inp[12]) ? 14'b00000010100100 : 14'b00100010100100;
									assign node1456 = (inp[8]) ? node1482 : node1457;
										assign node1457 = (inp[10]) ? node1467 : node1458;
											assign node1458 = (inp[4]) ? node1464 : node1459;
												assign node1459 = (inp[12]) ? 14'b01000010000100 : node1460;
													assign node1460 = (inp[7]) ? 14'b00000010000010 : 14'b00000000000001;
												assign node1464 = (inp[7]) ? 14'b00100010000110 : 14'b00100110000110;
											assign node1467 = (inp[4]) ? node1475 : node1468;
												assign node1468 = (inp[7]) ? node1472 : node1469;
													assign node1469 = (inp[12]) ? 14'b01100110000000 : 14'b01100110000010;
													assign node1472 = (inp[12]) ? 14'b01100010000000 : 14'b01100010000010;
												assign node1475 = (inp[7]) ? node1479 : node1476;
													assign node1476 = (inp[12]) ? 14'b00100110000000 : 14'b00100110000010;
													assign node1479 = (inp[12]) ? 14'b00100010000000 : 14'b00100010000010;
										assign node1482 = (inp[12]) ? node1490 : node1483;
											assign node1483 = (inp[4]) ? node1487 : node1484;
												assign node1484 = (inp[7]) ? 14'b00000010000000 : 14'b00000000000001;
												assign node1487 = (inp[7]) ? 14'b00100010000100 : 14'b00100110000100;
											assign node1490 = (inp[7]) ? node1494 : node1491;
												assign node1491 = (inp[4]) ? 14'b00000110000100 : 14'b01000110000100;
												assign node1494 = (inp[4]) ? 14'b00000010000100 : 14'b01000010000100;
						assign node1497 = (inp[4]) ? node1661 : node1498;
							assign node1498 = (inp[10]) ? node1610 : node1499;
								assign node1499 = (inp[7]) ? node1555 : node1500;
									assign node1500 = (inp[12]) ? node1528 : node1501;
										assign node1501 = (inp[8]) ? node1513 : node1502;
											assign node1502 = (inp[9]) ? node1506 : node1503;
												assign node1503 = (inp[3]) ? 14'b01100110100110 : 14'b01110110100110;
												assign node1506 = (inp[3]) ? node1510 : node1507;
													assign node1507 = (inp[1]) ? 14'b01110110000110 : 14'b01100100000110;
													assign node1510 = (inp[1]) ? 14'b01100110000110 : 14'b01110110010110;
											assign node1513 = (inp[9]) ? node1521 : node1514;
												assign node1514 = (inp[1]) ? node1518 : node1515;
													assign node1515 = (inp[11]) ? 14'b00000000000001 : 14'b01110110110100;
													assign node1518 = (inp[3]) ? 14'b01100110100100 : 14'b01110110100100;
												assign node1521 = (inp[1]) ? node1525 : node1522;
													assign node1522 = (inp[3]) ? 14'b01110110010100 : 14'b01100100000100;
													assign node1525 = (inp[3]) ? 14'b01100110000100 : 14'b01110110000100;
										assign node1528 = (inp[8]) ? node1542 : node1529;
											assign node1529 = (inp[1]) ? node1537 : node1530;
												assign node1530 = (inp[3]) ? node1534 : node1531;
													assign node1531 = (inp[9]) ? 14'b01100100000100 : 14'b00000000000001;
													assign node1534 = (inp[9]) ? 14'b01110110010100 : 14'b01110110110100;
												assign node1537 = (inp[3]) ? node1539 : 14'b01110110100100;
													assign node1539 = (inp[9]) ? 14'b01100110000100 : 14'b01100110100100;
											assign node1542 = (inp[1]) ? node1548 : node1543;
												assign node1543 = (inp[3]) ? 14'b01010110110000 : node1544;
													assign node1544 = (inp[9]) ? 14'b01000100000000 : 14'b00000000000001;
												assign node1548 = (inp[3]) ? node1552 : node1549;
													assign node1549 = (inp[9]) ? 14'b01010110000000 : 14'b01010110100000;
													assign node1552 = (inp[9]) ? 14'b01000110000000 : 14'b01000110100000;
									assign node1555 = (inp[3]) ? node1581 : node1556;
										assign node1556 = (inp[1]) ? node1566 : node1557;
											assign node1557 = (inp[9]) ? node1559 : 14'b00000000000001;
												assign node1559 = (inp[12]) ? node1563 : node1560;
													assign node1560 = (inp[8]) ? 14'b01100000000100 : 14'b01100000000110;
													assign node1563 = (inp[8]) ? 14'b01000000000000 : 14'b01100000000100;
											assign node1566 = (inp[12]) ? node1574 : node1567;
												assign node1567 = (inp[9]) ? node1571 : node1568;
													assign node1568 = (inp[11]) ? 14'b01110010100100 : 14'b01110010100110;
													assign node1571 = (inp[8]) ? 14'b01110010000100 : 14'b01110010000110;
												assign node1574 = (inp[8]) ? node1578 : node1575;
													assign node1575 = (inp[9]) ? 14'b01110010000100 : 14'b01110010100100;
													assign node1578 = (inp[9]) ? 14'b01010010000000 : 14'b01010010100000;
										assign node1581 = (inp[1]) ? node1597 : node1582;
											assign node1582 = (inp[9]) ? node1590 : node1583;
												assign node1583 = (inp[12]) ? node1587 : node1584;
													assign node1584 = (inp[8]) ? 14'b01110010110100 : 14'b01110010110110;
													assign node1587 = (inp[8]) ? 14'b01010010110000 : 14'b01110010110100;
												assign node1590 = (inp[12]) ? node1594 : node1591;
													assign node1591 = (inp[8]) ? 14'b01110010010100 : 14'b01110010010110;
													assign node1594 = (inp[8]) ? 14'b01010010010000 : 14'b01110010010100;
											assign node1597 = (inp[9]) ? node1603 : node1598;
												assign node1598 = (inp[12]) ? node1600 : 14'b01100010100100;
													assign node1600 = (inp[8]) ? 14'b01000010100000 : 14'b01100010100100;
												assign node1603 = (inp[12]) ? node1607 : node1604;
													assign node1604 = (inp[8]) ? 14'b01100010000100 : 14'b01100010000110;
													assign node1607 = (inp[8]) ? 14'b01000010000000 : 14'b01100010000100;
								assign node1610 = (inp[8]) ? node1612 : 14'b00000000000001;
									assign node1612 = (inp[12]) ? node1634 : node1613;
										assign node1613 = (inp[1]) ? node1619 : node1614;
											assign node1614 = (inp[9]) ? node1616 : 14'b00000000000001;
												assign node1616 = (inp[3]) ? 14'b01110110010100 : 14'b01100100000100;
											assign node1619 = (inp[7]) ? node1627 : node1620;
												assign node1620 = (inp[9]) ? node1624 : node1621;
													assign node1621 = (inp[3]) ? 14'b01100110100100 : 14'b01110110100100;
													assign node1624 = (inp[3]) ? 14'b01100110000100 : 14'b01110110000100;
												assign node1627 = (inp[3]) ? node1631 : node1628;
													assign node1628 = (inp[9]) ? 14'b01110010000100 : 14'b01110010100100;
													assign node1631 = (inp[9]) ? 14'b01100010000100 : 14'b01100010100100;
										assign node1634 = (inp[7]) ? node1650 : node1635;
											assign node1635 = (inp[9]) ? node1643 : node1636;
												assign node1636 = (inp[1]) ? node1640 : node1637;
													assign node1637 = (inp[3]) ? 14'b01010110110000 : 14'b00000000000001;
													assign node1640 = (inp[3]) ? 14'b01000110100000 : 14'b01010110100000;
												assign node1643 = (inp[1]) ? node1647 : node1644;
													assign node1644 = (inp[3]) ? 14'b01010110010000 : 14'b01000100000000;
													assign node1647 = (inp[3]) ? 14'b01000110000000 : 14'b01010110000000;
											assign node1650 = (inp[3]) ? node1656 : node1651;
												assign node1651 = (inp[9]) ? node1653 : 14'b00000000000001;
													assign node1653 = (inp[1]) ? 14'b01010010000000 : 14'b01000000000000;
												assign node1656 = (inp[1]) ? 14'b01000010100000 : node1657;
													assign node1657 = (inp[9]) ? 14'b01010010010000 : 14'b01010010110000;
							assign node1661 = (inp[8]) ? 14'b00000000000001 : node1662;
								assign node1662 = (inp[7]) ? 14'b00000000000001 : node1663;
									assign node1663 = (inp[12]) ? node1681 : node1664;
										assign node1664 = (inp[10]) ? node1666 : 14'b00000000000001;
											assign node1666 = (inp[9]) ? node1674 : node1667;
												assign node1667 = (inp[1]) ? node1671 : node1668;
													assign node1668 = (inp[3]) ? 14'b00010110110010 : 14'b00000000000001;
													assign node1671 = (inp[3]) ? 14'b00000110100010 : 14'b00010110100010;
												assign node1674 = (inp[3]) ? node1678 : node1675;
													assign node1675 = (inp[1]) ? 14'b00010110000010 : 14'b00000100000010;
													assign node1678 = (inp[1]) ? 14'b00000110000010 : 14'b00010110010010;
										assign node1681 = (inp[10]) ? node1697 : node1682;
											assign node1682 = (inp[3]) ? node1690 : node1683;
												assign node1683 = (inp[1]) ? node1687 : node1684;
													assign node1684 = (inp[9]) ? 14'b00000100000100 : 14'b00000000000001;
													assign node1687 = (inp[9]) ? 14'b00010110000100 : 14'b00010110100100;
												assign node1690 = (inp[1]) ? node1694 : node1691;
													assign node1691 = (inp[9]) ? 14'b00010110010100 : 14'b00010110110100;
													assign node1694 = (inp[9]) ? 14'b00000110000100 : 14'b00000110100100;
											assign node1697 = (inp[9]) ? node1703 : node1698;
												assign node1698 = (inp[1]) ? node1700 : 14'b00010110110000;
													assign node1700 = (inp[3]) ? 14'b00000110100000 : 14'b00010110100000;
												assign node1703 = (inp[1]) ? node1707 : node1704;
													assign node1704 = (inp[3]) ? 14'b00010110010000 : 14'b00000100000000;
													assign node1707 = (inp[3]) ? 14'b00000110000000 : 14'b00010110000000;
					assign node1712 = (inp[3]) ? node2002 : node1713;
						assign node1713 = (inp[2]) ? node1883 : node1714;
							assign node1714 = (inp[4]) ? node1792 : node1715;
								assign node1715 = (inp[12]) ? node1747 : node1716;
									assign node1716 = (inp[7]) ? node1724 : node1717;
										assign node1717 = (inp[8]) ? 14'b00000000000001 : node1718;
											assign node1718 = (inp[10]) ? node1720 : 14'b00000000000001;
												assign node1720 = (inp[9]) ? 14'b01110100000010 : 14'b01110100110010;
										assign node1724 = (inp[8]) ? node1740 : node1725;
											assign node1725 = (inp[10]) ? node1733 : node1726;
												assign node1726 = (inp[1]) ? node1730 : node1727;
													assign node1727 = (inp[9]) ? 14'b00010000010010 : 14'b00010000110010;
													assign node1730 = (inp[9]) ? 14'b00010000000010 : 14'b00010000100010;
												assign node1733 = (inp[9]) ? node1737 : node1734;
													assign node1734 = (inp[1]) ? 14'b01110000100010 : 14'b01110000110010;
													assign node1737 = (inp[1]) ? 14'b01110000000010 : 14'b01110000010010;
											assign node1740 = (inp[9]) ? node1744 : node1741;
												assign node1741 = (inp[1]) ? 14'b00010000100000 : 14'b00010000110000;
												assign node1744 = (inp[1]) ? 14'b00010000000000 : 14'b00010000010000;
									assign node1747 = (inp[8]) ? node1779 : node1748;
										assign node1748 = (inp[10]) ? node1764 : node1749;
											assign node1749 = (inp[7]) ? node1757 : node1750;
												assign node1750 = (inp[9]) ? node1754 : node1751;
													assign node1751 = (inp[1]) ? 14'b01010000100100 : 14'b01010000110100;
													assign node1754 = (inp[11]) ? 14'b01010000000100 : 14'b01010000010100;
												assign node1757 = (inp[9]) ? node1761 : node1758;
													assign node1758 = (inp[1]) ? 14'b00010000100000 : 14'b00010000110000;
													assign node1761 = (inp[1]) ? 14'b00010000000000 : 14'b00010000010000;
											assign node1764 = (inp[9]) ? node1772 : node1765;
												assign node1765 = (inp[1]) ? node1769 : node1766;
													assign node1766 = (inp[7]) ? 14'b01110000110000 : 14'b01110100110000;
													assign node1769 = (inp[7]) ? 14'b01110000100000 : 14'b01110100100000;
												assign node1772 = (inp[1]) ? node1776 : node1773;
													assign node1773 = (inp[7]) ? 14'b01110000010000 : 14'b01110100010000;
													assign node1776 = (inp[7]) ? 14'b01110000000000 : 14'b01110100000000;
										assign node1779 = (inp[7]) ? node1785 : node1780;
											assign node1780 = (inp[1]) ? node1782 : 14'b01010100010100;
												assign node1782 = (inp[9]) ? 14'b01010100000100 : 14'b01010100100100;
											assign node1785 = (inp[1]) ? node1789 : node1786;
												assign node1786 = (inp[9]) ? 14'b01010000010100 : 14'b01010000110100;
												assign node1789 = (inp[9]) ? 14'b01010000000100 : 14'b01010000100100;
								assign node1792 = (inp[9]) ? node1836 : node1793;
									assign node1793 = (inp[7]) ? node1815 : node1794;
										assign node1794 = (inp[8]) ? node1808 : node1795;
											assign node1795 = (inp[12]) ? node1803 : node1796;
												assign node1796 = (inp[1]) ? node1800 : node1797;
													assign node1797 = (inp[10]) ? 14'b00110100110010 : 14'b00110100110110;
													assign node1800 = (inp[10]) ? 14'b00110100100010 : 14'b00110100100110;
												assign node1803 = (inp[10]) ? 14'b00110100110000 : node1804;
													assign node1804 = (inp[1]) ? 14'b00110100100100 : 14'b00110100110100;
											assign node1808 = (inp[1]) ? node1812 : node1809;
												assign node1809 = (inp[12]) ? 14'b00010100110100 : 14'b00110100110100;
												assign node1812 = (inp[12]) ? 14'b00010100100100 : 14'b00110100100100;
										assign node1815 = (inp[1]) ? node1827 : node1816;
											assign node1816 = (inp[8]) ? node1824 : node1817;
												assign node1817 = (inp[12]) ? node1821 : node1818;
													assign node1818 = (inp[10]) ? 14'b00110000110010 : 14'b00110000110110;
													assign node1821 = (inp[10]) ? 14'b00110000110000 : 14'b00110000110100;
												assign node1824 = (inp[12]) ? 14'b00010000110100 : 14'b00110000110100;
											assign node1827 = (inp[8]) ? node1833 : node1828;
												assign node1828 = (inp[12]) ? node1830 : 14'b00110000100110;
													assign node1830 = (inp[10]) ? 14'b00110000100000 : 14'b00110000100100;
												assign node1833 = (inp[12]) ? 14'b00010000100100 : 14'b00110000100100;
									assign node1836 = (inp[1]) ? node1860 : node1837;
										assign node1837 = (inp[7]) ? node1849 : node1838;
											assign node1838 = (inp[8]) ? node1846 : node1839;
												assign node1839 = (inp[10]) ? node1843 : node1840;
													assign node1840 = (inp[12]) ? 14'b00110100010100 : 14'b00110100010110;
													assign node1843 = (inp[12]) ? 14'b00110100010000 : 14'b00110100010010;
												assign node1846 = (inp[12]) ? 14'b00010100010100 : 14'b00110100010100;
											assign node1849 = (inp[8]) ? node1857 : node1850;
												assign node1850 = (inp[10]) ? node1854 : node1851;
													assign node1851 = (inp[12]) ? 14'b00110000010100 : 14'b00110000010110;
													assign node1854 = (inp[12]) ? 14'b00110000010000 : 14'b00110000010010;
												assign node1857 = (inp[10]) ? 14'b00110000010100 : 14'b00010000010100;
										assign node1860 = (inp[7]) ? node1872 : node1861;
											assign node1861 = (inp[8]) ? node1869 : node1862;
												assign node1862 = (inp[12]) ? node1866 : node1863;
													assign node1863 = (inp[10]) ? 14'b00110100000010 : 14'b00110100000110;
													assign node1866 = (inp[10]) ? 14'b00110100000000 : 14'b00110100000100;
												assign node1869 = (inp[12]) ? 14'b00010100000100 : 14'b00110100000100;
											assign node1872 = (inp[8]) ? node1880 : node1873;
												assign node1873 = (inp[12]) ? node1877 : node1874;
													assign node1874 = (inp[10]) ? 14'b00110000000010 : 14'b00110000000110;
													assign node1877 = (inp[10]) ? 14'b00110000000000 : 14'b00110000000100;
												assign node1880 = (inp[12]) ? 14'b00010000000100 : 14'b00110000000100;
							assign node1883 = (inp[4]) ? node1977 : node1884;
								assign node1884 = (inp[10]) ? node1944 : node1885;
									assign node1885 = (inp[9]) ? node1913 : node1886;
										assign node1886 = (inp[7]) ? node1898 : node1887;
											assign node1887 = (inp[1]) ? node1893 : node1888;
												assign node1888 = (inp[8]) ? node1890 : 14'b01110100110100;
													assign node1890 = (inp[12]) ? 14'b01010100110000 : 14'b01110100110100;
												assign node1893 = (inp[11]) ? 14'b01110100100100 : node1894;
													assign node1894 = (inp[12]) ? 14'b01010100100000 : 14'b01110100100110;
											assign node1898 = (inp[1]) ? node1906 : node1899;
												assign node1899 = (inp[12]) ? node1903 : node1900;
													assign node1900 = (inp[8]) ? 14'b01110000110100 : 14'b01110000110110;
													assign node1903 = (inp[8]) ? 14'b01010000110000 : 14'b01110000110100;
												assign node1906 = (inp[12]) ? node1910 : node1907;
													assign node1907 = (inp[8]) ? 14'b01110000100100 : 14'b01110000100110;
													assign node1910 = (inp[8]) ? 14'b01010000100000 : 14'b01110000100100;
										assign node1913 = (inp[1]) ? node1929 : node1914;
											assign node1914 = (inp[12]) ? node1922 : node1915;
												assign node1915 = (inp[7]) ? node1919 : node1916;
													assign node1916 = (inp[8]) ? 14'b01110100010100 : 14'b01110100010110;
													assign node1919 = (inp[8]) ? 14'b01110000010100 : 14'b01110000010110;
												assign node1922 = (inp[8]) ? node1926 : node1923;
													assign node1923 = (inp[11]) ? 14'b01110000010100 : 14'b01110100010100;
													assign node1926 = (inp[7]) ? 14'b01010000010000 : 14'b01010100010000;
											assign node1929 = (inp[7]) ? node1937 : node1930;
												assign node1930 = (inp[8]) ? node1934 : node1931;
													assign node1931 = (inp[12]) ? 14'b01110100000100 : 14'b01110100000110;
													assign node1934 = (inp[12]) ? 14'b01010100000000 : 14'b01110100000100;
												assign node1937 = (inp[12]) ? node1941 : node1938;
													assign node1938 = (inp[8]) ? 14'b01110000000100 : 14'b01110000000110;
													assign node1941 = (inp[8]) ? 14'b01010000000000 : 14'b01110000000100;
									assign node1944 = (inp[8]) ? node1946 : 14'b00000000000001;
										assign node1946 = (inp[12]) ? node1962 : node1947;
											assign node1947 = (inp[9]) ? node1955 : node1948;
												assign node1948 = (inp[1]) ? node1952 : node1949;
													assign node1949 = (inp[7]) ? 14'b01110000110100 : 14'b01110100110100;
													assign node1952 = (inp[7]) ? 14'b01110000100100 : 14'b01110100100100;
												assign node1955 = (inp[7]) ? node1959 : node1956;
													assign node1956 = (inp[1]) ? 14'b01110100000100 : 14'b01110100010100;
													assign node1959 = (inp[1]) ? 14'b01110000000100 : 14'b01110000010100;
											assign node1962 = (inp[1]) ? node1970 : node1963;
												assign node1963 = (inp[7]) ? node1967 : node1964;
													assign node1964 = (inp[9]) ? 14'b01010100010000 : 14'b01010100110000;
													assign node1967 = (inp[9]) ? 14'b01010000010000 : 14'b01010000110000;
												assign node1970 = (inp[9]) ? node1974 : node1971;
													assign node1971 = (inp[11]) ? 14'b01010000100000 : 14'b01010100100000;
													assign node1974 = (inp[7]) ? 14'b01010000000000 : 14'b01010100000000;
								assign node1977 = (inp[8]) ? 14'b00000000000001 : node1978;
									assign node1978 = (inp[7]) ? 14'b00000000000001 : node1979;
										assign node1979 = (inp[12]) ? node1985 : node1980;
											assign node1980 = (inp[10]) ? node1982 : 14'b00000000000001;
												assign node1982 = (inp[9]) ? 14'b00010100000010 : 14'b00010100110010;
											assign node1985 = (inp[1]) ? node1993 : node1986;
												assign node1986 = (inp[9]) ? node1990 : node1987;
													assign node1987 = (inp[10]) ? 14'b00010100110000 : 14'b00010100110100;
													assign node1990 = (inp[10]) ? 14'b00010100010000 : 14'b00010100010100;
												assign node1993 = (inp[10]) ? node1997 : node1994;
													assign node1994 = (inp[9]) ? 14'b00010100000100 : 14'b00010100100100;
													assign node1997 = (inp[9]) ? 14'b00010100000000 : 14'b00010100100000;
						assign node2002 = (inp[2]) ? node2004 : 14'b00000000000001;
							assign node2004 = (inp[12]) ? 14'b00000000000001 : node2005;
								assign node2005 = (inp[9]) ? 14'b00000000000001 : node2006;
									assign node2006 = (inp[4]) ? node2016 : node2007;
										assign node2007 = (inp[7]) ? 14'b00000000000001 : node2008;
											assign node2008 = (inp[11]) ? node2010 : 14'b00000000000001;
												assign node2010 = (inp[1]) ? 14'b00000000000001 : node2011;
													assign node2011 = (inp[8]) ? 14'b00000000000001 : 14'b10000001001000;
										assign node2016 = (inp[1]) ? node2024 : node2017;
											assign node2017 = (inp[7]) ? 14'b00000000000001 : node2018;
												assign node2018 = (inp[10]) ? node2020 : 14'b10000001001010;
													assign node2020 = (inp[8]) ? 14'b10000001001010 : 14'b00000000000001;
											assign node2024 = (inp[7]) ? node2026 : 14'b00000000000001;
												assign node2026 = (inp[8]) ? 14'b10000000000000 : node2027;
													assign node2027 = (inp[10]) ? 14'b10000000000000 : 14'b00000000000001;
				assign node2033 = (inp[12]) ? node2289 : node2034;
					assign node2034 = (inp[2]) ? node2204 : node2035;
						assign node2035 = (inp[8]) ? node2113 : node2036;
							assign node2036 = (inp[10]) ? 14'b00000000000001 : node2037;
								assign node2037 = (inp[6]) ? node2081 : node2038;
									assign node2038 = (inp[7]) ? node2062 : node2039;
										assign node2039 = (inp[3]) ? node2051 : node2040;
											assign node2040 = (inp[1]) ? node2046 : node2041;
												assign node2041 = (inp[9]) ? node2043 : 14'b00000000000001;
													assign node2043 = (inp[4]) ? 14'b00000100000110 : 14'b01000100000110;
												assign node2046 = (inp[9]) ? node2048 : 14'b01010110100110;
													assign node2048 = (inp[4]) ? 14'b00010110000110 : 14'b01010110000110;
											assign node2051 = (inp[1]) ? node2057 : node2052;
												assign node2052 = (inp[9]) ? 14'b00010110010110 : node2053;
													assign node2053 = (inp[4]) ? 14'b00010110110110 : 14'b01010110110110;
												assign node2057 = (inp[4]) ? 14'b00000110000110 : node2058;
													assign node2058 = (inp[9]) ? 14'b01000110000110 : 14'b01000110100110;
										assign node2062 = (inp[1]) ? node2070 : node2063;
											assign node2063 = (inp[4]) ? node2067 : node2064;
												assign node2064 = (inp[9]) ? 14'b01010010010110 : 14'b01010010110110;
												assign node2067 = (inp[9]) ? 14'b00010010010110 : 14'b00010010110110;
											assign node2070 = (inp[9]) ? node2076 : node2071;
												assign node2071 = (inp[3]) ? 14'b01000010100110 : node2072;
													assign node2072 = (inp[11]) ? 14'b01010010100110 : 14'b00010010100110;
												assign node2076 = (inp[3]) ? node2078 : 14'b01010010000110;
													assign node2078 = (inp[4]) ? 14'b00000010000110 : 14'b01000010000110;
									assign node2081 = (inp[3]) ? 14'b00000000000001 : node2082;
										assign node2082 = (inp[9]) ? node2098 : node2083;
											assign node2083 = (inp[4]) ? node2091 : node2084;
												assign node2084 = (inp[7]) ? node2088 : node2085;
													assign node2085 = (inp[1]) ? 14'b01010100100110 : 14'b01010100110110;
													assign node2088 = (inp[1]) ? 14'b01010000100110 : 14'b01010000110110;
												assign node2091 = (inp[7]) ? node2095 : node2092;
													assign node2092 = (inp[1]) ? 14'b00010100100110 : 14'b00010100110110;
													assign node2095 = (inp[11]) ? 14'b00010000100110 : 14'b00010000110110;
											assign node2098 = (inp[4]) ? node2106 : node2099;
												assign node2099 = (inp[7]) ? node2103 : node2100;
													assign node2100 = (inp[1]) ? 14'b01010100000110 : 14'b01010100010110;
													assign node2103 = (inp[1]) ? 14'b01010000000110 : 14'b01010000010110;
												assign node2106 = (inp[1]) ? node2108 : 14'b00010100010110;
													assign node2108 = (inp[7]) ? 14'b00010000000110 : 14'b00010100000110;
							assign node2113 = (inp[6]) ? node2171 : node2114;
								assign node2114 = (inp[1]) ? node2140 : node2115;
									assign node2115 = (inp[3]) ? node2125 : node2116;
										assign node2116 = (inp[9]) ? node2118 : 14'b00000000000001;
											assign node2118 = (inp[4]) ? node2122 : node2119;
												assign node2119 = (inp[7]) ? 14'b01100000000000 : 14'b01100100000000;
												assign node2122 = (inp[7]) ? 14'b00100000000000 : 14'b00100100000000;
										assign node2125 = (inp[9]) ? node2133 : node2126;
											assign node2126 = (inp[7]) ? node2130 : node2127;
												assign node2127 = (inp[4]) ? 14'b00110110110000 : 14'b01110110110000;
												assign node2130 = (inp[4]) ? 14'b00110010110000 : 14'b01110010110000;
											assign node2133 = (inp[4]) ? node2137 : node2134;
												assign node2134 = (inp[7]) ? 14'b01110010010000 : 14'b01110110010000;
												assign node2137 = (inp[7]) ? 14'b00110010010000 : 14'b00110110010000;
									assign node2140 = (inp[3]) ? node2156 : node2141;
										assign node2141 = (inp[4]) ? node2149 : node2142;
											assign node2142 = (inp[7]) ? node2146 : node2143;
												assign node2143 = (inp[9]) ? 14'b01110110000000 : 14'b01110110100000;
												assign node2146 = (inp[9]) ? 14'b01110010000000 : 14'b01110010100000;
											assign node2149 = (inp[7]) ? node2153 : node2150;
												assign node2150 = (inp[9]) ? 14'b00110110000000 : 14'b00110110100000;
												assign node2153 = (inp[9]) ? 14'b00110010000000 : 14'b00110010100000;
										assign node2156 = (inp[9]) ? node2164 : node2157;
											assign node2157 = (inp[4]) ? node2161 : node2158;
												assign node2158 = (inp[7]) ? 14'b01100010100000 : 14'b01100110100000;
												assign node2161 = (inp[7]) ? 14'b00100010100000 : 14'b00100110100000;
											assign node2164 = (inp[7]) ? node2168 : node2165;
												assign node2165 = (inp[4]) ? 14'b00100110000000 : 14'b01100110000000;
												assign node2168 = (inp[4]) ? 14'b00100010000000 : 14'b01100010000000;
								assign node2171 = (inp[3]) ? 14'b00000000000001 : node2172;
									assign node2172 = (inp[7]) ? node2188 : node2173;
										assign node2173 = (inp[1]) ? node2181 : node2174;
											assign node2174 = (inp[9]) ? node2178 : node2175;
												assign node2175 = (inp[4]) ? 14'b00110100110000 : 14'b01110100110000;
												assign node2178 = (inp[4]) ? 14'b00110100010000 : 14'b01110100010000;
											assign node2181 = (inp[9]) ? node2185 : node2182;
												assign node2182 = (inp[4]) ? 14'b00110100100000 : 14'b01110100100000;
												assign node2185 = (inp[4]) ? 14'b00110100000000 : 14'b01110100000000;
										assign node2188 = (inp[1]) ? node2196 : node2189;
											assign node2189 = (inp[9]) ? node2193 : node2190;
												assign node2190 = (inp[4]) ? 14'b00110000110000 : 14'b01110000110000;
												assign node2193 = (inp[4]) ? 14'b00110000010000 : 14'b01110000010000;
											assign node2196 = (inp[4]) ? node2200 : node2197;
												assign node2197 = (inp[9]) ? 14'b01110000000000 : 14'b01110000100000;
												assign node2200 = (inp[9]) ? 14'b00110000000000 : 14'b00110000100000;
						assign node2204 = (inp[7]) ? 14'b00000000000001 : node2205;
							assign node2205 = (inp[4]) ? node2237 : node2206;
								assign node2206 = (inp[8]) ? node2228 : node2207;
									assign node2207 = (inp[10]) ? 14'b00000000000001 : node2208;
										assign node2208 = (inp[3]) ? node2220 : node2209;
											assign node2209 = (inp[9]) ? node2213 : node2210;
												assign node2210 = (inp[1]) ? 14'b01010110100010 : 14'b00000000000001;
												assign node2213 = (inp[6]) ? node2217 : node2214;
													assign node2214 = (inp[1]) ? 14'b01010110000010 : 14'b01000100000010;
													assign node2217 = (inp[1]) ? 14'b01010100000010 : 14'b01010100010010;
											assign node2220 = (inp[6]) ? 14'b00000000000001 : node2221;
												assign node2221 = (inp[1]) ? node2223 : 14'b01010110010010;
													assign node2223 = (inp[9]) ? 14'b01000110000010 : 14'b01000110100010;
									assign node2228 = (inp[3]) ? node2230 : 14'b00000000000001;
										assign node2230 = (inp[6]) ? node2232 : 14'b00000000000001;
											assign node2232 = (inp[9]) ? 14'b00000000000001 : node2233;
												assign node2233 = (inp[1]) ? 14'b00000000000001 : 14'b10000001001000;
								assign node2237 = (inp[8]) ? node2263 : node2238;
									assign node2238 = (inp[10]) ? 14'b00000000000001 : node2239;
										assign node2239 = (inp[6]) ? node2253 : node2240;
											assign node2240 = (inp[3]) ? node2248 : node2241;
												assign node2241 = (inp[1]) ? node2245 : node2242;
													assign node2242 = (inp[9]) ? 14'b01000000000010 : 14'b00000000000001;
													assign node2245 = (inp[9]) ? 14'b01010010000010 : 14'b01010010100010;
												assign node2248 = (inp[1]) ? 14'b01000010000010 : node2249;
													assign node2249 = (inp[9]) ? 14'b01010010010010 : 14'b01010010110010;
											assign node2253 = (inp[3]) ? 14'b00000000000001 : node2254;
												assign node2254 = (inp[9]) ? node2258 : node2255;
													assign node2255 = (inp[1]) ? 14'b01010000100010 : 14'b01010000110010;
													assign node2258 = (inp[11]) ? 14'b01010000000010 : 14'b01010000010010;
									assign node2263 = (inp[6]) ? node2279 : node2264;
										assign node2264 = (inp[9]) ? node2272 : node2265;
											assign node2265 = (inp[1]) ? node2269 : node2266;
												assign node2266 = (inp[3]) ? 14'b00010110110000 : 14'b00000000000001;
												assign node2269 = (inp[3]) ? 14'b00000110100000 : 14'b00010110100000;
											assign node2272 = (inp[3]) ? node2276 : node2273;
												assign node2273 = (inp[1]) ? 14'b00010110000000 : 14'b00000100000000;
												assign node2276 = (inp[1]) ? 14'b00000110000000 : 14'b00010110010000;
										assign node2279 = (inp[3]) ? 14'b00000000000001 : node2280;
											assign node2280 = (inp[1]) ? node2284 : node2281;
												assign node2281 = (inp[9]) ? 14'b00010100010000 : 14'b00010100110000;
												assign node2284 = (inp[9]) ? 14'b00010100000000 : 14'b00010100100000;
					assign node2289 = (inp[10]) ? node2407 : node2290;
						assign node2290 = (inp[8]) ? node2386 : node2291;
							assign node2291 = (inp[4]) ? node2359 : node2292;
								assign node2292 = (inp[7]) ? node2336 : node2293;
									assign node2293 = (inp[3]) ? node2321 : node2294;
										assign node2294 = (inp[6]) ? node2306 : node2295;
											assign node2295 = (inp[1]) ? node2301 : node2296;
												assign node2296 = (inp[9]) ? node2298 : 14'b00000000000001;
													assign node2298 = (inp[2]) ? 14'b01000100000000 : 14'b01000100000100;
												assign node2301 = (inp[2]) ? 14'b01010110000000 : node2302;
													assign node2302 = (inp[9]) ? 14'b01010110000100 : 14'b01010110100100;
											assign node2306 = (inp[1]) ? node2314 : node2307;
												assign node2307 = (inp[9]) ? node2311 : node2308;
													assign node2308 = (inp[11]) ? 14'b01010100110000 : 14'b01010100110100;
													assign node2311 = (inp[2]) ? 14'b01010100010000 : 14'b01010100010100;
												assign node2314 = (inp[9]) ? node2318 : node2315;
													assign node2315 = (inp[2]) ? 14'b01010100100000 : 14'b01010100100100;
													assign node2318 = (inp[2]) ? 14'b01010100000000 : 14'b01010100000100;
										assign node2321 = (inp[6]) ? 14'b00000000000001 : node2322;
											assign node2322 = (inp[1]) ? node2328 : node2323;
												assign node2323 = (inp[9]) ? 14'b01010110010000 : node2324;
													assign node2324 = (inp[2]) ? 14'b01010110110000 : 14'b01010110110100;
												assign node2328 = (inp[9]) ? node2332 : node2329;
													assign node2329 = (inp[2]) ? 14'b01000110100000 : 14'b01000110100100;
													assign node2332 = (inp[2]) ? 14'b01000110000000 : 14'b01000110000100;
									assign node2336 = (inp[2]) ? node2338 : 14'b00000000000001;
										assign node2338 = (inp[6]) ? node2350 : node2339;
											assign node2339 = (inp[3]) ? node2347 : node2340;
												assign node2340 = (inp[1]) ? node2344 : node2341;
													assign node2341 = (inp[9]) ? 14'b01000000000000 : 14'b00000000000001;
													assign node2344 = (inp[9]) ? 14'b01010010000000 : 14'b01010010100000;
												assign node2347 = (inp[9]) ? 14'b01000010000000 : 14'b01010010110000;
											assign node2350 = (inp[3]) ? 14'b00000000000001 : node2351;
												assign node2351 = (inp[9]) ? node2355 : node2352;
													assign node2352 = (inp[1]) ? 14'b01010000100000 : 14'b01010000110000;
													assign node2355 = (inp[1]) ? 14'b01010000000000 : 14'b01010000010000;
								assign node2359 = (inp[2]) ? 14'b00000000000001 : node2360;
									assign node2360 = (inp[7]) ? node2362 : 14'b00000000000001;
										assign node2362 = (inp[6]) ? node2378 : node2363;
											assign node2363 = (inp[9]) ? node2371 : node2364;
												assign node2364 = (inp[1]) ? node2368 : node2365;
													assign node2365 = (inp[3]) ? 14'b00010010110100 : 14'b00000000000001;
													assign node2368 = (inp[3]) ? 14'b00000010100100 : 14'b00010010100100;
												assign node2371 = (inp[1]) ? node2375 : node2372;
													assign node2372 = (inp[3]) ? 14'b00010010010100 : 14'b00000000000100;
													assign node2375 = (inp[3]) ? 14'b00000010000100 : 14'b00010010000100;
											assign node2378 = (inp[3]) ? 14'b00000000000001 : node2379;
												assign node2379 = (inp[9]) ? node2381 : 14'b00010000100100;
													assign node2381 = (inp[1]) ? 14'b00010000000100 : 14'b00010000010100;
							assign node2386 = (inp[1]) ? 14'b00000000000001 : node2387;
								assign node2387 = (inp[9]) ? 14'b00000000000001 : node2388;
									assign node2388 = (inp[6]) ? node2398 : node2389;
										assign node2389 = (inp[3]) ? 14'b00000000000001 : node2390;
											assign node2390 = (inp[2]) ? node2392 : 14'b00000000000001;
												assign node2392 = (inp[7]) ? node2394 : 14'b00000000000001;
													assign node2394 = (inp[4]) ? 14'b10001001000010 : 14'b10001000001000;
										assign node2398 = (inp[3]) ? node2400 : 14'b00000000000001;
											assign node2400 = (inp[2]) ? 14'b00000000000001 : node2401;
												assign node2401 = (inp[7]) ? 14'b00000000000001 : 14'b10001000000010;
						assign node2407 = (inp[1]) ? 14'b00000000000001 : node2408;
							assign node2408 = (inp[9]) ? 14'b00000000000001 : node2409;
								assign node2409 = (inp[8]) ? node2411 : 14'b00000000000001;
									assign node2411 = (inp[3]) ? node2421 : node2412;
										assign node2412 = (inp[2]) ? node2414 : 14'b00000000000001;
											assign node2414 = (inp[7]) ? node2416 : 14'b00000000000001;
												assign node2416 = (inp[6]) ? 14'b00000000000001 : node2417;
													assign node2417 = (inp[4]) ? 14'b10001001000010 : 14'b10001000001000;
										assign node2421 = (inp[4]) ? 14'b00000000000001 : node2422;
											assign node2422 = (inp[7]) ? 14'b00000000000001 : node2423;
												assign node2423 = (inp[6]) ? node2425 : 14'b00000000000001;
													assign node2425 = (inp[2]) ? 14'b00000000000001 : 14'b10001000000010;
			assign node2432 = (inp[1]) ? node3002 : node2433;
				assign node2433 = (inp[3]) ? node2855 : node2434;
					assign node2434 = (inp[5]) ? node2720 : node2435;
						assign node2435 = (inp[2]) ? node2599 : node2436;
							assign node2436 = (inp[4]) ? node2512 : node2437;
								assign node2437 = (inp[12]) ? node2471 : node2438;
									assign node2438 = (inp[8]) ? node2462 : node2439;
										assign node2439 = (inp[10]) ? node2447 : node2440;
											assign node2440 = (inp[7]) ? node2442 : 14'b00000000000001;
												assign node2442 = (inp[6]) ? node2444 : 14'b00000010010010;
													assign node2444 = (inp[11]) ? 14'b00000000110010 : 14'b00000000010010;
											assign node2447 = (inp[7]) ? node2455 : node2448;
												assign node2448 = (inp[6]) ? node2452 : node2449;
													assign node2449 = (inp[9]) ? 14'b01100110010010 : 14'b01100110110010;
													assign node2452 = (inp[9]) ? 14'b01100100010010 : 14'b01100100110010;
												assign node2455 = (inp[9]) ? node2459 : node2456;
													assign node2456 = (inp[6]) ? 14'b01100000110010 : 14'b01100010110010;
													assign node2459 = (inp[6]) ? 14'b01100000010010 : 14'b01100010010010;
										assign node2462 = (inp[7]) ? node2464 : 14'b00000000000001;
											assign node2464 = (inp[6]) ? node2468 : node2465;
												assign node2465 = (inp[9]) ? 14'b00000010010000 : 14'b00000010110000;
												assign node2468 = (inp[9]) ? 14'b00000000010000 : 14'b00000000110000;
									assign node2471 = (inp[6]) ? node2493 : node2472;
										assign node2472 = (inp[9]) ? node2482 : node2473;
											assign node2473 = (inp[8]) ? node2479 : node2474;
												assign node2474 = (inp[10]) ? node2476 : 14'b01000010110100;
													assign node2476 = (inp[7]) ? 14'b01100010110000 : 14'b01100110110000;
												assign node2479 = (inp[7]) ? 14'b01000010110100 : 14'b01000110110100;
											assign node2482 = (inp[8]) ? node2490 : node2483;
												assign node2483 = (inp[10]) ? node2487 : node2484;
													assign node2484 = (inp[11]) ? 14'b01000010010100 : 14'b00000010010000;
													assign node2487 = (inp[7]) ? 14'b01100010010000 : 14'b01100110010000;
												assign node2490 = (inp[7]) ? 14'b01000010010100 : 14'b01000110010100;
										assign node2493 = (inp[9]) ? node2505 : node2494;
											assign node2494 = (inp[8]) ? node2502 : node2495;
												assign node2495 = (inp[10]) ? node2499 : node2496;
													assign node2496 = (inp[7]) ? 14'b00000000110000 : 14'b01000000110100;
													assign node2499 = (inp[7]) ? 14'b01100000110000 : 14'b01100100110000;
												assign node2502 = (inp[7]) ? 14'b01000000110100 : 14'b01000100110100;
											assign node2505 = (inp[8]) ? node2509 : node2506;
												assign node2506 = (inp[7]) ? 14'b01100000010000 : 14'b01000000010100;
												assign node2509 = (inp[7]) ? 14'b01000000010100 : 14'b01000100010100;
								assign node2512 = (inp[7]) ? node2558 : node2513;
									assign node2513 = (inp[9]) ? node2535 : node2514;
										assign node2514 = (inp[8]) ? node2528 : node2515;
											assign node2515 = (inp[6]) ? node2523 : node2516;
												assign node2516 = (inp[10]) ? node2520 : node2517;
													assign node2517 = (inp[12]) ? 14'b00100110110100 : 14'b00100110110110;
													assign node2520 = (inp[12]) ? 14'b00100110110000 : 14'b00100110110010;
												assign node2523 = (inp[12]) ? node2525 : 14'b00100100110010;
													assign node2525 = (inp[10]) ? 14'b00100100110000 : 14'b00100100110100;
											assign node2528 = (inp[6]) ? node2532 : node2529;
												assign node2529 = (inp[12]) ? 14'b00000110110100 : 14'b00100110110100;
												assign node2532 = (inp[12]) ? 14'b00000100110100 : 14'b00100100110100;
										assign node2535 = (inp[6]) ? node2547 : node2536;
											assign node2536 = (inp[8]) ? node2544 : node2537;
												assign node2537 = (inp[12]) ? node2541 : node2538;
													assign node2538 = (inp[10]) ? 14'b00100110010010 : 14'b00100110010110;
													assign node2541 = (inp[10]) ? 14'b00100110010000 : 14'b00100110010100;
												assign node2544 = (inp[12]) ? 14'b00000110010100 : 14'b00100110010100;
											assign node2547 = (inp[8]) ? node2555 : node2548;
												assign node2548 = (inp[10]) ? node2552 : node2549;
													assign node2549 = (inp[12]) ? 14'b00100100010100 : 14'b00100100010110;
													assign node2552 = (inp[12]) ? 14'b00100100010000 : 14'b00100100010010;
												assign node2555 = (inp[12]) ? 14'b00000100010100 : 14'b00100100010100;
									assign node2558 = (inp[6]) ? node2578 : node2559;
										assign node2559 = (inp[9]) ? node2569 : node2560;
											assign node2560 = (inp[8]) ? node2566 : node2561;
												assign node2561 = (inp[10]) ? node2563 : 14'b00100010110100;
													assign node2563 = (inp[12]) ? 14'b00100010110000 : 14'b00100010110010;
												assign node2566 = (inp[12]) ? 14'b00000010110100 : 14'b00100010110100;
											assign node2569 = (inp[8]) ? node2575 : node2570;
												assign node2570 = (inp[10]) ? node2572 : 14'b00100010010100;
													assign node2572 = (inp[12]) ? 14'b00100010010000 : 14'b00100010010010;
												assign node2575 = (inp[12]) ? 14'b00000010010100 : 14'b00100010010100;
										assign node2578 = (inp[9]) ? node2588 : node2579;
											assign node2579 = (inp[12]) ? node2585 : node2580;
												assign node2580 = (inp[8]) ? 14'b00100000110100 : node2581;
													assign node2581 = (inp[10]) ? 14'b00100000110010 : 14'b00100000110110;
												assign node2585 = (inp[8]) ? 14'b00000000110100 : 14'b00100000110100;
											assign node2588 = (inp[8]) ? node2596 : node2589;
												assign node2589 = (inp[12]) ? node2593 : node2590;
													assign node2590 = (inp[11]) ? 14'b00100000010110 : 14'b00100000010010;
													assign node2593 = (inp[10]) ? 14'b00100000010000 : 14'b00100000010100;
												assign node2596 = (inp[12]) ? 14'b00000000010100 : 14'b00100000010100;
							assign node2599 = (inp[4]) ? node2691 : node2600;
								assign node2600 = (inp[10]) ? node2662 : node2601;
									assign node2601 = (inp[7]) ? node2633 : node2602;
										assign node2602 = (inp[9]) ? node2618 : node2603;
											assign node2603 = (inp[8]) ? node2611 : node2604;
												assign node2604 = (inp[12]) ? node2608 : node2605;
													assign node2605 = (inp[6]) ? 14'b01100100110110 : 14'b01100110110110;
													assign node2608 = (inp[6]) ? 14'b01100100110100 : 14'b01100110110100;
												assign node2611 = (inp[12]) ? node2615 : node2612;
													assign node2612 = (inp[6]) ? 14'b01100100110100 : 14'b01100110110100;
													assign node2615 = (inp[6]) ? 14'b01000100110000 : 14'b01000110110000;
											assign node2618 = (inp[6]) ? node2626 : node2619;
												assign node2619 = (inp[8]) ? node2623 : node2620;
													assign node2620 = (inp[12]) ? 14'b01100110010100 : 14'b01100110010110;
													assign node2623 = (inp[12]) ? 14'b01000110010000 : 14'b01100110010100;
												assign node2626 = (inp[8]) ? node2630 : node2627;
													assign node2627 = (inp[12]) ? 14'b01100100010100 : 14'b01100100010110;
													assign node2630 = (inp[12]) ? 14'b01000100010000 : 14'b01100100010100;
										assign node2633 = (inp[6]) ? node2649 : node2634;
											assign node2634 = (inp[9]) ? node2642 : node2635;
												assign node2635 = (inp[8]) ? node2639 : node2636;
													assign node2636 = (inp[12]) ? 14'b01100010110100 : 14'b01100010110110;
													assign node2639 = (inp[12]) ? 14'b01000010110000 : 14'b01100010110100;
												assign node2642 = (inp[8]) ? node2646 : node2643;
													assign node2643 = (inp[12]) ? 14'b01100010010100 : 14'b01100010010110;
													assign node2646 = (inp[12]) ? 14'b01000010010000 : 14'b01100010010100;
											assign node2649 = (inp[9]) ? node2657 : node2650;
												assign node2650 = (inp[8]) ? node2654 : node2651;
													assign node2651 = (inp[12]) ? 14'b01100000110100 : 14'b01100000110110;
													assign node2654 = (inp[12]) ? 14'b01000000110000 : 14'b01100000110100;
												assign node2657 = (inp[8]) ? node2659 : 14'b01100000010100;
													assign node2659 = (inp[12]) ? 14'b01000000010000 : 14'b01100000010100;
									assign node2662 = (inp[8]) ? node2664 : 14'b00000000000001;
										assign node2664 = (inp[12]) ? node2678 : node2665;
											assign node2665 = (inp[6]) ? node2671 : node2666;
												assign node2666 = (inp[9]) ? 14'b01100110010100 : node2667;
													assign node2667 = (inp[7]) ? 14'b01100010110100 : 14'b01100110110100;
												assign node2671 = (inp[9]) ? node2675 : node2672;
													assign node2672 = (inp[7]) ? 14'b01100000110100 : 14'b01100100110100;
													assign node2675 = (inp[7]) ? 14'b01100000010100 : 14'b01100100010100;
											assign node2678 = (inp[6]) ? node2686 : node2679;
												assign node2679 = (inp[7]) ? node2683 : node2680;
													assign node2680 = (inp[11]) ? 14'b01000110010000 : 14'b01000110110000;
													assign node2683 = (inp[9]) ? 14'b01000010010000 : 14'b01000010110000;
												assign node2686 = (inp[7]) ? 14'b01000000110000 : node2687;
													assign node2687 = (inp[9]) ? 14'b01000100010000 : 14'b01000100110000;
								assign node2691 = (inp[7]) ? 14'b00000000000001 : node2692;
									assign node2692 = (inp[8]) ? 14'b00000000000001 : node2693;
										assign node2693 = (inp[12]) ? node2703 : node2694;
											assign node2694 = (inp[10]) ? node2696 : 14'b00000000000001;
												assign node2696 = (inp[6]) ? node2700 : node2697;
													assign node2697 = (inp[9]) ? 14'b00000110010010 : 14'b00000110110010;
													assign node2700 = (inp[11]) ? 14'b00000100010010 : 14'b00000100110010;
											assign node2703 = (inp[9]) ? node2711 : node2704;
												assign node2704 = (inp[10]) ? node2708 : node2705;
													assign node2705 = (inp[6]) ? 14'b00000100110100 : 14'b00000110110100;
													assign node2708 = (inp[6]) ? 14'b00000100110000 : 14'b00000110110000;
												assign node2711 = (inp[10]) ? node2715 : node2712;
													assign node2712 = (inp[6]) ? 14'b00000100010100 : 14'b00000110010100;
													assign node2715 = (inp[6]) ? 14'b00000100010000 : 14'b00000110010000;
						assign node2720 = (inp[12]) ? node2816 : node2721;
							assign node2721 = (inp[2]) ? node2783 : node2722;
								assign node2722 = (inp[8]) ? node2752 : node2723;
									assign node2723 = (inp[10]) ? 14'b00000000000001 : node2724;
										assign node2724 = (inp[4]) ? node2738 : node2725;
											assign node2725 = (inp[7]) ? node2733 : node2726;
												assign node2726 = (inp[6]) ? node2730 : node2727;
													assign node2727 = (inp[9]) ? 14'b01000110010110 : 14'b01000110110110;
													assign node2730 = (inp[9]) ? 14'b01000100010110 : 14'b01000100110110;
												assign node2733 = (inp[6]) ? 14'b01000000110110 : node2734;
													assign node2734 = (inp[9]) ? 14'b01000010010110 : 14'b01000010110110;
											assign node2738 = (inp[9]) ? node2744 : node2739;
												assign node2739 = (inp[7]) ? 14'b00000010110110 : node2740;
													assign node2740 = (inp[6]) ? 14'b00000100110110 : 14'b00000110110110;
												assign node2744 = (inp[6]) ? node2748 : node2745;
													assign node2745 = (inp[7]) ? 14'b00000010010110 : 14'b00000110010110;
													assign node2748 = (inp[7]) ? 14'b00000000010110 : 14'b00000100010110;
									assign node2752 = (inp[4]) ? node2768 : node2753;
										assign node2753 = (inp[9]) ? node2761 : node2754;
											assign node2754 = (inp[7]) ? node2758 : node2755;
												assign node2755 = (inp[6]) ? 14'b01100100110000 : 14'b01100110110000;
												assign node2758 = (inp[6]) ? 14'b01100000110000 : 14'b01100010110000;
											assign node2761 = (inp[7]) ? node2765 : node2762;
												assign node2762 = (inp[6]) ? 14'b01100100010000 : 14'b01100110010000;
												assign node2765 = (inp[6]) ? 14'b01100000010000 : 14'b01100010010000;
										assign node2768 = (inp[7]) ? node2776 : node2769;
											assign node2769 = (inp[6]) ? node2773 : node2770;
												assign node2770 = (inp[9]) ? 14'b00100110010000 : 14'b00100110110000;
												assign node2773 = (inp[9]) ? 14'b00100100010000 : 14'b00100100110000;
											assign node2776 = (inp[9]) ? node2780 : node2777;
												assign node2777 = (inp[6]) ? 14'b00100000110000 : 14'b00100010110000;
												assign node2780 = (inp[6]) ? 14'b00100000010000 : 14'b00100010010000;
								assign node2783 = (inp[7]) ? 14'b00000000000001 : node2784;
									assign node2784 = (inp[10]) ? node2806 : node2785;
										assign node2785 = (inp[8]) ? node2799 : node2786;
											assign node2786 = (inp[4]) ? node2794 : node2787;
												assign node2787 = (inp[9]) ? node2791 : node2788;
													assign node2788 = (inp[6]) ? 14'b01000100110010 : 14'b01000110110010;
													assign node2791 = (inp[6]) ? 14'b01000100010010 : 14'b01000110010010;
												assign node2794 = (inp[9]) ? node2796 : 14'b01000010110010;
													assign node2796 = (inp[6]) ? 14'b01000000010010 : 14'b01000010010010;
											assign node2799 = (inp[4]) ? node2801 : 14'b00000000000001;
												assign node2801 = (inp[6]) ? node2803 : 14'b00000110110000;
													assign node2803 = (inp[9]) ? 14'b00000100010000 : 14'b00000100110000;
										assign node2806 = (inp[4]) ? node2808 : 14'b00000000000001;
											assign node2808 = (inp[8]) ? node2810 : 14'b00000000000001;
												assign node2810 = (inp[6]) ? node2812 : 14'b00000110010000;
													assign node2812 = (inp[9]) ? 14'b00000100010000 : 14'b00000100110000;
							assign node2816 = (inp[10]) ? 14'b00000000000001 : node2817;
								assign node2817 = (inp[8]) ? 14'b00000000000001 : node2818;
									assign node2818 = (inp[4]) ? node2842 : node2819;
										assign node2819 = (inp[7]) ? node2835 : node2820;
											assign node2820 = (inp[9]) ? node2828 : node2821;
												assign node2821 = (inp[2]) ? node2825 : node2822;
													assign node2822 = (inp[6]) ? 14'b01000100110100 : 14'b01000110110100;
													assign node2825 = (inp[6]) ? 14'b01000100110000 : 14'b01000110110000;
												assign node2828 = (inp[6]) ? node2832 : node2829;
													assign node2829 = (inp[2]) ? 14'b01000110010000 : 14'b01000110010100;
													assign node2832 = (inp[2]) ? 14'b01000100010000 : 14'b01000100010100;
											assign node2835 = (inp[2]) ? node2837 : 14'b00000000000001;
												assign node2837 = (inp[6]) ? 14'b01000000010000 : node2838;
													assign node2838 = (inp[9]) ? 14'b01000010010000 : 14'b01000010110000;
										assign node2842 = (inp[7]) ? node2844 : 14'b00000000000001;
											assign node2844 = (inp[2]) ? 14'b00000000000001 : node2845;
												assign node2845 = (inp[6]) ? node2849 : node2846;
													assign node2846 = (inp[9]) ? 14'b00000010010100 : 14'b00000010110100;
													assign node2849 = (inp[9]) ? 14'b00000000010100 : 14'b00000000110100;
					assign node2855 = (inp[6]) ? node2877 : node2856;
						assign node2856 = (inp[7]) ? 14'b00000000000001 : node2857;
							assign node2857 = (inp[12]) ? 14'b00000000000001 : node2858;
								assign node2858 = (inp[4]) ? 14'b00000000000001 : node2859;
									assign node2859 = (inp[2]) ? node2861 : 14'b00000000000001;
										assign node2861 = (inp[9]) ? 14'b00000000000001 : node2862;
											assign node2862 = (inp[10]) ? node2868 : node2863;
												assign node2863 = (inp[5]) ? node2865 : 14'b00000000000001;
													assign node2865 = (inp[8]) ? 14'b10000001000000 : 14'b00000000000001;
												assign node2868 = (inp[8]) ? 14'b00000000000001 : node2869;
													assign node2869 = (inp[5]) ? 14'b00000000000001 : 14'b10000001000000;
						assign node2877 = (inp[9]) ? 14'b00000000000001 : node2878;
							assign node2878 = (inp[2]) ? node2954 : node2879;
								assign node2879 = (inp[5]) ? node2927 : node2880;
									assign node2880 = (inp[4]) ? node2904 : node2881;
										assign node2881 = (inp[12]) ? node2893 : node2882;
											assign node2882 = (inp[8]) ? node2890 : node2883;
												assign node2883 = (inp[10]) ? node2887 : node2884;
													assign node2884 = (inp[7]) ? 14'b00000000100010 : 14'b00000000000001;
													assign node2887 = (inp[7]) ? 14'b01100000100010 : 14'b01100100100010;
												assign node2890 = (inp[7]) ? 14'b00000000100000 : 14'b00000000000001;
											assign node2893 = (inp[10]) ? node2899 : node2894;
												assign node2894 = (inp[7]) ? 14'b01000000100100 : node2895;
													assign node2895 = (inp[8]) ? 14'b01000100100100 : 14'b01000000100100;
												assign node2899 = (inp[8]) ? node2901 : 14'b01100100100000;
													assign node2901 = (inp[11]) ? 14'b01000100100100 : 14'b01000000100100;
										assign node2904 = (inp[7]) ? node2916 : node2905;
											assign node2905 = (inp[8]) ? node2913 : node2906;
												assign node2906 = (inp[10]) ? node2910 : node2907;
													assign node2907 = (inp[12]) ? 14'b00100100100100 : 14'b00100100100110;
													assign node2910 = (inp[12]) ? 14'b00100100100000 : 14'b00100100100010;
												assign node2913 = (inp[12]) ? 14'b00000100100100 : 14'b00100100100100;
											assign node2916 = (inp[10]) ? node2922 : node2917;
												assign node2917 = (inp[12]) ? 14'b00100000100100 : node2918;
													assign node2918 = (inp[8]) ? 14'b00100000100100 : 14'b00100000100110;
												assign node2922 = (inp[8]) ? node2924 : 14'b00100000100000;
													assign node2924 = (inp[12]) ? 14'b00000000100100 : 14'b00100000100100;
									assign node2927 = (inp[12]) ? node2945 : node2928;
										assign node2928 = (inp[8]) ? node2938 : node2929;
											assign node2929 = (inp[10]) ? 14'b00000000000001 : node2930;
												assign node2930 = (inp[4]) ? node2934 : node2931;
													assign node2931 = (inp[7]) ? 14'b01000000100110 : 14'b01000100100110;
													assign node2934 = (inp[7]) ? 14'b00000000100110 : 14'b00000100100110;
											assign node2938 = (inp[4]) ? node2942 : node2939;
												assign node2939 = (inp[7]) ? 14'b01100000100000 : 14'b01100100100000;
												assign node2942 = (inp[7]) ? 14'b00100000100000 : 14'b00100100100000;
										assign node2945 = (inp[10]) ? 14'b00000000000001 : node2946;
											assign node2946 = (inp[8]) ? 14'b00000000000001 : node2947;
												assign node2947 = (inp[11]) ? 14'b00000000000001 : node2948;
													assign node2948 = (inp[7]) ? 14'b00000000000000 : 14'b01000100100100;
								assign node2954 = (inp[4]) ? node2988 : node2955;
									assign node2955 = (inp[10]) ? node2979 : node2956;
										assign node2956 = (inp[5]) ? node2970 : node2957;
											assign node2957 = (inp[12]) ? node2965 : node2958;
												assign node2958 = (inp[7]) ? node2962 : node2959;
													assign node2959 = (inp[8]) ? 14'b01100100100100 : 14'b01100100100110;
													assign node2962 = (inp[8]) ? 14'b01100000100100 : 14'b01100000100110;
												assign node2965 = (inp[8]) ? node2967 : 14'b01100000100100;
													assign node2967 = (inp[7]) ? 14'b01000000100000 : 14'b01000100100000;
											assign node2970 = (inp[8]) ? 14'b00000000000001 : node2971;
												assign node2971 = (inp[7]) ? node2975 : node2972;
													assign node2972 = (inp[12]) ? 14'b01000100100000 : 14'b01000100100010;
													assign node2975 = (inp[12]) ? 14'b01000000100000 : 14'b00000000000001;
										assign node2979 = (inp[8]) ? node2981 : 14'b00000000000001;
											assign node2981 = (inp[5]) ? 14'b00000000000001 : node2982;
												assign node2982 = (inp[12]) ? node2984 : 14'b01100000100100;
													assign node2984 = (inp[7]) ? 14'b01000000100000 : 14'b01000100100000;
									assign node2988 = (inp[7]) ? 14'b00000000000001 : node2989;
										assign node2989 = (inp[8]) ? 14'b00000000000001 : node2990;
											assign node2990 = (inp[5]) ? node2996 : node2991;
												assign node2991 = (inp[12]) ? node2993 : 14'b00000100100010;
													assign node2993 = (inp[10]) ? 14'b00000100100000 : 14'b00000100100100;
												assign node2996 = (inp[10]) ? 14'b00000000000001 : 14'b01000000100010;
				assign node3002 = (inp[8]) ? node3032 : node3003;
					assign node3003 = (inp[12]) ? 14'b00000000000001 : node3004;
						assign node3004 = (inp[6]) ? 14'b00000000000001 : node3005;
							assign node3005 = (inp[7]) ? 14'b00000000000001 : node3006;
								assign node3006 = (inp[5]) ? 14'b00000000000001 : node3007;
									assign node3007 = (inp[9]) ? node3019 : node3008;
										assign node3008 = (inp[2]) ? node3010 : 14'b00000000000001;
											assign node3010 = (inp[3]) ? 14'b00000000000001 : node3011;
												assign node3011 = (inp[10]) ? node3015 : node3012;
													assign node3012 = (inp[4]) ? 14'b10000001000010 : 14'b00000000000001;
													assign node3015 = (inp[4]) ? 14'b00000000000001 : 14'b10000000001010;
										assign node3019 = (inp[4]) ? 14'b00000000000001 : node3020;
											assign node3020 = (inp[10]) ? 14'b00000000000001 : node3021;
												assign node3021 = (inp[3]) ? node3023 : 14'b00000000000001;
													assign node3023 = (inp[2]) ? 14'b00000000000001 : 14'b10000000000010;
					assign node3032 = (inp[5]) ? node3054 : node3033;
						assign node3033 = (inp[7]) ? 14'b00000000000001 : node3034;
							assign node3034 = (inp[6]) ? 14'b00000000000001 : node3035;
								assign node3035 = (inp[12]) ? 14'b00000000000001 : node3036;
									assign node3036 = (inp[3]) ? node3044 : node3037;
										assign node3037 = (inp[2]) ? node3039 : 14'b00000000000001;
											assign node3039 = (inp[9]) ? 14'b00000000000001 : node3040;
												assign node3040 = (inp[4]) ? 14'b10000001000010 : 14'b00000000000001;
										assign node3044 = (inp[9]) ? node3046 : 14'b00000000000001;
											assign node3046 = (inp[4]) ? 14'b00000000000001 : node3047;
												assign node3047 = (inp[2]) ? 14'b00000000000001 : 14'b10000000000010;
						assign node3054 = (inp[12]) ? node3068 : node3055;
							assign node3055 = (inp[9]) ? 14'b00000000000001 : node3056;
								assign node3056 = (inp[4]) ? 14'b00000000000001 : node3057;
									assign node3057 = (inp[7]) ? 14'b00000000000001 : node3058;
										assign node3058 = (inp[3]) ? 14'b00000000000001 : node3059;
											assign node3059 = (inp[2]) ? node3061 : 14'b00000000000001;
												assign node3061 = (inp[6]) ? 14'b00000000000001 : 14'b10000000001010;
							assign node3068 = (inp[2]) ? node3080 : node3069;
								assign node3069 = (inp[9]) ? 14'b00000000000001 : node3070;
									assign node3070 = (inp[3]) ? 14'b00000000000001 : node3071;
										assign node3071 = (inp[7]) ? 14'b00000000000001 : node3072;
											assign node3072 = (inp[6]) ? 14'b00000000000001 : node3073;
												assign node3073 = (inp[4]) ? 14'b00000000000001 : 14'b10001001001000;
								assign node3080 = (inp[3]) ? node3082 : 14'b00000000000001;
									assign node3082 = (inp[9]) ? node3084 : 14'b00000000000001;
										assign node3084 = (inp[7]) ? node3086 : 14'b00000000000001;
											assign node3086 = (inp[4]) ? node3090 : node3087;
												assign node3087 = (inp[6]) ? 14'b10001001000000 : 14'b10001000000000;
												assign node3090 = (inp[6]) ? 14'b10001001001010 : 14'b10001000001010;

endmodule