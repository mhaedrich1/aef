module dtc_split5_bm58 (
	input  wire [12-1:0] inp,
	output wire [3-1:0] outp
);

	wire [3-1:0] node2;
	wire [3-1:0] node3;
	wire [3-1:0] node4;
	wire [3-1:0] node5;
	wire [3-1:0] node6;
	wire [3-1:0] node7;
	wire [3-1:0] node8;
	wire [3-1:0] node9;
	wire [3-1:0] node10;
	wire [3-1:0] node16;
	wire [3-1:0] node18;
	wire [3-1:0] node19;
	wire [3-1:0] node21;
	wire [3-1:0] node24;
	wire [3-1:0] node28;
	wire [3-1:0] node29;
	wire [3-1:0] node30;
	wire [3-1:0] node31;
	wire [3-1:0] node32;
	wire [3-1:0] node33;
	wire [3-1:0] node38;
	wire [3-1:0] node39;
	wire [3-1:0] node41;
	wire [3-1:0] node46;
	wire [3-1:0] node47;
	wire [3-1:0] node48;
	wire [3-1:0] node49;
	wire [3-1:0] node51;
	wire [3-1:0] node54;
	wire [3-1:0] node56;
	wire [3-1:0] node59;
	wire [3-1:0] node60;
	wire [3-1:0] node63;
	wire [3-1:0] node64;
	wire [3-1:0] node67;
	wire [3-1:0] node70;
	wire [3-1:0] node71;
	wire [3-1:0] node72;
	wire [3-1:0] node75;
	wire [3-1:0] node76;
	wire [3-1:0] node80;
	wire [3-1:0] node81;
	wire [3-1:0] node84;
	wire [3-1:0] node86;
	wire [3-1:0] node89;
	wire [3-1:0] node90;
	wire [3-1:0] node92;
	wire [3-1:0] node93;
	wire [3-1:0] node94;
	wire [3-1:0] node95;
	wire [3-1:0] node96;
	wire [3-1:0] node97;
	wire [3-1:0] node102;
	wire [3-1:0] node104;
	wire [3-1:0] node108;
	wire [3-1:0] node110;
	wire [3-1:0] node111;
	wire [3-1:0] node112;
	wire [3-1:0] node116;
	wire [3-1:0] node118;
	wire [3-1:0] node121;
	wire [3-1:0] node122;
	wire [3-1:0] node123;
	wire [3-1:0] node124;
	wire [3-1:0] node125;
	wire [3-1:0] node126;
	wire [3-1:0] node127;
	wire [3-1:0] node131;
	wire [3-1:0] node135;
	wire [3-1:0] node136;
	wire [3-1:0] node138;
	wire [3-1:0] node139;
	wire [3-1:0] node144;
	wire [3-1:0] node145;
	wire [3-1:0] node146;
	wire [3-1:0] node147;
	wire [3-1:0] node151;
	wire [3-1:0] node152;
	wire [3-1:0] node156;
	wire [3-1:0] node157;
	wire [3-1:0] node160;
	wire [3-1:0] node163;
	wire [3-1:0] node164;
	wire [3-1:0] node165;
	wire [3-1:0] node166;
	wire [3-1:0] node167;
	wire [3-1:0] node169;
	wire [3-1:0] node172;
	wire [3-1:0] node175;
	wire [3-1:0] node178;
	wire [3-1:0] node179;
	wire [3-1:0] node180;
	wire [3-1:0] node183;
	wire [3-1:0] node186;
	wire [3-1:0] node189;
	wire [3-1:0] node190;
	wire [3-1:0] node191;
	wire [3-1:0] node194;
	wire [3-1:0] node198;
	wire [3-1:0] node200;
	wire [3-1:0] node201;
	wire [3-1:0] node202;
	wire [3-1:0] node203;
	wire [3-1:0] node204;
	wire [3-1:0] node205;
	wire [3-1:0] node206;
	wire [3-1:0] node212;
	wire [3-1:0] node213;
	wire [3-1:0] node214;
	wire [3-1:0] node216;
	wire [3-1:0] node220;
	wire [3-1:0] node221;
	wire [3-1:0] node222;
	wire [3-1:0] node227;
	wire [3-1:0] node228;
	wire [3-1:0] node230;
	wire [3-1:0] node231;
	wire [3-1:0] node232;
	wire [3-1:0] node237;
	wire [3-1:0] node238;
	wire [3-1:0] node239;
	wire [3-1:0] node240;
	wire [3-1:0] node241;
	wire [3-1:0] node246;
	wire [3-1:0] node248;
	wire [3-1:0] node251;
	wire [3-1:0] node252;
	wire [3-1:0] node253;
	wire [3-1:0] node256;
	wire [3-1:0] node260;
	wire [3-1:0] node262;
	wire [3-1:0] node263;
	wire [3-1:0] node264;
	wire [3-1:0] node265;
	wire [3-1:0] node268;
	wire [3-1:0] node269;
	wire [3-1:0] node273;
	wire [3-1:0] node275;
	wire [3-1:0] node276;
	wire [3-1:0] node280;
	wire [3-1:0] node282;
	wire [3-1:0] node284;
	wire [3-1:0] node286;
	wire [3-1:0] node287;

	assign outp = (inp[6]) ? node2 : 3'b000;
		assign node2 = (inp[0]) ? node198 : node3;
			assign node3 = (inp[4]) ? node89 : node4;
				assign node4 = (inp[9]) ? node28 : node5;
					assign node5 = (inp[1]) ? 3'b000 : node6;
						assign node6 = (inp[11]) ? node16 : node7;
							assign node7 = (inp[10]) ? 3'b100 : node8;
								assign node8 = (inp[8]) ? 3'b100 : node9;
									assign node9 = (inp[3]) ? 3'b000 : node10;
										assign node10 = (inp[7]) ? 3'b000 : 3'b100;
							assign node16 = (inp[8]) ? node18 : 3'b000;
								assign node18 = (inp[3]) ? node24 : node19;
									assign node19 = (inp[5]) ? node21 : 3'b100;
										assign node21 = (inp[7]) ? 3'b000 : 3'b100;
									assign node24 = (inp[10]) ? 3'b100 : 3'b000;
					assign node28 = (inp[8]) ? node46 : node29;
						assign node29 = (inp[1]) ? 3'b100 : node30;
							assign node30 = (inp[10]) ? node38 : node31;
								assign node31 = (inp[11]) ? 3'b100 : node32;
									assign node32 = (inp[2]) ? 3'b000 : node33;
										assign node33 = (inp[3]) ? 3'b100 : 3'b000;
								assign node38 = (inp[2]) ? 3'b000 : node39;
									assign node39 = (inp[3]) ? node41 : 3'b000;
										assign node41 = (inp[11]) ? 3'b100 : 3'b000;
						assign node46 = (inp[3]) ? node70 : node47;
							assign node47 = (inp[2]) ? node59 : node48;
								assign node48 = (inp[1]) ? node54 : node49;
									assign node49 = (inp[10]) ? node51 : 3'b000;
										assign node51 = (inp[11]) ? 3'b000 : 3'b100;
									assign node54 = (inp[11]) ? node56 : 3'b000;
										assign node56 = (inp[10]) ? 3'b000 : 3'b100;
								assign node59 = (inp[11]) ? node63 : node60;
									assign node60 = (inp[1]) ? 3'b000 : 3'b100;
									assign node63 = (inp[10]) ? node67 : node64;
										assign node64 = (inp[1]) ? 3'b100 : 3'b000;
										assign node67 = (inp[1]) ? 3'b000 : 3'b100;
							assign node70 = (inp[11]) ? node80 : node71;
								assign node71 = (inp[1]) ? node75 : node72;
									assign node72 = (inp[10]) ? 3'b100 : 3'b000;
									assign node75 = (inp[2]) ? 3'b000 : node76;
										assign node76 = (inp[10]) ? 3'b000 : 3'b100;
								assign node80 = (inp[1]) ? node84 : node81;
									assign node81 = (inp[2]) ? 3'b100 : 3'b000;
									assign node84 = (inp[10]) ? node86 : 3'b100;
										assign node86 = (inp[2]) ? 3'b000 : 3'b100;
				assign node89 = (inp[9]) ? node121 : node90;
					assign node90 = (inp[1]) ? node92 : 3'b100;
						assign node92 = (inp[11]) ? node108 : node93;
							assign node93 = (inp[8]) ? 3'b100 : node94;
								assign node94 = (inp[3]) ? node102 : node95;
									assign node95 = (inp[2]) ? 3'b100 : node96;
										assign node96 = (inp[10]) ? 3'b100 : node97;
											assign node97 = (inp[7]) ? 3'b000 : 3'b100;
									assign node102 = (inp[10]) ? node104 : 3'b000;
										assign node104 = (inp[7]) ? 3'b000 : 3'b100;
							assign node108 = (inp[8]) ? node110 : 3'b000;
								assign node110 = (inp[3]) ? node116 : node111;
									assign node111 = (inp[2]) ? 3'b100 : node112;
										assign node112 = (inp[7]) ? 3'b000 : 3'b100;
									assign node116 = (inp[10]) ? node118 : 3'b000;
										assign node118 = (inp[2]) ? 3'b100 : 3'b000;
					assign node121 = (inp[8]) ? node163 : node122;
						assign node122 = (inp[1]) ? node144 : node123;
							assign node123 = (inp[7]) ? node135 : node124;
								assign node124 = (inp[10]) ? 3'b101 : node125;
									assign node125 = (inp[11]) ? node131 : node126;
										assign node126 = (inp[3]) ? 3'b001 : node127;
											assign node127 = (inp[2]) ? 3'b101 : 3'b001;
										assign node131 = (inp[2]) ? 3'b001 : 3'b100;
								assign node135 = (inp[11]) ? 3'b001 : node136;
									assign node136 = (inp[10]) ? node138 : 3'b001;
										assign node138 = (inp[2]) ? 3'b101 : node139;
											assign node139 = (inp[3]) ? 3'b101 : 3'b001;
							assign node144 = (inp[10]) ? node156 : node145;
								assign node145 = (inp[3]) ? node151 : node146;
									assign node146 = (inp[2]) ? 3'b100 : node147;
										assign node147 = (inp[5]) ? 3'b000 : 3'b100;
									assign node151 = (inp[11]) ? 3'b000 : node152;
										assign node152 = (inp[7]) ? 3'b000 : 3'b100;
								assign node156 = (inp[11]) ? node160 : node157;
									assign node157 = (inp[2]) ? 3'b101 : 3'b001;
									assign node160 = (inp[2]) ? 3'b001 : 3'b100;
						assign node163 = (inp[10]) ? node189 : node164;
							assign node164 = (inp[3]) ? node178 : node165;
								assign node165 = (inp[2]) ? node175 : node166;
									assign node166 = (inp[1]) ? node172 : node167;
										assign node167 = (inp[11]) ? node169 : 3'b000;
											assign node169 = (inp[7]) ? 3'b000 : 3'b100;
										assign node172 = (inp[11]) ? 3'b001 : 3'b101;
									assign node175 = (inp[1]) ? 3'b100 : 3'b101;
								assign node178 = (inp[2]) ? node186 : node179;
									assign node179 = (inp[1]) ? node183 : node180;
										assign node180 = (inp[11]) ? 3'b000 : 3'b100;
										assign node183 = (inp[11]) ? 3'b101 : 3'b001;
									assign node186 = (inp[1]) ? 3'b000 : 3'b001;
							assign node189 = (inp[2]) ? 3'b000 : node190;
								assign node190 = (inp[7]) ? node194 : node191;
									assign node191 = (inp[11]) ? 3'b110 : 3'b111;
									assign node194 = (inp[11]) ? 3'b010 : 3'b011;
			assign node198 = (inp[9]) ? node200 : 3'b000;
				assign node200 = (inp[1]) ? node260 : node201;
					assign node201 = (inp[8]) ? node227 : node202;
						assign node202 = (inp[4]) ? node212 : node203;
							assign node203 = (inp[11]) ? 3'b000 : node204;
								assign node204 = (inp[10]) ? 3'b100 : node205;
									assign node205 = (inp[7]) ? 3'b000 : node206;
										assign node206 = (inp[3]) ? 3'b000 : 3'b100;
							assign node212 = (inp[10]) ? node220 : node213;
								assign node213 = (inp[11]) ? 3'b100 : node214;
									assign node214 = (inp[3]) ? node216 : 3'b000;
										assign node216 = (inp[2]) ? 3'b000 : 3'b100;
								assign node220 = (inp[11]) ? 3'b000 : node221;
									assign node221 = (inp[2]) ? 3'b100 : node222;
										assign node222 = (inp[3]) ? 3'b000 : 3'b100;
						assign node227 = (inp[4]) ? node237 : node228;
							assign node228 = (inp[11]) ? node230 : 3'b100;
								assign node230 = (inp[10]) ? 3'b100 : node231;
									assign node231 = (inp[3]) ? 3'b000 : node232;
										assign node232 = (inp[7]) ? 3'b000 : 3'b100;
							assign node237 = (inp[10]) ? node251 : node238;
								assign node238 = (inp[3]) ? node246 : node239;
									assign node239 = (inp[2]) ? 3'b101 : node240;
										assign node240 = (inp[11]) ? 3'b100 : node241;
											assign node241 = (inp[7]) ? 3'b001 : 3'b101;
									assign node246 = (inp[11]) ? node248 : 3'b001;
										assign node248 = (inp[2]) ? 3'b001 : 3'b000;
								assign node251 = (inp[2]) ? 3'b000 : node252;
									assign node252 = (inp[11]) ? node256 : node253;
										assign node253 = (inp[7]) ? 3'b001 : 3'b101;
										assign node256 = (inp[7]) ? 3'b000 : 3'b100;
					assign node260 = (inp[4]) ? node262 : 3'b000;
						assign node262 = (inp[11]) ? node280 : node263;
							assign node263 = (inp[10]) ? node273 : node264;
								assign node264 = (inp[3]) ? node268 : node265;
									assign node265 = (inp[2]) ? 3'b100 : 3'b000;
									assign node268 = (inp[2]) ? 3'b000 : node269;
										assign node269 = (inp[8]) ? 3'b100 : 3'b000;
								assign node273 = (inp[8]) ? node275 : 3'b100;
									assign node275 = (inp[2]) ? 3'b000 : node276;
										assign node276 = (inp[3]) ? 3'b001 : 3'b101;
							assign node280 = (inp[8]) ? node282 : 3'b000;
								assign node282 = (inp[5]) ? node284 : 3'b000;
									assign node284 = (inp[10]) ? node286 : 3'b100;
										assign node286 = (inp[2]) ? 3'b000 : node287;
											assign node287 = (inp[7]) ? 3'b000 : 3'b100;

endmodule