module dtc_split66_bm28 (
	input  wire [7-1:0] inp,
	output wire [10-1:0] outp
);

	wire [10-1:0] node1;
	wire [10-1:0] node2;
	wire [10-1:0] node3;
	wire [10-1:0] node4;
	wire [10-1:0] node5;
	wire [10-1:0] node8;
	wire [10-1:0] node9;
	wire [10-1:0] node12;
	wire [10-1:0] node15;
	wire [10-1:0] node16;
	wire [10-1:0] node17;
	wire [10-1:0] node20;
	wire [10-1:0] node23;
	wire [10-1:0] node26;
	wire [10-1:0] node27;
	wire [10-1:0] node29;
	wire [10-1:0] node31;
	wire [10-1:0] node34;
	wire [10-1:0] node35;
	wire [10-1:0] node38;
	wire [10-1:0] node39;
	wire [10-1:0] node43;
	wire [10-1:0] node44;
	wire [10-1:0] node45;
	wire [10-1:0] node46;
	wire [10-1:0] node47;
	wire [10-1:0] node51;
	wire [10-1:0] node52;
	wire [10-1:0] node56;
	wire [10-1:0] node57;
	wire [10-1:0] node59;
	wire [10-1:0] node63;
	wire [10-1:0] node64;
	wire [10-1:0] node65;
	wire [10-1:0] node67;
	wire [10-1:0] node70;
	wire [10-1:0] node72;
	wire [10-1:0] node75;
	wire [10-1:0] node76;
	wire [10-1:0] node77;
	wire [10-1:0] node80;
	wire [10-1:0] node83;
	wire [10-1:0] node85;
	wire [10-1:0] node88;
	wire [10-1:0] node89;
	wire [10-1:0] node90;
	wire [10-1:0] node91;
	wire [10-1:0] node92;
	wire [10-1:0] node95;
	wire [10-1:0] node96;
	wire [10-1:0] node100;
	wire [10-1:0] node101;
	wire [10-1:0] node103;
	wire [10-1:0] node106;
	wire [10-1:0] node107;
	wire [10-1:0] node110;
	wire [10-1:0] node113;
	wire [10-1:0] node114;
	wire [10-1:0] node115;
	wire [10-1:0] node117;
	wire [10-1:0] node120;
	wire [10-1:0] node123;
	wire [10-1:0] node124;
	wire [10-1:0] node127;
	wire [10-1:0] node130;
	wire [10-1:0] node131;
	wire [10-1:0] node132;
	wire [10-1:0] node133;
	wire [10-1:0] node136;
	wire [10-1:0] node139;
	wire [10-1:0] node141;
	wire [10-1:0] node142;
	wire [10-1:0] node145;
	wire [10-1:0] node148;
	wire [10-1:0] node149;
	wire [10-1:0] node150;
	wire [10-1:0] node151;
	wire [10-1:0] node154;
	wire [10-1:0] node158;
	wire [10-1:0] node159;
	wire [10-1:0] node160;
	wire [10-1:0] node164;
	wire [10-1:0] node166;

	assign outp = (inp[4]) ? node88 : node1;
		assign node1 = (inp[2]) ? node43 : node2;
			assign node2 = (inp[5]) ? node26 : node3;
				assign node3 = (inp[3]) ? node15 : node4;
					assign node4 = (inp[6]) ? node8 : node5;
						assign node5 = (inp[0]) ? 10'b0011110001 : 10'b0001010101;
						assign node8 = (inp[1]) ? node12 : node9;
							assign node9 = (inp[0]) ? 10'b0011011000 : 10'b0111111000;
							assign node12 = (inp[0]) ? 10'b0001110000 : 10'b0111010000;
					assign node15 = (inp[1]) ? node23 : node16;
						assign node16 = (inp[6]) ? node20 : node17;
							assign node17 = (inp[0]) ? 10'b0101000001 : 10'b0001100101;
							assign node20 = (inp[0]) ? 10'b0011000000 : 10'b0111100000;
						assign node23 = (inp[0]) ? 10'b0001001001 : 10'b0001001100;
				assign node26 = (inp[3]) ? node34 : node27;
					assign node27 = (inp[6]) ? node29 : 10'b0010110000;
						assign node29 = (inp[1]) ? node31 : 10'b0110011001;
							assign node31 = (inp[0]) ? 10'b0000010001 : 10'b0100110001;
					assign node34 = (inp[0]) ? node38 : node35;
						assign node35 = (inp[6]) ? 10'b0100101000 : 10'b0110101001;
						assign node38 = (inp[1]) ? 10'b0000001000 : node39;
							assign node39 = (inp[6]) ? 10'b0000100001 : 10'b0100000000;
			assign node43 = (inp[3]) ? node63 : node44;
				assign node44 = (inp[5]) ? node56 : node45;
					assign node45 = (inp[6]) ? node51 : node46;
						assign node46 = (inp[0]) ? 10'b1010100001 : node47;
							assign node47 = (inp[1]) ? 10'b1000000101 : 10'b1000101101;
						assign node51 = (inp[0]) ? 10'b1000100000 : node52;
							assign node52 = (inp[1]) ? 10'b1110000000 : 10'b1110101000;
					assign node56 = (inp[1]) ? 10'b1101101000 : node57;
						assign node57 = (inp[6]) ? node59 : 10'b1101000000;
							assign node59 = (inp[0]) ? 10'b1001100001 : 10'b1111000001;
				assign node63 = (inp[5]) ? node75 : node64;
					assign node64 = (inp[6]) ? node70 : node65;
						assign node65 = (inp[1]) ? node67 : 10'b1101011000;
							assign node67 = (inp[0]) ? 10'b1011110000 : 10'b1001010100;
						assign node70 = (inp[0]) ? node72 : 10'b1101110001;
							assign node72 = (inp[1]) ? 10'b1001010001 : 10'b1001111001;
					assign node75 = (inp[6]) ? node83 : node76;
						assign node76 = (inp[1]) ? node80 : node77;
							assign node77 = (inp[0]) ? 10'b1010111001 : 10'b1000011101;
							assign node80 = (inp[0]) ? 10'b1010010001 : 10'b1110110001;
						assign node83 = (inp[1]) ? node85 : 10'b1110011000;
							assign node85 = (inp[0]) ? 10'b1000010000 : 10'b1100110000;
		assign node88 = (inp[3]) ? node130 : node89;
			assign node89 = (inp[2]) ? node113 : node90;
				assign node90 = (inp[5]) ? node100 : node91;
					assign node91 = (inp[6]) ? node95 : node92;
						assign node92 = (inp[1]) ? 10'b1000010111 : 10'b1000111111;
						assign node95 = (inp[1]) ? 10'b1000110010 : node96;
							assign node96 = (inp[0]) ? 10'b1010011010 : 10'b1110111010;
					assign node100 = (inp[1]) ? node106 : node101;
						assign node101 = (inp[6]) ? node103 : 10'b1001110110;
							assign node103 = (inp[0]) ? 10'b1001110011 : 10'b1111010011;
						assign node106 = (inp[0]) ? node110 : node107;
							assign node107 = (inp[6]) ? 10'b1101111010 : 10'b1111111011;
							assign node110 = (inp[6]) ? 10'b1001011010 : 10'b1011011011;
				assign node113 = (inp[5]) ? node123 : node114;
					assign node114 = (inp[1]) ? node120 : node115;
						assign node115 = (inp[6]) ? node117 : 10'b0101010011;
							assign node117 = (inp[0]) ? 10'b0011010010 : 10'b0111110010;
						assign node120 = (inp[6]) ? 10'b0001011011 : 10'b0001011110;
					assign node123 = (inp[1]) ? node127 : node124;
						assign node124 = (inp[0]) ? 10'b0000110011 : 10'b0110010011;
						assign node127 = (inp[6]) ? 10'b0100111010 : 10'b0110111011;
			assign node130 = (inp[2]) ? node148 : node131;
				assign node131 = (inp[5]) ? node139 : node132;
					assign node132 = (inp[1]) ? node136 : node133;
						assign node133 = (inp[6]) ? 10'b1010000010 : 10'b1100000011;
						assign node136 = (inp[0]) ? 10'b1010101010 : 10'b1000001110;
					assign node139 = (inp[6]) ? node141 : 10'b1011000011;
						assign node141 = (inp[1]) ? node145 : node142;
							assign node142 = (inp[0]) ? 10'b1001101010 : 10'b1111001010;
							assign node145 = (inp[0]) ? 10'b1001000010 : 10'b1101100010;
				assign node148 = (inp[5]) ? node158 : node149;
					assign node149 = (inp[6]) ? 10'b0101100011 : node150;
						assign node150 = (inp[1]) ? node154 : node151;
							assign node151 = (inp[0]) ? 10'b0101001010 : 10'b0001101110;
							assign node154 = (inp[0]) ? 10'b0011100010 : 10'b0001000110;
					assign node158 = (inp[6]) ? node164 : node159;
						assign node159 = (inp[1]) ? 10'b0110100011 : node160;
							assign node160 = (inp[0]) ? 10'b0010101011 : 10'b0000001111;
						assign node164 = (inp[0]) ? node166 : 10'b0110001010;
							assign node166 = (inp[1]) ? 10'b0000000010 : 10'b0000101010;

endmodule