module dtc_split33_bm56 (
	input  wire [12-1:0] inp,
	output wire [3-1:0] outp
);

	wire [3-1:0] node1;
	wire [3-1:0] node2;
	wire [3-1:0] node3;
	wire [3-1:0] node4;
	wire [3-1:0] node5;
	wire [3-1:0] node6;
	wire [3-1:0] node7;
	wire [3-1:0] node8;
	wire [3-1:0] node10;
	wire [3-1:0] node13;
	wire [3-1:0] node14;
	wire [3-1:0] node18;
	wire [3-1:0] node21;
	wire [3-1:0] node22;
	wire [3-1:0] node23;
	wire [3-1:0] node24;
	wire [3-1:0] node29;
	wire [3-1:0] node30;
	wire [3-1:0] node33;
	wire [3-1:0] node36;
	wire [3-1:0] node37;
	wire [3-1:0] node38;
	wire [3-1:0] node39;
	wire [3-1:0] node40;
	wire [3-1:0] node44;
	wire [3-1:0] node46;
	wire [3-1:0] node49;
	wire [3-1:0] node50;
	wire [3-1:0] node51;
	wire [3-1:0] node54;
	wire [3-1:0] node57;
	wire [3-1:0] node60;
	wire [3-1:0] node61;
	wire [3-1:0] node62;
	wire [3-1:0] node63;
	wire [3-1:0] node66;
	wire [3-1:0] node69;
	wire [3-1:0] node71;
	wire [3-1:0] node74;
	wire [3-1:0] node75;
	wire [3-1:0] node76;
	wire [3-1:0] node79;
	wire [3-1:0] node82;
	wire [3-1:0] node85;
	wire [3-1:0] node86;
	wire [3-1:0] node87;
	wire [3-1:0] node88;
	wire [3-1:0] node89;
	wire [3-1:0] node91;
	wire [3-1:0] node94;
	wire [3-1:0] node95;
	wire [3-1:0] node99;
	wire [3-1:0] node101;
	wire [3-1:0] node102;
	wire [3-1:0] node106;
	wire [3-1:0] node107;
	wire [3-1:0] node108;
	wire [3-1:0] node109;
	wire [3-1:0] node113;
	wire [3-1:0] node114;
	wire [3-1:0] node118;
	wire [3-1:0] node119;
	wire [3-1:0] node121;
	wire [3-1:0] node124;
	wire [3-1:0] node125;
	wire [3-1:0] node129;
	wire [3-1:0] node130;
	wire [3-1:0] node131;
	wire [3-1:0] node132;
	wire [3-1:0] node134;
	wire [3-1:0] node137;
	wire [3-1:0] node140;
	wire [3-1:0] node141;
	wire [3-1:0] node142;
	wire [3-1:0] node146;
	wire [3-1:0] node147;
	wire [3-1:0] node150;
	wire [3-1:0] node153;
	wire [3-1:0] node154;
	wire [3-1:0] node155;
	wire [3-1:0] node156;
	wire [3-1:0] node161;
	wire [3-1:0] node162;
	wire [3-1:0] node164;
	wire [3-1:0] node167;
	wire [3-1:0] node168;
	wire [3-1:0] node172;
	wire [3-1:0] node173;
	wire [3-1:0] node174;
	wire [3-1:0] node175;
	wire [3-1:0] node176;
	wire [3-1:0] node177;
	wire [3-1:0] node178;
	wire [3-1:0] node182;
	wire [3-1:0] node185;
	wire [3-1:0] node186;
	wire [3-1:0] node187;
	wire [3-1:0] node191;
	wire [3-1:0] node194;
	wire [3-1:0] node195;
	wire [3-1:0] node196;
	wire [3-1:0] node198;
	wire [3-1:0] node201;
	wire [3-1:0] node203;
	wire [3-1:0] node206;
	wire [3-1:0] node207;
	wire [3-1:0] node208;
	wire [3-1:0] node211;
	wire [3-1:0] node214;
	wire [3-1:0] node215;
	wire [3-1:0] node219;
	wire [3-1:0] node220;
	wire [3-1:0] node221;
	wire [3-1:0] node223;
	wire [3-1:0] node225;
	wire [3-1:0] node228;
	wire [3-1:0] node229;
	wire [3-1:0] node230;
	wire [3-1:0] node233;
	wire [3-1:0] node236;
	wire [3-1:0] node238;
	wire [3-1:0] node241;
	wire [3-1:0] node242;
	wire [3-1:0] node244;
	wire [3-1:0] node245;
	wire [3-1:0] node248;
	wire [3-1:0] node251;
	wire [3-1:0] node252;
	wire [3-1:0] node254;
	wire [3-1:0] node257;
	wire [3-1:0] node259;
	wire [3-1:0] node262;
	wire [3-1:0] node263;
	wire [3-1:0] node264;
	wire [3-1:0] node265;
	wire [3-1:0] node266;
	wire [3-1:0] node267;
	wire [3-1:0] node271;
	wire [3-1:0] node272;
	wire [3-1:0] node276;
	wire [3-1:0] node277;
	wire [3-1:0] node279;
	wire [3-1:0] node283;
	wire [3-1:0] node284;
	wire [3-1:0] node285;
	wire [3-1:0] node287;
	wire [3-1:0] node290;
	wire [3-1:0] node291;
	wire [3-1:0] node295;
	wire [3-1:0] node296;
	wire [3-1:0] node297;
	wire [3-1:0] node300;
	wire [3-1:0] node304;
	wire [3-1:0] node305;
	wire [3-1:0] node306;
	wire [3-1:0] node308;
	wire [3-1:0] node309;
	wire [3-1:0] node313;
	wire [3-1:0] node314;
	wire [3-1:0] node316;
	wire [3-1:0] node319;
	wire [3-1:0] node321;
	wire [3-1:0] node324;
	wire [3-1:0] node325;
	wire [3-1:0] node326;
	wire [3-1:0] node327;
	wire [3-1:0] node330;
	wire [3-1:0] node334;
	wire [3-1:0] node335;
	wire [3-1:0] node336;
	wire [3-1:0] node340;
	wire [3-1:0] node341;
	wire [3-1:0] node345;
	wire [3-1:0] node346;
	wire [3-1:0] node347;
	wire [3-1:0] node348;
	wire [3-1:0] node349;
	wire [3-1:0] node350;
	wire [3-1:0] node351;
	wire [3-1:0] node352;
	wire [3-1:0] node356;
	wire [3-1:0] node358;
	wire [3-1:0] node361;
	wire [3-1:0] node362;
	wire [3-1:0] node363;
	wire [3-1:0] node367;
	wire [3-1:0] node370;
	wire [3-1:0] node371;
	wire [3-1:0] node372;
	wire [3-1:0] node375;
	wire [3-1:0] node376;
	wire [3-1:0] node380;
	wire [3-1:0] node381;
	wire [3-1:0] node382;
	wire [3-1:0] node385;
	wire [3-1:0] node388;
	wire [3-1:0] node390;
	wire [3-1:0] node393;
	wire [3-1:0] node394;
	wire [3-1:0] node395;
	wire [3-1:0] node396;
	wire [3-1:0] node398;
	wire [3-1:0] node401;
	wire [3-1:0] node403;
	wire [3-1:0] node406;
	wire [3-1:0] node407;
	wire [3-1:0] node410;
	wire [3-1:0] node412;
	wire [3-1:0] node415;
	wire [3-1:0] node416;
	wire [3-1:0] node418;
	wire [3-1:0] node421;
	wire [3-1:0] node422;
	wire [3-1:0] node424;
	wire [3-1:0] node428;
	wire [3-1:0] node429;
	wire [3-1:0] node430;
	wire [3-1:0] node431;
	wire [3-1:0] node432;
	wire [3-1:0] node433;
	wire [3-1:0] node437;
	wire [3-1:0] node438;
	wire [3-1:0] node442;
	wire [3-1:0] node443;
	wire [3-1:0] node444;
	wire [3-1:0] node447;
	wire [3-1:0] node450;
	wire [3-1:0] node452;
	wire [3-1:0] node455;
	wire [3-1:0] node456;
	wire [3-1:0] node457;
	wire [3-1:0] node459;
	wire [3-1:0] node462;
	wire [3-1:0] node465;
	wire [3-1:0] node466;
	wire [3-1:0] node467;
	wire [3-1:0] node471;
	wire [3-1:0] node472;
	wire [3-1:0] node475;
	wire [3-1:0] node478;
	wire [3-1:0] node479;
	wire [3-1:0] node480;
	wire [3-1:0] node482;
	wire [3-1:0] node484;
	wire [3-1:0] node487;
	wire [3-1:0] node488;
	wire [3-1:0] node489;
	wire [3-1:0] node492;
	wire [3-1:0] node495;
	wire [3-1:0] node496;
	wire [3-1:0] node500;
	wire [3-1:0] node501;
	wire [3-1:0] node502;
	wire [3-1:0] node504;
	wire [3-1:0] node507;
	wire [3-1:0] node509;
	wire [3-1:0] node512;
	wire [3-1:0] node513;
	wire [3-1:0] node515;
	wire [3-1:0] node518;
	wire [3-1:0] node520;
	wire [3-1:0] node523;
	wire [3-1:0] node524;
	wire [3-1:0] node525;
	wire [3-1:0] node526;
	wire [3-1:0] node527;
	wire [3-1:0] node528;
	wire [3-1:0] node529;
	wire [3-1:0] node533;
	wire [3-1:0] node534;
	wire [3-1:0] node538;
	wire [3-1:0] node540;
	wire [3-1:0] node541;
	wire [3-1:0] node545;
	wire [3-1:0] node546;
	wire [3-1:0] node547;
	wire [3-1:0] node548;
	wire [3-1:0] node552;
	wire [3-1:0] node553;
	wire [3-1:0] node557;
	wire [3-1:0] node558;
	wire [3-1:0] node559;
	wire [3-1:0] node563;
	wire [3-1:0] node564;
	wire [3-1:0] node568;
	wire [3-1:0] node569;
	wire [3-1:0] node570;
	wire [3-1:0] node571;
	wire [3-1:0] node574;
	wire [3-1:0] node576;
	wire [3-1:0] node579;
	wire [3-1:0] node580;
	wire [3-1:0] node581;
	wire [3-1:0] node584;
	wire [3-1:0] node587;
	wire [3-1:0] node588;
	wire [3-1:0] node592;
	wire [3-1:0] node593;
	wire [3-1:0] node594;
	wire [3-1:0] node595;
	wire [3-1:0] node600;
	wire [3-1:0] node601;
	wire [3-1:0] node603;
	wire [3-1:0] node607;
	wire [3-1:0] node608;
	wire [3-1:0] node609;
	wire [3-1:0] node610;
	wire [3-1:0] node611;
	wire [3-1:0] node612;
	wire [3-1:0] node615;
	wire [3-1:0] node618;
	wire [3-1:0] node619;
	wire [3-1:0] node623;
	wire [3-1:0] node624;
	wire [3-1:0] node626;
	wire [3-1:0] node629;
	wire [3-1:0] node630;
	wire [3-1:0] node634;
	wire [3-1:0] node635;
	wire [3-1:0] node636;
	wire [3-1:0] node637;
	wire [3-1:0] node640;
	wire [3-1:0] node643;
	wire [3-1:0] node645;
	wire [3-1:0] node648;
	wire [3-1:0] node649;
	wire [3-1:0] node650;
	wire [3-1:0] node654;
	wire [3-1:0] node656;
	wire [3-1:0] node659;
	wire [3-1:0] node660;
	wire [3-1:0] node661;
	wire [3-1:0] node662;
	wire [3-1:0] node663;
	wire [3-1:0] node666;
	wire [3-1:0] node669;
	wire [3-1:0] node671;
	wire [3-1:0] node674;
	wire [3-1:0] node675;
	wire [3-1:0] node676;
	wire [3-1:0] node680;
	wire [3-1:0] node682;
	wire [3-1:0] node685;
	wire [3-1:0] node686;
	wire [3-1:0] node688;
	wire [3-1:0] node691;
	wire [3-1:0] node692;
	wire [3-1:0] node693;
	wire [3-1:0] node696;
	wire [3-1:0] node700;
	wire [3-1:0] node701;
	wire [3-1:0] node702;
	wire [3-1:0] node703;
	wire [3-1:0] node704;
	wire [3-1:0] node705;
	wire [3-1:0] node706;
	wire [3-1:0] node707;
	wire [3-1:0] node708;
	wire [3-1:0] node711;
	wire [3-1:0] node714;
	wire [3-1:0] node715;
	wire [3-1:0] node719;
	wire [3-1:0] node720;
	wire [3-1:0] node722;
	wire [3-1:0] node725;
	wire [3-1:0] node727;
	wire [3-1:0] node730;
	wire [3-1:0] node731;
	wire [3-1:0] node732;
	wire [3-1:0] node734;
	wire [3-1:0] node737;
	wire [3-1:0] node738;
	wire [3-1:0] node741;
	wire [3-1:0] node744;
	wire [3-1:0] node745;
	wire [3-1:0] node747;
	wire [3-1:0] node750;
	wire [3-1:0] node753;
	wire [3-1:0] node754;
	wire [3-1:0] node755;
	wire [3-1:0] node756;
	wire [3-1:0] node758;
	wire [3-1:0] node761;
	wire [3-1:0] node762;
	wire [3-1:0] node765;
	wire [3-1:0] node768;
	wire [3-1:0] node769;
	wire [3-1:0] node770;
	wire [3-1:0] node773;
	wire [3-1:0] node776;
	wire [3-1:0] node778;
	wire [3-1:0] node781;
	wire [3-1:0] node782;
	wire [3-1:0] node783;
	wire [3-1:0] node785;
	wire [3-1:0] node789;
	wire [3-1:0] node790;
	wire [3-1:0] node791;
	wire [3-1:0] node795;
	wire [3-1:0] node798;
	wire [3-1:0] node799;
	wire [3-1:0] node800;
	wire [3-1:0] node801;
	wire [3-1:0] node802;
	wire [3-1:0] node803;
	wire [3-1:0] node807;
	wire [3-1:0] node810;
	wire [3-1:0] node812;
	wire [3-1:0] node813;
	wire [3-1:0] node817;
	wire [3-1:0] node818;
	wire [3-1:0] node819;
	wire [3-1:0] node820;
	wire [3-1:0] node823;
	wire [3-1:0] node826;
	wire [3-1:0] node827;
	wire [3-1:0] node831;
	wire [3-1:0] node832;
	wire [3-1:0] node834;
	wire [3-1:0] node837;
	wire [3-1:0] node838;
	wire [3-1:0] node841;
	wire [3-1:0] node844;
	wire [3-1:0] node845;
	wire [3-1:0] node846;
	wire [3-1:0] node847;
	wire [3-1:0] node848;
	wire [3-1:0] node851;
	wire [3-1:0] node854;
	wire [3-1:0] node855;
	wire [3-1:0] node858;
	wire [3-1:0] node861;
	wire [3-1:0] node862;
	wire [3-1:0] node863;
	wire [3-1:0] node866;
	wire [3-1:0] node869;
	wire [3-1:0] node872;
	wire [3-1:0] node873;
	wire [3-1:0] node874;
	wire [3-1:0] node876;
	wire [3-1:0] node879;
	wire [3-1:0] node880;
	wire [3-1:0] node883;
	wire [3-1:0] node886;
	wire [3-1:0] node887;
	wire [3-1:0] node888;
	wire [3-1:0] node891;
	wire [3-1:0] node894;
	wire [3-1:0] node895;
	wire [3-1:0] node899;
	wire [3-1:0] node900;
	wire [3-1:0] node901;
	wire [3-1:0] node902;
	wire [3-1:0] node903;
	wire [3-1:0] node905;
	wire [3-1:0] node907;
	wire [3-1:0] node910;
	wire [3-1:0] node911;
	wire [3-1:0] node913;
	wire [3-1:0] node916;
	wire [3-1:0] node917;
	wire [3-1:0] node921;
	wire [3-1:0] node922;
	wire [3-1:0] node923;
	wire [3-1:0] node925;
	wire [3-1:0] node929;
	wire [3-1:0] node930;
	wire [3-1:0] node931;
	wire [3-1:0] node934;
	wire [3-1:0] node937;
	wire [3-1:0] node939;
	wire [3-1:0] node942;
	wire [3-1:0] node943;
	wire [3-1:0] node944;
	wire [3-1:0] node945;
	wire [3-1:0] node946;
	wire [3-1:0] node950;
	wire [3-1:0] node952;
	wire [3-1:0] node955;
	wire [3-1:0] node956;
	wire [3-1:0] node959;
	wire [3-1:0] node961;
	wire [3-1:0] node964;
	wire [3-1:0] node965;
	wire [3-1:0] node966;
	wire [3-1:0] node967;
	wire [3-1:0] node972;
	wire [3-1:0] node973;
	wire [3-1:0] node975;
	wire [3-1:0] node978;
	wire [3-1:0] node979;
	wire [3-1:0] node983;
	wire [3-1:0] node984;
	wire [3-1:0] node985;
	wire [3-1:0] node986;
	wire [3-1:0] node987;
	wire [3-1:0] node988;
	wire [3-1:0] node991;
	wire [3-1:0] node994;
	wire [3-1:0] node995;
	wire [3-1:0] node999;
	wire [3-1:0] node1000;
	wire [3-1:0] node1003;
	wire [3-1:0] node1004;
	wire [3-1:0] node1008;
	wire [3-1:0] node1009;
	wire [3-1:0] node1010;
	wire [3-1:0] node1012;
	wire [3-1:0] node1016;
	wire [3-1:0] node1017;
	wire [3-1:0] node1019;
	wire [3-1:0] node1022;
	wire [3-1:0] node1024;
	wire [3-1:0] node1027;
	wire [3-1:0] node1028;
	wire [3-1:0] node1029;
	wire [3-1:0] node1030;
	wire [3-1:0] node1031;
	wire [3-1:0] node1034;
	wire [3-1:0] node1037;
	wire [3-1:0] node1039;
	wire [3-1:0] node1042;
	wire [3-1:0] node1043;
	wire [3-1:0] node1044;
	wire [3-1:0] node1048;
	wire [3-1:0] node1051;
	wire [3-1:0] node1052;
	wire [3-1:0] node1053;
	wire [3-1:0] node1054;
	wire [3-1:0] node1058;
	wire [3-1:0] node1060;
	wire [3-1:0] node1063;
	wire [3-1:0] node1064;
	wire [3-1:0] node1065;
	wire [3-1:0] node1068;
	wire [3-1:0] node1072;
	wire [3-1:0] node1073;
	wire [3-1:0] node1074;
	wire [3-1:0] node1075;
	wire [3-1:0] node1076;
	wire [3-1:0] node1077;
	wire [3-1:0] node1078;
	wire [3-1:0] node1079;
	wire [3-1:0] node1082;
	wire [3-1:0] node1085;
	wire [3-1:0] node1086;
	wire [3-1:0] node1090;
	wire [3-1:0] node1091;
	wire [3-1:0] node1092;
	wire [3-1:0] node1095;
	wire [3-1:0] node1098;
	wire [3-1:0] node1099;
	wire [3-1:0] node1102;
	wire [3-1:0] node1105;
	wire [3-1:0] node1106;
	wire [3-1:0] node1107;
	wire [3-1:0] node1108;
	wire [3-1:0] node1112;
	wire [3-1:0] node1113;
	wire [3-1:0] node1116;
	wire [3-1:0] node1119;
	wire [3-1:0] node1120;
	wire [3-1:0] node1121;
	wire [3-1:0] node1124;
	wire [3-1:0] node1127;
	wire [3-1:0] node1130;
	wire [3-1:0] node1131;
	wire [3-1:0] node1132;
	wire [3-1:0] node1133;
	wire [3-1:0] node1134;
	wire [3-1:0] node1137;
	wire [3-1:0] node1140;
	wire [3-1:0] node1143;
	wire [3-1:0] node1144;
	wire [3-1:0] node1145;
	wire [3-1:0] node1149;
	wire [3-1:0] node1150;
	wire [3-1:0] node1154;
	wire [3-1:0] node1155;
	wire [3-1:0] node1156;
	wire [3-1:0] node1157;
	wire [3-1:0] node1162;
	wire [3-1:0] node1163;
	wire [3-1:0] node1166;
	wire [3-1:0] node1168;
	wire [3-1:0] node1171;
	wire [3-1:0] node1172;
	wire [3-1:0] node1173;
	wire [3-1:0] node1174;
	wire [3-1:0] node1175;
	wire [3-1:0] node1176;
	wire [3-1:0] node1179;
	wire [3-1:0] node1183;
	wire [3-1:0] node1184;
	wire [3-1:0] node1185;
	wire [3-1:0] node1189;
	wire [3-1:0] node1190;
	wire [3-1:0] node1193;
	wire [3-1:0] node1196;
	wire [3-1:0] node1197;
	wire [3-1:0] node1198;
	wire [3-1:0] node1199;
	wire [3-1:0] node1202;
	wire [3-1:0] node1205;
	wire [3-1:0] node1206;
	wire [3-1:0] node1209;
	wire [3-1:0] node1212;
	wire [3-1:0] node1213;
	wire [3-1:0] node1215;
	wire [3-1:0] node1218;
	wire [3-1:0] node1219;
	wire [3-1:0] node1223;
	wire [3-1:0] node1224;
	wire [3-1:0] node1225;
	wire [3-1:0] node1226;
	wire [3-1:0] node1227;
	wire [3-1:0] node1231;
	wire [3-1:0] node1233;
	wire [3-1:0] node1236;
	wire [3-1:0] node1237;
	wire [3-1:0] node1238;
	wire [3-1:0] node1242;
	wire [3-1:0] node1245;
	wire [3-1:0] node1246;
	wire [3-1:0] node1247;
	wire [3-1:0] node1248;
	wire [3-1:0] node1252;
	wire [3-1:0] node1253;
	wire [3-1:0] node1256;
	wire [3-1:0] node1259;
	wire [3-1:0] node1260;
	wire [3-1:0] node1261;
	wire [3-1:0] node1265;
	wire [3-1:0] node1267;
	wire [3-1:0] node1270;
	wire [3-1:0] node1271;
	wire [3-1:0] node1272;
	wire [3-1:0] node1273;
	wire [3-1:0] node1274;
	wire [3-1:0] node1275;
	wire [3-1:0] node1276;
	wire [3-1:0] node1279;
	wire [3-1:0] node1282;
	wire [3-1:0] node1283;
	wire [3-1:0] node1287;
	wire [3-1:0] node1288;
	wire [3-1:0] node1289;
	wire [3-1:0] node1293;
	wire [3-1:0] node1295;
	wire [3-1:0] node1298;
	wire [3-1:0] node1299;
	wire [3-1:0] node1300;
	wire [3-1:0] node1303;
	wire [3-1:0] node1306;
	wire [3-1:0] node1308;
	wire [3-1:0] node1309;
	wire [3-1:0] node1312;
	wire [3-1:0] node1315;
	wire [3-1:0] node1316;
	wire [3-1:0] node1317;
	wire [3-1:0] node1318;
	wire [3-1:0] node1320;
	wire [3-1:0] node1324;
	wire [3-1:0] node1325;
	wire [3-1:0] node1328;
	wire [3-1:0] node1329;
	wire [3-1:0] node1333;
	wire [3-1:0] node1334;
	wire [3-1:0] node1335;
	wire [3-1:0] node1336;
	wire [3-1:0] node1339;
	wire [3-1:0] node1342;
	wire [3-1:0] node1343;
	wire [3-1:0] node1346;
	wire [3-1:0] node1349;
	wire [3-1:0] node1350;
	wire [3-1:0] node1353;
	wire [3-1:0] node1354;
	wire [3-1:0] node1358;
	wire [3-1:0] node1359;
	wire [3-1:0] node1360;
	wire [3-1:0] node1361;
	wire [3-1:0] node1362;
	wire [3-1:0] node1364;
	wire [3-1:0] node1367;
	wire [3-1:0] node1369;
	wire [3-1:0] node1372;
	wire [3-1:0] node1373;
	wire [3-1:0] node1374;
	wire [3-1:0] node1377;
	wire [3-1:0] node1380;
	wire [3-1:0] node1381;
	wire [3-1:0] node1385;
	wire [3-1:0] node1386;
	wire [3-1:0] node1387;
	wire [3-1:0] node1388;
	wire [3-1:0] node1392;
	wire [3-1:0] node1394;
	wire [3-1:0] node1397;
	wire [3-1:0] node1398;
	wire [3-1:0] node1399;
	wire [3-1:0] node1402;
	wire [3-1:0] node1405;
	wire [3-1:0] node1408;
	wire [3-1:0] node1409;
	wire [3-1:0] node1410;
	wire [3-1:0] node1412;
	wire [3-1:0] node1413;
	wire [3-1:0] node1416;
	wire [3-1:0] node1419;
	wire [3-1:0] node1420;
	wire [3-1:0] node1423;
	wire [3-1:0] node1425;
	wire [3-1:0] node1428;
	wire [3-1:0] node1429;
	wire [3-1:0] node1430;
	wire [3-1:0] node1431;
	wire [3-1:0] node1434;
	wire [3-1:0] node1437;
	wire [3-1:0] node1438;
	wire [3-1:0] node1442;
	wire [3-1:0] node1443;
	wire [3-1:0] node1445;

	assign outp = (inp[3]) ? node700 : node1;
		assign node1 = (inp[4]) ? node345 : node2;
			assign node2 = (inp[8]) ? node172 : node3;
				assign node3 = (inp[5]) ? node85 : node4;
					assign node4 = (inp[2]) ? node36 : node5;
						assign node5 = (inp[10]) ? node21 : node6;
							assign node6 = (inp[9]) ? node18 : node7;
								assign node7 = (inp[7]) ? node13 : node8;
									assign node8 = (inp[11]) ? node10 : 3'b111;
										assign node10 = (inp[1]) ? 3'b111 : 3'b011;
									assign node13 = (inp[0]) ? 3'b010 : node14;
										assign node14 = (inp[6]) ? 3'b110 : 3'b010;
								assign node18 = (inp[7]) ? 3'b111 : 3'b010;
							assign node21 = (inp[6]) ? node29 : node22;
								assign node22 = (inp[1]) ? 3'b110 : node23;
									assign node23 = (inp[0]) ? 3'b010 : node24;
										assign node24 = (inp[7]) ? 3'b010 : 3'b011;
								assign node29 = (inp[7]) ? node33 : node30;
									assign node30 = (inp[9]) ? 3'b010 : 3'b011;
									assign node33 = (inp[9]) ? 3'b011 : 3'b010;
						assign node36 = (inp[9]) ? node60 : node37;
							assign node37 = (inp[7]) ? node49 : node38;
								assign node38 = (inp[0]) ? node44 : node39;
									assign node39 = (inp[1]) ? 3'b111 : node40;
										assign node40 = (inp[11]) ? 3'b111 : 3'b011;
									assign node44 = (inp[11]) ? node46 : 3'b110;
										assign node46 = (inp[1]) ? 3'b110 : 3'b010;
								assign node49 = (inp[0]) ? node57 : node50;
									assign node50 = (inp[1]) ? node54 : node51;
										assign node51 = (inp[11]) ? 3'b110 : 3'b110;
										assign node54 = (inp[6]) ? 3'b110 : 3'b010;
									assign node57 = (inp[1]) ? 3'b011 : 3'b111;
							assign node60 = (inp[6]) ? node74 : node61;
								assign node61 = (inp[10]) ? node69 : node62;
									assign node62 = (inp[11]) ? node66 : node63;
										assign node63 = (inp[1]) ? 3'b010 : 3'b111;
										assign node66 = (inp[0]) ? 3'b010 : 3'b011;
									assign node69 = (inp[0]) ? node71 : 3'b110;
										assign node71 = (inp[1]) ? 3'b110 : 3'b010;
								assign node74 = (inp[10]) ? node82 : node75;
									assign node75 = (inp[11]) ? node79 : node76;
										assign node76 = (inp[1]) ? 3'b110 : 3'b010;
										assign node79 = (inp[0]) ? 3'b110 : 3'b111;
									assign node82 = (inp[1]) ? 3'b011 : 3'b111;
					assign node85 = (inp[10]) ? node129 : node86;
						assign node86 = (inp[6]) ? node106 : node87;
							assign node87 = (inp[11]) ? node99 : node88;
								assign node88 = (inp[1]) ? node94 : node89;
									assign node89 = (inp[7]) ? node91 : 3'b110;
										assign node91 = (inp[0]) ? 3'b111 : 3'b110;
									assign node94 = (inp[0]) ? 3'b010 : node95;
										assign node95 = (inp[2]) ? 3'b010 : 3'b011;
								assign node99 = (inp[9]) ? node101 : 3'b011;
									assign node101 = (inp[7]) ? 3'b011 : node102;
										assign node102 = (inp[0]) ? 3'b011 : 3'b010;
							assign node106 = (inp[11]) ? node118 : node107;
								assign node107 = (inp[1]) ? node113 : node108;
									assign node108 = (inp[2]) ? 3'b010 : node109;
										assign node109 = (inp[9]) ? 3'b010 : 3'b010;
									assign node113 = (inp[9]) ? 3'b101 : node114;
										assign node114 = (inp[0]) ? 3'b100 : 3'b101;
								assign node118 = (inp[1]) ? node124 : node119;
									assign node119 = (inp[9]) ? node121 : 3'b101;
										assign node121 = (inp[2]) ? 3'b101 : 3'b100;
									assign node124 = (inp[9]) ? 3'b100 : node125;
										assign node125 = (inp[7]) ? 3'b100 : 3'b101;
						assign node129 = (inp[6]) ? node153 : node130;
							assign node130 = (inp[1]) ? node140 : node131;
								assign node131 = (inp[11]) ? node137 : node132;
									assign node132 = (inp[7]) ? node134 : 3'b010;
										assign node134 = (inp[9]) ? 3'b011 : 3'b010;
									assign node137 = (inp[2]) ? 3'b100 : 3'b101;
								assign node140 = (inp[7]) ? node146 : node141;
									assign node141 = (inp[9]) ? 3'b100 : node142;
										assign node142 = (inp[11]) ? 3'b101 : 3'b100;
									assign node146 = (inp[0]) ? node150 : node147;
										assign node147 = (inp[9]) ? 3'b101 : 3'b100;
										assign node150 = (inp[9]) ? 3'b100 : 3'b101;
							assign node153 = (inp[1]) ? node161 : node154;
								assign node154 = (inp[11]) ? 3'b001 : node155;
									assign node155 = (inp[2]) ? 3'b101 : node156;
										assign node156 = (inp[9]) ? 3'b101 : 3'b100;
								assign node161 = (inp[2]) ? node167 : node162;
									assign node162 = (inp[11]) ? node164 : 3'b001;
										assign node164 = (inp[0]) ? 3'b001 : 3'b000;
									assign node167 = (inp[11]) ? 3'b000 : node168;
										assign node168 = (inp[0]) ? 3'b000 : 3'b000;
				assign node172 = (inp[5]) ? node262 : node173;
					assign node173 = (inp[11]) ? node219 : node174;
						assign node174 = (inp[7]) ? node194 : node175;
							assign node175 = (inp[9]) ? node185 : node176;
								assign node176 = (inp[2]) ? node182 : node177;
									assign node177 = (inp[6]) ? 3'b001 : node178;
										assign node178 = (inp[0]) ? 3'b001 : 3'b101;
									assign node182 = (inp[0]) ? 3'b000 : 3'b001;
								assign node185 = (inp[2]) ? node191 : node186;
									assign node186 = (inp[1]) ? 3'b000 : node187;
										assign node187 = (inp[0]) ? 3'b100 : 3'b000;
									assign node191 = (inp[0]) ? 3'b001 : 3'b000;
							assign node194 = (inp[6]) ? node206 : node195;
								assign node195 = (inp[9]) ? node201 : node196;
									assign node196 = (inp[10]) ? node198 : 3'b101;
										assign node198 = (inp[1]) ? 3'b100 : 3'b000;
									assign node201 = (inp[1]) ? node203 : 3'b100;
										assign node203 = (inp[10]) ? 3'b101 : 3'b001;
								assign node206 = (inp[9]) ? node214 : node207;
									assign node207 = (inp[0]) ? node211 : node208;
										assign node208 = (inp[1]) ? 3'b000 : 3'b000;
										assign node211 = (inp[2]) ? 3'b001 : 3'b000;
									assign node214 = (inp[2]) ? 3'b000 : node215;
										assign node215 = (inp[10]) ? 3'b001 : 3'b001;
						assign node219 = (inp[6]) ? node241 : node220;
							assign node220 = (inp[10]) ? node228 : node221;
								assign node221 = (inp[0]) ? node223 : 3'b000;
									assign node223 = (inp[2]) ? node225 : 3'b000;
										assign node225 = (inp[1]) ? 3'b001 : 3'b000;
								assign node228 = (inp[0]) ? node236 : node229;
									assign node229 = (inp[2]) ? node233 : node230;
										assign node230 = (inp[7]) ? 3'b100 : 3'b100;
										assign node233 = (inp[9]) ? 3'b100 : 3'b101;
									assign node236 = (inp[7]) ? node238 : 3'b100;
										assign node238 = (inp[2]) ? 3'b100 : 3'b101;
							assign node241 = (inp[10]) ? node251 : node242;
								assign node242 = (inp[9]) ? node244 : 3'b101;
									assign node244 = (inp[7]) ? node248 : node245;
										assign node245 = (inp[0]) ? 3'b101 : 3'b100;
										assign node248 = (inp[0]) ? 3'b100 : 3'b101;
								assign node251 = (inp[1]) ? node257 : node252;
									assign node252 = (inp[0]) ? node254 : 3'b001;
										assign node254 = (inp[2]) ? 3'b000 : 3'b001;
									assign node257 = (inp[0]) ? node259 : 3'b000;
										assign node259 = (inp[7]) ? 3'b001 : 3'b000;
					assign node262 = (inp[6]) ? node304 : node263;
						assign node263 = (inp[10]) ? node283 : node264;
							assign node264 = (inp[11]) ? node276 : node265;
								assign node265 = (inp[1]) ? node271 : node266;
									assign node266 = (inp[2]) ? 3'b100 : node267;
										assign node267 = (inp[0]) ? 3'b100 : 3'b100;
									assign node271 = (inp[2]) ? 3'b000 : node272;
										assign node272 = (inp[9]) ? 3'b001 : 3'b000;
								assign node276 = (inp[7]) ? 3'b000 : node277;
									assign node277 = (inp[9]) ? node279 : 3'b001;
										assign node279 = (inp[0]) ? 3'b001 : 3'b000;
							assign node283 = (inp[11]) ? node295 : node284;
								assign node284 = (inp[1]) ? node290 : node285;
									assign node285 = (inp[7]) ? node287 : 3'b000;
										assign node287 = (inp[0]) ? 3'b001 : 3'b000;
									assign node290 = (inp[2]) ? 3'b110 : node291;
										assign node291 = (inp[7]) ? 3'b111 : 3'b110;
								assign node295 = (inp[2]) ? 3'b111 : node296;
									assign node296 = (inp[7]) ? node300 : node297;
										assign node297 = (inp[0]) ? 3'b110 : 3'b110;
										assign node300 = (inp[0]) ? 3'b110 : 3'b111;
						assign node304 = (inp[10]) ? node324 : node305;
							assign node305 = (inp[1]) ? node313 : node306;
								assign node306 = (inp[11]) ? node308 : 3'b000;
									assign node308 = (inp[2]) ? 3'b110 : node309;
										assign node309 = (inp[7]) ? 3'b110 : 3'b111;
								assign node313 = (inp[11]) ? node319 : node314;
									assign node314 = (inp[2]) ? node316 : 3'b111;
										assign node316 = (inp[0]) ? 3'b110 : 3'b111;
									assign node319 = (inp[7]) ? node321 : 3'b110;
										assign node321 = (inp[9]) ? 3'b110 : 3'b111;
							assign node324 = (inp[1]) ? node334 : node325;
								assign node325 = (inp[11]) ? 3'b010 : node326;
									assign node326 = (inp[0]) ? node330 : node327;
										assign node327 = (inp[2]) ? 3'b110 : 3'b110;
										assign node330 = (inp[9]) ? 3'b110 : 3'b111;
								assign node334 = (inp[2]) ? node340 : node335;
									assign node335 = (inp[0]) ? 3'b010 : node336;
										assign node336 = (inp[9]) ? 3'b011 : 3'b010;
									assign node340 = (inp[9]) ? 3'b010 : node341;
										assign node341 = (inp[7]) ? 3'b011 : 3'b010;
			assign node345 = (inp[8]) ? node523 : node346;
				assign node346 = (inp[5]) ? node428 : node347;
					assign node347 = (inp[6]) ? node393 : node348;
						assign node348 = (inp[10]) ? node370 : node349;
							assign node349 = (inp[11]) ? node361 : node350;
								assign node350 = (inp[1]) ? node356 : node351;
									assign node351 = (inp[2]) ? 3'b100 : node352;
										assign node352 = (inp[9]) ? 3'b100 : 3'b100;
									assign node356 = (inp[7]) ? node358 : 3'b000;
										assign node358 = (inp[0]) ? 3'b000 : 3'b001;
								assign node361 = (inp[2]) ? node367 : node362;
									assign node362 = (inp[0]) ? 3'b000 : node363;
										assign node363 = (inp[9]) ? 3'b001 : 3'b000;
									assign node367 = (inp[0]) ? 3'b001 : 3'b000;
							assign node370 = (inp[1]) ? node380 : node371;
								assign node371 = (inp[11]) ? node375 : node372;
									assign node372 = (inp[9]) ? 3'b000 : 3'b001;
									assign node375 = (inp[0]) ? 3'b101 : node376;
										assign node376 = (inp[9]) ? 3'b100 : 3'b101;
								assign node380 = (inp[0]) ? node388 : node381;
									assign node381 = (inp[7]) ? node385 : node382;
										assign node382 = (inp[9]) ? 3'b100 : 3'b101;
										assign node385 = (inp[9]) ? 3'b101 : 3'b100;
									assign node388 = (inp[2]) ? node390 : 3'b101;
										assign node390 = (inp[7]) ? 3'b101 : 3'b100;
						assign node393 = (inp[10]) ? node415 : node394;
							assign node394 = (inp[11]) ? node406 : node395;
								assign node395 = (inp[1]) ? node401 : node396;
									assign node396 = (inp[7]) ? node398 : 3'b001;
										assign node398 = (inp[2]) ? 3'b001 : 3'b000;
									assign node401 = (inp[7]) ? node403 : 3'b100;
										assign node403 = (inp[2]) ? 3'b101 : 3'b100;
								assign node406 = (inp[9]) ? node410 : node407;
									assign node407 = (inp[7]) ? 3'b100 : 3'b101;
									assign node410 = (inp[2]) ? node412 : 3'b100;
										assign node412 = (inp[7]) ? 3'b101 : 3'b100;
							assign node415 = (inp[0]) ? node421 : node416;
								assign node416 = (inp[9]) ? node418 : 3'b000;
									assign node418 = (inp[7]) ? 3'b001 : 3'b000;
								assign node421 = (inp[11]) ? 3'b000 : node422;
									assign node422 = (inp[1]) ? node424 : 3'b100;
										assign node424 = (inp[7]) ? 3'b000 : 3'b001;
					assign node428 = (inp[6]) ? node478 : node429;
						assign node429 = (inp[10]) ? node455 : node430;
							assign node430 = (inp[1]) ? node442 : node431;
								assign node431 = (inp[11]) ? node437 : node432;
									assign node432 = (inp[7]) ? 3'b100 : node433;
										assign node433 = (inp[9]) ? 3'b100 : 3'b101;
									assign node437 = (inp[7]) ? 3'b000 : node438;
										assign node438 = (inp[9]) ? 3'b000 : 3'b001;
								assign node442 = (inp[9]) ? node450 : node443;
									assign node443 = (inp[7]) ? node447 : node444;
										assign node444 = (inp[2]) ? 3'b000 : 3'b001;
										assign node447 = (inp[2]) ? 3'b001 : 3'b000;
									assign node450 = (inp[0]) ? node452 : 3'b000;
										assign node452 = (inp[2]) ? 3'b001 : 3'b000;
							assign node455 = (inp[11]) ? node465 : node456;
								assign node456 = (inp[1]) ? node462 : node457;
									assign node457 = (inp[2]) ? node459 : 3'b001;
										assign node459 = (inp[0]) ? 3'b001 : 3'b000;
									assign node462 = (inp[9]) ? 3'b111 : 3'b110;
								assign node465 = (inp[9]) ? node471 : node466;
									assign node466 = (inp[7]) ? 3'b111 : node467;
										assign node467 = (inp[2]) ? 3'b110 : 3'b111;
									assign node471 = (inp[7]) ? node475 : node472;
										assign node472 = (inp[0]) ? 3'b111 : 3'b110;
										assign node475 = (inp[1]) ? 3'b110 : 3'b110;
						assign node478 = (inp[10]) ? node500 : node479;
							assign node479 = (inp[11]) ? node487 : node480;
								assign node480 = (inp[1]) ? node482 : 3'b000;
									assign node482 = (inp[9]) ? node484 : 3'b110;
										assign node484 = (inp[2]) ? 3'b110 : 3'b111;
								assign node487 = (inp[1]) ? node495 : node488;
									assign node488 = (inp[7]) ? node492 : node489;
										assign node489 = (inp[0]) ? 3'b111 : 3'b110;
										assign node492 = (inp[2]) ? 3'b110 : 3'b111;
									assign node495 = (inp[9]) ? 3'b110 : node496;
										assign node496 = (inp[2]) ? 3'b110 : 3'b110;
							assign node500 = (inp[1]) ? node512 : node501;
								assign node501 = (inp[11]) ? node507 : node502;
									assign node502 = (inp[9]) ? node504 : 3'b110;
										assign node504 = (inp[2]) ? 3'b111 : 3'b110;
									assign node507 = (inp[9]) ? node509 : 3'b010;
										assign node509 = (inp[7]) ? 3'b010 : 3'b011;
								assign node512 = (inp[9]) ? node518 : node513;
									assign node513 = (inp[2]) ? node515 : 3'b011;
										assign node515 = (inp[7]) ? 3'b011 : 3'b010;
									assign node518 = (inp[2]) ? node520 : 3'b010;
										assign node520 = (inp[7]) ? 3'b010 : 3'b011;
				assign node523 = (inp[5]) ? node607 : node524;
					assign node524 = (inp[9]) ? node568 : node525;
						assign node525 = (inp[7]) ? node545 : node526;
							assign node526 = (inp[0]) ? node538 : node527;
								assign node527 = (inp[2]) ? node533 : node528;
									assign node528 = (inp[10]) ? 3'b011 : node529;
										assign node529 = (inp[6]) ? 3'b111 : 3'b011;
									assign node533 = (inp[1]) ? 3'b010 : node534;
										assign node534 = (inp[11]) ? 3'b110 : 3'b110;
								assign node538 = (inp[1]) ? node540 : 3'b110;
									assign node540 = (inp[10]) ? 3'b010 : node541;
										assign node541 = (inp[6]) ? 3'b110 : 3'b010;
							assign node545 = (inp[0]) ? node557 : node546;
								assign node546 = (inp[2]) ? node552 : node547;
									assign node547 = (inp[11]) ? 3'b010 : node548;
										assign node548 = (inp[6]) ? 3'b110 : 3'b010;
									assign node552 = (inp[1]) ? 3'b111 : node553;
										assign node553 = (inp[10]) ? 3'b111 : 3'b011;
								assign node557 = (inp[1]) ? node563 : node558;
									assign node558 = (inp[2]) ? 3'b111 : node559;
										assign node559 = (inp[10]) ? 3'b111 : 3'b011;
									assign node563 = (inp[2]) ? 3'b011 : node564;
										assign node564 = (inp[10]) ? 3'b111 : 3'b011;
						assign node568 = (inp[7]) ? node592 : node569;
							assign node569 = (inp[0]) ? node579 : node570;
								assign node570 = (inp[2]) ? node574 : node571;
									assign node571 = (inp[1]) ? 3'b110 : 3'b010;
									assign node574 = (inp[6]) ? node576 : 3'b011;
										assign node576 = (inp[11]) ? 3'b011 : 3'b111;
								assign node579 = (inp[2]) ? node587 : node580;
									assign node580 = (inp[10]) ? node584 : node581;
										assign node581 = (inp[6]) ? 3'b011 : 3'b011;
										assign node584 = (inp[11]) ? 3'b011 : 3'b011;
									assign node587 = (inp[1]) ? 3'b111 : node588;
										assign node588 = (inp[6]) ? 3'b011 : 3'b111;
							assign node592 = (inp[2]) ? node600 : node593;
								assign node593 = (inp[0]) ? 3'b110 : node594;
									assign node594 = (inp[11]) ? 3'b111 : node595;
										assign node595 = (inp[1]) ? 3'b111 : 3'b011;
								assign node600 = (inp[6]) ? 3'b110 : node601;
									assign node601 = (inp[10]) ? node603 : 3'b010;
										assign node603 = (inp[0]) ? 3'b110 : 3'b010;
					assign node607 = (inp[10]) ? node659 : node608;
						assign node608 = (inp[6]) ? node634 : node609;
							assign node609 = (inp[11]) ? node623 : node610;
								assign node610 = (inp[1]) ? node618 : node611;
									assign node611 = (inp[9]) ? node615 : node612;
										assign node612 = (inp[2]) ? 3'b110 : 3'b110;
										assign node615 = (inp[0]) ? 3'b110 : 3'b111;
									assign node618 = (inp[2]) ? 3'b010 : node619;
										assign node619 = (inp[7]) ? 3'b010 : 3'b011;
								assign node623 = (inp[1]) ? node629 : node624;
									assign node624 = (inp[7]) ? node626 : 3'b010;
										assign node626 = (inp[9]) ? 3'b010 : 3'b011;
									assign node629 = (inp[7]) ? 3'b011 : node630;
										assign node630 = (inp[2]) ? 3'b011 : 3'b010;
							assign node634 = (inp[1]) ? node648 : node635;
								assign node635 = (inp[11]) ? node643 : node636;
									assign node636 = (inp[9]) ? node640 : node637;
										assign node637 = (inp[7]) ? 3'b011 : 3'b010;
										assign node640 = (inp[7]) ? 3'b010 : 3'b011;
									assign node643 = (inp[7]) ? node645 : 3'b101;
										assign node645 = (inp[0]) ? 3'b100 : 3'b101;
								assign node648 = (inp[2]) ? node654 : node649;
									assign node649 = (inp[9]) ? 3'b101 : node650;
										assign node650 = (inp[7]) ? 3'b100 : 3'b100;
									assign node654 = (inp[11]) ? node656 : 3'b100;
										assign node656 = (inp[9]) ? 3'b100 : 3'b101;
						assign node659 = (inp[6]) ? node685 : node660;
							assign node660 = (inp[1]) ? node674 : node661;
								assign node661 = (inp[11]) ? node669 : node662;
									assign node662 = (inp[2]) ? node666 : node663;
										assign node663 = (inp[0]) ? 3'b011 : 3'b010;
										assign node666 = (inp[9]) ? 3'b010 : 3'b011;
									assign node669 = (inp[2]) ? node671 : 3'b101;
										assign node671 = (inp[9]) ? 3'b100 : 3'b100;
								assign node674 = (inp[11]) ? node680 : node675;
									assign node675 = (inp[0]) ? 3'b101 : node676;
										assign node676 = (inp[7]) ? 3'b101 : 3'b101;
									assign node680 = (inp[0]) ? node682 : 3'b101;
										assign node682 = (inp[9]) ? 3'b100 : 3'b100;
							assign node685 = (inp[11]) ? node691 : node686;
								assign node686 = (inp[1]) ? node688 : 3'b101;
									assign node688 = (inp[0]) ? 3'b001 : 3'b000;
								assign node691 = (inp[0]) ? 3'b000 : node692;
									assign node692 = (inp[2]) ? node696 : node693;
										assign node693 = (inp[1]) ? 3'b001 : 3'b000;
										assign node696 = (inp[7]) ? 3'b000 : 3'b001;
		assign node700 = (inp[9]) ? node1072 : node701;
			assign node701 = (inp[7]) ? node899 : node702;
				assign node702 = (inp[2]) ? node798 : node703;
					assign node703 = (inp[0]) ? node753 : node704;
						assign node704 = (inp[10]) ? node730 : node705;
							assign node705 = (inp[6]) ? node719 : node706;
								assign node706 = (inp[5]) ? node714 : node707;
									assign node707 = (inp[11]) ? node711 : node708;
										assign node708 = (inp[1]) ? 3'b001 : 3'b101;
										assign node711 = (inp[4]) ? 3'b001 : 3'b001;
									assign node714 = (inp[4]) ? 3'b001 : node715;
										assign node715 = (inp[8]) ? 3'b011 : 3'b001;
								assign node719 = (inp[11]) ? node725 : node720;
									assign node720 = (inp[1]) ? node722 : 3'b011;
										assign node722 = (inp[8]) ? 3'b111 : 3'b101;
									assign node725 = (inp[4]) ? node727 : 3'b101;
										assign node727 = (inp[8]) ? 3'b101 : 3'b111;
							assign node730 = (inp[6]) ? node744 : node731;
								assign node731 = (inp[11]) ? node737 : node732;
									assign node732 = (inp[1]) ? node734 : 3'b011;
										assign node734 = (inp[4]) ? 3'b111 : 3'b101;
									assign node737 = (inp[5]) ? node741 : node738;
										assign node738 = (inp[4]) ? 3'b101 : 3'b101;
										assign node741 = (inp[1]) ? 3'b101 : 3'b111;
								assign node744 = (inp[4]) ? node750 : node745;
									assign node745 = (inp[11]) ? node747 : 3'b101;
										assign node747 = (inp[8]) ? 3'b011 : 3'b001;
									assign node750 = (inp[8]) ? 3'b001 : 3'b011;
						assign node753 = (inp[4]) ? node781 : node754;
							assign node754 = (inp[8]) ? node768 : node755;
								assign node755 = (inp[1]) ? node761 : node756;
									assign node756 = (inp[5]) ? node758 : 3'b101;
										assign node758 = (inp[11]) ? 3'b101 : 3'b001;
									assign node761 = (inp[11]) ? node765 : node762;
										assign node762 = (inp[10]) ? 3'b001 : 3'b001;
										assign node765 = (inp[10]) ? 3'b001 : 3'b101;
								assign node768 = (inp[6]) ? node776 : node769;
									assign node769 = (inp[5]) ? node773 : node770;
										assign node770 = (inp[11]) ? 3'b000 : 3'b001;
										assign node773 = (inp[11]) ? 3'b110 : 3'b010;
									assign node776 = (inp[10]) ? node778 : 3'b110;
										assign node778 = (inp[11]) ? 3'b010 : 3'b110;
							assign node781 = (inp[8]) ? node789 : node782;
								assign node782 = (inp[10]) ? 3'b010 : node783;
									assign node783 = (inp[1]) ? node785 : 3'b001;
										assign node785 = (inp[6]) ? 3'b110 : 3'b000;
								assign node789 = (inp[5]) ? node795 : node790;
									assign node790 = (inp[10]) ? 3'b000 : node791;
										assign node791 = (inp[1]) ? 3'b010 : 3'b110;
									assign node795 = (inp[10]) ? 3'b100 : 3'b000;
					assign node798 = (inp[0]) ? node844 : node799;
						assign node799 = (inp[4]) ? node817 : node800;
							assign node800 = (inp[8]) ? node810 : node801;
								assign node801 = (inp[10]) ? node807 : node802;
									assign node802 = (inp[6]) ? 3'b101 : node803;
										assign node803 = (inp[5]) ? 3'b101 : 3'b011;
									assign node807 = (inp[1]) ? 3'b101 : 3'b001;
								assign node810 = (inp[1]) ? node812 : 3'b001;
									assign node812 = (inp[5]) ? 3'b010 : node813;
										assign node813 = (inp[6]) ? 3'b110 : 3'b000;
							assign node817 = (inp[8]) ? node831 : node818;
								assign node818 = (inp[10]) ? node826 : node819;
									assign node819 = (inp[5]) ? node823 : node820;
										assign node820 = (inp[6]) ? 3'b001 : 3'b101;
										assign node823 = (inp[1]) ? 3'b010 : 3'b010;
									assign node826 = (inp[5]) ? 3'b110 : node827;
										assign node827 = (inp[6]) ? 3'b010 : 3'b110;
								assign node831 = (inp[5]) ? node837 : node832;
									assign node832 = (inp[11]) ? node834 : 3'b110;
										assign node834 = (inp[1]) ? 3'b000 : 3'b100;
									assign node837 = (inp[1]) ? node841 : node838;
										assign node838 = (inp[10]) ? 3'b000 : 3'b000;
										assign node841 = (inp[10]) ? 3'b000 : 3'b100;
						assign node844 = (inp[5]) ? node872 : node845;
							assign node845 = (inp[10]) ? node861 : node846;
								assign node846 = (inp[6]) ? node854 : node847;
									assign node847 = (inp[1]) ? node851 : node848;
										assign node848 = (inp[11]) ? 3'b000 : 3'b100;
										assign node851 = (inp[11]) ? 3'b000 : 3'b000;
									assign node854 = (inp[11]) ? node858 : node855;
										assign node855 = (inp[1]) ? 3'b100 : 3'b010;
										assign node858 = (inp[1]) ? 3'b110 : 3'b100;
								assign node861 = (inp[1]) ? node869 : node862;
									assign node862 = (inp[8]) ? node866 : node863;
										assign node863 = (inp[4]) ? 3'b000 : 3'b010;
										assign node866 = (inp[4]) ? 3'b010 : 3'b000;
									assign node869 = (inp[6]) ? 3'b000 : 3'b100;
							assign node872 = (inp[11]) ? node886 : node873;
								assign node873 = (inp[10]) ? node879 : node874;
									assign node874 = (inp[4]) ? node876 : 3'b110;
										assign node876 = (inp[8]) ? 3'b100 : 3'b110;
									assign node879 = (inp[1]) ? node883 : node880;
										assign node880 = (inp[4]) ? 3'b100 : 3'b000;
										assign node883 = (inp[6]) ? 3'b010 : 3'b100;
								assign node886 = (inp[4]) ? node894 : node887;
									assign node887 = (inp[8]) ? node891 : node888;
										assign node888 = (inp[10]) ? 3'b100 : 3'b000;
										assign node891 = (inp[10]) ? 3'b010 : 3'b110;
									assign node894 = (inp[8]) ? 3'b000 : node895;
										assign node895 = (inp[10]) ? 3'b110 : 3'b010;
				assign node899 = (inp[2]) ? node983 : node900;
					assign node900 = (inp[0]) ? node942 : node901;
						assign node901 = (inp[11]) ? node921 : node902;
							assign node902 = (inp[8]) ? node910 : node903;
								assign node903 = (inp[1]) ? node905 : 3'b110;
									assign node905 = (inp[5]) ? node907 : 3'b010;
										assign node907 = (inp[6]) ? 3'b110 : 3'b010;
								assign node910 = (inp[4]) ? node916 : node911;
									assign node911 = (inp[5]) ? node913 : 3'b110;
										assign node913 = (inp[1]) ? 3'b110 : 3'b010;
									assign node916 = (inp[10]) ? 3'b100 : node917;
										assign node917 = (inp[1]) ? 3'b100 : 3'b110;
							assign node921 = (inp[10]) ? node929 : node922;
								assign node922 = (inp[6]) ? 3'b110 : node923;
									assign node923 = (inp[1]) ? node925 : 3'b000;
										assign node925 = (inp[8]) ? 3'b010 : 3'b000;
								assign node929 = (inp[6]) ? node937 : node930;
									assign node930 = (inp[5]) ? node934 : node931;
										assign node931 = (inp[1]) ? 3'b100 : 3'b100;
										assign node934 = (inp[1]) ? 3'b100 : 3'b110;
									assign node937 = (inp[5]) ? node939 : 3'b000;
										assign node939 = (inp[4]) ? 3'b010 : 3'b000;
						assign node942 = (inp[4]) ? node964 : node943;
							assign node943 = (inp[8]) ? node955 : node944;
								assign node944 = (inp[1]) ? node950 : node945;
									assign node945 = (inp[5]) ? 3'b000 : node946;
										assign node946 = (inp[6]) ? 3'b000 : 3'b010;
									assign node950 = (inp[10]) ? node952 : 3'b100;
										assign node952 = (inp[6]) ? 3'b000 : 3'b100;
								assign node955 = (inp[5]) ? node959 : node956;
									assign node956 = (inp[10]) ? 3'b111 : 3'b000;
									assign node959 = (inp[6]) ? node961 : 3'b011;
										assign node961 = (inp[10]) ? 3'b011 : 3'b111;
							assign node964 = (inp[8]) ? node972 : node965;
								assign node965 = (inp[10]) ? 3'b111 : node966;
									assign node966 = (inp[6]) ? 3'b111 : node967;
										assign node967 = (inp[11]) ? 3'b000 : 3'b011;
								assign node972 = (inp[5]) ? node978 : node973;
									assign node973 = (inp[10]) ? node975 : 3'b011;
										assign node975 = (inp[11]) ? 3'b001 : 3'b101;
									assign node978 = (inp[1]) ? 3'b101 : node979;
										assign node979 = (inp[6]) ? 3'b001 : 3'b001;
					assign node983 = (inp[0]) ? node1027 : node984;
						assign node984 = (inp[8]) ? node1008 : node985;
							assign node985 = (inp[4]) ? node999 : node986;
								assign node986 = (inp[11]) ? node994 : node987;
									assign node987 = (inp[6]) ? node991 : node988;
										assign node988 = (inp[10]) ? 3'b010 : 3'b010;
										assign node991 = (inp[10]) ? 3'b100 : 3'b000;
									assign node994 = (inp[1]) ? 3'b000 : node995;
										assign node995 = (inp[6]) ? 3'b000 : 3'b100;
								assign node999 = (inp[10]) ? node1003 : node1000;
									assign node1000 = (inp[1]) ? 3'b111 : 3'b011;
									assign node1003 = (inp[1]) ? 3'b011 : node1004;
										assign node1004 = (inp[5]) ? 3'b011 : 3'b011;
							assign node1008 = (inp[4]) ? node1016 : node1009;
								assign node1009 = (inp[6]) ? 3'b111 : node1010;
									assign node1010 = (inp[10]) ? node1012 : 3'b011;
										assign node1012 = (inp[1]) ? 3'b111 : 3'b011;
								assign node1016 = (inp[11]) ? node1022 : node1017;
									assign node1017 = (inp[5]) ? node1019 : 3'b011;
										assign node1019 = (inp[10]) ? 3'b001 : 3'b101;
									assign node1022 = (inp[5]) ? node1024 : 3'b101;
										assign node1024 = (inp[1]) ? 3'b001 : 3'b101;
						assign node1027 = (inp[8]) ? node1051 : node1028;
							assign node1028 = (inp[4]) ? node1042 : node1029;
								assign node1029 = (inp[10]) ? node1037 : node1030;
									assign node1030 = (inp[5]) ? node1034 : node1031;
										assign node1031 = (inp[1]) ? 3'b101 : 3'b011;
										assign node1034 = (inp[6]) ? 3'b101 : 3'b001;
									assign node1037 = (inp[6]) ? node1039 : 3'b101;
										assign node1039 = (inp[11]) ? 3'b001 : 3'b101;
								assign node1042 = (inp[6]) ? node1048 : node1043;
									assign node1043 = (inp[5]) ? 3'b111 : node1044;
										assign node1044 = (inp[11]) ? 3'b111 : 3'b001;
									assign node1048 = (inp[10]) ? 3'b011 : 3'b001;
							assign node1051 = (inp[4]) ? node1063 : node1052;
								assign node1052 = (inp[10]) ? node1058 : node1053;
									assign node1053 = (inp[11]) ? 3'b001 : node1054;
										assign node1054 = (inp[5]) ? 3'b011 : 3'b111;
									assign node1058 = (inp[6]) ? node1060 : 3'b111;
										assign node1060 = (inp[1]) ? 3'b011 : 3'b111;
								assign node1063 = (inp[1]) ? 3'b101 : node1064;
									assign node1064 = (inp[5]) ? node1068 : node1065;
										assign node1065 = (inp[6]) ? 3'b101 : 3'b011;
										assign node1068 = (inp[10]) ? 3'b001 : 3'b001;
			assign node1072 = (inp[7]) ? node1270 : node1073;
				assign node1073 = (inp[2]) ? node1171 : node1074;
					assign node1074 = (inp[0]) ? node1130 : node1075;
						assign node1075 = (inp[1]) ? node1105 : node1076;
							assign node1076 = (inp[5]) ? node1090 : node1077;
								assign node1077 = (inp[10]) ? node1085 : node1078;
									assign node1078 = (inp[8]) ? node1082 : node1079;
										assign node1079 = (inp[6]) ? 3'b010 : 3'b110;
										assign node1082 = (inp[4]) ? 3'b010 : 3'b000;
									assign node1085 = (inp[11]) ? 3'b100 : node1086;
										assign node1086 = (inp[6]) ? 3'b100 : 3'b010;
								assign node1090 = (inp[11]) ? node1098 : node1091;
									assign node1091 = (inp[8]) ? node1095 : node1092;
										assign node1092 = (inp[10]) ? 3'b000 : 3'b000;
										assign node1095 = (inp[4]) ? 3'b000 : 3'b110;
									assign node1098 = (inp[4]) ? node1102 : node1099;
										assign node1099 = (inp[8]) ? 3'b110 : 3'b000;
										assign node1102 = (inp[8]) ? 3'b000 : 3'b010;
							assign node1105 = (inp[10]) ? node1119 : node1106;
								assign node1106 = (inp[6]) ? node1112 : node1107;
									assign node1107 = (inp[11]) ? 3'b000 : node1108;
										assign node1108 = (inp[5]) ? 3'b010 : 3'b000;
									assign node1112 = (inp[8]) ? node1116 : node1113;
										assign node1113 = (inp[4]) ? 3'b110 : 3'b100;
										assign node1116 = (inp[4]) ? 3'b100 : 3'b110;
								assign node1119 = (inp[6]) ? node1127 : node1120;
									assign node1120 = (inp[4]) ? node1124 : node1121;
										assign node1121 = (inp[8]) ? 3'b110 : 3'b100;
										assign node1124 = (inp[8]) ? 3'b100 : 3'b110;
									assign node1127 = (inp[11]) ? 3'b000 : 3'b010;
						assign node1130 = (inp[8]) ? node1154 : node1131;
							assign node1131 = (inp[4]) ? node1143 : node1132;
								assign node1132 = (inp[6]) ? node1140 : node1133;
									assign node1133 = (inp[5]) ? node1137 : node1134;
										assign node1134 = (inp[11]) ? 3'b010 : 3'b110;
										assign node1137 = (inp[10]) ? 3'b100 : 3'b000;
									assign node1140 = (inp[10]) ? 3'b000 : 3'b100;
								assign node1143 = (inp[11]) ? node1149 : node1144;
									assign node1144 = (inp[5]) ? 3'b011 : node1145;
										assign node1145 = (inp[6]) ? 3'b000 : 3'b000;
									assign node1149 = (inp[10]) ? 3'b111 : node1150;
										assign node1150 = (inp[1]) ? 3'b011 : 3'b111;
							assign node1154 = (inp[4]) ? node1162 : node1155;
								assign node1155 = (inp[1]) ? 3'b111 : node1156;
									assign node1156 = (inp[5]) ? 3'b011 : node1157;
										assign node1157 = (inp[10]) ? 3'b011 : 3'b111;
								assign node1162 = (inp[10]) ? node1166 : node1163;
									assign node1163 = (inp[1]) ? 3'b011 : 3'b111;
									assign node1166 = (inp[1]) ? node1168 : 3'b101;
										assign node1168 = (inp[6]) ? 3'b001 : 3'b101;
					assign node1171 = (inp[0]) ? node1223 : node1172;
						assign node1172 = (inp[4]) ? node1196 : node1173;
							assign node1173 = (inp[8]) ? node1183 : node1174;
								assign node1174 = (inp[1]) ? 3'b100 : node1175;
									assign node1175 = (inp[5]) ? node1179 : node1176;
										assign node1176 = (inp[10]) ? 3'b000 : 3'b010;
										assign node1179 = (inp[10]) ? 3'b000 : 3'b100;
								assign node1183 = (inp[5]) ? node1189 : node1184;
									assign node1184 = (inp[6]) ? 3'b111 : node1185;
										assign node1185 = (inp[10]) ? 3'b111 : 3'b100;
									assign node1189 = (inp[10]) ? node1193 : node1190;
										assign node1190 = (inp[11]) ? 3'b011 : 3'b111;
										assign node1193 = (inp[11]) ? 3'b011 : 3'b011;
							assign node1196 = (inp[8]) ? node1212 : node1197;
								assign node1197 = (inp[5]) ? node1205 : node1198;
									assign node1198 = (inp[6]) ? node1202 : node1199;
										assign node1199 = (inp[10]) ? 3'b000 : 3'b100;
										assign node1202 = (inp[10]) ? 3'b011 : 3'b111;
									assign node1205 = (inp[11]) ? node1209 : node1206;
										assign node1206 = (inp[1]) ? 3'b011 : 3'b011;
										assign node1209 = (inp[10]) ? 3'b111 : 3'b011;
								assign node1212 = (inp[5]) ? node1218 : node1213;
									assign node1213 = (inp[10]) ? node1215 : 3'b011;
										assign node1215 = (inp[11]) ? 3'b001 : 3'b011;
									assign node1218 = (inp[1]) ? 3'b001 : node1219;
										assign node1219 = (inp[11]) ? 3'b001 : 3'b101;
						assign node1223 = (inp[1]) ? node1245 : node1224;
							assign node1224 = (inp[4]) ? node1236 : node1225;
								assign node1225 = (inp[10]) ? node1231 : node1226;
									assign node1226 = (inp[5]) ? 3'b111 : node1227;
										assign node1227 = (inp[11]) ? 3'b001 : 3'b001;
									assign node1231 = (inp[8]) ? node1233 : 3'b101;
										assign node1233 = (inp[11]) ? 3'b111 : 3'b111;
								assign node1236 = (inp[8]) ? node1242 : node1237;
									assign node1237 = (inp[5]) ? 3'b011 : node1238;
										assign node1238 = (inp[11]) ? 3'b111 : 3'b001;
									assign node1242 = (inp[6]) ? 3'b101 : 3'b001;
							assign node1245 = (inp[5]) ? node1259 : node1246;
								assign node1246 = (inp[6]) ? node1252 : node1247;
									assign node1247 = (inp[10]) ? 3'b111 : node1248;
										assign node1248 = (inp[4]) ? 3'b001 : 3'b011;
									assign node1252 = (inp[10]) ? node1256 : node1253;
										assign node1253 = (inp[11]) ? 3'b111 : 3'b101;
										assign node1256 = (inp[8]) ? 3'b001 : 3'b001;
								assign node1259 = (inp[10]) ? node1265 : node1260;
									assign node1260 = (inp[6]) ? 3'b111 : node1261;
										assign node1261 = (inp[11]) ? 3'b011 : 3'b001;
									assign node1265 = (inp[6]) ? node1267 : 3'b101;
										assign node1267 = (inp[4]) ? 3'b001 : 3'b001;
				assign node1270 = (inp[2]) ? node1358 : node1271;
					assign node1271 = (inp[0]) ? node1315 : node1272;
						assign node1272 = (inp[11]) ? node1298 : node1273;
							assign node1273 = (inp[4]) ? node1287 : node1274;
								assign node1274 = (inp[10]) ? node1282 : node1275;
									assign node1275 = (inp[6]) ? node1279 : node1276;
										assign node1276 = (inp[1]) ? 3'b011 : 3'b111;
										assign node1279 = (inp[1]) ? 3'b101 : 3'b011;
									assign node1282 = (inp[6]) ? 3'b101 : node1283;
										assign node1283 = (inp[5]) ? 3'b011 : 3'b001;
								assign node1287 = (inp[8]) ? node1293 : node1288;
									assign node1288 = (inp[6]) ? 3'b111 : node1289;
										assign node1289 = (inp[10]) ? 3'b001 : 3'b101;
									assign node1293 = (inp[6]) ? node1295 : 3'b101;
										assign node1295 = (inp[10]) ? 3'b101 : 3'b001;
							assign node1298 = (inp[1]) ? node1306 : node1299;
								assign node1299 = (inp[10]) ? node1303 : node1300;
									assign node1300 = (inp[6]) ? 3'b111 : 3'b011;
									assign node1303 = (inp[5]) ? 3'b011 : 3'b001;
								assign node1306 = (inp[6]) ? node1308 : 3'b101;
									assign node1308 = (inp[10]) ? node1312 : node1309;
										assign node1309 = (inp[4]) ? 3'b101 : 3'b101;
										assign node1312 = (inp[5]) ? 3'b011 : 3'b011;
						assign node1315 = (inp[8]) ? node1333 : node1316;
							assign node1316 = (inp[4]) ? node1324 : node1317;
								assign node1317 = (inp[1]) ? 3'b001 : node1318;
									assign node1318 = (inp[11]) ? node1320 : 3'b101;
										assign node1320 = (inp[6]) ? 3'b001 : 3'b101;
								assign node1324 = (inp[5]) ? node1328 : node1325;
									assign node1325 = (inp[6]) ? 3'b110 : 3'b001;
									assign node1328 = (inp[10]) ? 3'b110 : node1329;
										assign node1329 = (inp[11]) ? 3'b110 : 3'b010;
							assign node1333 = (inp[4]) ? node1349 : node1334;
								assign node1334 = (inp[5]) ? node1342 : node1335;
									assign node1335 = (inp[10]) ? node1339 : node1336;
										assign node1336 = (inp[11]) ? 3'b110 : 3'b001;
										assign node1339 = (inp[11]) ? 3'b010 : 3'b110;
									assign node1342 = (inp[11]) ? node1346 : node1343;
										assign node1343 = (inp[1]) ? 3'b010 : 3'b010;
										assign node1346 = (inp[1]) ? 3'b010 : 3'b110;
								assign node1349 = (inp[5]) ? node1353 : node1350;
									assign node1350 = (inp[6]) ? 3'b000 : 3'b010;
									assign node1353 = (inp[1]) ? 3'b100 : node1354;
										assign node1354 = (inp[10]) ? 3'b100 : 3'b000;
					assign node1358 = (inp[0]) ? node1408 : node1359;
						assign node1359 = (inp[4]) ? node1385 : node1360;
							assign node1360 = (inp[8]) ? node1372 : node1361;
								assign node1361 = (inp[10]) ? node1367 : node1362;
									assign node1362 = (inp[5]) ? node1364 : 3'b011;
										assign node1364 = (inp[6]) ? 3'b101 : 3'b001;
									assign node1367 = (inp[11]) ? node1369 : 3'b101;
										assign node1369 = (inp[6]) ? 3'b001 : 3'b101;
								assign node1372 = (inp[5]) ? node1380 : node1373;
									assign node1373 = (inp[6]) ? node1377 : node1374;
										assign node1374 = (inp[1]) ? 3'b110 : 3'b001;
										assign node1377 = (inp[11]) ? 3'b110 : 3'b010;
									assign node1380 = (inp[10]) ? 3'b110 : node1381;
										assign node1381 = (inp[6]) ? 3'b110 : 3'b010;
							assign node1385 = (inp[8]) ? node1397 : node1386;
								assign node1386 = (inp[5]) ? node1392 : node1387;
									assign node1387 = (inp[10]) ? 3'b110 : node1388;
										assign node1388 = (inp[1]) ? 3'b110 : 3'b001;
									assign node1392 = (inp[11]) ? node1394 : 3'b110;
										assign node1394 = (inp[10]) ? 3'b010 : 3'b110;
								assign node1397 = (inp[5]) ? node1405 : node1398;
									assign node1398 = (inp[6]) ? node1402 : node1399;
										assign node1399 = (inp[1]) ? 3'b010 : 3'b010;
										assign node1402 = (inp[1]) ? 3'b100 : 3'b010;
									assign node1405 = (inp[11]) ? 3'b000 : 3'b100;
						assign node1408 = (inp[11]) ? node1428 : node1409;
							assign node1409 = (inp[4]) ? node1419 : node1410;
								assign node1410 = (inp[8]) ? node1412 : 3'b100;
									assign node1412 = (inp[6]) ? node1416 : node1413;
										assign node1413 = (inp[5]) ? 3'b110 : 3'b100;
										assign node1416 = (inp[5]) ? 3'b110 : 3'b110;
								assign node1419 = (inp[8]) ? node1423 : node1420;
									assign node1420 = (inp[1]) ? 3'b110 : 3'b010;
									assign node1423 = (inp[5]) ? node1425 : 3'b100;
										assign node1425 = (inp[10]) ? 3'b000 : 3'b100;
							assign node1428 = (inp[10]) ? node1442 : node1429;
								assign node1429 = (inp[6]) ? node1437 : node1430;
									assign node1430 = (inp[1]) ? node1434 : node1431;
										assign node1431 = (inp[4]) ? 3'b000 : 3'b010;
										assign node1434 = (inp[5]) ? 3'b000 : 3'b010;
									assign node1437 = (inp[5]) ? 3'b110 : node1438;
										assign node1438 = (inp[4]) ? 3'b100 : 3'b100;
								assign node1442 = (inp[6]) ? 3'b010 : node1443;
									assign node1443 = (inp[8]) ? node1445 : 3'b110;
										assign node1445 = (inp[4]) ? 3'b100 : 3'b110;

endmodule