module dtc_split25_bm90 (
	input  wire [12-1:0] inp,
	output wire [3-1:0] outp
);

	wire [3-1:0] node1;
	wire [3-1:0] node2;
	wire [3-1:0] node3;
	wire [3-1:0] node5;
	wire [3-1:0] node7;
	wire [3-1:0] node9;
	wire [3-1:0] node11;
	wire [3-1:0] node13;
	wire [3-1:0] node16;
	wire [3-1:0] node17;
	wire [3-1:0] node19;
	wire [3-1:0] node20;
	wire [3-1:0] node21;
	wire [3-1:0] node23;
	wire [3-1:0] node27;
	wire [3-1:0] node28;
	wire [3-1:0] node29;
	wire [3-1:0] node33;
	wire [3-1:0] node34;
	wire [3-1:0] node37;
	wire [3-1:0] node38;
	wire [3-1:0] node43;
	wire [3-1:0] node44;
	wire [3-1:0] node45;
	wire [3-1:0] node46;
	wire [3-1:0] node47;
	wire [3-1:0] node48;
	wire [3-1:0] node49;
	wire [3-1:0] node50;
	wire [3-1:0] node52;
	wire [3-1:0] node57;
	wire [3-1:0] node58;
	wire [3-1:0] node59;
	wire [3-1:0] node63;
	wire [3-1:0] node66;
	wire [3-1:0] node67;
	wire [3-1:0] node68;
	wire [3-1:0] node70;
	wire [3-1:0] node72;
	wire [3-1:0] node76;
	wire [3-1:0] node78;
	wire [3-1:0] node81;
	wire [3-1:0] node82;
	wire [3-1:0] node83;
	wire [3-1:0] node84;
	wire [3-1:0] node88;
	wire [3-1:0] node89;
	wire [3-1:0] node90;
	wire [3-1:0] node95;
	wire [3-1:0] node96;
	wire [3-1:0] node97;
	wire [3-1:0] node98;
	wire [3-1:0] node99;
	wire [3-1:0] node102;
	wire [3-1:0] node106;
	wire [3-1:0] node108;
	wire [3-1:0] node111;
	wire [3-1:0] node112;
	wire [3-1:0] node114;
	wire [3-1:0] node115;
	wire [3-1:0] node120;
	wire [3-1:0] node121;
	wire [3-1:0] node122;
	wire [3-1:0] node123;
	wire [3-1:0] node124;
	wire [3-1:0] node125;
	wire [3-1:0] node128;
	wire [3-1:0] node131;
	wire [3-1:0] node132;
	wire [3-1:0] node136;
	wire [3-1:0] node139;
	wire [3-1:0] node140;
	wire [3-1:0] node141;
	wire [3-1:0] node142;
	wire [3-1:0] node143;
	wire [3-1:0] node148;
	wire [3-1:0] node150;
	wire [3-1:0] node153;
	wire [3-1:0] node154;
	wire [3-1:0] node157;
	wire [3-1:0] node158;
	wire [3-1:0] node161;
	wire [3-1:0] node162;
	wire [3-1:0] node166;
	wire [3-1:0] node167;
	wire [3-1:0] node169;
	wire [3-1:0] node170;
	wire [3-1:0] node171;
	wire [3-1:0] node175;
	wire [3-1:0] node177;
	wire [3-1:0] node180;
	wire [3-1:0] node181;
	wire [3-1:0] node182;
	wire [3-1:0] node184;
	wire [3-1:0] node185;
	wire [3-1:0] node189;
	wire [3-1:0] node190;
	wire [3-1:0] node192;
	wire [3-1:0] node196;
	wire [3-1:0] node197;
	wire [3-1:0] node201;
	wire [3-1:0] node202;
	wire [3-1:0] node203;
	wire [3-1:0] node204;
	wire [3-1:0] node205;
	wire [3-1:0] node207;
	wire [3-1:0] node209;
	wire [3-1:0] node210;
	wire [3-1:0] node215;
	wire [3-1:0] node216;
	wire [3-1:0] node217;
	wire [3-1:0] node218;
	wire [3-1:0] node220;
	wire [3-1:0] node223;
	wire [3-1:0] node226;
	wire [3-1:0] node228;
	wire [3-1:0] node231;
	wire [3-1:0] node232;
	wire [3-1:0] node235;
	wire [3-1:0] node236;
	wire [3-1:0] node239;
	wire [3-1:0] node242;
	wire [3-1:0] node243;
	wire [3-1:0] node244;
	wire [3-1:0] node246;
	wire [3-1:0] node247;
	wire [3-1:0] node248;
	wire [3-1:0] node252;
	wire [3-1:0] node254;
	wire [3-1:0] node257;
	wire [3-1:0] node259;
	wire [3-1:0] node261;
	wire [3-1:0] node262;
	wire [3-1:0] node265;
	wire [3-1:0] node268;
	wire [3-1:0] node269;
	wire [3-1:0] node271;
	wire [3-1:0] node272;
	wire [3-1:0] node275;
	wire [3-1:0] node276;
	wire [3-1:0] node280;
	wire [3-1:0] node281;
	wire [3-1:0] node283;
	wire [3-1:0] node286;
	wire [3-1:0] node287;
	wire [3-1:0] node290;
	wire [3-1:0] node293;
	wire [3-1:0] node294;
	wire [3-1:0] node295;
	wire [3-1:0] node296;
	wire [3-1:0] node297;
	wire [3-1:0] node298;
	wire [3-1:0] node301;
	wire [3-1:0] node304;
	wire [3-1:0] node305;
	wire [3-1:0] node309;
	wire [3-1:0] node310;
	wire [3-1:0] node311;
	wire [3-1:0] node312;
	wire [3-1:0] node315;
	wire [3-1:0] node318;
	wire [3-1:0] node322;
	wire [3-1:0] node323;
	wire [3-1:0] node325;
	wire [3-1:0] node328;
	wire [3-1:0] node329;
	wire [3-1:0] node333;
	wire [3-1:0] node334;
	wire [3-1:0] node335;
	wire [3-1:0] node336;
	wire [3-1:0] node337;
	wire [3-1:0] node340;
	wire [3-1:0] node341;
	wire [3-1:0] node346;
	wire [3-1:0] node348;
	wire [3-1:0] node351;
	wire [3-1:0] node352;
	wire [3-1:0] node353;
	wire [3-1:0] node355;
	wire [3-1:0] node358;
	wire [3-1:0] node359;
	wire [3-1:0] node361;
	wire [3-1:0] node365;
	wire [3-1:0] node366;
	wire [3-1:0] node367;
	wire [3-1:0] node370;
	wire [3-1:0] node372;
	wire [3-1:0] node375;
	wire [3-1:0] node377;
	wire [3-1:0] node380;
	wire [3-1:0] node381;
	wire [3-1:0] node382;
	wire [3-1:0] node383;
	wire [3-1:0] node384;
	wire [3-1:0] node385;
	wire [3-1:0] node386;
	wire [3-1:0] node387;
	wire [3-1:0] node388;
	wire [3-1:0] node390;
	wire [3-1:0] node394;
	wire [3-1:0] node395;
	wire [3-1:0] node398;
	wire [3-1:0] node401;
	wire [3-1:0] node402;
	wire [3-1:0] node403;
	wire [3-1:0] node406;
	wire [3-1:0] node408;
	wire [3-1:0] node411;
	wire [3-1:0] node412;
	wire [3-1:0] node414;
	wire [3-1:0] node417;
	wire [3-1:0] node420;
	wire [3-1:0] node422;
	wire [3-1:0] node423;
	wire [3-1:0] node426;
	wire [3-1:0] node427;
	wire [3-1:0] node431;
	wire [3-1:0] node433;
	wire [3-1:0] node434;
	wire [3-1:0] node437;
	wire [3-1:0] node438;
	wire [3-1:0] node439;
	wire [3-1:0] node443;
	wire [3-1:0] node445;
	wire [3-1:0] node448;
	wire [3-1:0] node449;
	wire [3-1:0] node450;
	wire [3-1:0] node451;
	wire [3-1:0] node452;
	wire [3-1:0] node453;
	wire [3-1:0] node454;
	wire [3-1:0] node460;
	wire [3-1:0] node461;
	wire [3-1:0] node464;
	wire [3-1:0] node465;
	wire [3-1:0] node469;
	wire [3-1:0] node471;
	wire [3-1:0] node474;
	wire [3-1:0] node475;
	wire [3-1:0] node476;
	wire [3-1:0] node478;
	wire [3-1:0] node479;
	wire [3-1:0] node481;
	wire [3-1:0] node485;
	wire [3-1:0] node486;
	wire [3-1:0] node488;
	wire [3-1:0] node490;
	wire [3-1:0] node494;
	wire [3-1:0] node495;
	wire [3-1:0] node497;
	wire [3-1:0] node500;
	wire [3-1:0] node501;
	wire [3-1:0] node503;
	wire [3-1:0] node504;
	wire [3-1:0] node508;
	wire [3-1:0] node509;
	wire [3-1:0] node513;
	wire [3-1:0] node514;
	wire [3-1:0] node515;
	wire [3-1:0] node516;
	wire [3-1:0] node517;
	wire [3-1:0] node519;
	wire [3-1:0] node521;
	wire [3-1:0] node524;
	wire [3-1:0] node525;
	wire [3-1:0] node528;
	wire [3-1:0] node529;
	wire [3-1:0] node530;
	wire [3-1:0] node535;
	wire [3-1:0] node536;
	wire [3-1:0] node537;
	wire [3-1:0] node539;
	wire [3-1:0] node542;
	wire [3-1:0] node544;
	wire [3-1:0] node545;
	wire [3-1:0] node549;
	wire [3-1:0] node550;
	wire [3-1:0] node551;
	wire [3-1:0] node555;
	wire [3-1:0] node558;
	wire [3-1:0] node559;
	wire [3-1:0] node560;
	wire [3-1:0] node561;
	wire [3-1:0] node562;
	wire [3-1:0] node565;
	wire [3-1:0] node569;
	wire [3-1:0] node571;
	wire [3-1:0] node573;
	wire [3-1:0] node574;
	wire [3-1:0] node578;
	wire [3-1:0] node579;
	wire [3-1:0] node580;
	wire [3-1:0] node582;
	wire [3-1:0] node585;
	wire [3-1:0] node586;
	wire [3-1:0] node589;
	wire [3-1:0] node590;
	wire [3-1:0] node594;
	wire [3-1:0] node595;
	wire [3-1:0] node597;
	wire [3-1:0] node601;
	wire [3-1:0] node602;
	wire [3-1:0] node603;
	wire [3-1:0] node605;
	wire [3-1:0] node608;
	wire [3-1:0] node609;
	wire [3-1:0] node610;
	wire [3-1:0] node612;
	wire [3-1:0] node615;
	wire [3-1:0] node617;
	wire [3-1:0] node620;
	wire [3-1:0] node621;
	wire [3-1:0] node625;
	wire [3-1:0] node626;
	wire [3-1:0] node627;
	wire [3-1:0] node628;
	wire [3-1:0] node629;
	wire [3-1:0] node632;
	wire [3-1:0] node634;
	wire [3-1:0] node637;
	wire [3-1:0] node639;
	wire [3-1:0] node642;
	wire [3-1:0] node644;
	wire [3-1:0] node647;
	wire [3-1:0] node648;
	wire [3-1:0] node650;
	wire [3-1:0] node651;
	wire [3-1:0] node654;
	wire [3-1:0] node657;
	wire [3-1:0] node658;
	wire [3-1:0] node661;
	wire [3-1:0] node662;
	wire [3-1:0] node663;
	wire [3-1:0] node666;
	wire [3-1:0] node669;
	wire [3-1:0] node672;
	wire [3-1:0] node673;
	wire [3-1:0] node674;
	wire [3-1:0] node675;
	wire [3-1:0] node676;
	wire [3-1:0] node677;
	wire [3-1:0] node679;
	wire [3-1:0] node680;
	wire [3-1:0] node681;
	wire [3-1:0] node685;
	wire [3-1:0] node688;
	wire [3-1:0] node689;
	wire [3-1:0] node690;
	wire [3-1:0] node693;
	wire [3-1:0] node697;
	wire [3-1:0] node698;
	wire [3-1:0] node699;
	wire [3-1:0] node701;
	wire [3-1:0] node704;
	wire [3-1:0] node705;
	wire [3-1:0] node706;
	wire [3-1:0] node711;
	wire [3-1:0] node712;
	wire [3-1:0] node715;
	wire [3-1:0] node718;
	wire [3-1:0] node719;
	wire [3-1:0] node720;
	wire [3-1:0] node721;
	wire [3-1:0] node724;
	wire [3-1:0] node727;
	wire [3-1:0] node728;
	wire [3-1:0] node732;
	wire [3-1:0] node733;
	wire [3-1:0] node734;
	wire [3-1:0] node737;
	wire [3-1:0] node738;
	wire [3-1:0] node741;
	wire [3-1:0] node742;
	wire [3-1:0] node746;
	wire [3-1:0] node747;
	wire [3-1:0] node751;
	wire [3-1:0] node752;
	wire [3-1:0] node753;
	wire [3-1:0] node755;
	wire [3-1:0] node756;
	wire [3-1:0] node759;
	wire [3-1:0] node763;
	wire [3-1:0] node764;
	wire [3-1:0] node765;
	wire [3-1:0] node768;
	wire [3-1:0] node770;
	wire [3-1:0] node771;
	wire [3-1:0] node772;
	wire [3-1:0] node777;
	wire [3-1:0] node778;
	wire [3-1:0] node779;
	wire [3-1:0] node781;
	wire [3-1:0] node784;
	wire [3-1:0] node785;
	wire [3-1:0] node789;
	wire [3-1:0] node791;
	wire [3-1:0] node792;
	wire [3-1:0] node795;
	wire [3-1:0] node796;
	wire [3-1:0] node800;
	wire [3-1:0] node801;
	wire [3-1:0] node803;
	wire [3-1:0] node804;
	wire [3-1:0] node805;
	wire [3-1:0] node806;
	wire [3-1:0] node808;
	wire [3-1:0] node810;
	wire [3-1:0] node813;
	wire [3-1:0] node815;
	wire [3-1:0] node817;
	wire [3-1:0] node820;
	wire [3-1:0] node824;
	wire [3-1:0] node825;
	wire [3-1:0] node826;
	wire [3-1:0] node828;
	wire [3-1:0] node829;
	wire [3-1:0] node833;
	wire [3-1:0] node834;
	wire [3-1:0] node835;
	wire [3-1:0] node836;
	wire [3-1:0] node840;
	wire [3-1:0] node843;
	wire [3-1:0] node844;
	wire [3-1:0] node845;
	wire [3-1:0] node846;
	wire [3-1:0] node852;
	wire [3-1:0] node853;
	wire [3-1:0] node854;
	wire [3-1:0] node855;
	wire [3-1:0] node856;
	wire [3-1:0] node857;
	wire [3-1:0] node861;
	wire [3-1:0] node864;
	wire [3-1:0] node866;
	wire [3-1:0] node867;
	wire [3-1:0] node871;
	wire [3-1:0] node872;
	wire [3-1:0] node873;
	wire [3-1:0] node877;
	wire [3-1:0] node880;
	wire [3-1:0] node881;
	wire [3-1:0] node882;
	wire [3-1:0] node883;
	wire [3-1:0] node887;
	wire [3-1:0] node889;
	wire [3-1:0] node892;
	wire [3-1:0] node894;
	wire [3-1:0] node895;
	wire [3-1:0] node898;
	wire [3-1:0] node899;
	wire [3-1:0] node902;

	assign outp = (inp[0]) ? node380 : node1;
		assign node1 = (inp[6]) ? node43 : node2;
			assign node2 = (inp[3]) ? node16 : node3;
				assign node3 = (inp[7]) ? node5 : 3'b011;
					assign node5 = (inp[4]) ? node7 : 3'b011;
						assign node7 = (inp[8]) ? node9 : 3'b111;
							assign node9 = (inp[5]) ? node11 : 3'b111;
								assign node11 = (inp[1]) ? node13 : 3'b111;
									assign node13 = (inp[2]) ? 3'b011 : 3'b111;
				assign node16 = (inp[9]) ? 3'b111 : node17;
					assign node17 = (inp[7]) ? node19 : 3'b111;
						assign node19 = (inp[1]) ? node27 : node20;
							assign node20 = (inp[4]) ? 3'b111 : node21;
								assign node21 = (inp[8]) ? node23 : 3'b111;
									assign node23 = (inp[5]) ? 3'b111 : 3'b011;
							assign node27 = (inp[4]) ? node33 : node28;
								assign node28 = (inp[11]) ? 3'b001 : node29;
									assign node29 = (inp[10]) ? 3'b101 : 3'b001;
								assign node33 = (inp[2]) ? node37 : node34;
									assign node34 = (inp[8]) ? 3'b011 : 3'b111;
									assign node37 = (inp[10]) ? 3'b011 : node38;
										assign node38 = (inp[8]) ? 3'b101 : 3'b011;
			assign node43 = (inp[7]) ? node201 : node44;
				assign node44 = (inp[3]) ? node120 : node45;
					assign node45 = (inp[4]) ? node81 : node46;
						assign node46 = (inp[10]) ? node66 : node47;
							assign node47 = (inp[8]) ? node57 : node48;
								assign node48 = (inp[11]) ? 3'b001 : node49;
									assign node49 = (inp[9]) ? 3'b001 : node50;
										assign node50 = (inp[5]) ? node52 : 3'b101;
											assign node52 = (inp[2]) ? 3'b101 : 3'b001;
								assign node57 = (inp[2]) ? node63 : node58;
									assign node58 = (inp[9]) ? 3'b101 : node59;
										assign node59 = (inp[11]) ? 3'b101 : 3'b001;
									assign node63 = (inp[1]) ? 3'b010 : 3'b101;
							assign node66 = (inp[1]) ? node76 : node67;
								assign node67 = (inp[5]) ? 3'b001 : node68;
									assign node68 = (inp[11]) ? node70 : 3'b101;
										assign node70 = (inp[8]) ? node72 : 3'b001;
											assign node72 = (inp[2]) ? 3'b101 : 3'b001;
								assign node76 = (inp[5]) ? node78 : 3'b101;
									assign node78 = (inp[11]) ? 3'b110 : 3'b101;
						assign node81 = (inp[10]) ? node95 : node82;
							assign node82 = (inp[1]) ? node88 : node83;
								assign node83 = (inp[9]) ? 3'b011 : node84;
									assign node84 = (inp[11]) ? 3'b101 : 3'b001;
								assign node88 = (inp[5]) ? 3'b101 : node89;
									assign node89 = (inp[9]) ? 3'b111 : node90;
										assign node90 = (inp[8]) ? 3'b011 : 3'b111;
							assign node95 = (inp[8]) ? node111 : node96;
								assign node96 = (inp[11]) ? node106 : node97;
									assign node97 = (inp[9]) ? 3'b101 : node98;
										assign node98 = (inp[2]) ? node102 : node99;
											assign node99 = (inp[1]) ? 3'b001 : 3'b101;
											assign node102 = (inp[5]) ? 3'b011 : 3'b001;
									assign node106 = (inp[5]) ? node108 : 3'b101;
										assign node108 = (inp[2]) ? 3'b011 : 3'b111;
								assign node111 = (inp[11]) ? 3'b001 : node112;
									assign node112 = (inp[5]) ? node114 : 3'b011;
										assign node114 = (inp[2]) ? 3'b101 : node115;
											assign node115 = (inp[9]) ? 3'b001 : 3'b011;
					assign node120 = (inp[9]) ? node166 : node121;
						assign node121 = (inp[1]) ? node139 : node122;
							assign node122 = (inp[5]) ? node136 : node123;
								assign node123 = (inp[11]) ? node131 : node124;
									assign node124 = (inp[10]) ? node128 : node125;
										assign node125 = (inp[8]) ? 3'b111 : 3'b101;
										assign node128 = (inp[4]) ? 3'b111 : 3'b011;
									assign node131 = (inp[10]) ? 3'b101 : node132;
										assign node132 = (inp[2]) ? 3'b001 : 3'b101;
								assign node136 = (inp[4]) ? 3'b111 : 3'b011;
							assign node139 = (inp[11]) ? node153 : node140;
								assign node140 = (inp[2]) ? node148 : node141;
									assign node141 = (inp[5]) ? 3'b101 : node142;
										assign node142 = (inp[4]) ? 3'b101 : node143;
											assign node143 = (inp[10]) ? 3'b101 : 3'b001;
									assign node148 = (inp[10]) ? node150 : 3'b001;
										assign node150 = (inp[4]) ? 3'b010 : 3'b001;
								assign node153 = (inp[8]) ? node157 : node154;
									assign node154 = (inp[5]) ? 3'b010 : 3'b001;
									assign node157 = (inp[10]) ? node161 : node158;
										assign node158 = (inp[4]) ? 3'b110 : 3'b010;
										assign node161 = (inp[5]) ? 3'b001 : node162;
											assign node162 = (inp[4]) ? 3'b110 : 3'b001;
						assign node166 = (inp[1]) ? node180 : node167;
							assign node167 = (inp[2]) ? node169 : 3'b111;
								assign node169 = (inp[5]) ? node175 : node170;
									assign node170 = (inp[8]) ? 3'b101 : node171;
										assign node171 = (inp[11]) ? 3'b111 : 3'b101;
									assign node175 = (inp[4]) ? node177 : 3'b111;
										assign node177 = (inp[10]) ? 3'b111 : 3'b011;
							assign node180 = (inp[10]) ? node196 : node181;
								assign node181 = (inp[4]) ? node189 : node182;
									assign node182 = (inp[2]) ? node184 : 3'b111;
										assign node184 = (inp[8]) ? 3'b101 : node185;
											assign node185 = (inp[11]) ? 3'b001 : 3'b011;
									assign node189 = (inp[8]) ? 3'b011 : node190;
										assign node190 = (inp[11]) ? node192 : 3'b111;
											assign node192 = (inp[2]) ? 3'b011 : 3'b111;
								assign node196 = (inp[5]) ? 3'b111 : node197;
									assign node197 = (inp[2]) ? 3'b111 : 3'b011;
				assign node201 = (inp[3]) ? node293 : node202;
					assign node202 = (inp[4]) ? node242 : node203;
						assign node203 = (inp[9]) ? node215 : node204;
							assign node204 = (inp[8]) ? 3'b000 : node205;
								assign node205 = (inp[2]) ? node207 : 3'b100;
									assign node207 = (inp[11]) ? node209 : 3'b000;
										assign node209 = (inp[10]) ? 3'b100 : node210;
											assign node210 = (inp[5]) ? 3'b000 : 3'b100;
							assign node215 = (inp[10]) ? node231 : node216;
								assign node216 = (inp[5]) ? node226 : node217;
									assign node217 = (inp[8]) ? node223 : node218;
										assign node218 = (inp[2]) ? node220 : 3'b110;
											assign node220 = (inp[11]) ? 3'b100 : 3'b000;
										assign node223 = (inp[2]) ? 3'b010 : 3'b000;
									assign node226 = (inp[11]) ? node228 : 3'b011;
										assign node228 = (inp[1]) ? 3'b001 : 3'b000;
								assign node231 = (inp[1]) ? node235 : node232;
									assign node232 = (inp[2]) ? 3'b100 : 3'b101;
									assign node235 = (inp[8]) ? node239 : node236;
										assign node236 = (inp[2]) ? 3'b010 : 3'b110;
										assign node239 = (inp[2]) ? 3'b100 : 3'b110;
						assign node242 = (inp[1]) ? node268 : node243;
							assign node243 = (inp[9]) ? node257 : node244;
								assign node244 = (inp[11]) ? node246 : 3'b110;
									assign node246 = (inp[10]) ? node252 : node247;
										assign node247 = (inp[2]) ? 3'b010 : node248;
											assign node248 = (inp[5]) ? 3'b011 : 3'b111;
										assign node252 = (inp[5]) ? node254 : 3'b111;
											assign node254 = (inp[8]) ? 3'b111 : 3'b001;
								assign node257 = (inp[10]) ? node259 : 3'b101;
									assign node259 = (inp[2]) ? node261 : 3'b011;
										assign node261 = (inp[5]) ? node265 : node262;
											assign node262 = (inp[8]) ? 3'b001 : 3'b101;
											assign node265 = (inp[8]) ? 3'b101 : 3'b011;
							assign node268 = (inp[8]) ? node280 : node269;
								assign node269 = (inp[9]) ? node271 : 3'b010;
									assign node271 = (inp[2]) ? node275 : node272;
										assign node272 = (inp[11]) ? 3'b001 : 3'b101;
										assign node275 = (inp[5]) ? 3'b001 : node276;
											assign node276 = (inp[10]) ? 3'b110 : 3'b010;
								assign node280 = (inp[5]) ? node286 : node281;
									assign node281 = (inp[9]) ? node283 : 3'b100;
										assign node283 = (inp[10]) ? 3'b010 : 3'b100;
									assign node286 = (inp[10]) ? node290 : node287;
										assign node287 = (inp[9]) ? 3'b010 : 3'b000;
										assign node290 = (inp[11]) ? 3'b010 : 3'b110;
					assign node293 = (inp[4]) ? node333 : node294;
						assign node294 = (inp[1]) ? node322 : node295;
							assign node295 = (inp[8]) ? node309 : node296;
								assign node296 = (inp[10]) ? node304 : node297;
									assign node297 = (inp[2]) ? node301 : node298;
										assign node298 = (inp[9]) ? 3'b111 : 3'b101;
										assign node301 = (inp[9]) ? 3'b101 : 3'b110;
									assign node304 = (inp[9]) ? 3'b011 : node305;
										assign node305 = (inp[2]) ? 3'b010 : 3'b011;
								assign node309 = (inp[11]) ? 3'b011 : node310;
									assign node310 = (inp[9]) ? node318 : node311;
										assign node311 = (inp[10]) ? node315 : node312;
											assign node312 = (inp[2]) ? 3'b010 : 3'b001;
											assign node315 = (inp[5]) ? 3'b001 : 3'b101;
										assign node318 = (inp[10]) ? 3'b011 : 3'b001;
							assign node322 = (inp[2]) ? node328 : node323;
								assign node323 = (inp[11]) ? node325 : 3'b110;
									assign node325 = (inp[5]) ? 3'b101 : 3'b001;
								assign node328 = (inp[5]) ? 3'b010 : node329;
									assign node329 = (inp[8]) ? 3'b000 : 3'b010;
						assign node333 = (inp[1]) ? node351 : node334;
							assign node334 = (inp[9]) ? node346 : node335;
								assign node335 = (inp[2]) ? 3'b001 : node336;
									assign node336 = (inp[11]) ? node340 : node337;
										assign node337 = (inp[5]) ? 3'b011 : 3'b101;
										assign node340 = (inp[8]) ? 3'b111 : node341;
											assign node341 = (inp[5]) ? 3'b101 : 3'b111;
								assign node346 = (inp[2]) ? node348 : 3'b111;
									assign node348 = (inp[10]) ? 3'b111 : 3'b011;
							assign node351 = (inp[9]) ? node365 : node352;
								assign node352 = (inp[2]) ? node358 : node353;
									assign node353 = (inp[11]) ? node355 : 3'b001;
										assign node355 = (inp[8]) ? 3'b001 : 3'b101;
									assign node358 = (inp[5]) ? 3'b110 : node359;
										assign node359 = (inp[8]) ? node361 : 3'b001;
											assign node361 = (inp[10]) ? 3'b110 : 3'b010;
								assign node365 = (inp[10]) ? node375 : node366;
									assign node366 = (inp[2]) ? node370 : node367;
										assign node367 = (inp[11]) ? 3'b111 : 3'b101;
										assign node370 = (inp[5]) ? node372 : 3'b001;
											assign node372 = (inp[11]) ? 3'b101 : 3'b001;
									assign node375 = (inp[2]) ? node377 : 3'b011;
										assign node377 = (inp[8]) ? 3'b101 : 3'b011;
		assign node380 = (inp[6]) ? node672 : node381;
			assign node381 = (inp[3]) ? node513 : node382;
				assign node382 = (inp[4]) ? node448 : node383;
					assign node383 = (inp[9]) ? node431 : node384;
						assign node384 = (inp[10]) ? node420 : node385;
							assign node385 = (inp[8]) ? node401 : node386;
								assign node386 = (inp[1]) ? node394 : node387;
									assign node387 = (inp[5]) ? 3'b100 : node388;
										assign node388 = (inp[11]) ? node390 : 3'b100;
											assign node390 = (inp[2]) ? 3'b100 : 3'b000;
									assign node394 = (inp[2]) ? node398 : node395;
										assign node395 = (inp[7]) ? 3'b110 : 3'b100;
										assign node398 = (inp[7]) ? 3'b010 : 3'b000;
								assign node401 = (inp[2]) ? node411 : node402;
									assign node402 = (inp[5]) ? node406 : node403;
										assign node403 = (inp[11]) ? 3'b010 : 3'b000;
										assign node406 = (inp[11]) ? node408 : 3'b110;
											assign node408 = (inp[1]) ? 3'b100 : 3'b110;
									assign node411 = (inp[5]) ? node417 : node412;
										assign node412 = (inp[7]) ? node414 : 3'b100;
											assign node414 = (inp[1]) ? 3'b100 : 3'b110;
										assign node417 = (inp[7]) ? 3'b000 : 3'b010;
							assign node420 = (inp[5]) ? node422 : 3'b000;
								assign node422 = (inp[11]) ? node426 : node423;
									assign node423 = (inp[1]) ? 3'b010 : 3'b100;
									assign node426 = (inp[1]) ? 3'b110 : node427;
										assign node427 = (inp[8]) ? 3'b010 : 3'b110;
						assign node431 = (inp[1]) ? node433 : 3'b110;
							assign node433 = (inp[5]) ? node437 : node434;
								assign node434 = (inp[8]) ? 3'b100 : 3'b010;
								assign node437 = (inp[2]) ? node443 : node438;
									assign node438 = (inp[10]) ? 3'b110 : node439;
										assign node439 = (inp[7]) ? 3'b100 : 3'b110;
									assign node443 = (inp[10]) ? node445 : 3'b110;
										assign node445 = (inp[11]) ? 3'b010 : 3'b000;
					assign node448 = (inp[9]) ? node474 : node449;
						assign node449 = (inp[2]) ? node469 : node450;
							assign node450 = (inp[7]) ? node460 : node451;
								assign node451 = (inp[8]) ? 3'b001 : node452;
									assign node452 = (inp[10]) ? 3'b110 : node453;
										assign node453 = (inp[1]) ? 3'b001 : node454;
											assign node454 = (inp[11]) ? 3'b110 : 3'b000;
								assign node460 = (inp[1]) ? node464 : node461;
									assign node461 = (inp[10]) ? 3'b101 : 3'b001;
									assign node464 = (inp[8]) ? 3'b000 : node465;
										assign node465 = (inp[5]) ? 3'b001 : 3'b000;
							assign node469 = (inp[7]) ? node471 : 3'b001;
								assign node471 = (inp[1]) ? 3'b000 : 3'b001;
						assign node474 = (inp[1]) ? node494 : node475;
							assign node475 = (inp[7]) ? node485 : node476;
								assign node476 = (inp[11]) ? node478 : 3'b110;
									assign node478 = (inp[8]) ? 3'b110 : node479;
										assign node479 = (inp[5]) ? node481 : 3'b001;
											assign node481 = (inp[2]) ? 3'b110 : 3'b001;
								assign node485 = (inp[10]) ? 3'b101 : node486;
									assign node486 = (inp[2]) ? node488 : 3'b001;
										assign node488 = (inp[8]) ? node490 : 3'b001;
											assign node490 = (inp[5]) ? 3'b101 : 3'b001;
							assign node494 = (inp[2]) ? node500 : node495;
								assign node495 = (inp[5]) ? node497 : 3'b110;
									assign node497 = (inp[8]) ? 3'b110 : 3'b001;
								assign node500 = (inp[7]) ? node508 : node501;
									assign node501 = (inp[10]) ? node503 : 3'b110;
										assign node503 = (inp[8]) ? 3'b001 : node504;
											assign node504 = (inp[11]) ? 3'b001 : 3'b110;
									assign node508 = (inp[5]) ? 3'b010 : node509;
										assign node509 = (inp[8]) ? 3'b100 : 3'b010;
				assign node513 = (inp[9]) ? node601 : node514;
					assign node514 = (inp[1]) ? node558 : node515;
						assign node515 = (inp[7]) ? node535 : node516;
							assign node516 = (inp[4]) ? node524 : node517;
								assign node517 = (inp[2]) ? node519 : 3'b111;
									assign node519 = (inp[11]) ? node521 : 3'b111;
										assign node521 = (inp[8]) ? 3'b011 : 3'b111;
								assign node524 = (inp[2]) ? node528 : node525;
									assign node525 = (inp[5]) ? 3'b111 : 3'b011;
									assign node528 = (inp[11]) ? 3'b011 : node529;
										assign node529 = (inp[8]) ? 3'b101 : node530;
											assign node530 = (inp[5]) ? 3'b011 : 3'b101;
							assign node535 = (inp[4]) ? node549 : node536;
								assign node536 = (inp[11]) ? node542 : node537;
									assign node537 = (inp[2]) ? node539 : 3'b110;
										assign node539 = (inp[10]) ? 3'b110 : 3'b010;
									assign node542 = (inp[8]) ? node544 : 3'b000;
										assign node544 = (inp[5]) ? 3'b000 : node545;
											assign node545 = (inp[10]) ? 3'b110 : 3'b010;
								assign node549 = (inp[8]) ? node555 : node550;
									assign node550 = (inp[2]) ? 3'b011 : node551;
										assign node551 = (inp[10]) ? 3'b111 : 3'b011;
									assign node555 = (inp[10]) ? 3'b001 : 3'b110;
						assign node558 = (inp[5]) ? node578 : node559;
							assign node559 = (inp[8]) ? node569 : node560;
								assign node560 = (inp[4]) ? 3'b001 : node561;
									assign node561 = (inp[10]) ? node565 : node562;
										assign node562 = (inp[7]) ? 3'b100 : 3'b110;
										assign node565 = (inp[2]) ? 3'b110 : 3'b010;
								assign node569 = (inp[4]) ? node571 : 3'b000;
									assign node571 = (inp[2]) ? node573 : 3'b010;
										assign node573 = (inp[11]) ? 3'b000 : node574;
											assign node574 = (inp[7]) ? 3'b000 : 3'b010;
							assign node578 = (inp[11]) ? node594 : node579;
								assign node579 = (inp[7]) ? node585 : node580;
									assign node580 = (inp[2]) ? node582 : 3'b101;
										assign node582 = (inp[4]) ? 3'b110 : 3'b010;
									assign node585 = (inp[4]) ? node589 : node586;
										assign node586 = (inp[2]) ? 3'b100 : 3'b110;
										assign node589 = (inp[10]) ? 3'b000 : node590;
											assign node590 = (inp[2]) ? 3'b010 : 3'b110;
								assign node594 = (inp[4]) ? 3'b110 : node595;
									assign node595 = (inp[10]) ? node597 : 3'b011;
										assign node597 = (inp[8]) ? 3'b110 : 3'b010;
					assign node601 = (inp[7]) ? node625 : node602;
						assign node602 = (inp[2]) ? node608 : node603;
							assign node603 = (inp[1]) ? node605 : 3'b111;
								assign node605 = (inp[4]) ? 3'b111 : 3'b011;
							assign node608 = (inp[4]) ? node620 : node609;
								assign node609 = (inp[1]) ? node615 : node610;
									assign node610 = (inp[8]) ? node612 : 3'b111;
										assign node612 = (inp[5]) ? 3'b111 : 3'b011;
									assign node615 = (inp[11]) ? node617 : 3'b101;
										assign node617 = (inp[5]) ? 3'b001 : 3'b101;
								assign node620 = (inp[5]) ? 3'b111 : node621;
									assign node621 = (inp[1]) ? 3'b011 : 3'b111;
						assign node625 = (inp[1]) ? node647 : node626;
							assign node626 = (inp[4]) ? node642 : node627;
								assign node627 = (inp[10]) ? node637 : node628;
									assign node628 = (inp[8]) ? node632 : node629;
										assign node629 = (inp[2]) ? 3'b101 : 3'b011;
										assign node632 = (inp[2]) ? node634 : 3'b101;
											assign node634 = (inp[5]) ? 3'b101 : 3'b001;
									assign node637 = (inp[5]) ? node639 : 3'b011;
										assign node639 = (inp[2]) ? 3'b011 : 3'b111;
								assign node642 = (inp[2]) ? node644 : 3'b111;
									assign node644 = (inp[10]) ? 3'b111 : 3'b011;
							assign node647 = (inp[8]) ? node657 : node648;
								assign node648 = (inp[10]) ? node650 : 3'b001;
									assign node650 = (inp[5]) ? node654 : node651;
										assign node651 = (inp[11]) ? 3'b101 : 3'b001;
										assign node654 = (inp[11]) ? 3'b001 : 3'b101;
								assign node657 = (inp[10]) ? node661 : node658;
									assign node658 = (inp[11]) ? 3'b110 : 3'b010;
									assign node661 = (inp[11]) ? node669 : node662;
										assign node662 = (inp[4]) ? node666 : node663;
											assign node663 = (inp[5]) ? 3'b110 : 3'b100;
											assign node666 = (inp[2]) ? 3'b001 : 3'b111;
										assign node669 = (inp[4]) ? 3'b101 : 3'b001;
			assign node672 = (inp[7]) ? node800 : node673;
				assign node673 = (inp[1]) ? node751 : node674;
					assign node674 = (inp[3]) ? node718 : node675;
						assign node675 = (inp[9]) ? node697 : node676;
							assign node676 = (inp[4]) ? node688 : node677;
								assign node677 = (inp[2]) ? node679 : 3'b110;
									assign node679 = (inp[10]) ? node685 : node680;
										assign node680 = (inp[8]) ? 3'b000 : node681;
											assign node681 = (inp[5]) ? 3'b100 : 3'b000;
										assign node685 = (inp[8]) ? 3'b100 : 3'b010;
								assign node688 = (inp[2]) ? 3'b110 : node689;
									assign node689 = (inp[5]) ? node693 : node690;
										assign node690 = (inp[8]) ? 3'b110 : 3'b100;
										assign node693 = (inp[10]) ? 3'b101 : 3'b100;
							assign node697 = (inp[8]) ? node711 : node698;
								assign node698 = (inp[11]) ? node704 : node699;
									assign node699 = (inp[2]) ? node701 : 3'b000;
										assign node701 = (inp[4]) ? 3'b110 : 3'b100;
									assign node704 = (inp[4]) ? 3'b110 : node705;
										assign node705 = (inp[2]) ? 3'b000 : node706;
											assign node706 = (inp[10]) ? 3'b110 : 3'b010;
								assign node711 = (inp[5]) ? node715 : node712;
									assign node712 = (inp[2]) ? 3'b010 : 3'b110;
									assign node715 = (inp[2]) ? 3'b110 : 3'b010;
						assign node718 = (inp[9]) ? node732 : node719;
							assign node719 = (inp[2]) ? node727 : node720;
								assign node720 = (inp[5]) ? node724 : node721;
									assign node721 = (inp[4]) ? 3'b010 : 3'b100;
									assign node724 = (inp[4]) ? 3'b001 : 3'b010;
								assign node727 = (inp[8]) ? 3'b100 : node728;
									assign node728 = (inp[4]) ? 3'b110 : 3'b100;
							assign node732 = (inp[4]) ? node746 : node733;
								assign node733 = (inp[10]) ? node737 : node734;
									assign node734 = (inp[5]) ? 3'b100 : 3'b000;
									assign node737 = (inp[11]) ? node741 : node738;
										assign node738 = (inp[2]) ? 3'b100 : 3'b101;
										assign node741 = (inp[8]) ? 3'b001 : node742;
											assign node742 = (inp[5]) ? 3'b101 : 3'b001;
								assign node746 = (inp[2]) ? 3'b101 : node747;
									assign node747 = (inp[10]) ? 3'b111 : 3'b101;
					assign node751 = (inp[3]) ? node763 : node752;
						assign node752 = (inp[8]) ? 3'b000 : node753;
							assign node753 = (inp[5]) ? node755 : 3'b000;
								assign node755 = (inp[2]) ? node759 : node756;
									assign node756 = (inp[4]) ? 3'b010 : 3'b100;
									assign node759 = (inp[10]) ? 3'b100 : 3'b000;
						assign node763 = (inp[9]) ? node777 : node764;
							assign node764 = (inp[8]) ? node768 : node765;
								assign node765 = (inp[4]) ? 3'b010 : 3'b000;
								assign node768 = (inp[4]) ? node770 : 3'b000;
									assign node770 = (inp[10]) ? 3'b100 : node771;
										assign node771 = (inp[2]) ? 3'b000 : node772;
											assign node772 = (inp[11]) ? 3'b000 : 3'b100;
							assign node777 = (inp[2]) ? node789 : node778;
								assign node778 = (inp[4]) ? node784 : node779;
									assign node779 = (inp[11]) ? node781 : 3'b110;
										assign node781 = (inp[10]) ? 3'b110 : 3'b010;
									assign node784 = (inp[5]) ? 3'b101 : node785;
										assign node785 = (inp[10]) ? 3'b001 : 3'b101;
								assign node789 = (inp[11]) ? node791 : 3'b010;
									assign node791 = (inp[5]) ? node795 : node792;
										assign node792 = (inp[8]) ? 3'b100 : 3'b110;
										assign node795 = (inp[10]) ? 3'b110 : node796;
											assign node796 = (inp[8]) ? 3'b010 : 3'b110;
				assign node800 = (inp[3]) ? node824 : node801;
					assign node801 = (inp[9]) ? node803 : 3'b000;
						assign node803 = (inp[1]) ? 3'b000 : node804;
							assign node804 = (inp[5]) ? node820 : node805;
								assign node805 = (inp[4]) ? node813 : node806;
									assign node806 = (inp[10]) ? node808 : 3'b000;
										assign node808 = (inp[11]) ? node810 : 3'b000;
											assign node810 = (inp[2]) ? 3'b000 : 3'b100;
									assign node813 = (inp[8]) ? node815 : 3'b100;
										assign node815 = (inp[10]) ? node817 : 3'b000;
											assign node817 = (inp[2]) ? 3'b000 : 3'b100;
								assign node820 = (inp[2]) ? 3'b000 : 3'b010;
					assign node824 = (inp[9]) ? node852 : node825;
						assign node825 = (inp[4]) ? node833 : node826;
							assign node826 = (inp[5]) ? node828 : 3'b000;
								assign node828 = (inp[1]) ? 3'b000 : node829;
									assign node829 = (inp[10]) ? 3'b100 : 3'b000;
							assign node833 = (inp[8]) ? node843 : node834;
								assign node834 = (inp[2]) ? node840 : node835;
									assign node835 = (inp[10]) ? 3'b100 : node836;
										assign node836 = (inp[11]) ? 3'b110 : 3'b100;
									assign node840 = (inp[10]) ? 3'b100 : 3'b000;
								assign node843 = (inp[1]) ? 3'b000 : node844;
									assign node844 = (inp[5]) ? 3'b100 : node845;
										assign node845 = (inp[11]) ? 3'b100 : node846;
											assign node846 = (inp[10]) ? 3'b010 : 3'b000;
						assign node852 = (inp[8]) ? node880 : node853;
							assign node853 = (inp[11]) ? node871 : node854;
								assign node854 = (inp[5]) ? node864 : node855;
									assign node855 = (inp[2]) ? node861 : node856;
										assign node856 = (inp[1]) ? 3'b010 : node857;
											assign node857 = (inp[10]) ? 3'b001 : 3'b011;
										assign node861 = (inp[4]) ? 3'b110 : 3'b010;
									assign node864 = (inp[4]) ? node866 : 3'b101;
										assign node866 = (inp[2]) ? 3'b110 : node867;
											assign node867 = (inp[1]) ? 3'b110 : 3'b101;
								assign node871 = (inp[1]) ? node877 : node872;
									assign node872 = (inp[10]) ? 3'b001 : node873;
										assign node873 = (inp[4]) ? 3'b001 : 3'b000;
									assign node877 = (inp[5]) ? 3'b100 : 3'b000;
							assign node880 = (inp[4]) ? node892 : node881;
								assign node881 = (inp[1]) ? node887 : node882;
									assign node882 = (inp[2]) ? 3'b100 : node883;
										assign node883 = (inp[5]) ? 3'b110 : 3'b010;
									assign node887 = (inp[11]) ? node889 : 3'b000;
										assign node889 = (inp[5]) ? 3'b100 : 3'b000;
								assign node892 = (inp[1]) ? node894 : 3'b010;
									assign node894 = (inp[10]) ? node898 : node895;
										assign node895 = (inp[2]) ? 3'b000 : 3'b100;
										assign node898 = (inp[11]) ? node902 : node899;
											assign node899 = (inp[2]) ? 3'b000 : 3'b010;
											assign node902 = (inp[2]) ? 3'b010 : 3'b010;

endmodule