module dtc_split75_bm30 (
	input  wire [14-1:0] inp,
	output wire [8-1:0] outp
);

	wire [8-1:0] node1;
	wire [8-1:0] node2;
	wire [8-1:0] node3;
	wire [8-1:0] node4;
	wire [8-1:0] node5;
	wire [8-1:0] node6;
	wire [8-1:0] node7;
	wire [8-1:0] node9;
	wire [8-1:0] node11;
	wire [8-1:0] node14;
	wire [8-1:0] node15;
	wire [8-1:0] node18;
	wire [8-1:0] node19;
	wire [8-1:0] node21;
	wire [8-1:0] node24;
	wire [8-1:0] node25;
	wire [8-1:0] node29;
	wire [8-1:0] node30;
	wire [8-1:0] node31;
	wire [8-1:0] node33;
	wire [8-1:0] node36;
	wire [8-1:0] node38;
	wire [8-1:0] node39;
	wire [8-1:0] node42;
	wire [8-1:0] node45;
	wire [8-1:0] node46;
	wire [8-1:0] node49;
	wire [8-1:0] node50;
	wire [8-1:0] node51;
	wire [8-1:0] node52;
	wire [8-1:0] node56;
	wire [8-1:0] node57;
	wire [8-1:0] node61;
	wire [8-1:0] node62;
	wire [8-1:0] node64;
	wire [8-1:0] node67;
	wire [8-1:0] node68;
	wire [8-1:0] node72;
	wire [8-1:0] node73;
	wire [8-1:0] node74;
	wire [8-1:0] node75;
	wire [8-1:0] node77;
	wire [8-1:0] node80;
	wire [8-1:0] node81;
	wire [8-1:0] node83;
	wire [8-1:0] node86;
	wire [8-1:0] node88;
	wire [8-1:0] node91;
	wire [8-1:0] node92;
	wire [8-1:0] node93;
	wire [8-1:0] node95;
	wire [8-1:0] node98;
	wire [8-1:0] node99;
	wire [8-1:0] node101;
	wire [8-1:0] node104;
	wire [8-1:0] node106;
	wire [8-1:0] node109;
	wire [8-1:0] node110;
	wire [8-1:0] node112;
	wire [8-1:0] node115;
	wire [8-1:0] node116;
	wire [8-1:0] node118;
	wire [8-1:0] node121;
	wire [8-1:0] node123;
	wire [8-1:0] node127;
	wire [8-1:0] node128;
	wire [8-1:0] node129;
	wire [8-1:0] node130;
	wire [8-1:0] node133;
	wire [8-1:0] node134;
	wire [8-1:0] node135;
	wire [8-1:0] node137;
	wire [8-1:0] node140;
	wire [8-1:0] node142;
	wire [8-1:0] node145;
	wire [8-1:0] node146;
	wire [8-1:0] node147;
	wire [8-1:0] node151;
	wire [8-1:0] node152;
	wire [8-1:0] node156;
	wire [8-1:0] node157;
	wire [8-1:0] node158;
	wire [8-1:0] node159;
	wire [8-1:0] node161;
	wire [8-1:0] node164;
	wire [8-1:0] node165;
	wire [8-1:0] node169;
	wire [8-1:0] node170;
	wire [8-1:0] node172;
	wire [8-1:0] node173;
	wire [8-1:0] node176;
	wire [8-1:0] node179;
	wire [8-1:0] node180;
	wire [8-1:0] node181;
	wire [8-1:0] node184;
	wire [8-1:0] node188;
	wire [8-1:0] node189;
	wire [8-1:0] node190;
	wire [8-1:0] node192;
	wire [8-1:0] node195;
	wire [8-1:0] node197;
	wire [8-1:0] node198;
	wire [8-1:0] node201;
	wire [8-1:0] node204;
	wire [8-1:0] node205;
	wire [8-1:0] node207;
	wire [8-1:0] node210;
	wire [8-1:0] node211;
	wire [8-1:0] node212;
	wire [8-1:0] node215;
	wire [8-1:0] node219;
	wire [8-1:0] node220;
	wire [8-1:0] node221;
	wire [8-1:0] node222;
	wire [8-1:0] node223;
	wire [8-1:0] node225;
	wire [8-1:0] node228;
	wire [8-1:0] node230;
	wire [8-1:0] node231;
	wire [8-1:0] node234;
	wire [8-1:0] node237;
	wire [8-1:0] node238;
	wire [8-1:0] node239;
	wire [8-1:0] node243;
	wire [8-1:0] node244;
	wire [8-1:0] node245;
	wire [8-1:0] node248;
	wire [8-1:0] node252;
	wire [8-1:0] node253;
	wire [8-1:0] node254;
	wire [8-1:0] node256;
	wire [8-1:0] node257;
	wire [8-1:0] node260;
	wire [8-1:0] node263;
	wire [8-1:0] node264;
	wire [8-1:0] node265;
	wire [8-1:0] node268;
	wire [8-1:0] node272;
	wire [8-1:0] node273;
	wire [8-1:0] node275;
	wire [8-1:0] node276;
	wire [8-1:0] node277;
	wire [8-1:0] node280;
	wire [8-1:0] node283;
	wire [8-1:0] node284;
	wire [8-1:0] node287;
	wire [8-1:0] node290;
	wire [8-1:0] node291;
	wire [8-1:0] node292;
	wire [8-1:0] node293;
	wire [8-1:0] node296;
	wire [8-1:0] node299;
	wire [8-1:0] node300;
	wire [8-1:0] node303;
	wire [8-1:0] node307;
	wire [8-1:0] node308;
	wire [8-1:0] node309;
	wire [8-1:0] node310;
	wire [8-1:0] node313;
	wire [8-1:0] node314;
	wire [8-1:0] node315;
	wire [8-1:0] node318;
	wire [8-1:0] node321;
	wire [8-1:0] node323;
	wire [8-1:0] node326;
	wire [8-1:0] node327;
	wire [8-1:0] node328;
	wire [8-1:0] node332;
	wire [8-1:0] node333;
	wire [8-1:0] node334;
	wire [8-1:0] node337;
	wire [8-1:0] node341;
	wire [8-1:0] node342;
	wire [8-1:0] node343;
	wire [8-1:0] node346;
	wire [8-1:0] node347;
	wire [8-1:0] node348;
	wire [8-1:0] node350;
	wire [8-1:0] node353;
	wire [8-1:0] node355;
	wire [8-1:0] node358;
	wire [8-1:0] node359;
	wire [8-1:0] node362;
	wire [8-1:0] node363;
	wire [8-1:0] node366;
	wire [8-1:0] node369;
	wire [8-1:0] node370;
	wire [8-1:0] node371;
	wire [8-1:0] node372;
	wire [8-1:0] node375;
	wire [8-1:0] node376;
	wire [8-1:0] node379;
	wire [8-1:0] node382;
	wire [8-1:0] node383;
	wire [8-1:0] node384;
	wire [8-1:0] node387;
	wire [8-1:0] node390;
	wire [8-1:0] node392;
	wire [8-1:0] node395;
	wire [8-1:0] node398;
	wire [8-1:0] node399;
	wire [8-1:0] node400;
	wire [8-1:0] node401;
	wire [8-1:0] node402;
	wire [8-1:0] node403;
	wire [8-1:0] node404;
	wire [8-1:0] node405;
	wire [8-1:0] node406;
	wire [8-1:0] node410;
	wire [8-1:0] node411;
	wire [8-1:0] node415;
	wire [8-1:0] node416;
	wire [8-1:0] node417;
	wire [8-1:0] node419;
	wire [8-1:0] node421;
	wire [8-1:0] node424;
	wire [8-1:0] node426;
	wire [8-1:0] node429;
	wire [8-1:0] node430;
	wire [8-1:0] node431;
	wire [8-1:0] node435;
	wire [8-1:0] node436;
	wire [8-1:0] node439;
	wire [8-1:0] node442;
	wire [8-1:0] node443;
	wire [8-1:0] node444;
	wire [8-1:0] node446;
	wire [8-1:0] node447;
	wire [8-1:0] node451;
	wire [8-1:0] node452;
	wire [8-1:0] node453;
	wire [8-1:0] node456;
	wire [8-1:0] node460;
	wire [8-1:0] node461;
	wire [8-1:0] node462;
	wire [8-1:0] node465;
	wire [8-1:0] node468;
	wire [8-1:0] node469;
	wire [8-1:0] node470;
	wire [8-1:0] node471;
	wire [8-1:0] node475;
	wire [8-1:0] node476;
	wire [8-1:0] node480;
	wire [8-1:0] node481;
	wire [8-1:0] node483;
	wire [8-1:0] node486;
	wire [8-1:0] node487;
	wire [8-1:0] node491;
	wire [8-1:0] node492;
	wire [8-1:0] node493;
	wire [8-1:0] node494;
	wire [8-1:0] node495;
	wire [8-1:0] node498;
	wire [8-1:0] node499;
	wire [8-1:0] node503;
	wire [8-1:0] node504;
	wire [8-1:0] node506;
	wire [8-1:0] node509;
	wire [8-1:0] node511;
	wire [8-1:0] node514;
	wire [8-1:0] node515;
	wire [8-1:0] node516;
	wire [8-1:0] node517;
	wire [8-1:0] node521;
	wire [8-1:0] node522;
	wire [8-1:0] node526;
	wire [8-1:0] node527;
	wire [8-1:0] node529;
	wire [8-1:0] node531;
	wire [8-1:0] node534;
	wire [8-1:0] node535;
	wire [8-1:0] node539;
	wire [8-1:0] node540;
	wire [8-1:0] node541;
	wire [8-1:0] node542;
	wire [8-1:0] node545;
	wire [8-1:0] node546;
	wire [8-1:0] node547;
	wire [8-1:0] node552;
	wire [8-1:0] node553;
	wire [8-1:0] node554;
	wire [8-1:0] node555;
	wire [8-1:0] node559;
	wire [8-1:0] node562;
	wire [8-1:0] node563;
	wire [8-1:0] node566;
	wire [8-1:0] node569;
	wire [8-1:0] node570;
	wire [8-1:0] node571;
	wire [8-1:0] node574;
	wire [8-1:0] node575;
	wire [8-1:0] node579;
	wire [8-1:0] node580;
	wire [8-1:0] node581;
	wire [8-1:0] node582;
	wire [8-1:0] node585;
	wire [8-1:0] node589;
	wire [8-1:0] node590;
	wire [8-1:0] node594;
	wire [8-1:0] node595;
	wire [8-1:0] node596;
	wire [8-1:0] node597;
	wire [8-1:0] node599;
	wire [8-1:0] node601;
	wire [8-1:0] node604;
	wire [8-1:0] node605;
	wire [8-1:0] node606;
	wire [8-1:0] node610;
	wire [8-1:0] node611;
	wire [8-1:0] node614;
	wire [8-1:0] node616;
	wire [8-1:0] node619;
	wire [8-1:0] node620;
	wire [8-1:0] node621;
	wire [8-1:0] node623;
	wire [8-1:0] node626;
	wire [8-1:0] node628;
	wire [8-1:0] node631;
	wire [8-1:0] node632;
	wire [8-1:0] node633;
	wire [8-1:0] node635;
	wire [8-1:0] node638;
	wire [8-1:0] node639;
	wire [8-1:0] node642;
	wire [8-1:0] node645;
	wire [8-1:0] node648;
	wire [8-1:0] node649;
	wire [8-1:0] node650;
	wire [8-1:0] node651;
	wire [8-1:0] node652;
	wire [8-1:0] node655;
	wire [8-1:0] node658;
	wire [8-1:0] node659;
	wire [8-1:0] node660;
	wire [8-1:0] node664;
	wire [8-1:0] node665;
	wire [8-1:0] node668;
	wire [8-1:0] node669;
	wire [8-1:0] node673;
	wire [8-1:0] node674;
	wire [8-1:0] node675;
	wire [8-1:0] node678;
	wire [8-1:0] node681;
	wire [8-1:0] node682;
	wire [8-1:0] node683;
	wire [8-1:0] node685;
	wire [8-1:0] node689;
	wire [8-1:0] node690;
	wire [8-1:0] node692;
	wire [8-1:0] node696;
	wire [8-1:0] node697;
	wire [8-1:0] node698;
	wire [8-1:0] node699;
	wire [8-1:0] node701;
	wire [8-1:0] node704;
	wire [8-1:0] node706;
	wire [8-1:0] node707;
	wire [8-1:0] node711;
	wire [8-1:0] node712;
	wire [8-1:0] node714;
	wire [8-1:0] node715;
	wire [8-1:0] node719;
	wire [8-1:0] node720;
	wire [8-1:0] node723;
	wire [8-1:0] node724;
	wire [8-1:0] node728;
	wire [8-1:0] node729;
	wire [8-1:0] node731;
	wire [8-1:0] node732;
	wire [8-1:0] node735;
	wire [8-1:0] node736;
	wire [8-1:0] node739;
	wire [8-1:0] node742;
	wire [8-1:0] node743;
	wire [8-1:0] node745;
	wire [8-1:0] node748;
	wire [8-1:0] node749;
	wire [8-1:0] node750;
	wire [8-1:0] node753;
	wire [8-1:0] node756;
	wire [8-1:0] node759;
	wire [8-1:0] node760;
	wire [8-1:0] node761;
	wire [8-1:0] node762;
	wire [8-1:0] node763;
	wire [8-1:0] node764;
	wire [8-1:0] node765;
	wire [8-1:0] node767;
	wire [8-1:0] node770;
	wire [8-1:0] node772;
	wire [8-1:0] node775;
	wire [8-1:0] node777;
	wire [8-1:0] node780;
	wire [8-1:0] node781;
	wire [8-1:0] node782;
	wire [8-1:0] node784;
	wire [8-1:0] node787;
	wire [8-1:0] node789;
	wire [8-1:0] node792;
	wire [8-1:0] node794;
	wire [8-1:0] node797;
	wire [8-1:0] node798;
	wire [8-1:0] node799;
	wire [8-1:0] node800;
	wire [8-1:0] node804;
	wire [8-1:0] node805;
	wire [8-1:0] node809;
	wire [8-1:0] node811;
	wire [8-1:0] node814;
	wire [8-1:0] node815;
	wire [8-1:0] node816;
	wire [8-1:0] node817;
	wire [8-1:0] node818;
	wire [8-1:0] node819;
	wire [8-1:0] node823;
	wire [8-1:0] node825;
	wire [8-1:0] node828;
	wire [8-1:0] node829;
	wire [8-1:0] node830;
	wire [8-1:0] node833;
	wire [8-1:0] node836;
	wire [8-1:0] node837;
	wire [8-1:0] node840;
	wire [8-1:0] node843;
	wire [8-1:0] node844;
	wire [8-1:0] node845;
	wire [8-1:0] node846;
	wire [8-1:0] node847;
	wire [8-1:0] node850;
	wire [8-1:0] node853;
	wire [8-1:0] node854;
	wire [8-1:0] node857;
	wire [8-1:0] node860;
	wire [8-1:0] node861;
	wire [8-1:0] node862;
	wire [8-1:0] node865;
	wire [8-1:0] node868;
	wire [8-1:0] node869;
	wire [8-1:0] node873;
	wire [8-1:0] node874;
	wire [8-1:0] node875;
	wire [8-1:0] node876;
	wire [8-1:0] node880;
	wire [8-1:0] node881;
	wire [8-1:0] node884;
	wire [8-1:0] node887;
	wire [8-1:0] node889;
	wire [8-1:0] node890;
	wire [8-1:0] node893;
	wire [8-1:0] node896;
	wire [8-1:0] node897;
	wire [8-1:0] node898;
	wire [8-1:0] node899;
	wire [8-1:0] node900;
	wire [8-1:0] node903;
	wire [8-1:0] node906;
	wire [8-1:0] node908;
	wire [8-1:0] node911;
	wire [8-1:0] node912;
	wire [8-1:0] node913;
	wire [8-1:0] node914;
	wire [8-1:0] node917;
	wire [8-1:0] node921;
	wire [8-1:0] node922;
	wire [8-1:0] node923;
	wire [8-1:0] node926;
	wire [8-1:0] node930;
	wire [8-1:0] node931;
	wire [8-1:0] node932;
	wire [8-1:0] node934;
	wire [8-1:0] node937;
	wire [8-1:0] node938;
	wire [8-1:0] node940;
	wire [8-1:0] node943;
	wire [8-1:0] node946;
	wire [8-1:0] node947;
	wire [8-1:0] node948;
	wire [8-1:0] node949;
	wire [8-1:0] node953;
	wire [8-1:0] node956;
	wire [8-1:0] node957;
	wire [8-1:0] node960;
	wire [8-1:0] node963;
	wire [8-1:0] node964;
	wire [8-1:0] node965;
	wire [8-1:0] node966;
	wire [8-1:0] node967;
	wire [8-1:0] node968;
	wire [8-1:0] node972;
	wire [8-1:0] node973;
	wire [8-1:0] node976;
	wire [8-1:0] node979;
	wire [8-1:0] node980;
	wire [8-1:0] node981;
	wire [8-1:0] node984;
	wire [8-1:0] node987;
	wire [8-1:0] node988;
	wire [8-1:0] node991;
	wire [8-1:0] node994;
	wire [8-1:0] node995;
	wire [8-1:0] node996;
	wire [8-1:0] node997;
	wire [8-1:0] node999;
	wire [8-1:0] node1002;
	wire [8-1:0] node1003;
	wire [8-1:0] node1007;
	wire [8-1:0] node1008;
	wire [8-1:0] node1010;
	wire [8-1:0] node1014;
	wire [8-1:0] node1015;
	wire [8-1:0] node1016;
	wire [8-1:0] node1019;
	wire [8-1:0] node1022;
	wire [8-1:0] node1023;
	wire [8-1:0] node1025;
	wire [8-1:0] node1026;
	wire [8-1:0] node1030;
	wire [8-1:0] node1031;
	wire [8-1:0] node1035;
	wire [8-1:0] node1036;
	wire [8-1:0] node1037;
	wire [8-1:0] node1038;
	wire [8-1:0] node1039;
	wire [8-1:0] node1040;
	wire [8-1:0] node1043;
	wire [8-1:0] node1045;
	wire [8-1:0] node1048;
	wire [8-1:0] node1050;
	wire [8-1:0] node1051;
	wire [8-1:0] node1055;
	wire [8-1:0] node1056;
	wire [8-1:0] node1058;
	wire [8-1:0] node1061;
	wire [8-1:0] node1062;
	wire [8-1:0] node1066;
	wire [8-1:0] node1067;
	wire [8-1:0] node1068;
	wire [8-1:0] node1069;
	wire [8-1:0] node1073;
	wire [8-1:0] node1074;
	wire [8-1:0] node1077;
	wire [8-1:0] node1078;
	wire [8-1:0] node1082;
	wire [8-1:0] node1083;
	wire [8-1:0] node1084;
	wire [8-1:0] node1086;
	wire [8-1:0] node1089;
	wire [8-1:0] node1091;
	wire [8-1:0] node1094;
	wire [8-1:0] node1095;
	wire [8-1:0] node1096;
	wire [8-1:0] node1100;
	wire [8-1:0] node1101;
	wire [8-1:0] node1105;
	wire [8-1:0] node1106;
	wire [8-1:0] node1107;
	wire [8-1:0] node1108;
	wire [8-1:0] node1109;
	wire [8-1:0] node1112;
	wire [8-1:0] node1115;
	wire [8-1:0] node1116;
	wire [8-1:0] node1119;
	wire [8-1:0] node1122;
	wire [8-1:0] node1123;
	wire [8-1:0] node1126;
	wire [8-1:0] node1129;
	wire [8-1:0] node1130;
	wire [8-1:0] node1131;
	wire [8-1:0] node1132;
	wire [8-1:0] node1133;
	wire [8-1:0] node1137;
	wire [8-1:0] node1140;
	wire [8-1:0] node1141;
	wire [8-1:0] node1145;
	wire [8-1:0] node1146;
	wire [8-1:0] node1147;
	wire [8-1:0] node1150;
	wire [8-1:0] node1151;
	wire [8-1:0] node1155;
	wire [8-1:0] node1156;
	wire [8-1:0] node1157;
	wire [8-1:0] node1160;
	wire [8-1:0] node1164;
	wire [8-1:0] node1165;
	wire [8-1:0] node1166;
	wire [8-1:0] node1167;
	wire [8-1:0] node1168;
	wire [8-1:0] node1170;
	wire [8-1:0] node1171;
	wire [8-1:0] node1175;
	wire [8-1:0] node1176;
	wire [8-1:0] node1178;
	wire [8-1:0] node1181;
	wire [8-1:0] node1182;
	wire [8-1:0] node1183;
	wire [8-1:0] node1186;
	wire [8-1:0] node1190;
	wire [8-1:0] node1191;
	wire [8-1:0] node1192;
	wire [8-1:0] node1193;
	wire [8-1:0] node1194;
	wire [8-1:0] node1197;
	wire [8-1:0] node1198;
	wire [8-1:0] node1202;
	wire [8-1:0] node1203;
	wire [8-1:0] node1204;
	wire [8-1:0] node1206;
	wire [8-1:0] node1210;
	wire [8-1:0] node1211;
	wire [8-1:0] node1215;
	wire [8-1:0] node1216;
	wire [8-1:0] node1217;
	wire [8-1:0] node1218;
	wire [8-1:0] node1221;
	wire [8-1:0] node1224;
	wire [8-1:0] node1225;
	wire [8-1:0] node1228;
	wire [8-1:0] node1231;
	wire [8-1:0] node1232;
	wire [8-1:0] node1236;
	wire [8-1:0] node1237;
	wire [8-1:0] node1238;
	wire [8-1:0] node1239;
	wire [8-1:0] node1241;
	wire [8-1:0] node1242;
	wire [8-1:0] node1245;
	wire [8-1:0] node1248;
	wire [8-1:0] node1249;
	wire [8-1:0] node1252;
	wire [8-1:0] node1255;
	wire [8-1:0] node1256;
	wire [8-1:0] node1257;
	wire [8-1:0] node1258;
	wire [8-1:0] node1261;
	wire [8-1:0] node1265;
	wire [8-1:0] node1266;
	wire [8-1:0] node1269;
	wire [8-1:0] node1272;
	wire [8-1:0] node1273;
	wire [8-1:0] node1274;
	wire [8-1:0] node1275;
	wire [8-1:0] node1280;
	wire [8-1:0] node1281;
	wire [8-1:0] node1285;
	wire [8-1:0] node1286;
	wire [8-1:0] node1287;
	wire [8-1:0] node1288;
	wire [8-1:0] node1289;
	wire [8-1:0] node1290;
	wire [8-1:0] node1292;
	wire [8-1:0] node1296;
	wire [8-1:0] node1298;
	wire [8-1:0] node1301;
	wire [8-1:0] node1302;
	wire [8-1:0] node1303;
	wire [8-1:0] node1304;
	wire [8-1:0] node1305;
	wire [8-1:0] node1308;
	wire [8-1:0] node1311;
	wire [8-1:0] node1312;
	wire [8-1:0] node1315;
	wire [8-1:0] node1318;
	wire [8-1:0] node1320;
	wire [8-1:0] node1322;
	wire [8-1:0] node1325;
	wire [8-1:0] node1326;
	wire [8-1:0] node1327;
	wire [8-1:0] node1330;
	wire [8-1:0] node1333;
	wire [8-1:0] node1335;
	wire [8-1:0] node1338;
	wire [8-1:0] node1339;
	wire [8-1:0] node1340;
	wire [8-1:0] node1342;
	wire [8-1:0] node1345;
	wire [8-1:0] node1346;
	wire [8-1:0] node1347;
	wire [8-1:0] node1351;
	wire [8-1:0] node1352;
	wire [8-1:0] node1356;
	wire [8-1:0] node1357;
	wire [8-1:0] node1358;
	wire [8-1:0] node1359;
	wire [8-1:0] node1362;
	wire [8-1:0] node1365;
	wire [8-1:0] node1366;
	wire [8-1:0] node1369;
	wire [8-1:0] node1372;
	wire [8-1:0] node1373;
	wire [8-1:0] node1374;
	wire [8-1:0] node1377;
	wire [8-1:0] node1380;
	wire [8-1:0] node1381;
	wire [8-1:0] node1384;
	wire [8-1:0] node1387;
	wire [8-1:0] node1388;
	wire [8-1:0] node1389;
	wire [8-1:0] node1391;
	wire [8-1:0] node1392;
	wire [8-1:0] node1395;
	wire [8-1:0] node1398;
	wire [8-1:0] node1400;
	wire [8-1:0] node1403;
	wire [8-1:0] node1404;
	wire [8-1:0] node1406;
	wire [8-1:0] node1410;
	wire [8-1:0] node1411;
	wire [8-1:0] node1412;
	wire [8-1:0] node1413;
	wire [8-1:0] node1414;
	wire [8-1:0] node1415;
	wire [8-1:0] node1416;
	wire [8-1:0] node1419;
	wire [8-1:0] node1422;
	wire [8-1:0] node1424;
	wire [8-1:0] node1425;
	wire [8-1:0] node1427;
	wire [8-1:0] node1430;
	wire [8-1:0] node1433;
	wire [8-1:0] node1434;
	wire [8-1:0] node1435;
	wire [8-1:0] node1438;
	wire [8-1:0] node1441;
	wire [8-1:0] node1442;
	wire [8-1:0] node1443;
	wire [8-1:0] node1447;
	wire [8-1:0] node1448;
	wire [8-1:0] node1452;
	wire [8-1:0] node1453;
	wire [8-1:0] node1454;
	wire [8-1:0] node1455;
	wire [8-1:0] node1457;
	wire [8-1:0] node1458;
	wire [8-1:0] node1461;
	wire [8-1:0] node1464;
	wire [8-1:0] node1465;
	wire [8-1:0] node1467;
	wire [8-1:0] node1470;
	wire [8-1:0] node1473;
	wire [8-1:0] node1474;
	wire [8-1:0] node1476;
	wire [8-1:0] node1479;
	wire [8-1:0] node1480;
	wire [8-1:0] node1481;
	wire [8-1:0] node1484;
	wire [8-1:0] node1487;
	wire [8-1:0] node1488;
	wire [8-1:0] node1491;
	wire [8-1:0] node1494;
	wire [8-1:0] node1495;
	wire [8-1:0] node1496;
	wire [8-1:0] node1497;
	wire [8-1:0] node1499;
	wire [8-1:0] node1502;
	wire [8-1:0] node1503;
	wire [8-1:0] node1506;
	wire [8-1:0] node1509;
	wire [8-1:0] node1510;
	wire [8-1:0] node1512;
	wire [8-1:0] node1515;
	wire [8-1:0] node1516;
	wire [8-1:0] node1520;
	wire [8-1:0] node1521;
	wire [8-1:0] node1522;
	wire [8-1:0] node1524;
	wire [8-1:0] node1527;
	wire [8-1:0] node1529;
	wire [8-1:0] node1532;
	wire [8-1:0] node1535;
	wire [8-1:0] node1536;
	wire [8-1:0] node1537;
	wire [8-1:0] node1538;
	wire [8-1:0] node1539;
	wire [8-1:0] node1542;
	wire [8-1:0] node1545;
	wire [8-1:0] node1546;
	wire [8-1:0] node1548;
	wire [8-1:0] node1549;
	wire [8-1:0] node1553;
	wire [8-1:0] node1554;
	wire [8-1:0] node1558;
	wire [8-1:0] node1559;
	wire [8-1:0] node1560;
	wire [8-1:0] node1562;
	wire [8-1:0] node1565;
	wire [8-1:0] node1567;
	wire [8-1:0] node1570;
	wire [8-1:0] node1571;
	wire [8-1:0] node1574;
	wire [8-1:0] node1575;
	wire [8-1:0] node1576;
	wire [8-1:0] node1581;
	wire [8-1:0] node1582;
	wire [8-1:0] node1583;
	wire [8-1:0] node1584;
	wire [8-1:0] node1586;
	wire [8-1:0] node1589;
	wire [8-1:0] node1590;
	wire [8-1:0] node1592;
	wire [8-1:0] node1595;
	wire [8-1:0] node1597;
	wire [8-1:0] node1600;
	wire [8-1:0] node1601;
	wire [8-1:0] node1603;
	wire [8-1:0] node1606;
	wire [8-1:0] node1607;
	wire [8-1:0] node1610;
	wire [8-1:0] node1611;
	wire [8-1:0] node1614;
	wire [8-1:0] node1617;
	wire [8-1:0] node1618;
	wire [8-1:0] node1619;
	wire [8-1:0] node1620;
	wire [8-1:0] node1622;
	wire [8-1:0] node1626;
	wire [8-1:0] node1627;
	wire [8-1:0] node1628;
	wire [8-1:0] node1633;
	wire [8-1:0] node1634;
	wire [8-1:0] node1636;
	wire [8-1:0] node1639;
	wire [8-1:0] node1640;
	wire [8-1:0] node1644;
	wire [8-1:0] node1645;
	wire [8-1:0] node1646;
	wire [8-1:0] node1647;
	wire [8-1:0] node1648;
	wire [8-1:0] node1649;
	wire [8-1:0] node1652;
	wire [8-1:0] node1654;
	wire [8-1:0] node1657;
	wire [8-1:0] node1659;
	wire [8-1:0] node1662;
	wire [8-1:0] node1663;
	wire [8-1:0] node1665;
	wire [8-1:0] node1668;
	wire [8-1:0] node1669;
	wire [8-1:0] node1671;
	wire [8-1:0] node1674;
	wire [8-1:0] node1676;
	wire [8-1:0] node1679;
	wire [8-1:0] node1680;
	wire [8-1:0] node1681;
	wire [8-1:0] node1682;
	wire [8-1:0] node1683;
	wire [8-1:0] node1684;
	wire [8-1:0] node1687;
	wire [8-1:0] node1690;
	wire [8-1:0] node1691;
	wire [8-1:0] node1694;
	wire [8-1:0] node1697;
	wire [8-1:0] node1698;
	wire [8-1:0] node1699;
	wire [8-1:0] node1702;
	wire [8-1:0] node1705;
	wire [8-1:0] node1706;
	wire [8-1:0] node1709;
	wire [8-1:0] node1712;
	wire [8-1:0] node1713;
	wire [8-1:0] node1715;
	wire [8-1:0] node1717;
	wire [8-1:0] node1720;
	wire [8-1:0] node1721;
	wire [8-1:0] node1722;
	wire [8-1:0] node1725;
	wire [8-1:0] node1728;
	wire [8-1:0] node1730;
	wire [8-1:0] node1733;
	wire [8-1:0] node1734;
	wire [8-1:0] node1735;
	wire [8-1:0] node1736;
	wire [8-1:0] node1737;
	wire [8-1:0] node1740;
	wire [8-1:0] node1743;
	wire [8-1:0] node1744;
	wire [8-1:0] node1747;
	wire [8-1:0] node1750;
	wire [8-1:0] node1751;
	wire [8-1:0] node1752;
	wire [8-1:0] node1755;
	wire [8-1:0] node1758;
	wire [8-1:0] node1759;
	wire [8-1:0] node1762;
	wire [8-1:0] node1765;
	wire [8-1:0] node1766;
	wire [8-1:0] node1767;
	wire [8-1:0] node1768;
	wire [8-1:0] node1771;
	wire [8-1:0] node1775;
	wire [8-1:0] node1776;
	wire [8-1:0] node1778;
	wire [8-1:0] node1781;
	wire [8-1:0] node1782;
	wire [8-1:0] node1785;
	wire [8-1:0] node1788;
	wire [8-1:0] node1789;
	wire [8-1:0] node1790;
	wire [8-1:0] node1791;
	wire [8-1:0] node1792;
	wire [8-1:0] node1793;
	wire [8-1:0] node1795;
	wire [8-1:0] node1798;
	wire [8-1:0] node1800;
	wire [8-1:0] node1803;
	wire [8-1:0] node1804;
	wire [8-1:0] node1807;
	wire [8-1:0] node1810;
	wire [8-1:0] node1811;
	wire [8-1:0] node1812;
	wire [8-1:0] node1814;
	wire [8-1:0] node1817;
	wire [8-1:0] node1819;
	wire [8-1:0] node1822;
	wire [8-1:0] node1825;
	wire [8-1:0] node1826;
	wire [8-1:0] node1827;
	wire [8-1:0] node1828;
	wire [8-1:0] node1829;
	wire [8-1:0] node1834;
	wire [8-1:0] node1835;
	wire [8-1:0] node1838;
	wire [8-1:0] node1839;
	wire [8-1:0] node1843;
	wire [8-1:0] node1844;
	wire [8-1:0] node1845;
	wire [8-1:0] node1848;
	wire [8-1:0] node1851;
	wire [8-1:0] node1854;
	wire [8-1:0] node1855;
	wire [8-1:0] node1856;
	wire [8-1:0] node1857;
	wire [8-1:0] node1858;
	wire [8-1:0] node1859;
	wire [8-1:0] node1863;
	wire [8-1:0] node1864;
	wire [8-1:0] node1868;
	wire [8-1:0] node1869;
	wire [8-1:0] node1870;
	wire [8-1:0] node1873;
	wire [8-1:0] node1876;
	wire [8-1:0] node1878;
	wire [8-1:0] node1881;
	wire [8-1:0] node1882;
	wire [8-1:0] node1885;
	wire [8-1:0] node1888;
	wire [8-1:0] node1889;
	wire [8-1:0] node1890;
	wire [8-1:0] node1891;
	wire [8-1:0] node1893;
	wire [8-1:0] node1896;
	wire [8-1:0] node1897;
	wire [8-1:0] node1901;
	wire [8-1:0] node1902;
	wire [8-1:0] node1903;
	wire [8-1:0] node1906;
	wire [8-1:0] node1909;
	wire [8-1:0] node1910;
	wire [8-1:0] node1913;
	wire [8-1:0] node1916;
	wire [8-1:0] node1919;
	wire [8-1:0] node1920;
	wire [8-1:0] node1921;
	wire [8-1:0] node1922;
	wire [8-1:0] node1923;
	wire [8-1:0] node1924;
	wire [8-1:0] node1925;
	wire [8-1:0] node1926;
	wire [8-1:0] node1930;
	wire [8-1:0] node1932;
	wire [8-1:0] node1935;
	wire [8-1:0] node1936;
	wire [8-1:0] node1937;
	wire [8-1:0] node1941;
	wire [8-1:0] node1943;
	wire [8-1:0] node1946;
	wire [8-1:0] node1947;
	wire [8-1:0] node1948;
	wire [8-1:0] node1949;
	wire [8-1:0] node1950;
	wire [8-1:0] node1951;
	wire [8-1:0] node1954;
	wire [8-1:0] node1956;
	wire [8-1:0] node1959;
	wire [8-1:0] node1961;
	wire [8-1:0] node1964;
	wire [8-1:0] node1965;
	wire [8-1:0] node1966;
	wire [8-1:0] node1970;
	wire [8-1:0] node1971;
	wire [8-1:0] node1972;
	wire [8-1:0] node1976;
	wire [8-1:0] node1978;
	wire [8-1:0] node1981;
	wire [8-1:0] node1982;
	wire [8-1:0] node1983;
	wire [8-1:0] node1987;
	wire [8-1:0] node1988;
	wire [8-1:0] node1990;
	wire [8-1:0] node1993;
	wire [8-1:0] node1995;
	wire [8-1:0] node1998;
	wire [8-1:0] node1999;
	wire [8-1:0] node2000;
	wire [8-1:0] node2001;
	wire [8-1:0] node2003;
	wire [8-1:0] node2006;
	wire [8-1:0] node2007;
	wire [8-1:0] node2011;
	wire [8-1:0] node2012;
	wire [8-1:0] node2016;
	wire [8-1:0] node2017;
	wire [8-1:0] node2018;
	wire [8-1:0] node2020;
	wire [8-1:0] node2023;
	wire [8-1:0] node2025;
	wire [8-1:0] node2026;
	wire [8-1:0] node2029;
	wire [8-1:0] node2032;
	wire [8-1:0] node2033;
	wire [8-1:0] node2034;
	wire [8-1:0] node2036;
	wire [8-1:0] node2039;
	wire [8-1:0] node2041;
	wire [8-1:0] node2044;
	wire [8-1:0] node2046;
	wire [8-1:0] node2049;
	wire [8-1:0] node2050;
	wire [8-1:0] node2051;
	wire [8-1:0] node2052;
	wire [8-1:0] node2054;
	wire [8-1:0] node2057;
	wire [8-1:0] node2059;
	wire [8-1:0] node2062;
	wire [8-1:0] node2063;
	wire [8-1:0] node2064;
	wire [8-1:0] node2065;
	wire [8-1:0] node2067;
	wire [8-1:0] node2070;
	wire [8-1:0] node2072;
	wire [8-1:0] node2075;
	wire [8-1:0] node2076;
	wire [8-1:0] node2080;
	wire [8-1:0] node2081;
	wire [8-1:0] node2082;
	wire [8-1:0] node2083;
	wire [8-1:0] node2087;
	wire [8-1:0] node2089;
	wire [8-1:0] node2092;
	wire [8-1:0] node2093;
	wire [8-1:0] node2097;
	wire [8-1:0] node2098;
	wire [8-1:0] node2099;
	wire [8-1:0] node2100;
	wire [8-1:0] node2101;
	wire [8-1:0] node2105;
	wire [8-1:0] node2106;
	wire [8-1:0] node2110;
	wire [8-1:0] node2112;
	wire [8-1:0] node2115;
	wire [8-1:0] node2116;
	wire [8-1:0] node2120;
	wire [8-1:0] node2121;
	wire [8-1:0] node2122;
	wire [8-1:0] node2123;
	wire [8-1:0] node2124;
	wire [8-1:0] node2125;
	wire [8-1:0] node2127;
	wire [8-1:0] node2130;
	wire [8-1:0] node2131;
	wire [8-1:0] node2133;
	wire [8-1:0] node2136;
	wire [8-1:0] node2138;
	wire [8-1:0] node2141;
	wire [8-1:0] node2142;
	wire [8-1:0] node2143;
	wire [8-1:0] node2145;
	wire [8-1:0] node2148;
	wire [8-1:0] node2149;
	wire [8-1:0] node2152;
	wire [8-1:0] node2153;
	wire [8-1:0] node2156;
	wire [8-1:0] node2159;
	wire [8-1:0] node2160;
	wire [8-1:0] node2162;
	wire [8-1:0] node2165;
	wire [8-1:0] node2166;
	wire [8-1:0] node2169;
	wire [8-1:0] node2170;
	wire [8-1:0] node2173;
	wire [8-1:0] node2176;
	wire [8-1:0] node2177;
	wire [8-1:0] node2178;
	wire [8-1:0] node2179;
	wire [8-1:0] node2180;
	wire [8-1:0] node2181;
	wire [8-1:0] node2182;
	wire [8-1:0] node2185;
	wire [8-1:0] node2189;
	wire [8-1:0] node2190;
	wire [8-1:0] node2193;
	wire [8-1:0] node2196;
	wire [8-1:0] node2197;
	wire [8-1:0] node2198;
	wire [8-1:0] node2201;
	wire [8-1:0] node2204;
	wire [8-1:0] node2206;
	wire [8-1:0] node2209;
	wire [8-1:0] node2210;
	wire [8-1:0] node2211;
	wire [8-1:0] node2212;
	wire [8-1:0] node2215;
	wire [8-1:0] node2218;
	wire [8-1:0] node2219;
	wire [8-1:0] node2222;
	wire [8-1:0] node2225;
	wire [8-1:0] node2226;
	wire [8-1:0] node2227;
	wire [8-1:0] node2231;
	wire [8-1:0] node2232;
	wire [8-1:0] node2236;
	wire [8-1:0] node2237;
	wire [8-1:0] node2238;
	wire [8-1:0] node2239;
	wire [8-1:0] node2240;
	wire [8-1:0] node2243;
	wire [8-1:0] node2246;
	wire [8-1:0] node2247;
	wire [8-1:0] node2250;
	wire [8-1:0] node2253;
	wire [8-1:0] node2254;
	wire [8-1:0] node2255;
	wire [8-1:0] node2256;
	wire [8-1:0] node2259;
	wire [8-1:0] node2262;
	wire [8-1:0] node2263;
	wire [8-1:0] node2267;
	wire [8-1:0] node2268;
	wire [8-1:0] node2269;
	wire [8-1:0] node2272;
	wire [8-1:0] node2276;
	wire [8-1:0] node2277;
	wire [8-1:0] node2278;
	wire [8-1:0] node2279;
	wire [8-1:0] node2280;
	wire [8-1:0] node2284;
	wire [8-1:0] node2285;
	wire [8-1:0] node2289;
	wire [8-1:0] node2290;
	wire [8-1:0] node2293;
	wire [8-1:0] node2296;
	wire [8-1:0] node2297;
	wire [8-1:0] node2298;
	wire [8-1:0] node2301;
	wire [8-1:0] node2304;
	wire [8-1:0] node2305;
	wire [8-1:0] node2309;
	wire [8-1:0] node2310;
	wire [8-1:0] node2311;
	wire [8-1:0] node2312;
	wire [8-1:0] node2313;
	wire [8-1:0] node2316;
	wire [8-1:0] node2317;
	wire [8-1:0] node2320;
	wire [8-1:0] node2323;
	wire [8-1:0] node2324;
	wire [8-1:0] node2325;
	wire [8-1:0] node2328;
	wire [8-1:0] node2329;
	wire [8-1:0] node2332;
	wire [8-1:0] node2335;
	wire [8-1:0] node2336;
	wire [8-1:0] node2339;
	wire [8-1:0] node2340;
	wire [8-1:0] node2343;
	wire [8-1:0] node2346;
	wire [8-1:0] node2347;
	wire [8-1:0] node2348;
	wire [8-1:0] node2349;
	wire [8-1:0] node2350;
	wire [8-1:0] node2351;
	wire [8-1:0] node2354;
	wire [8-1:0] node2357;
	wire [8-1:0] node2358;
	wire [8-1:0] node2362;
	wire [8-1:0] node2363;
	wire [8-1:0] node2364;
	wire [8-1:0] node2367;
	wire [8-1:0] node2370;
	wire [8-1:0] node2371;
	wire [8-1:0] node2375;
	wire [8-1:0] node2376;
	wire [8-1:0] node2377;
	wire [8-1:0] node2378;
	wire [8-1:0] node2381;
	wire [8-1:0] node2384;
	wire [8-1:0] node2387;
	wire [8-1:0] node2388;
	wire [8-1:0] node2389;
	wire [8-1:0] node2392;
	wire [8-1:0] node2395;
	wire [8-1:0] node2397;
	wire [8-1:0] node2400;
	wire [8-1:0] node2401;
	wire [8-1:0] node2402;
	wire [8-1:0] node2403;
	wire [8-1:0] node2404;
	wire [8-1:0] node2408;
	wire [8-1:0] node2411;
	wire [8-1:0] node2412;
	wire [8-1:0] node2413;
	wire [8-1:0] node2417;
	wire [8-1:0] node2418;
	wire [8-1:0] node2421;
	wire [8-1:0] node2424;
	wire [8-1:0] node2425;
	wire [8-1:0] node2426;
	wire [8-1:0] node2429;
	wire [8-1:0] node2430;
	wire [8-1:0] node2434;
	wire [8-1:0] node2435;
	wire [8-1:0] node2436;
	wire [8-1:0] node2439;
	wire [8-1:0] node2443;
	wire [8-1:0] node2444;
	wire [8-1:0] node2445;
	wire [8-1:0] node2446;
	wire [8-1:0] node2447;
	wire [8-1:0] node2450;
	wire [8-1:0] node2451;
	wire [8-1:0] node2454;
	wire [8-1:0] node2457;
	wire [8-1:0] node2458;
	wire [8-1:0] node2459;
	wire [8-1:0] node2460;
	wire [8-1:0] node2463;
	wire [8-1:0] node2466;
	wire [8-1:0] node2467;
	wire [8-1:0] node2470;
	wire [8-1:0] node2473;
	wire [8-1:0] node2474;
	wire [8-1:0] node2475;
	wire [8-1:0] node2479;
	wire [8-1:0] node2481;
	wire [8-1:0] node2484;
	wire [8-1:0] node2485;
	wire [8-1:0] node2486;
	wire [8-1:0] node2488;
	wire [8-1:0] node2490;
	wire [8-1:0] node2493;
	wire [8-1:0] node2494;
	wire [8-1:0] node2495;
	wire [8-1:0] node2499;
	wire [8-1:0] node2501;
	wire [8-1:0] node2504;
	wire [8-1:0] node2505;
	wire [8-1:0] node2506;
	wire [8-1:0] node2509;
	wire [8-1:0] node2512;
	wire [8-1:0] node2513;
	wire [8-1:0] node2516;
	wire [8-1:0] node2519;
	wire [8-1:0] node2520;
	wire [8-1:0] node2521;
	wire [8-1:0] node2522;
	wire [8-1:0] node2525;
	wire [8-1:0] node2526;
	wire [8-1:0] node2529;
	wire [8-1:0] node2532;
	wire [8-1:0] node2533;
	wire [8-1:0] node2534;
	wire [8-1:0] node2535;
	wire [8-1:0] node2538;
	wire [8-1:0] node2541;
	wire [8-1:0] node2544;
	wire [8-1:0] node2545;
	wire [8-1:0] node2547;
	wire [8-1:0] node2550;
	wire [8-1:0] node2551;
	wire [8-1:0] node2554;
	wire [8-1:0] node2557;
	wire [8-1:0] node2558;
	wire [8-1:0] node2559;
	wire [8-1:0] node2561;
	wire [8-1:0] node2562;
	wire [8-1:0] node2566;
	wire [8-1:0] node2567;
	wire [8-1:0] node2569;
	wire [8-1:0] node2572;
	wire [8-1:0] node2575;
	wire [8-1:0] node2576;
	wire [8-1:0] node2577;
	wire [8-1:0] node2580;
	wire [8-1:0] node2583;
	wire [8-1:0] node2584;
	wire [8-1:0] node2587;
	wire [8-1:0] node2590;
	wire [8-1:0] node2591;
	wire [8-1:0] node2592;
	wire [8-1:0] node2593;
	wire [8-1:0] node2594;
	wire [8-1:0] node2596;
	wire [8-1:0] node2599;
	wire [8-1:0] node2600;
	wire [8-1:0] node2603;
	wire [8-1:0] node2604;
	wire [8-1:0] node2607;
	wire [8-1:0] node2610;
	wire [8-1:0] node2611;
	wire [8-1:0] node2612;
	wire [8-1:0] node2614;
	wire [8-1:0] node2617;
	wire [8-1:0] node2619;
	wire [8-1:0] node2622;
	wire [8-1:0] node2623;
	wire [8-1:0] node2624;
	wire [8-1:0] node2627;
	wire [8-1:0] node2628;
	wire [8-1:0] node2631;
	wire [8-1:0] node2634;
	wire [8-1:0] node2635;
	wire [8-1:0] node2638;
	wire [8-1:0] node2639;
	wire [8-1:0] node2642;
	wire [8-1:0] node2645;
	wire [8-1:0] node2646;
	wire [8-1:0] node2647;
	wire [8-1:0] node2648;
	wire [8-1:0] node2649;
	wire [8-1:0] node2650;
	wire [8-1:0] node2653;
	wire [8-1:0] node2655;
	wire [8-1:0] node2658;
	wire [8-1:0] node2659;
	wire [8-1:0] node2662;
	wire [8-1:0] node2665;
	wire [8-1:0] node2666;
	wire [8-1:0] node2667;
	wire [8-1:0] node2669;
	wire [8-1:0] node2673;
	wire [8-1:0] node2674;
	wire [8-1:0] node2677;
	wire [8-1:0] node2680;
	wire [8-1:0] node2681;
	wire [8-1:0] node2682;
	wire [8-1:0] node2683;
	wire [8-1:0] node2684;
	wire [8-1:0] node2688;
	wire [8-1:0] node2690;
	wire [8-1:0] node2693;
	wire [8-1:0] node2694;
	wire [8-1:0] node2695;
	wire [8-1:0] node2698;
	wire [8-1:0] node2701;
	wire [8-1:0] node2702;
	wire [8-1:0] node2705;
	wire [8-1:0] node2708;
	wire [8-1:0] node2709;
	wire [8-1:0] node2710;
	wire [8-1:0] node2713;
	wire [8-1:0] node2714;
	wire [8-1:0] node2717;
	wire [8-1:0] node2720;
	wire [8-1:0] node2721;
	wire [8-1:0] node2724;
	wire [8-1:0] node2725;
	wire [8-1:0] node2729;
	wire [8-1:0] node2730;
	wire [8-1:0] node2731;
	wire [8-1:0] node2732;
	wire [8-1:0] node2733;
	wire [8-1:0] node2736;
	wire [8-1:0] node2739;
	wire [8-1:0] node2740;
	wire [8-1:0] node2743;
	wire [8-1:0] node2746;
	wire [8-1:0] node2747;
	wire [8-1:0] node2748;
	wire [8-1:0] node2749;
	wire [8-1:0] node2753;
	wire [8-1:0] node2755;
	wire [8-1:0] node2758;
	wire [8-1:0] node2759;
	wire [8-1:0] node2762;
	wire [8-1:0] node2765;
	wire [8-1:0] node2766;
	wire [8-1:0] node2767;
	wire [8-1:0] node2768;
	wire [8-1:0] node2770;
	wire [8-1:0] node2773;
	wire [8-1:0] node2774;
	wire [8-1:0] node2777;
	wire [8-1:0] node2780;
	wire [8-1:0] node2781;
	wire [8-1:0] node2782;
	wire [8-1:0] node2785;
	wire [8-1:0] node2788;
	wire [8-1:0] node2790;
	wire [8-1:0] node2793;
	wire [8-1:0] node2794;
	wire [8-1:0] node2795;
	wire [8-1:0] node2796;
	wire [8-1:0] node2799;
	wire [8-1:0] node2802;
	wire [8-1:0] node2803;
	wire [8-1:0] node2806;
	wire [8-1:0] node2809;
	wire [8-1:0] node2810;
	wire [8-1:0] node2811;
	wire [8-1:0] node2816;
	wire [8-1:0] node2817;
	wire [8-1:0] node2818;
	wire [8-1:0] node2819;
	wire [8-1:0] node2820;
	wire [8-1:0] node2822;
	wire [8-1:0] node2825;
	wire [8-1:0] node2826;
	wire [8-1:0] node2829;
	wire [8-1:0] node2832;
	wire [8-1:0] node2833;
	wire [8-1:0] node2834;
	wire [8-1:0] node2835;
	wire [8-1:0] node2838;
	wire [8-1:0] node2841;
	wire [8-1:0] node2843;
	wire [8-1:0] node2846;
	wire [8-1:0] node2847;
	wire [8-1:0] node2848;
	wire [8-1:0] node2851;
	wire [8-1:0] node2854;
	wire [8-1:0] node2855;
	wire [8-1:0] node2858;
	wire [8-1:0] node2861;
	wire [8-1:0] node2862;
	wire [8-1:0] node2863;
	wire [8-1:0] node2864;
	wire [8-1:0] node2867;
	wire [8-1:0] node2868;
	wire [8-1:0] node2871;
	wire [8-1:0] node2874;
	wire [8-1:0] node2875;
	wire [8-1:0] node2876;
	wire [8-1:0] node2879;
	wire [8-1:0] node2881;
	wire [8-1:0] node2884;
	wire [8-1:0] node2886;
	wire [8-1:0] node2888;
	wire [8-1:0] node2891;
	wire [8-1:0] node2892;
	wire [8-1:0] node2893;
	wire [8-1:0] node2894;
	wire [8-1:0] node2898;
	wire [8-1:0] node2899;
	wire [8-1:0] node2902;
	wire [8-1:0] node2905;
	wire [8-1:0] node2907;
	wire [8-1:0] node2908;
	wire [8-1:0] node2910;
	wire [8-1:0] node2913;
	wire [8-1:0] node2916;
	wire [8-1:0] node2917;
	wire [8-1:0] node2918;
	wire [8-1:0] node2919;
	wire [8-1:0] node2920;
	wire [8-1:0] node2924;
	wire [8-1:0] node2925;
	wire [8-1:0] node2928;
	wire [8-1:0] node2929;
	wire [8-1:0] node2932;
	wire [8-1:0] node2935;
	wire [8-1:0] node2936;
	wire [8-1:0] node2937;
	wire [8-1:0] node2938;
	wire [8-1:0] node2939;
	wire [8-1:0] node2942;
	wire [8-1:0] node2945;
	wire [8-1:0] node2946;
	wire [8-1:0] node2950;
	wire [8-1:0] node2951;
	wire [8-1:0] node2954;
	wire [8-1:0] node2957;
	wire [8-1:0] node2958;
	wire [8-1:0] node2959;
	wire [8-1:0] node2961;
	wire [8-1:0] node2964;
	wire [8-1:0] node2966;
	wire [8-1:0] node2969;
	wire [8-1:0] node2970;
	wire [8-1:0] node2972;
	wire [8-1:0] node2975;
	wire [8-1:0] node2978;
	wire [8-1:0] node2979;
	wire [8-1:0] node2980;
	wire [8-1:0] node2981;
	wire [8-1:0] node2982;
	wire [8-1:0] node2986;
	wire [8-1:0] node2989;
	wire [8-1:0] node2990;
	wire [8-1:0] node2991;
	wire [8-1:0] node2993;
	wire [8-1:0] node2997;
	wire [8-1:0] node2999;
	wire [8-1:0] node3002;
	wire [8-1:0] node3003;
	wire [8-1:0] node3004;
	wire [8-1:0] node3005;
	wire [8-1:0] node3008;
	wire [8-1:0] node3011;
	wire [8-1:0] node3012;
	wire [8-1:0] node3015;
	wire [8-1:0] node3018;
	wire [8-1:0] node3019;
	wire [8-1:0] node3021;
	wire [8-1:0] node3024;
	wire [8-1:0] node3025;
	wire [8-1:0] node3028;
	wire [8-1:0] node3031;
	wire [8-1:0] node3032;
	wire [8-1:0] node3033;
	wire [8-1:0] node3034;
	wire [8-1:0] node3035;
	wire [8-1:0] node3036;
	wire [8-1:0] node3037;
	wire [8-1:0] node3038;
	wire [8-1:0] node3040;
	wire [8-1:0] node3043;
	wire [8-1:0] node3044;
	wire [8-1:0] node3048;
	wire [8-1:0] node3049;
	wire [8-1:0] node3050;
	wire [8-1:0] node3053;
	wire [8-1:0] node3056;
	wire [8-1:0] node3059;
	wire [8-1:0] node3060;
	wire [8-1:0] node3061;
	wire [8-1:0] node3064;
	wire [8-1:0] node3065;
	wire [8-1:0] node3069;
	wire [8-1:0] node3070;
	wire [8-1:0] node3072;
	wire [8-1:0] node3074;
	wire [8-1:0] node3078;
	wire [8-1:0] node3079;
	wire [8-1:0] node3080;
	wire [8-1:0] node3081;
	wire [8-1:0] node3083;
	wire [8-1:0] node3086;
	wire [8-1:0] node3087;
	wire [8-1:0] node3088;
	wire [8-1:0] node3089;
	wire [8-1:0] node3094;
	wire [8-1:0] node3097;
	wire [8-1:0] node3098;
	wire [8-1:0] node3099;
	wire [8-1:0] node3100;
	wire [8-1:0] node3102;
	wire [8-1:0] node3106;
	wire [8-1:0] node3109;
	wire [8-1:0] node3110;
	wire [8-1:0] node3111;
	wire [8-1:0] node3115;
	wire [8-1:0] node3118;
	wire [8-1:0] node3119;
	wire [8-1:0] node3120;
	wire [8-1:0] node3121;
	wire [8-1:0] node3124;
	wire [8-1:0] node3127;
	wire [8-1:0] node3130;
	wire [8-1:0] node3131;
	wire [8-1:0] node3132;
	wire [8-1:0] node3133;
	wire [8-1:0] node3134;
	wire [8-1:0] node3139;
	wire [8-1:0] node3140;
	wire [8-1:0] node3144;
	wire [8-1:0] node3146;
	wire [8-1:0] node3149;
	wire [8-1:0] node3150;
	wire [8-1:0] node3151;
	wire [8-1:0] node3152;
	wire [8-1:0] node3153;
	wire [8-1:0] node3154;
	wire [8-1:0] node3157;
	wire [8-1:0] node3158;
	wire [8-1:0] node3162;
	wire [8-1:0] node3163;
	wire [8-1:0] node3164;
	wire [8-1:0] node3168;
	wire [8-1:0] node3171;
	wire [8-1:0] node3173;
	wire [8-1:0] node3176;
	wire [8-1:0] node3177;
	wire [8-1:0] node3178;
	wire [8-1:0] node3179;
	wire [8-1:0] node3182;
	wire [8-1:0] node3184;
	wire [8-1:0] node3187;
	wire [8-1:0] node3190;
	wire [8-1:0] node3191;
	wire [8-1:0] node3193;
	wire [8-1:0] node3195;
	wire [8-1:0] node3198;
	wire [8-1:0] node3200;
	wire [8-1:0] node3203;
	wire [8-1:0] node3204;
	wire [8-1:0] node3205;
	wire [8-1:0] node3206;
	wire [8-1:0] node3207;
	wire [8-1:0] node3210;
	wire [8-1:0] node3212;
	wire [8-1:0] node3215;
	wire [8-1:0] node3218;
	wire [8-1:0] node3219;
	wire [8-1:0] node3221;
	wire [8-1:0] node3223;
	wire [8-1:0] node3226;
	wire [8-1:0] node3228;
	wire [8-1:0] node3231;
	wire [8-1:0] node3232;
	wire [8-1:0] node3233;
	wire [8-1:0] node3236;
	wire [8-1:0] node3238;
	wire [8-1:0] node3241;
	wire [8-1:0] node3243;
	wire [8-1:0] node3245;
	wire [8-1:0] node3248;
	wire [8-1:0] node3249;
	wire [8-1:0] node3251;
	wire [8-1:0] node3253;
	wire [8-1:0] node3256;
	wire [8-1:0] node3257;
	wire [8-1:0] node3258;
	wire [8-1:0] node3259;
	wire [8-1:0] node3260;
	wire [8-1:0] node3261;
	wire [8-1:0] node3265;
	wire [8-1:0] node3268;
	wire [8-1:0] node3269;
	wire [8-1:0] node3272;
	wire [8-1:0] node3275;
	wire [8-1:0] node3276;
	wire [8-1:0] node3277;
	wire [8-1:0] node3278;
	wire [8-1:0] node3282;
	wire [8-1:0] node3283;
	wire [8-1:0] node3287;
	wire [8-1:0] node3288;
	wire [8-1:0] node3292;
	wire [8-1:0] node3293;
	wire [8-1:0] node3294;
	wire [8-1:0] node3295;
	wire [8-1:0] node3298;
	wire [8-1:0] node3301;
	wire [8-1:0] node3302;
	wire [8-1:0] node3306;
	wire [8-1:0] node3307;
	wire [8-1:0] node3308;
	wire [8-1:0] node3312;
	wire [8-1:0] node3313;
	wire [8-1:0] node3316;
	wire [8-1:0] node3319;
	wire [8-1:0] node3320;
	wire [8-1:0] node3321;
	wire [8-1:0] node3322;
	wire [8-1:0] node3323;
	wire [8-1:0] node3324;
	wire [8-1:0] node3325;
	wire [8-1:0] node3326;
	wire [8-1:0] node3329;
	wire [8-1:0] node3330;
	wire [8-1:0] node3333;
	wire [8-1:0] node3336;
	wire [8-1:0] node3337;
	wire [8-1:0] node3338;
	wire [8-1:0] node3341;
	wire [8-1:0] node3342;
	wire [8-1:0] node3346;
	wire [8-1:0] node3347;
	wire [8-1:0] node3350;
	wire [8-1:0] node3353;
	wire [8-1:0] node3354;
	wire [8-1:0] node3355;
	wire [8-1:0] node3356;
	wire [8-1:0] node3358;
	wire [8-1:0] node3361;
	wire [8-1:0] node3363;
	wire [8-1:0] node3366;
	wire [8-1:0] node3367;
	wire [8-1:0] node3368;
	wire [8-1:0] node3371;
	wire [8-1:0] node3374;
	wire [8-1:0] node3375;
	wire [8-1:0] node3378;
	wire [8-1:0] node3381;
	wire [8-1:0] node3382;
	wire [8-1:0] node3383;
	wire [8-1:0] node3386;
	wire [8-1:0] node3388;
	wire [8-1:0] node3391;
	wire [8-1:0] node3392;
	wire [8-1:0] node3395;
	wire [8-1:0] node3396;
	wire [8-1:0] node3400;
	wire [8-1:0] node3401;
	wire [8-1:0] node3402;
	wire [8-1:0] node3403;
	wire [8-1:0] node3405;
	wire [8-1:0] node3407;
	wire [8-1:0] node3410;
	wire [8-1:0] node3411;
	wire [8-1:0] node3415;
	wire [8-1:0] node3416;
	wire [8-1:0] node3417;
	wire [8-1:0] node3418;
	wire [8-1:0] node3422;
	wire [8-1:0] node3423;
	wire [8-1:0] node3427;
	wire [8-1:0] node3428;
	wire [8-1:0] node3431;
	wire [8-1:0] node3434;
	wire [8-1:0] node3435;
	wire [8-1:0] node3436;
	wire [8-1:0] node3438;
	wire [8-1:0] node3439;
	wire [8-1:0] node3443;
	wire [8-1:0] node3444;
	wire [8-1:0] node3447;
	wire [8-1:0] node3450;
	wire [8-1:0] node3451;
	wire [8-1:0] node3452;
	wire [8-1:0] node3454;
	wire [8-1:0] node3457;
	wire [8-1:0] node3460;
	wire [8-1:0] node3461;
	wire [8-1:0] node3464;
	wire [8-1:0] node3467;
	wire [8-1:0] node3468;
	wire [8-1:0] node3469;
	wire [8-1:0] node3470;
	wire [8-1:0] node3473;
	wire [8-1:0] node3474;
	wire [8-1:0] node3475;
	wire [8-1:0] node3478;
	wire [8-1:0] node3481;
	wire [8-1:0] node3482;
	wire [8-1:0] node3483;
	wire [8-1:0] node3487;
	wire [8-1:0] node3490;
	wire [8-1:0] node3491;
	wire [8-1:0] node3492;
	wire [8-1:0] node3495;
	wire [8-1:0] node3498;
	wire [8-1:0] node3499;
	wire [8-1:0] node3501;
	wire [8-1:0] node3505;
	wire [8-1:0] node3506;
	wire [8-1:0] node3507;
	wire [8-1:0] node3510;
	wire [8-1:0] node3511;
	wire [8-1:0] node3512;
	wire [8-1:0] node3513;
	wire [8-1:0] node3517;
	wire [8-1:0] node3520;
	wire [8-1:0] node3521;
	wire [8-1:0] node3525;
	wire [8-1:0] node3526;
	wire [8-1:0] node3528;
	wire [8-1:0] node3529;
	wire [8-1:0] node3532;
	wire [8-1:0] node3535;
	wire [8-1:0] node3536;
	wire [8-1:0] node3540;
	wire [8-1:0] node3541;
	wire [8-1:0] node3542;
	wire [8-1:0] node3543;
	wire [8-1:0] node3544;
	wire [8-1:0] node3546;
	wire [8-1:0] node3547;
	wire [8-1:0] node3551;
	wire [8-1:0] node3552;
	wire [8-1:0] node3555;
	wire [8-1:0] node3556;
	wire [8-1:0] node3560;
	wire [8-1:0] node3561;
	wire [8-1:0] node3562;
	wire [8-1:0] node3564;
	wire [8-1:0] node3565;
	wire [8-1:0] node3568;
	wire [8-1:0] node3571;
	wire [8-1:0] node3572;
	wire [8-1:0] node3574;
	wire [8-1:0] node3578;
	wire [8-1:0] node3579;
	wire [8-1:0] node3581;
	wire [8-1:0] node3583;
	wire [8-1:0] node3586;
	wire [8-1:0] node3587;
	wire [8-1:0] node3589;
	wire [8-1:0] node3592;
	wire [8-1:0] node3594;
	wire [8-1:0] node3597;
	wire [8-1:0] node3598;
	wire [8-1:0] node3599;
	wire [8-1:0] node3600;
	wire [8-1:0] node3602;
	wire [8-1:0] node3605;
	wire [8-1:0] node3606;
	wire [8-1:0] node3609;
	wire [8-1:0] node3610;
	wire [8-1:0] node3613;
	wire [8-1:0] node3616;
	wire [8-1:0] node3617;
	wire [8-1:0] node3619;
	wire [8-1:0] node3622;
	wire [8-1:0] node3624;
	wire [8-1:0] node3627;
	wire [8-1:0] node3628;
	wire [8-1:0] node3630;
	wire [8-1:0] node3631;
	wire [8-1:0] node3634;
	wire [8-1:0] node3637;
	wire [8-1:0] node3638;
	wire [8-1:0] node3639;
	wire [8-1:0] node3643;
	wire [8-1:0] node3644;
	wire [8-1:0] node3645;
	wire [8-1:0] node3650;
	wire [8-1:0] node3651;
	wire [8-1:0] node3652;
	wire [8-1:0] node3654;
	wire [8-1:0] node3655;
	wire [8-1:0] node3659;
	wire [8-1:0] node3660;
	wire [8-1:0] node3661;
	wire [8-1:0] node3662;
	wire [8-1:0] node3665;
	wire [8-1:0] node3666;
	wire [8-1:0] node3670;
	wire [8-1:0] node3673;
	wire [8-1:0] node3674;
	wire [8-1:0] node3676;
	wire [8-1:0] node3678;
	wire [8-1:0] node3681;
	wire [8-1:0] node3682;
	wire [8-1:0] node3685;
	wire [8-1:0] node3688;
	wire [8-1:0] node3689;
	wire [8-1:0] node3690;
	wire [8-1:0] node3691;
	wire [8-1:0] node3695;
	wire [8-1:0] node3696;
	wire [8-1:0] node3697;
	wire [8-1:0] node3700;
	wire [8-1:0] node3704;
	wire [8-1:0] node3705;
	wire [8-1:0] node3706;
	wire [8-1:0] node3707;
	wire [8-1:0] node3710;
	wire [8-1:0] node3711;
	wire [8-1:0] node3715;
	wire [8-1:0] node3716;
	wire [8-1:0] node3720;
	wire [8-1:0] node3721;
	wire [8-1:0] node3722;
	wire [8-1:0] node3723;
	wire [8-1:0] node3727;
	wire [8-1:0] node3730;
	wire [8-1:0] node3731;
	wire [8-1:0] node3732;
	wire [8-1:0] node3736;
	wire [8-1:0] node3739;
	wire [8-1:0] node3740;
	wire [8-1:0] node3741;
	wire [8-1:0] node3742;
	wire [8-1:0] node3743;
	wire [8-1:0] node3744;
	wire [8-1:0] node3745;
	wire [8-1:0] node3746;
	wire [8-1:0] node3748;
	wire [8-1:0] node3751;
	wire [8-1:0] node3754;
	wire [8-1:0] node3756;
	wire [8-1:0] node3757;
	wire [8-1:0] node3761;
	wire [8-1:0] node3762;
	wire [8-1:0] node3763;
	wire [8-1:0] node3766;
	wire [8-1:0] node3768;
	wire [8-1:0] node3771;
	wire [8-1:0] node3772;
	wire [8-1:0] node3775;
	wire [8-1:0] node3776;
	wire [8-1:0] node3780;
	wire [8-1:0] node3781;
	wire [8-1:0] node3782;
	wire [8-1:0] node3784;
	wire [8-1:0] node3787;
	wire [8-1:0] node3789;
	wire [8-1:0] node3792;
	wire [8-1:0] node3793;
	wire [8-1:0] node3794;
	wire [8-1:0] node3797;
	wire [8-1:0] node3800;
	wire [8-1:0] node3801;
	wire [8-1:0] node3804;
	wire [8-1:0] node3807;
	wire [8-1:0] node3808;
	wire [8-1:0] node3809;
	wire [8-1:0] node3810;
	wire [8-1:0] node3811;
	wire [8-1:0] node3813;
	wire [8-1:0] node3817;
	wire [8-1:0] node3818;
	wire [8-1:0] node3821;
	wire [8-1:0] node3822;
	wire [8-1:0] node3826;
	wire [8-1:0] node3827;
	wire [8-1:0] node3829;
	wire [8-1:0] node3831;
	wire [8-1:0] node3834;
	wire [8-1:0] node3835;
	wire [8-1:0] node3837;
	wire [8-1:0] node3840;
	wire [8-1:0] node3843;
	wire [8-1:0] node3844;
	wire [8-1:0] node3845;
	wire [8-1:0] node3846;
	wire [8-1:0] node3850;
	wire [8-1:0] node3853;
	wire [8-1:0] node3854;
	wire [8-1:0] node3855;
	wire [8-1:0] node3859;
	wire [8-1:0] node3860;
	wire [8-1:0] node3863;
	wire [8-1:0] node3864;
	wire [8-1:0] node3867;
	wire [8-1:0] node3870;
	wire [8-1:0] node3871;
	wire [8-1:0] node3872;
	wire [8-1:0] node3875;
	wire [8-1:0] node3876;
	wire [8-1:0] node3877;
	wire [8-1:0] node3880;
	wire [8-1:0] node3883;
	wire [8-1:0] node3884;
	wire [8-1:0] node3887;
	wire [8-1:0] node3890;
	wire [8-1:0] node3891;
	wire [8-1:0] node3894;
	wire [8-1:0] node3895;
	wire [8-1:0] node3898;
	wire [8-1:0] node3901;
	wire [8-1:0] node3902;
	wire [8-1:0] node3903;
	wire [8-1:0] node3904;
	wire [8-1:0] node3905;
	wire [8-1:0] node3906;
	wire [8-1:0] node3907;
	wire [8-1:0] node3910;
	wire [8-1:0] node3913;
	wire [8-1:0] node3914;
	wire [8-1:0] node3917;
	wire [8-1:0] node3920;
	wire [8-1:0] node3921;
	wire [8-1:0] node3922;
	wire [8-1:0] node3925;
	wire [8-1:0] node3928;
	wire [8-1:0] node3929;
	wire [8-1:0] node3932;
	wire [8-1:0] node3935;
	wire [8-1:0] node3938;
	wire [8-1:0] node3939;
	wire [8-1:0] node3940;
	wire [8-1:0] node3941;
	wire [8-1:0] node3942;
	wire [8-1:0] node3943;
	wire [8-1:0] node3946;
	wire [8-1:0] node3949;
	wire [8-1:0] node3950;
	wire [8-1:0] node3953;
	wire [8-1:0] node3956;
	wire [8-1:0] node3957;
	wire [8-1:0] node3958;
	wire [8-1:0] node3961;
	wire [8-1:0] node3964;
	wire [8-1:0] node3965;
	wire [8-1:0] node3968;
	wire [8-1:0] node3971;
	wire [8-1:0] node3974;
	wire [8-1:0] node3975;
	wire [8-1:0] node3976;
	wire [8-1:0] node3977;
	wire [8-1:0] node3979;
	wire [8-1:0] node3982;
	wire [8-1:0] node3983;
	wire [8-1:0] node3987;
	wire [8-1:0] node3988;
	wire [8-1:0] node3989;
	wire [8-1:0] node3994;
	wire [8-1:0] node3997;
	wire [8-1:0] node3998;
	wire [8-1:0] node3999;
	wire [8-1:0] node4000;
	wire [8-1:0] node4001;
	wire [8-1:0] node4002;
	wire [8-1:0] node4005;
	wire [8-1:0] node4008;
	wire [8-1:0] node4009;
	wire [8-1:0] node4012;
	wire [8-1:0] node4015;
	wire [8-1:0] node4016;
	wire [8-1:0] node4017;
	wire [8-1:0] node4020;
	wire [8-1:0] node4023;
	wire [8-1:0] node4024;
	wire [8-1:0] node4027;
	wire [8-1:0] node4030;
	wire [8-1:0] node4031;
	wire [8-1:0] node4032;
	wire [8-1:0] node4033;
	wire [8-1:0] node4036;
	wire [8-1:0] node4039;
	wire [8-1:0] node4040;
	wire [8-1:0] node4043;
	wire [8-1:0] node4046;
	wire [8-1:0] node4047;
	wire [8-1:0] node4049;
	wire [8-1:0] node4052;
	wire [8-1:0] node4053;
	wire [8-1:0] node4056;
	wire [8-1:0] node4059;
	wire [8-1:0] node4062;
	wire [8-1:0] node4063;
	wire [8-1:0] node4064;
	wire [8-1:0] node4065;
	wire [8-1:0] node4066;
	wire [8-1:0] node4067;
	wire [8-1:0] node4068;
	wire [8-1:0] node4069;
	wire [8-1:0] node4070;
	wire [8-1:0] node4071;
	wire [8-1:0] node4072;
	wire [8-1:0] node4073;
	wire [8-1:0] node4078;
	wire [8-1:0] node4079;
	wire [8-1:0] node4083;
	wire [8-1:0] node4084;
	wire [8-1:0] node4086;
	wire [8-1:0] node4087;
	wire [8-1:0] node4090;
	wire [8-1:0] node4093;
	wire [8-1:0] node4094;
	wire [8-1:0] node4095;
	wire [8-1:0] node4098;
	wire [8-1:0] node4101;
	wire [8-1:0] node4102;
	wire [8-1:0] node4103;
	wire [8-1:0] node4106;
	wire [8-1:0] node4110;
	wire [8-1:0] node4111;
	wire [8-1:0] node4112;
	wire [8-1:0] node4113;
	wire [8-1:0] node4116;
	wire [8-1:0] node4118;
	wire [8-1:0] node4121;
	wire [8-1:0] node4122;
	wire [8-1:0] node4123;
	wire [8-1:0] node4127;
	wire [8-1:0] node4130;
	wire [8-1:0] node4131;
	wire [8-1:0] node4132;
	wire [8-1:0] node4135;
	wire [8-1:0] node4137;
	wire [8-1:0] node4140;
	wire [8-1:0] node4141;
	wire [8-1:0] node4144;
	wire [8-1:0] node4145;
	wire [8-1:0] node4146;
	wire [8-1:0] node4150;
	wire [8-1:0] node4151;
	wire [8-1:0] node4154;
	wire [8-1:0] node4157;
	wire [8-1:0] node4158;
	wire [8-1:0] node4160;
	wire [8-1:0] node4162;
	wire [8-1:0] node4165;
	wire [8-1:0] node4166;
	wire [8-1:0] node4168;
	wire [8-1:0] node4171;
	wire [8-1:0] node4173;
	wire [8-1:0] node4174;
	wire [8-1:0] node4177;
	wire [8-1:0] node4180;
	wire [8-1:0] node4181;
	wire [8-1:0] node4182;
	wire [8-1:0] node4183;
	wire [8-1:0] node4184;
	wire [8-1:0] node4185;
	wire [8-1:0] node4188;
	wire [8-1:0] node4192;
	wire [8-1:0] node4193;
	wire [8-1:0] node4197;
	wire [8-1:0] node4198;
	wire [8-1:0] node4199;
	wire [8-1:0] node4204;
	wire [8-1:0] node4205;
	wire [8-1:0] node4206;
	wire [8-1:0] node4207;
	wire [8-1:0] node4208;
	wire [8-1:0] node4211;
	wire [8-1:0] node4213;
	wire [8-1:0] node4216;
	wire [8-1:0] node4217;
	wire [8-1:0] node4218;
	wire [8-1:0] node4219;
	wire [8-1:0] node4223;
	wire [8-1:0] node4224;
	wire [8-1:0] node4228;
	wire [8-1:0] node4230;
	wire [8-1:0] node4233;
	wire [8-1:0] node4234;
	wire [8-1:0] node4235;
	wire [8-1:0] node4238;
	wire [8-1:0] node4239;
	wire [8-1:0] node4243;
	wire [8-1:0] node4244;
	wire [8-1:0] node4245;
	wire [8-1:0] node4248;
	wire [8-1:0] node4252;
	wire [8-1:0] node4253;
	wire [8-1:0] node4254;
	wire [8-1:0] node4255;
	wire [8-1:0] node4256;
	wire [8-1:0] node4260;
	wire [8-1:0] node4262;
	wire [8-1:0] node4263;
	wire [8-1:0] node4266;
	wire [8-1:0] node4269;
	wire [8-1:0] node4270;
	wire [8-1:0] node4271;
	wire [8-1:0] node4274;
	wire [8-1:0] node4277;
	wire [8-1:0] node4278;
	wire [8-1:0] node4281;
	wire [8-1:0] node4284;
	wire [8-1:0] node4285;
	wire [8-1:0] node4286;
	wire [8-1:0] node4289;
	wire [8-1:0] node4291;
	wire [8-1:0] node4294;
	wire [8-1:0] node4295;
	wire [8-1:0] node4299;
	wire [8-1:0] node4300;
	wire [8-1:0] node4301;
	wire [8-1:0] node4302;
	wire [8-1:0] node4303;
	wire [8-1:0] node4304;
	wire [8-1:0] node4305;
	wire [8-1:0] node4308;
	wire [8-1:0] node4311;
	wire [8-1:0] node4312;
	wire [8-1:0] node4314;
	wire [8-1:0] node4316;
	wire [8-1:0] node4319;
	wire [8-1:0] node4320;
	wire [8-1:0] node4321;
	wire [8-1:0] node4326;
	wire [8-1:0] node4327;
	wire [8-1:0] node4328;
	wire [8-1:0] node4331;
	wire [8-1:0] node4333;
	wire [8-1:0] node4336;
	wire [8-1:0] node4337;
	wire [8-1:0] node4338;
	wire [8-1:0] node4342;
	wire [8-1:0] node4343;
	wire [8-1:0] node4346;
	wire [8-1:0] node4347;
	wire [8-1:0] node4351;
	wire [8-1:0] node4352;
	wire [8-1:0] node4353;
	wire [8-1:0] node4354;
	wire [8-1:0] node4356;
	wire [8-1:0] node4359;
	wire [8-1:0] node4360;
	wire [8-1:0] node4364;
	wire [8-1:0] node4366;
	wire [8-1:0] node4367;
	wire [8-1:0] node4368;
	wire [8-1:0] node4371;
	wire [8-1:0] node4374;
	wire [8-1:0] node4375;
	wire [8-1:0] node4379;
	wire [8-1:0] node4380;
	wire [8-1:0] node4381;
	wire [8-1:0] node4382;
	wire [8-1:0] node4383;
	wire [8-1:0] node4387;
	wire [8-1:0] node4388;
	wire [8-1:0] node4392;
	wire [8-1:0] node4393;
	wire [8-1:0] node4394;
	wire [8-1:0] node4398;
	wire [8-1:0] node4401;
	wire [8-1:0] node4402;
	wire [8-1:0] node4403;
	wire [8-1:0] node4406;
	wire [8-1:0] node4409;
	wire [8-1:0] node4412;
	wire [8-1:0] node4413;
	wire [8-1:0] node4414;
	wire [8-1:0] node4415;
	wire [8-1:0] node4416;
	wire [8-1:0] node4419;
	wire [8-1:0] node4422;
	wire [8-1:0] node4423;
	wire [8-1:0] node4424;
	wire [8-1:0] node4428;
	wire [8-1:0] node4429;
	wire [8-1:0] node4433;
	wire [8-1:0] node4434;
	wire [8-1:0] node4435;
	wire [8-1:0] node4437;
	wire [8-1:0] node4440;
	wire [8-1:0] node4442;
	wire [8-1:0] node4445;
	wire [8-1:0] node4447;
	wire [8-1:0] node4448;
	wire [8-1:0] node4451;
	wire [8-1:0] node4454;
	wire [8-1:0] node4455;
	wire [8-1:0] node4456;
	wire [8-1:0] node4457;
	wire [8-1:0] node4458;
	wire [8-1:0] node4460;
	wire [8-1:0] node4463;
	wire [8-1:0] node4466;
	wire [8-1:0] node4469;
	wire [8-1:0] node4470;
	wire [8-1:0] node4471;
	wire [8-1:0] node4475;
	wire [8-1:0] node4477;
	wire [8-1:0] node4478;
	wire [8-1:0] node4482;
	wire [8-1:0] node4483;
	wire [8-1:0] node4484;
	wire [8-1:0] node4486;
	wire [8-1:0] node4490;
	wire [8-1:0] node4491;
	wire [8-1:0] node4492;
	wire [8-1:0] node4494;
	wire [8-1:0] node4497;
	wire [8-1:0] node4498;
	wire [8-1:0] node4501;
	wire [8-1:0] node4504;
	wire [8-1:0] node4505;
	wire [8-1:0] node4508;
	wire [8-1:0] node4511;
	wire [8-1:0] node4512;
	wire [8-1:0] node4513;
	wire [8-1:0] node4514;
	wire [8-1:0] node4515;
	wire [8-1:0] node4516;
	wire [8-1:0] node4517;
	wire [8-1:0] node4521;
	wire [8-1:0] node4522;
	wire [8-1:0] node4526;
	wire [8-1:0] node4527;
	wire [8-1:0] node4531;
	wire [8-1:0] node4532;
	wire [8-1:0] node4533;
	wire [8-1:0] node4536;
	wire [8-1:0] node4537;
	wire [8-1:0] node4541;
	wire [8-1:0] node4542;
	wire [8-1:0] node4546;
	wire [8-1:0] node4547;
	wire [8-1:0] node4548;
	wire [8-1:0] node4549;
	wire [8-1:0] node4550;
	wire [8-1:0] node4551;
	wire [8-1:0] node4554;
	wire [8-1:0] node4558;
	wire [8-1:0] node4559;
	wire [8-1:0] node4560;
	wire [8-1:0] node4563;
	wire [8-1:0] node4566;
	wire [8-1:0] node4567;
	wire [8-1:0] node4571;
	wire [8-1:0] node4572;
	wire [8-1:0] node4574;
	wire [8-1:0] node4575;
	wire [8-1:0] node4579;
	wire [8-1:0] node4580;
	wire [8-1:0] node4581;
	wire [8-1:0] node4585;
	wire [8-1:0] node4588;
	wire [8-1:0] node4589;
	wire [8-1:0] node4590;
	wire [8-1:0] node4591;
	wire [8-1:0] node4592;
	wire [8-1:0] node4596;
	wire [8-1:0] node4597;
	wire [8-1:0] node4601;
	wire [8-1:0] node4602;
	wire [8-1:0] node4605;
	wire [8-1:0] node4608;
	wire [8-1:0] node4609;
	wire [8-1:0] node4610;
	wire [8-1:0] node4612;
	wire [8-1:0] node4615;
	wire [8-1:0] node4616;
	wire [8-1:0] node4619;
	wire [8-1:0] node4622;
	wire [8-1:0] node4623;
	wire [8-1:0] node4626;
	wire [8-1:0] node4628;
	wire [8-1:0] node4631;
	wire [8-1:0] node4632;
	wire [8-1:0] node4633;
	wire [8-1:0] node4634;
	wire [8-1:0] node4635;
	wire [8-1:0] node4636;
	wire [8-1:0] node4638;
	wire [8-1:0] node4641;
	wire [8-1:0] node4642;
	wire [8-1:0] node4645;
	wire [8-1:0] node4648;
	wire [8-1:0] node4649;
	wire [8-1:0] node4650;
	wire [8-1:0] node4654;
	wire [8-1:0] node4656;
	wire [8-1:0] node4659;
	wire [8-1:0] node4660;
	wire [8-1:0] node4661;
	wire [8-1:0] node4663;
	wire [8-1:0] node4666;
	wire [8-1:0] node4669;
	wire [8-1:0] node4670;
	wire [8-1:0] node4673;
	wire [8-1:0] node4674;
	wire [8-1:0] node4677;
	wire [8-1:0] node4680;
	wire [8-1:0] node4681;
	wire [8-1:0] node4682;
	wire [8-1:0] node4683;
	wire [8-1:0] node4684;
	wire [8-1:0] node4687;
	wire [8-1:0] node4690;
	wire [8-1:0] node4692;
	wire [8-1:0] node4695;
	wire [8-1:0] node4696;
	wire [8-1:0] node4698;
	wire [8-1:0] node4701;
	wire [8-1:0] node4702;
	wire [8-1:0] node4705;
	wire [8-1:0] node4708;
	wire [8-1:0] node4709;
	wire [8-1:0] node4710;
	wire [8-1:0] node4711;
	wire [8-1:0] node4715;
	wire [8-1:0] node4717;
	wire [8-1:0] node4720;
	wire [8-1:0] node4721;
	wire [8-1:0] node4723;
	wire [8-1:0] node4727;
	wire [8-1:0] node4728;
	wire [8-1:0] node4729;
	wire [8-1:0] node4730;
	wire [8-1:0] node4731;
	wire [8-1:0] node4736;
	wire [8-1:0] node4737;
	wire [8-1:0] node4738;
	wire [8-1:0] node4741;
	wire [8-1:0] node4744;
	wire [8-1:0] node4747;
	wire [8-1:0] node4748;
	wire [8-1:0] node4749;
	wire [8-1:0] node4752;
	wire [8-1:0] node4755;
	wire [8-1:0] node4758;
	wire [8-1:0] node4759;
	wire [8-1:0] node4760;
	wire [8-1:0] node4761;
	wire [8-1:0] node4762;
	wire [8-1:0] node4763;
	wire [8-1:0] node4764;
	wire [8-1:0] node4766;
	wire [8-1:0] node4769;
	wire [8-1:0] node4771;
	wire [8-1:0] node4774;
	wire [8-1:0] node4775;
	wire [8-1:0] node4776;
	wire [8-1:0] node4779;
	wire [8-1:0] node4782;
	wire [8-1:0] node4784;
	wire [8-1:0] node4786;
	wire [8-1:0] node4789;
	wire [8-1:0] node4790;
	wire [8-1:0] node4791;
	wire [8-1:0] node4793;
	wire [8-1:0] node4797;
	wire [8-1:0] node4798;
	wire [8-1:0] node4799;
	wire [8-1:0] node4800;
	wire [8-1:0] node4804;
	wire [8-1:0] node4806;
	wire [8-1:0] node4809;
	wire [8-1:0] node4810;
	wire [8-1:0] node4811;
	wire [8-1:0] node4815;
	wire [8-1:0] node4818;
	wire [8-1:0] node4819;
	wire [8-1:0] node4820;
	wire [8-1:0] node4821;
	wire [8-1:0] node4822;
	wire [8-1:0] node4825;
	wire [8-1:0] node4828;
	wire [8-1:0] node4829;
	wire [8-1:0] node4830;
	wire [8-1:0] node4834;
	wire [8-1:0] node4835;
	wire [8-1:0] node4838;
	wire [8-1:0] node4839;
	wire [8-1:0] node4843;
	wire [8-1:0] node4844;
	wire [8-1:0] node4845;
	wire [8-1:0] node4848;
	wire [8-1:0] node4851;
	wire [8-1:0] node4852;
	wire [8-1:0] node4853;
	wire [8-1:0] node4855;
	wire [8-1:0] node4859;
	wire [8-1:0] node4861;
	wire [8-1:0] node4862;
	wire [8-1:0] node4866;
	wire [8-1:0] node4867;
	wire [8-1:0] node4868;
	wire [8-1:0] node4869;
	wire [8-1:0] node4870;
	wire [8-1:0] node4872;
	wire [8-1:0] node4876;
	wire [8-1:0] node4877;
	wire [8-1:0] node4879;
	wire [8-1:0] node4882;
	wire [8-1:0] node4885;
	wire [8-1:0] node4886;
	wire [8-1:0] node4887;
	wire [8-1:0] node4891;
	wire [8-1:0] node4892;
	wire [8-1:0] node4893;
	wire [8-1:0] node4896;
	wire [8-1:0] node4899;
	wire [8-1:0] node4900;
	wire [8-1:0] node4903;
	wire [8-1:0] node4906;
	wire [8-1:0] node4907;
	wire [8-1:0] node4908;
	wire [8-1:0] node4909;
	wire [8-1:0] node4911;
	wire [8-1:0] node4914;
	wire [8-1:0] node4917;
	wire [8-1:0] node4920;
	wire [8-1:0] node4921;
	wire [8-1:0] node4922;
	wire [8-1:0] node4926;
	wire [8-1:0] node4927;
	wire [8-1:0] node4931;
	wire [8-1:0] node4932;
	wire [8-1:0] node4933;
	wire [8-1:0] node4934;
	wire [8-1:0] node4935;
	wire [8-1:0] node4936;
	wire [8-1:0] node4940;
	wire [8-1:0] node4942;
	wire [8-1:0] node4945;
	wire [8-1:0] node4946;
	wire [8-1:0] node4947;
	wire [8-1:0] node4949;
	wire [8-1:0] node4952;
	wire [8-1:0] node4954;
	wire [8-1:0] node4957;
	wire [8-1:0] node4958;
	wire [8-1:0] node4960;
	wire [8-1:0] node4963;
	wire [8-1:0] node4964;
	wire [8-1:0] node4967;
	wire [8-1:0] node4968;
	wire [8-1:0] node4972;
	wire [8-1:0] node4973;
	wire [8-1:0] node4974;
	wire [8-1:0] node4976;
	wire [8-1:0] node4979;
	wire [8-1:0] node4980;
	wire [8-1:0] node4984;
	wire [8-1:0] node4985;
	wire [8-1:0] node4986;
	wire [8-1:0] node4988;
	wire [8-1:0] node4990;
	wire [8-1:0] node4993;
	wire [8-1:0] node4994;
	wire [8-1:0] node4996;
	wire [8-1:0] node5000;
	wire [8-1:0] node5001;
	wire [8-1:0] node5002;
	wire [8-1:0] node5005;
	wire [8-1:0] node5006;
	wire [8-1:0] node5010;
	wire [8-1:0] node5013;
	wire [8-1:0] node5014;
	wire [8-1:0] node5015;
	wire [8-1:0] node5016;
	wire [8-1:0] node5017;
	wire [8-1:0] node5018;
	wire [8-1:0] node5022;
	wire [8-1:0] node5023;
	wire [8-1:0] node5026;
	wire [8-1:0] node5029;
	wire [8-1:0] node5031;
	wire [8-1:0] node5032;
	wire [8-1:0] node5036;
	wire [8-1:0] node5037;
	wire [8-1:0] node5038;
	wire [8-1:0] node5039;
	wire [8-1:0] node5042;
	wire [8-1:0] node5043;
	wire [8-1:0] node5047;
	wire [8-1:0] node5049;
	wire [8-1:0] node5050;
	wire [8-1:0] node5053;
	wire [8-1:0] node5056;
	wire [8-1:0] node5057;
	wire [8-1:0] node5061;
	wire [8-1:0] node5062;
	wire [8-1:0] node5063;
	wire [8-1:0] node5064;
	wire [8-1:0] node5065;
	wire [8-1:0] node5069;
	wire [8-1:0] node5070;
	wire [8-1:0] node5074;
	wire [8-1:0] node5075;
	wire [8-1:0] node5076;
	wire [8-1:0] node5079;
	wire [8-1:0] node5081;
	wire [8-1:0] node5084;
	wire [8-1:0] node5085;
	wire [8-1:0] node5088;
	wire [8-1:0] node5089;
	wire [8-1:0] node5093;
	wire [8-1:0] node5094;
	wire [8-1:0] node5095;
	wire [8-1:0] node5097;
	wire [8-1:0] node5100;
	wire [8-1:0] node5101;
	wire [8-1:0] node5102;
	wire [8-1:0] node5106;
	wire [8-1:0] node5107;
	wire [8-1:0] node5111;
	wire [8-1:0] node5112;
	wire [8-1:0] node5113;
	wire [8-1:0] node5114;
	wire [8-1:0] node5118;
	wire [8-1:0] node5119;
	wire [8-1:0] node5122;
	wire [8-1:0] node5125;
	wire [8-1:0] node5128;
	wire [8-1:0] node5129;
	wire [8-1:0] node5130;
	wire [8-1:0] node5131;
	wire [8-1:0] node5132;
	wire [8-1:0] node5133;
	wire [8-1:0] node5134;
	wire [8-1:0] node5135;
	wire [8-1:0] node5139;
	wire [8-1:0] node5140;
	wire [8-1:0] node5144;
	wire [8-1:0] node5145;
	wire [8-1:0] node5149;
	wire [8-1:0] node5150;
	wire [8-1:0] node5151;
	wire [8-1:0] node5152;
	wire [8-1:0] node5157;
	wire [8-1:0] node5158;
	wire [8-1:0] node5162;
	wire [8-1:0] node5163;
	wire [8-1:0] node5164;
	wire [8-1:0] node5165;
	wire [8-1:0] node5169;
	wire [8-1:0] node5170;
	wire [8-1:0] node5174;
	wire [8-1:0] node5175;
	wire [8-1:0] node5179;
	wire [8-1:0] node5180;
	wire [8-1:0] node5181;
	wire [8-1:0] node5182;
	wire [8-1:0] node5183;
	wire [8-1:0] node5186;
	wire [8-1:0] node5189;
	wire [8-1:0] node5190;
	wire [8-1:0] node5194;
	wire [8-1:0] node5195;
	wire [8-1:0] node5196;
	wire [8-1:0] node5197;
	wire [8-1:0] node5200;
	wire [8-1:0] node5203;
	wire [8-1:0] node5204;
	wire [8-1:0] node5207;
	wire [8-1:0] node5209;
	wire [8-1:0] node5212;
	wire [8-1:0] node5213;
	wire [8-1:0] node5214;
	wire [8-1:0] node5216;
	wire [8-1:0] node5219;
	wire [8-1:0] node5222;
	wire [8-1:0] node5225;
	wire [8-1:0] node5226;
	wire [8-1:0] node5227;
	wire [8-1:0] node5228;
	wire [8-1:0] node5231;
	wire [8-1:0] node5232;
	wire [8-1:0] node5233;
	wire [8-1:0] node5236;
	wire [8-1:0] node5239;
	wire [8-1:0] node5240;
	wire [8-1:0] node5243;
	wire [8-1:0] node5246;
	wire [8-1:0] node5247;
	wire [8-1:0] node5248;
	wire [8-1:0] node5251;
	wire [8-1:0] node5252;
	wire [8-1:0] node5256;
	wire [8-1:0] node5257;
	wire [8-1:0] node5260;
	wire [8-1:0] node5261;
	wire [8-1:0] node5265;
	wire [8-1:0] node5266;
	wire [8-1:0] node5267;
	wire [8-1:0] node5268;
	wire [8-1:0] node5272;
	wire [8-1:0] node5273;
	wire [8-1:0] node5276;
	wire [8-1:0] node5279;
	wire [8-1:0] node5280;
	wire [8-1:0] node5281;
	wire [8-1:0] node5283;
	wire [8-1:0] node5286;
	wire [8-1:0] node5287;
	wire [8-1:0] node5291;
	wire [8-1:0] node5292;
	wire [8-1:0] node5294;
	wire [8-1:0] node5297;
	wire [8-1:0] node5298;
	wire [8-1:0] node5301;
	wire [8-1:0] node5304;
	wire [8-1:0] node5305;
	wire [8-1:0] node5306;
	wire [8-1:0] node5307;
	wire [8-1:0] node5308;
	wire [8-1:0] node5309;
	wire [8-1:0] node5310;
	wire [8-1:0] node5313;
	wire [8-1:0] node5316;
	wire [8-1:0] node5317;
	wire [8-1:0] node5318;
	wire [8-1:0] node5321;
	wire [8-1:0] node5325;
	wire [8-1:0] node5326;
	wire [8-1:0] node5327;
	wire [8-1:0] node5329;
	wire [8-1:0] node5332;
	wire [8-1:0] node5333;
	wire [8-1:0] node5336;
	wire [8-1:0] node5339;
	wire [8-1:0] node5341;
	wire [8-1:0] node5344;
	wire [8-1:0] node5345;
	wire [8-1:0] node5346;
	wire [8-1:0] node5347;
	wire [8-1:0] node5350;
	wire [8-1:0] node5353;
	wire [8-1:0] node5354;
	wire [8-1:0] node5358;
	wire [8-1:0] node5359;
	wire [8-1:0] node5360;
	wire [8-1:0] node5363;
	wire [8-1:0] node5366;
	wire [8-1:0] node5367;
	wire [8-1:0] node5370;
	wire [8-1:0] node5373;
	wire [8-1:0] node5374;
	wire [8-1:0] node5376;
	wire [8-1:0] node5377;
	wire [8-1:0] node5380;
	wire [8-1:0] node5383;
	wire [8-1:0] node5384;
	wire [8-1:0] node5388;
	wire [8-1:0] node5389;
	wire [8-1:0] node5390;
	wire [8-1:0] node5391;
	wire [8-1:0] node5392;
	wire [8-1:0] node5394;
	wire [8-1:0] node5397;
	wire [8-1:0] node5399;
	wire [8-1:0] node5400;
	wire [8-1:0] node5404;
	wire [8-1:0] node5405;
	wire [8-1:0] node5407;
	wire [8-1:0] node5410;
	wire [8-1:0] node5413;
	wire [8-1:0] node5414;
	wire [8-1:0] node5415;
	wire [8-1:0] node5416;
	wire [8-1:0] node5419;
	wire [8-1:0] node5422;
	wire [8-1:0] node5423;
	wire [8-1:0] node5426;
	wire [8-1:0] node5427;
	wire [8-1:0] node5431;
	wire [8-1:0] node5432;
	wire [8-1:0] node5433;
	wire [8-1:0] node5435;
	wire [8-1:0] node5438;
	wire [8-1:0] node5439;
	wire [8-1:0] node5442;
	wire [8-1:0] node5445;
	wire [8-1:0] node5448;
	wire [8-1:0] node5449;
	wire [8-1:0] node5450;
	wire [8-1:0] node5451;
	wire [8-1:0] node5453;
	wire [8-1:0] node5454;
	wire [8-1:0] node5458;
	wire [8-1:0] node5459;
	wire [8-1:0] node5460;
	wire [8-1:0] node5465;
	wire [8-1:0] node5466;
	wire [8-1:0] node5467;
	wire [8-1:0] node5468;
	wire [8-1:0] node5472;
	wire [8-1:0] node5474;
	wire [8-1:0] node5477;
	wire [8-1:0] node5478;
	wire [8-1:0] node5479;
	wire [8-1:0] node5482;
	wire [8-1:0] node5485;
	wire [8-1:0] node5488;
	wire [8-1:0] node5489;
	wire [8-1:0] node5490;
	wire [8-1:0] node5493;
	wire [8-1:0] node5496;
	wire [8-1:0] node5499;
	wire [8-1:0] node5500;
	wire [8-1:0] node5501;
	wire [8-1:0] node5502;
	wire [8-1:0] node5503;
	wire [8-1:0] node5504;
	wire [8-1:0] node5505;
	wire [8-1:0] node5506;
	wire [8-1:0] node5507;
	wire [8-1:0] node5508;
	wire [8-1:0] node5512;
	wire [8-1:0] node5513;
	wire [8-1:0] node5517;
	wire [8-1:0] node5518;
	wire [8-1:0] node5522;
	wire [8-1:0] node5523;
	wire [8-1:0] node5524;
	wire [8-1:0] node5525;
	wire [8-1:0] node5529;
	wire [8-1:0] node5531;
	wire [8-1:0] node5532;
	wire [8-1:0] node5536;
	wire [8-1:0] node5537;
	wire [8-1:0] node5541;
	wire [8-1:0] node5542;
	wire [8-1:0] node5543;
	wire [8-1:0] node5544;
	wire [8-1:0] node5548;
	wire [8-1:0] node5549;
	wire [8-1:0] node5553;
	wire [8-1:0] node5554;
	wire [8-1:0] node5558;
	wire [8-1:0] node5559;
	wire [8-1:0] node5560;
	wire [8-1:0] node5561;
	wire [8-1:0] node5562;
	wire [8-1:0] node5563;
	wire [8-1:0] node5567;
	wire [8-1:0] node5568;
	wire [8-1:0] node5572;
	wire [8-1:0] node5573;
	wire [8-1:0] node5577;
	wire [8-1:0] node5578;
	wire [8-1:0] node5579;
	wire [8-1:0] node5580;
	wire [8-1:0] node5584;
	wire [8-1:0] node5585;
	wire [8-1:0] node5589;
	wire [8-1:0] node5590;
	wire [8-1:0] node5594;
	wire [8-1:0] node5595;
	wire [8-1:0] node5596;
	wire [8-1:0] node5597;
	wire [8-1:0] node5601;
	wire [8-1:0] node5602;
	wire [8-1:0] node5606;
	wire [8-1:0] node5607;
	wire [8-1:0] node5611;
	wire [8-1:0] node5612;
	wire [8-1:0] node5613;
	wire [8-1:0] node5614;
	wire [8-1:0] node5615;
	wire [8-1:0] node5616;
	wire [8-1:0] node5620;
	wire [8-1:0] node5621;
	wire [8-1:0] node5625;
	wire [8-1:0] node5626;
	wire [8-1:0] node5630;
	wire [8-1:0] node5631;
	wire [8-1:0] node5632;
	wire [8-1:0] node5633;
	wire [8-1:0] node5637;
	wire [8-1:0] node5638;
	wire [8-1:0] node5642;
	wire [8-1:0] node5643;
	wire [8-1:0] node5647;
	wire [8-1:0] node5648;
	wire [8-1:0] node5649;
	wire [8-1:0] node5650;
	wire [8-1:0] node5654;
	wire [8-1:0] node5655;
	wire [8-1:0] node5659;
	wire [8-1:0] node5660;
	wire [8-1:0] node5664;
	wire [8-1:0] node5665;
	wire [8-1:0] node5666;
	wire [8-1:0] node5667;
	wire [8-1:0] node5668;
	wire [8-1:0] node5669;
	wire [8-1:0] node5670;
	wire [8-1:0] node5671;
	wire [8-1:0] node5672;
	wire [8-1:0] node5676;
	wire [8-1:0] node5677;
	wire [8-1:0] node5680;
	wire [8-1:0] node5683;
	wire [8-1:0] node5685;
	wire [8-1:0] node5686;
	wire [8-1:0] node5689;
	wire [8-1:0] node5692;
	wire [8-1:0] node5693;
	wire [8-1:0] node5694;
	wire [8-1:0] node5697;
	wire [8-1:0] node5698;
	wire [8-1:0] node5702;
	wire [8-1:0] node5705;
	wire [8-1:0] node5706;
	wire [8-1:0] node5707;
	wire [8-1:0] node5708;
	wire [8-1:0] node5709;
	wire [8-1:0] node5713;
	wire [8-1:0] node5714;
	wire [8-1:0] node5717;
	wire [8-1:0] node5720;
	wire [8-1:0] node5721;
	wire [8-1:0] node5722;
	wire [8-1:0] node5725;
	wire [8-1:0] node5728;
	wire [8-1:0] node5730;
	wire [8-1:0] node5733;
	wire [8-1:0] node5734;
	wire [8-1:0] node5735;
	wire [8-1:0] node5736;
	wire [8-1:0] node5739;
	wire [8-1:0] node5743;
	wire [8-1:0] node5744;
	wire [8-1:0] node5747;
	wire [8-1:0] node5750;
	wire [8-1:0] node5751;
	wire [8-1:0] node5752;
	wire [8-1:0] node5753;
	wire [8-1:0] node5754;
	wire [8-1:0] node5756;
	wire [8-1:0] node5760;
	wire [8-1:0] node5761;
	wire [8-1:0] node5764;
	wire [8-1:0] node5765;
	wire [8-1:0] node5768;
	wire [8-1:0] node5771;
	wire [8-1:0] node5772;
	wire [8-1:0] node5773;
	wire [8-1:0] node5775;
	wire [8-1:0] node5778;
	wire [8-1:0] node5781;
	wire [8-1:0] node5782;
	wire [8-1:0] node5783;
	wire [8-1:0] node5787;
	wire [8-1:0] node5790;
	wire [8-1:0] node5791;
	wire [8-1:0] node5792;
	wire [8-1:0] node5793;
	wire [8-1:0] node5796;
	wire [8-1:0] node5797;
	wire [8-1:0] node5801;
	wire [8-1:0] node5802;
	wire [8-1:0] node5805;
	wire [8-1:0] node5808;
	wire [8-1:0] node5809;
	wire [8-1:0] node5810;
	wire [8-1:0] node5811;
	wire [8-1:0] node5814;
	wire [8-1:0] node5817;
	wire [8-1:0] node5820;
	wire [8-1:0] node5821;
	wire [8-1:0] node5822;
	wire [8-1:0] node5825;
	wire [8-1:0] node5829;
	wire [8-1:0] node5830;
	wire [8-1:0] node5831;
	wire [8-1:0] node5832;
	wire [8-1:0] node5833;
	wire [8-1:0] node5835;
	wire [8-1:0] node5837;
	wire [8-1:0] node5840;
	wire [8-1:0] node5841;
	wire [8-1:0] node5842;
	wire [8-1:0] node5845;
	wire [8-1:0] node5848;
	wire [8-1:0] node5850;
	wire [8-1:0] node5853;
	wire [8-1:0] node5854;
	wire [8-1:0] node5855;
	wire [8-1:0] node5857;
	wire [8-1:0] node5860;
	wire [8-1:0] node5863;
	wire [8-1:0] node5864;
	wire [8-1:0] node5865;
	wire [8-1:0] node5869;
	wire [8-1:0] node5871;
	wire [8-1:0] node5874;
	wire [8-1:0] node5875;
	wire [8-1:0] node5876;
	wire [8-1:0] node5878;
	wire [8-1:0] node5881;
	wire [8-1:0] node5882;
	wire [8-1:0] node5883;
	wire [8-1:0] node5887;
	wire [8-1:0] node5888;
	wire [8-1:0] node5892;
	wire [8-1:0] node5893;
	wire [8-1:0] node5894;
	wire [8-1:0] node5897;
	wire [8-1:0] node5900;
	wire [8-1:0] node5902;
	wire [8-1:0] node5903;
	wire [8-1:0] node5906;
	wire [8-1:0] node5909;
	wire [8-1:0] node5910;
	wire [8-1:0] node5911;
	wire [8-1:0] node5912;
	wire [8-1:0] node5913;
	wire [8-1:0] node5916;
	wire [8-1:0] node5919;
	wire [8-1:0] node5921;
	wire [8-1:0] node5924;
	wire [8-1:0] node5925;
	wire [8-1:0] node5926;
	wire [8-1:0] node5929;
	wire [8-1:0] node5932;
	wire [8-1:0] node5933;
	wire [8-1:0] node5936;
	wire [8-1:0] node5939;
	wire [8-1:0] node5940;
	wire [8-1:0] node5941;
	wire [8-1:0] node5942;
	wire [8-1:0] node5944;
	wire [8-1:0] node5947;
	wire [8-1:0] node5948;
	wire [8-1:0] node5951;
	wire [8-1:0] node5954;
	wire [8-1:0] node5955;
	wire [8-1:0] node5956;
	wire [8-1:0] node5959;
	wire [8-1:0] node5963;
	wire [8-1:0] node5964;
	wire [8-1:0] node5965;
	wire [8-1:0] node5967;
	wire [8-1:0] node5970;
	wire [8-1:0] node5971;
	wire [8-1:0] node5975;
	wire [8-1:0] node5976;
	wire [8-1:0] node5978;
	wire [8-1:0] node5981;
	wire [8-1:0] node5984;
	wire [8-1:0] node5985;
	wire [8-1:0] node5986;
	wire [8-1:0] node5987;
	wire [8-1:0] node5988;
	wire [8-1:0] node5989;
	wire [8-1:0] node5990;
	wire [8-1:0] node5993;
	wire [8-1:0] node5996;
	wire [8-1:0] node5997;
	wire [8-1:0] node6000;
	wire [8-1:0] node6003;
	wire [8-1:0] node6004;
	wire [8-1:0] node6005;
	wire [8-1:0] node6008;
	wire [8-1:0] node6011;
	wire [8-1:0] node6012;
	wire [8-1:0] node6015;
	wire [8-1:0] node6018;
	wire [8-1:0] node6019;
	wire [8-1:0] node6020;
	wire [8-1:0] node6022;
	wire [8-1:0] node6023;
	wire [8-1:0] node6026;
	wire [8-1:0] node6029;
	wire [8-1:0] node6032;
	wire [8-1:0] node6033;
	wire [8-1:0] node6034;
	wire [8-1:0] node6037;
	wire [8-1:0] node6040;
	wire [8-1:0] node6041;
	wire [8-1:0] node6044;
	wire [8-1:0] node6047;
	wire [8-1:0] node6048;
	wire [8-1:0] node6049;
	wire [8-1:0] node6050;
	wire [8-1:0] node6051;
	wire [8-1:0] node6054;
	wire [8-1:0] node6057;
	wire [8-1:0] node6058;
	wire [8-1:0] node6061;
	wire [8-1:0] node6064;
	wire [8-1:0] node6066;
	wire [8-1:0] node6067;
	wire [8-1:0] node6070;
	wire [8-1:0] node6073;
	wire [8-1:0] node6074;
	wire [8-1:0] node6075;
	wire [8-1:0] node6076;
	wire [8-1:0] node6079;
	wire [8-1:0] node6082;
	wire [8-1:0] node6084;
	wire [8-1:0] node6085;
	wire [8-1:0] node6088;
	wire [8-1:0] node6091;
	wire [8-1:0] node6092;
	wire [8-1:0] node6093;
	wire [8-1:0] node6096;
	wire [8-1:0] node6099;
	wire [8-1:0] node6100;
	wire [8-1:0] node6103;
	wire [8-1:0] node6106;
	wire [8-1:0] node6107;
	wire [8-1:0] node6108;
	wire [8-1:0] node6109;
	wire [8-1:0] node6110;
	wire [8-1:0] node6111;
	wire [8-1:0] node6114;
	wire [8-1:0] node6116;
	wire [8-1:0] node6119;
	wire [8-1:0] node6120;
	wire [8-1:0] node6122;
	wire [8-1:0] node6125;
	wire [8-1:0] node6126;
	wire [8-1:0] node6129;
	wire [8-1:0] node6132;
	wire [8-1:0] node6133;
	wire [8-1:0] node6135;
	wire [8-1:0] node6137;
	wire [8-1:0] node6140;
	wire [8-1:0] node6141;
	wire [8-1:0] node6142;
	wire [8-1:0] node6145;
	wire [8-1:0] node6148;
	wire [8-1:0] node6149;
	wire [8-1:0] node6153;
	wire [8-1:0] node6154;
	wire [8-1:0] node6155;
	wire [8-1:0] node6156;
	wire [8-1:0] node6158;
	wire [8-1:0] node6161;
	wire [8-1:0] node6163;
	wire [8-1:0] node6166;
	wire [8-1:0] node6168;
	wire [8-1:0] node6171;
	wire [8-1:0] node6172;
	wire [8-1:0] node6173;
	wire [8-1:0] node6175;
	wire [8-1:0] node6178;
	wire [8-1:0] node6179;
	wire [8-1:0] node6183;
	wire [8-1:0] node6184;
	wire [8-1:0] node6186;
	wire [8-1:0] node6189;
	wire [8-1:0] node6191;
	wire [8-1:0] node6194;
	wire [8-1:0] node6195;
	wire [8-1:0] node6196;
	wire [8-1:0] node6197;
	wire [8-1:0] node6198;
	wire [8-1:0] node6199;
	wire [8-1:0] node6203;
	wire [8-1:0] node6204;
	wire [8-1:0] node6207;
	wire [8-1:0] node6210;
	wire [8-1:0] node6211;
	wire [8-1:0] node6214;
	wire [8-1:0] node6216;
	wire [8-1:0] node6219;
	wire [8-1:0] node6220;
	wire [8-1:0] node6221;
	wire [8-1:0] node6222;
	wire [8-1:0] node6226;
	wire [8-1:0] node6227;
	wire [8-1:0] node6230;
	wire [8-1:0] node6233;
	wire [8-1:0] node6234;
	wire [8-1:0] node6235;
	wire [8-1:0] node6238;
	wire [8-1:0] node6241;
	wire [8-1:0] node6243;
	wire [8-1:0] node6246;
	wire [8-1:0] node6247;
	wire [8-1:0] node6248;
	wire [8-1:0] node6250;
	wire [8-1:0] node6252;
	wire [8-1:0] node6255;
	wire [8-1:0] node6256;
	wire [8-1:0] node6259;
	wire [8-1:0] node6262;
	wire [8-1:0] node6263;
	wire [8-1:0] node6264;
	wire [8-1:0] node6267;
	wire [8-1:0] node6270;
	wire [8-1:0] node6271;
	wire [8-1:0] node6272;
	wire [8-1:0] node6275;
	wire [8-1:0] node6278;
	wire [8-1:0] node6279;
	wire [8-1:0] node6282;
	wire [8-1:0] node6285;
	wire [8-1:0] node6286;
	wire [8-1:0] node6287;
	wire [8-1:0] node6288;
	wire [8-1:0] node6289;
	wire [8-1:0] node6290;
	wire [8-1:0] node6292;
	wire [8-1:0] node6294;
	wire [8-1:0] node6297;
	wire [8-1:0] node6298;
	wire [8-1:0] node6300;
	wire [8-1:0] node6302;
	wire [8-1:0] node6305;
	wire [8-1:0] node6307;
	wire [8-1:0] node6309;
	wire [8-1:0] node6312;
	wire [8-1:0] node6313;
	wire [8-1:0] node6314;
	wire [8-1:0] node6316;
	wire [8-1:0] node6319;
	wire [8-1:0] node6321;
	wire [8-1:0] node6324;
	wire [8-1:0] node6325;
	wire [8-1:0] node6327;
	wire [8-1:0] node6330;
	wire [8-1:0] node6332;
	wire [8-1:0] node6335;
	wire [8-1:0] node6336;
	wire [8-1:0] node6337;
	wire [8-1:0] node6338;
	wire [8-1:0] node6340;
	wire [8-1:0] node6343;
	wire [8-1:0] node6346;
	wire [8-1:0] node6347;
	wire [8-1:0] node6348;
	wire [8-1:0] node6352;
	wire [8-1:0] node6353;
	wire [8-1:0] node6357;
	wire [8-1:0] node6358;
	wire [8-1:0] node6359;
	wire [8-1:0] node6360;
	wire [8-1:0] node6364;
	wire [8-1:0] node6365;
	wire [8-1:0] node6369;
	wire [8-1:0] node6370;
	wire [8-1:0] node6372;
	wire [8-1:0] node6375;
	wire [8-1:0] node6378;
	wire [8-1:0] node6379;
	wire [8-1:0] node6380;
	wire [8-1:0] node6381;
	wire [8-1:0] node6382;
	wire [8-1:0] node6383;
	wire [8-1:0] node6384;
	wire [8-1:0] node6387;
	wire [8-1:0] node6390;
	wire [8-1:0] node6391;
	wire [8-1:0] node6393;
	wire [8-1:0] node6396;
	wire [8-1:0] node6397;
	wire [8-1:0] node6401;
	wire [8-1:0] node6402;
	wire [8-1:0] node6403;
	wire [8-1:0] node6404;
	wire [8-1:0] node6407;
	wire [8-1:0] node6410;
	wire [8-1:0] node6411;
	wire [8-1:0] node6414;
	wire [8-1:0] node6417;
	wire [8-1:0] node6420;
	wire [8-1:0] node6421;
	wire [8-1:0] node6422;
	wire [8-1:0] node6423;
	wire [8-1:0] node6426;
	wire [8-1:0] node6429;
	wire [8-1:0] node6431;
	wire [8-1:0] node6434;
	wire [8-1:0] node6435;
	wire [8-1:0] node6438;
	wire [8-1:0] node6439;
	wire [8-1:0] node6442;
	wire [8-1:0] node6445;
	wire [8-1:0] node6446;
	wire [8-1:0] node6447;
	wire [8-1:0] node6448;
	wire [8-1:0] node6451;
	wire [8-1:0] node6452;
	wire [8-1:0] node6453;
	wire [8-1:0] node6456;
	wire [8-1:0] node6460;
	wire [8-1:0] node6461;
	wire [8-1:0] node6462;
	wire [8-1:0] node6466;
	wire [8-1:0] node6468;
	wire [8-1:0] node6471;
	wire [8-1:0] node6472;
	wire [8-1:0] node6473;
	wire [8-1:0] node6474;
	wire [8-1:0] node6477;
	wire [8-1:0] node6480;
	wire [8-1:0] node6481;
	wire [8-1:0] node6484;
	wire [8-1:0] node6487;
	wire [8-1:0] node6488;
	wire [8-1:0] node6491;
	wire [8-1:0] node6492;
	wire [8-1:0] node6495;
	wire [8-1:0] node6498;
	wire [8-1:0] node6499;
	wire [8-1:0] node6500;
	wire [8-1:0] node6501;
	wire [8-1:0] node6502;
	wire [8-1:0] node6503;
	wire [8-1:0] node6507;
	wire [8-1:0] node6508;
	wire [8-1:0] node6512;
	wire [8-1:0] node6513;
	wire [8-1:0] node6514;
	wire [8-1:0] node6515;
	wire [8-1:0] node6519;
	wire [8-1:0] node6520;
	wire [8-1:0] node6524;
	wire [8-1:0] node6525;
	wire [8-1:0] node6528;
	wire [8-1:0] node6529;
	wire [8-1:0] node6533;
	wire [8-1:0] node6534;
	wire [8-1:0] node6535;
	wire [8-1:0] node6538;
	wire [8-1:0] node6539;
	wire [8-1:0] node6543;
	wire [8-1:0] node6544;
	wire [8-1:0] node6545;
	wire [8-1:0] node6549;
	wire [8-1:0] node6550;
	wire [8-1:0] node6554;
	wire [8-1:0] node6555;
	wire [8-1:0] node6556;
	wire [8-1:0] node6557;
	wire [8-1:0] node6558;
	wire [8-1:0] node6559;
	wire [8-1:0] node6562;
	wire [8-1:0] node6566;
	wire [8-1:0] node6568;
	wire [8-1:0] node6569;
	wire [8-1:0] node6573;
	wire [8-1:0] node6574;
	wire [8-1:0] node6575;
	wire [8-1:0] node6579;
	wire [8-1:0] node6580;
	wire [8-1:0] node6583;
	wire [8-1:0] node6586;
	wire [8-1:0] node6587;
	wire [8-1:0] node6588;
	wire [8-1:0] node6589;
	wire [8-1:0] node6591;
	wire [8-1:0] node6595;
	wire [8-1:0] node6596;
	wire [8-1:0] node6599;
	wire [8-1:0] node6602;
	wire [8-1:0] node6603;
	wire [8-1:0] node6606;
	wire [8-1:0] node6608;
	wire [8-1:0] node6611;
	wire [8-1:0] node6612;
	wire [8-1:0] node6613;
	wire [8-1:0] node6614;
	wire [8-1:0] node6615;
	wire [8-1:0] node6616;
	wire [8-1:0] node6617;
	wire [8-1:0] node6619;
	wire [8-1:0] node6622;
	wire [8-1:0] node6624;
	wire [8-1:0] node6627;
	wire [8-1:0] node6629;
	wire [8-1:0] node6632;
	wire [8-1:0] node6633;
	wire [8-1:0] node6634;
	wire [8-1:0] node6638;
	wire [8-1:0] node6639;
	wire [8-1:0] node6640;
	wire [8-1:0] node6644;
	wire [8-1:0] node6645;
	wire [8-1:0] node6649;
	wire [8-1:0] node6650;
	wire [8-1:0] node6651;
	wire [8-1:0] node6655;
	wire [8-1:0] node6656;
	wire [8-1:0] node6657;
	wire [8-1:0] node6661;
	wire [8-1:0] node6662;
	wire [8-1:0] node6666;
	wire [8-1:0] node6667;
	wire [8-1:0] node6668;
	wire [8-1:0] node6669;
	wire [8-1:0] node6672;
	wire [8-1:0] node6673;
	wire [8-1:0] node6674;
	wire [8-1:0] node6678;
	wire [8-1:0] node6679;
	wire [8-1:0] node6683;
	wire [8-1:0] node6684;
	wire [8-1:0] node6685;
	wire [8-1:0] node6687;
	wire [8-1:0] node6690;
	wire [8-1:0] node6691;
	wire [8-1:0] node6695;
	wire [8-1:0] node6696;
	wire [8-1:0] node6698;
	wire [8-1:0] node6701;
	wire [8-1:0] node6702;
	wire [8-1:0] node6705;
	wire [8-1:0] node6708;
	wire [8-1:0] node6709;
	wire [8-1:0] node6710;
	wire [8-1:0] node6711;
	wire [8-1:0] node6715;
	wire [8-1:0] node6716;
	wire [8-1:0] node6717;
	wire [8-1:0] node6721;
	wire [8-1:0] node6722;
	wire [8-1:0] node6726;
	wire [8-1:0] node6727;
	wire [8-1:0] node6728;
	wire [8-1:0] node6731;
	wire [8-1:0] node6733;
	wire [8-1:0] node6736;
	wire [8-1:0] node6739;
	wire [8-1:0] node6740;
	wire [8-1:0] node6741;
	wire [8-1:0] node6742;
	wire [8-1:0] node6743;
	wire [8-1:0] node6744;
	wire [8-1:0] node6748;
	wire [8-1:0] node6749;
	wire [8-1:0] node6752;
	wire [8-1:0] node6755;
	wire [8-1:0] node6756;
	wire [8-1:0] node6760;
	wire [8-1:0] node6761;
	wire [8-1:0] node6762;
	wire [8-1:0] node6763;
	wire [8-1:0] node6767;
	wire [8-1:0] node6768;
	wire [8-1:0] node6771;
	wire [8-1:0] node6774;
	wire [8-1:0] node6775;
	wire [8-1:0] node6779;
	wire [8-1:0] node6780;
	wire [8-1:0] node6781;
	wire [8-1:0] node6782;
	wire [8-1:0] node6783;
	wire [8-1:0] node6786;
	wire [8-1:0] node6787;
	wire [8-1:0] node6790;
	wire [8-1:0] node6793;
	wire [8-1:0] node6794;
	wire [8-1:0] node6797;
	wire [8-1:0] node6800;
	wire [8-1:0] node6801;
	wire [8-1:0] node6802;
	wire [8-1:0] node6803;
	wire [8-1:0] node6806;
	wire [8-1:0] node6809;
	wire [8-1:0] node6810;
	wire [8-1:0] node6813;
	wire [8-1:0] node6816;
	wire [8-1:0] node6817;
	wire [8-1:0] node6820;
	wire [8-1:0] node6823;
	wire [8-1:0] node6824;
	wire [8-1:0] node6825;
	wire [8-1:0] node6826;
	wire [8-1:0] node6829;
	wire [8-1:0] node6832;
	wire [8-1:0] node6833;
	wire [8-1:0] node6836;
	wire [8-1:0] node6839;
	wire [8-1:0] node6840;
	wire [8-1:0] node6843;
	wire [8-1:0] node6846;
	wire [8-1:0] node6847;
	wire [8-1:0] node6848;
	wire [8-1:0] node6849;
	wire [8-1:0] node6852;
	wire [8-1:0] node6853;
	wire [8-1:0] node6854;
	wire [8-1:0] node6855;
	wire [8-1:0] node6856;
	wire [8-1:0] node6857;
	wire [8-1:0] node6858;
	wire [8-1:0] node6859;
	wire [8-1:0] node6863;
	wire [8-1:0] node6865;
	wire [8-1:0] node6868;
	wire [8-1:0] node6869;
	wire [8-1:0] node6873;
	wire [8-1:0] node6874;
	wire [8-1:0] node6876;
	wire [8-1:0] node6879;
	wire [8-1:0] node6881;
	wire [8-1:0] node6884;
	wire [8-1:0] node6885;
	wire [8-1:0] node6887;
	wire [8-1:0] node6890;
	wire [8-1:0] node6891;
	wire [8-1:0] node6893;
	wire [8-1:0] node6896;
	wire [8-1:0] node6897;
	wire [8-1:0] node6901;
	wire [8-1:0] node6902;
	wire [8-1:0] node6903;
	wire [8-1:0] node6904;
	wire [8-1:0] node6908;
	wire [8-1:0] node6910;
	wire [8-1:0] node6913;
	wire [8-1:0] node6914;
	wire [8-1:0] node6916;
	wire [8-1:0] node6919;
	wire [8-1:0] node6920;
	wire [8-1:0] node6922;
	wire [8-1:0] node6925;
	wire [8-1:0] node6927;
	wire [8-1:0] node6930;
	wire [8-1:0] node6931;
	wire [8-1:0] node6932;
	wire [8-1:0] node6933;
	wire [8-1:0] node6934;
	wire [8-1:0] node6936;
	wire [8-1:0] node6938;
	wire [8-1:0] node6941;
	wire [8-1:0] node6943;
	wire [8-1:0] node6946;
	wire [8-1:0] node6947;
	wire [8-1:0] node6949;
	wire [8-1:0] node6952;
	wire [8-1:0] node6953;
	wire [8-1:0] node6957;
	wire [8-1:0] node6958;
	wire [8-1:0] node6959;
	wire [8-1:0] node6960;
	wire [8-1:0] node6964;
	wire [8-1:0] node6965;
	wire [8-1:0] node6969;
	wire [8-1:0] node6971;
	wire [8-1:0] node6974;
	wire [8-1:0] node6975;
	wire [8-1:0] node6976;
	wire [8-1:0] node6977;
	wire [8-1:0] node6978;
	wire [8-1:0] node6980;
	wire [8-1:0] node6984;
	wire [8-1:0] node6985;
	wire [8-1:0] node6986;
	wire [8-1:0] node6990;
	wire [8-1:0] node6993;
	wire [8-1:0] node6994;
	wire [8-1:0] node6995;
	wire [8-1:0] node6998;
	wire [8-1:0] node6999;
	wire [8-1:0] node7003;
	wire [8-1:0] node7005;
	wire [8-1:0] node7008;
	wire [8-1:0] node7009;
	wire [8-1:0] node7010;
	wire [8-1:0] node7011;
	wire [8-1:0] node7012;
	wire [8-1:0] node7016;
	wire [8-1:0] node7019;
	wire [8-1:0] node7020;
	wire [8-1:0] node7024;
	wire [8-1:0] node7025;
	wire [8-1:0] node7026;
	wire [8-1:0] node7030;
	wire [8-1:0] node7031;
	wire [8-1:0] node7035;
	wire [8-1:0] node7036;
	wire [8-1:0] node7037;
	wire [8-1:0] node7038;
	wire [8-1:0] node7039;
	wire [8-1:0] node7042;
	wire [8-1:0] node7043;
	wire [8-1:0] node7044;
	wire [8-1:0] node7049;
	wire [8-1:0] node7050;
	wire [8-1:0] node7051;
	wire [8-1:0] node7052;
	wire [8-1:0] node7057;
	wire [8-1:0] node7058;
	wire [8-1:0] node7059;
	wire [8-1:0] node7060;
	wire [8-1:0] node7064;
	wire [8-1:0] node7068;
	wire [8-1:0] node7069;
	wire [8-1:0] node7070;
	wire [8-1:0] node7071;
	wire [8-1:0] node7072;
	wire [8-1:0] node7077;
	wire [8-1:0] node7078;
	wire [8-1:0] node7079;
	wire [8-1:0] node7080;
	wire [8-1:0] node7084;
	wire [8-1:0] node7088;
	wire [8-1:0] node7089;
	wire [8-1:0] node7090;
	wire [8-1:0] node7091;
	wire [8-1:0] node7092;
	wire [8-1:0] node7094;
	wire [8-1:0] node7098;
	wire [8-1:0] node7100;
	wire [8-1:0] node7103;
	wire [8-1:0] node7104;
	wire [8-1:0] node7106;
	wire [8-1:0] node7109;
	wire [8-1:0] node7111;
	wire [8-1:0] node7114;
	wire [8-1:0] node7117;
	wire [8-1:0] node7118;
	wire [8-1:0] node7119;
	wire [8-1:0] node7120;
	wire [8-1:0] node7121;
	wire [8-1:0] node7122;
	wire [8-1:0] node7127;
	wire [8-1:0] node7128;
	wire [8-1:0] node7129;
	wire [8-1:0] node7130;
	wire [8-1:0] node7134;
	wire [8-1:0] node7138;
	wire [8-1:0] node7139;
	wire [8-1:0] node7140;
	wire [8-1:0] node7141;
	wire [8-1:0] node7142;
	wire [8-1:0] node7144;
	wire [8-1:0] node7147;
	wire [8-1:0] node7150;
	wire [8-1:0] node7152;
	wire [8-1:0] node7155;
	wire [8-1:0] node7156;
	wire [8-1:0] node7158;
	wire [8-1:0] node7161;
	wire [8-1:0] node7163;
	wire [8-1:0] node7166;
	wire [8-1:0] node7169;
	wire [8-1:0] node7170;
	wire [8-1:0] node7171;
	wire [8-1:0] node7172;
	wire [8-1:0] node7173;
	wire [8-1:0] node7174;
	wire [8-1:0] node7176;
	wire [8-1:0] node7179;
	wire [8-1:0] node7181;
	wire [8-1:0] node7184;
	wire [8-1:0] node7185;
	wire [8-1:0] node7187;
	wire [8-1:0] node7190;
	wire [8-1:0] node7192;
	wire [8-1:0] node7195;
	wire [8-1:0] node7196;
	wire [8-1:0] node7198;
	wire [8-1:0] node7201;
	wire [8-1:0] node7202;
	wire [8-1:0] node7204;
	wire [8-1:0] node7207;
	wire [8-1:0] node7209;
	wire [8-1:0] node7212;
	wire [8-1:0] node7213;
	wire [8-1:0] node7214;
	wire [8-1:0] node7216;
	wire [8-1:0] node7219;
	wire [8-1:0] node7220;
	wire [8-1:0] node7222;
	wire [8-1:0] node7225;
	wire [8-1:0] node7227;
	wire [8-1:0] node7230;
	wire [8-1:0] node7231;
	wire [8-1:0] node7233;
	wire [8-1:0] node7236;
	wire [8-1:0] node7237;
	wire [8-1:0] node7239;
	wire [8-1:0] node7242;
	wire [8-1:0] node7244;
	wire [8-1:0] node7247;
	wire [8-1:0] node7248;
	wire [8-1:0] node7251;
	wire [8-1:0] node7254;
	wire [8-1:0] node7255;
	wire [8-1:0] node7256;
	wire [8-1:0] node7258;
	wire [8-1:0] node7259;
	wire [8-1:0] node7260;
	wire [8-1:0] node7261;
	wire [8-1:0] node7262;
	wire [8-1:0] node7263;
	wire [8-1:0] node7266;
	wire [8-1:0] node7267;
	wire [8-1:0] node7271;
	wire [8-1:0] node7272;
	wire [8-1:0] node7276;
	wire [8-1:0] node7277;
	wire [8-1:0] node7278;
	wire [8-1:0] node7282;
	wire [8-1:0] node7283;
	wire [8-1:0] node7284;
	wire [8-1:0] node7288;
	wire [8-1:0] node7291;
	wire [8-1:0] node7292;
	wire [8-1:0] node7294;
	wire [8-1:0] node7297;
	wire [8-1:0] node7298;
	wire [8-1:0] node7299;
	wire [8-1:0] node7303;
	wire [8-1:0] node7305;
	wire [8-1:0] node7308;
	wire [8-1:0] node7309;
	wire [8-1:0] node7310;
	wire [8-1:0] node7311;
	wire [8-1:0] node7312;
	wire [8-1:0] node7313;
	wire [8-1:0] node7317;
	wire [8-1:0] node7319;
	wire [8-1:0] node7322;
	wire [8-1:0] node7323;
	wire [8-1:0] node7324;
	wire [8-1:0] node7327;
	wire [8-1:0] node7329;
	wire [8-1:0] node7332;
	wire [8-1:0] node7333;
	wire [8-1:0] node7337;
	wire [8-1:0] node7338;
	wire [8-1:0] node7340;
	wire [8-1:0] node7343;
	wire [8-1:0] node7344;
	wire [8-1:0] node7345;
	wire [8-1:0] node7349;
	wire [8-1:0] node7350;
	wire [8-1:0] node7354;
	wire [8-1:0] node7355;
	wire [8-1:0] node7356;
	wire [8-1:0] node7357;
	wire [8-1:0] node7358;
	wire [8-1:0] node7362;
	wire [8-1:0] node7364;
	wire [8-1:0] node7367;
	wire [8-1:0] node7369;
	wire [8-1:0] node7372;
	wire [8-1:0] node7373;
	wire [8-1:0] node7374;
	wire [8-1:0] node7376;
	wire [8-1:0] node7377;
	wire [8-1:0] node7381;
	wire [8-1:0] node7384;
	wire [8-1:0] node7385;
	wire [8-1:0] node7387;
	wire [8-1:0] node7390;
	wire [8-1:0] node7391;
	wire [8-1:0] node7394;
	wire [8-1:0] node7397;
	wire [8-1:0] node7398;
	wire [8-1:0] node7399;
	wire [8-1:0] node7400;
	wire [8-1:0] node7402;
	wire [8-1:0] node7403;
	wire [8-1:0] node7407;
	wire [8-1:0] node7408;
	wire [8-1:0] node7409;
	wire [8-1:0] node7411;
	wire [8-1:0] node7414;
	wire [8-1:0] node7417;
	wire [8-1:0] node7419;
	wire [8-1:0] node7420;
	wire [8-1:0] node7424;
	wire [8-1:0] node7425;
	wire [8-1:0] node7426;
	wire [8-1:0] node7427;
	wire [8-1:0] node7429;
	wire [8-1:0] node7432;
	wire [8-1:0] node7434;
	wire [8-1:0] node7437;
	wire [8-1:0] node7440;
	wire [8-1:0] node7441;
	wire [8-1:0] node7442;
	wire [8-1:0] node7443;
	wire [8-1:0] node7446;
	wire [8-1:0] node7448;
	wire [8-1:0] node7451;
	wire [8-1:0] node7452;
	wire [8-1:0] node7454;
	wire [8-1:0] node7457;
	wire [8-1:0] node7458;
	wire [8-1:0] node7462;
	wire [8-1:0] node7465;
	wire [8-1:0] node7466;
	wire [8-1:0] node7467;
	wire [8-1:0] node7468;
	wire [8-1:0] node7469;
	wire [8-1:0] node7473;
	wire [8-1:0] node7474;
	wire [8-1:0] node7475;
	wire [8-1:0] node7478;
	wire [8-1:0] node7482;
	wire [8-1:0] node7483;
	wire [8-1:0] node7484;
	wire [8-1:0] node7485;
	wire [8-1:0] node7488;
	wire [8-1:0] node7492;
	wire [8-1:0] node7493;
	wire [8-1:0] node7494;
	wire [8-1:0] node7495;
	wire [8-1:0] node7498;
	wire [8-1:0] node7501;
	wire [8-1:0] node7502;
	wire [8-1:0] node7505;
	wire [8-1:0] node7509;
	wire [8-1:0] node7510;
	wire [8-1:0] node7511;
	wire [8-1:0] node7512;
	wire [8-1:0] node7513;
	wire [8-1:0] node7515;
	wire [8-1:0] node7518;
	wire [8-1:0] node7519;
	wire [8-1:0] node7521;
	wire [8-1:0] node7525;
	wire [8-1:0] node7526;
	wire [8-1:0] node7528;
	wire [8-1:0] node7531;
	wire [8-1:0] node7534;
	wire [8-1:0] node7535;
	wire [8-1:0] node7536;
	wire [8-1:0] node7538;
	wire [8-1:0] node7541;
	wire [8-1:0] node7543;
	wire [8-1:0] node7546;
	wire [8-1:0] node7548;
	wire [8-1:0] node7549;
	wire [8-1:0] node7551;
	wire [8-1:0] node7554;
	wire [8-1:0] node7557;
	wire [8-1:0] node7558;
	wire [8-1:0] node7561;
	wire [8-1:0] node7564;
	wire [8-1:0] node7565;
	wire [8-1:0] node7567;
	wire [8-1:0] node7568;
	wire [8-1:0] node7569;
	wire [8-1:0] node7570;
	wire [8-1:0] node7571;
	wire [8-1:0] node7573;
	wire [8-1:0] node7576;
	wire [8-1:0] node7577;
	wire [8-1:0] node7579;
	wire [8-1:0] node7582;
	wire [8-1:0] node7584;
	wire [8-1:0] node7587;
	wire [8-1:0] node7588;
	wire [8-1:0] node7589;
	wire [8-1:0] node7591;
	wire [8-1:0] node7594;
	wire [8-1:0] node7595;
	wire [8-1:0] node7599;
	wire [8-1:0] node7600;
	wire [8-1:0] node7602;
	wire [8-1:0] node7605;
	wire [8-1:0] node7607;
	wire [8-1:0] node7608;
	wire [8-1:0] node7612;
	wire [8-1:0] node7613;
	wire [8-1:0] node7614;
	wire [8-1:0] node7615;
	wire [8-1:0] node7619;
	wire [8-1:0] node7620;
	wire [8-1:0] node7622;
	wire [8-1:0] node7625;
	wire [8-1:0] node7626;
	wire [8-1:0] node7630;
	wire [8-1:0] node7631;
	wire [8-1:0] node7632;
	wire [8-1:0] node7634;
	wire [8-1:0] node7637;
	wire [8-1:0] node7640;
	wire [8-1:0] node7641;
	wire [8-1:0] node7642;
	wire [8-1:0] node7645;
	wire [8-1:0] node7649;
	wire [8-1:0] node7650;
	wire [8-1:0] node7651;
	wire [8-1:0] node7652;
	wire [8-1:0] node7654;
	wire [8-1:0] node7657;
	wire [8-1:0] node7658;
	wire [8-1:0] node7662;
	wire [8-1:0] node7663;
	wire [8-1:0] node7667;
	wire [8-1:0] node7668;
	wire [8-1:0] node7669;
	wire [8-1:0] node7671;
	wire [8-1:0] node7673;
	wire [8-1:0] node7676;
	wire [8-1:0] node7678;
	wire [8-1:0] node7681;
	wire [8-1:0] node7682;
	wire [8-1:0] node7683;
	wire [8-1:0] node7687;
	wire [8-1:0] node7688;
	wire [8-1:0] node7690;
	wire [8-1:0] node7693;
	wire [8-1:0] node7694;
	wire [8-1:0] node7698;
	wire [8-1:0] node7699;
	wire [8-1:0] node7700;
	wire [8-1:0] node7701;
	wire [8-1:0] node7703;
	wire [8-1:0] node7704;
	wire [8-1:0] node7708;
	wire [8-1:0] node7709;
	wire [8-1:0] node7710;
	wire [8-1:0] node7712;
	wire [8-1:0] node7715;
	wire [8-1:0] node7718;
	wire [8-1:0] node7720;
	wire [8-1:0] node7721;
	wire [8-1:0] node7725;
	wire [8-1:0] node7726;
	wire [8-1:0] node7727;
	wire [8-1:0] node7728;
	wire [8-1:0] node7730;
	wire [8-1:0] node7733;
	wire [8-1:0] node7734;
	wire [8-1:0] node7736;
	wire [8-1:0] node7739;
	wire [8-1:0] node7741;
	wire [8-1:0] node7744;
	wire [8-1:0] node7745;
	wire [8-1:0] node7748;
	wire [8-1:0] node7751;
	wire [8-1:0] node7752;
	wire [8-1:0] node7754;
	wire [8-1:0] node7755;
	wire [8-1:0] node7759;
	wire [8-1:0] node7760;
	wire [8-1:0] node7761;
	wire [8-1:0] node7765;
	wire [8-1:0] node7766;
	wire [8-1:0] node7767;
	wire [8-1:0] node7770;
	wire [8-1:0] node7774;
	wire [8-1:0] node7775;
	wire [8-1:0] node7776;
	wire [8-1:0] node7777;
	wire [8-1:0] node7778;
	wire [8-1:0] node7780;
	wire [8-1:0] node7783;
	wire [8-1:0] node7784;
	wire [8-1:0] node7786;
	wire [8-1:0] node7789;
	wire [8-1:0] node7791;
	wire [8-1:0] node7794;
	wire [8-1:0] node7795;
	wire [8-1:0] node7796;
	wire [8-1:0] node7798;
	wire [8-1:0] node7801;
	wire [8-1:0] node7803;
	wire [8-1:0] node7805;
	wire [8-1:0] node7808;
	wire [8-1:0] node7809;
	wire [8-1:0] node7811;
	wire [8-1:0] node7814;
	wire [8-1:0] node7815;
	wire [8-1:0] node7819;
	wire [8-1:0] node7820;
	wire [8-1:0] node7821;
	wire [8-1:0] node7824;
	wire [8-1:0] node7827;
	wire [8-1:0] node7828;
	wire [8-1:0] node7831;
	wire [8-1:0] node7834;
	wire [8-1:0] node7835;
	wire [8-1:0] node7836;
	wire [8-1:0] node7838;
	wire [8-1:0] node7839;
	wire [8-1:0] node7843;
	wire [8-1:0] node7844;
	wire [8-1:0] node7845;
	wire [8-1:0] node7847;
	wire [8-1:0] node7850;
	wire [8-1:0] node7852;
	wire [8-1:0] node7855;
	wire [8-1:0] node7858;
	wire [8-1:0] node7859;
	wire [8-1:0] node7860;
	wire [8-1:0] node7861;
	wire [8-1:0] node7865;
	wire [8-1:0] node7866;
	wire [8-1:0] node7867;
	wire [8-1:0] node7870;
	wire [8-1:0] node7874;
	wire [8-1:0] node7875;
	wire [8-1:0] node7876;
	wire [8-1:0] node7879;
	wire [8-1:0] node7880;
	wire [8-1:0] node7882;
	wire [8-1:0] node7886;

	assign outp = (inp[7]) ? node4062 : node1;
		assign node1 = (inp[13]) ? node1919 : node2;
			assign node2 = (inp[4]) ? node398 : node3;
				assign node3 = (inp[11]) ? node127 : node4;
					assign node4 = (inp[0]) ? node72 : node5;
						assign node5 = (inp[1]) ? node29 : node6;
							assign node6 = (inp[8]) ? node14 : node7;
								assign node7 = (inp[2]) ? node9 : 8'b01111111;
									assign node9 = (inp[6]) ? node11 : 8'b00101111;
										assign node11 = (inp[5]) ? 8'b01111111 : 8'b00101111;
								assign node14 = (inp[5]) ? node18 : node15;
									assign node15 = (inp[2]) ? 8'b00101011 : 8'b00111011;
									assign node18 = (inp[10]) ? node24 : node19;
										assign node19 = (inp[2]) ? node21 : 8'b00111011;
											assign node21 = (inp[6]) ? 8'b00111011 : 8'b00101011;
										assign node24 = (inp[6]) ? 8'b01111111 : node25;
											assign node25 = (inp[2]) ? 8'b00101111 : 8'b01111111;
							assign node29 = (inp[2]) ? node45 : node30;
								assign node30 = (inp[8]) ? node36 : node31;
									assign node31 = (inp[3]) ? node33 : 8'b00111110;
										assign node33 = (inp[5]) ? 8'b01111111 : 8'b00111110;
									assign node36 = (inp[5]) ? node38 : 8'b00111010;
										assign node38 = (inp[3]) ? node42 : node39;
											assign node39 = (inp[10]) ? 8'b00111110 : 8'b00111010;
											assign node42 = (inp[10]) ? 8'b01111111 : 8'b00111011;
								assign node45 = (inp[5]) ? node49 : node46;
									assign node46 = (inp[8]) ? 8'b00101010 : 8'b00101110;
									assign node49 = (inp[3]) ? node61 : node50;
										assign node50 = (inp[6]) ? node56 : node51;
											assign node51 = (inp[10]) ? 8'b00101110 : node52;
												assign node52 = (inp[8]) ? 8'b00101010 : 8'b00101110;
											assign node56 = (inp[10]) ? 8'b00111110 : node57;
												assign node57 = (inp[8]) ? 8'b00111010 : 8'b00111110;
										assign node61 = (inp[6]) ? node67 : node62;
											assign node62 = (inp[8]) ? node64 : 8'b00101111;
												assign node64 = (inp[10]) ? 8'b00101111 : 8'b00101011;
											assign node67 = (inp[10]) ? 8'b01111111 : node68;
												assign node68 = (inp[8]) ? 8'b00111011 : 8'b01111111;
						assign node72 = (inp[5]) ? 8'b01111111 : node73;
							assign node73 = (inp[10]) ? node91 : node74;
								assign node74 = (inp[1]) ? node80 : node75;
									assign node75 = (inp[6]) ? node77 : 8'b01111111;
										assign node77 = (inp[2]) ? 8'b00101111 : 8'b01111111;
									assign node80 = (inp[3]) ? node86 : node81;
										assign node81 = (inp[2]) ? node83 : 8'b01111111;
											assign node83 = (inp[6]) ? 8'b00101111 : 8'b01111111;
										assign node86 = (inp[2]) ? node88 : 8'b00111110;
											assign node88 = (inp[6]) ? 8'b00101110 : 8'b00111110;
								assign node91 = (inp[8]) ? node109 : node92;
									assign node92 = (inp[6]) ? node98 : node93;
										assign node93 = (inp[3]) ? node95 : 8'b01111111;
											assign node95 = (inp[1]) ? 8'b00111110 : 8'b01111111;
										assign node98 = (inp[2]) ? node104 : node99;
											assign node99 = (inp[1]) ? node101 : 8'b01111111;
												assign node101 = (inp[3]) ? 8'b00111110 : 8'b01111111;
											assign node104 = (inp[3]) ? node106 : 8'b00101111;
												assign node106 = (inp[1]) ? 8'b00101110 : 8'b00101111;
									assign node109 = (inp[3]) ? node115 : node110;
										assign node110 = (inp[6]) ? node112 : 8'b00111011;
											assign node112 = (inp[2]) ? 8'b00101011 : 8'b00111011;
										assign node115 = (inp[1]) ? node121 : node116;
											assign node116 = (inp[2]) ? node118 : 8'b00111011;
												assign node118 = (inp[6]) ? 8'b00101011 : 8'b00111011;
											assign node121 = (inp[6]) ? node123 : 8'b00111010;
												assign node123 = (inp[2]) ? 8'b00101010 : 8'b00111010;
					assign node127 = (inp[8]) ? node219 : node128;
						assign node128 = (inp[1]) ? node156 : node129;
							assign node129 = (inp[2]) ? node133 : node130;
								assign node130 = (inp[12]) ? 8'b01111111 : 8'b00101111;
								assign node133 = (inp[12]) ? node145 : node134;
									assign node134 = (inp[0]) ? node140 : node135;
										assign node135 = (inp[6]) ? node137 : 8'b00111110;
											assign node137 = (inp[5]) ? 8'b00101110 : 8'b00111110;
										assign node140 = (inp[6]) ? node142 : 8'b00101110;
											assign node142 = (inp[5]) ? 8'b00101110 : 8'b00111110;
									assign node145 = (inp[5]) ? node151 : node146;
										assign node146 = (inp[6]) ? 8'b00101111 : node147;
											assign node147 = (inp[0]) ? 8'b00111110 : 8'b00101111;
										assign node151 = (inp[6]) ? 8'b00111110 : node152;
											assign node152 = (inp[0]) ? 8'b00111110 : 8'b00101111;
							assign node156 = (inp[12]) ? node188 : node157;
								assign node157 = (inp[2]) ? node169 : node158;
									assign node158 = (inp[5]) ? node164 : node159;
										assign node159 = (inp[0]) ? node161 : 8'b00101110;
											assign node161 = (inp[3]) ? 8'b00101110 : 8'b00101011;
										assign node164 = (inp[3]) ? 8'b00101011 : node165;
											assign node165 = (inp[0]) ? 8'b00101011 : 8'b00101110;
									assign node169 = (inp[5]) ? node179 : node170;
										assign node170 = (inp[0]) ? node172 : 8'b00111011;
											assign node172 = (inp[3]) ? node176 : node173;
												assign node173 = (inp[6]) ? 8'b00111010 : 8'b00101010;
												assign node176 = (inp[6]) ? 8'b00111011 : 8'b00101011;
										assign node179 = (inp[0]) ? 8'b00101010 : node180;
											assign node180 = (inp[6]) ? node184 : node181;
												assign node181 = (inp[3]) ? 8'b00111010 : 8'b00111011;
												assign node184 = (inp[3]) ? 8'b00101010 : 8'b00101011;
								assign node188 = (inp[0]) ? node204 : node189;
									assign node189 = (inp[2]) ? node195 : node190;
										assign node190 = (inp[3]) ? node192 : 8'b00111110;
											assign node192 = (inp[5]) ? 8'b00111011 : 8'b00111110;
										assign node195 = (inp[5]) ? node197 : 8'b00101110;
											assign node197 = (inp[6]) ? node201 : node198;
												assign node198 = (inp[3]) ? 8'b00101011 : 8'b00101110;
												assign node201 = (inp[3]) ? 8'b00111010 : 8'b00111011;
									assign node204 = (inp[2]) ? node210 : node205;
										assign node205 = (inp[3]) ? node207 : 8'b00111011;
											assign node207 = (inp[5]) ? 8'b00111011 : 8'b00111110;
										assign node210 = (inp[5]) ? 8'b00111010 : node211;
											assign node211 = (inp[6]) ? node215 : node212;
												assign node212 = (inp[3]) ? 8'b00111011 : 8'b00111010;
												assign node215 = (inp[3]) ? 8'b00101110 : 8'b00101011;
						assign node219 = (inp[12]) ? node307 : node220;
							assign node220 = (inp[2]) ? node252 : node221;
								assign node221 = (inp[0]) ? node237 : node222;
									assign node222 = (inp[1]) ? node228 : node223;
										assign node223 = (inp[10]) ? node225 : 8'b00101011;
											assign node225 = (inp[5]) ? 8'b00001111 : 8'b00101011;
										assign node228 = (inp[5]) ? node230 : 8'b00101010;
											assign node230 = (inp[3]) ? node234 : node231;
												assign node231 = (inp[10]) ? 8'b00001110 : 8'b00101010;
												assign node234 = (inp[10]) ? 8'b00001011 : 8'b00001111;
									assign node237 = (inp[1]) ? node243 : node238;
										assign node238 = (inp[5]) ? 8'b00001111 : node239;
											assign node239 = (inp[10]) ? 8'b00101011 : 8'b00001111;
										assign node243 = (inp[5]) ? 8'b00001011 : node244;
											assign node244 = (inp[3]) ? node248 : node245;
												assign node245 = (inp[10]) ? 8'b00001111 : 8'b00001011;
												assign node248 = (inp[10]) ? 8'b00101010 : 8'b00001110;
								assign node252 = (inp[1]) ? node272 : node253;
									assign node253 = (inp[0]) ? node263 : node254;
										assign node254 = (inp[5]) ? node256 : 8'b00111010;
											assign node256 = (inp[10]) ? node260 : node257;
												assign node257 = (inp[6]) ? 8'b00101010 : 8'b00111010;
												assign node260 = (inp[6]) ? 8'b00001110 : 8'b00011110;
										assign node263 = (inp[5]) ? 8'b00001110 : node264;
											assign node264 = (inp[10]) ? node268 : node265;
												assign node265 = (inp[6]) ? 8'b00011110 : 8'b00001110;
												assign node268 = (inp[6]) ? 8'b00111010 : 8'b00101010;
									assign node272 = (inp[5]) ? node290 : node273;
										assign node273 = (inp[0]) ? node275 : 8'b00011111;
											assign node275 = (inp[6]) ? node283 : node276;
												assign node276 = (inp[3]) ? node280 : node277;
													assign node277 = (inp[10]) ? 8'b00001110 : 8'b00001010;
													assign node280 = (inp[10]) ? 8'b00001111 : 8'b00001011;
												assign node283 = (inp[10]) ? node287 : node284;
													assign node284 = (inp[3]) ? 8'b00011011 : 8'b00011010;
													assign node287 = (inp[3]) ? 8'b00011111 : 8'b00011110;
										assign node290 = (inp[0]) ? 8'b00001010 : node291;
											assign node291 = (inp[6]) ? node299 : node292;
												assign node292 = (inp[3]) ? node296 : node293;
													assign node293 = (inp[10]) ? 8'b00011011 : 8'b00011111;
													assign node296 = (inp[10]) ? 8'b00011010 : 8'b00011110;
												assign node299 = (inp[10]) ? node303 : node300;
													assign node300 = (inp[3]) ? 8'b00001110 : 8'b00001111;
													assign node303 = (inp[3]) ? 8'b00001010 : 8'b00001011;
							assign node307 = (inp[2]) ? node341 : node308;
								assign node308 = (inp[5]) ? node326 : node309;
									assign node309 = (inp[0]) ? node313 : node310;
										assign node310 = (inp[1]) ? 8'b00111010 : 8'b00111011;
										assign node313 = (inp[10]) ? node321 : node314;
											assign node314 = (inp[3]) ? node318 : node315;
												assign node315 = (inp[1]) ? 8'b00011011 : 8'b00011111;
												assign node318 = (inp[1]) ? 8'b00011110 : 8'b00011111;
											assign node321 = (inp[1]) ? node323 : 8'b00111011;
												assign node323 = (inp[3]) ? 8'b00111010 : 8'b00011111;
									assign node326 = (inp[1]) ? node332 : node327;
										assign node327 = (inp[0]) ? 8'b00011111 : node328;
											assign node328 = (inp[10]) ? 8'b00011111 : 8'b00111011;
										assign node332 = (inp[0]) ? 8'b00011011 : node333;
											assign node333 = (inp[3]) ? node337 : node334;
												assign node334 = (inp[10]) ? 8'b00011110 : 8'b00111010;
												assign node337 = (inp[10]) ? 8'b00011011 : 8'b00011111;
								assign node341 = (inp[0]) ? node369 : node342;
									assign node342 = (inp[5]) ? node346 : node343;
										assign node343 = (inp[1]) ? 8'b00101010 : 8'b00101011;
										assign node346 = (inp[6]) ? node358 : node347;
											assign node347 = (inp[10]) ? node353 : node348;
												assign node348 = (inp[1]) ? node350 : 8'b00101011;
													assign node350 = (inp[3]) ? 8'b00001111 : 8'b00101010;
												assign node353 = (inp[1]) ? node355 : 8'b00001111;
													assign node355 = (inp[3]) ? 8'b00001011 : 8'b00001110;
											assign node358 = (inp[1]) ? node362 : node359;
												assign node359 = (inp[10]) ? 8'b00011110 : 8'b00111010;
												assign node362 = (inp[3]) ? node366 : node363;
													assign node363 = (inp[10]) ? 8'b00011011 : 8'b00011111;
													assign node366 = (inp[10]) ? 8'b00011010 : 8'b00011110;
									assign node369 = (inp[5]) ? node395 : node370;
										assign node370 = (inp[6]) ? node382 : node371;
											assign node371 = (inp[1]) ? node375 : node372;
												assign node372 = (inp[10]) ? 8'b00111010 : 8'b00011110;
												assign node375 = (inp[10]) ? node379 : node376;
													assign node376 = (inp[3]) ? 8'b00011011 : 8'b00011010;
													assign node379 = (inp[3]) ? 8'b00011111 : 8'b00011110;
											assign node382 = (inp[10]) ? node390 : node383;
												assign node383 = (inp[3]) ? node387 : node384;
													assign node384 = (inp[1]) ? 8'b00001011 : 8'b00001111;
													assign node387 = (inp[1]) ? 8'b00001110 : 8'b00001111;
												assign node390 = (inp[1]) ? node392 : 8'b00101011;
													assign node392 = (inp[3]) ? 8'b00101010 : 8'b00001111;
										assign node395 = (inp[1]) ? 8'b00011010 : 8'b00011110;
				assign node398 = (inp[9]) ? node1164 : node399;
					assign node399 = (inp[8]) ? node759 : node400;
						assign node400 = (inp[10]) ? node594 : node401;
							assign node401 = (inp[1]) ? node491 : node402;
								assign node402 = (inp[3]) ? node442 : node403;
									assign node403 = (inp[2]) ? node415 : node404;
										assign node404 = (inp[6]) ? node410 : node405;
											assign node405 = (inp[12]) ? 8'b00000010 : node406;
												assign node406 = (inp[11]) ? 8'b11110111 : 8'b10000010;
											assign node410 = (inp[12]) ? 8'b00011010 : node411;
												assign node411 = (inp[11]) ? 8'b00001010 : 8'b00011010;
										assign node415 = (inp[11]) ? node429 : node416;
											assign node416 = (inp[0]) ? node424 : node417;
												assign node417 = (inp[12]) ? node419 : 8'b10000010;
													assign node419 = (inp[5]) ? node421 : 8'b00000010;
														assign node421 = (inp[6]) ? 8'b10010000 : 8'b00000010;
												assign node424 = (inp[6]) ? node426 : 8'b10010000;
													assign node426 = (inp[5]) ? 8'b10010000 : 8'b00000010;
											assign node429 = (inp[12]) ? node435 : node430;
												assign node430 = (inp[5]) ? 8'b10100101 : node431;
													assign node431 = (inp[6]) ? 8'b11110111 : 8'b10100101;
												assign node435 = (inp[5]) ? node439 : node436;
													assign node436 = (inp[6]) ? 8'b00000010 : 8'b11110101;
													assign node439 = (inp[6]) ? 8'b11110101 : 8'b00000010;
									assign node442 = (inp[11]) ? node460 : node443;
										assign node443 = (inp[0]) ? node451 : node444;
											assign node444 = (inp[6]) ? node446 : 8'b00001011;
												assign node446 = (inp[5]) ? 8'b00011011 : node447;
													assign node447 = (inp[2]) ? 8'b00001011 : 8'b00011011;
											assign node451 = (inp[5]) ? 8'b00011011 : node452;
												assign node452 = (inp[6]) ? node456 : node453;
													assign node453 = (inp[2]) ? 8'b00011011 : 8'b00001011;
													assign node456 = (inp[2]) ? 8'b00001011 : 8'b00011011;
										assign node460 = (inp[2]) ? node468 : node461;
											assign node461 = (inp[12]) ? node465 : node462;
												assign node462 = (inp[6]) ? 8'b00001011 : 8'b00011010;
												assign node465 = (inp[6]) ? 8'b00011011 : 8'b00001011;
											assign node468 = (inp[12]) ? node480 : node469;
												assign node469 = (inp[5]) ? node475 : node470;
													assign node470 = (inp[6]) ? 8'b00011010 : node471;
														assign node471 = (inp[0]) ? 8'b00001010 : 8'b00011010;
													assign node475 = (inp[0]) ? 8'b00001010 : node476;
														assign node476 = (inp[6]) ? 8'b00001010 : 8'b00011010;
												assign node480 = (inp[5]) ? node486 : node481;
													assign node481 = (inp[0]) ? node483 : 8'b00001011;
														assign node483 = (inp[6]) ? 8'b00001011 : 8'b00011010;
													assign node486 = (inp[0]) ? 8'b00011010 : node487;
														assign node487 = (inp[6]) ? 8'b00011010 : 8'b00001011;
								assign node491 = (inp[11]) ? node539 : node492;
									assign node492 = (inp[6]) ? node514 : node493;
										assign node493 = (inp[0]) ? node503 : node494;
											assign node494 = (inp[3]) ? node498 : node495;
												assign node495 = (inp[12]) ? 8'b00000010 : 8'b10000010;
												assign node498 = (inp[5]) ? 8'b10000001 : node499;
													assign node499 = (inp[12]) ? 8'b00000010 : 8'b10000010;
											assign node503 = (inp[2]) ? node509 : node504;
												assign node504 = (inp[3]) ? node506 : 8'b10000001;
													assign node506 = (inp[12]) ? 8'b10000001 : 8'b10000010;
												assign node509 = (inp[3]) ? node511 : 8'b10010001;
													assign node511 = (inp[5]) ? 8'b10010001 : 8'b10010000;
										assign node514 = (inp[2]) ? node526 : node515;
											assign node515 = (inp[5]) ? node521 : node516;
												assign node516 = (inp[3]) ? 8'b00011010 : node517;
													assign node517 = (inp[0]) ? 8'b10011001 : 8'b00011010;
												assign node521 = (inp[3]) ? 8'b10011001 : node522;
													assign node522 = (inp[0]) ? 8'b10011001 : 8'b00011010;
											assign node526 = (inp[5]) ? node534 : node527;
												assign node527 = (inp[12]) ? node529 : 8'b10000010;
													assign node529 = (inp[0]) ? node531 : 8'b00000010;
														assign node531 = (inp[3]) ? 8'b00000010 : 8'b10000001;
												assign node534 = (inp[3]) ? 8'b10010001 : node535;
													assign node535 = (inp[0]) ? 8'b10010001 : 8'b10010000;
									assign node539 = (inp[2]) ? node569 : node540;
										assign node540 = (inp[5]) ? node552 : node541;
											assign node541 = (inp[6]) ? node545 : node542;
												assign node542 = (inp[12]) ? 8'b00000010 : 8'b11110111;
												assign node545 = (inp[12]) ? 8'b00011010 : node546;
													assign node546 = (inp[3]) ? 8'b00001010 : node547;
														assign node547 = (inp[0]) ? 8'b10101101 : 8'b00001010;
											assign node552 = (inp[3]) ? node562 : node553;
												assign node553 = (inp[6]) ? node559 : node554;
													assign node554 = (inp[12]) ? 8'b00000010 : node555;
														assign node555 = (inp[0]) ? 8'b10110100 : 8'b11110111;
													assign node559 = (inp[12]) ? 8'b00011010 : 8'b00001010;
												assign node562 = (inp[6]) ? node566 : node563;
													assign node563 = (inp[12]) ? 8'b10100101 : 8'b10110100;
													assign node566 = (inp[12]) ? 8'b11111101 : 8'b10101101;
										assign node569 = (inp[0]) ? node579 : node570;
											assign node570 = (inp[5]) ? node574 : node571;
												assign node571 = (inp[12]) ? 8'b00000010 : 8'b11110111;
												assign node574 = (inp[3]) ? 8'b10100101 : node575;
													assign node575 = (inp[12]) ? 8'b11110101 : 8'b10100101;
											assign node579 = (inp[12]) ? node589 : node580;
												assign node580 = (inp[5]) ? 8'b10100100 : node581;
													assign node581 = (inp[6]) ? node585 : node582;
														assign node582 = (inp[3]) ? 8'b10100101 : 8'b10100100;
														assign node585 = (inp[3]) ? 8'b11110111 : 8'b10110100;
												assign node589 = (inp[5]) ? 8'b10110100 : node590;
													assign node590 = (inp[3]) ? 8'b11110101 : 8'b10110100;
							assign node594 = (inp[11]) ? node648 : node595;
								assign node595 = (inp[3]) ? node619 : node596;
									assign node596 = (inp[0]) ? node604 : node597;
										assign node597 = (inp[6]) ? node599 : 8'b00001110;
											assign node599 = (inp[2]) ? node601 : 8'b00011110;
												assign node601 = (inp[5]) ? 8'b00011110 : 8'b00001110;
										assign node604 = (inp[1]) ? node610 : node605;
											assign node605 = (inp[2]) ? 8'b00011110 : node606;
												assign node606 = (inp[6]) ? 8'b00011110 : 8'b00001110;
											assign node610 = (inp[2]) ? node614 : node611;
												assign node611 = (inp[6]) ? 8'b00011111 : 8'b00001111;
												assign node614 = (inp[6]) ? node616 : 8'b00011111;
													assign node616 = (inp[5]) ? 8'b00011111 : 8'b00001111;
									assign node619 = (inp[1]) ? node631 : node620;
										assign node620 = (inp[6]) ? node626 : node621;
											assign node621 = (inp[2]) ? node623 : 8'b00001111;
												assign node623 = (inp[0]) ? 8'b00011111 : 8'b00001111;
											assign node626 = (inp[2]) ? node628 : 8'b00011111;
												assign node628 = (inp[5]) ? 8'b00011111 : 8'b00001111;
										assign node631 = (inp[5]) ? node645 : node632;
											assign node632 = (inp[0]) ? node638 : node633;
												assign node633 = (inp[6]) ? node635 : 8'b00001110;
													assign node635 = (inp[2]) ? 8'b00001110 : 8'b00011110;
												assign node638 = (inp[2]) ? node642 : node639;
													assign node639 = (inp[6]) ? 8'b00011110 : 8'b00001110;
													assign node642 = (inp[6]) ? 8'b00001110 : 8'b00011110;
											assign node645 = (inp[6]) ? 8'b00011111 : 8'b00001111;
								assign node648 = (inp[1]) ? node696 : node649;
									assign node649 = (inp[3]) ? node673 : node650;
										assign node650 = (inp[2]) ? node658 : node651;
											assign node651 = (inp[6]) ? node655 : node652;
												assign node652 = (inp[12]) ? 8'b00001110 : 8'b00011011;
												assign node655 = (inp[12]) ? 8'b00011110 : 8'b00001110;
											assign node658 = (inp[12]) ? node664 : node659;
												assign node659 = (inp[5]) ? 8'b00001011 : node660;
													assign node660 = (inp[6]) ? 8'b00011011 : 8'b00001011;
												assign node664 = (inp[5]) ? node668 : node665;
													assign node665 = (inp[6]) ? 8'b00001110 : 8'b00011011;
													assign node668 = (inp[6]) ? 8'b00011011 : node669;
														assign node669 = (inp[0]) ? 8'b00011011 : 8'b00001110;
										assign node673 = (inp[2]) ? node681 : node674;
											assign node674 = (inp[12]) ? node678 : node675;
												assign node675 = (inp[6]) ? 8'b00001111 : 8'b00011110;
												assign node678 = (inp[6]) ? 8'b00011111 : 8'b00001111;
											assign node681 = (inp[12]) ? node689 : node682;
												assign node682 = (inp[5]) ? 8'b00001110 : node683;
													assign node683 = (inp[0]) ? node685 : 8'b00011110;
														assign node685 = (inp[6]) ? 8'b00011110 : 8'b00001110;
												assign node689 = (inp[0]) ? 8'b00011110 : node690;
													assign node690 = (inp[6]) ? node692 : 8'b00001111;
														assign node692 = (inp[5]) ? 8'b00011110 : 8'b00001111;
									assign node696 = (inp[12]) ? node728 : node697;
										assign node697 = (inp[6]) ? node711 : node698;
											assign node698 = (inp[0]) ? node704 : node699;
												assign node699 = (inp[3]) ? node701 : 8'b00011011;
													assign node701 = (inp[5]) ? 8'b00011010 : 8'b00011011;
												assign node704 = (inp[2]) ? node706 : 8'b00011010;
													assign node706 = (inp[5]) ? 8'b00001010 : node707;
														assign node707 = (inp[3]) ? 8'b00001011 : 8'b00001010;
											assign node711 = (inp[2]) ? node719 : node712;
												assign node712 = (inp[0]) ? node714 : 8'b00001110;
													assign node714 = (inp[5]) ? 8'b00001011 : node715;
														assign node715 = (inp[3]) ? 8'b00001110 : 8'b00001011;
												assign node719 = (inp[5]) ? node723 : node720;
													assign node720 = (inp[0]) ? 8'b00011010 : 8'b00011011;
													assign node723 = (inp[0]) ? 8'b00001010 : node724;
														assign node724 = (inp[3]) ? 8'b00001010 : 8'b00001011;
										assign node728 = (inp[0]) ? node742 : node729;
											assign node729 = (inp[6]) ? node731 : 8'b00001110;
												assign node731 = (inp[5]) ? node735 : node732;
													assign node732 = (inp[2]) ? 8'b00001110 : 8'b00011110;
													assign node735 = (inp[2]) ? node739 : node736;
														assign node736 = (inp[3]) ? 8'b00011011 : 8'b00011110;
														assign node739 = (inp[3]) ? 8'b00011010 : 8'b00011011;
											assign node742 = (inp[3]) ? node748 : node743;
												assign node743 = (inp[6]) ? node745 : 8'b00001011;
													assign node745 = (inp[2]) ? 8'b00011010 : 8'b00011011;
												assign node748 = (inp[5]) ? node756 : node749;
													assign node749 = (inp[2]) ? node753 : node750;
														assign node750 = (inp[6]) ? 8'b00011110 : 8'b00001110;
														assign node753 = (inp[6]) ? 8'b00001110 : 8'b00011011;
													assign node756 = (inp[2]) ? 8'b00011010 : 8'b00001011;
						assign node759 = (inp[5]) ? node963 : node760;
							assign node760 = (inp[0]) ? node814 : node761;
								assign node761 = (inp[12]) ? node797 : node762;
									assign node762 = (inp[11]) ? node780 : node763;
										assign node763 = (inp[1]) ? node775 : node764;
											assign node764 = (inp[3]) ? node770 : node765;
												assign node765 = (inp[6]) ? node767 : 8'b10000010;
													assign node767 = (inp[2]) ? 8'b10000010 : 8'b00011010;
												assign node770 = (inp[6]) ? node772 : 8'b00001011;
													assign node772 = (inp[2]) ? 8'b00001011 : 8'b00011011;
											assign node775 = (inp[6]) ? node777 : 8'b10000010;
												assign node777 = (inp[2]) ? 8'b10000010 : 8'b00011010;
										assign node780 = (inp[2]) ? node792 : node781;
											assign node781 = (inp[6]) ? node787 : node782;
												assign node782 = (inp[3]) ? node784 : 8'b11110111;
													assign node784 = (inp[1]) ? 8'b11110111 : 8'b00011010;
												assign node787 = (inp[3]) ? node789 : 8'b00001010;
													assign node789 = (inp[1]) ? 8'b00001010 : 8'b00001011;
											assign node792 = (inp[3]) ? node794 : 8'b11110111;
												assign node794 = (inp[1]) ? 8'b11110111 : 8'b00011010;
									assign node797 = (inp[2]) ? node809 : node798;
										assign node798 = (inp[6]) ? node804 : node799;
											assign node799 = (inp[1]) ? 8'b00000010 : node800;
												assign node800 = (inp[3]) ? 8'b00001011 : 8'b00000010;
											assign node804 = (inp[1]) ? 8'b00011010 : node805;
												assign node805 = (inp[3]) ? 8'b00011011 : 8'b00011010;
										assign node809 = (inp[3]) ? node811 : 8'b00000010;
											assign node811 = (inp[1]) ? 8'b00000010 : 8'b00001011;
								assign node814 = (inp[10]) ? node896 : node815;
									assign node815 = (inp[11]) ? node843 : node816;
										assign node816 = (inp[6]) ? node828 : node817;
											assign node817 = (inp[2]) ? node823 : node818;
												assign node818 = (inp[3]) ? 8'b10000100 : node819;
													assign node819 = (inp[1]) ? 8'b10000101 : 8'b10000100;
												assign node823 = (inp[1]) ? node825 : 8'b10011101;
													assign node825 = (inp[3]) ? 8'b10010100 : 8'b10010101;
											assign node828 = (inp[2]) ? node836 : node829;
												assign node829 = (inp[1]) ? node833 : node830;
													assign node830 = (inp[3]) ? 8'b10011101 : 8'b10011100;
													assign node833 = (inp[3]) ? 8'b10011100 : 8'b10011101;
												assign node836 = (inp[1]) ? node840 : node837;
													assign node837 = (inp[3]) ? 8'b10001101 : 8'b10000100;
													assign node840 = (inp[3]) ? 8'b10000100 : 8'b10000101;
										assign node843 = (inp[3]) ? node873 : node844;
											assign node844 = (inp[6]) ? node860 : node845;
												assign node845 = (inp[1]) ? node853 : node846;
													assign node846 = (inp[2]) ? node850 : node847;
														assign node847 = (inp[12]) ? 8'b10100100 : 8'b10110001;
														assign node850 = (inp[12]) ? 8'b10110001 : 8'b10100001;
													assign node853 = (inp[2]) ? node857 : node854;
														assign node854 = (inp[12]) ? 8'b10100001 : 8'b10110000;
														assign node857 = (inp[12]) ? 8'b10110000 : 8'b10100000;
												assign node860 = (inp[2]) ? node868 : node861;
													assign node861 = (inp[1]) ? node865 : node862;
														assign node862 = (inp[12]) ? 8'b10111100 : 8'b10101100;
														assign node865 = (inp[12]) ? 8'b10111001 : 8'b10101001;
													assign node868 = (inp[12]) ? 8'b10100100 : node869;
														assign node869 = (inp[1]) ? 8'b10110000 : 8'b10110001;
											assign node873 = (inp[1]) ? node887 : node874;
												assign node874 = (inp[2]) ? node880 : node875;
													assign node875 = (inp[12]) ? 8'b10101101 : node876;
														assign node876 = (inp[6]) ? 8'b10101101 : 8'b10111100;
													assign node880 = (inp[6]) ? node884 : node881;
														assign node881 = (inp[12]) ? 8'b10111100 : 8'b10101100;
														assign node884 = (inp[12]) ? 8'b10101101 : 8'b10111100;
												assign node887 = (inp[6]) ? node889 : 8'b10110001;
													assign node889 = (inp[2]) ? node893 : node890;
														assign node890 = (inp[12]) ? 8'b10111100 : 8'b10101100;
														assign node893 = (inp[12]) ? 8'b10100100 : 8'b10110001;
									assign node896 = (inp[1]) ? node930 : node897;
										assign node897 = (inp[3]) ? node911 : node898;
											assign node898 = (inp[2]) ? node906 : node899;
												assign node899 = (inp[6]) ? node903 : node900;
													assign node900 = (inp[12]) ? 8'b00000010 : 8'b10000010;
													assign node903 = (inp[12]) ? 8'b00011010 : 8'b00001010;
												assign node906 = (inp[11]) ? node908 : 8'b10010000;
													assign node908 = (inp[12]) ? 8'b00000010 : 8'b11110111;
											assign node911 = (inp[11]) ? node921 : node912;
												assign node912 = (inp[12]) ? 8'b00001011 : node913;
													assign node913 = (inp[2]) ? node917 : node914;
														assign node914 = (inp[6]) ? 8'b00011011 : 8'b00001011;
														assign node917 = (inp[6]) ? 8'b00001011 : 8'b00011011;
												assign node921 = (inp[2]) ? 8'b00011010 : node922;
													assign node922 = (inp[12]) ? node926 : node923;
														assign node923 = (inp[6]) ? 8'b00001011 : 8'b00011010;
														assign node926 = (inp[6]) ? 8'b00011011 : 8'b00001011;
										assign node930 = (inp[3]) ? node946 : node931;
											assign node931 = (inp[11]) ? node937 : node932;
												assign node932 = (inp[2]) ? node934 : 8'b10011001;
													assign node934 = (inp[6]) ? 8'b10000001 : 8'b10010001;
												assign node937 = (inp[12]) ? node943 : node938;
													assign node938 = (inp[2]) ? node940 : 8'b10110100;
														assign node940 = (inp[6]) ? 8'b10110100 : 8'b10100100;
													assign node943 = (inp[2]) ? 8'b10100101 : 8'b11111101;
											assign node946 = (inp[6]) ? node956 : node947;
												assign node947 = (inp[2]) ? node953 : node948;
													assign node948 = (inp[12]) ? 8'b00000010 : node949;
														assign node949 = (inp[11]) ? 8'b11110111 : 8'b10000010;
													assign node953 = (inp[11]) ? 8'b11110101 : 8'b10010000;
												assign node956 = (inp[2]) ? node960 : node957;
													assign node957 = (inp[11]) ? 8'b00001010 : 8'b00011010;
													assign node960 = (inp[12]) ? 8'b00000010 : 8'b10000010;
							assign node963 = (inp[11]) ? node1035 : node964;
								assign node964 = (inp[6]) ? node994 : node965;
									assign node965 = (inp[3]) ? node979 : node966;
										assign node966 = (inp[0]) ? node972 : node967;
											assign node967 = (inp[10]) ? 8'b10000100 : node968;
												assign node968 = (inp[12]) ? 8'b00000010 : 8'b10000010;
											assign node972 = (inp[1]) ? node976 : node973;
												assign node973 = (inp[2]) ? 8'b10010100 : 8'b10000100;
												assign node976 = (inp[2]) ? 8'b10010101 : 8'b10000101;
										assign node979 = (inp[1]) ? node987 : node980;
											assign node980 = (inp[0]) ? node984 : node981;
												assign node981 = (inp[10]) ? 8'b10001101 : 8'b00001011;
												assign node984 = (inp[2]) ? 8'b10011101 : 8'b10001101;
											assign node987 = (inp[0]) ? node991 : node988;
												assign node988 = (inp[10]) ? 8'b10000101 : 8'b10000001;
												assign node991 = (inp[2]) ? 8'b10010101 : 8'b10000101;
									assign node994 = (inp[2]) ? node1014 : node995;
										assign node995 = (inp[10]) ? node1007 : node996;
											assign node996 = (inp[0]) ? node1002 : node997;
												assign node997 = (inp[3]) ? node999 : 8'b00011010;
													assign node999 = (inp[1]) ? 8'b10011001 : 8'b00011011;
												assign node1002 = (inp[3]) ? 8'b10011101 : node1003;
													assign node1003 = (inp[1]) ? 8'b10011101 : 8'b10011100;
											assign node1007 = (inp[3]) ? 8'b10011101 : node1008;
												assign node1008 = (inp[0]) ? node1010 : 8'b10011100;
													assign node1010 = (inp[1]) ? 8'b10011101 : 8'b10011100;
										assign node1014 = (inp[3]) ? node1022 : node1015;
											assign node1015 = (inp[0]) ? node1019 : node1016;
												assign node1016 = (inp[10]) ? 8'b10010100 : 8'b10010000;
												assign node1019 = (inp[1]) ? 8'b10010101 : 8'b10010100;
											assign node1022 = (inp[1]) ? node1030 : node1023;
												assign node1023 = (inp[12]) ? node1025 : 8'b10011101;
													assign node1025 = (inp[10]) ? 8'b10011101 : node1026;
														assign node1026 = (inp[0]) ? 8'b10011101 : 8'b00011011;
												assign node1030 = (inp[0]) ? 8'b10010101 : node1031;
													assign node1031 = (inp[10]) ? 8'b10010101 : 8'b10010001;
								assign node1035 = (inp[2]) ? node1105 : node1036;
									assign node1036 = (inp[6]) ? node1066 : node1037;
										assign node1037 = (inp[12]) ? node1055 : node1038;
											assign node1038 = (inp[3]) ? node1048 : node1039;
												assign node1039 = (inp[10]) ? node1043 : node1040;
													assign node1040 = (inp[0]) ? 8'b10110001 : 8'b11110111;
													assign node1043 = (inp[0]) ? node1045 : 8'b10110001;
														assign node1045 = (inp[1]) ? 8'b10110000 : 8'b10110001;
												assign node1048 = (inp[1]) ? node1050 : 8'b10111100;
													assign node1050 = (inp[0]) ? 8'b10110000 : node1051;
														assign node1051 = (inp[10]) ? 8'b10110000 : 8'b10110100;
											assign node1055 = (inp[3]) ? node1061 : node1056;
												assign node1056 = (inp[1]) ? node1058 : 8'b10100100;
													assign node1058 = (inp[0]) ? 8'b10100001 : 8'b10100100;
												assign node1061 = (inp[0]) ? 8'b10101101 : node1062;
													assign node1062 = (inp[10]) ? 8'b10101101 : 8'b00001011;
										assign node1066 = (inp[12]) ? node1082 : node1067;
											assign node1067 = (inp[10]) ? node1073 : node1068;
												assign node1068 = (inp[0]) ? 8'b10101001 : node1069;
													assign node1069 = (inp[1]) ? 8'b00001010 : 8'b00001011;
												assign node1073 = (inp[1]) ? node1077 : node1074;
													assign node1074 = (inp[3]) ? 8'b10101101 : 8'b10101100;
													assign node1077 = (inp[3]) ? 8'b10101001 : node1078;
														assign node1078 = (inp[0]) ? 8'b10101001 : 8'b10101100;
											assign node1082 = (inp[3]) ? node1094 : node1083;
												assign node1083 = (inp[10]) ? node1089 : node1084;
													assign node1084 = (inp[0]) ? node1086 : 8'b00011010;
														assign node1086 = (inp[1]) ? 8'b10111001 : 8'b10111100;
													assign node1089 = (inp[1]) ? node1091 : 8'b10111100;
														assign node1091 = (inp[0]) ? 8'b10111001 : 8'b10111100;
												assign node1094 = (inp[1]) ? node1100 : node1095;
													assign node1095 = (inp[10]) ? 8'b11111101 : node1096;
														assign node1096 = (inp[0]) ? 8'b11111101 : 8'b00011011;
													assign node1100 = (inp[10]) ? 8'b10111001 : node1101;
														assign node1101 = (inp[0]) ? 8'b10111001 : 8'b11111101;
									assign node1105 = (inp[3]) ? node1129 : node1106;
										assign node1106 = (inp[0]) ? node1122 : node1107;
											assign node1107 = (inp[10]) ? node1115 : node1108;
												assign node1108 = (inp[6]) ? node1112 : node1109;
													assign node1109 = (inp[12]) ? 8'b00000010 : 8'b11110111;
													assign node1112 = (inp[12]) ? 8'b11110101 : 8'b10100101;
												assign node1115 = (inp[6]) ? node1119 : node1116;
													assign node1116 = (inp[12]) ? 8'b10100100 : 8'b10110001;
													assign node1119 = (inp[12]) ? 8'b10110001 : 8'b10100001;
											assign node1122 = (inp[12]) ? node1126 : node1123;
												assign node1123 = (inp[1]) ? 8'b10100000 : 8'b10100001;
												assign node1126 = (inp[1]) ? 8'b10110000 : 8'b10110001;
										assign node1129 = (inp[1]) ? node1145 : node1130;
											assign node1130 = (inp[10]) ? node1140 : node1131;
												assign node1131 = (inp[0]) ? node1137 : node1132;
													assign node1132 = (inp[12]) ? 8'b00001011 : node1133;
														assign node1133 = (inp[6]) ? 8'b00001010 : 8'b00011010;
													assign node1137 = (inp[12]) ? 8'b10111100 : 8'b10101100;
												assign node1140 = (inp[12]) ? 8'b10111100 : node1141;
													assign node1141 = (inp[6]) ? 8'b10101100 : 8'b10111100;
											assign node1145 = (inp[12]) ? node1155 : node1146;
												assign node1146 = (inp[10]) ? node1150 : node1147;
													assign node1147 = (inp[0]) ? 8'b10100000 : 8'b10100100;
													assign node1150 = (inp[6]) ? 8'b10100000 : node1151;
														assign node1151 = (inp[0]) ? 8'b10100000 : 8'b10110000;
												assign node1155 = (inp[0]) ? 8'b10110000 : node1156;
													assign node1156 = (inp[6]) ? node1160 : node1157;
														assign node1157 = (inp[10]) ? 8'b10100001 : 8'b10100101;
														assign node1160 = (inp[10]) ? 8'b10110000 : 8'b10110100;
					assign node1164 = (inp[11]) ? node1410 : node1165;
						assign node1165 = (inp[3]) ? node1285 : node1166;
							assign node1166 = (inp[0]) ? node1190 : node1167;
								assign node1167 = (inp[10]) ? node1175 : node1168;
									assign node1168 = (inp[6]) ? node1170 : 8'b00101010;
										assign node1170 = (inp[5]) ? 8'b00111010 : node1171;
											assign node1171 = (inp[2]) ? 8'b00101010 : 8'b00111010;
									assign node1175 = (inp[6]) ? node1181 : node1176;
										assign node1176 = (inp[8]) ? node1178 : 8'b00101110;
											assign node1178 = (inp[5]) ? 8'b00101110 : 8'b00101010;
										assign node1181 = (inp[5]) ? 8'b00111110 : node1182;
											assign node1182 = (inp[2]) ? node1186 : node1183;
												assign node1183 = (inp[8]) ? 8'b00111010 : 8'b00111110;
												assign node1186 = (inp[8]) ? 8'b00101010 : 8'b00101110;
								assign node1190 = (inp[1]) ? node1236 : node1191;
									assign node1191 = (inp[10]) ? node1215 : node1192;
										assign node1192 = (inp[8]) ? node1202 : node1193;
											assign node1193 = (inp[6]) ? node1197 : node1194;
												assign node1194 = (inp[2]) ? 8'b00111010 : 8'b00101010;
												assign node1197 = (inp[5]) ? 8'b00111010 : node1198;
													assign node1198 = (inp[2]) ? 8'b00101010 : 8'b00111010;
											assign node1202 = (inp[5]) ? node1210 : node1203;
												assign node1203 = (inp[12]) ? 8'b00111110 : node1204;
													assign node1204 = (inp[6]) ? node1206 : 8'b00101110;
														assign node1206 = (inp[2]) ? 8'b00101110 : 8'b00111110;
												assign node1210 = (inp[6]) ? 8'b00111110 : node1211;
													assign node1211 = (inp[2]) ? 8'b00111110 : 8'b00101110;
										assign node1215 = (inp[5]) ? node1231 : node1216;
											assign node1216 = (inp[8]) ? node1224 : node1217;
												assign node1217 = (inp[6]) ? node1221 : node1218;
													assign node1218 = (inp[2]) ? 8'b00111110 : 8'b00101110;
													assign node1221 = (inp[2]) ? 8'b00101110 : 8'b00111110;
												assign node1224 = (inp[6]) ? node1228 : node1225;
													assign node1225 = (inp[2]) ? 8'b00111010 : 8'b00101010;
													assign node1228 = (inp[2]) ? 8'b00101010 : 8'b00111010;
											assign node1231 = (inp[6]) ? 8'b00111110 : node1232;
												assign node1232 = (inp[2]) ? 8'b00111110 : 8'b00101110;
									assign node1236 = (inp[5]) ? node1272 : node1237;
										assign node1237 = (inp[10]) ? node1255 : node1238;
											assign node1238 = (inp[8]) ? node1248 : node1239;
												assign node1239 = (inp[12]) ? node1241 : 8'b00111011;
													assign node1241 = (inp[6]) ? node1245 : node1242;
														assign node1242 = (inp[2]) ? 8'b00111011 : 8'b00101011;
														assign node1245 = (inp[2]) ? 8'b00101011 : 8'b00111011;
												assign node1248 = (inp[2]) ? node1252 : node1249;
													assign node1249 = (inp[6]) ? 8'b01111111 : 8'b00101111;
													assign node1252 = (inp[6]) ? 8'b00101111 : 8'b01111111;
											assign node1255 = (inp[8]) ? node1265 : node1256;
												assign node1256 = (inp[12]) ? 8'b01111111 : node1257;
													assign node1257 = (inp[6]) ? node1261 : node1258;
														assign node1258 = (inp[2]) ? 8'b01111111 : 8'b00101111;
														assign node1261 = (inp[2]) ? 8'b00101111 : 8'b01111111;
												assign node1265 = (inp[6]) ? node1269 : node1266;
													assign node1266 = (inp[2]) ? 8'b00111011 : 8'b00101011;
													assign node1269 = (inp[2]) ? 8'b00101011 : 8'b00111011;
										assign node1272 = (inp[8]) ? node1280 : node1273;
											assign node1273 = (inp[10]) ? 8'b01111111 : node1274;
												assign node1274 = (inp[6]) ? 8'b00111011 : node1275;
													assign node1275 = (inp[2]) ? 8'b00111011 : 8'b00101011;
											assign node1280 = (inp[2]) ? 8'b01111111 : node1281;
												assign node1281 = (inp[6]) ? 8'b01111111 : 8'b00101111;
							assign node1285 = (inp[5]) ? node1387 : node1286;
								assign node1286 = (inp[1]) ? node1338 : node1287;
									assign node1287 = (inp[0]) ? node1301 : node1288;
										assign node1288 = (inp[8]) ? node1296 : node1289;
											assign node1289 = (inp[10]) ? 8'b00101111 : node1290;
												assign node1290 = (inp[6]) ? node1292 : 8'b00101011;
													assign node1292 = (inp[2]) ? 8'b00101011 : 8'b00111011;
											assign node1296 = (inp[6]) ? node1298 : 8'b00101011;
												assign node1298 = (inp[2]) ? 8'b00101011 : 8'b00111011;
										assign node1301 = (inp[8]) ? node1325 : node1302;
											assign node1302 = (inp[10]) ? node1318 : node1303;
												assign node1303 = (inp[12]) ? node1311 : node1304;
													assign node1304 = (inp[6]) ? node1308 : node1305;
														assign node1305 = (inp[2]) ? 8'b00111011 : 8'b00101011;
														assign node1308 = (inp[2]) ? 8'b00101011 : 8'b00111011;
													assign node1311 = (inp[2]) ? node1315 : node1312;
														assign node1312 = (inp[6]) ? 8'b00111011 : 8'b00101011;
														assign node1315 = (inp[6]) ? 8'b00101011 : 8'b00111011;
												assign node1318 = (inp[12]) ? node1320 : 8'b01111111;
													assign node1320 = (inp[6]) ? node1322 : 8'b00101111;
														assign node1322 = (inp[2]) ? 8'b00101111 : 8'b01111111;
											assign node1325 = (inp[10]) ? node1333 : node1326;
												assign node1326 = (inp[6]) ? node1330 : node1327;
													assign node1327 = (inp[2]) ? 8'b01111111 : 8'b00101111;
													assign node1330 = (inp[2]) ? 8'b00101111 : 8'b01111111;
												assign node1333 = (inp[2]) ? node1335 : 8'b00101011;
													assign node1335 = (inp[6]) ? 8'b00101011 : 8'b00111011;
									assign node1338 = (inp[0]) ? node1356 : node1339;
										assign node1339 = (inp[10]) ? node1345 : node1340;
											assign node1340 = (inp[6]) ? node1342 : 8'b00101010;
												assign node1342 = (inp[2]) ? 8'b00101010 : 8'b00111010;
											assign node1345 = (inp[8]) ? node1351 : node1346;
												assign node1346 = (inp[2]) ? 8'b00101110 : node1347;
													assign node1347 = (inp[6]) ? 8'b00111110 : 8'b00101110;
												assign node1351 = (inp[2]) ? 8'b00101010 : node1352;
													assign node1352 = (inp[6]) ? 8'b00111010 : 8'b00101010;
										assign node1356 = (inp[8]) ? node1372 : node1357;
											assign node1357 = (inp[10]) ? node1365 : node1358;
												assign node1358 = (inp[2]) ? node1362 : node1359;
													assign node1359 = (inp[6]) ? 8'b00111010 : 8'b00101010;
													assign node1362 = (inp[6]) ? 8'b00101010 : 8'b00111010;
												assign node1365 = (inp[2]) ? node1369 : node1366;
													assign node1366 = (inp[6]) ? 8'b00111110 : 8'b00101110;
													assign node1369 = (inp[6]) ? 8'b00101110 : 8'b00111110;
											assign node1372 = (inp[10]) ? node1380 : node1373;
												assign node1373 = (inp[2]) ? node1377 : node1374;
													assign node1374 = (inp[6]) ? 8'b00111110 : 8'b00101110;
													assign node1377 = (inp[6]) ? 8'b00101110 : 8'b00111110;
												assign node1380 = (inp[2]) ? node1384 : node1381;
													assign node1381 = (inp[6]) ? 8'b00111010 : 8'b00101010;
													assign node1384 = (inp[6]) ? 8'b00101010 : 8'b00111010;
								assign node1387 = (inp[6]) ? node1403 : node1388;
									assign node1388 = (inp[10]) ? node1398 : node1389;
										assign node1389 = (inp[0]) ? node1391 : 8'b00101011;
											assign node1391 = (inp[8]) ? node1395 : node1392;
												assign node1392 = (inp[2]) ? 8'b00111011 : 8'b00101011;
												assign node1395 = (inp[2]) ? 8'b01111111 : 8'b00101111;
										assign node1398 = (inp[2]) ? node1400 : 8'b00101111;
											assign node1400 = (inp[0]) ? 8'b01111111 : 8'b00101111;
									assign node1403 = (inp[10]) ? 8'b01111111 : node1404;
										assign node1404 = (inp[0]) ? node1406 : 8'b00111011;
											assign node1406 = (inp[8]) ? 8'b01111111 : 8'b00111011;
						assign node1410 = (inp[8]) ? node1644 : node1411;
							assign node1411 = (inp[10]) ? node1535 : node1412;
								assign node1412 = (inp[1]) ? node1452 : node1413;
									assign node1413 = (inp[3]) ? node1433 : node1414;
										assign node1414 = (inp[2]) ? node1422 : node1415;
											assign node1415 = (inp[12]) ? node1419 : node1416;
												assign node1416 = (inp[6]) ? 8'b00101010 : 8'b00011111;
												assign node1419 = (inp[6]) ? 8'b00111010 : 8'b00101010;
											assign node1422 = (inp[0]) ? node1424 : 8'b00011111;
												assign node1424 = (inp[12]) ? node1430 : node1425;
													assign node1425 = (inp[6]) ? node1427 : 8'b00001111;
														assign node1427 = (inp[5]) ? 8'b00001111 : 8'b00011111;
													assign node1430 = (inp[6]) ? 8'b00101010 : 8'b00011111;
										assign node1433 = (inp[2]) ? node1441 : node1434;
											assign node1434 = (inp[6]) ? node1438 : node1435;
												assign node1435 = (inp[12]) ? 8'b00101011 : 8'b00111010;
												assign node1438 = (inp[12]) ? 8'b00111011 : 8'b00101011;
											assign node1441 = (inp[12]) ? node1447 : node1442;
												assign node1442 = (inp[5]) ? 8'b00101010 : node1443;
													assign node1443 = (inp[6]) ? 8'b00111010 : 8'b00101010;
												assign node1447 = (inp[0]) ? 8'b00111010 : node1448;
													assign node1448 = (inp[6]) ? 8'b00111010 : 8'b00101011;
									assign node1452 = (inp[5]) ? node1494 : node1453;
										assign node1453 = (inp[12]) ? node1473 : node1454;
											assign node1454 = (inp[6]) ? node1464 : node1455;
												assign node1455 = (inp[0]) ? node1457 : 8'b00011111;
													assign node1457 = (inp[2]) ? node1461 : node1458;
														assign node1458 = (inp[3]) ? 8'b00011111 : 8'b00011110;
														assign node1461 = (inp[3]) ? 8'b00001111 : 8'b00001110;
												assign node1464 = (inp[2]) ? node1470 : node1465;
													assign node1465 = (inp[0]) ? node1467 : 8'b00101010;
														assign node1467 = (inp[3]) ? 8'b00101010 : 8'b00001111;
													assign node1470 = (inp[0]) ? 8'b00011110 : 8'b00011111;
											assign node1473 = (inp[0]) ? node1479 : node1474;
												assign node1474 = (inp[6]) ? node1476 : 8'b00101010;
													assign node1476 = (inp[2]) ? 8'b00101010 : 8'b00111010;
												assign node1479 = (inp[3]) ? node1487 : node1480;
													assign node1480 = (inp[6]) ? node1484 : node1481;
														assign node1481 = (inp[2]) ? 8'b00011110 : 8'b00001111;
														assign node1484 = (inp[2]) ? 8'b00001111 : 8'b00011111;
													assign node1487 = (inp[6]) ? node1491 : node1488;
														assign node1488 = (inp[2]) ? 8'b00011111 : 8'b00101010;
														assign node1491 = (inp[2]) ? 8'b00101010 : 8'b00111010;
										assign node1494 = (inp[2]) ? node1520 : node1495;
											assign node1495 = (inp[0]) ? node1509 : node1496;
												assign node1496 = (inp[3]) ? node1502 : node1497;
													assign node1497 = (inp[12]) ? node1499 : 8'b00011111;
														assign node1499 = (inp[6]) ? 8'b00111010 : 8'b00101010;
													assign node1502 = (inp[6]) ? node1506 : node1503;
														assign node1503 = (inp[12]) ? 8'b00001111 : 8'b00011110;
														assign node1506 = (inp[12]) ? 8'b00011111 : 8'b00001111;
												assign node1509 = (inp[3]) ? node1515 : node1510;
													assign node1510 = (inp[6]) ? node1512 : 8'b00001111;
														assign node1512 = (inp[12]) ? 8'b00011111 : 8'b00001111;
													assign node1515 = (inp[12]) ? 8'b00001111 : node1516;
														assign node1516 = (inp[6]) ? 8'b00001111 : 8'b00011110;
											assign node1520 = (inp[0]) ? node1532 : node1521;
												assign node1521 = (inp[3]) ? node1527 : node1522;
													assign node1522 = (inp[12]) ? node1524 : 8'b00011111;
														assign node1524 = (inp[6]) ? 8'b00011111 : 8'b00101010;
													assign node1527 = (inp[6]) ? node1529 : 8'b00001111;
														assign node1529 = (inp[12]) ? 8'b00011110 : 8'b00001110;
												assign node1532 = (inp[12]) ? 8'b00011110 : 8'b00001110;
								assign node1535 = (inp[1]) ? node1581 : node1536;
									assign node1536 = (inp[3]) ? node1558 : node1537;
										assign node1537 = (inp[2]) ? node1545 : node1538;
											assign node1538 = (inp[12]) ? node1542 : node1539;
												assign node1539 = (inp[6]) ? 8'b00101110 : 8'b00111011;
												assign node1542 = (inp[6]) ? 8'b00111110 : 8'b00101110;
											assign node1545 = (inp[12]) ? node1553 : node1546;
												assign node1546 = (inp[5]) ? node1548 : 8'b00111011;
													assign node1548 = (inp[0]) ? 8'b00101011 : node1549;
														assign node1549 = (inp[6]) ? 8'b00101011 : 8'b00111011;
												assign node1553 = (inp[0]) ? 8'b00111011 : node1554;
													assign node1554 = (inp[6]) ? 8'b00111011 : 8'b00101110;
										assign node1558 = (inp[12]) ? node1570 : node1559;
											assign node1559 = (inp[6]) ? node1565 : node1560;
												assign node1560 = (inp[2]) ? node1562 : 8'b00111110;
													assign node1562 = (inp[0]) ? 8'b00101110 : 8'b00111110;
												assign node1565 = (inp[2]) ? node1567 : 8'b00101111;
													assign node1567 = (inp[5]) ? 8'b00101110 : 8'b00111110;
											assign node1570 = (inp[2]) ? node1574 : node1571;
												assign node1571 = (inp[6]) ? 8'b01111111 : 8'b00101111;
												assign node1574 = (inp[5]) ? 8'b00111110 : node1575;
													assign node1575 = (inp[6]) ? 8'b00101111 : node1576;
														assign node1576 = (inp[0]) ? 8'b00111110 : 8'b00101111;
									assign node1581 = (inp[0]) ? node1617 : node1582;
										assign node1582 = (inp[12]) ? node1600 : node1583;
											assign node1583 = (inp[6]) ? node1589 : node1584;
												assign node1584 = (inp[5]) ? node1586 : 8'b00111011;
													assign node1586 = (inp[3]) ? 8'b00111010 : 8'b00111011;
												assign node1589 = (inp[2]) ? node1595 : node1590;
													assign node1590 = (inp[5]) ? node1592 : 8'b00101110;
														assign node1592 = (inp[3]) ? 8'b00101011 : 8'b00101110;
													assign node1595 = (inp[5]) ? node1597 : 8'b00111011;
														assign node1597 = (inp[3]) ? 8'b00101010 : 8'b00101011;
											assign node1600 = (inp[6]) ? node1606 : node1601;
												assign node1601 = (inp[5]) ? node1603 : 8'b00101110;
													assign node1603 = (inp[3]) ? 8'b00101011 : 8'b00101110;
												assign node1606 = (inp[5]) ? node1610 : node1607;
													assign node1607 = (inp[2]) ? 8'b00101110 : 8'b00111110;
													assign node1610 = (inp[3]) ? node1614 : node1611;
														assign node1611 = (inp[2]) ? 8'b00111011 : 8'b00111110;
														assign node1614 = (inp[2]) ? 8'b00111010 : 8'b00111011;
										assign node1617 = (inp[12]) ? node1633 : node1618;
											assign node1618 = (inp[2]) ? node1626 : node1619;
												assign node1619 = (inp[6]) ? 8'b00101011 : node1620;
													assign node1620 = (inp[3]) ? node1622 : 8'b00111010;
														assign node1622 = (inp[5]) ? 8'b00111010 : 8'b00111011;
												assign node1626 = (inp[5]) ? 8'b00101010 : node1627;
													assign node1627 = (inp[6]) ? 8'b00111010 : node1628;
														assign node1628 = (inp[3]) ? 8'b00101011 : 8'b00101010;
											assign node1633 = (inp[2]) ? node1639 : node1634;
												assign node1634 = (inp[6]) ? node1636 : 8'b00101011;
													assign node1636 = (inp[3]) ? 8'b00111110 : 8'b00111011;
												assign node1639 = (inp[5]) ? 8'b00111010 : node1640;
													assign node1640 = (inp[3]) ? 8'b00111011 : 8'b00101011;
							assign node1644 = (inp[5]) ? node1788 : node1645;
								assign node1645 = (inp[0]) ? node1679 : node1646;
									assign node1646 = (inp[12]) ? node1662 : node1647;
										assign node1647 = (inp[2]) ? node1657 : node1648;
											assign node1648 = (inp[6]) ? node1652 : node1649;
												assign node1649 = (inp[1]) ? 8'b00011111 : 8'b00111010;
												assign node1652 = (inp[3]) ? node1654 : 8'b00101010;
													assign node1654 = (inp[1]) ? 8'b00101010 : 8'b00101011;
											assign node1657 = (inp[3]) ? node1659 : 8'b00011111;
												assign node1659 = (inp[1]) ? 8'b00011111 : 8'b00111010;
										assign node1662 = (inp[6]) ? node1668 : node1663;
											assign node1663 = (inp[3]) ? node1665 : 8'b00101010;
												assign node1665 = (inp[1]) ? 8'b00101010 : 8'b00101011;
											assign node1668 = (inp[2]) ? node1674 : node1669;
												assign node1669 = (inp[3]) ? node1671 : 8'b00111010;
													assign node1671 = (inp[10]) ? 8'b00111010 : 8'b00111011;
												assign node1674 = (inp[3]) ? node1676 : 8'b00101010;
													assign node1676 = (inp[1]) ? 8'b00101010 : 8'b00101011;
									assign node1679 = (inp[10]) ? node1733 : node1680;
										assign node1680 = (inp[3]) ? node1712 : node1681;
											assign node1681 = (inp[1]) ? node1697 : node1682;
												assign node1682 = (inp[12]) ? node1690 : node1683;
													assign node1683 = (inp[6]) ? node1687 : node1684;
														assign node1684 = (inp[2]) ? 8'b00001011 : 8'b00011011;
														assign node1687 = (inp[2]) ? 8'b00011011 : 8'b00001110;
													assign node1690 = (inp[2]) ? node1694 : node1691;
														assign node1691 = (inp[6]) ? 8'b00011110 : 8'b00001110;
														assign node1694 = (inp[6]) ? 8'b00001110 : 8'b00011011;
												assign node1697 = (inp[12]) ? node1705 : node1698;
													assign node1698 = (inp[2]) ? node1702 : node1699;
														assign node1699 = (inp[6]) ? 8'b00001011 : 8'b00011010;
														assign node1702 = (inp[6]) ? 8'b00011010 : 8'b00001010;
													assign node1705 = (inp[6]) ? node1709 : node1706;
														assign node1706 = (inp[2]) ? 8'b00011010 : 8'b00001011;
														assign node1709 = (inp[2]) ? 8'b00001011 : 8'b00011011;
											assign node1712 = (inp[2]) ? node1720 : node1713;
												assign node1713 = (inp[1]) ? node1715 : 8'b00001111;
													assign node1715 = (inp[6]) ? node1717 : 8'b00001110;
														assign node1717 = (inp[12]) ? 8'b00011110 : 8'b00001110;
												assign node1720 = (inp[1]) ? node1728 : node1721;
													assign node1721 = (inp[6]) ? node1725 : node1722;
														assign node1722 = (inp[12]) ? 8'b00011110 : 8'b00001110;
														assign node1725 = (inp[12]) ? 8'b00001111 : 8'b00011110;
													assign node1728 = (inp[6]) ? node1730 : 8'b00011011;
														assign node1730 = (inp[12]) ? 8'b00001110 : 8'b00011011;
										assign node1733 = (inp[1]) ? node1765 : node1734;
											assign node1734 = (inp[3]) ? node1750 : node1735;
												assign node1735 = (inp[6]) ? node1743 : node1736;
													assign node1736 = (inp[12]) ? node1740 : node1737;
														assign node1737 = (inp[2]) ? 8'b00001111 : 8'b00011111;
														assign node1740 = (inp[2]) ? 8'b00011111 : 8'b00101010;
													assign node1743 = (inp[12]) ? node1747 : node1744;
														assign node1744 = (inp[2]) ? 8'b00011111 : 8'b00101010;
														assign node1747 = (inp[2]) ? 8'b00101010 : 8'b00111010;
												assign node1750 = (inp[12]) ? node1758 : node1751;
													assign node1751 = (inp[6]) ? node1755 : node1752;
														assign node1752 = (inp[2]) ? 8'b00101010 : 8'b00111010;
														assign node1755 = (inp[2]) ? 8'b00111010 : 8'b00101011;
													assign node1758 = (inp[2]) ? node1762 : node1759;
														assign node1759 = (inp[6]) ? 8'b00111011 : 8'b00101011;
														assign node1762 = (inp[6]) ? 8'b00101011 : 8'b00111010;
											assign node1765 = (inp[3]) ? node1775 : node1766;
												assign node1766 = (inp[12]) ? 8'b00001111 : node1767;
													assign node1767 = (inp[6]) ? node1771 : node1768;
														assign node1768 = (inp[2]) ? 8'b00001110 : 8'b00011110;
														assign node1771 = (inp[2]) ? 8'b00011110 : 8'b00001111;
												assign node1775 = (inp[6]) ? node1781 : node1776;
													assign node1776 = (inp[2]) ? node1778 : 8'b00011111;
														assign node1778 = (inp[12]) ? 8'b00011111 : 8'b00001111;
													assign node1781 = (inp[2]) ? node1785 : node1782;
														assign node1782 = (inp[12]) ? 8'b00111010 : 8'b00101010;
														assign node1785 = (inp[12]) ? 8'b00101010 : 8'b00011111;
								assign node1788 = (inp[1]) ? node1854 : node1789;
									assign node1789 = (inp[10]) ? node1825 : node1790;
										assign node1790 = (inp[0]) ? node1810 : node1791;
											assign node1791 = (inp[3]) ? node1803 : node1792;
												assign node1792 = (inp[12]) ? node1798 : node1793;
													assign node1793 = (inp[6]) ? node1795 : 8'b00011111;
														assign node1795 = (inp[2]) ? 8'b00001111 : 8'b00101010;
													assign node1798 = (inp[6]) ? node1800 : 8'b00101010;
														assign node1800 = (inp[2]) ? 8'b00011111 : 8'b00111010;
												assign node1803 = (inp[12]) ? node1807 : node1804;
													assign node1804 = (inp[2]) ? 8'b00101010 : 8'b00101011;
													assign node1807 = (inp[6]) ? 8'b00111011 : 8'b00101011;
											assign node1810 = (inp[6]) ? node1822 : node1811;
												assign node1811 = (inp[3]) ? node1817 : node1812;
													assign node1812 = (inp[12]) ? node1814 : 8'b00011011;
														assign node1814 = (inp[2]) ? 8'b00011011 : 8'b00001110;
													assign node1817 = (inp[2]) ? node1819 : 8'b00001111;
														assign node1819 = (inp[12]) ? 8'b00011110 : 8'b00001110;
												assign node1822 = (inp[12]) ? 8'b00011110 : 8'b00001110;
										assign node1825 = (inp[3]) ? node1843 : node1826;
											assign node1826 = (inp[2]) ? node1834 : node1827;
												assign node1827 = (inp[0]) ? 8'b00011110 : node1828;
													assign node1828 = (inp[12]) ? 8'b00001110 : node1829;
														assign node1829 = (inp[6]) ? 8'b00001110 : 8'b00011011;
												assign node1834 = (inp[12]) ? node1838 : node1835;
													assign node1835 = (inp[6]) ? 8'b00001011 : 8'b00011011;
													assign node1838 = (inp[0]) ? 8'b00011011 : node1839;
														assign node1839 = (inp[6]) ? 8'b00011011 : 8'b00001110;
											assign node1843 = (inp[2]) ? node1851 : node1844;
												assign node1844 = (inp[6]) ? node1848 : node1845;
													assign node1845 = (inp[12]) ? 8'b00001111 : 8'b00011110;
													assign node1848 = (inp[12]) ? 8'b00011111 : 8'b00001111;
												assign node1851 = (inp[0]) ? 8'b00001110 : 8'b00011110;
									assign node1854 = (inp[2]) ? node1888 : node1855;
										assign node1855 = (inp[0]) ? node1881 : node1856;
											assign node1856 = (inp[3]) ? node1868 : node1857;
												assign node1857 = (inp[10]) ? node1863 : node1858;
													assign node1858 = (inp[6]) ? 8'b00101010 : node1859;
														assign node1859 = (inp[12]) ? 8'b00101010 : 8'b00011111;
													assign node1863 = (inp[12]) ? 8'b00001110 : node1864;
														assign node1864 = (inp[6]) ? 8'b00001110 : 8'b00011011;
												assign node1868 = (inp[10]) ? node1876 : node1869;
													assign node1869 = (inp[12]) ? node1873 : node1870;
														assign node1870 = (inp[6]) ? 8'b00001111 : 8'b00011110;
														assign node1873 = (inp[6]) ? 8'b00011111 : 8'b00001111;
													assign node1876 = (inp[12]) ? node1878 : 8'b00001011;
														assign node1878 = (inp[6]) ? 8'b00011011 : 8'b00001011;
											assign node1881 = (inp[12]) ? node1885 : node1882;
												assign node1882 = (inp[6]) ? 8'b00001011 : 8'b00011010;
												assign node1885 = (inp[6]) ? 8'b00011011 : 8'b00001011;
										assign node1888 = (inp[0]) ? node1916 : node1889;
											assign node1889 = (inp[10]) ? node1901 : node1890;
												assign node1890 = (inp[3]) ? node1896 : node1891;
													assign node1891 = (inp[6]) ? node1893 : 8'b00101010;
														assign node1893 = (inp[12]) ? 8'b00011111 : 8'b00001111;
													assign node1896 = (inp[12]) ? 8'b00011110 : node1897;
														assign node1897 = (inp[6]) ? 8'b00001110 : 8'b00011110;
												assign node1901 = (inp[3]) ? node1909 : node1902;
													assign node1902 = (inp[6]) ? node1906 : node1903;
														assign node1903 = (inp[12]) ? 8'b00001110 : 8'b00011011;
														assign node1906 = (inp[12]) ? 8'b00011011 : 8'b00001011;
													assign node1909 = (inp[6]) ? node1913 : node1910;
														assign node1910 = (inp[12]) ? 8'b00001011 : 8'b00011010;
														assign node1913 = (inp[12]) ? 8'b00011010 : 8'b00001010;
											assign node1916 = (inp[12]) ? 8'b00011010 : 8'b00001010;
			assign node1919 = (inp[5]) ? node3031 : node1920;
				assign node1920 = (inp[0]) ? node2120 : node1921;
					assign node1921 = (inp[8]) ? node2049 : node1922;
						assign node1922 = (inp[4]) ? node1946 : node1923;
							assign node1923 = (inp[1]) ? node1935 : node1924;
								assign node1924 = (inp[2]) ? node1930 : node1925;
									assign node1925 = (inp[12]) ? 8'b00011111 : node1926;
										assign node1926 = (inp[11]) ? 8'b00001111 : 8'b00011111;
									assign node1930 = (inp[11]) ? node1932 : 8'b00001111;
										assign node1932 = (inp[12]) ? 8'b00001111 : 8'b00011110;
								assign node1935 = (inp[2]) ? node1941 : node1936;
									assign node1936 = (inp[12]) ? 8'b00011110 : node1937;
										assign node1937 = (inp[11]) ? 8'b00001110 : 8'b00011110;
									assign node1941 = (inp[11]) ? node1943 : 8'b00001110;
										assign node1943 = (inp[12]) ? 8'b00001110 : 8'b00011011;
							assign node1946 = (inp[10]) ? node1998 : node1947;
								assign node1947 = (inp[12]) ? node1981 : node1948;
									assign node1948 = (inp[11]) ? node1964 : node1949;
										assign node1949 = (inp[2]) ? node1959 : node1950;
											assign node1950 = (inp[6]) ? node1954 : node1951;
												assign node1951 = (inp[3]) ? 8'b00001011 : 8'b10000010;
												assign node1954 = (inp[3]) ? node1956 : 8'b00011010;
													assign node1956 = (inp[1]) ? 8'b00011010 : 8'b00011011;
											assign node1959 = (inp[3]) ? node1961 : 8'b10000010;
												assign node1961 = (inp[1]) ? 8'b10000010 : 8'b00001011;
										assign node1964 = (inp[6]) ? node1970 : node1965;
											assign node1965 = (inp[1]) ? 8'b11110111 : node1966;
												assign node1966 = (inp[3]) ? 8'b00011010 : 8'b11110111;
											assign node1970 = (inp[2]) ? node1976 : node1971;
												assign node1971 = (inp[1]) ? 8'b00001010 : node1972;
													assign node1972 = (inp[3]) ? 8'b00001011 : 8'b00001010;
												assign node1976 = (inp[3]) ? node1978 : 8'b11110111;
													assign node1978 = (inp[1]) ? 8'b11110111 : 8'b00011010;
									assign node1981 = (inp[6]) ? node1987 : node1982;
										assign node1982 = (inp[1]) ? 8'b00000010 : node1983;
											assign node1983 = (inp[3]) ? 8'b00001011 : 8'b00000010;
										assign node1987 = (inp[2]) ? node1993 : node1988;
											assign node1988 = (inp[3]) ? node1990 : 8'b00011010;
												assign node1990 = (inp[1]) ? 8'b00011010 : 8'b00011011;
											assign node1993 = (inp[3]) ? node1995 : 8'b00000010;
												assign node1995 = (inp[1]) ? 8'b00000010 : 8'b00001011;
								assign node1998 = (inp[3]) ? node2016 : node1999;
									assign node1999 = (inp[12]) ? node2011 : node2000;
										assign node2000 = (inp[11]) ? node2006 : node2001;
											assign node2001 = (inp[6]) ? node2003 : 8'b00001110;
												assign node2003 = (inp[2]) ? 8'b00001110 : 8'b00011110;
											assign node2006 = (inp[2]) ? 8'b00011011 : node2007;
												assign node2007 = (inp[6]) ? 8'b00001110 : 8'b00011011;
										assign node2011 = (inp[2]) ? 8'b00001110 : node2012;
											assign node2012 = (inp[6]) ? 8'b00011110 : 8'b00001110;
									assign node2016 = (inp[1]) ? node2032 : node2017;
										assign node2017 = (inp[6]) ? node2023 : node2018;
											assign node2018 = (inp[11]) ? node2020 : 8'b00001111;
												assign node2020 = (inp[12]) ? 8'b00001111 : 8'b00011110;
											assign node2023 = (inp[11]) ? node2025 : 8'b00011111;
												assign node2025 = (inp[12]) ? node2029 : node2026;
													assign node2026 = (inp[2]) ? 8'b00011110 : 8'b00001111;
													assign node2029 = (inp[2]) ? 8'b00001111 : 8'b00011111;
										assign node2032 = (inp[2]) ? node2044 : node2033;
											assign node2033 = (inp[6]) ? node2039 : node2034;
												assign node2034 = (inp[11]) ? node2036 : 8'b00001110;
													assign node2036 = (inp[12]) ? 8'b00001110 : 8'b00011011;
												assign node2039 = (inp[11]) ? node2041 : 8'b00011110;
													assign node2041 = (inp[12]) ? 8'b00011110 : 8'b00001110;
											assign node2044 = (inp[11]) ? node2046 : 8'b00001110;
												assign node2046 = (inp[12]) ? 8'b00001110 : 8'b00011011;
						assign node2049 = (inp[1]) ? node2097 : node2050;
							assign node2050 = (inp[4]) ? node2062 : node2051;
								assign node2051 = (inp[2]) ? node2057 : node2052;
									assign node2052 = (inp[11]) ? node2054 : 8'b00011011;
										assign node2054 = (inp[12]) ? 8'b00011011 : 8'b00001011;
									assign node2057 = (inp[11]) ? node2059 : 8'b00001011;
										assign node2059 = (inp[12]) ? 8'b00001011 : 8'b00011010;
								assign node2062 = (inp[3]) ? node2080 : node2063;
									assign node2063 = (inp[12]) ? node2075 : node2064;
										assign node2064 = (inp[11]) ? node2070 : node2065;
											assign node2065 = (inp[6]) ? node2067 : 8'b10000010;
												assign node2067 = (inp[2]) ? 8'b10000010 : 8'b00011010;
											assign node2070 = (inp[6]) ? node2072 : 8'b11110111;
												assign node2072 = (inp[2]) ? 8'b11110111 : 8'b00001010;
										assign node2075 = (inp[2]) ? 8'b00000010 : node2076;
											assign node2076 = (inp[6]) ? 8'b00011010 : 8'b00000010;
									assign node2080 = (inp[12]) ? node2092 : node2081;
										assign node2081 = (inp[11]) ? node2087 : node2082;
											assign node2082 = (inp[2]) ? 8'b00001011 : node2083;
												assign node2083 = (inp[6]) ? 8'b00011011 : 8'b00001011;
											assign node2087 = (inp[6]) ? node2089 : 8'b00011010;
												assign node2089 = (inp[2]) ? 8'b00011010 : 8'b00001011;
										assign node2092 = (inp[2]) ? 8'b00001011 : node2093;
											assign node2093 = (inp[6]) ? 8'b00011011 : 8'b00001011;
							assign node2097 = (inp[2]) ? node2115 : node2098;
								assign node2098 = (inp[6]) ? node2110 : node2099;
									assign node2099 = (inp[4]) ? node2105 : node2100;
										assign node2100 = (inp[12]) ? 8'b00011010 : node2101;
											assign node2101 = (inp[11]) ? 8'b00001010 : 8'b00011010;
										assign node2105 = (inp[12]) ? 8'b00000010 : node2106;
											assign node2106 = (inp[11]) ? 8'b11110111 : 8'b10000010;
									assign node2110 = (inp[11]) ? node2112 : 8'b00011010;
										assign node2112 = (inp[12]) ? 8'b00011010 : 8'b00001010;
								assign node2115 = (inp[12]) ? 8'b00000010 : node2116;
									assign node2116 = (inp[11]) ? 8'b11110111 : 8'b10000010;
					assign node2120 = (inp[9]) ? node2590 : node2121;
						assign node2121 = (inp[11]) ? node2309 : node2122;
							assign node2122 = (inp[4]) ? node2176 : node2123;
								assign node2123 = (inp[8]) ? node2141 : node2124;
									assign node2124 = (inp[1]) ? node2130 : node2125;
										assign node2125 = (inp[2]) ? node2127 : 8'b11111101;
											assign node2127 = (inp[6]) ? 8'b10101101 : 8'b11111101;
										assign node2130 = (inp[3]) ? node2136 : node2131;
											assign node2131 = (inp[6]) ? node2133 : 8'b11111101;
												assign node2133 = (inp[2]) ? 8'b10101101 : 8'b11111101;
											assign node2136 = (inp[6]) ? node2138 : 8'b10111100;
												assign node2138 = (inp[2]) ? 8'b10101100 : 8'b10111100;
									assign node2141 = (inp[10]) ? node2159 : node2142;
										assign node2142 = (inp[2]) ? node2148 : node2143;
											assign node2143 = (inp[3]) ? node2145 : 8'b11111101;
												assign node2145 = (inp[1]) ? 8'b10111100 : 8'b11111101;
											assign node2148 = (inp[1]) ? node2152 : node2149;
												assign node2149 = (inp[6]) ? 8'b10101101 : 8'b11111101;
												assign node2152 = (inp[3]) ? node2156 : node2153;
													assign node2153 = (inp[12]) ? 8'b10100101 : 8'b11110101;
													assign node2156 = (inp[6]) ? 8'b10100100 : 8'b10110100;
										assign node2159 = (inp[2]) ? node2165 : node2160;
											assign node2160 = (inp[3]) ? node2162 : 8'b10111001;
												assign node2162 = (inp[1]) ? 8'b10111000 : 8'b10111001;
											assign node2165 = (inp[1]) ? node2169 : node2166;
												assign node2166 = (inp[6]) ? 8'b10101001 : 8'b10111001;
												assign node2169 = (inp[6]) ? node2173 : node2170;
													assign node2170 = (inp[3]) ? 8'b10110000 : 8'b10110001;
													assign node2173 = (inp[3]) ? 8'b10100000 : 8'b10100001;
								assign node2176 = (inp[3]) ? node2236 : node2177;
									assign node2177 = (inp[1]) ? node2209 : node2178;
										assign node2178 = (inp[10]) ? node2196 : node2179;
											assign node2179 = (inp[8]) ? node2189 : node2180;
												assign node2180 = (inp[12]) ? 8'b10100000 : node2181;
													assign node2181 = (inp[2]) ? node2185 : node2182;
														assign node2182 = (inp[6]) ? 8'b10111000 : 8'b10100000;
														assign node2185 = (inp[6]) ? 8'b10100000 : 8'b10110000;
												assign node2189 = (inp[6]) ? node2193 : node2190;
													assign node2190 = (inp[2]) ? 8'b10110100 : 8'b10100100;
													assign node2193 = (inp[2]) ? 8'b10100100 : 8'b10111100;
											assign node2196 = (inp[8]) ? node2204 : node2197;
												assign node2197 = (inp[6]) ? node2201 : node2198;
													assign node2198 = (inp[2]) ? 8'b10111100 : 8'b10101100;
													assign node2201 = (inp[2]) ? 8'b10101100 : 8'b10111100;
												assign node2204 = (inp[12]) ? node2206 : 8'b10100000;
													assign node2206 = (inp[6]) ? 8'b10111000 : 8'b10110000;
										assign node2209 = (inp[2]) ? node2225 : node2210;
											assign node2210 = (inp[6]) ? node2218 : node2211;
												assign node2211 = (inp[8]) ? node2215 : node2212;
													assign node2212 = (inp[10]) ? 8'b10101101 : 8'b10100001;
													assign node2215 = (inp[10]) ? 8'b10100001 : 8'b10100101;
												assign node2218 = (inp[8]) ? node2222 : node2219;
													assign node2219 = (inp[10]) ? 8'b11111101 : 8'b10111001;
													assign node2222 = (inp[10]) ? 8'b10111001 : 8'b11111101;
											assign node2225 = (inp[6]) ? node2231 : node2226;
												assign node2226 = (inp[10]) ? 8'b11111101 : node2227;
													assign node2227 = (inp[8]) ? 8'b11110101 : 8'b10110001;
												assign node2231 = (inp[10]) ? 8'b10100001 : node2232;
													assign node2232 = (inp[8]) ? 8'b10100101 : 8'b10100001;
									assign node2236 = (inp[1]) ? node2276 : node2237;
										assign node2237 = (inp[6]) ? node2253 : node2238;
											assign node2238 = (inp[2]) ? node2246 : node2239;
												assign node2239 = (inp[8]) ? node2243 : node2240;
													assign node2240 = (inp[10]) ? 8'b10101101 : 8'b10101001;
													assign node2243 = (inp[10]) ? 8'b10101001 : 8'b10101101;
												assign node2246 = (inp[8]) ? node2250 : node2247;
													assign node2247 = (inp[10]) ? 8'b11111101 : 8'b10111001;
													assign node2250 = (inp[10]) ? 8'b10111001 : 8'b11111101;
											assign node2253 = (inp[2]) ? node2267 : node2254;
												assign node2254 = (inp[12]) ? node2262 : node2255;
													assign node2255 = (inp[8]) ? node2259 : node2256;
														assign node2256 = (inp[10]) ? 8'b11111101 : 8'b10111001;
														assign node2259 = (inp[10]) ? 8'b10111001 : 8'b11111101;
													assign node2262 = (inp[10]) ? 8'b10111001 : node2263;
														assign node2263 = (inp[8]) ? 8'b11111101 : 8'b10111001;
												assign node2267 = (inp[12]) ? 8'b10101101 : node2268;
													assign node2268 = (inp[8]) ? node2272 : node2269;
														assign node2269 = (inp[10]) ? 8'b10101101 : 8'b10101001;
														assign node2272 = (inp[10]) ? 8'b10101001 : 8'b10101101;
										assign node2276 = (inp[6]) ? node2296 : node2277;
											assign node2277 = (inp[2]) ? node2289 : node2278;
												assign node2278 = (inp[12]) ? node2284 : node2279;
													assign node2279 = (inp[8]) ? 8'b10100000 : node2280;
														assign node2280 = (inp[10]) ? 8'b10101100 : 8'b10100000;
													assign node2284 = (inp[10]) ? 8'b10100000 : node2285;
														assign node2285 = (inp[8]) ? 8'b10100100 : 8'b10100000;
												assign node2289 = (inp[10]) ? node2293 : node2290;
													assign node2290 = (inp[12]) ? 8'b10110100 : 8'b10110000;
													assign node2293 = (inp[8]) ? 8'b10110000 : 8'b10111100;
											assign node2296 = (inp[2]) ? node2304 : node2297;
												assign node2297 = (inp[8]) ? node2301 : node2298;
													assign node2298 = (inp[10]) ? 8'b10111100 : 8'b10111000;
													assign node2301 = (inp[10]) ? 8'b10111000 : 8'b10111100;
												assign node2304 = (inp[8]) ? 8'b10100000 : node2305;
													assign node2305 = (inp[10]) ? 8'b10101100 : 8'b10100000;
							assign node2309 = (inp[8]) ? node2443 : node2310;
								assign node2310 = (inp[4]) ? node2346 : node2311;
									assign node2311 = (inp[1]) ? node2323 : node2312;
										assign node2312 = (inp[2]) ? node2316 : node2313;
											assign node2313 = (inp[12]) ? 8'b11111101 : 8'b10101101;
											assign node2316 = (inp[12]) ? node2320 : node2317;
												assign node2317 = (inp[6]) ? 8'b10111100 : 8'b10101100;
												assign node2320 = (inp[6]) ? 8'b10101101 : 8'b10111100;
										assign node2323 = (inp[3]) ? node2335 : node2324;
											assign node2324 = (inp[2]) ? node2328 : node2325;
												assign node2325 = (inp[12]) ? 8'b10111001 : 8'b10101001;
												assign node2328 = (inp[12]) ? node2332 : node2329;
													assign node2329 = (inp[6]) ? 8'b10111000 : 8'b10101000;
													assign node2332 = (inp[6]) ? 8'b10101001 : 8'b10111000;
											assign node2335 = (inp[2]) ? node2339 : node2336;
												assign node2336 = (inp[12]) ? 8'b10111100 : 8'b10101100;
												assign node2339 = (inp[12]) ? node2343 : node2340;
													assign node2340 = (inp[6]) ? 8'b10111001 : 8'b10101001;
													assign node2343 = (inp[6]) ? 8'b10101100 : 8'b10111001;
									assign node2346 = (inp[10]) ? node2400 : node2347;
										assign node2347 = (inp[1]) ? node2375 : node2348;
											assign node2348 = (inp[3]) ? node2362 : node2349;
												assign node2349 = (inp[6]) ? node2357 : node2350;
													assign node2350 = (inp[12]) ? node2354 : node2351;
														assign node2351 = (inp[2]) ? 8'b10000101 : 8'b10010101;
														assign node2354 = (inp[2]) ? 8'b10010101 : 8'b10100000;
													assign node2357 = (inp[2]) ? 8'b10100000 : node2358;
														assign node2358 = (inp[12]) ? 8'b10111000 : 8'b10101000;
												assign node2362 = (inp[2]) ? node2370 : node2363;
													assign node2363 = (inp[6]) ? node2367 : node2364;
														assign node2364 = (inp[12]) ? 8'b10101001 : 8'b10111000;
														assign node2367 = (inp[12]) ? 8'b10111001 : 8'b10101001;
													assign node2370 = (inp[6]) ? 8'b10111000 : node2371;
														assign node2371 = (inp[12]) ? 8'b10111000 : 8'b10101000;
											assign node2375 = (inp[3]) ? node2387 : node2376;
												assign node2376 = (inp[6]) ? node2384 : node2377;
													assign node2377 = (inp[2]) ? node2381 : node2378;
														assign node2378 = (inp[12]) ? 8'b10000101 : 8'b10010100;
														assign node2381 = (inp[12]) ? 8'b10010100 : 8'b10000100;
													assign node2384 = (inp[2]) ? 8'b10000101 : 8'b10011101;
												assign node2387 = (inp[12]) ? node2395 : node2388;
													assign node2388 = (inp[2]) ? node2392 : node2389;
														assign node2389 = (inp[6]) ? 8'b10101000 : 8'b10010101;
														assign node2392 = (inp[6]) ? 8'b10010101 : 8'b10000101;
													assign node2395 = (inp[6]) ? node2397 : 8'b10100000;
														assign node2397 = (inp[2]) ? 8'b10100000 : 8'b10111000;
										assign node2400 = (inp[3]) ? node2424 : node2401;
											assign node2401 = (inp[1]) ? node2411 : node2402;
												assign node2402 = (inp[2]) ? node2408 : node2403;
													assign node2403 = (inp[6]) ? 8'b10101100 : node2404;
														assign node2404 = (inp[12]) ? 8'b10101100 : 8'b10111001;
													assign node2408 = (inp[12]) ? 8'b10111001 : 8'b10101001;
												assign node2411 = (inp[12]) ? node2417 : node2412;
													assign node2412 = (inp[6]) ? 8'b10111000 : node2413;
														assign node2413 = (inp[2]) ? 8'b10101000 : 8'b10111000;
													assign node2417 = (inp[6]) ? node2421 : node2418;
														assign node2418 = (inp[2]) ? 8'b10111000 : 8'b10101001;
														assign node2421 = (inp[2]) ? 8'b10101001 : 8'b10111001;
											assign node2424 = (inp[1]) ? node2434 : node2425;
												assign node2425 = (inp[2]) ? node2429 : node2426;
													assign node2426 = (inp[12]) ? 8'b10101101 : 8'b10111100;
													assign node2429 = (inp[12]) ? 8'b10111100 : node2430;
														assign node2430 = (inp[6]) ? 8'b10111100 : 8'b10101100;
												assign node2434 = (inp[6]) ? 8'b10101100 : node2435;
													assign node2435 = (inp[2]) ? node2439 : node2436;
														assign node2436 = (inp[12]) ? 8'b10101100 : 8'b10111001;
														assign node2439 = (inp[12]) ? 8'b10111001 : 8'b10101001;
								assign node2443 = (inp[10]) ? node2519 : node2444;
									assign node2444 = (inp[1]) ? node2484 : node2445;
										assign node2445 = (inp[4]) ? node2457 : node2446;
											assign node2446 = (inp[2]) ? node2450 : node2447;
												assign node2447 = (inp[12]) ? 8'b10011101 : 8'b10001101;
												assign node2450 = (inp[12]) ? node2454 : node2451;
													assign node2451 = (inp[6]) ? 8'b10011100 : 8'b10001100;
													assign node2454 = (inp[6]) ? 8'b10001101 : 8'b10011100;
											assign node2457 = (inp[3]) ? node2473 : node2458;
												assign node2458 = (inp[6]) ? node2466 : node2459;
													assign node2459 = (inp[2]) ? node2463 : node2460;
														assign node2460 = (inp[12]) ? 8'b10000100 : 8'b10010001;
														assign node2463 = (inp[12]) ? 8'b10010001 : 8'b10000001;
													assign node2466 = (inp[2]) ? node2470 : node2467;
														assign node2467 = (inp[12]) ? 8'b10011100 : 8'b10001100;
														assign node2470 = (inp[12]) ? 8'b10000100 : 8'b10010001;
												assign node2473 = (inp[12]) ? node2479 : node2474;
													assign node2474 = (inp[6]) ? 8'b10011100 : node2475;
														assign node2475 = (inp[2]) ? 8'b10001100 : 8'b10011100;
													assign node2479 = (inp[2]) ? node2481 : 8'b10001101;
														assign node2481 = (inp[6]) ? 8'b10001101 : 8'b10011100;
										assign node2484 = (inp[2]) ? node2504 : node2485;
											assign node2485 = (inp[3]) ? node2493 : node2486;
												assign node2486 = (inp[12]) ? node2488 : 8'b10001001;
													assign node2488 = (inp[4]) ? node2490 : 8'b10011001;
														assign node2490 = (inp[6]) ? 8'b10011001 : 8'b10000001;
												assign node2493 = (inp[12]) ? node2499 : node2494;
													assign node2494 = (inp[6]) ? 8'b10001100 : node2495;
														assign node2495 = (inp[4]) ? 8'b10010001 : 8'b10001100;
													assign node2499 = (inp[4]) ? node2501 : 8'b10011100;
														assign node2501 = (inp[6]) ? 8'b10011100 : 8'b10000100;
											assign node2504 = (inp[3]) ? node2512 : node2505;
												assign node2505 = (inp[6]) ? node2509 : node2506;
													assign node2506 = (inp[12]) ? 8'b10010000 : 8'b10000000;
													assign node2509 = (inp[12]) ? 8'b10000001 : 8'b10010000;
												assign node2512 = (inp[12]) ? node2516 : node2513;
													assign node2513 = (inp[6]) ? 8'b10010001 : 8'b10000001;
													assign node2516 = (inp[6]) ? 8'b10000100 : 8'b10010001;
									assign node2519 = (inp[1]) ? node2557 : node2520;
										assign node2520 = (inp[4]) ? node2532 : node2521;
											assign node2521 = (inp[2]) ? node2525 : node2522;
												assign node2522 = (inp[12]) ? 8'b10111001 : 8'b10101001;
												assign node2525 = (inp[12]) ? node2529 : node2526;
													assign node2526 = (inp[6]) ? 8'b10111000 : 8'b10101000;
													assign node2529 = (inp[6]) ? 8'b10101001 : 8'b10111000;
											assign node2532 = (inp[3]) ? node2544 : node2533;
												assign node2533 = (inp[6]) ? node2541 : node2534;
													assign node2534 = (inp[12]) ? node2538 : node2535;
														assign node2535 = (inp[2]) ? 8'b10000101 : 8'b10010101;
														assign node2538 = (inp[2]) ? 8'b10010101 : 8'b10100000;
													assign node2541 = (inp[2]) ? 8'b10100000 : 8'b10101000;
												assign node2544 = (inp[2]) ? node2550 : node2545;
													assign node2545 = (inp[6]) ? node2547 : 8'b10101001;
														assign node2547 = (inp[12]) ? 8'b10111001 : 8'b10101001;
													assign node2550 = (inp[6]) ? node2554 : node2551;
														assign node2551 = (inp[12]) ? 8'b10111000 : 8'b10101000;
														assign node2554 = (inp[12]) ? 8'b10101001 : 8'b10111000;
										assign node2557 = (inp[2]) ? node2575 : node2558;
											assign node2558 = (inp[3]) ? node2566 : node2559;
												assign node2559 = (inp[12]) ? node2561 : 8'b10001101;
													assign node2561 = (inp[6]) ? 8'b10011101 : node2562;
														assign node2562 = (inp[4]) ? 8'b10000101 : 8'b10011101;
												assign node2566 = (inp[6]) ? node2572 : node2567;
													assign node2567 = (inp[4]) ? node2569 : 8'b10101000;
														assign node2569 = (inp[12]) ? 8'b10100000 : 8'b10010101;
													assign node2572 = (inp[12]) ? 8'b10111000 : 8'b10101000;
											assign node2575 = (inp[3]) ? node2583 : node2576;
												assign node2576 = (inp[6]) ? node2580 : node2577;
													assign node2577 = (inp[12]) ? 8'b10010100 : 8'b10000100;
													assign node2580 = (inp[12]) ? 8'b10000101 : 8'b10010100;
												assign node2583 = (inp[12]) ? node2587 : node2584;
													assign node2584 = (inp[6]) ? 8'b10010101 : 8'b10000101;
													assign node2587 = (inp[6]) ? 8'b10100000 : 8'b10010101;
						assign node2590 = (inp[8]) ? node2816 : node2591;
							assign node2591 = (inp[4]) ? node2645 : node2592;
								assign node2592 = (inp[1]) ? node2610 : node2593;
									assign node2593 = (inp[11]) ? node2599 : node2594;
										assign node2594 = (inp[6]) ? node2596 : 8'b00011111;
											assign node2596 = (inp[2]) ? 8'b00001111 : 8'b00011111;
										assign node2599 = (inp[2]) ? node2603 : node2600;
											assign node2600 = (inp[12]) ? 8'b00011111 : 8'b00001111;
											assign node2603 = (inp[6]) ? node2607 : node2604;
												assign node2604 = (inp[12]) ? 8'b00011110 : 8'b00001110;
												assign node2607 = (inp[12]) ? 8'b00001111 : 8'b00011110;
									assign node2610 = (inp[11]) ? node2622 : node2611;
										assign node2611 = (inp[3]) ? node2617 : node2612;
											assign node2612 = (inp[6]) ? node2614 : 8'b00011111;
												assign node2614 = (inp[2]) ? 8'b00001111 : 8'b00011111;
											assign node2617 = (inp[2]) ? node2619 : 8'b00011110;
												assign node2619 = (inp[6]) ? 8'b00001110 : 8'b00011110;
										assign node2622 = (inp[3]) ? node2634 : node2623;
											assign node2623 = (inp[2]) ? node2627 : node2624;
												assign node2624 = (inp[12]) ? 8'b00011011 : 8'b00001011;
												assign node2627 = (inp[12]) ? node2631 : node2628;
													assign node2628 = (inp[6]) ? 8'b00011010 : 8'b00001010;
													assign node2631 = (inp[6]) ? 8'b00001011 : 8'b00011010;
											assign node2634 = (inp[2]) ? node2638 : node2635;
												assign node2635 = (inp[12]) ? 8'b00011110 : 8'b00001110;
												assign node2638 = (inp[6]) ? node2642 : node2639;
													assign node2639 = (inp[12]) ? 8'b00011011 : 8'b00001011;
													assign node2642 = (inp[12]) ? 8'b00001110 : 8'b00011011;
								assign node2645 = (inp[10]) ? node2729 : node2646;
									assign node2646 = (inp[3]) ? node2680 : node2647;
										assign node2647 = (inp[11]) ? node2665 : node2648;
											assign node2648 = (inp[1]) ? node2658 : node2649;
												assign node2649 = (inp[2]) ? node2653 : node2650;
													assign node2650 = (inp[12]) ? 8'b00000010 : 8'b00011010;
													assign node2653 = (inp[6]) ? node2655 : 8'b10010000;
														assign node2655 = (inp[12]) ? 8'b00000010 : 8'b10000010;
												assign node2658 = (inp[2]) ? node2662 : node2659;
													assign node2659 = (inp[6]) ? 8'b10011001 : 8'b10000001;
													assign node2662 = (inp[6]) ? 8'b10000001 : 8'b10010001;
											assign node2665 = (inp[1]) ? node2673 : node2666;
												assign node2666 = (inp[12]) ? 8'b11110101 : node2667;
													assign node2667 = (inp[2]) ? node2669 : 8'b11110111;
														assign node2669 = (inp[6]) ? 8'b11110111 : 8'b10100101;
												assign node2673 = (inp[2]) ? node2677 : node2674;
													assign node2674 = (inp[12]) ? 8'b10100101 : 8'b10101101;
													assign node2677 = (inp[12]) ? 8'b10110100 : 8'b10100100;
										assign node2680 = (inp[1]) ? node2708 : node2681;
											assign node2681 = (inp[11]) ? node2693 : node2682;
												assign node2682 = (inp[12]) ? node2688 : node2683;
													assign node2683 = (inp[6]) ? 8'b00001011 : node2684;
														assign node2684 = (inp[2]) ? 8'b00011011 : 8'b00001011;
													assign node2688 = (inp[2]) ? node2690 : 8'b00011011;
														assign node2690 = (inp[6]) ? 8'b00001011 : 8'b00011011;
												assign node2693 = (inp[12]) ? node2701 : node2694;
													assign node2694 = (inp[6]) ? node2698 : node2695;
														assign node2695 = (inp[2]) ? 8'b00001010 : 8'b00011010;
														assign node2698 = (inp[2]) ? 8'b00011010 : 8'b00001011;
													assign node2701 = (inp[2]) ? node2705 : node2702;
														assign node2702 = (inp[6]) ? 8'b00011011 : 8'b00001011;
														assign node2705 = (inp[6]) ? 8'b00001011 : 8'b00011010;
											assign node2708 = (inp[6]) ? node2720 : node2709;
												assign node2709 = (inp[11]) ? node2713 : node2710;
													assign node2710 = (inp[2]) ? 8'b10010000 : 8'b10000010;
													assign node2713 = (inp[2]) ? node2717 : node2714;
														assign node2714 = (inp[12]) ? 8'b00000010 : 8'b11110111;
														assign node2717 = (inp[12]) ? 8'b11110101 : 8'b10100101;
												assign node2720 = (inp[2]) ? node2724 : node2721;
													assign node2721 = (inp[12]) ? 8'b00011010 : 8'b00001010;
													assign node2724 = (inp[12]) ? 8'b00000010 : node2725;
														assign node2725 = (inp[11]) ? 8'b11110111 : 8'b10000010;
									assign node2729 = (inp[11]) ? node2765 : node2730;
										assign node2730 = (inp[2]) ? node2746 : node2731;
											assign node2731 = (inp[6]) ? node2739 : node2732;
												assign node2732 = (inp[1]) ? node2736 : node2733;
													assign node2733 = (inp[3]) ? 8'b00001111 : 8'b00001110;
													assign node2736 = (inp[3]) ? 8'b00001110 : 8'b00001111;
												assign node2739 = (inp[1]) ? node2743 : node2740;
													assign node2740 = (inp[3]) ? 8'b00011111 : 8'b00011110;
													assign node2743 = (inp[3]) ? 8'b00011110 : 8'b00011111;
											assign node2746 = (inp[6]) ? node2758 : node2747;
												assign node2747 = (inp[12]) ? node2753 : node2748;
													assign node2748 = (inp[1]) ? 8'b00011111 : node2749;
														assign node2749 = (inp[3]) ? 8'b00011111 : 8'b00011110;
													assign node2753 = (inp[3]) ? node2755 : 8'b00011111;
														assign node2755 = (inp[1]) ? 8'b00011110 : 8'b00011111;
												assign node2758 = (inp[3]) ? node2762 : node2759;
													assign node2759 = (inp[1]) ? 8'b00001111 : 8'b00001110;
													assign node2762 = (inp[1]) ? 8'b00001110 : 8'b00001111;
										assign node2765 = (inp[1]) ? node2793 : node2766;
											assign node2766 = (inp[3]) ? node2780 : node2767;
												assign node2767 = (inp[12]) ? node2773 : node2768;
													assign node2768 = (inp[2]) ? node2770 : 8'b00011011;
														assign node2770 = (inp[6]) ? 8'b00011011 : 8'b00001011;
													assign node2773 = (inp[2]) ? node2777 : node2774;
														assign node2774 = (inp[6]) ? 8'b00011110 : 8'b00001110;
														assign node2777 = (inp[6]) ? 8'b00001110 : 8'b00011011;
												assign node2780 = (inp[6]) ? node2788 : node2781;
													assign node2781 = (inp[12]) ? node2785 : node2782;
														assign node2782 = (inp[2]) ? 8'b00001110 : 8'b00011110;
														assign node2785 = (inp[2]) ? 8'b00011110 : 8'b00001111;
													assign node2788 = (inp[12]) ? node2790 : 8'b00001111;
														assign node2790 = (inp[2]) ? 8'b00001111 : 8'b00011111;
											assign node2793 = (inp[6]) ? node2809 : node2794;
												assign node2794 = (inp[3]) ? node2802 : node2795;
													assign node2795 = (inp[2]) ? node2799 : node2796;
														assign node2796 = (inp[12]) ? 8'b00001011 : 8'b00011010;
														assign node2799 = (inp[12]) ? 8'b00011010 : 8'b00001010;
													assign node2802 = (inp[12]) ? node2806 : node2803;
														assign node2803 = (inp[2]) ? 8'b00001011 : 8'b00011011;
														assign node2806 = (inp[2]) ? 8'b00011011 : 8'b00001110;
												assign node2809 = (inp[3]) ? 8'b00011011 : node2810;
													assign node2810 = (inp[2]) ? 8'b00001011 : node2811;
														assign node2811 = (inp[12]) ? 8'b00011011 : 8'b00001011;
							assign node2816 = (inp[10]) ? node2916 : node2817;
								assign node2817 = (inp[11]) ? node2861 : node2818;
									assign node2818 = (inp[4]) ? node2832 : node2819;
										assign node2819 = (inp[1]) ? node2825 : node2820;
											assign node2820 = (inp[6]) ? node2822 : 8'b10011101;
												assign node2822 = (inp[2]) ? 8'b10001101 : 8'b10011101;
											assign node2825 = (inp[3]) ? node2829 : node2826;
												assign node2826 = (inp[2]) ? 8'b10010101 : 8'b10011101;
												assign node2829 = (inp[2]) ? 8'b10010100 : 8'b10011100;
										assign node2832 = (inp[6]) ? node2846 : node2833;
											assign node2833 = (inp[2]) ? node2841 : node2834;
												assign node2834 = (inp[1]) ? node2838 : node2835;
													assign node2835 = (inp[3]) ? 8'b10001101 : 8'b10000100;
													assign node2838 = (inp[3]) ? 8'b10000100 : 8'b10000101;
												assign node2841 = (inp[1]) ? node2843 : 8'b10010100;
													assign node2843 = (inp[3]) ? 8'b10010100 : 8'b10010101;
											assign node2846 = (inp[2]) ? node2854 : node2847;
												assign node2847 = (inp[1]) ? node2851 : node2848;
													assign node2848 = (inp[3]) ? 8'b10011101 : 8'b10011100;
													assign node2851 = (inp[3]) ? 8'b10011100 : 8'b10011101;
												assign node2854 = (inp[3]) ? node2858 : node2855;
													assign node2855 = (inp[1]) ? 8'b10000101 : 8'b10000100;
													assign node2858 = (inp[1]) ? 8'b10000100 : 8'b10001101;
									assign node2861 = (inp[1]) ? node2891 : node2862;
										assign node2862 = (inp[4]) ? node2874 : node2863;
											assign node2863 = (inp[2]) ? node2867 : node2864;
												assign node2864 = (inp[12]) ? 8'b11111101 : 8'b10101101;
												assign node2867 = (inp[12]) ? node2871 : node2868;
													assign node2868 = (inp[6]) ? 8'b10111100 : 8'b10101100;
													assign node2871 = (inp[6]) ? 8'b10101101 : 8'b10111100;
											assign node2874 = (inp[3]) ? node2884 : node2875;
												assign node2875 = (inp[2]) ? node2879 : node2876;
													assign node2876 = (inp[12]) ? 8'b10100100 : 8'b10101100;
													assign node2879 = (inp[6]) ? node2881 : 8'b10110001;
														assign node2881 = (inp[12]) ? 8'b10100100 : 8'b10110001;
												assign node2884 = (inp[6]) ? node2886 : 8'b10111100;
													assign node2886 = (inp[2]) ? node2888 : 8'b11111101;
														assign node2888 = (inp[12]) ? 8'b10101101 : 8'b10111100;
										assign node2891 = (inp[3]) ? node2905 : node2892;
											assign node2892 = (inp[6]) ? node2898 : node2893;
												assign node2893 = (inp[12]) ? 8'b10110000 : node2894;
													assign node2894 = (inp[2]) ? 8'b10100000 : 8'b10110000;
												assign node2898 = (inp[2]) ? node2902 : node2899;
													assign node2899 = (inp[12]) ? 8'b10111001 : 8'b10101001;
													assign node2902 = (inp[12]) ? 8'b10100001 : 8'b10110000;
											assign node2905 = (inp[12]) ? node2907 : 8'b10110001;
												assign node2907 = (inp[2]) ? node2913 : node2908;
													assign node2908 = (inp[4]) ? node2910 : 8'b10111100;
														assign node2910 = (inp[6]) ? 8'b10111100 : 8'b10100100;
													assign node2913 = (inp[6]) ? 8'b10100100 : 8'b10110001;
								assign node2916 = (inp[1]) ? node2978 : node2917;
									assign node2917 = (inp[4]) ? node2935 : node2918;
										assign node2918 = (inp[2]) ? node2924 : node2919;
											assign node2919 = (inp[12]) ? 8'b00011011 : node2920;
												assign node2920 = (inp[11]) ? 8'b00001011 : 8'b00011011;
											assign node2924 = (inp[11]) ? node2928 : node2925;
												assign node2925 = (inp[6]) ? 8'b00001011 : 8'b00011011;
												assign node2928 = (inp[12]) ? node2932 : node2929;
													assign node2929 = (inp[6]) ? 8'b00011010 : 8'b00001010;
													assign node2932 = (inp[6]) ? 8'b00001011 : 8'b00011010;
										assign node2935 = (inp[3]) ? node2957 : node2936;
											assign node2936 = (inp[12]) ? node2950 : node2937;
												assign node2937 = (inp[11]) ? node2945 : node2938;
													assign node2938 = (inp[6]) ? node2942 : node2939;
														assign node2939 = (inp[2]) ? 8'b10010000 : 8'b10000010;
														assign node2942 = (inp[2]) ? 8'b10000010 : 8'b00011010;
													assign node2945 = (inp[6]) ? 8'b11110111 : node2946;
														assign node2946 = (inp[2]) ? 8'b10100101 : 8'b11110111;
												assign node2950 = (inp[2]) ? node2954 : node2951;
													assign node2951 = (inp[6]) ? 8'b00011010 : 8'b00000010;
													assign node2954 = (inp[11]) ? 8'b00000010 : 8'b10010000;
											assign node2957 = (inp[11]) ? node2969 : node2958;
												assign node2958 = (inp[12]) ? node2964 : node2959;
													assign node2959 = (inp[2]) ? node2961 : 8'b00001011;
														assign node2961 = (inp[6]) ? 8'b00001011 : 8'b00011011;
													assign node2964 = (inp[2]) ? node2966 : 8'b00011011;
														assign node2966 = (inp[6]) ? 8'b00001011 : 8'b00011011;
												assign node2969 = (inp[12]) ? node2975 : node2970;
													assign node2970 = (inp[2]) ? node2972 : 8'b00011010;
														assign node2972 = (inp[6]) ? 8'b00011010 : 8'b00001010;
													assign node2975 = (inp[2]) ? 8'b00011010 : 8'b00001011;
									assign node2978 = (inp[11]) ? node3002 : node2979;
										assign node2979 = (inp[3]) ? node2989 : node2980;
											assign node2980 = (inp[2]) ? node2986 : node2981;
												assign node2981 = (inp[6]) ? 8'b10011001 : node2982;
													assign node2982 = (inp[4]) ? 8'b10000001 : 8'b10011001;
												assign node2986 = (inp[6]) ? 8'b10000001 : 8'b10010001;
											assign node2989 = (inp[2]) ? node2997 : node2990;
												assign node2990 = (inp[6]) ? 8'b00011010 : node2991;
													assign node2991 = (inp[4]) ? node2993 : 8'b00011010;
														assign node2993 = (inp[12]) ? 8'b00000010 : 8'b10000010;
												assign node2997 = (inp[6]) ? node2999 : 8'b10010000;
													assign node2999 = (inp[12]) ? 8'b00000010 : 8'b10000010;
										assign node3002 = (inp[3]) ? node3018 : node3003;
											assign node3003 = (inp[2]) ? node3011 : node3004;
												assign node3004 = (inp[6]) ? node3008 : node3005;
													assign node3005 = (inp[4]) ? 8'b10100101 : 8'b10101101;
													assign node3008 = (inp[12]) ? 8'b11111101 : 8'b10101101;
												assign node3011 = (inp[12]) ? node3015 : node3012;
													assign node3012 = (inp[6]) ? 8'b10110100 : 8'b10100100;
													assign node3015 = (inp[6]) ? 8'b10100101 : 8'b10110100;
											assign node3018 = (inp[6]) ? node3024 : node3019;
												assign node3019 = (inp[2]) ? node3021 : 8'b11110111;
													assign node3021 = (inp[12]) ? 8'b11110101 : 8'b10100101;
												assign node3024 = (inp[2]) ? node3028 : node3025;
													assign node3025 = (inp[12]) ? 8'b00011010 : 8'b00001010;
													assign node3028 = (inp[12]) ? 8'b00000010 : 8'b11110111;
				assign node3031 = (inp[11]) ? node3319 : node3032;
					assign node3032 = (inp[0]) ? node3248 : node3033;
						assign node3033 = (inp[9]) ? node3149 : node3034;
							assign node3034 = (inp[8]) ? node3078 : node3035;
								assign node3035 = (inp[3]) ? node3059 : node3036;
									assign node3036 = (inp[4]) ? node3048 : node3037;
										assign node3037 = (inp[1]) ? node3043 : node3038;
											assign node3038 = (inp[2]) ? node3040 : 8'b00011111;
												assign node3040 = (inp[6]) ? 8'b00011111 : 8'b00001111;
											assign node3043 = (inp[6]) ? 8'b00011110 : node3044;
												assign node3044 = (inp[2]) ? 8'b00001110 : 8'b00011110;
										assign node3048 = (inp[10]) ? node3056 : node3049;
											assign node3049 = (inp[6]) ? node3053 : node3050;
												assign node3050 = (inp[12]) ? 8'b00000010 : 8'b10000010;
												assign node3053 = (inp[2]) ? 8'b10010000 : 8'b00011010;
											assign node3056 = (inp[6]) ? 8'b00011110 : 8'b00001110;
									assign node3059 = (inp[6]) ? node3069 : node3060;
										assign node3060 = (inp[4]) ? node3064 : node3061;
											assign node3061 = (inp[2]) ? 8'b00001111 : 8'b00011111;
											assign node3064 = (inp[10]) ? 8'b00001111 : node3065;
												assign node3065 = (inp[1]) ? 8'b10000001 : 8'b00001011;
										assign node3069 = (inp[10]) ? 8'b00011111 : node3070;
											assign node3070 = (inp[4]) ? node3072 : 8'b00011111;
												assign node3072 = (inp[1]) ? node3074 : 8'b00011011;
													assign node3074 = (inp[12]) ? 8'b10011001 : 8'b10010001;
								assign node3078 = (inp[10]) ? node3118 : node3079;
									assign node3079 = (inp[1]) ? node3097 : node3080;
										assign node3080 = (inp[4]) ? node3086 : node3081;
											assign node3081 = (inp[2]) ? node3083 : 8'b00011011;
												assign node3083 = (inp[6]) ? 8'b00011011 : 8'b00001011;
											assign node3086 = (inp[3]) ? node3094 : node3087;
												assign node3087 = (inp[2]) ? 8'b10010000 : node3088;
													assign node3088 = (inp[6]) ? 8'b00011010 : node3089;
														assign node3089 = (inp[12]) ? 8'b00000010 : 8'b10000010;
												assign node3094 = (inp[6]) ? 8'b00011011 : 8'b00001011;
										assign node3097 = (inp[3]) ? node3109 : node3098;
											assign node3098 = (inp[2]) ? node3106 : node3099;
												assign node3099 = (inp[6]) ? 8'b00011010 : node3100;
													assign node3100 = (inp[4]) ? node3102 : 8'b00011010;
														assign node3102 = (inp[12]) ? 8'b00000010 : 8'b10000010;
												assign node3106 = (inp[6]) ? 8'b10010000 : 8'b00000010;
											assign node3109 = (inp[2]) ? node3115 : node3110;
												assign node3110 = (inp[6]) ? 8'b10011001 : node3111;
													assign node3111 = (inp[4]) ? 8'b10000001 : 8'b10011001;
												assign node3115 = (inp[6]) ? 8'b10010001 : 8'b10000001;
									assign node3118 = (inp[6]) ? node3130 : node3119;
										assign node3119 = (inp[1]) ? node3127 : node3120;
											assign node3120 = (inp[4]) ? node3124 : node3121;
												assign node3121 = (inp[2]) ? 8'b10001101 : 8'b10011101;
												assign node3124 = (inp[3]) ? 8'b10001101 : 8'b10000100;
											assign node3127 = (inp[3]) ? 8'b10000101 : 8'b10000100;
										assign node3130 = (inp[3]) ? node3144 : node3131;
											assign node3131 = (inp[2]) ? node3139 : node3132;
												assign node3132 = (inp[12]) ? 8'b10011100 : node3133;
													assign node3133 = (inp[4]) ? 8'b10011100 : node3134;
														assign node3134 = (inp[1]) ? 8'b10011100 : 8'b10011101;
												assign node3139 = (inp[1]) ? 8'b10010100 : node3140;
													assign node3140 = (inp[4]) ? 8'b10010100 : 8'b10011101;
											assign node3144 = (inp[2]) ? node3146 : 8'b10011101;
												assign node3146 = (inp[1]) ? 8'b10010101 : 8'b10011101;
							assign node3149 = (inp[6]) ? node3203 : node3150;
								assign node3150 = (inp[3]) ? node3176 : node3151;
									assign node3151 = (inp[4]) ? node3171 : node3152;
										assign node3152 = (inp[2]) ? node3162 : node3153;
											assign node3153 = (inp[1]) ? node3157 : node3154;
												assign node3154 = (inp[8]) ? 8'b10111001 : 8'b11111101;
												assign node3157 = (inp[10]) ? 8'b10111100 : node3158;
													assign node3158 = (inp[8]) ? 8'b10111000 : 8'b10111100;
											assign node3162 = (inp[1]) ? node3168 : node3163;
												assign node3163 = (inp[10]) ? 8'b10101101 : node3164;
													assign node3164 = (inp[8]) ? 8'b10101001 : 8'b10101101;
												assign node3168 = (inp[8]) ? 8'b10100000 : 8'b10101100;
										assign node3171 = (inp[10]) ? node3173 : 8'b10100000;
											assign node3173 = (inp[8]) ? 8'b10100100 : 8'b10101100;
									assign node3176 = (inp[10]) ? node3190 : node3177;
										assign node3177 = (inp[4]) ? node3187 : node3178;
											assign node3178 = (inp[8]) ? node3182 : node3179;
												assign node3179 = (inp[2]) ? 8'b10101101 : 8'b11111101;
												assign node3182 = (inp[2]) ? node3184 : 8'b10111001;
													assign node3184 = (inp[1]) ? 8'b10100001 : 8'b10101001;
											assign node3187 = (inp[1]) ? 8'b10100001 : 8'b10101001;
										assign node3190 = (inp[4]) ? node3198 : node3191;
											assign node3191 = (inp[2]) ? node3193 : 8'b11111101;
												assign node3193 = (inp[1]) ? node3195 : 8'b10101101;
													assign node3195 = (inp[8]) ? 8'b10100101 : 8'b10101101;
											assign node3198 = (inp[1]) ? node3200 : 8'b10101101;
												assign node3200 = (inp[8]) ? 8'b10100101 : 8'b10101101;
								assign node3203 = (inp[10]) ? node3231 : node3204;
									assign node3204 = (inp[3]) ? node3218 : node3205;
										assign node3205 = (inp[4]) ? node3215 : node3206;
											assign node3206 = (inp[8]) ? node3210 : node3207;
												assign node3207 = (inp[1]) ? 8'b10111100 : 8'b11111101;
												assign node3210 = (inp[1]) ? node3212 : 8'b10111001;
													assign node3212 = (inp[2]) ? 8'b10110000 : 8'b10111000;
											assign node3215 = (inp[2]) ? 8'b10110000 : 8'b10111000;
										assign node3218 = (inp[8]) ? node3226 : node3219;
											assign node3219 = (inp[4]) ? node3221 : 8'b11111101;
												assign node3221 = (inp[1]) ? node3223 : 8'b10111001;
													assign node3223 = (inp[2]) ? 8'b10110001 : 8'b10111001;
											assign node3226 = (inp[2]) ? node3228 : 8'b10111001;
												assign node3228 = (inp[1]) ? 8'b10110001 : 8'b10111001;
									assign node3231 = (inp[3]) ? node3241 : node3232;
										assign node3232 = (inp[4]) ? node3236 : node3233;
											assign node3233 = (inp[1]) ? 8'b10111100 : 8'b11111101;
											assign node3236 = (inp[2]) ? node3238 : 8'b10111100;
												assign node3238 = (inp[8]) ? 8'b10110100 : 8'b10111100;
										assign node3241 = (inp[1]) ? node3243 : 8'b11111101;
											assign node3243 = (inp[2]) ? node3245 : 8'b11111101;
												assign node3245 = (inp[8]) ? 8'b11110101 : 8'b11111101;
						assign node3248 = (inp[4]) ? node3256 : node3249;
							assign node3249 = (inp[8]) ? node3251 : 8'b11111101;
								assign node3251 = (inp[1]) ? node3253 : 8'b11111101;
									assign node3253 = (inp[2]) ? 8'b11110101 : 8'b11111101;
							assign node3256 = (inp[8]) ? node3292 : node3257;
								assign node3257 = (inp[10]) ? node3275 : node3258;
									assign node3258 = (inp[2]) ? node3268 : node3259;
										assign node3259 = (inp[6]) ? node3265 : node3260;
											assign node3260 = (inp[1]) ? 8'b10100001 : node3261;
												assign node3261 = (inp[3]) ? 8'b10101001 : 8'b10100000;
											assign node3265 = (inp[1]) ? 8'b10111001 : 8'b10111000;
										assign node3268 = (inp[3]) ? node3272 : node3269;
											assign node3269 = (inp[1]) ? 8'b10110001 : 8'b10110000;
											assign node3272 = (inp[1]) ? 8'b10110001 : 8'b10111001;
									assign node3275 = (inp[3]) ? node3287 : node3276;
										assign node3276 = (inp[1]) ? node3282 : node3277;
											assign node3277 = (inp[2]) ? 8'b10111100 : node3278;
												assign node3278 = (inp[6]) ? 8'b10111100 : 8'b10101100;
											assign node3282 = (inp[2]) ? 8'b11111101 : node3283;
												assign node3283 = (inp[6]) ? 8'b11111101 : 8'b10101101;
										assign node3287 = (inp[6]) ? 8'b11111101 : node3288;
											assign node3288 = (inp[2]) ? 8'b11111101 : 8'b10101101;
								assign node3292 = (inp[6]) ? node3306 : node3293;
									assign node3293 = (inp[2]) ? node3301 : node3294;
										assign node3294 = (inp[3]) ? node3298 : node3295;
											assign node3295 = (inp[1]) ? 8'b10100101 : 8'b10100100;
											assign node3298 = (inp[1]) ? 8'b10100101 : 8'b10101101;
										assign node3301 = (inp[1]) ? 8'b11110101 : node3302;
											assign node3302 = (inp[3]) ? 8'b11111101 : 8'b10110100;
									assign node3306 = (inp[2]) ? node3312 : node3307;
										assign node3307 = (inp[3]) ? 8'b11111101 : node3308;
											assign node3308 = (inp[1]) ? 8'b11111101 : 8'b10111100;
										assign node3312 = (inp[3]) ? node3316 : node3313;
											assign node3313 = (inp[1]) ? 8'b11110101 : 8'b10110100;
											assign node3316 = (inp[1]) ? 8'b11110101 : 8'b11111101;
					assign node3319 = (inp[8]) ? node3739 : node3320;
						assign node3320 = (inp[9]) ? node3540 : node3321;
							assign node3321 = (inp[0]) ? node3467 : node3322;
								assign node3322 = (inp[10]) ? node3400 : node3323;
									assign node3323 = (inp[4]) ? node3353 : node3324;
										assign node3324 = (inp[1]) ? node3336 : node3325;
											assign node3325 = (inp[2]) ? node3329 : node3326;
												assign node3326 = (inp[12]) ? 8'b00011111 : 8'b00001111;
												assign node3329 = (inp[12]) ? node3333 : node3330;
													assign node3330 = (inp[6]) ? 8'b00001110 : 8'b00011110;
													assign node3333 = (inp[6]) ? 8'b00011110 : 8'b00001111;
											assign node3336 = (inp[3]) ? node3346 : node3337;
												assign node3337 = (inp[2]) ? node3341 : node3338;
													assign node3338 = (inp[12]) ? 8'b00011110 : 8'b00001110;
													assign node3341 = (inp[6]) ? 8'b00011011 : node3342;
														assign node3342 = (inp[12]) ? 8'b00001110 : 8'b00011011;
												assign node3346 = (inp[2]) ? node3350 : node3347;
													assign node3347 = (inp[12]) ? 8'b00011011 : 8'b00001011;
													assign node3350 = (inp[12]) ? 8'b00011010 : 8'b00001010;
										assign node3353 = (inp[1]) ? node3381 : node3354;
											assign node3354 = (inp[3]) ? node3366 : node3355;
												assign node3355 = (inp[2]) ? node3361 : node3356;
													assign node3356 = (inp[6]) ? node3358 : 8'b00000010;
														assign node3358 = (inp[12]) ? 8'b00011010 : 8'b00001010;
													assign node3361 = (inp[6]) ? node3363 : 8'b11110111;
														assign node3363 = (inp[12]) ? 8'b11110101 : 8'b10100101;
												assign node3366 = (inp[2]) ? node3374 : node3367;
													assign node3367 = (inp[12]) ? node3371 : node3368;
														assign node3368 = (inp[6]) ? 8'b00001011 : 8'b00011010;
														assign node3371 = (inp[6]) ? 8'b00011011 : 8'b00001011;
													assign node3374 = (inp[6]) ? node3378 : node3375;
														assign node3375 = (inp[12]) ? 8'b00001011 : 8'b00011010;
														assign node3378 = (inp[12]) ? 8'b00011010 : 8'b00001010;
											assign node3381 = (inp[3]) ? node3391 : node3382;
												assign node3382 = (inp[6]) ? node3386 : node3383;
													assign node3383 = (inp[12]) ? 8'b00000010 : 8'b11110111;
													assign node3386 = (inp[2]) ? node3388 : 8'b00001010;
														assign node3388 = (inp[12]) ? 8'b11110101 : 8'b10100101;
												assign node3391 = (inp[6]) ? node3395 : node3392;
													assign node3392 = (inp[12]) ? 8'b10100101 : 8'b10110100;
													assign node3395 = (inp[2]) ? 8'b10100100 : node3396;
														assign node3396 = (inp[12]) ? 8'b11111101 : 8'b10101101;
									assign node3400 = (inp[1]) ? node3434 : node3401;
										assign node3401 = (inp[3]) ? node3415 : node3402;
											assign node3402 = (inp[12]) ? node3410 : node3403;
												assign node3403 = (inp[4]) ? node3405 : 8'b00011110;
													assign node3405 = (inp[6]) ? node3407 : 8'b00011011;
														assign node3407 = (inp[2]) ? 8'b00001011 : 8'b00001110;
												assign node3410 = (inp[6]) ? 8'b00011110 : node3411;
													assign node3411 = (inp[4]) ? 8'b00001110 : 8'b00001111;
											assign node3415 = (inp[2]) ? node3427 : node3416;
												assign node3416 = (inp[12]) ? node3422 : node3417;
													assign node3417 = (inp[6]) ? 8'b00001111 : node3418;
														assign node3418 = (inp[4]) ? 8'b00011110 : 8'b00001111;
													assign node3422 = (inp[6]) ? 8'b00011111 : node3423;
														assign node3423 = (inp[4]) ? 8'b00001111 : 8'b00011111;
												assign node3427 = (inp[4]) ? node3431 : node3428;
													assign node3428 = (inp[12]) ? 8'b00001111 : 8'b00011110;
													assign node3431 = (inp[12]) ? 8'b00011110 : 8'b00001110;
										assign node3434 = (inp[3]) ? node3450 : node3435;
											assign node3435 = (inp[2]) ? node3443 : node3436;
												assign node3436 = (inp[12]) ? node3438 : 8'b00001110;
													assign node3438 = (inp[6]) ? 8'b00011110 : node3439;
														assign node3439 = (inp[4]) ? 8'b00001110 : 8'b00011110;
												assign node3443 = (inp[6]) ? node3447 : node3444;
													assign node3444 = (inp[12]) ? 8'b00001110 : 8'b00011011;
													assign node3447 = (inp[12]) ? 8'b00011011 : 8'b00001011;
											assign node3450 = (inp[2]) ? node3460 : node3451;
												assign node3451 = (inp[12]) ? node3457 : node3452;
													assign node3452 = (inp[4]) ? node3454 : 8'b00001011;
														assign node3454 = (inp[6]) ? 8'b00001011 : 8'b00011010;
													assign node3457 = (inp[6]) ? 8'b00011011 : 8'b00001011;
												assign node3460 = (inp[6]) ? node3464 : node3461;
													assign node3461 = (inp[12]) ? 8'b00001011 : 8'b00011010;
													assign node3464 = (inp[12]) ? 8'b00011010 : 8'b00001010;
								assign node3467 = (inp[12]) ? node3505 : node3468;
									assign node3468 = (inp[2]) ? node3490 : node3469;
										assign node3469 = (inp[4]) ? node3473 : node3470;
											assign node3470 = (inp[1]) ? 8'b10101001 : 8'b10101101;
											assign node3473 = (inp[6]) ? node3481 : node3474;
												assign node3474 = (inp[1]) ? node3478 : node3475;
													assign node3475 = (inp[10]) ? 8'b10111100 : 8'b10111000;
													assign node3478 = (inp[10]) ? 8'b10111000 : 8'b10010100;
												assign node3481 = (inp[1]) ? node3487 : node3482;
													assign node3482 = (inp[10]) ? 8'b10101100 : node3483;
														assign node3483 = (inp[3]) ? 8'b10101001 : 8'b10101000;
													assign node3487 = (inp[10]) ? 8'b10101001 : 8'b10001101;
										assign node3490 = (inp[10]) ? node3498 : node3491;
											assign node3491 = (inp[4]) ? node3495 : node3492;
												assign node3492 = (inp[1]) ? 8'b10101000 : 8'b10101100;
												assign node3495 = (inp[1]) ? 8'b10000100 : 8'b10101000;
											assign node3498 = (inp[1]) ? 8'b10101000 : node3499;
												assign node3499 = (inp[4]) ? node3501 : 8'b10101100;
													assign node3501 = (inp[3]) ? 8'b10101100 : 8'b10101001;
									assign node3505 = (inp[2]) ? node3525 : node3506;
										assign node3506 = (inp[4]) ? node3510 : node3507;
											assign node3507 = (inp[1]) ? 8'b10111001 : 8'b11111101;
											assign node3510 = (inp[6]) ? node3520 : node3511;
												assign node3511 = (inp[10]) ? node3517 : node3512;
													assign node3512 = (inp[1]) ? 8'b10000101 : node3513;
														assign node3513 = (inp[3]) ? 8'b10101001 : 8'b10100000;
													assign node3517 = (inp[1]) ? 8'b10101001 : 8'b10101100;
												assign node3520 = (inp[10]) ? 8'b10111001 : node3521;
													assign node3521 = (inp[1]) ? 8'b10011101 : 8'b10111001;
										assign node3525 = (inp[1]) ? node3535 : node3526;
											assign node3526 = (inp[4]) ? node3528 : 8'b10111100;
												assign node3528 = (inp[3]) ? node3532 : node3529;
													assign node3529 = (inp[10]) ? 8'b10111001 : 8'b10010101;
													assign node3532 = (inp[10]) ? 8'b10111100 : 8'b10111000;
											assign node3535 = (inp[10]) ? 8'b10111000 : node3536;
												assign node3536 = (inp[4]) ? 8'b10010100 : 8'b10111000;
							assign node3540 = (inp[12]) ? node3650 : node3541;
								assign node3541 = (inp[6]) ? node3597 : node3542;
									assign node3542 = (inp[4]) ? node3560 : node3543;
										assign node3543 = (inp[2]) ? node3551 : node3544;
											assign node3544 = (inp[1]) ? node3546 : 8'b10101101;
												assign node3546 = (inp[3]) ? 8'b10101001 : node3547;
													assign node3547 = (inp[0]) ? 8'b10101001 : 8'b10101100;
											assign node3551 = (inp[1]) ? node3555 : node3552;
												assign node3552 = (inp[0]) ? 8'b10101100 : 8'b10111100;
												assign node3555 = (inp[0]) ? 8'b10101000 : node3556;
													assign node3556 = (inp[3]) ? 8'b10111000 : 8'b10111001;
										assign node3560 = (inp[10]) ? node3578 : node3561;
											assign node3561 = (inp[3]) ? node3571 : node3562;
												assign node3562 = (inp[0]) ? node3564 : 8'b10010101;
													assign node3564 = (inp[1]) ? node3568 : node3565;
														assign node3565 = (inp[2]) ? 8'b10000101 : 8'b10010101;
														assign node3568 = (inp[2]) ? 8'b10000100 : 8'b10010100;
												assign node3571 = (inp[1]) ? 8'b10010100 : node3572;
													assign node3572 = (inp[0]) ? node3574 : 8'b10111000;
														assign node3574 = (inp[2]) ? 8'b10101000 : 8'b10111000;
											assign node3578 = (inp[3]) ? node3586 : node3579;
												assign node3579 = (inp[1]) ? node3581 : 8'b10111001;
													assign node3581 = (inp[0]) ? node3583 : 8'b10111001;
														assign node3583 = (inp[2]) ? 8'b10101000 : 8'b10111000;
												assign node3586 = (inp[1]) ? node3592 : node3587;
													assign node3587 = (inp[0]) ? node3589 : 8'b10111100;
														assign node3589 = (inp[2]) ? 8'b10101100 : 8'b10111100;
													assign node3592 = (inp[2]) ? node3594 : 8'b10111000;
														assign node3594 = (inp[0]) ? 8'b10101000 : 8'b10111000;
									assign node3597 = (inp[2]) ? node3627 : node3598;
										assign node3598 = (inp[3]) ? node3616 : node3599;
											assign node3599 = (inp[4]) ? node3605 : node3600;
												assign node3600 = (inp[1]) ? node3602 : 8'b10101101;
													assign node3602 = (inp[0]) ? 8'b10101001 : 8'b10101100;
												assign node3605 = (inp[0]) ? node3609 : node3606;
													assign node3606 = (inp[10]) ? 8'b10101100 : 8'b10101000;
													assign node3609 = (inp[1]) ? node3613 : node3610;
														assign node3610 = (inp[10]) ? 8'b10101100 : 8'b10101000;
														assign node3613 = (inp[10]) ? 8'b10101001 : 8'b10001101;
											assign node3616 = (inp[1]) ? node3622 : node3617;
												assign node3617 = (inp[4]) ? node3619 : 8'b10101101;
													assign node3619 = (inp[10]) ? 8'b10101101 : 8'b10101001;
												assign node3622 = (inp[4]) ? node3624 : 8'b10101001;
													assign node3624 = (inp[10]) ? 8'b10101001 : 8'b10001101;
										assign node3627 = (inp[1]) ? node3637 : node3628;
											assign node3628 = (inp[4]) ? node3630 : 8'b10101100;
												assign node3630 = (inp[3]) ? node3634 : node3631;
													assign node3631 = (inp[10]) ? 8'b10101001 : 8'b10000101;
													assign node3634 = (inp[10]) ? 8'b10101100 : 8'b10101000;
											assign node3637 = (inp[4]) ? node3643 : node3638;
												assign node3638 = (inp[0]) ? 8'b10101000 : node3639;
													assign node3639 = (inp[3]) ? 8'b10101000 : 8'b10101001;
												assign node3643 = (inp[10]) ? 8'b10101000 : node3644;
													assign node3644 = (inp[3]) ? 8'b10000100 : node3645;
														assign node3645 = (inp[0]) ? 8'b10000100 : 8'b10000101;
								assign node3650 = (inp[1]) ? node3688 : node3651;
									assign node3651 = (inp[4]) ? node3659 : node3652;
										assign node3652 = (inp[2]) ? node3654 : 8'b11111101;
											assign node3654 = (inp[6]) ? 8'b10111100 : node3655;
												assign node3655 = (inp[0]) ? 8'b10111100 : 8'b10101101;
										assign node3659 = (inp[10]) ? node3673 : node3660;
											assign node3660 = (inp[3]) ? node3670 : node3661;
												assign node3661 = (inp[2]) ? node3665 : node3662;
													assign node3662 = (inp[6]) ? 8'b10111000 : 8'b10100000;
													assign node3665 = (inp[0]) ? 8'b10010101 : node3666;
														assign node3666 = (inp[6]) ? 8'b10010101 : 8'b10100000;
												assign node3670 = (inp[2]) ? 8'b10111000 : 8'b10111001;
											assign node3673 = (inp[6]) ? node3681 : node3674;
												assign node3674 = (inp[0]) ? node3676 : 8'b10101100;
													assign node3676 = (inp[2]) ? node3678 : 8'b10101100;
														assign node3678 = (inp[3]) ? 8'b10111100 : 8'b10111001;
												assign node3681 = (inp[2]) ? node3685 : node3682;
													assign node3682 = (inp[3]) ? 8'b11111101 : 8'b10111100;
													assign node3685 = (inp[3]) ? 8'b10111100 : 8'b10111001;
									assign node3688 = (inp[4]) ? node3704 : node3689;
										assign node3689 = (inp[2]) ? node3695 : node3690;
											assign node3690 = (inp[3]) ? 8'b10111001 : node3691;
												assign node3691 = (inp[0]) ? 8'b10111001 : 8'b10111100;
											assign node3695 = (inp[0]) ? 8'b10111000 : node3696;
												assign node3696 = (inp[6]) ? node3700 : node3697;
													assign node3697 = (inp[3]) ? 8'b10101001 : 8'b10101100;
													assign node3700 = (inp[3]) ? 8'b10111000 : 8'b10111001;
										assign node3704 = (inp[10]) ? node3720 : node3705;
											assign node3705 = (inp[3]) ? node3715 : node3706;
												assign node3706 = (inp[2]) ? node3710 : node3707;
													assign node3707 = (inp[6]) ? 8'b10111000 : 8'b10100000;
													assign node3710 = (inp[6]) ? 8'b10010101 : node3711;
														assign node3711 = (inp[0]) ? 8'b10010100 : 8'b10100000;
												assign node3715 = (inp[2]) ? 8'b10010100 : node3716;
													assign node3716 = (inp[6]) ? 8'b10011101 : 8'b10000101;
											assign node3720 = (inp[6]) ? node3730 : node3721;
												assign node3721 = (inp[2]) ? node3727 : node3722;
													assign node3722 = (inp[3]) ? 8'b10101001 : node3723;
														assign node3723 = (inp[0]) ? 8'b10101001 : 8'b10101100;
													assign node3727 = (inp[0]) ? 8'b10111000 : 8'b10101001;
												assign node3730 = (inp[2]) ? node3736 : node3731;
													assign node3731 = (inp[0]) ? 8'b10111001 : node3732;
														assign node3732 = (inp[3]) ? 8'b10111001 : 8'b10111100;
													assign node3736 = (inp[0]) ? 8'b10111000 : 8'b10111001;
						assign node3739 = (inp[2]) ? node3901 : node3740;
							assign node3740 = (inp[0]) ? node3870 : node3741;
								assign node3741 = (inp[10]) ? node3807 : node3742;
									assign node3742 = (inp[9]) ? node3780 : node3743;
										assign node3743 = (inp[3]) ? node3761 : node3744;
											assign node3744 = (inp[6]) ? node3754 : node3745;
												assign node3745 = (inp[4]) ? node3751 : node3746;
													assign node3746 = (inp[1]) ? node3748 : 8'b00001011;
														assign node3748 = (inp[12]) ? 8'b00011010 : 8'b00001010;
													assign node3751 = (inp[12]) ? 8'b00000010 : 8'b11110111;
												assign node3754 = (inp[12]) ? node3756 : 8'b00001010;
													assign node3756 = (inp[1]) ? 8'b00011010 : node3757;
														assign node3757 = (inp[4]) ? 8'b00011010 : 8'b00011011;
											assign node3761 = (inp[1]) ? node3771 : node3762;
												assign node3762 = (inp[4]) ? node3766 : node3763;
													assign node3763 = (inp[12]) ? 8'b00011011 : 8'b00001011;
													assign node3766 = (inp[12]) ? node3768 : 8'b00011010;
														assign node3768 = (inp[6]) ? 8'b00011011 : 8'b00001011;
												assign node3771 = (inp[4]) ? node3775 : node3772;
													assign node3772 = (inp[12]) ? 8'b11111101 : 8'b10101101;
													assign node3775 = (inp[6]) ? 8'b11111101 : node3776;
														assign node3776 = (inp[12]) ? 8'b10100101 : 8'b10110100;
										assign node3780 = (inp[1]) ? node3792 : node3781;
											assign node3781 = (inp[12]) ? node3787 : node3782;
												assign node3782 = (inp[4]) ? node3784 : 8'b10101001;
													assign node3784 = (inp[3]) ? 8'b10111000 : 8'b10010101;
												assign node3787 = (inp[4]) ? node3789 : 8'b10111001;
													assign node3789 = (inp[6]) ? 8'b10111001 : 8'b10101001;
											assign node3792 = (inp[3]) ? node3800 : node3793;
												assign node3793 = (inp[6]) ? node3797 : node3794;
													assign node3794 = (inp[4]) ? 8'b10010101 : 8'b10101000;
													assign node3797 = (inp[4]) ? 8'b10101000 : 8'b10111000;
												assign node3800 = (inp[6]) ? node3804 : node3801;
													assign node3801 = (inp[12]) ? 8'b10000101 : 8'b10010100;
													assign node3804 = (inp[12]) ? 8'b10011101 : 8'b10001101;
									assign node3807 = (inp[9]) ? node3843 : node3808;
										assign node3808 = (inp[3]) ? node3826 : node3809;
											assign node3809 = (inp[12]) ? node3817 : node3810;
												assign node3810 = (inp[1]) ? 8'b10101100 : node3811;
													assign node3811 = (inp[4]) ? node3813 : 8'b10101101;
														assign node3813 = (inp[6]) ? 8'b10101100 : 8'b10110001;
												assign node3817 = (inp[1]) ? node3821 : node3818;
													assign node3818 = (inp[6]) ? 8'b10111100 : 8'b11111101;
													assign node3821 = (inp[6]) ? 8'b10111100 : node3822;
														assign node3822 = (inp[4]) ? 8'b10100100 : 8'b10111100;
											assign node3826 = (inp[1]) ? node3834 : node3827;
												assign node3827 = (inp[12]) ? node3829 : 8'b10101101;
													assign node3829 = (inp[4]) ? node3831 : 8'b11111101;
														assign node3831 = (inp[6]) ? 8'b11111101 : 8'b10101101;
												assign node3834 = (inp[6]) ? node3840 : node3835;
													assign node3835 = (inp[4]) ? node3837 : 8'b10111001;
														assign node3837 = (inp[12]) ? 8'b10100001 : 8'b10110000;
													assign node3840 = (inp[12]) ? 8'b10111001 : 8'b10101001;
										assign node3843 = (inp[3]) ? node3853 : node3844;
											assign node3844 = (inp[6]) ? node3850 : node3845;
												assign node3845 = (inp[12]) ? 8'b10000100 : node3846;
													assign node3846 = (inp[4]) ? 8'b10010001 : 8'b10001100;
												assign node3850 = (inp[12]) ? 8'b10011100 : 8'b10001100;
											assign node3853 = (inp[1]) ? node3859 : node3854;
												assign node3854 = (inp[12]) ? 8'b10011101 : node3855;
													assign node3855 = (inp[4]) ? 8'b10011100 : 8'b10001101;
												assign node3859 = (inp[4]) ? node3863 : node3860;
													assign node3860 = (inp[12]) ? 8'b10011001 : 8'b10001001;
													assign node3863 = (inp[6]) ? node3867 : node3864;
														assign node3864 = (inp[12]) ? 8'b10000001 : 8'b10010000;
														assign node3867 = (inp[12]) ? 8'b10011001 : 8'b10001001;
								assign node3870 = (inp[1]) ? node3890 : node3871;
									assign node3871 = (inp[4]) ? node3875 : node3872;
										assign node3872 = (inp[12]) ? 8'b10011101 : 8'b10001101;
										assign node3875 = (inp[3]) ? node3883 : node3876;
											assign node3876 = (inp[6]) ? node3880 : node3877;
												assign node3877 = (inp[12]) ? 8'b10000100 : 8'b10010001;
												assign node3880 = (inp[12]) ? 8'b10011100 : 8'b10001100;
											assign node3883 = (inp[12]) ? node3887 : node3884;
												assign node3884 = (inp[6]) ? 8'b10001101 : 8'b10011100;
												assign node3887 = (inp[6]) ? 8'b10011101 : 8'b10001101;
									assign node3890 = (inp[4]) ? node3894 : node3891;
										assign node3891 = (inp[12]) ? 8'b10011001 : 8'b10001001;
										assign node3894 = (inp[6]) ? node3898 : node3895;
											assign node3895 = (inp[12]) ? 8'b10000001 : 8'b10010000;
											assign node3898 = (inp[12]) ? 8'b10011001 : 8'b10001001;
							assign node3901 = (inp[1]) ? node3997 : node3902;
								assign node3902 = (inp[4]) ? node3938 : node3903;
									assign node3903 = (inp[0]) ? node3935 : node3904;
										assign node3904 = (inp[10]) ? node3920 : node3905;
											assign node3905 = (inp[9]) ? node3913 : node3906;
												assign node3906 = (inp[12]) ? node3910 : node3907;
													assign node3907 = (inp[6]) ? 8'b00001010 : 8'b00011010;
													assign node3910 = (inp[6]) ? 8'b00011010 : 8'b00001011;
												assign node3913 = (inp[12]) ? node3917 : node3914;
													assign node3914 = (inp[6]) ? 8'b10101000 : 8'b10111000;
													assign node3917 = (inp[6]) ? 8'b10111000 : 8'b10101001;
											assign node3920 = (inp[9]) ? node3928 : node3921;
												assign node3921 = (inp[6]) ? node3925 : node3922;
													assign node3922 = (inp[12]) ? 8'b10101101 : 8'b10111100;
													assign node3925 = (inp[12]) ? 8'b10111100 : 8'b10101100;
												assign node3928 = (inp[6]) ? node3932 : node3929;
													assign node3929 = (inp[12]) ? 8'b10001101 : 8'b10011100;
													assign node3932 = (inp[12]) ? 8'b10011100 : 8'b10001100;
										assign node3935 = (inp[12]) ? 8'b10011100 : 8'b10001100;
									assign node3938 = (inp[3]) ? node3974 : node3939;
										assign node3939 = (inp[0]) ? node3971 : node3940;
											assign node3940 = (inp[9]) ? node3956 : node3941;
												assign node3941 = (inp[10]) ? node3949 : node3942;
													assign node3942 = (inp[6]) ? node3946 : node3943;
														assign node3943 = (inp[12]) ? 8'b00000010 : 8'b11110111;
														assign node3946 = (inp[12]) ? 8'b11110101 : 8'b10100101;
													assign node3949 = (inp[12]) ? node3953 : node3950;
														assign node3950 = (inp[6]) ? 8'b10100001 : 8'b10110001;
														assign node3953 = (inp[6]) ? 8'b10110001 : 8'b10100100;
												assign node3956 = (inp[12]) ? node3964 : node3957;
													assign node3957 = (inp[10]) ? node3961 : node3958;
														assign node3958 = (inp[6]) ? 8'b10000101 : 8'b10010101;
														assign node3961 = (inp[6]) ? 8'b10000001 : 8'b10010001;
													assign node3964 = (inp[6]) ? node3968 : node3965;
														assign node3965 = (inp[10]) ? 8'b10000100 : 8'b10100000;
														assign node3968 = (inp[10]) ? 8'b10010001 : 8'b10010101;
											assign node3971 = (inp[12]) ? 8'b10010001 : 8'b10000001;
										assign node3974 = (inp[0]) ? node3994 : node3975;
											assign node3975 = (inp[10]) ? node3987 : node3976;
												assign node3976 = (inp[9]) ? node3982 : node3977;
													assign node3977 = (inp[6]) ? node3979 : 8'b00011010;
														assign node3979 = (inp[12]) ? 8'b00011010 : 8'b00001010;
													assign node3982 = (inp[12]) ? 8'b10101001 : node3983;
														assign node3983 = (inp[6]) ? 8'b10101000 : 8'b10111000;
												assign node3987 = (inp[9]) ? 8'b10011100 : node3988;
													assign node3988 = (inp[6]) ? 8'b10111100 : node3989;
														assign node3989 = (inp[12]) ? 8'b10101101 : 8'b10111100;
											assign node3994 = (inp[12]) ? 8'b10011100 : 8'b10001100;
								assign node3997 = (inp[0]) ? node4059 : node3998;
									assign node3998 = (inp[9]) ? node4030 : node3999;
										assign node3999 = (inp[10]) ? node4015 : node4000;
											assign node4000 = (inp[3]) ? node4008 : node4001;
												assign node4001 = (inp[6]) ? node4005 : node4002;
													assign node4002 = (inp[12]) ? 8'b00000010 : 8'b11110111;
													assign node4005 = (inp[12]) ? 8'b11110101 : 8'b10100101;
												assign node4008 = (inp[12]) ? node4012 : node4009;
													assign node4009 = (inp[6]) ? 8'b10100100 : 8'b10110100;
													assign node4012 = (inp[6]) ? 8'b10110100 : 8'b10100101;
											assign node4015 = (inp[3]) ? node4023 : node4016;
												assign node4016 = (inp[6]) ? node4020 : node4017;
													assign node4017 = (inp[12]) ? 8'b10100100 : 8'b10110001;
													assign node4020 = (inp[12]) ? 8'b10110001 : 8'b10100001;
												assign node4023 = (inp[12]) ? node4027 : node4024;
													assign node4024 = (inp[6]) ? 8'b10100000 : 8'b10110000;
													assign node4027 = (inp[6]) ? 8'b10110000 : 8'b10100001;
										assign node4030 = (inp[10]) ? node4046 : node4031;
											assign node4031 = (inp[3]) ? node4039 : node4032;
												assign node4032 = (inp[12]) ? node4036 : node4033;
													assign node4033 = (inp[6]) ? 8'b10000101 : 8'b10010101;
													assign node4036 = (inp[6]) ? 8'b10010101 : 8'b10100000;
												assign node4039 = (inp[6]) ? node4043 : node4040;
													assign node4040 = (inp[12]) ? 8'b10000101 : 8'b10010100;
													assign node4043 = (inp[12]) ? 8'b10010100 : 8'b10000100;
											assign node4046 = (inp[3]) ? node4052 : node4047;
												assign node4047 = (inp[6]) ? node4049 : 8'b10000100;
													assign node4049 = (inp[12]) ? 8'b10010001 : 8'b10000001;
												assign node4052 = (inp[6]) ? node4056 : node4053;
													assign node4053 = (inp[12]) ? 8'b10000001 : 8'b10010000;
													assign node4056 = (inp[12]) ? 8'b10010000 : 8'b10000000;
									assign node4059 = (inp[12]) ? 8'b10010000 : 8'b10000000;
		assign node4062 = (inp[4]) ? node6846 : node4063;
			assign node4063 = (inp[13]) ? node5499 : node4064;
				assign node4064 = (inp[9]) ? node4758 : node4065;
					assign node4065 = (inp[11]) ? node4299 : node4066;
						assign node4066 = (inp[6]) ? node4180 : node4067;
							assign node4067 = (inp[0]) ? node4157 : node4068;
								assign node4068 = (inp[2]) ? node4110 : node4069;
									assign node4069 = (inp[5]) ? node4083 : node4070;
										assign node4070 = (inp[8]) ? node4078 : node4071;
											assign node4071 = (inp[10]) ? 8'b00111010 : node4072;
												assign node4072 = (inp[3]) ? 8'b00111110 : node4073;
													assign node4073 = (inp[1]) ? 8'b00111110 : 8'b01111111;
											assign node4078 = (inp[3]) ? 8'b00111010 : node4079;
												assign node4079 = (inp[1]) ? 8'b00111010 : 8'b00111011;
										assign node4083 = (inp[10]) ? node4093 : node4084;
											assign node4084 = (inp[8]) ? node4086 : 8'b01111111;
												assign node4086 = (inp[1]) ? node4090 : node4087;
													assign node4087 = (inp[3]) ? 8'b00111010 : 8'b00111011;
													assign node4090 = (inp[3]) ? 8'b00111011 : 8'b00111010;
											assign node4093 = (inp[8]) ? node4101 : node4094;
												assign node4094 = (inp[1]) ? node4098 : node4095;
													assign node4095 = (inp[3]) ? 8'b00111010 : 8'b00111011;
													assign node4098 = (inp[3]) ? 8'b00111011 : 8'b00111010;
												assign node4101 = (inp[12]) ? 8'b00111110 : node4102;
													assign node4102 = (inp[3]) ? node4106 : node4103;
														assign node4103 = (inp[1]) ? 8'b00111110 : 8'b01111111;
														assign node4106 = (inp[1]) ? 8'b01111111 : 8'b00111110;
									assign node4110 = (inp[8]) ? node4130 : node4111;
										assign node4111 = (inp[10]) ? node4121 : node4112;
											assign node4112 = (inp[3]) ? node4116 : node4113;
												assign node4113 = (inp[1]) ? 8'b00101110 : 8'b00101111;
												assign node4116 = (inp[1]) ? node4118 : 8'b00101110;
													assign node4118 = (inp[5]) ? 8'b00101111 : 8'b00101110;
											assign node4121 = (inp[5]) ? node4127 : node4122;
												assign node4122 = (inp[1]) ? 8'b00101010 : node4123;
													assign node4123 = (inp[12]) ? 8'b00101010 : 8'b00101011;
												assign node4127 = (inp[1]) ? 8'b00101011 : 8'b00101010;
										assign node4130 = (inp[10]) ? node4140 : node4131;
											assign node4131 = (inp[1]) ? node4135 : node4132;
												assign node4132 = (inp[3]) ? 8'b00101010 : 8'b00101011;
												assign node4135 = (inp[3]) ? node4137 : 8'b00101010;
													assign node4137 = (inp[5]) ? 8'b00101011 : 8'b00101010;
											assign node4140 = (inp[5]) ? node4144 : node4141;
												assign node4141 = (inp[3]) ? 8'b00101010 : 8'b00101011;
												assign node4144 = (inp[12]) ? node4150 : node4145;
													assign node4145 = (inp[1]) ? 8'b00101111 : node4146;
														assign node4146 = (inp[3]) ? 8'b00101110 : 8'b00101111;
													assign node4150 = (inp[1]) ? node4154 : node4151;
														assign node4151 = (inp[3]) ? 8'b00101110 : 8'b00101111;
														assign node4154 = (inp[3]) ? 8'b00101111 : 8'b00101110;
								assign node4157 = (inp[10]) ? node4165 : node4158;
									assign node4158 = (inp[3]) ? node4160 : 8'b01111111;
										assign node4160 = (inp[1]) ? node4162 : 8'b00111110;
											assign node4162 = (inp[5]) ? 8'b01111111 : 8'b00111110;
									assign node4165 = (inp[3]) ? node4171 : node4166;
										assign node4166 = (inp[8]) ? node4168 : 8'b00111011;
											assign node4168 = (inp[5]) ? 8'b01111111 : 8'b00111011;
										assign node4171 = (inp[5]) ? node4173 : 8'b00111010;
											assign node4173 = (inp[1]) ? node4177 : node4174;
												assign node4174 = (inp[8]) ? 8'b00111110 : 8'b00111010;
												assign node4177 = (inp[8]) ? 8'b01111111 : 8'b00111011;
							assign node4180 = (inp[5]) ? node4204 : node4181;
								assign node4181 = (inp[10]) ? node4197 : node4182;
									assign node4182 = (inp[3]) ? node4192 : node4183;
										assign node4183 = (inp[0]) ? 8'b00101111 : node4184;
											assign node4184 = (inp[1]) ? node4188 : node4185;
												assign node4185 = (inp[8]) ? 8'b00101011 : 8'b00101111;
												assign node4188 = (inp[8]) ? 8'b00101010 : 8'b00101110;
										assign node4192 = (inp[0]) ? 8'b00101110 : node4193;
											assign node4193 = (inp[8]) ? 8'b00101010 : 8'b00101110;
									assign node4197 = (inp[3]) ? 8'b00101010 : node4198;
										assign node4198 = (inp[0]) ? 8'b00101011 : node4199;
											assign node4199 = (inp[1]) ? 8'b00101010 : 8'b00101011;
								assign node4204 = (inp[2]) ? node4252 : node4205;
									assign node4205 = (inp[10]) ? node4233 : node4206;
										assign node4206 = (inp[8]) ? node4216 : node4207;
											assign node4207 = (inp[1]) ? node4211 : node4208;
												assign node4208 = (inp[3]) ? 8'b00101110 : 8'b00101111;
												assign node4211 = (inp[12]) ? node4213 : 8'b00101111;
													assign node4213 = (inp[3]) ? 8'b00101111 : 8'b00101110;
											assign node4216 = (inp[0]) ? node4228 : node4217;
												assign node4217 = (inp[12]) ? node4223 : node4218;
													assign node4218 = (inp[3]) ? 8'b00101011 : node4219;
														assign node4219 = (inp[1]) ? 8'b00101010 : 8'b00101011;
													assign node4223 = (inp[1]) ? 8'b00101011 : node4224;
														assign node4224 = (inp[3]) ? 8'b00101010 : 8'b00101011;
												assign node4228 = (inp[3]) ? node4230 : 8'b00101111;
													assign node4230 = (inp[1]) ? 8'b00101111 : 8'b00101110;
										assign node4233 = (inp[8]) ? node4243 : node4234;
											assign node4234 = (inp[1]) ? node4238 : node4235;
												assign node4235 = (inp[3]) ? 8'b00101010 : 8'b00101011;
												assign node4238 = (inp[0]) ? 8'b00101011 : node4239;
													assign node4239 = (inp[3]) ? 8'b00101011 : 8'b00101010;
											assign node4243 = (inp[0]) ? 8'b00101111 : node4244;
												assign node4244 = (inp[1]) ? node4248 : node4245;
													assign node4245 = (inp[3]) ? 8'b00101110 : 8'b00101111;
													assign node4248 = (inp[3]) ? 8'b00101111 : 8'b00101110;
									assign node4252 = (inp[0]) ? node4284 : node4253;
										assign node4253 = (inp[3]) ? node4269 : node4254;
											assign node4254 = (inp[1]) ? node4260 : node4255;
												assign node4255 = (inp[8]) ? 8'b00111011 : node4256;
													assign node4256 = (inp[10]) ? 8'b00111011 : 8'b01111111;
												assign node4260 = (inp[12]) ? node4262 : 8'b00111010;
													assign node4262 = (inp[10]) ? node4266 : node4263;
														assign node4263 = (inp[8]) ? 8'b00111010 : 8'b00111110;
														assign node4266 = (inp[8]) ? 8'b00111110 : 8'b00111010;
											assign node4269 = (inp[1]) ? node4277 : node4270;
												assign node4270 = (inp[8]) ? node4274 : node4271;
													assign node4271 = (inp[10]) ? 8'b00111010 : 8'b00111110;
													assign node4274 = (inp[10]) ? 8'b00111110 : 8'b00111010;
												assign node4277 = (inp[8]) ? node4281 : node4278;
													assign node4278 = (inp[10]) ? 8'b00111011 : 8'b01111111;
													assign node4281 = (inp[10]) ? 8'b01111111 : 8'b00111011;
										assign node4284 = (inp[1]) ? node4294 : node4285;
											assign node4285 = (inp[3]) ? node4289 : node4286;
												assign node4286 = (inp[8]) ? 8'b01111111 : 8'b00111011;
												assign node4289 = (inp[10]) ? node4291 : 8'b00111110;
													assign node4291 = (inp[8]) ? 8'b00111110 : 8'b00111010;
											assign node4294 = (inp[8]) ? 8'b01111111 : node4295;
												assign node4295 = (inp[10]) ? 8'b00111011 : 8'b01111111;
						assign node4299 = (inp[8]) ? node4511 : node4300;
							assign node4300 = (inp[10]) ? node4412 : node4301;
								assign node4301 = (inp[1]) ? node4351 : node4302;
									assign node4302 = (inp[3]) ? node4326 : node4303;
										assign node4303 = (inp[2]) ? node4311 : node4304;
											assign node4304 = (inp[6]) ? node4308 : node4305;
												assign node4305 = (inp[12]) ? 8'b01111111 : 8'b00101111;
												assign node4308 = (inp[12]) ? 8'b00101111 : 8'b00111110;
											assign node4311 = (inp[5]) ? node4319 : node4312;
												assign node4312 = (inp[12]) ? node4314 : 8'b00111110;
													assign node4314 = (inp[0]) ? node4316 : 8'b00101111;
														assign node4316 = (inp[6]) ? 8'b00101111 : 8'b00111110;
												assign node4319 = (inp[12]) ? 8'b00111110 : node4320;
													assign node4320 = (inp[6]) ? 8'b00101110 : node4321;
														assign node4321 = (inp[0]) ? 8'b00101110 : 8'b00111110;
										assign node4326 = (inp[12]) ? node4336 : node4327;
											assign node4327 = (inp[6]) ? node4331 : node4328;
												assign node4328 = (inp[2]) ? 8'b00111011 : 8'b00101110;
												assign node4331 = (inp[2]) ? node4333 : 8'b00111011;
													assign node4333 = (inp[5]) ? 8'b00101011 : 8'b00111011;
											assign node4336 = (inp[5]) ? node4342 : node4337;
												assign node4337 = (inp[6]) ? 8'b00101110 : node4338;
													assign node4338 = (inp[0]) ? 8'b00111110 : 8'b00101110;
												assign node4342 = (inp[2]) ? node4346 : node4343;
													assign node4343 = (inp[6]) ? 8'b00101110 : 8'b00111110;
													assign node4346 = (inp[0]) ? 8'b00111011 : node4347;
														assign node4347 = (inp[6]) ? 8'b00111011 : 8'b00101110;
									assign node4351 = (inp[0]) ? node4379 : node4352;
										assign node4352 = (inp[6]) ? node4364 : node4353;
											assign node4353 = (inp[2]) ? node4359 : node4354;
												assign node4354 = (inp[12]) ? node4356 : 8'b00101110;
													assign node4356 = (inp[3]) ? 8'b00111011 : 8'b00111110;
												assign node4359 = (inp[12]) ? 8'b00101110 : node4360;
													assign node4360 = (inp[3]) ? 8'b00111010 : 8'b00111011;
											assign node4364 = (inp[5]) ? node4366 : 8'b00111011;
												assign node4366 = (inp[3]) ? node4374 : node4367;
													assign node4367 = (inp[12]) ? node4371 : node4368;
														assign node4368 = (inp[2]) ? 8'b00101011 : 8'b00111011;
														assign node4371 = (inp[2]) ? 8'b00111011 : 8'b00101110;
													assign node4374 = (inp[2]) ? 8'b00111010 : node4375;
														assign node4375 = (inp[12]) ? 8'b00101011 : 8'b00111010;
										assign node4379 = (inp[5]) ? node4401 : node4380;
											assign node4380 = (inp[3]) ? node4392 : node4381;
												assign node4381 = (inp[12]) ? node4387 : node4382;
													assign node4382 = (inp[6]) ? 8'b00111010 : node4383;
														assign node4383 = (inp[2]) ? 8'b00101010 : 8'b00101011;
													assign node4387 = (inp[6]) ? 8'b00101011 : node4388;
														assign node4388 = (inp[2]) ? 8'b00111010 : 8'b00111011;
												assign node4392 = (inp[12]) ? node4398 : node4393;
													assign node4393 = (inp[6]) ? 8'b00111011 : node4394;
														assign node4394 = (inp[2]) ? 8'b00101011 : 8'b00101110;
													assign node4398 = (inp[6]) ? 8'b00101110 : 8'b00111011;
											assign node4401 = (inp[2]) ? node4409 : node4402;
												assign node4402 = (inp[6]) ? node4406 : node4403;
													assign node4403 = (inp[12]) ? 8'b00111011 : 8'b00101011;
													assign node4406 = (inp[12]) ? 8'b00101011 : 8'b00111010;
												assign node4409 = (inp[12]) ? 8'b00111010 : 8'b00101010;
								assign node4412 = (inp[1]) ? node4454 : node4413;
									assign node4413 = (inp[3]) ? node4433 : node4414;
										assign node4414 = (inp[2]) ? node4422 : node4415;
											assign node4415 = (inp[6]) ? node4419 : node4416;
												assign node4416 = (inp[12]) ? 8'b00111011 : 8'b00101011;
												assign node4419 = (inp[12]) ? 8'b00101011 : 8'b00111010;
											assign node4422 = (inp[12]) ? node4428 : node4423;
												assign node4423 = (inp[5]) ? 8'b00101010 : node4424;
													assign node4424 = (inp[0]) ? 8'b00101010 : 8'b00111010;
												assign node4428 = (inp[5]) ? 8'b00111010 : node4429;
													assign node4429 = (inp[6]) ? 8'b00101011 : 8'b00111010;
										assign node4433 = (inp[12]) ? node4445 : node4434;
											assign node4434 = (inp[6]) ? node4440 : node4435;
												assign node4435 = (inp[2]) ? node4437 : 8'b00101010;
													assign node4437 = (inp[0]) ? 8'b00001111 : 8'b00011111;
												assign node4440 = (inp[2]) ? node4442 : 8'b00011111;
													assign node4442 = (inp[5]) ? 8'b00001111 : 8'b00011111;
											assign node4445 = (inp[5]) ? node4447 : 8'b00101010;
												assign node4447 = (inp[2]) ? node4451 : node4448;
													assign node4448 = (inp[6]) ? 8'b00101010 : 8'b00111010;
													assign node4451 = (inp[0]) ? 8'b00011111 : 8'b00101010;
									assign node4454 = (inp[6]) ? node4482 : node4455;
										assign node4455 = (inp[0]) ? node4469 : node4456;
											assign node4456 = (inp[12]) ? node4466 : node4457;
												assign node4457 = (inp[2]) ? node4463 : node4458;
													assign node4458 = (inp[5]) ? node4460 : 8'b00101010;
														assign node4460 = (inp[3]) ? 8'b00001111 : 8'b00101010;
													assign node4463 = (inp[3]) ? 8'b00011110 : 8'b00011111;
												assign node4466 = (inp[2]) ? 8'b00101010 : 8'b00111010;
											assign node4469 = (inp[12]) ? node4475 : node4470;
												assign node4470 = (inp[2]) ? 8'b00001110 : node4471;
													assign node4471 = (inp[3]) ? 8'b00101010 : 8'b00001111;
												assign node4475 = (inp[2]) ? node4477 : 8'b00011111;
													assign node4477 = (inp[5]) ? 8'b00011110 : node4478;
														assign node4478 = (inp[3]) ? 8'b00011111 : 8'b00011110;
										assign node4482 = (inp[2]) ? node4490 : node4483;
											assign node4483 = (inp[12]) ? 8'b00001111 : node4484;
												assign node4484 = (inp[0]) ? node4486 : 8'b00011111;
													assign node4486 = (inp[3]) ? 8'b00011111 : 8'b00011110;
											assign node4490 = (inp[3]) ? node4504 : node4491;
												assign node4491 = (inp[0]) ? node4497 : node4492;
													assign node4492 = (inp[5]) ? node4494 : 8'b00011111;
														assign node4494 = (inp[12]) ? 8'b00011111 : 8'b00001111;
													assign node4497 = (inp[5]) ? node4501 : node4498;
														assign node4498 = (inp[12]) ? 8'b00001111 : 8'b00011110;
														assign node4501 = (inp[12]) ? 8'b00011110 : 8'b00001110;
												assign node4504 = (inp[5]) ? node4508 : node4505;
													assign node4505 = (inp[12]) ? 8'b00101010 : 8'b00011111;
													assign node4508 = (inp[12]) ? 8'b00011110 : 8'b00001110;
							assign node4511 = (inp[5]) ? node4631 : node4512;
								assign node4512 = (inp[0]) ? node4546 : node4513;
									assign node4513 = (inp[12]) ? node4531 : node4514;
										assign node4514 = (inp[6]) ? node4526 : node4515;
											assign node4515 = (inp[2]) ? node4521 : node4516;
												assign node4516 = (inp[3]) ? 8'b00101010 : node4517;
													assign node4517 = (inp[1]) ? 8'b00101010 : 8'b00101011;
												assign node4521 = (inp[1]) ? 8'b00011111 : node4522;
													assign node4522 = (inp[10]) ? 8'b00011111 : 8'b00111010;
											assign node4526 = (inp[3]) ? 8'b00011111 : node4527;
												assign node4527 = (inp[1]) ? 8'b00011111 : 8'b00111010;
										assign node4531 = (inp[2]) ? node4541 : node4532;
											assign node4532 = (inp[6]) ? node4536 : node4533;
												assign node4533 = (inp[1]) ? 8'b00111010 : 8'b00111011;
												assign node4536 = (inp[3]) ? 8'b00101010 : node4537;
													assign node4537 = (inp[1]) ? 8'b00101010 : 8'b00101011;
											assign node4541 = (inp[1]) ? 8'b00101010 : node4542;
												assign node4542 = (inp[3]) ? 8'b00101010 : 8'b00101011;
									assign node4546 = (inp[10]) ? node4588 : node4547;
										assign node4547 = (inp[1]) ? node4571 : node4548;
											assign node4548 = (inp[3]) ? node4558 : node4549;
												assign node4549 = (inp[6]) ? 8'b00001111 : node4550;
													assign node4550 = (inp[12]) ? node4554 : node4551;
														assign node4551 = (inp[2]) ? 8'b00001110 : 8'b00001111;
														assign node4554 = (inp[2]) ? 8'b00011110 : 8'b00011111;
												assign node4558 = (inp[2]) ? node4566 : node4559;
													assign node4559 = (inp[6]) ? node4563 : node4560;
														assign node4560 = (inp[12]) ? 8'b00011110 : 8'b00001110;
														assign node4563 = (inp[12]) ? 8'b00001110 : 8'b00011011;
													assign node4566 = (inp[6]) ? 8'b00011011 : node4567;
														assign node4567 = (inp[12]) ? 8'b00011011 : 8'b00001011;
											assign node4571 = (inp[3]) ? node4579 : node4572;
												assign node4572 = (inp[12]) ? node4574 : 8'b00011010;
													assign node4574 = (inp[6]) ? 8'b00001011 : node4575;
														assign node4575 = (inp[2]) ? 8'b00011010 : 8'b00011011;
												assign node4579 = (inp[12]) ? node4585 : node4580;
													assign node4580 = (inp[6]) ? 8'b00011011 : node4581;
														assign node4581 = (inp[2]) ? 8'b00001011 : 8'b00001110;
													assign node4585 = (inp[2]) ? 8'b00001110 : 8'b00011110;
										assign node4588 = (inp[1]) ? node4608 : node4589;
											assign node4589 = (inp[3]) ? node4601 : node4590;
												assign node4590 = (inp[12]) ? node4596 : node4591;
													assign node4591 = (inp[6]) ? 8'b00111010 : node4592;
														assign node4592 = (inp[2]) ? 8'b00101010 : 8'b00101011;
													assign node4596 = (inp[6]) ? 8'b00101011 : node4597;
														assign node4597 = (inp[2]) ? 8'b00111010 : 8'b00111011;
												assign node4601 = (inp[6]) ? node4605 : node4602;
													assign node4602 = (inp[12]) ? 8'b00011111 : 8'b00101010;
													assign node4605 = (inp[2]) ? 8'b00101010 : 8'b00011111;
											assign node4608 = (inp[3]) ? node4622 : node4609;
												assign node4609 = (inp[2]) ? node4615 : node4610;
													assign node4610 = (inp[6]) ? node4612 : 8'b00001111;
														assign node4612 = (inp[12]) ? 8'b00001111 : 8'b00011110;
													assign node4615 = (inp[6]) ? node4619 : node4616;
														assign node4616 = (inp[12]) ? 8'b00011110 : 8'b00001110;
														assign node4619 = (inp[12]) ? 8'b00001111 : 8'b00011110;
												assign node4622 = (inp[2]) ? node4626 : node4623;
													assign node4623 = (inp[12]) ? 8'b00111010 : 8'b00101010;
													assign node4626 = (inp[12]) ? node4628 : 8'b00011111;
														assign node4628 = (inp[6]) ? 8'b00101010 : 8'b00011111;
								assign node4631 = (inp[0]) ? node4727 : node4632;
									assign node4632 = (inp[10]) ? node4680 : node4633;
										assign node4633 = (inp[1]) ? node4659 : node4634;
											assign node4634 = (inp[3]) ? node4648 : node4635;
												assign node4635 = (inp[12]) ? node4641 : node4636;
													assign node4636 = (inp[2]) ? node4638 : 8'b00111010;
														assign node4638 = (inp[6]) ? 8'b00101010 : 8'b00111010;
													assign node4641 = (inp[2]) ? node4645 : node4642;
														assign node4642 = (inp[6]) ? 8'b00101011 : 8'b00111011;
														assign node4645 = (inp[6]) ? 8'b00111010 : 8'b00101011;
												assign node4648 = (inp[6]) ? node4654 : node4649;
													assign node4649 = (inp[2]) ? 8'b00101010 : node4650;
														assign node4650 = (inp[12]) ? 8'b00111010 : 8'b00101010;
													assign node4654 = (inp[2]) ? node4656 : 8'b00011111;
														assign node4656 = (inp[12]) ? 8'b00011111 : 8'b00001111;
											assign node4659 = (inp[3]) ? node4669 : node4660;
												assign node4660 = (inp[6]) ? node4666 : node4661;
													assign node4661 = (inp[2]) ? node4663 : 8'b00101010;
														assign node4663 = (inp[12]) ? 8'b00101010 : 8'b00011111;
													assign node4666 = (inp[2]) ? 8'b00001111 : 8'b00011111;
												assign node4669 = (inp[2]) ? node4673 : node4670;
													assign node4670 = (inp[12]) ? 8'b00011111 : 8'b00001111;
													assign node4673 = (inp[6]) ? node4677 : node4674;
														assign node4674 = (inp[12]) ? 8'b00001111 : 8'b00011110;
														assign node4677 = (inp[12]) ? 8'b00011110 : 8'b00001110;
										assign node4680 = (inp[3]) ? node4708 : node4681;
											assign node4681 = (inp[1]) ? node4695 : node4682;
												assign node4682 = (inp[6]) ? node4690 : node4683;
													assign node4683 = (inp[12]) ? node4687 : node4684;
														assign node4684 = (inp[2]) ? 8'b00011110 : 8'b00001111;
														assign node4687 = (inp[2]) ? 8'b00001111 : 8'b00011111;
													assign node4690 = (inp[2]) ? node4692 : 8'b00011110;
														assign node4692 = (inp[12]) ? 8'b00011110 : 8'b00001110;
												assign node4695 = (inp[2]) ? node4701 : node4696;
													assign node4696 = (inp[12]) ? node4698 : 8'b00001110;
														assign node4698 = (inp[6]) ? 8'b00001110 : 8'b00011110;
													assign node4701 = (inp[6]) ? node4705 : node4702;
														assign node4702 = (inp[12]) ? 8'b00001110 : 8'b00011011;
														assign node4705 = (inp[12]) ? 8'b00011011 : 8'b00001011;
											assign node4708 = (inp[1]) ? node4720 : node4709;
												assign node4709 = (inp[12]) ? node4715 : node4710;
													assign node4710 = (inp[6]) ? 8'b00011011 : node4711;
														assign node4711 = (inp[2]) ? 8'b00011011 : 8'b00001110;
													assign node4715 = (inp[2]) ? node4717 : 8'b00001110;
														assign node4717 = (inp[6]) ? 8'b00011011 : 8'b00001110;
												assign node4720 = (inp[6]) ? 8'b00011010 : node4721;
													assign node4721 = (inp[12]) ? node4723 : 8'b00001011;
														assign node4723 = (inp[2]) ? 8'b00001011 : 8'b00011011;
									assign node4727 = (inp[1]) ? node4747 : node4728;
										assign node4728 = (inp[3]) ? node4736 : node4729;
											assign node4729 = (inp[12]) ? 8'b00011110 : node4730;
												assign node4730 = (inp[2]) ? 8'b00001110 : node4731;
													assign node4731 = (inp[6]) ? 8'b00011110 : 8'b00001111;
											assign node4736 = (inp[2]) ? node4744 : node4737;
												assign node4737 = (inp[6]) ? node4741 : node4738;
													assign node4738 = (inp[12]) ? 8'b00011110 : 8'b00001110;
													assign node4741 = (inp[12]) ? 8'b00001110 : 8'b00011011;
												assign node4744 = (inp[12]) ? 8'b00011011 : 8'b00001011;
										assign node4747 = (inp[2]) ? node4755 : node4748;
											assign node4748 = (inp[6]) ? node4752 : node4749;
												assign node4749 = (inp[12]) ? 8'b00011011 : 8'b00001011;
												assign node4752 = (inp[12]) ? 8'b00001011 : 8'b00011010;
											assign node4755 = (inp[12]) ? 8'b00011010 : 8'b00001010;
					assign node4758 = (inp[8]) ? node5128 : node4759;
						assign node4759 = (inp[10]) ? node4931 : node4760;
							assign node4760 = (inp[11]) ? node4818 : node4761;
								assign node4761 = (inp[6]) ? node4789 : node4762;
									assign node4762 = (inp[2]) ? node4774 : node4763;
										assign node4763 = (inp[3]) ? node4769 : node4764;
											assign node4764 = (inp[1]) ? node4766 : 8'b00011111;
												assign node4766 = (inp[0]) ? 8'b00011111 : 8'b00011110;
											assign node4769 = (inp[1]) ? node4771 : 8'b00011110;
												assign node4771 = (inp[5]) ? 8'b00011111 : 8'b00011110;
										assign node4774 = (inp[0]) ? node4782 : node4775;
											assign node4775 = (inp[1]) ? node4779 : node4776;
												assign node4776 = (inp[3]) ? 8'b00001110 : 8'b00001111;
												assign node4779 = (inp[3]) ? 8'b00001111 : 8'b00001110;
											assign node4782 = (inp[3]) ? node4784 : 8'b00011111;
												assign node4784 = (inp[1]) ? node4786 : 8'b00011110;
													assign node4786 = (inp[5]) ? 8'b00011111 : 8'b00011110;
									assign node4789 = (inp[5]) ? node4797 : node4790;
										assign node4790 = (inp[3]) ? 8'b00001110 : node4791;
											assign node4791 = (inp[1]) ? node4793 : 8'b00001111;
												assign node4793 = (inp[0]) ? 8'b00001111 : 8'b00001110;
										assign node4797 = (inp[2]) ? node4809 : node4798;
											assign node4798 = (inp[0]) ? node4804 : node4799;
												assign node4799 = (inp[3]) ? 8'b00001111 : node4800;
													assign node4800 = (inp[1]) ? 8'b00001110 : 8'b00001111;
												assign node4804 = (inp[3]) ? node4806 : 8'b00001111;
													assign node4806 = (inp[1]) ? 8'b00001111 : 8'b00001110;
											assign node4809 = (inp[3]) ? node4815 : node4810;
												assign node4810 = (inp[0]) ? 8'b00011111 : node4811;
													assign node4811 = (inp[12]) ? 8'b00011111 : 8'b00011110;
												assign node4815 = (inp[1]) ? 8'b00011111 : 8'b00011110;
								assign node4818 = (inp[1]) ? node4866 : node4819;
									assign node4819 = (inp[3]) ? node4843 : node4820;
										assign node4820 = (inp[2]) ? node4828 : node4821;
											assign node4821 = (inp[6]) ? node4825 : node4822;
												assign node4822 = (inp[12]) ? 8'b00011111 : 8'b00001111;
												assign node4825 = (inp[12]) ? 8'b00001111 : 8'b00011110;
											assign node4828 = (inp[12]) ? node4834 : node4829;
												assign node4829 = (inp[0]) ? 8'b00001110 : node4830;
													assign node4830 = (inp[6]) ? 8'b00001110 : 8'b00011110;
												assign node4834 = (inp[5]) ? node4838 : node4835;
													assign node4835 = (inp[6]) ? 8'b00001111 : 8'b00011110;
													assign node4838 = (inp[6]) ? 8'b00011110 : node4839;
														assign node4839 = (inp[0]) ? 8'b00011110 : 8'b00001111;
										assign node4843 = (inp[2]) ? node4851 : node4844;
											assign node4844 = (inp[6]) ? node4848 : node4845;
												assign node4845 = (inp[12]) ? 8'b00011110 : 8'b00001110;
												assign node4848 = (inp[12]) ? 8'b00001110 : 8'b00011011;
											assign node4851 = (inp[12]) ? node4859 : node4852;
												assign node4852 = (inp[0]) ? 8'b00001011 : node4853;
													assign node4853 = (inp[6]) ? node4855 : 8'b00011011;
														assign node4855 = (inp[5]) ? 8'b00001011 : 8'b00011011;
												assign node4859 = (inp[5]) ? node4861 : 8'b00001110;
													assign node4861 = (inp[6]) ? 8'b00011011 : node4862;
														assign node4862 = (inp[0]) ? 8'b00011011 : 8'b00001110;
									assign node4866 = (inp[0]) ? node4906 : node4867;
										assign node4867 = (inp[12]) ? node4885 : node4868;
											assign node4868 = (inp[2]) ? node4876 : node4869;
												assign node4869 = (inp[6]) ? 8'b00011011 : node4870;
													assign node4870 = (inp[5]) ? node4872 : 8'b00001110;
														assign node4872 = (inp[3]) ? 8'b00001011 : 8'b00001110;
												assign node4876 = (inp[6]) ? node4882 : node4877;
													assign node4877 = (inp[3]) ? node4879 : 8'b00011011;
														assign node4879 = (inp[5]) ? 8'b00011010 : 8'b00011011;
													assign node4882 = (inp[3]) ? 8'b00001010 : 8'b00001011;
											assign node4885 = (inp[5]) ? node4891 : node4886;
												assign node4886 = (inp[2]) ? 8'b00001110 : node4887;
													assign node4887 = (inp[6]) ? 8'b00001110 : 8'b00011110;
												assign node4891 = (inp[3]) ? node4899 : node4892;
													assign node4892 = (inp[6]) ? node4896 : node4893;
														assign node4893 = (inp[2]) ? 8'b00001110 : 8'b00011110;
														assign node4896 = (inp[2]) ? 8'b00011011 : 8'b00001110;
													assign node4899 = (inp[2]) ? node4903 : node4900;
														assign node4900 = (inp[6]) ? 8'b00001011 : 8'b00011011;
														assign node4903 = (inp[6]) ? 8'b00011010 : 8'b00001011;
										assign node4906 = (inp[2]) ? node4920 : node4907;
											assign node4907 = (inp[12]) ? node4917 : node4908;
												assign node4908 = (inp[6]) ? node4914 : node4909;
													assign node4909 = (inp[3]) ? node4911 : 8'b00001011;
														assign node4911 = (inp[5]) ? 8'b00001011 : 8'b00001110;
													assign node4914 = (inp[3]) ? 8'b00011011 : 8'b00011010;
												assign node4917 = (inp[6]) ? 8'b00001011 : 8'b00011011;
											assign node4920 = (inp[12]) ? node4926 : node4921;
												assign node4921 = (inp[5]) ? 8'b00001010 : node4922;
													assign node4922 = (inp[3]) ? 8'b00001011 : 8'b00011010;
												assign node4926 = (inp[5]) ? 8'b00011010 : node4927;
													assign node4927 = (inp[6]) ? 8'b00001011 : 8'b00011010;
							assign node4931 = (inp[1]) ? node5013 : node4932;
								assign node4932 = (inp[3]) ? node4972 : node4933;
									assign node4933 = (inp[11]) ? node4945 : node4934;
										assign node4934 = (inp[6]) ? node4940 : node4935;
											assign node4935 = (inp[0]) ? 8'b00011011 : node4936;
												assign node4936 = (inp[2]) ? 8'b00001011 : 8'b00011011;
											assign node4940 = (inp[2]) ? node4942 : 8'b00001011;
												assign node4942 = (inp[5]) ? 8'b00011011 : 8'b00001011;
										assign node4945 = (inp[12]) ? node4957 : node4946;
											assign node4946 = (inp[6]) ? node4952 : node4947;
												assign node4947 = (inp[2]) ? node4949 : 8'b00001011;
													assign node4949 = (inp[0]) ? 8'b00001010 : 8'b00011010;
												assign node4952 = (inp[2]) ? node4954 : 8'b00011010;
													assign node4954 = (inp[5]) ? 8'b00001010 : 8'b00011010;
											assign node4957 = (inp[5]) ? node4963 : node4958;
												assign node4958 = (inp[0]) ? node4960 : 8'b00001011;
													assign node4960 = (inp[2]) ? 8'b00001011 : 8'b00011011;
												assign node4963 = (inp[2]) ? node4967 : node4964;
													assign node4964 = (inp[0]) ? 8'b00001011 : 8'b00011011;
													assign node4967 = (inp[6]) ? 8'b00011010 : node4968;
														assign node4968 = (inp[0]) ? 8'b00011010 : 8'b00001011;
									assign node4972 = (inp[2]) ? node4984 : node4973;
										assign node4973 = (inp[6]) ? node4979 : node4974;
											assign node4974 = (inp[11]) ? node4976 : 8'b00011010;
												assign node4976 = (inp[12]) ? 8'b00011010 : 8'b00001010;
											assign node4979 = (inp[12]) ? 8'b00000010 : node4980;
												assign node4980 = (inp[11]) ? 8'b11110111 : 8'b10000010;
										assign node4984 = (inp[11]) ? node5000 : node4985;
											assign node4985 = (inp[0]) ? node4993 : node4986;
												assign node4986 = (inp[12]) ? node4988 : 8'b10000010;
													assign node4988 = (inp[5]) ? node4990 : 8'b00000010;
														assign node4990 = (inp[6]) ? 8'b10010000 : 8'b00000010;
												assign node4993 = (inp[5]) ? 8'b10010000 : node4994;
													assign node4994 = (inp[6]) ? node4996 : 8'b10010000;
														assign node4996 = (inp[12]) ? 8'b00000010 : 8'b10000010;
											assign node5000 = (inp[12]) ? node5010 : node5001;
												assign node5001 = (inp[5]) ? node5005 : node5002;
													assign node5002 = (inp[6]) ? 8'b11110111 : 8'b10100101;
													assign node5005 = (inp[6]) ? 8'b10100101 : node5006;
														assign node5006 = (inp[0]) ? 8'b10100101 : 8'b11110111;
												assign node5010 = (inp[5]) ? 8'b11110101 : 8'b00000010;
								assign node5013 = (inp[11]) ? node5061 : node5014;
									assign node5014 = (inp[5]) ? node5036 : node5015;
										assign node5015 = (inp[6]) ? node5029 : node5016;
											assign node5016 = (inp[2]) ? node5022 : node5017;
												assign node5017 = (inp[3]) ? 8'b00011010 : node5018;
													assign node5018 = (inp[0]) ? 8'b10011001 : 8'b00011010;
												assign node5022 = (inp[0]) ? node5026 : node5023;
													assign node5023 = (inp[12]) ? 8'b00000010 : 8'b10000010;
													assign node5026 = (inp[3]) ? 8'b10010000 : 8'b10010001;
											assign node5029 = (inp[12]) ? node5031 : 8'b10000010;
												assign node5031 = (inp[3]) ? 8'b00000010 : node5032;
													assign node5032 = (inp[0]) ? 8'b10000001 : 8'b00000010;
										assign node5036 = (inp[0]) ? node5056 : node5037;
											assign node5037 = (inp[3]) ? node5047 : node5038;
												assign node5038 = (inp[2]) ? node5042 : node5039;
													assign node5039 = (inp[6]) ? 8'b00000010 : 8'b00011010;
													assign node5042 = (inp[6]) ? 8'b10010000 : node5043;
														assign node5043 = (inp[12]) ? 8'b00000010 : 8'b10000010;
												assign node5047 = (inp[12]) ? node5049 : 8'b10011001;
													assign node5049 = (inp[2]) ? node5053 : node5050;
														assign node5050 = (inp[6]) ? 8'b10000001 : 8'b10011001;
														assign node5053 = (inp[6]) ? 8'b10010001 : 8'b10000001;
											assign node5056 = (inp[2]) ? 8'b10010001 : node5057;
												assign node5057 = (inp[6]) ? 8'b10000001 : 8'b10011001;
									assign node5061 = (inp[5]) ? node5093 : node5062;
										assign node5062 = (inp[0]) ? node5074 : node5063;
											assign node5063 = (inp[12]) ? node5069 : node5064;
												assign node5064 = (inp[6]) ? 8'b11110111 : node5065;
													assign node5065 = (inp[2]) ? 8'b11110111 : 8'b00001010;
												assign node5069 = (inp[2]) ? 8'b00000010 : node5070;
													assign node5070 = (inp[6]) ? 8'b00000010 : 8'b00011010;
											assign node5074 = (inp[2]) ? node5084 : node5075;
												assign node5075 = (inp[3]) ? node5079 : node5076;
													assign node5076 = (inp[12]) ? 8'b11111101 : 8'b10101101;
													assign node5079 = (inp[6]) ? node5081 : 8'b00001010;
														assign node5081 = (inp[12]) ? 8'b00000010 : 8'b11110111;
												assign node5084 = (inp[3]) ? node5088 : node5085;
													assign node5085 = (inp[6]) ? 8'b10100101 : 8'b10100100;
													assign node5088 = (inp[6]) ? 8'b11110111 : node5089;
														assign node5089 = (inp[12]) ? 8'b11110101 : 8'b10100101;
										assign node5093 = (inp[2]) ? node5111 : node5094;
											assign node5094 = (inp[6]) ? node5100 : node5095;
												assign node5095 = (inp[12]) ? node5097 : 8'b10101101;
													assign node5097 = (inp[0]) ? 8'b11111101 : 8'b00011010;
												assign node5100 = (inp[12]) ? node5106 : node5101;
													assign node5101 = (inp[0]) ? 8'b10110100 : node5102;
														assign node5102 = (inp[3]) ? 8'b10110100 : 8'b11110111;
													assign node5106 = (inp[3]) ? 8'b10100101 : node5107;
														assign node5107 = (inp[0]) ? 8'b10100101 : 8'b00000010;
											assign node5111 = (inp[0]) ? node5125 : node5112;
												assign node5112 = (inp[3]) ? node5118 : node5113;
													assign node5113 = (inp[6]) ? 8'b11110101 : node5114;
														assign node5114 = (inp[12]) ? 8'b00000010 : 8'b11110111;
													assign node5118 = (inp[6]) ? node5122 : node5119;
														assign node5119 = (inp[12]) ? 8'b10100101 : 8'b10110100;
														assign node5122 = (inp[12]) ? 8'b10110100 : 8'b10100100;
												assign node5125 = (inp[12]) ? 8'b10110100 : 8'b10100100;
						assign node5128 = (inp[5]) ? node5304 : node5129;
							assign node5129 = (inp[0]) ? node5179 : node5130;
								assign node5130 = (inp[12]) ? node5162 : node5131;
									assign node5131 = (inp[11]) ? node5149 : node5132;
										assign node5132 = (inp[6]) ? node5144 : node5133;
											assign node5133 = (inp[2]) ? node5139 : node5134;
												assign node5134 = (inp[1]) ? 8'b00011010 : node5135;
													assign node5135 = (inp[3]) ? 8'b00011010 : 8'b00011011;
												assign node5139 = (inp[3]) ? 8'b10000010 : node5140;
													assign node5140 = (inp[1]) ? 8'b10000010 : 8'b00001011;
											assign node5144 = (inp[3]) ? 8'b10000010 : node5145;
												assign node5145 = (inp[1]) ? 8'b10000010 : 8'b00001011;
										assign node5149 = (inp[2]) ? node5157 : node5150;
											assign node5150 = (inp[6]) ? 8'b11110111 : node5151;
												assign node5151 = (inp[1]) ? 8'b00001010 : node5152;
													assign node5152 = (inp[3]) ? 8'b00001010 : 8'b00001011;
											assign node5157 = (inp[1]) ? 8'b11110111 : node5158;
												assign node5158 = (inp[3]) ? 8'b11110111 : 8'b00011010;
									assign node5162 = (inp[3]) ? node5174 : node5163;
										assign node5163 = (inp[1]) ? node5169 : node5164;
											assign node5164 = (inp[2]) ? 8'b00001011 : node5165;
												assign node5165 = (inp[6]) ? 8'b00001011 : 8'b00011011;
											assign node5169 = (inp[6]) ? 8'b00000010 : node5170;
												assign node5170 = (inp[2]) ? 8'b00000010 : 8'b00011010;
										assign node5174 = (inp[2]) ? 8'b00000010 : node5175;
											assign node5175 = (inp[6]) ? 8'b00000010 : 8'b00011010;
								assign node5179 = (inp[10]) ? node5225 : node5180;
									assign node5180 = (inp[11]) ? node5194 : node5181;
										assign node5181 = (inp[6]) ? node5189 : node5182;
											assign node5182 = (inp[3]) ? node5186 : node5183;
												assign node5183 = (inp[1]) ? 8'b10010101 : 8'b10011101;
												assign node5186 = (inp[2]) ? 8'b10010100 : 8'b10011100;
											assign node5189 = (inp[3]) ? 8'b10000100 : node5190;
												assign node5190 = (inp[1]) ? 8'b10000101 : 8'b10001101;
										assign node5194 = (inp[1]) ? node5212 : node5195;
											assign node5195 = (inp[3]) ? node5203 : node5196;
												assign node5196 = (inp[12]) ? node5200 : node5197;
													assign node5197 = (inp[6]) ? 8'b10111100 : 8'b10101101;
													assign node5200 = (inp[6]) ? 8'b10101101 : 8'b11111101;
												assign node5203 = (inp[2]) ? node5207 : node5204;
													assign node5204 = (inp[6]) ? 8'b10110001 : 8'b10101100;
													assign node5207 = (inp[12]) ? node5209 : 8'b10110001;
														assign node5209 = (inp[6]) ? 8'b10100100 : 8'b10110001;
											assign node5212 = (inp[6]) ? node5222 : node5213;
												assign node5213 = (inp[12]) ? node5219 : node5214;
													assign node5214 = (inp[2]) ? node5216 : 8'b10101100;
														assign node5216 = (inp[3]) ? 8'b10100001 : 8'b10100000;
													assign node5219 = (inp[2]) ? 8'b10110001 : 8'b10111001;
												assign node5222 = (inp[3]) ? 8'b10110001 : 8'b10110000;
									assign node5225 = (inp[1]) ? node5265 : node5226;
										assign node5226 = (inp[3]) ? node5246 : node5227;
											assign node5227 = (inp[11]) ? node5231 : node5228;
												assign node5228 = (inp[6]) ? 8'b00001011 : 8'b00011011;
												assign node5231 = (inp[2]) ? node5239 : node5232;
													assign node5232 = (inp[6]) ? node5236 : node5233;
														assign node5233 = (inp[12]) ? 8'b00011011 : 8'b00001011;
														assign node5236 = (inp[12]) ? 8'b00001011 : 8'b00011010;
													assign node5239 = (inp[12]) ? node5243 : node5240;
														assign node5240 = (inp[6]) ? 8'b00011010 : 8'b00001010;
														assign node5243 = (inp[6]) ? 8'b00001011 : 8'b00011010;
											assign node5246 = (inp[2]) ? node5256 : node5247;
												assign node5247 = (inp[6]) ? node5251 : node5248;
													assign node5248 = (inp[12]) ? 8'b00011010 : 8'b00001010;
													assign node5251 = (inp[12]) ? 8'b00000010 : node5252;
														assign node5252 = (inp[11]) ? 8'b11110111 : 8'b10000010;
												assign node5256 = (inp[11]) ? node5260 : node5257;
													assign node5257 = (inp[12]) ? 8'b00000010 : 8'b10010000;
													assign node5260 = (inp[6]) ? 8'b11110111 : node5261;
														assign node5261 = (inp[12]) ? 8'b11110101 : 8'b10100101;
										assign node5265 = (inp[3]) ? node5279 : node5266;
											assign node5266 = (inp[11]) ? node5272 : node5267;
												assign node5267 = (inp[6]) ? 8'b10000001 : node5268;
													assign node5268 = (inp[2]) ? 8'b10010001 : 8'b10011001;
												assign node5272 = (inp[2]) ? node5276 : node5273;
													assign node5273 = (inp[6]) ? 8'b10100101 : 8'b11111101;
													assign node5276 = (inp[6]) ? 8'b10110100 : 8'b10100100;
											assign node5279 = (inp[2]) ? node5291 : node5280;
												assign node5280 = (inp[6]) ? node5286 : node5281;
													assign node5281 = (inp[11]) ? node5283 : 8'b00011010;
														assign node5283 = (inp[12]) ? 8'b00011010 : 8'b00001010;
													assign node5286 = (inp[12]) ? 8'b00000010 : node5287;
														assign node5287 = (inp[11]) ? 8'b11110111 : 8'b10000010;
												assign node5291 = (inp[11]) ? node5297 : node5292;
													assign node5292 = (inp[6]) ? node5294 : 8'b10010000;
														assign node5294 = (inp[12]) ? 8'b00000010 : 8'b10000010;
													assign node5297 = (inp[6]) ? node5301 : node5298;
														assign node5298 = (inp[12]) ? 8'b11110101 : 8'b10100101;
														assign node5301 = (inp[12]) ? 8'b00000010 : 8'b11110111;
							assign node5304 = (inp[11]) ? node5388 : node5305;
								assign node5305 = (inp[0]) ? node5373 : node5306;
									assign node5306 = (inp[10]) ? node5344 : node5307;
										assign node5307 = (inp[6]) ? node5325 : node5308;
											assign node5308 = (inp[2]) ? node5316 : node5309;
												assign node5309 = (inp[1]) ? node5313 : node5310;
													assign node5310 = (inp[3]) ? 8'b00011010 : 8'b00011011;
													assign node5313 = (inp[3]) ? 8'b10011001 : 8'b00011010;
												assign node5316 = (inp[12]) ? 8'b00000010 : node5317;
													assign node5317 = (inp[3]) ? node5321 : node5318;
														assign node5318 = (inp[1]) ? 8'b10000010 : 8'b00001011;
														assign node5321 = (inp[1]) ? 8'b10000001 : 8'b10000010;
											assign node5325 = (inp[2]) ? node5339 : node5326;
												assign node5326 = (inp[12]) ? node5332 : node5327;
													assign node5327 = (inp[3]) ? node5329 : 8'b10000010;
														assign node5329 = (inp[1]) ? 8'b10000001 : 8'b10000010;
													assign node5332 = (inp[3]) ? node5336 : node5333;
														assign node5333 = (inp[1]) ? 8'b00000010 : 8'b00001011;
														assign node5336 = (inp[1]) ? 8'b10000001 : 8'b00000010;
												assign node5339 = (inp[1]) ? node5341 : 8'b10010000;
													assign node5341 = (inp[3]) ? 8'b10010001 : 8'b10010000;
										assign node5344 = (inp[6]) ? node5358 : node5345;
											assign node5345 = (inp[2]) ? node5353 : node5346;
												assign node5346 = (inp[1]) ? node5350 : node5347;
													assign node5347 = (inp[3]) ? 8'b10011100 : 8'b10011101;
													assign node5350 = (inp[3]) ? 8'b10011101 : 8'b10011100;
												assign node5353 = (inp[1]) ? 8'b10000100 : node5354;
													assign node5354 = (inp[3]) ? 8'b10000100 : 8'b10001101;
											assign node5358 = (inp[2]) ? node5366 : node5359;
												assign node5359 = (inp[1]) ? node5363 : node5360;
													assign node5360 = (inp[3]) ? 8'b10000100 : 8'b10001101;
													assign node5363 = (inp[3]) ? 8'b10000101 : 8'b10000100;
												assign node5366 = (inp[1]) ? node5370 : node5367;
													assign node5367 = (inp[3]) ? 8'b10010100 : 8'b10011101;
													assign node5370 = (inp[3]) ? 8'b10010101 : 8'b10010100;
									assign node5373 = (inp[2]) ? node5383 : node5374;
										assign node5374 = (inp[6]) ? node5376 : 8'b10011101;
											assign node5376 = (inp[3]) ? node5380 : node5377;
												assign node5377 = (inp[1]) ? 8'b10000101 : 8'b10001101;
												assign node5380 = (inp[1]) ? 8'b10000101 : 8'b10000100;
										assign node5383 = (inp[1]) ? 8'b10010101 : node5384;
											assign node5384 = (inp[3]) ? 8'b10010100 : 8'b10011101;
								assign node5388 = (inp[1]) ? node5448 : node5389;
									assign node5389 = (inp[3]) ? node5413 : node5390;
										assign node5390 = (inp[0]) ? node5404 : node5391;
											assign node5391 = (inp[10]) ? node5397 : node5392;
												assign node5392 = (inp[12]) ? node5394 : 8'b00011010;
													assign node5394 = (inp[6]) ? 8'b00011010 : 8'b00001011;
												assign node5397 = (inp[12]) ? node5399 : 8'b10111100;
													assign node5399 = (inp[6]) ? 8'b10101101 : node5400;
														assign node5400 = (inp[2]) ? 8'b10101101 : 8'b11111101;
											assign node5404 = (inp[2]) ? node5410 : node5405;
												assign node5405 = (inp[6]) ? node5407 : 8'b11111101;
													assign node5407 = (inp[12]) ? 8'b10101101 : 8'b10111100;
												assign node5410 = (inp[12]) ? 8'b10111100 : 8'b10101100;
										assign node5413 = (inp[2]) ? node5431 : node5414;
											assign node5414 = (inp[6]) ? node5422 : node5415;
												assign node5415 = (inp[10]) ? node5419 : node5416;
													assign node5416 = (inp[0]) ? 8'b10111100 : 8'b00011010;
													assign node5419 = (inp[12]) ? 8'b10111100 : 8'b10101100;
												assign node5422 = (inp[12]) ? node5426 : node5423;
													assign node5423 = (inp[0]) ? 8'b10110001 : 8'b11110111;
													assign node5426 = (inp[10]) ? 8'b10100100 : node5427;
														assign node5427 = (inp[0]) ? 8'b10100100 : 8'b00000010;
											assign node5431 = (inp[0]) ? node5445 : node5432;
												assign node5432 = (inp[6]) ? node5438 : node5433;
													assign node5433 = (inp[10]) ? node5435 : 8'b00000010;
														assign node5435 = (inp[12]) ? 8'b10100100 : 8'b10110001;
													assign node5438 = (inp[12]) ? node5442 : node5439;
														assign node5439 = (inp[10]) ? 8'b10100001 : 8'b10100101;
														assign node5442 = (inp[10]) ? 8'b10110001 : 8'b11110101;
												assign node5445 = (inp[12]) ? 8'b10110001 : 8'b10100001;
									assign node5448 = (inp[0]) ? node5488 : node5449;
										assign node5449 = (inp[10]) ? node5465 : node5450;
											assign node5450 = (inp[3]) ? node5458 : node5451;
												assign node5451 = (inp[12]) ? node5453 : 8'b11110111;
													assign node5453 = (inp[6]) ? 8'b00000010 : node5454;
														assign node5454 = (inp[2]) ? 8'b00000010 : 8'b00011010;
												assign node5458 = (inp[2]) ? 8'b10110100 : node5459;
													assign node5459 = (inp[6]) ? 8'b10100101 : node5460;
														assign node5460 = (inp[12]) ? 8'b11111101 : 8'b10101101;
											assign node5465 = (inp[6]) ? node5477 : node5466;
												assign node5466 = (inp[3]) ? node5472 : node5467;
													assign node5467 = (inp[2]) ? 8'b10100100 : node5468;
														assign node5468 = (inp[12]) ? 8'b10111100 : 8'b10101100;
													assign node5472 = (inp[2]) ? node5474 : 8'b10111001;
														assign node5474 = (inp[12]) ? 8'b10100001 : 8'b10110000;
												assign node5477 = (inp[2]) ? node5485 : node5478;
													assign node5478 = (inp[12]) ? node5482 : node5479;
														assign node5479 = (inp[3]) ? 8'b10110000 : 8'b10110001;
														assign node5482 = (inp[3]) ? 8'b10100001 : 8'b10100100;
													assign node5485 = (inp[12]) ? 8'b10110001 : 8'b10100001;
										assign node5488 = (inp[2]) ? node5496 : node5489;
											assign node5489 = (inp[6]) ? node5493 : node5490;
												assign node5490 = (inp[12]) ? 8'b10111001 : 8'b10101001;
												assign node5493 = (inp[12]) ? 8'b10100001 : 8'b10110000;
											assign node5496 = (inp[12]) ? 8'b10110000 : 8'b10100000;
				assign node5499 = (inp[0]) ? node6285 : node5500;
					assign node5500 = (inp[5]) ? node5664 : node5501;
						assign node5501 = (inp[12]) ? node5611 : node5502;
							assign node5502 = (inp[11]) ? node5558 : node5503;
								assign node5503 = (inp[2]) ? node5541 : node5504;
									assign node5504 = (inp[6]) ? node5522 : node5505;
										assign node5505 = (inp[8]) ? node5517 : node5506;
											assign node5506 = (inp[10]) ? node5512 : node5507;
												assign node5507 = (inp[1]) ? 8'b00011110 : node5508;
													assign node5508 = (inp[3]) ? 8'b00011110 : 8'b00011111;
												assign node5512 = (inp[1]) ? 8'b00011010 : node5513;
													assign node5513 = (inp[3]) ? 8'b00011010 : 8'b00011011;
											assign node5517 = (inp[3]) ? 8'b00011010 : node5518;
												assign node5518 = (inp[1]) ? 8'b00011010 : 8'b00011011;
										assign node5522 = (inp[3]) ? node5536 : node5523;
											assign node5523 = (inp[1]) ? node5529 : node5524;
												assign node5524 = (inp[10]) ? 8'b00001011 : node5525;
													assign node5525 = (inp[8]) ? 8'b00001011 : 8'b00001111;
												assign node5529 = (inp[9]) ? node5531 : 8'b00001110;
													assign node5531 = (inp[8]) ? 8'b10000010 : node5532;
														assign node5532 = (inp[10]) ? 8'b10000010 : 8'b00001110;
											assign node5536 = (inp[10]) ? 8'b10000010 : node5537;
												assign node5537 = (inp[8]) ? 8'b10000010 : 8'b00001110;
									assign node5541 = (inp[8]) ? node5553 : node5542;
										assign node5542 = (inp[10]) ? node5548 : node5543;
											assign node5543 = (inp[1]) ? 8'b00001110 : node5544;
												assign node5544 = (inp[3]) ? 8'b00001110 : 8'b00001111;
											assign node5548 = (inp[3]) ? 8'b10000010 : node5549;
												assign node5549 = (inp[1]) ? 8'b10000010 : 8'b00001011;
										assign node5553 = (inp[1]) ? 8'b10000010 : node5554;
											assign node5554 = (inp[3]) ? 8'b10000010 : 8'b00001011;
								assign node5558 = (inp[6]) ? node5594 : node5559;
									assign node5559 = (inp[2]) ? node5577 : node5560;
										assign node5560 = (inp[10]) ? node5572 : node5561;
											assign node5561 = (inp[8]) ? node5567 : node5562;
												assign node5562 = (inp[3]) ? 8'b00001110 : node5563;
													assign node5563 = (inp[1]) ? 8'b00001110 : 8'b00001111;
												assign node5567 = (inp[1]) ? 8'b00001010 : node5568;
													assign node5568 = (inp[3]) ? 8'b00001010 : 8'b00001011;
											assign node5572 = (inp[1]) ? 8'b00001010 : node5573;
												assign node5573 = (inp[3]) ? 8'b00001010 : 8'b00001011;
										assign node5577 = (inp[1]) ? node5589 : node5578;
											assign node5578 = (inp[3]) ? node5584 : node5579;
												assign node5579 = (inp[8]) ? 8'b00011010 : node5580;
													assign node5580 = (inp[10]) ? 8'b00011010 : 8'b00011110;
												assign node5584 = (inp[8]) ? 8'b11110111 : node5585;
													assign node5585 = (inp[10]) ? 8'b11110111 : 8'b00011011;
											assign node5589 = (inp[10]) ? 8'b11110111 : node5590;
												assign node5590 = (inp[8]) ? 8'b11110111 : 8'b00011011;
									assign node5594 = (inp[1]) ? node5606 : node5595;
										assign node5595 = (inp[3]) ? node5601 : node5596;
											assign node5596 = (inp[10]) ? 8'b00011010 : node5597;
												assign node5597 = (inp[8]) ? 8'b00011010 : 8'b00011110;
											assign node5601 = (inp[10]) ? 8'b11110111 : node5602;
												assign node5602 = (inp[8]) ? 8'b11110111 : 8'b00011011;
										assign node5606 = (inp[8]) ? 8'b11110111 : node5607;
											assign node5607 = (inp[10]) ? 8'b11110111 : 8'b00011011;
							assign node5611 = (inp[1]) ? node5647 : node5612;
								assign node5612 = (inp[3]) ? node5630 : node5613;
									assign node5613 = (inp[6]) ? node5625 : node5614;
										assign node5614 = (inp[2]) ? node5620 : node5615;
											assign node5615 = (inp[8]) ? 8'b00011011 : node5616;
												assign node5616 = (inp[10]) ? 8'b00011011 : 8'b00011111;
											assign node5620 = (inp[10]) ? 8'b00001011 : node5621;
												assign node5621 = (inp[8]) ? 8'b00001011 : 8'b00001111;
										assign node5625 = (inp[10]) ? 8'b00001011 : node5626;
											assign node5626 = (inp[8]) ? 8'b00001011 : 8'b00001111;
									assign node5630 = (inp[8]) ? node5642 : node5631;
										assign node5631 = (inp[10]) ? node5637 : node5632;
											assign node5632 = (inp[6]) ? 8'b00001110 : node5633;
												assign node5633 = (inp[2]) ? 8'b00001110 : 8'b00011110;
											assign node5637 = (inp[6]) ? 8'b00000010 : node5638;
												assign node5638 = (inp[2]) ? 8'b00000010 : 8'b00011010;
										assign node5642 = (inp[6]) ? 8'b00000010 : node5643;
											assign node5643 = (inp[2]) ? 8'b00000010 : 8'b00011010;
								assign node5647 = (inp[8]) ? node5659 : node5648;
									assign node5648 = (inp[10]) ? node5654 : node5649;
										assign node5649 = (inp[2]) ? 8'b00001110 : node5650;
											assign node5650 = (inp[6]) ? 8'b00001110 : 8'b00011110;
										assign node5654 = (inp[6]) ? 8'b00000010 : node5655;
											assign node5655 = (inp[2]) ? 8'b00000010 : 8'b00011010;
									assign node5659 = (inp[2]) ? 8'b00000010 : node5660;
										assign node5660 = (inp[6]) ? 8'b00000010 : 8'b00011010;
						assign node5664 = (inp[9]) ? node5984 : node5665;
							assign node5665 = (inp[8]) ? node5829 : node5666;
								assign node5666 = (inp[10]) ? node5750 : node5667;
									assign node5667 = (inp[11]) ? node5705 : node5668;
										assign node5668 = (inp[12]) ? node5692 : node5669;
											assign node5669 = (inp[6]) ? node5683 : node5670;
												assign node5670 = (inp[2]) ? node5676 : node5671;
													assign node5671 = (inp[3]) ? 8'b00011110 : node5672;
														assign node5672 = (inp[1]) ? 8'b00011110 : 8'b00011111;
													assign node5676 = (inp[3]) ? node5680 : node5677;
														assign node5677 = (inp[1]) ? 8'b00001110 : 8'b00001111;
														assign node5680 = (inp[1]) ? 8'b00001111 : 8'b00001110;
												assign node5683 = (inp[2]) ? node5685 : 8'b00001110;
													assign node5685 = (inp[1]) ? node5689 : node5686;
														assign node5686 = (inp[3]) ? 8'b00011110 : 8'b00011111;
														assign node5689 = (inp[3]) ? 8'b00011111 : 8'b00011110;
											assign node5692 = (inp[1]) ? node5702 : node5693;
												assign node5693 = (inp[3]) ? node5697 : node5694;
													assign node5694 = (inp[6]) ? 8'b00001111 : 8'b00011111;
													assign node5697 = (inp[2]) ? 8'b00001110 : node5698;
														assign node5698 = (inp[6]) ? 8'b00001110 : 8'b00011110;
												assign node5702 = (inp[3]) ? 8'b00001111 : 8'b00001110;
										assign node5705 = (inp[3]) ? node5733 : node5706;
											assign node5706 = (inp[1]) ? node5720 : node5707;
												assign node5707 = (inp[2]) ? node5713 : node5708;
													assign node5708 = (inp[6]) ? 8'b00001111 : node5709;
														assign node5709 = (inp[12]) ? 8'b00011111 : 8'b00001111;
													assign node5713 = (inp[6]) ? node5717 : node5714;
														assign node5714 = (inp[12]) ? 8'b00001111 : 8'b00011110;
														assign node5717 = (inp[12]) ? 8'b00011110 : 8'b00001110;
												assign node5720 = (inp[6]) ? node5728 : node5721;
													assign node5721 = (inp[12]) ? node5725 : node5722;
														assign node5722 = (inp[2]) ? 8'b00011011 : 8'b00001110;
														assign node5725 = (inp[2]) ? 8'b00001110 : 8'b00011110;
													assign node5728 = (inp[12]) ? node5730 : 8'b00011011;
														assign node5730 = (inp[2]) ? 8'b00011011 : 8'b00001110;
											assign node5733 = (inp[1]) ? node5743 : node5734;
												assign node5734 = (inp[12]) ? 8'b00001110 : node5735;
													assign node5735 = (inp[2]) ? node5739 : node5736;
														assign node5736 = (inp[6]) ? 8'b00011011 : 8'b00001110;
														assign node5739 = (inp[6]) ? 8'b00001011 : 8'b00011011;
												assign node5743 = (inp[2]) ? node5747 : node5744;
													assign node5744 = (inp[6]) ? 8'b00001011 : 8'b00011011;
													assign node5747 = (inp[12]) ? 8'b00011010 : 8'b00001010;
									assign node5750 = (inp[1]) ? node5790 : node5751;
										assign node5751 = (inp[3]) ? node5771 : node5752;
											assign node5752 = (inp[6]) ? node5760 : node5753;
												assign node5753 = (inp[2]) ? 8'b00001011 : node5754;
													assign node5754 = (inp[11]) ? node5756 : 8'b00011011;
														assign node5756 = (inp[12]) ? 8'b00011011 : 8'b00001011;
												assign node5760 = (inp[11]) ? node5764 : node5761;
													assign node5761 = (inp[2]) ? 8'b00011011 : 8'b00001011;
													assign node5764 = (inp[12]) ? node5768 : node5765;
														assign node5765 = (inp[2]) ? 8'b00001010 : 8'b00011010;
														assign node5768 = (inp[2]) ? 8'b00011010 : 8'b00001011;
											assign node5771 = (inp[2]) ? node5781 : node5772;
												assign node5772 = (inp[6]) ? node5778 : node5773;
													assign node5773 = (inp[11]) ? node5775 : 8'b00011010;
														assign node5775 = (inp[12]) ? 8'b00011010 : 8'b00001010;
													assign node5778 = (inp[12]) ? 8'b00000010 : 8'b10000010;
												assign node5781 = (inp[6]) ? node5787 : node5782;
													assign node5782 = (inp[12]) ? 8'b00000010 : node5783;
														assign node5783 = (inp[11]) ? 8'b11110111 : 8'b10000010;
													assign node5787 = (inp[11]) ? 8'b11110101 : 8'b10010000;
										assign node5790 = (inp[11]) ? node5808 : node5791;
											assign node5791 = (inp[3]) ? node5801 : node5792;
												assign node5792 = (inp[2]) ? node5796 : node5793;
													assign node5793 = (inp[6]) ? 8'b00000010 : 8'b00011010;
													assign node5796 = (inp[6]) ? 8'b10010000 : node5797;
														assign node5797 = (inp[12]) ? 8'b00000010 : 8'b10000010;
												assign node5801 = (inp[2]) ? node5805 : node5802;
													assign node5802 = (inp[6]) ? 8'b10000001 : 8'b10011001;
													assign node5805 = (inp[6]) ? 8'b10010001 : 8'b10000001;
											assign node5808 = (inp[3]) ? node5820 : node5809;
												assign node5809 = (inp[2]) ? node5817 : node5810;
													assign node5810 = (inp[6]) ? node5814 : node5811;
														assign node5811 = (inp[12]) ? 8'b00011010 : 8'b00001010;
														assign node5814 = (inp[12]) ? 8'b00000010 : 8'b11110111;
													assign node5817 = (inp[12]) ? 8'b11110101 : 8'b11110111;
												assign node5820 = (inp[6]) ? 8'b10110100 : node5821;
													assign node5821 = (inp[2]) ? node5825 : node5822;
														assign node5822 = (inp[12]) ? 8'b11111101 : 8'b10101101;
														assign node5825 = (inp[12]) ? 8'b10100101 : 8'b10110100;
								assign node5829 = (inp[10]) ? node5909 : node5830;
									assign node5830 = (inp[1]) ? node5874 : node5831;
										assign node5831 = (inp[3]) ? node5853 : node5832;
											assign node5832 = (inp[11]) ? node5840 : node5833;
												assign node5833 = (inp[12]) ? node5835 : 8'b00011011;
													assign node5835 = (inp[2]) ? node5837 : 8'b00001011;
														assign node5837 = (inp[6]) ? 8'b00011011 : 8'b00001011;
												assign node5840 = (inp[6]) ? node5848 : node5841;
													assign node5841 = (inp[12]) ? node5845 : node5842;
														assign node5842 = (inp[2]) ? 8'b00011010 : 8'b00001011;
														assign node5845 = (inp[2]) ? 8'b00001011 : 8'b00011011;
													assign node5848 = (inp[2]) ? node5850 : 8'b00011010;
														assign node5850 = (inp[12]) ? 8'b00011010 : 8'b00001010;
											assign node5853 = (inp[11]) ? node5863 : node5854;
												assign node5854 = (inp[6]) ? node5860 : node5855;
													assign node5855 = (inp[2]) ? node5857 : 8'b00011010;
														assign node5857 = (inp[12]) ? 8'b00000010 : 8'b10000010;
													assign node5860 = (inp[2]) ? 8'b10010000 : 8'b10000010;
												assign node5863 = (inp[12]) ? node5869 : node5864;
													assign node5864 = (inp[6]) ? 8'b11110111 : node5865;
														assign node5865 = (inp[2]) ? 8'b11110111 : 8'b00001010;
													assign node5869 = (inp[6]) ? node5871 : 8'b00000010;
														assign node5871 = (inp[2]) ? 8'b11110101 : 8'b00000010;
										assign node5874 = (inp[3]) ? node5892 : node5875;
											assign node5875 = (inp[2]) ? node5881 : node5876;
												assign node5876 = (inp[6]) ? node5878 : 8'b00001010;
													assign node5878 = (inp[12]) ? 8'b00000010 : 8'b10000010;
												assign node5881 = (inp[11]) ? node5887 : node5882;
													assign node5882 = (inp[6]) ? 8'b10010000 : node5883;
														assign node5883 = (inp[12]) ? 8'b00000010 : 8'b10000010;
													assign node5887 = (inp[6]) ? 8'b11110101 : node5888;
														assign node5888 = (inp[12]) ? 8'b00000010 : 8'b11110111;
											assign node5892 = (inp[11]) ? node5900 : node5893;
												assign node5893 = (inp[2]) ? node5897 : node5894;
													assign node5894 = (inp[6]) ? 8'b10000001 : 8'b10011001;
													assign node5897 = (inp[6]) ? 8'b10010001 : 8'b10000001;
												assign node5900 = (inp[2]) ? node5902 : 8'b11111101;
													assign node5902 = (inp[6]) ? node5906 : node5903;
														assign node5903 = (inp[12]) ? 8'b10100101 : 8'b10110100;
														assign node5906 = (inp[12]) ? 8'b10110100 : 8'b10100100;
									assign node5909 = (inp[11]) ? node5939 : node5910;
										assign node5910 = (inp[1]) ? node5924 : node5911;
											assign node5911 = (inp[3]) ? node5919 : node5912;
												assign node5912 = (inp[6]) ? node5916 : node5913;
													assign node5913 = (inp[2]) ? 8'b10001101 : 8'b10011101;
													assign node5916 = (inp[2]) ? 8'b10011101 : 8'b10001101;
												assign node5919 = (inp[6]) ? node5921 : 8'b10011100;
													assign node5921 = (inp[2]) ? 8'b10010100 : 8'b10000100;
											assign node5924 = (inp[3]) ? node5932 : node5925;
												assign node5925 = (inp[2]) ? node5929 : node5926;
													assign node5926 = (inp[6]) ? 8'b10000100 : 8'b10011100;
													assign node5929 = (inp[6]) ? 8'b10010100 : 8'b10000100;
												assign node5932 = (inp[6]) ? node5936 : node5933;
													assign node5933 = (inp[2]) ? 8'b10000101 : 8'b10011101;
													assign node5936 = (inp[2]) ? 8'b10010101 : 8'b10000101;
										assign node5939 = (inp[1]) ? node5963 : node5940;
											assign node5940 = (inp[3]) ? node5954 : node5941;
												assign node5941 = (inp[2]) ? node5947 : node5942;
													assign node5942 = (inp[6]) ? node5944 : 8'b10101101;
														assign node5944 = (inp[12]) ? 8'b10101101 : 8'b10111100;
													assign node5947 = (inp[12]) ? node5951 : node5948;
														assign node5948 = (inp[6]) ? 8'b10101100 : 8'b10111100;
														assign node5951 = (inp[6]) ? 8'b10111100 : 8'b10101101;
												assign node5954 = (inp[6]) ? 8'b10110001 : node5955;
													assign node5955 = (inp[2]) ? node5959 : node5956;
														assign node5956 = (inp[12]) ? 8'b10111100 : 8'b10101100;
														assign node5959 = (inp[12]) ? 8'b10100100 : 8'b10110001;
											assign node5963 = (inp[2]) ? node5975 : node5964;
												assign node5964 = (inp[6]) ? node5970 : node5965;
													assign node5965 = (inp[3]) ? node5967 : 8'b10111100;
														assign node5967 = (inp[12]) ? 8'b10111001 : 8'b10101001;
													assign node5970 = (inp[12]) ? 8'b10100100 : node5971;
														assign node5971 = (inp[3]) ? 8'b10110000 : 8'b10110001;
												assign node5975 = (inp[3]) ? node5981 : node5976;
													assign node5976 = (inp[6]) ? node5978 : 8'b10110001;
														assign node5978 = (inp[12]) ? 8'b10110001 : 8'b10100001;
													assign node5981 = (inp[6]) ? 8'b10110000 : 8'b10100001;
							assign node5984 = (inp[11]) ? node6106 : node5985;
								assign node5985 = (inp[2]) ? node6047 : node5986;
									assign node5986 = (inp[6]) ? node6018 : node5987;
										assign node5987 = (inp[3]) ? node6003 : node5988;
											assign node5988 = (inp[1]) ? node5996 : node5989;
												assign node5989 = (inp[10]) ? node5993 : node5990;
													assign node5990 = (inp[8]) ? 8'b10111001 : 8'b11111101;
													assign node5993 = (inp[8]) ? 8'b11111101 : 8'b10111001;
												assign node5996 = (inp[10]) ? node6000 : node5997;
													assign node5997 = (inp[8]) ? 8'b10111000 : 8'b10111100;
													assign node6000 = (inp[8]) ? 8'b10111100 : 8'b10111000;
											assign node6003 = (inp[1]) ? node6011 : node6004;
												assign node6004 = (inp[8]) ? node6008 : node6005;
													assign node6005 = (inp[10]) ? 8'b10111000 : 8'b10111100;
													assign node6008 = (inp[10]) ? 8'b10111100 : 8'b10111000;
												assign node6011 = (inp[8]) ? node6015 : node6012;
													assign node6012 = (inp[10]) ? 8'b10111001 : 8'b11111101;
													assign node6015 = (inp[10]) ? 8'b11111101 : 8'b10111001;
										assign node6018 = (inp[10]) ? node6032 : node6019;
											assign node6019 = (inp[8]) ? node6029 : node6020;
												assign node6020 = (inp[12]) ? node6022 : 8'b10101100;
													assign node6022 = (inp[3]) ? node6026 : node6023;
														assign node6023 = (inp[1]) ? 8'b10101100 : 8'b10101101;
														assign node6026 = (inp[1]) ? 8'b10101101 : 8'b10101100;
												assign node6029 = (inp[3]) ? 8'b10100000 : 8'b10101001;
											assign node6032 = (inp[8]) ? node6040 : node6033;
												assign node6033 = (inp[3]) ? node6037 : node6034;
													assign node6034 = (inp[1]) ? 8'b10100000 : 8'b10101001;
													assign node6037 = (inp[1]) ? 8'b10100001 : 8'b10100000;
												assign node6040 = (inp[3]) ? node6044 : node6041;
													assign node6041 = (inp[1]) ? 8'b10100100 : 8'b10101101;
													assign node6044 = (inp[1]) ? 8'b10100101 : 8'b10100100;
									assign node6047 = (inp[6]) ? node6073 : node6048;
										assign node6048 = (inp[3]) ? node6064 : node6049;
											assign node6049 = (inp[1]) ? node6057 : node6050;
												assign node6050 = (inp[8]) ? node6054 : node6051;
													assign node6051 = (inp[10]) ? 8'b10101001 : 8'b10101101;
													assign node6054 = (inp[10]) ? 8'b10101101 : 8'b10101001;
												assign node6057 = (inp[10]) ? node6061 : node6058;
													assign node6058 = (inp[8]) ? 8'b10100000 : 8'b10101100;
													assign node6061 = (inp[8]) ? 8'b10100100 : 8'b10100000;
											assign node6064 = (inp[1]) ? node6066 : 8'b10100000;
												assign node6066 = (inp[8]) ? node6070 : node6067;
													assign node6067 = (inp[10]) ? 8'b10100001 : 8'b10101101;
													assign node6070 = (inp[10]) ? 8'b10100101 : 8'b10100001;
										assign node6073 = (inp[1]) ? node6091 : node6074;
											assign node6074 = (inp[3]) ? node6082 : node6075;
												assign node6075 = (inp[10]) ? node6079 : node6076;
													assign node6076 = (inp[8]) ? 8'b10111001 : 8'b11111101;
													assign node6079 = (inp[8]) ? 8'b11111101 : 8'b10111001;
												assign node6082 = (inp[12]) ? node6084 : 8'b10110000;
													assign node6084 = (inp[8]) ? node6088 : node6085;
														assign node6085 = (inp[10]) ? 8'b10110000 : 8'b10111100;
														assign node6088 = (inp[10]) ? 8'b10110100 : 8'b10110000;
											assign node6091 = (inp[3]) ? node6099 : node6092;
												assign node6092 = (inp[8]) ? node6096 : node6093;
													assign node6093 = (inp[10]) ? 8'b10110000 : 8'b10111100;
													assign node6096 = (inp[10]) ? 8'b10110100 : 8'b10110000;
												assign node6099 = (inp[10]) ? node6103 : node6100;
													assign node6100 = (inp[8]) ? 8'b10110001 : 8'b11111101;
													assign node6103 = (inp[8]) ? 8'b11110101 : 8'b10110001;
								assign node6106 = (inp[8]) ? node6194 : node6107;
									assign node6107 = (inp[10]) ? node6153 : node6108;
										assign node6108 = (inp[1]) ? node6132 : node6109;
											assign node6109 = (inp[3]) ? node6119 : node6110;
												assign node6110 = (inp[2]) ? node6114 : node6111;
													assign node6111 = (inp[12]) ? 8'b11111101 : 8'b10101101;
													assign node6114 = (inp[6]) ? node6116 : 8'b10111100;
														assign node6116 = (inp[12]) ? 8'b10111100 : 8'b10101100;
												assign node6119 = (inp[6]) ? node6125 : node6120;
													assign node6120 = (inp[2]) ? node6122 : 8'b10101100;
														assign node6122 = (inp[12]) ? 8'b10101100 : 8'b10111001;
													assign node6125 = (inp[2]) ? node6129 : node6126;
														assign node6126 = (inp[12]) ? 8'b10101100 : 8'b10111001;
														assign node6129 = (inp[12]) ? 8'b10111001 : 8'b10101001;
											assign node6132 = (inp[3]) ? node6140 : node6133;
												assign node6133 = (inp[12]) ? node6135 : 8'b10111001;
													assign node6135 = (inp[2]) ? node6137 : 8'b10101100;
														assign node6137 = (inp[6]) ? 8'b10111001 : 8'b10101100;
												assign node6140 = (inp[6]) ? node6148 : node6141;
													assign node6141 = (inp[12]) ? node6145 : node6142;
														assign node6142 = (inp[2]) ? 8'b10111000 : 8'b10101001;
														assign node6145 = (inp[2]) ? 8'b10101001 : 8'b10111001;
													assign node6148 = (inp[12]) ? 8'b10111000 : node6149;
														assign node6149 = (inp[2]) ? 8'b10101000 : 8'b10111000;
										assign node6153 = (inp[1]) ? node6171 : node6154;
											assign node6154 = (inp[3]) ? node6166 : node6155;
												assign node6155 = (inp[6]) ? node6161 : node6156;
													assign node6156 = (inp[12]) ? node6158 : 8'b10101001;
														assign node6158 = (inp[2]) ? 8'b10101001 : 8'b10111001;
													assign node6161 = (inp[12]) ? node6163 : 8'b10111000;
														assign node6163 = (inp[2]) ? 8'b10111000 : 8'b10101001;
												assign node6166 = (inp[12]) ? node6168 : 8'b10010101;
													assign node6168 = (inp[6]) ? 8'b10100000 : 8'b10111000;
											assign node6171 = (inp[6]) ? node6183 : node6172;
												assign node6172 = (inp[12]) ? node6178 : node6173;
													assign node6173 = (inp[2]) ? node6175 : 8'b10001101;
														assign node6175 = (inp[3]) ? 8'b10010100 : 8'b10010101;
													assign node6178 = (inp[3]) ? 8'b10000101 : node6179;
														assign node6179 = (inp[2]) ? 8'b10100000 : 8'b10111000;
												assign node6183 = (inp[3]) ? node6189 : node6184;
													assign node6184 = (inp[2]) ? node6186 : 8'b10010101;
														assign node6186 = (inp[12]) ? 8'b10010101 : 8'b10000101;
													assign node6189 = (inp[2]) ? node6191 : 8'b10000101;
														assign node6191 = (inp[12]) ? 8'b10010100 : 8'b10000100;
									assign node6194 = (inp[2]) ? node6246 : node6195;
										assign node6195 = (inp[6]) ? node6219 : node6196;
											assign node6196 = (inp[12]) ? node6210 : node6197;
												assign node6197 = (inp[10]) ? node6203 : node6198;
													assign node6198 = (inp[3]) ? 8'b10001101 : node6199;
														assign node6199 = (inp[1]) ? 8'b10101000 : 8'b10101001;
													assign node6203 = (inp[1]) ? node6207 : node6204;
														assign node6204 = (inp[3]) ? 8'b10001100 : 8'b10001101;
														assign node6207 = (inp[3]) ? 8'b10001001 : 8'b10001100;
												assign node6210 = (inp[1]) ? node6214 : node6211;
													assign node6211 = (inp[3]) ? 8'b10011100 : 8'b10011101;
													assign node6214 = (inp[3]) ? node6216 : 8'b10111000;
														assign node6216 = (inp[10]) ? 8'b10011001 : 8'b10011101;
											assign node6219 = (inp[12]) ? node6233 : node6220;
												assign node6220 = (inp[1]) ? node6226 : node6221;
													assign node6221 = (inp[3]) ? 8'b10010101 : node6222;
														assign node6222 = (inp[10]) ? 8'b10011100 : 8'b10111000;
													assign node6226 = (inp[3]) ? node6230 : node6227;
														assign node6227 = (inp[10]) ? 8'b10010001 : 8'b10010101;
														assign node6230 = (inp[10]) ? 8'b10010000 : 8'b10010100;
												assign node6233 = (inp[10]) ? node6241 : node6234;
													assign node6234 = (inp[1]) ? node6238 : node6235;
														assign node6235 = (inp[3]) ? 8'b10100000 : 8'b10101001;
														assign node6238 = (inp[3]) ? 8'b10000101 : 8'b10100000;
													assign node6241 = (inp[1]) ? node6243 : 8'b10001101;
														assign node6243 = (inp[3]) ? 8'b10000001 : 8'b10000100;
										assign node6246 = (inp[10]) ? node6262 : node6247;
											assign node6247 = (inp[12]) ? node6255 : node6248;
												assign node6248 = (inp[6]) ? node6250 : 8'b10010101;
													assign node6250 = (inp[1]) ? node6252 : 8'b10000101;
														assign node6252 = (inp[3]) ? 8'b10000100 : 8'b10000101;
												assign node6255 = (inp[1]) ? node6259 : node6256;
													assign node6256 = (inp[3]) ? 8'b10100000 : 8'b10101001;
													assign node6259 = (inp[3]) ? 8'b10000101 : 8'b10100000;
											assign node6262 = (inp[3]) ? node6270 : node6263;
												assign node6263 = (inp[1]) ? node6267 : node6264;
													assign node6264 = (inp[12]) ? 8'b10001101 : 8'b10001100;
													assign node6267 = (inp[6]) ? 8'b10010001 : 8'b10000100;
												assign node6270 = (inp[1]) ? node6278 : node6271;
													assign node6271 = (inp[6]) ? node6275 : node6272;
														assign node6272 = (inp[12]) ? 8'b10000100 : 8'b10010001;
														assign node6275 = (inp[12]) ? 8'b10010001 : 8'b10000001;
													assign node6278 = (inp[12]) ? node6282 : node6279;
														assign node6279 = (inp[6]) ? 8'b10000000 : 8'b10010000;
														assign node6282 = (inp[6]) ? 8'b10010000 : 8'b10000001;
					assign node6285 = (inp[6]) ? node6611 : node6286;
						assign node6286 = (inp[11]) ? node6378 : node6287;
							assign node6287 = (inp[10]) ? node6335 : node6288;
								assign node6288 = (inp[3]) ? node6312 : node6289;
									assign node6289 = (inp[9]) ? node6297 : node6290;
										assign node6290 = (inp[8]) ? node6292 : 8'b11111101;
											assign node6292 = (inp[1]) ? node6294 : 8'b11111101;
												assign node6294 = (inp[2]) ? 8'b11110101 : 8'b11111101;
										assign node6297 = (inp[5]) ? node6305 : node6298;
											assign node6298 = (inp[8]) ? node6300 : 8'b00011111;
												assign node6300 = (inp[1]) ? node6302 : 8'b10011101;
													assign node6302 = (inp[2]) ? 8'b10010101 : 8'b10011101;
											assign node6305 = (inp[1]) ? node6307 : 8'b11111101;
												assign node6307 = (inp[2]) ? node6309 : 8'b11111101;
													assign node6309 = (inp[8]) ? 8'b11110101 : 8'b11111101;
									assign node6312 = (inp[5]) ? node6324 : node6313;
										assign node6313 = (inp[9]) ? node6319 : node6314;
											assign node6314 = (inp[8]) ? node6316 : 8'b10111100;
												assign node6316 = (inp[2]) ? 8'b10110100 : 8'b10111100;
											assign node6319 = (inp[8]) ? node6321 : 8'b00011110;
												assign node6321 = (inp[2]) ? 8'b10010100 : 8'b10011100;
										assign node6324 = (inp[1]) ? node6330 : node6325;
											assign node6325 = (inp[8]) ? node6327 : 8'b10111100;
												assign node6327 = (inp[2]) ? 8'b10110100 : 8'b10111100;
											assign node6330 = (inp[8]) ? node6332 : 8'b11111101;
												assign node6332 = (inp[2]) ? 8'b11110101 : 8'b11111101;
								assign node6335 = (inp[5]) ? node6357 : node6336;
									assign node6336 = (inp[9]) ? node6346 : node6337;
										assign node6337 = (inp[3]) ? node6343 : node6338;
											assign node6338 = (inp[2]) ? node6340 : 8'b10111001;
												assign node6340 = (inp[1]) ? 8'b10110001 : 8'b10111001;
											assign node6343 = (inp[2]) ? 8'b10110000 : 8'b10111000;
										assign node6346 = (inp[2]) ? node6352 : node6347;
											assign node6347 = (inp[3]) ? 8'b00011010 : node6348;
												assign node6348 = (inp[1]) ? 8'b10011001 : 8'b00011011;
											assign node6352 = (inp[3]) ? 8'b10010000 : node6353;
												assign node6353 = (inp[1]) ? 8'b10010001 : 8'b00011011;
									assign node6357 = (inp[8]) ? node6369 : node6358;
										assign node6358 = (inp[2]) ? node6364 : node6359;
											assign node6359 = (inp[1]) ? 8'b10111001 : node6360;
												assign node6360 = (inp[3]) ? 8'b10111000 : 8'b10111001;
											assign node6364 = (inp[1]) ? 8'b10110001 : node6365;
												assign node6365 = (inp[3]) ? 8'b10110000 : 8'b10111001;
										assign node6369 = (inp[1]) ? node6375 : node6370;
											assign node6370 = (inp[3]) ? node6372 : 8'b11111101;
												assign node6372 = (inp[2]) ? 8'b10110100 : 8'b10111100;
											assign node6375 = (inp[2]) ? 8'b11110101 : 8'b11111101;
							assign node6378 = (inp[12]) ? node6498 : node6379;
								assign node6379 = (inp[2]) ? node6445 : node6380;
									assign node6380 = (inp[3]) ? node6420 : node6381;
										assign node6381 = (inp[8]) ? node6401 : node6382;
											assign node6382 = (inp[9]) ? node6390 : node6383;
												assign node6383 = (inp[10]) ? node6387 : node6384;
													assign node6384 = (inp[1]) ? 8'b10101001 : 8'b10101101;
													assign node6387 = (inp[1]) ? 8'b10001101 : 8'b10101001;
												assign node6390 = (inp[5]) ? node6396 : node6391;
													assign node6391 = (inp[10]) ? node6393 : 8'b00001011;
														assign node6393 = (inp[1]) ? 8'b10101101 : 8'b00001011;
													assign node6396 = (inp[1]) ? 8'b10001101 : node6397;
														assign node6397 = (inp[10]) ? 8'b10101001 : 8'b10101101;
											assign node6401 = (inp[5]) ? node6417 : node6402;
												assign node6402 = (inp[9]) ? node6410 : node6403;
													assign node6403 = (inp[1]) ? node6407 : node6404;
														assign node6404 = (inp[10]) ? 8'b10101001 : 8'b10001101;
														assign node6407 = (inp[10]) ? 8'b10001101 : 8'b10001001;
													assign node6410 = (inp[1]) ? node6414 : node6411;
														assign node6411 = (inp[10]) ? 8'b00001011 : 8'b10101101;
														assign node6414 = (inp[10]) ? 8'b10101101 : 8'b10101001;
												assign node6417 = (inp[1]) ? 8'b10001001 : 8'b10001101;
										assign node6420 = (inp[10]) ? node6434 : node6421;
											assign node6421 = (inp[8]) ? node6429 : node6422;
												assign node6422 = (inp[5]) ? node6426 : node6423;
													assign node6423 = (inp[9]) ? 8'b00001110 : 8'b10101100;
													assign node6426 = (inp[1]) ? 8'b10101001 : 8'b10101100;
												assign node6429 = (inp[9]) ? node6431 : 8'b10001100;
													assign node6431 = (inp[5]) ? 8'b10001100 : 8'b10101100;
											assign node6434 = (inp[5]) ? node6438 : node6435;
												assign node6435 = (inp[9]) ? 8'b00001010 : 8'b10101000;
												assign node6438 = (inp[1]) ? node6442 : node6439;
													assign node6439 = (inp[8]) ? 8'b10001100 : 8'b10101000;
													assign node6442 = (inp[8]) ? 8'b10001001 : 8'b10001101;
									assign node6445 = (inp[3]) ? node6471 : node6446;
										assign node6446 = (inp[1]) ? node6460 : node6447;
											assign node6447 = (inp[8]) ? node6451 : node6448;
												assign node6448 = (inp[10]) ? 8'b10101000 : 8'b10101100;
												assign node6451 = (inp[5]) ? 8'b10001100 : node6452;
													assign node6452 = (inp[10]) ? node6456 : node6453;
														assign node6453 = (inp[9]) ? 8'b10101100 : 8'b10001100;
														assign node6456 = (inp[9]) ? 8'b00001010 : 8'b10101000;
											assign node6460 = (inp[10]) ? node6466 : node6461;
												assign node6461 = (inp[8]) ? 8'b10000000 : node6462;
													assign node6462 = (inp[9]) ? 8'b00001010 : 8'b10101000;
												assign node6466 = (inp[9]) ? node6468 : 8'b10000100;
													assign node6468 = (inp[5]) ? 8'b10000000 : 8'b10100100;
										assign node6471 = (inp[10]) ? node6487 : node6472;
											assign node6472 = (inp[8]) ? node6480 : node6473;
												assign node6473 = (inp[5]) ? node6477 : node6474;
													assign node6474 = (inp[9]) ? 8'b00001011 : 8'b10101001;
													assign node6477 = (inp[1]) ? 8'b10101000 : 8'b10101001;
												assign node6480 = (inp[5]) ? node6484 : node6481;
													assign node6481 = (inp[9]) ? 8'b10100001 : 8'b10000001;
													assign node6484 = (inp[1]) ? 8'b10000000 : 8'b10000001;
											assign node6487 = (inp[5]) ? node6491 : node6488;
												assign node6488 = (inp[9]) ? 8'b10100101 : 8'b10000101;
												assign node6491 = (inp[8]) ? node6495 : node6492;
													assign node6492 = (inp[1]) ? 8'b10000100 : 8'b10000101;
													assign node6495 = (inp[1]) ? 8'b10000000 : 8'b10000001;
								assign node6498 = (inp[2]) ? node6554 : node6499;
									assign node6499 = (inp[3]) ? node6533 : node6500;
										assign node6500 = (inp[9]) ? node6512 : node6501;
											assign node6501 = (inp[1]) ? node6507 : node6502;
												assign node6502 = (inp[10]) ? 8'b10111001 : node6503;
													assign node6503 = (inp[8]) ? 8'b10011101 : 8'b11111101;
												assign node6507 = (inp[10]) ? 8'b10011101 : node6508;
													assign node6508 = (inp[8]) ? 8'b10011001 : 8'b10111001;
											assign node6512 = (inp[5]) ? node6524 : node6513;
												assign node6513 = (inp[1]) ? node6519 : node6514;
													assign node6514 = (inp[10]) ? 8'b00011011 : node6515;
														assign node6515 = (inp[8]) ? 8'b11111101 : 8'b00011111;
													assign node6519 = (inp[10]) ? 8'b11111101 : node6520;
														assign node6520 = (inp[8]) ? 8'b10111001 : 8'b00011011;
												assign node6524 = (inp[1]) ? node6528 : node6525;
													assign node6525 = (inp[10]) ? 8'b10111001 : 8'b11111101;
													assign node6528 = (inp[8]) ? 8'b10011001 : node6529;
														assign node6529 = (inp[10]) ? 8'b10011101 : 8'b10111001;
										assign node6533 = (inp[5]) ? node6543 : node6534;
											assign node6534 = (inp[9]) ? node6538 : node6535;
												assign node6535 = (inp[10]) ? 8'b10111000 : 8'b10011100;
												assign node6538 = (inp[10]) ? 8'b00011010 : node6539;
													assign node6539 = (inp[8]) ? 8'b10111100 : 8'b00011110;
											assign node6543 = (inp[1]) ? node6549 : node6544;
												assign node6544 = (inp[10]) ? 8'b10111000 : node6545;
													assign node6545 = (inp[8]) ? 8'b10011100 : 8'b10111100;
												assign node6549 = (inp[10]) ? 8'b10011101 : node6550;
													assign node6550 = (inp[8]) ? 8'b10011001 : 8'b10111001;
									assign node6554 = (inp[3]) ? node6586 : node6555;
										assign node6555 = (inp[1]) ? node6573 : node6556;
											assign node6556 = (inp[10]) ? node6566 : node6557;
												assign node6557 = (inp[5]) ? 8'b10111100 : node6558;
													assign node6558 = (inp[8]) ? node6562 : node6559;
														assign node6559 = (inp[9]) ? 8'b00011110 : 8'b10111100;
														assign node6562 = (inp[9]) ? 8'b10111100 : 8'b10011100;
												assign node6566 = (inp[8]) ? node6568 : 8'b10111000;
													assign node6568 = (inp[9]) ? 8'b00011010 : node6569;
														assign node6569 = (inp[5]) ? 8'b10011100 : 8'b10111000;
											assign node6573 = (inp[10]) ? node6579 : node6574;
												assign node6574 = (inp[8]) ? 8'b10010000 : node6575;
													assign node6575 = (inp[5]) ? 8'b10111000 : 8'b00011010;
												assign node6579 = (inp[5]) ? node6583 : node6580;
													assign node6580 = (inp[9]) ? 8'b10110100 : 8'b10010100;
													assign node6583 = (inp[8]) ? 8'b10010000 : 8'b10010100;
										assign node6586 = (inp[10]) ? node6602 : node6587;
											assign node6587 = (inp[8]) ? node6595 : node6588;
												assign node6588 = (inp[9]) ? 8'b00011011 : node6589;
													assign node6589 = (inp[5]) ? node6591 : 8'b10111001;
														assign node6591 = (inp[1]) ? 8'b10111000 : 8'b10111001;
												assign node6595 = (inp[5]) ? node6599 : node6596;
													assign node6596 = (inp[1]) ? 8'b10010001 : 8'b10110001;
													assign node6599 = (inp[1]) ? 8'b10010000 : 8'b10010001;
											assign node6602 = (inp[9]) ? node6606 : node6603;
												assign node6603 = (inp[5]) ? 8'b10010100 : 8'b10010101;
												assign node6606 = (inp[5]) ? node6608 : 8'b11110101;
													assign node6608 = (inp[1]) ? 8'b10010100 : 8'b10010001;
						assign node6611 = (inp[5]) ? node6739 : node6612;
							assign node6612 = (inp[9]) ? node6666 : node6613;
								assign node6613 = (inp[3]) ? node6649 : node6614;
									assign node6614 = (inp[1]) ? node6632 : node6615;
										assign node6615 = (inp[10]) ? node6627 : node6616;
											assign node6616 = (inp[8]) ? node6622 : node6617;
												assign node6617 = (inp[11]) ? node6619 : 8'b10101101;
													assign node6619 = (inp[12]) ? 8'b10101101 : 8'b10111100;
												assign node6622 = (inp[12]) ? node6624 : 8'b10011100;
													assign node6624 = (inp[11]) ? 8'b10001101 : 8'b10101101;
											assign node6627 = (inp[11]) ? node6629 : 8'b10101001;
												assign node6629 = (inp[12]) ? 8'b10101001 : 8'b10111000;
										assign node6632 = (inp[11]) ? node6638 : node6633;
											assign node6633 = (inp[10]) ? 8'b10100001 : node6634;
												assign node6634 = (inp[8]) ? 8'b10100101 : 8'b10101101;
											assign node6638 = (inp[12]) ? node6644 : node6639;
												assign node6639 = (inp[10]) ? 8'b10010100 : node6640;
													assign node6640 = (inp[8]) ? 8'b10010000 : 8'b10111000;
												assign node6644 = (inp[10]) ? 8'b10000101 : node6645;
													assign node6645 = (inp[8]) ? 8'b10000001 : 8'b10101001;
									assign node6649 = (inp[11]) ? node6655 : node6650;
										assign node6650 = (inp[10]) ? 8'b10100000 : node6651;
											assign node6651 = (inp[8]) ? 8'b10100100 : 8'b10101100;
										assign node6655 = (inp[12]) ? node6661 : node6656;
											assign node6656 = (inp[10]) ? 8'b10010101 : node6657;
												assign node6657 = (inp[8]) ? 8'b10010001 : 8'b10111001;
											assign node6661 = (inp[10]) ? 8'b10100000 : node6662;
												assign node6662 = (inp[8]) ? 8'b10000100 : 8'b10101100;
								assign node6666 = (inp[8]) ? node6708 : node6667;
									assign node6667 = (inp[10]) ? node6683 : node6668;
										assign node6668 = (inp[11]) ? node6672 : node6669;
											assign node6669 = (inp[3]) ? 8'b00001110 : 8'b00001111;
											assign node6672 = (inp[12]) ? node6678 : node6673;
												assign node6673 = (inp[3]) ? 8'b00011011 : node6674;
													assign node6674 = (inp[1]) ? 8'b00011010 : 8'b00011110;
												assign node6678 = (inp[3]) ? 8'b00001110 : node6679;
													assign node6679 = (inp[1]) ? 8'b00001011 : 8'b00001111;
										assign node6683 = (inp[1]) ? node6695 : node6684;
											assign node6684 = (inp[3]) ? node6690 : node6685;
												assign node6685 = (inp[11]) ? node6687 : 8'b00001011;
													assign node6687 = (inp[12]) ? 8'b00001011 : 8'b00011010;
												assign node6690 = (inp[12]) ? 8'b00000010 : node6691;
													assign node6691 = (inp[11]) ? 8'b11110111 : 8'b10000010;
											assign node6695 = (inp[11]) ? node6701 : node6696;
												assign node6696 = (inp[3]) ? node6698 : 8'b10000001;
													assign node6698 = (inp[12]) ? 8'b00000010 : 8'b10000010;
												assign node6701 = (inp[3]) ? node6705 : node6702;
													assign node6702 = (inp[12]) ? 8'b10100101 : 8'b10110100;
													assign node6705 = (inp[12]) ? 8'b00000010 : 8'b11110111;
									assign node6708 = (inp[10]) ? node6726 : node6709;
										assign node6709 = (inp[11]) ? node6715 : node6710;
											assign node6710 = (inp[3]) ? 8'b10000100 : node6711;
												assign node6711 = (inp[1]) ? 8'b10000101 : 8'b10001101;
											assign node6715 = (inp[12]) ? node6721 : node6716;
												assign node6716 = (inp[3]) ? 8'b10110001 : node6717;
													assign node6717 = (inp[1]) ? 8'b10110000 : 8'b10111100;
												assign node6721 = (inp[3]) ? 8'b10100100 : node6722;
													assign node6722 = (inp[1]) ? 8'b10100001 : 8'b10101101;
										assign node6726 = (inp[3]) ? node6736 : node6727;
											assign node6727 = (inp[1]) ? node6731 : node6728;
												assign node6728 = (inp[11]) ? 8'b00011010 : 8'b00001011;
												assign node6731 = (inp[11]) ? node6733 : 8'b10000001;
													assign node6733 = (inp[12]) ? 8'b10100101 : 8'b10110100;
											assign node6736 = (inp[12]) ? 8'b00000010 : 8'b10000010;
							assign node6739 = (inp[11]) ? node6779 : node6740;
								assign node6740 = (inp[2]) ? node6760 : node6741;
									assign node6741 = (inp[8]) ? node6755 : node6742;
										assign node6742 = (inp[10]) ? node6748 : node6743;
											assign node6743 = (inp[1]) ? 8'b10101101 : node6744;
												assign node6744 = (inp[3]) ? 8'b10101100 : 8'b10101101;
											assign node6748 = (inp[3]) ? node6752 : node6749;
												assign node6749 = (inp[1]) ? 8'b10100001 : 8'b10101001;
												assign node6752 = (inp[1]) ? 8'b10100001 : 8'b10100000;
										assign node6755 = (inp[1]) ? 8'b10100101 : node6756;
											assign node6756 = (inp[3]) ? 8'b10100100 : 8'b10101101;
									assign node6760 = (inp[1]) ? node6774 : node6761;
										assign node6761 = (inp[3]) ? node6767 : node6762;
											assign node6762 = (inp[8]) ? 8'b11111101 : node6763;
												assign node6763 = (inp[10]) ? 8'b10111001 : 8'b11111101;
											assign node6767 = (inp[10]) ? node6771 : node6768;
												assign node6768 = (inp[8]) ? 8'b10110100 : 8'b10111100;
												assign node6771 = (inp[8]) ? 8'b10110100 : 8'b10110000;
										assign node6774 = (inp[8]) ? 8'b11110101 : node6775;
											assign node6775 = (inp[10]) ? 8'b10110001 : 8'b11111101;
								assign node6779 = (inp[8]) ? node6823 : node6780;
									assign node6780 = (inp[10]) ? node6800 : node6781;
										assign node6781 = (inp[1]) ? node6793 : node6782;
											assign node6782 = (inp[12]) ? node6786 : node6783;
												assign node6783 = (inp[2]) ? 8'b10101001 : 8'b10111001;
												assign node6786 = (inp[2]) ? node6790 : node6787;
													assign node6787 = (inp[3]) ? 8'b10101100 : 8'b10101101;
													assign node6790 = (inp[3]) ? 8'b10111001 : 8'b10111100;
											assign node6793 = (inp[2]) ? node6797 : node6794;
												assign node6794 = (inp[12]) ? 8'b10101001 : 8'b10111000;
												assign node6797 = (inp[12]) ? 8'b10111000 : 8'b10101000;
										assign node6800 = (inp[1]) ? node6816 : node6801;
											assign node6801 = (inp[3]) ? node6809 : node6802;
												assign node6802 = (inp[12]) ? node6806 : node6803;
													assign node6803 = (inp[2]) ? 8'b10101000 : 8'b10111000;
													assign node6806 = (inp[2]) ? 8'b10111000 : 8'b10101001;
												assign node6809 = (inp[2]) ? node6813 : node6810;
													assign node6810 = (inp[12]) ? 8'b10100000 : 8'b10010101;
													assign node6813 = (inp[12]) ? 8'b10010101 : 8'b10000101;
											assign node6816 = (inp[12]) ? node6820 : node6817;
												assign node6817 = (inp[2]) ? 8'b10000100 : 8'b10010100;
												assign node6820 = (inp[2]) ? 8'b10010100 : 8'b10000101;
									assign node6823 = (inp[1]) ? node6839 : node6824;
										assign node6824 = (inp[3]) ? node6832 : node6825;
											assign node6825 = (inp[12]) ? node6829 : node6826;
												assign node6826 = (inp[2]) ? 8'b10001100 : 8'b10011100;
												assign node6829 = (inp[2]) ? 8'b10011100 : 8'b10001101;
											assign node6832 = (inp[12]) ? node6836 : node6833;
												assign node6833 = (inp[2]) ? 8'b10000001 : 8'b10010001;
												assign node6836 = (inp[2]) ? 8'b10010001 : 8'b10000100;
										assign node6839 = (inp[2]) ? node6843 : node6840;
											assign node6840 = (inp[12]) ? 8'b10000001 : 8'b10010000;
											assign node6843 = (inp[12]) ? 8'b10010000 : 8'b10000000;
			assign node6846 = (inp[11]) ? node7254 : node6847;
				assign node6847 = (inp[5]) ? node7035 : node6848;
					assign node6848 = (inp[0]) ? node6852 : node6849;
						assign node6849 = (inp[12]) ? 8'b00000010 : 8'b10000010;
						assign node6852 = (inp[13]) ? node6930 : node6853;
							assign node6853 = (inp[10]) ? node6901 : node6854;
								assign node6854 = (inp[8]) ? node6884 : node6855;
									assign node6855 = (inp[6]) ? node6873 : node6856;
										assign node6856 = (inp[2]) ? node6868 : node6857;
											assign node6857 = (inp[12]) ? node6863 : node6858;
												assign node6858 = (inp[3]) ? 8'b10000010 : node6859;
													assign node6859 = (inp[1]) ? 8'b10000001 : 8'b10000010;
												assign node6863 = (inp[1]) ? node6865 : 8'b00000010;
													assign node6865 = (inp[9]) ? 8'b00000010 : 8'b10000001;
											assign node6868 = (inp[3]) ? 8'b10010000 : node6869;
												assign node6869 = (inp[1]) ? 8'b10010001 : 8'b10010000;
										assign node6873 = (inp[12]) ? node6879 : node6874;
											assign node6874 = (inp[1]) ? node6876 : 8'b10000010;
												assign node6876 = (inp[3]) ? 8'b10000010 : 8'b10000001;
											assign node6879 = (inp[1]) ? node6881 : 8'b00000010;
												assign node6881 = (inp[3]) ? 8'b00000010 : 8'b10000001;
									assign node6884 = (inp[1]) ? node6890 : node6885;
										assign node6885 = (inp[2]) ? node6887 : 8'b10000100;
											assign node6887 = (inp[6]) ? 8'b10000100 : 8'b10010100;
										assign node6890 = (inp[3]) ? node6896 : node6891;
											assign node6891 = (inp[2]) ? node6893 : 8'b10000101;
												assign node6893 = (inp[6]) ? 8'b10000101 : 8'b10010101;
											assign node6896 = (inp[6]) ? 8'b10000100 : node6897;
												assign node6897 = (inp[2]) ? 8'b10010100 : 8'b10000100;
								assign node6901 = (inp[2]) ? node6913 : node6902;
									assign node6902 = (inp[12]) ? node6908 : node6903;
										assign node6903 = (inp[3]) ? 8'b10000010 : node6904;
											assign node6904 = (inp[1]) ? 8'b10000001 : 8'b10000010;
										assign node6908 = (inp[1]) ? node6910 : 8'b00000010;
											assign node6910 = (inp[3]) ? 8'b00000010 : 8'b10000001;
									assign node6913 = (inp[6]) ? node6919 : node6914;
										assign node6914 = (inp[1]) ? node6916 : 8'b10010000;
											assign node6916 = (inp[3]) ? 8'b10010000 : 8'b10010001;
										assign node6919 = (inp[12]) ? node6925 : node6920;
											assign node6920 = (inp[1]) ? node6922 : 8'b10000010;
												assign node6922 = (inp[3]) ? 8'b10000010 : 8'b10000001;
											assign node6925 = (inp[1]) ? node6927 : 8'b00000010;
												assign node6927 = (inp[3]) ? 8'b00000010 : 8'b10000001;
							assign node6930 = (inp[9]) ? node6974 : node6931;
								assign node6931 = (inp[3]) ? node6957 : node6932;
									assign node6932 = (inp[1]) ? node6946 : node6933;
										assign node6933 = (inp[10]) ? node6941 : node6934;
											assign node6934 = (inp[8]) ? node6936 : 8'b10100000;
												assign node6936 = (inp[2]) ? node6938 : 8'b10100100;
													assign node6938 = (inp[6]) ? 8'b10100100 : 8'b10110100;
											assign node6941 = (inp[2]) ? node6943 : 8'b10100000;
												assign node6943 = (inp[6]) ? 8'b10100000 : 8'b10110000;
										assign node6946 = (inp[10]) ? node6952 : node6947;
											assign node6947 = (inp[8]) ? node6949 : 8'b10100001;
												assign node6949 = (inp[2]) ? 8'b11110101 : 8'b10100101;
											assign node6952 = (inp[6]) ? 8'b10100001 : node6953;
												assign node6953 = (inp[2]) ? 8'b10110001 : 8'b10100001;
									assign node6957 = (inp[6]) ? node6969 : node6958;
										assign node6958 = (inp[2]) ? node6964 : node6959;
											assign node6959 = (inp[10]) ? 8'b10100000 : node6960;
												assign node6960 = (inp[8]) ? 8'b10100100 : 8'b10100000;
											assign node6964 = (inp[10]) ? 8'b10110000 : node6965;
												assign node6965 = (inp[8]) ? 8'b10110100 : 8'b10110000;
										assign node6969 = (inp[8]) ? node6971 : 8'b10100000;
											assign node6971 = (inp[10]) ? 8'b10100000 : 8'b10100100;
								assign node6974 = (inp[6]) ? node7008 : node6975;
									assign node6975 = (inp[2]) ? node6993 : node6976;
										assign node6976 = (inp[8]) ? node6984 : node6977;
											assign node6977 = (inp[12]) ? 8'b00000010 : node6978;
												assign node6978 = (inp[1]) ? node6980 : 8'b10000010;
													assign node6980 = (inp[3]) ? 8'b10000010 : 8'b10000001;
											assign node6984 = (inp[10]) ? node6990 : node6985;
												assign node6985 = (inp[3]) ? 8'b10000100 : node6986;
													assign node6986 = (inp[1]) ? 8'b10000101 : 8'b10000100;
												assign node6990 = (inp[1]) ? 8'b10000001 : 8'b00000010;
										assign node6993 = (inp[10]) ? node7003 : node6994;
											assign node6994 = (inp[8]) ? node6998 : node6995;
												assign node6995 = (inp[3]) ? 8'b10010000 : 8'b10010001;
												assign node6998 = (inp[3]) ? 8'b10010100 : node6999;
													assign node6999 = (inp[1]) ? 8'b10010101 : 8'b10010100;
											assign node7003 = (inp[1]) ? node7005 : 8'b10010000;
												assign node7005 = (inp[3]) ? 8'b10010000 : 8'b10010001;
									assign node7008 = (inp[10]) ? node7024 : node7009;
										assign node7009 = (inp[8]) ? node7019 : node7010;
											assign node7010 = (inp[3]) ? node7016 : node7011;
												assign node7011 = (inp[1]) ? 8'b10000001 : node7012;
													assign node7012 = (inp[12]) ? 8'b00000010 : 8'b10000010;
												assign node7016 = (inp[12]) ? 8'b00000010 : 8'b10000010;
											assign node7019 = (inp[3]) ? 8'b10000100 : node7020;
												assign node7020 = (inp[1]) ? 8'b10000101 : 8'b10000100;
										assign node7024 = (inp[12]) ? node7030 : node7025;
											assign node7025 = (inp[3]) ? 8'b10000010 : node7026;
												assign node7026 = (inp[1]) ? 8'b10000001 : 8'b10000010;
											assign node7030 = (inp[3]) ? 8'b00000010 : node7031;
												assign node7031 = (inp[1]) ? 8'b10000001 : 8'b00000010;
					assign node7035 = (inp[8]) ? node7117 : node7036;
						assign node7036 = (inp[1]) ? node7068 : node7037;
							assign node7037 = (inp[13]) ? node7049 : node7038;
								assign node7038 = (inp[2]) ? node7042 : node7039;
									assign node7039 = (inp[12]) ? 8'b00000010 : 8'b10000010;
									assign node7042 = (inp[0]) ? 8'b10010000 : node7043;
										assign node7043 = (inp[6]) ? 8'b10010000 : node7044;
											assign node7044 = (inp[12]) ? 8'b00000010 : 8'b10000010;
								assign node7049 = (inp[2]) ? node7057 : node7050;
									assign node7050 = (inp[0]) ? 8'b10100000 : node7051;
										assign node7051 = (inp[9]) ? 8'b10100000 : node7052;
											assign node7052 = (inp[12]) ? 8'b00000010 : 8'b10000010;
									assign node7057 = (inp[0]) ? 8'b10110000 : node7058;
										assign node7058 = (inp[6]) ? node7064 : node7059;
											assign node7059 = (inp[9]) ? 8'b10100000 : node7060;
												assign node7060 = (inp[12]) ? 8'b00000010 : 8'b10000010;
											assign node7064 = (inp[9]) ? 8'b10110000 : 8'b10010000;
							assign node7068 = (inp[2]) ? node7088 : node7069;
								assign node7069 = (inp[13]) ? node7077 : node7070;
									assign node7070 = (inp[3]) ? 8'b10000001 : node7071;
										assign node7071 = (inp[0]) ? 8'b10000001 : node7072;
											assign node7072 = (inp[12]) ? 8'b00000010 : 8'b10000010;
									assign node7077 = (inp[0]) ? 8'b10100001 : node7078;
										assign node7078 = (inp[3]) ? node7084 : node7079;
											assign node7079 = (inp[9]) ? 8'b10100000 : node7080;
												assign node7080 = (inp[12]) ? 8'b00000010 : 8'b10000010;
											assign node7084 = (inp[9]) ? 8'b10100001 : 8'b10000001;
								assign node7088 = (inp[0]) ? node7114 : node7089;
									assign node7089 = (inp[6]) ? node7103 : node7090;
										assign node7090 = (inp[3]) ? node7098 : node7091;
											assign node7091 = (inp[12]) ? 8'b00000010 : node7092;
												assign node7092 = (inp[13]) ? node7094 : 8'b10000010;
													assign node7094 = (inp[9]) ? 8'b10100000 : 8'b10000010;
											assign node7098 = (inp[13]) ? node7100 : 8'b10000001;
												assign node7100 = (inp[9]) ? 8'b10100001 : 8'b10000001;
										assign node7103 = (inp[3]) ? node7109 : node7104;
											assign node7104 = (inp[9]) ? node7106 : 8'b10010000;
												assign node7106 = (inp[13]) ? 8'b10110000 : 8'b10010000;
											assign node7109 = (inp[13]) ? node7111 : 8'b10010001;
												assign node7111 = (inp[9]) ? 8'b10110001 : 8'b10010001;
									assign node7114 = (inp[13]) ? 8'b10110001 : 8'b10010001;
						assign node7117 = (inp[13]) ? node7169 : node7118;
							assign node7118 = (inp[2]) ? node7138 : node7119;
								assign node7119 = (inp[1]) ? node7127 : node7120;
									assign node7120 = (inp[10]) ? 8'b10000100 : node7121;
										assign node7121 = (inp[0]) ? 8'b10000100 : node7122;
											assign node7122 = (inp[12]) ? 8'b00000010 : 8'b10000010;
									assign node7127 = (inp[0]) ? 8'b10000101 : node7128;
										assign node7128 = (inp[10]) ? node7134 : node7129;
											assign node7129 = (inp[3]) ? 8'b10000001 : node7130;
												assign node7130 = (inp[12]) ? 8'b00000010 : 8'b10000010;
											assign node7134 = (inp[3]) ? 8'b10000101 : 8'b10000100;
								assign node7138 = (inp[0]) ? node7166 : node7139;
									assign node7139 = (inp[10]) ? node7155 : node7140;
										assign node7140 = (inp[6]) ? node7150 : node7141;
											assign node7141 = (inp[9]) ? node7147 : node7142;
												assign node7142 = (inp[1]) ? node7144 : 8'b10000010;
													assign node7144 = (inp[3]) ? 8'b10000001 : 8'b10000010;
												assign node7147 = (inp[12]) ? 8'b00000010 : 8'b10000010;
											assign node7150 = (inp[1]) ? node7152 : 8'b10010000;
												assign node7152 = (inp[3]) ? 8'b10010001 : 8'b10010000;
										assign node7155 = (inp[6]) ? node7161 : node7156;
											assign node7156 = (inp[1]) ? node7158 : 8'b10000100;
												assign node7158 = (inp[3]) ? 8'b10000101 : 8'b10000100;
											assign node7161 = (inp[1]) ? node7163 : 8'b10010100;
												assign node7163 = (inp[3]) ? 8'b10010101 : 8'b10010100;
									assign node7166 = (inp[1]) ? 8'b10010101 : 8'b10010100;
							assign node7169 = (inp[0]) ? node7247 : node7170;
								assign node7170 = (inp[10]) ? node7212 : node7171;
									assign node7171 = (inp[9]) ? node7195 : node7172;
										assign node7172 = (inp[6]) ? node7184 : node7173;
											assign node7173 = (inp[12]) ? node7179 : node7174;
												assign node7174 = (inp[3]) ? node7176 : 8'b10000010;
													assign node7176 = (inp[1]) ? 8'b10000001 : 8'b10000010;
												assign node7179 = (inp[1]) ? node7181 : 8'b00000010;
													assign node7181 = (inp[3]) ? 8'b10000001 : 8'b00000010;
											assign node7184 = (inp[2]) ? node7190 : node7185;
												assign node7185 = (inp[3]) ? node7187 : 8'b00000010;
													assign node7187 = (inp[1]) ? 8'b10000001 : 8'b10000010;
												assign node7190 = (inp[1]) ? node7192 : 8'b10010000;
													assign node7192 = (inp[3]) ? 8'b10010001 : 8'b10010000;
										assign node7195 = (inp[3]) ? node7201 : node7196;
											assign node7196 = (inp[6]) ? node7198 : 8'b10100000;
												assign node7198 = (inp[2]) ? 8'b10110000 : 8'b10100000;
											assign node7201 = (inp[1]) ? node7207 : node7202;
												assign node7202 = (inp[6]) ? node7204 : 8'b10100000;
													assign node7204 = (inp[12]) ? 8'b10110000 : 8'b10100000;
												assign node7207 = (inp[6]) ? node7209 : 8'b10100001;
													assign node7209 = (inp[2]) ? 8'b10110001 : 8'b10100001;
									assign node7212 = (inp[9]) ? node7230 : node7213;
										assign node7213 = (inp[6]) ? node7219 : node7214;
											assign node7214 = (inp[1]) ? node7216 : 8'b10000100;
												assign node7216 = (inp[3]) ? 8'b10000101 : 8'b10000100;
											assign node7219 = (inp[2]) ? node7225 : node7220;
												assign node7220 = (inp[3]) ? node7222 : 8'b10000100;
													assign node7222 = (inp[1]) ? 8'b10000101 : 8'b10000100;
												assign node7225 = (inp[3]) ? node7227 : 8'b10010100;
													assign node7227 = (inp[1]) ? 8'b10010101 : 8'b10010100;
										assign node7230 = (inp[6]) ? node7236 : node7231;
											assign node7231 = (inp[3]) ? node7233 : 8'b10100100;
												assign node7233 = (inp[1]) ? 8'b10100101 : 8'b10100100;
											assign node7236 = (inp[2]) ? node7242 : node7237;
												assign node7237 = (inp[3]) ? node7239 : 8'b10100100;
													assign node7239 = (inp[12]) ? 8'b10100100 : 8'b10100101;
												assign node7242 = (inp[1]) ? node7244 : 8'b10110100;
													assign node7244 = (inp[3]) ? 8'b11110101 : 8'b10110100;
								assign node7247 = (inp[1]) ? node7251 : node7248;
									assign node7248 = (inp[2]) ? 8'b10110100 : 8'b10100100;
									assign node7251 = (inp[2]) ? 8'b11110101 : 8'b10100101;
				assign node7254 = (inp[12]) ? node7564 : node7255;
					assign node7255 = (inp[5]) ? node7397 : node7256;
						assign node7256 = (inp[0]) ? node7258 : 8'b11110111;
							assign node7258 = (inp[2]) ? node7308 : node7259;
								assign node7259 = (inp[10]) ? node7291 : node7260;
									assign node7260 = (inp[8]) ? node7276 : node7261;
										assign node7261 = (inp[3]) ? node7271 : node7262;
											assign node7262 = (inp[1]) ? node7266 : node7263;
												assign node7263 = (inp[13]) ? 8'b10010101 : 8'b11110111;
												assign node7266 = (inp[9]) ? 8'b10110100 : node7267;
													assign node7267 = (inp[13]) ? 8'b10010100 : 8'b10110100;
											assign node7271 = (inp[9]) ? 8'b11110111 : node7272;
												assign node7272 = (inp[13]) ? 8'b10010101 : 8'b11110111;
										assign node7276 = (inp[1]) ? node7282 : node7277;
											assign node7277 = (inp[9]) ? 8'b10110001 : node7278;
												assign node7278 = (inp[13]) ? 8'b10010001 : 8'b10110001;
											assign node7282 = (inp[3]) ? node7288 : node7283;
												assign node7283 = (inp[9]) ? 8'b10110000 : node7284;
													assign node7284 = (inp[13]) ? 8'b10010000 : 8'b10110000;
												assign node7288 = (inp[13]) ? 8'b10010001 : 8'b10110001;
									assign node7291 = (inp[13]) ? node7297 : node7292;
										assign node7292 = (inp[1]) ? node7294 : 8'b11110111;
											assign node7294 = (inp[3]) ? 8'b11110111 : 8'b10110100;
										assign node7297 = (inp[9]) ? node7303 : node7298;
											assign node7298 = (inp[3]) ? 8'b10010101 : node7299;
												assign node7299 = (inp[1]) ? 8'b10010100 : 8'b10010101;
											assign node7303 = (inp[1]) ? node7305 : 8'b11110111;
												assign node7305 = (inp[3]) ? 8'b11110111 : 8'b10110100;
								assign node7308 = (inp[6]) ? node7354 : node7309;
									assign node7309 = (inp[3]) ? node7337 : node7310;
										assign node7310 = (inp[1]) ? node7322 : node7311;
											assign node7311 = (inp[8]) ? node7317 : node7312;
												assign node7312 = (inp[9]) ? 8'b10100101 : node7313;
													assign node7313 = (inp[13]) ? 8'b10000101 : 8'b10100101;
												assign node7317 = (inp[10]) ? node7319 : 8'b10100001;
													assign node7319 = (inp[13]) ? 8'b10000101 : 8'b10100101;
											assign node7322 = (inp[9]) ? node7332 : node7323;
												assign node7323 = (inp[13]) ? node7327 : node7324;
													assign node7324 = (inp[10]) ? 8'b10100100 : 8'b10100000;
													assign node7327 = (inp[8]) ? node7329 : 8'b10000100;
														assign node7329 = (inp[10]) ? 8'b10000100 : 8'b10000000;
												assign node7332 = (inp[10]) ? 8'b10100100 : node7333;
													assign node7333 = (inp[8]) ? 8'b10100000 : 8'b10100100;
										assign node7337 = (inp[13]) ? node7343 : node7338;
											assign node7338 = (inp[8]) ? node7340 : 8'b10100101;
												assign node7340 = (inp[10]) ? 8'b10100101 : 8'b10100001;
											assign node7343 = (inp[9]) ? node7349 : node7344;
												assign node7344 = (inp[10]) ? 8'b10000101 : node7345;
													assign node7345 = (inp[8]) ? 8'b10000001 : 8'b10000101;
												assign node7349 = (inp[10]) ? 8'b10100101 : node7350;
													assign node7350 = (inp[8]) ? 8'b10100001 : 8'b10100101;
									assign node7354 = (inp[8]) ? node7372 : node7355;
										assign node7355 = (inp[9]) ? node7367 : node7356;
											assign node7356 = (inp[13]) ? node7362 : node7357;
												assign node7357 = (inp[3]) ? 8'b11110111 : node7358;
													assign node7358 = (inp[1]) ? 8'b10110100 : 8'b11110111;
												assign node7362 = (inp[1]) ? node7364 : 8'b10010101;
													assign node7364 = (inp[3]) ? 8'b10010101 : 8'b10010100;
											assign node7367 = (inp[1]) ? node7369 : 8'b11110111;
												assign node7369 = (inp[3]) ? 8'b11110111 : 8'b10110100;
										assign node7372 = (inp[10]) ? node7384 : node7373;
											assign node7373 = (inp[9]) ? node7381 : node7374;
												assign node7374 = (inp[13]) ? node7376 : 8'b10110001;
													assign node7376 = (inp[3]) ? 8'b10010001 : node7377;
														assign node7377 = (inp[1]) ? 8'b10010000 : 8'b10010001;
												assign node7381 = (inp[1]) ? 8'b10110000 : 8'b10110001;
											assign node7384 = (inp[13]) ? node7390 : node7385;
												assign node7385 = (inp[1]) ? node7387 : 8'b11110111;
													assign node7387 = (inp[3]) ? 8'b11110111 : 8'b10110100;
												assign node7390 = (inp[9]) ? node7394 : node7391;
													assign node7391 = (inp[3]) ? 8'b10010101 : 8'b10010100;
													assign node7394 = (inp[1]) ? 8'b10110100 : 8'b11110111;
						assign node7397 = (inp[1]) ? node7465 : node7398;
							assign node7398 = (inp[2]) ? node7424 : node7399;
								assign node7399 = (inp[8]) ? node7407 : node7400;
									assign node7400 = (inp[13]) ? node7402 : 8'b11110111;
										assign node7402 = (inp[9]) ? 8'b10010101 : node7403;
											assign node7403 = (inp[0]) ? 8'b10010101 : 8'b11110111;
									assign node7407 = (inp[10]) ? node7417 : node7408;
										assign node7408 = (inp[0]) ? node7414 : node7409;
											assign node7409 = (inp[9]) ? node7411 : 8'b11110111;
												assign node7411 = (inp[13]) ? 8'b10010101 : 8'b11110111;
											assign node7414 = (inp[13]) ? 8'b10010001 : 8'b10110001;
										assign node7417 = (inp[13]) ? node7419 : 8'b10110001;
											assign node7419 = (inp[0]) ? 8'b10010001 : node7420;
												assign node7420 = (inp[9]) ? 8'b10010001 : 8'b10110001;
								assign node7424 = (inp[13]) ? node7440 : node7425;
									assign node7425 = (inp[0]) ? node7437 : node7426;
										assign node7426 = (inp[6]) ? node7432 : node7427;
											assign node7427 = (inp[10]) ? node7429 : 8'b11110111;
												assign node7429 = (inp[8]) ? 8'b10110001 : 8'b11110111;
											assign node7432 = (inp[8]) ? node7434 : 8'b10100101;
												assign node7434 = (inp[10]) ? 8'b10100001 : 8'b10100101;
										assign node7437 = (inp[8]) ? 8'b10100001 : 8'b10100101;
									assign node7440 = (inp[0]) ? node7462 : node7441;
										assign node7441 = (inp[6]) ? node7451 : node7442;
											assign node7442 = (inp[9]) ? node7446 : node7443;
												assign node7443 = (inp[8]) ? 8'b10110001 : 8'b11110111;
												assign node7446 = (inp[8]) ? node7448 : 8'b10010101;
													assign node7448 = (inp[10]) ? 8'b10010001 : 8'b10010101;
											assign node7451 = (inp[9]) ? node7457 : node7452;
												assign node7452 = (inp[8]) ? node7454 : 8'b10100101;
													assign node7454 = (inp[10]) ? 8'b10100001 : 8'b10100101;
												assign node7457 = (inp[3]) ? 8'b10000101 : node7458;
													assign node7458 = (inp[10]) ? 8'b10000001 : 8'b10000101;
										assign node7462 = (inp[8]) ? 8'b10000001 : 8'b10000101;
							assign node7465 = (inp[13]) ? node7509 : node7466;
								assign node7466 = (inp[8]) ? node7482 : node7467;
									assign node7467 = (inp[2]) ? node7473 : node7468;
										assign node7468 = (inp[0]) ? 8'b10110100 : node7469;
											assign node7469 = (inp[3]) ? 8'b10110100 : 8'b11110111;
										assign node7473 = (inp[0]) ? 8'b10100100 : node7474;
											assign node7474 = (inp[6]) ? node7478 : node7475;
												assign node7475 = (inp[3]) ? 8'b10110100 : 8'b11110111;
												assign node7478 = (inp[3]) ? 8'b10100100 : 8'b10100101;
									assign node7482 = (inp[2]) ? node7492 : node7483;
										assign node7483 = (inp[0]) ? 8'b10110000 : node7484;
											assign node7484 = (inp[10]) ? node7488 : node7485;
												assign node7485 = (inp[3]) ? 8'b10110100 : 8'b11110111;
												assign node7488 = (inp[3]) ? 8'b10110000 : 8'b10110001;
										assign node7492 = (inp[0]) ? 8'b10100000 : node7493;
											assign node7493 = (inp[3]) ? node7501 : node7494;
												assign node7494 = (inp[10]) ? node7498 : node7495;
													assign node7495 = (inp[6]) ? 8'b10100101 : 8'b11110111;
													assign node7498 = (inp[6]) ? 8'b10100001 : 8'b10110001;
												assign node7501 = (inp[6]) ? node7505 : node7502;
													assign node7502 = (inp[10]) ? 8'b10110000 : 8'b10110100;
													assign node7505 = (inp[10]) ? 8'b10100000 : 8'b10100100;
								assign node7509 = (inp[0]) ? node7557 : node7510;
									assign node7510 = (inp[9]) ? node7534 : node7511;
										assign node7511 = (inp[3]) ? node7525 : node7512;
											assign node7512 = (inp[6]) ? node7518 : node7513;
												assign node7513 = (inp[8]) ? node7515 : 8'b11110111;
													assign node7515 = (inp[10]) ? 8'b10110001 : 8'b11110111;
												assign node7518 = (inp[2]) ? 8'b10100101 : node7519;
													assign node7519 = (inp[10]) ? node7521 : 8'b11110111;
														assign node7521 = (inp[8]) ? 8'b10110001 : 8'b11110111;
											assign node7525 = (inp[6]) ? node7531 : node7526;
												assign node7526 = (inp[8]) ? node7528 : 8'b10110100;
													assign node7528 = (inp[10]) ? 8'b10110000 : 8'b10110100;
												assign node7531 = (inp[2]) ? 8'b10100100 : 8'b10110100;
										assign node7534 = (inp[3]) ? node7546 : node7535;
											assign node7535 = (inp[2]) ? node7541 : node7536;
												assign node7536 = (inp[8]) ? node7538 : 8'b10010101;
													assign node7538 = (inp[10]) ? 8'b10010001 : 8'b10010101;
												assign node7541 = (inp[6]) ? node7543 : 8'b10010101;
													assign node7543 = (inp[10]) ? 8'b10000001 : 8'b10000101;
											assign node7546 = (inp[8]) ? node7548 : 8'b10010100;
												assign node7548 = (inp[10]) ? node7554 : node7549;
													assign node7549 = (inp[6]) ? node7551 : 8'b10010100;
														assign node7551 = (inp[2]) ? 8'b10000100 : 8'b10010100;
													assign node7554 = (inp[6]) ? 8'b10000000 : 8'b10010000;
									assign node7557 = (inp[2]) ? node7561 : node7558;
										assign node7558 = (inp[8]) ? 8'b10010000 : 8'b10010100;
										assign node7561 = (inp[8]) ? 8'b10000000 : 8'b10000100;
					assign node7564 = (inp[5]) ? node7698 : node7565;
						assign node7565 = (inp[0]) ? node7567 : 8'b00000010;
							assign node7567 = (inp[6]) ? node7649 : node7568;
								assign node7568 = (inp[2]) ? node7612 : node7569;
									assign node7569 = (inp[1]) ? node7587 : node7570;
										assign node7570 = (inp[8]) ? node7576 : node7571;
											assign node7571 = (inp[13]) ? node7573 : 8'b00000010;
												assign node7573 = (inp[9]) ? 8'b00000010 : 8'b10100000;
											assign node7576 = (inp[10]) ? node7582 : node7577;
												assign node7577 = (inp[13]) ? node7579 : 8'b10100100;
													assign node7579 = (inp[9]) ? 8'b10100100 : 8'b10000100;
												assign node7582 = (inp[13]) ? node7584 : 8'b00000010;
													assign node7584 = (inp[9]) ? 8'b00000010 : 8'b10100000;
										assign node7587 = (inp[3]) ? node7599 : node7588;
											assign node7588 = (inp[9]) ? node7594 : node7589;
												assign node7589 = (inp[13]) ? node7591 : 8'b10100101;
													assign node7591 = (inp[8]) ? 8'b10000001 : 8'b10000101;
												assign node7594 = (inp[10]) ? 8'b10100101 : node7595;
													assign node7595 = (inp[8]) ? 8'b10100001 : 8'b10100101;
											assign node7599 = (inp[13]) ? node7605 : node7600;
												assign node7600 = (inp[8]) ? node7602 : 8'b00000010;
													assign node7602 = (inp[10]) ? 8'b00000010 : 8'b10100100;
												assign node7605 = (inp[8]) ? node7607 : 8'b10100000;
													assign node7607 = (inp[10]) ? 8'b10100000 : node7608;
														assign node7608 = (inp[9]) ? 8'b10100100 : 8'b10000100;
									assign node7612 = (inp[13]) ? node7630 : node7613;
										assign node7613 = (inp[1]) ? node7619 : node7614;
											assign node7614 = (inp[10]) ? 8'b11110101 : node7615;
												assign node7615 = (inp[8]) ? 8'b10110001 : 8'b11110101;
											assign node7619 = (inp[3]) ? node7625 : node7620;
												assign node7620 = (inp[8]) ? node7622 : 8'b10110100;
													assign node7622 = (inp[10]) ? 8'b10110100 : 8'b10110000;
												assign node7625 = (inp[10]) ? 8'b11110101 : node7626;
													assign node7626 = (inp[8]) ? 8'b10110001 : 8'b11110101;
										assign node7630 = (inp[9]) ? node7640 : node7631;
											assign node7631 = (inp[1]) ? node7637 : node7632;
												assign node7632 = (inp[8]) ? node7634 : 8'b10010101;
													assign node7634 = (inp[10]) ? 8'b10010101 : 8'b10010001;
												assign node7637 = (inp[3]) ? 8'b10010101 : 8'b10010100;
											assign node7640 = (inp[10]) ? 8'b11110101 : node7641;
												assign node7641 = (inp[8]) ? node7645 : node7642;
													assign node7642 = (inp[3]) ? 8'b11110101 : 8'b10110100;
													assign node7645 = (inp[1]) ? 8'b10110000 : 8'b10110001;
								assign node7649 = (inp[1]) ? node7667 : node7650;
									assign node7650 = (inp[10]) ? node7662 : node7651;
										assign node7651 = (inp[8]) ? node7657 : node7652;
											assign node7652 = (inp[13]) ? node7654 : 8'b00000010;
												assign node7654 = (inp[9]) ? 8'b00000010 : 8'b10100000;
											assign node7657 = (inp[9]) ? 8'b10100100 : node7658;
												assign node7658 = (inp[13]) ? 8'b10000100 : 8'b10100100;
										assign node7662 = (inp[9]) ? 8'b00000010 : node7663;
											assign node7663 = (inp[13]) ? 8'b10100000 : 8'b00000010;
									assign node7667 = (inp[3]) ? node7681 : node7668;
										assign node7668 = (inp[10]) ? node7676 : node7669;
											assign node7669 = (inp[8]) ? node7671 : 8'b10100101;
												assign node7671 = (inp[13]) ? node7673 : 8'b10100001;
													assign node7673 = (inp[9]) ? 8'b10100001 : 8'b10000001;
											assign node7676 = (inp[13]) ? node7678 : 8'b10100101;
												assign node7678 = (inp[9]) ? 8'b10100101 : 8'b10000101;
										assign node7681 = (inp[8]) ? node7687 : node7682;
											assign node7682 = (inp[9]) ? 8'b00000010 : node7683;
												assign node7683 = (inp[13]) ? 8'b10100000 : 8'b00000010;
											assign node7687 = (inp[10]) ? node7693 : node7688;
												assign node7688 = (inp[13]) ? node7690 : 8'b10100100;
													assign node7690 = (inp[9]) ? 8'b10100100 : 8'b10000100;
												assign node7693 = (inp[9]) ? 8'b00000010 : node7694;
													assign node7694 = (inp[13]) ? 8'b10100000 : 8'b00000010;
						assign node7698 = (inp[2]) ? node7774 : node7699;
							assign node7699 = (inp[1]) ? node7725 : node7700;
								assign node7700 = (inp[8]) ? node7708 : node7701;
									assign node7701 = (inp[13]) ? node7703 : 8'b00000010;
										assign node7703 = (inp[9]) ? 8'b10100000 : node7704;
											assign node7704 = (inp[0]) ? 8'b10100000 : 8'b00000010;
									assign node7708 = (inp[10]) ? node7718 : node7709;
										assign node7709 = (inp[0]) ? node7715 : node7710;
											assign node7710 = (inp[9]) ? node7712 : 8'b00000010;
												assign node7712 = (inp[13]) ? 8'b10100000 : 8'b00000010;
											assign node7715 = (inp[13]) ? 8'b10000100 : 8'b10100100;
										assign node7718 = (inp[13]) ? node7720 : 8'b10100100;
											assign node7720 = (inp[9]) ? 8'b10000100 : node7721;
												assign node7721 = (inp[0]) ? 8'b10000100 : 8'b10100100;
								assign node7725 = (inp[3]) ? node7751 : node7726;
									assign node7726 = (inp[0]) ? node7744 : node7727;
										assign node7727 = (inp[10]) ? node7733 : node7728;
											assign node7728 = (inp[13]) ? node7730 : 8'b00000010;
												assign node7730 = (inp[9]) ? 8'b10100000 : 8'b00000010;
											assign node7733 = (inp[8]) ? node7739 : node7734;
												assign node7734 = (inp[13]) ? node7736 : 8'b00000010;
													assign node7736 = (inp[9]) ? 8'b10100000 : 8'b00000010;
												assign node7739 = (inp[9]) ? node7741 : 8'b10100100;
													assign node7741 = (inp[13]) ? 8'b10000100 : 8'b10100100;
										assign node7744 = (inp[8]) ? node7748 : node7745;
											assign node7745 = (inp[13]) ? 8'b10000101 : 8'b10100101;
											assign node7748 = (inp[13]) ? 8'b10000001 : 8'b10100001;
									assign node7751 = (inp[8]) ? node7759 : node7752;
										assign node7752 = (inp[13]) ? node7754 : 8'b10100101;
											assign node7754 = (inp[0]) ? 8'b10000101 : node7755;
												assign node7755 = (inp[9]) ? 8'b10000101 : 8'b10100101;
										assign node7759 = (inp[13]) ? node7765 : node7760;
											assign node7760 = (inp[10]) ? 8'b10100001 : node7761;
												assign node7761 = (inp[0]) ? 8'b10100001 : 8'b10100101;
											assign node7765 = (inp[0]) ? 8'b10000001 : node7766;
												assign node7766 = (inp[9]) ? node7770 : node7767;
													assign node7767 = (inp[10]) ? 8'b10100001 : 8'b10100101;
													assign node7770 = (inp[10]) ? 8'b10000001 : 8'b10000101;
							assign node7774 = (inp[6]) ? node7834 : node7775;
								assign node7775 = (inp[0]) ? node7819 : node7776;
									assign node7776 = (inp[1]) ? node7794 : node7777;
										assign node7777 = (inp[10]) ? node7783 : node7778;
											assign node7778 = (inp[13]) ? node7780 : 8'b00000010;
												assign node7780 = (inp[9]) ? 8'b10100000 : 8'b00000010;
											assign node7783 = (inp[8]) ? node7789 : node7784;
												assign node7784 = (inp[13]) ? node7786 : 8'b00000010;
													assign node7786 = (inp[9]) ? 8'b10100000 : 8'b00000010;
												assign node7789 = (inp[9]) ? node7791 : 8'b10100100;
													assign node7791 = (inp[13]) ? 8'b10000100 : 8'b10100100;
										assign node7794 = (inp[3]) ? node7808 : node7795;
											assign node7795 = (inp[13]) ? node7801 : node7796;
												assign node7796 = (inp[8]) ? node7798 : 8'b00000010;
													assign node7798 = (inp[10]) ? 8'b10100100 : 8'b00000010;
												assign node7801 = (inp[9]) ? node7803 : 8'b00000010;
													assign node7803 = (inp[10]) ? node7805 : 8'b10100000;
														assign node7805 = (inp[8]) ? 8'b10000100 : 8'b10100000;
											assign node7808 = (inp[10]) ? node7814 : node7809;
												assign node7809 = (inp[9]) ? node7811 : 8'b10100101;
													assign node7811 = (inp[13]) ? 8'b10000101 : 8'b10100101;
												assign node7814 = (inp[8]) ? 8'b10100001 : node7815;
													assign node7815 = (inp[9]) ? 8'b10000101 : 8'b10100101;
									assign node7819 = (inp[1]) ? node7827 : node7820;
										assign node7820 = (inp[13]) ? node7824 : node7821;
											assign node7821 = (inp[8]) ? 8'b10110001 : 8'b11110101;
											assign node7824 = (inp[8]) ? 8'b10010001 : 8'b10010101;
										assign node7827 = (inp[8]) ? node7831 : node7828;
											assign node7828 = (inp[13]) ? 8'b10010100 : 8'b10110100;
											assign node7831 = (inp[13]) ? 8'b10010000 : 8'b10110000;
								assign node7834 = (inp[8]) ? node7858 : node7835;
									assign node7835 = (inp[1]) ? node7843 : node7836;
										assign node7836 = (inp[13]) ? node7838 : 8'b11110101;
											assign node7838 = (inp[9]) ? 8'b10010101 : node7839;
												assign node7839 = (inp[0]) ? 8'b10010101 : 8'b11110101;
										assign node7843 = (inp[0]) ? node7855 : node7844;
											assign node7844 = (inp[3]) ? node7850 : node7845;
												assign node7845 = (inp[9]) ? node7847 : 8'b11110101;
													assign node7847 = (inp[13]) ? 8'b10010101 : 8'b11110101;
												assign node7850 = (inp[13]) ? node7852 : 8'b10110100;
													assign node7852 = (inp[9]) ? 8'b10010100 : 8'b10110100;
											assign node7855 = (inp[13]) ? 8'b10010100 : 8'b10110100;
									assign node7858 = (inp[1]) ? node7874 : node7859;
										assign node7859 = (inp[13]) ? node7865 : node7860;
											assign node7860 = (inp[0]) ? 8'b10110001 : node7861;
												assign node7861 = (inp[10]) ? 8'b10110001 : 8'b11110101;
											assign node7865 = (inp[0]) ? 8'b10010001 : node7866;
												assign node7866 = (inp[9]) ? node7870 : node7867;
													assign node7867 = (inp[10]) ? 8'b10110001 : 8'b11110101;
													assign node7870 = (inp[10]) ? 8'b10010001 : 8'b10010101;
										assign node7874 = (inp[0]) ? node7886 : node7875;
											assign node7875 = (inp[10]) ? node7879 : node7876;
												assign node7876 = (inp[3]) ? 8'b10110100 : 8'b11110101;
												assign node7879 = (inp[3]) ? 8'b10110000 : node7880;
													assign node7880 = (inp[9]) ? node7882 : 8'b10110001;
														assign node7882 = (inp[13]) ? 8'b10010001 : 8'b10110001;
											assign node7886 = (inp[13]) ? 8'b10010000 : 8'b10110000;

endmodule