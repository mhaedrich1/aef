module dtc_split33_bm25 (
	input  wire [14-1:0] inp,
	output wire [14-1:0] outp
);

	wire [14-1:0] node1;
	wire [14-1:0] node2;
	wire [14-1:0] node3;
	wire [14-1:0] node4;
	wire [14-1:0] node5;
	wire [14-1:0] node6;
	wire [14-1:0] node7;
	wire [14-1:0] node8;
	wire [14-1:0] node9;
	wire [14-1:0] node10;
	wire [14-1:0] node11;
	wire [14-1:0] node14;
	wire [14-1:0] node17;
	wire [14-1:0] node19;
	wire [14-1:0] node22;
	wire [14-1:0] node23;
	wire [14-1:0] node24;
	wire [14-1:0] node27;
	wire [14-1:0] node31;
	wire [14-1:0] node32;
	wire [14-1:0] node33;
	wire [14-1:0] node34;
	wire [14-1:0] node37;
	wire [14-1:0] node40;
	wire [14-1:0] node41;
	wire [14-1:0] node45;
	wire [14-1:0] node46;
	wire [14-1:0] node47;
	wire [14-1:0] node50;
	wire [14-1:0] node53;
	wire [14-1:0] node54;
	wire [14-1:0] node58;
	wire [14-1:0] node59;
	wire [14-1:0] node60;
	wire [14-1:0] node61;
	wire [14-1:0] node62;
	wire [14-1:0] node66;
	wire [14-1:0] node67;
	wire [14-1:0] node70;
	wire [14-1:0] node73;
	wire [14-1:0] node74;
	wire [14-1:0] node75;
	wire [14-1:0] node78;
	wire [14-1:0] node81;
	wire [14-1:0] node84;
	wire [14-1:0] node85;
	wire [14-1:0] node86;
	wire [14-1:0] node87;
	wire [14-1:0] node90;
	wire [14-1:0] node93;
	wire [14-1:0] node94;
	wire [14-1:0] node98;
	wire [14-1:0] node99;
	wire [14-1:0] node100;
	wire [14-1:0] node103;
	wire [14-1:0] node106;
	wire [14-1:0] node107;
	wire [14-1:0] node110;
	wire [14-1:0] node113;
	wire [14-1:0] node114;
	wire [14-1:0] node115;
	wire [14-1:0] node116;
	wire [14-1:0] node117;
	wire [14-1:0] node118;
	wire [14-1:0] node121;
	wire [14-1:0] node124;
	wire [14-1:0] node125;
	wire [14-1:0] node128;
	wire [14-1:0] node131;
	wire [14-1:0] node132;
	wire [14-1:0] node134;
	wire [14-1:0] node137;
	wire [14-1:0] node138;
	wire [14-1:0] node142;
	wire [14-1:0] node143;
	wire [14-1:0] node144;
	wire [14-1:0] node145;
	wire [14-1:0] node148;
	wire [14-1:0] node151;
	wire [14-1:0] node152;
	wire [14-1:0] node155;
	wire [14-1:0] node158;
	wire [14-1:0] node159;
	wire [14-1:0] node160;
	wire [14-1:0] node163;
	wire [14-1:0] node166;
	wire [14-1:0] node167;
	wire [14-1:0] node171;
	wire [14-1:0] node172;
	wire [14-1:0] node173;
	wire [14-1:0] node174;
	wire [14-1:0] node175;
	wire [14-1:0] node179;
	wire [14-1:0] node180;
	wire [14-1:0] node184;
	wire [14-1:0] node185;
	wire [14-1:0] node187;
	wire [14-1:0] node190;
	wire [14-1:0] node192;
	wire [14-1:0] node195;
	wire [14-1:0] node196;
	wire [14-1:0] node197;
	wire [14-1:0] node199;
	wire [14-1:0] node202;
	wire [14-1:0] node203;
	wire [14-1:0] node206;
	wire [14-1:0] node209;
	wire [14-1:0] node210;
	wire [14-1:0] node212;
	wire [14-1:0] node215;
	wire [14-1:0] node217;
	wire [14-1:0] node220;
	wire [14-1:0] node221;
	wire [14-1:0] node222;
	wire [14-1:0] node223;
	wire [14-1:0] node224;
	wire [14-1:0] node225;
	wire [14-1:0] node226;
	wire [14-1:0] node229;
	wire [14-1:0] node232;
	wire [14-1:0] node233;
	wire [14-1:0] node236;
	wire [14-1:0] node239;
	wire [14-1:0] node240;
	wire [14-1:0] node241;
	wire [14-1:0] node244;
	wire [14-1:0] node247;
	wire [14-1:0] node248;
	wire [14-1:0] node251;
	wire [14-1:0] node254;
	wire [14-1:0] node255;
	wire [14-1:0] node256;
	wire [14-1:0] node258;
	wire [14-1:0] node262;
	wire [14-1:0] node263;
	wire [14-1:0] node265;
	wire [14-1:0] node268;
	wire [14-1:0] node269;
	wire [14-1:0] node273;
	wire [14-1:0] node274;
	wire [14-1:0] node275;
	wire [14-1:0] node276;
	wire [14-1:0] node277;
	wire [14-1:0] node281;
	wire [14-1:0] node282;
	wire [14-1:0] node285;
	wire [14-1:0] node288;
	wire [14-1:0] node289;
	wire [14-1:0] node290;
	wire [14-1:0] node293;
	wire [14-1:0] node296;
	wire [14-1:0] node297;
	wire [14-1:0] node300;
	wire [14-1:0] node303;
	wire [14-1:0] node304;
	wire [14-1:0] node305;
	wire [14-1:0] node306;
	wire [14-1:0] node309;
	wire [14-1:0] node312;
	wire [14-1:0] node314;
	wire [14-1:0] node317;
	wire [14-1:0] node319;
	wire [14-1:0] node320;
	wire [14-1:0] node323;
	wire [14-1:0] node326;
	wire [14-1:0] node327;
	wire [14-1:0] node328;
	wire [14-1:0] node329;
	wire [14-1:0] node330;
	wire [14-1:0] node332;
	wire [14-1:0] node335;
	wire [14-1:0] node337;
	wire [14-1:0] node340;
	wire [14-1:0] node342;
	wire [14-1:0] node343;
	wire [14-1:0] node347;
	wire [14-1:0] node348;
	wire [14-1:0] node349;
	wire [14-1:0] node350;
	wire [14-1:0] node354;
	wire [14-1:0] node355;
	wire [14-1:0] node358;
	wire [14-1:0] node361;
	wire [14-1:0] node362;
	wire [14-1:0] node363;
	wire [14-1:0] node366;
	wire [14-1:0] node369;
	wire [14-1:0] node370;
	wire [14-1:0] node373;
	wire [14-1:0] node376;
	wire [14-1:0] node377;
	wire [14-1:0] node378;
	wire [14-1:0] node379;
	wire [14-1:0] node380;
	wire [14-1:0] node384;
	wire [14-1:0] node387;
	wire [14-1:0] node388;
	wire [14-1:0] node390;
	wire [14-1:0] node393;
	wire [14-1:0] node396;
	wire [14-1:0] node397;
	wire [14-1:0] node398;
	wire [14-1:0] node400;
	wire [14-1:0] node404;
	wire [14-1:0] node405;
	wire [14-1:0] node406;
	wire [14-1:0] node409;
	wire [14-1:0] node412;
	wire [14-1:0] node414;
	wire [14-1:0] node417;
	wire [14-1:0] node418;
	wire [14-1:0] node419;
	wire [14-1:0] node420;
	wire [14-1:0] node421;
	wire [14-1:0] node422;
	wire [14-1:0] node423;
	wire [14-1:0] node424;
	wire [14-1:0] node427;
	wire [14-1:0] node430;
	wire [14-1:0] node431;
	wire [14-1:0] node434;
	wire [14-1:0] node437;
	wire [14-1:0] node438;
	wire [14-1:0] node440;
	wire [14-1:0] node443;
	wire [14-1:0] node444;
	wire [14-1:0] node447;
	wire [14-1:0] node450;
	wire [14-1:0] node451;
	wire [14-1:0] node452;
	wire [14-1:0] node454;
	wire [14-1:0] node457;
	wire [14-1:0] node458;
	wire [14-1:0] node462;
	wire [14-1:0] node463;
	wire [14-1:0] node464;
	wire [14-1:0] node467;
	wire [14-1:0] node470;
	wire [14-1:0] node471;
	wire [14-1:0] node474;
	wire [14-1:0] node477;
	wire [14-1:0] node478;
	wire [14-1:0] node479;
	wire [14-1:0] node480;
	wire [14-1:0] node481;
	wire [14-1:0] node484;
	wire [14-1:0] node487;
	wire [14-1:0] node488;
	wire [14-1:0] node492;
	wire [14-1:0] node493;
	wire [14-1:0] node494;
	wire [14-1:0] node497;
	wire [14-1:0] node500;
	wire [14-1:0] node502;
	wire [14-1:0] node505;
	wire [14-1:0] node506;
	wire [14-1:0] node507;
	wire [14-1:0] node509;
	wire [14-1:0] node512;
	wire [14-1:0] node513;
	wire [14-1:0] node517;
	wire [14-1:0] node518;
	wire [14-1:0] node519;
	wire [14-1:0] node523;
	wire [14-1:0] node525;
	wire [14-1:0] node528;
	wire [14-1:0] node529;
	wire [14-1:0] node530;
	wire [14-1:0] node531;
	wire [14-1:0] node532;
	wire [14-1:0] node533;
	wire [14-1:0] node536;
	wire [14-1:0] node539;
	wire [14-1:0] node540;
	wire [14-1:0] node544;
	wire [14-1:0] node545;
	wire [14-1:0] node547;
	wire [14-1:0] node550;
	wire [14-1:0] node551;
	wire [14-1:0] node554;
	wire [14-1:0] node557;
	wire [14-1:0] node558;
	wire [14-1:0] node559;
	wire [14-1:0] node561;
	wire [14-1:0] node564;
	wire [14-1:0] node565;
	wire [14-1:0] node568;
	wire [14-1:0] node571;
	wire [14-1:0] node572;
	wire [14-1:0] node573;
	wire [14-1:0] node576;
	wire [14-1:0] node579;
	wire [14-1:0] node580;
	wire [14-1:0] node584;
	wire [14-1:0] node585;
	wire [14-1:0] node586;
	wire [14-1:0] node587;
	wire [14-1:0] node588;
	wire [14-1:0] node592;
	wire [14-1:0] node595;
	wire [14-1:0] node596;
	wire [14-1:0] node597;
	wire [14-1:0] node600;
	wire [14-1:0] node603;
	wire [14-1:0] node604;
	wire [14-1:0] node608;
	wire [14-1:0] node609;
	wire [14-1:0] node610;
	wire [14-1:0] node612;
	wire [14-1:0] node615;
	wire [14-1:0] node617;
	wire [14-1:0] node620;
	wire [14-1:0] node621;
	wire [14-1:0] node622;
	wire [14-1:0] node625;
	wire [14-1:0] node628;
	wire [14-1:0] node631;
	wire [14-1:0] node632;
	wire [14-1:0] node633;
	wire [14-1:0] node634;
	wire [14-1:0] node635;
	wire [14-1:0] node636;
	wire [14-1:0] node637;
	wire [14-1:0] node640;
	wire [14-1:0] node643;
	wire [14-1:0] node644;
	wire [14-1:0] node647;
	wire [14-1:0] node650;
	wire [14-1:0] node651;
	wire [14-1:0] node652;
	wire [14-1:0] node655;
	wire [14-1:0] node658;
	wire [14-1:0] node659;
	wire [14-1:0] node663;
	wire [14-1:0] node664;
	wire [14-1:0] node665;
	wire [14-1:0] node666;
	wire [14-1:0] node669;
	wire [14-1:0] node672;
	wire [14-1:0] node673;
	wire [14-1:0] node677;
	wire [14-1:0] node678;
	wire [14-1:0] node679;
	wire [14-1:0] node682;
	wire [14-1:0] node685;
	wire [14-1:0] node686;
	wire [14-1:0] node689;
	wire [14-1:0] node692;
	wire [14-1:0] node693;
	wire [14-1:0] node694;
	wire [14-1:0] node695;
	wire [14-1:0] node696;
	wire [14-1:0] node699;
	wire [14-1:0] node702;
	wire [14-1:0] node703;
	wire [14-1:0] node706;
	wire [14-1:0] node709;
	wire [14-1:0] node710;
	wire [14-1:0] node711;
	wire [14-1:0] node716;
	wire [14-1:0] node717;
	wire [14-1:0] node718;
	wire [14-1:0] node719;
	wire [14-1:0] node723;
	wire [14-1:0] node724;
	wire [14-1:0] node727;
	wire [14-1:0] node730;
	wire [14-1:0] node731;
	wire [14-1:0] node733;
	wire [14-1:0] node736;
	wire [14-1:0] node738;
	wire [14-1:0] node741;
	wire [14-1:0] node742;
	wire [14-1:0] node743;
	wire [14-1:0] node744;
	wire [14-1:0] node745;
	wire [14-1:0] node748;
	wire [14-1:0] node749;
	wire [14-1:0] node753;
	wire [14-1:0] node755;
	wire [14-1:0] node756;
	wire [14-1:0] node760;
	wire [14-1:0] node761;
	wire [14-1:0] node762;
	wire [14-1:0] node763;
	wire [14-1:0] node766;
	wire [14-1:0] node769;
	wire [14-1:0] node771;
	wire [14-1:0] node774;
	wire [14-1:0] node775;
	wire [14-1:0] node776;
	wire [14-1:0] node779;
	wire [14-1:0] node782;
	wire [14-1:0] node783;
	wire [14-1:0] node786;
	wire [14-1:0] node789;
	wire [14-1:0] node790;
	wire [14-1:0] node791;
	wire [14-1:0] node792;
	wire [14-1:0] node793;
	wire [14-1:0] node796;
	wire [14-1:0] node799;
	wire [14-1:0] node800;
	wire [14-1:0] node804;
	wire [14-1:0] node805;
	wire [14-1:0] node806;
	wire [14-1:0] node809;
	wire [14-1:0] node812;
	wire [14-1:0] node813;
	wire [14-1:0] node816;
	wire [14-1:0] node819;
	wire [14-1:0] node820;
	wire [14-1:0] node821;
	wire [14-1:0] node823;
	wire [14-1:0] node826;
	wire [14-1:0] node827;
	wire [14-1:0] node830;
	wire [14-1:0] node833;
	wire [14-1:0] node834;
	wire [14-1:0] node835;
	wire [14-1:0] node838;
	wire [14-1:0] node841;
	wire [14-1:0] node842;
	wire [14-1:0] node845;
	wire [14-1:0] node848;
	wire [14-1:0] node849;
	wire [14-1:0] node850;
	wire [14-1:0] node851;
	wire [14-1:0] node852;
	wire [14-1:0] node853;
	wire [14-1:0] node854;
	wire [14-1:0] node855;
	wire [14-1:0] node856;
	wire [14-1:0] node860;
	wire [14-1:0] node862;
	wire [14-1:0] node865;
	wire [14-1:0] node867;
	wire [14-1:0] node868;
	wire [14-1:0] node871;
	wire [14-1:0] node874;
	wire [14-1:0] node875;
	wire [14-1:0] node876;
	wire [14-1:0] node879;
	wire [14-1:0] node880;
	wire [14-1:0] node884;
	wire [14-1:0] node885;
	wire [14-1:0] node886;
	wire [14-1:0] node889;
	wire [14-1:0] node892;
	wire [14-1:0] node893;
	wire [14-1:0] node897;
	wire [14-1:0] node898;
	wire [14-1:0] node899;
	wire [14-1:0] node900;
	wire [14-1:0] node901;
	wire [14-1:0] node904;
	wire [14-1:0] node907;
	wire [14-1:0] node908;
	wire [14-1:0] node911;
	wire [14-1:0] node914;
	wire [14-1:0] node915;
	wire [14-1:0] node916;
	wire [14-1:0] node919;
	wire [14-1:0] node922;
	wire [14-1:0] node923;
	wire [14-1:0] node927;
	wire [14-1:0] node928;
	wire [14-1:0] node929;
	wire [14-1:0] node931;
	wire [14-1:0] node934;
	wire [14-1:0] node935;
	wire [14-1:0] node939;
	wire [14-1:0] node940;
	wire [14-1:0] node942;
	wire [14-1:0] node945;
	wire [14-1:0] node946;
	wire [14-1:0] node950;
	wire [14-1:0] node951;
	wire [14-1:0] node952;
	wire [14-1:0] node953;
	wire [14-1:0] node954;
	wire [14-1:0] node955;
	wire [14-1:0] node958;
	wire [14-1:0] node961;
	wire [14-1:0] node962;
	wire [14-1:0] node966;
	wire [14-1:0] node967;
	wire [14-1:0] node968;
	wire [14-1:0] node971;
	wire [14-1:0] node974;
	wire [14-1:0] node975;
	wire [14-1:0] node978;
	wire [14-1:0] node981;
	wire [14-1:0] node982;
	wire [14-1:0] node983;
	wire [14-1:0] node984;
	wire [14-1:0] node987;
	wire [14-1:0] node990;
	wire [14-1:0] node991;
	wire [14-1:0] node995;
	wire [14-1:0] node996;
	wire [14-1:0] node997;
	wire [14-1:0] node1000;
	wire [14-1:0] node1003;
	wire [14-1:0] node1004;
	wire [14-1:0] node1008;
	wire [14-1:0] node1009;
	wire [14-1:0] node1010;
	wire [14-1:0] node1011;
	wire [14-1:0] node1013;
	wire [14-1:0] node1016;
	wire [14-1:0] node1017;
	wire [14-1:0] node1021;
	wire [14-1:0] node1022;
	wire [14-1:0] node1023;
	wire [14-1:0] node1026;
	wire [14-1:0] node1029;
	wire [14-1:0] node1030;
	wire [14-1:0] node1033;
	wire [14-1:0] node1036;
	wire [14-1:0] node1037;
	wire [14-1:0] node1038;
	wire [14-1:0] node1040;
	wire [14-1:0] node1043;
	wire [14-1:0] node1044;
	wire [14-1:0] node1047;
	wire [14-1:0] node1050;
	wire [14-1:0] node1051;
	wire [14-1:0] node1054;
	wire [14-1:0] node1056;
	wire [14-1:0] node1059;
	wire [14-1:0] node1060;
	wire [14-1:0] node1061;
	wire [14-1:0] node1062;
	wire [14-1:0] node1063;
	wire [14-1:0] node1064;
	wire [14-1:0] node1065;
	wire [14-1:0] node1068;
	wire [14-1:0] node1071;
	wire [14-1:0] node1072;
	wire [14-1:0] node1076;
	wire [14-1:0] node1077;
	wire [14-1:0] node1079;
	wire [14-1:0] node1082;
	wire [14-1:0] node1083;
	wire [14-1:0] node1087;
	wire [14-1:0] node1088;
	wire [14-1:0] node1089;
	wire [14-1:0] node1091;
	wire [14-1:0] node1095;
	wire [14-1:0] node1096;
	wire [14-1:0] node1097;
	wire [14-1:0] node1101;
	wire [14-1:0] node1104;
	wire [14-1:0] node1105;
	wire [14-1:0] node1106;
	wire [14-1:0] node1107;
	wire [14-1:0] node1109;
	wire [14-1:0] node1112;
	wire [14-1:0] node1113;
	wire [14-1:0] node1116;
	wire [14-1:0] node1119;
	wire [14-1:0] node1120;
	wire [14-1:0] node1121;
	wire [14-1:0] node1124;
	wire [14-1:0] node1127;
	wire [14-1:0] node1130;
	wire [14-1:0] node1131;
	wire [14-1:0] node1132;
	wire [14-1:0] node1133;
	wire [14-1:0] node1136;
	wire [14-1:0] node1139;
	wire [14-1:0] node1141;
	wire [14-1:0] node1144;
	wire [14-1:0] node1145;
	wire [14-1:0] node1146;
	wire [14-1:0] node1150;
	wire [14-1:0] node1151;
	wire [14-1:0] node1154;
	wire [14-1:0] node1157;
	wire [14-1:0] node1158;
	wire [14-1:0] node1159;
	wire [14-1:0] node1160;
	wire [14-1:0] node1161;
	wire [14-1:0] node1162;
	wire [14-1:0] node1165;
	wire [14-1:0] node1168;
	wire [14-1:0] node1169;
	wire [14-1:0] node1172;
	wire [14-1:0] node1175;
	wire [14-1:0] node1176;
	wire [14-1:0] node1177;
	wire [14-1:0] node1180;
	wire [14-1:0] node1183;
	wire [14-1:0] node1185;
	wire [14-1:0] node1188;
	wire [14-1:0] node1189;
	wire [14-1:0] node1190;
	wire [14-1:0] node1191;
	wire [14-1:0] node1194;
	wire [14-1:0] node1197;
	wire [14-1:0] node1198;
	wire [14-1:0] node1201;
	wire [14-1:0] node1204;
	wire [14-1:0] node1205;
	wire [14-1:0] node1206;
	wire [14-1:0] node1210;
	wire [14-1:0] node1212;
	wire [14-1:0] node1215;
	wire [14-1:0] node1216;
	wire [14-1:0] node1217;
	wire [14-1:0] node1218;
	wire [14-1:0] node1221;
	wire [14-1:0] node1222;
	wire [14-1:0] node1226;
	wire [14-1:0] node1227;
	wire [14-1:0] node1230;
	wire [14-1:0] node1231;
	wire [14-1:0] node1234;
	wire [14-1:0] node1237;
	wire [14-1:0] node1238;
	wire [14-1:0] node1239;
	wire [14-1:0] node1241;
	wire [14-1:0] node1244;
	wire [14-1:0] node1245;
	wire [14-1:0] node1248;
	wire [14-1:0] node1251;
	wire [14-1:0] node1252;
	wire [14-1:0] node1253;
	wire [14-1:0] node1257;
	wire [14-1:0] node1259;
	wire [14-1:0] node1262;
	wire [14-1:0] node1263;
	wire [14-1:0] node1264;
	wire [14-1:0] node1265;
	wire [14-1:0] node1266;
	wire [14-1:0] node1267;
	wire [14-1:0] node1268;
	wire [14-1:0] node1270;
	wire [14-1:0] node1273;
	wire [14-1:0] node1276;
	wire [14-1:0] node1278;
	wire [14-1:0] node1279;
	wire [14-1:0] node1283;
	wire [14-1:0] node1284;
	wire [14-1:0] node1285;
	wire [14-1:0] node1287;
	wire [14-1:0] node1290;
	wire [14-1:0] node1291;
	wire [14-1:0] node1295;
	wire [14-1:0] node1296;
	wire [14-1:0] node1297;
	wire [14-1:0] node1300;
	wire [14-1:0] node1303;
	wire [14-1:0] node1304;
	wire [14-1:0] node1307;
	wire [14-1:0] node1310;
	wire [14-1:0] node1311;
	wire [14-1:0] node1312;
	wire [14-1:0] node1313;
	wire [14-1:0] node1314;
	wire [14-1:0] node1317;
	wire [14-1:0] node1320;
	wire [14-1:0] node1321;
	wire [14-1:0] node1324;
	wire [14-1:0] node1327;
	wire [14-1:0] node1328;
	wire [14-1:0] node1329;
	wire [14-1:0] node1332;
	wire [14-1:0] node1335;
	wire [14-1:0] node1336;
	wire [14-1:0] node1339;
	wire [14-1:0] node1342;
	wire [14-1:0] node1343;
	wire [14-1:0] node1344;
	wire [14-1:0] node1345;
	wire [14-1:0] node1348;
	wire [14-1:0] node1351;
	wire [14-1:0] node1352;
	wire [14-1:0] node1355;
	wire [14-1:0] node1358;
	wire [14-1:0] node1359;
	wire [14-1:0] node1362;
	wire [14-1:0] node1364;
	wire [14-1:0] node1367;
	wire [14-1:0] node1368;
	wire [14-1:0] node1369;
	wire [14-1:0] node1370;
	wire [14-1:0] node1371;
	wire [14-1:0] node1372;
	wire [14-1:0] node1376;
	wire [14-1:0] node1379;
	wire [14-1:0] node1381;
	wire [14-1:0] node1383;
	wire [14-1:0] node1386;
	wire [14-1:0] node1387;
	wire [14-1:0] node1388;
	wire [14-1:0] node1390;
	wire [14-1:0] node1393;
	wire [14-1:0] node1394;
	wire [14-1:0] node1397;
	wire [14-1:0] node1400;
	wire [14-1:0] node1401;
	wire [14-1:0] node1403;
	wire [14-1:0] node1406;
	wire [14-1:0] node1407;
	wire [14-1:0] node1411;
	wire [14-1:0] node1412;
	wire [14-1:0] node1413;
	wire [14-1:0] node1414;
	wire [14-1:0] node1415;
	wire [14-1:0] node1418;
	wire [14-1:0] node1421;
	wire [14-1:0] node1422;
	wire [14-1:0] node1427;
	wire [14-1:0] node1428;
	wire [14-1:0] node1429;
	wire [14-1:0] node1431;
	wire [14-1:0] node1434;
	wire [14-1:0] node1437;
	wire [14-1:0] node1438;
	wire [14-1:0] node1441;
	wire [14-1:0] node1442;
	wire [14-1:0] node1445;
	wire [14-1:0] node1448;
	wire [14-1:0] node1449;
	wire [14-1:0] node1450;
	wire [14-1:0] node1451;
	wire [14-1:0] node1452;
	wire [14-1:0] node1453;
	wire [14-1:0] node1454;
	wire [14-1:0] node1457;
	wire [14-1:0] node1460;
	wire [14-1:0] node1461;
	wire [14-1:0] node1465;
	wire [14-1:0] node1466;
	wire [14-1:0] node1467;
	wire [14-1:0] node1472;
	wire [14-1:0] node1473;
	wire [14-1:0] node1474;
	wire [14-1:0] node1475;
	wire [14-1:0] node1478;
	wire [14-1:0] node1481;
	wire [14-1:0] node1482;
	wire [14-1:0] node1485;
	wire [14-1:0] node1488;
	wire [14-1:0] node1489;
	wire [14-1:0] node1491;
	wire [14-1:0] node1494;
	wire [14-1:0] node1496;
	wire [14-1:0] node1499;
	wire [14-1:0] node1500;
	wire [14-1:0] node1501;
	wire [14-1:0] node1502;
	wire [14-1:0] node1503;
	wire [14-1:0] node1506;
	wire [14-1:0] node1510;
	wire [14-1:0] node1511;
	wire [14-1:0] node1512;
	wire [14-1:0] node1515;
	wire [14-1:0] node1518;
	wire [14-1:0] node1519;
	wire [14-1:0] node1522;
	wire [14-1:0] node1525;
	wire [14-1:0] node1526;
	wire [14-1:0] node1527;
	wire [14-1:0] node1530;
	wire [14-1:0] node1531;
	wire [14-1:0] node1534;
	wire [14-1:0] node1537;
	wire [14-1:0] node1538;
	wire [14-1:0] node1540;
	wire [14-1:0] node1543;
	wire [14-1:0] node1546;
	wire [14-1:0] node1547;
	wire [14-1:0] node1548;
	wire [14-1:0] node1549;
	wire [14-1:0] node1550;
	wire [14-1:0] node1551;
	wire [14-1:0] node1555;
	wire [14-1:0] node1556;
	wire [14-1:0] node1559;
	wire [14-1:0] node1562;
	wire [14-1:0] node1563;
	wire [14-1:0] node1565;
	wire [14-1:0] node1568;
	wire [14-1:0] node1570;
	wire [14-1:0] node1573;
	wire [14-1:0] node1574;
	wire [14-1:0] node1575;
	wire [14-1:0] node1576;
	wire [14-1:0] node1579;
	wire [14-1:0] node1582;
	wire [14-1:0] node1583;
	wire [14-1:0] node1586;
	wire [14-1:0] node1589;
	wire [14-1:0] node1590;
	wire [14-1:0] node1591;
	wire [14-1:0] node1595;
	wire [14-1:0] node1596;
	wire [14-1:0] node1599;
	wire [14-1:0] node1602;
	wire [14-1:0] node1603;
	wire [14-1:0] node1604;
	wire [14-1:0] node1605;
	wire [14-1:0] node1606;
	wire [14-1:0] node1610;
	wire [14-1:0] node1611;
	wire [14-1:0] node1614;
	wire [14-1:0] node1617;
	wire [14-1:0] node1619;
	wire [14-1:0] node1620;
	wire [14-1:0] node1624;
	wire [14-1:0] node1625;
	wire [14-1:0] node1626;
	wire [14-1:0] node1628;
	wire [14-1:0] node1631;
	wire [14-1:0] node1633;
	wire [14-1:0] node1636;
	wire [14-1:0] node1637;
	wire [14-1:0] node1638;
	wire [14-1:0] node1641;
	wire [14-1:0] node1644;
	wire [14-1:0] node1645;
	wire [14-1:0] node1648;
	wire [14-1:0] node1651;
	wire [14-1:0] node1652;
	wire [14-1:0] node1653;
	wire [14-1:0] node1654;
	wire [14-1:0] node1655;
	wire [14-1:0] node1656;
	wire [14-1:0] node1657;
	wire [14-1:0] node1658;
	wire [14-1:0] node1659;
	wire [14-1:0] node1660;
	wire [14-1:0] node1663;
	wire [14-1:0] node1666;
	wire [14-1:0] node1669;
	wire [14-1:0] node1670;
	wire [14-1:0] node1671;
	wire [14-1:0] node1675;
	wire [14-1:0] node1677;
	wire [14-1:0] node1680;
	wire [14-1:0] node1681;
	wire [14-1:0] node1682;
	wire [14-1:0] node1683;
	wire [14-1:0] node1687;
	wire [14-1:0] node1690;
	wire [14-1:0] node1691;
	wire [14-1:0] node1692;
	wire [14-1:0] node1696;
	wire [14-1:0] node1697;
	wire [14-1:0] node1700;
	wire [14-1:0] node1703;
	wire [14-1:0] node1704;
	wire [14-1:0] node1705;
	wire [14-1:0] node1706;
	wire [14-1:0] node1707;
	wire [14-1:0] node1710;
	wire [14-1:0] node1713;
	wire [14-1:0] node1715;
	wire [14-1:0] node1718;
	wire [14-1:0] node1719;
	wire [14-1:0] node1720;
	wire [14-1:0] node1723;
	wire [14-1:0] node1726;
	wire [14-1:0] node1727;
	wire [14-1:0] node1730;
	wire [14-1:0] node1733;
	wire [14-1:0] node1734;
	wire [14-1:0] node1736;
	wire [14-1:0] node1738;
	wire [14-1:0] node1741;
	wire [14-1:0] node1742;
	wire [14-1:0] node1743;
	wire [14-1:0] node1746;
	wire [14-1:0] node1749;
	wire [14-1:0] node1750;
	wire [14-1:0] node1754;
	wire [14-1:0] node1755;
	wire [14-1:0] node1756;
	wire [14-1:0] node1757;
	wire [14-1:0] node1758;
	wire [14-1:0] node1759;
	wire [14-1:0] node1764;
	wire [14-1:0] node1765;
	wire [14-1:0] node1766;
	wire [14-1:0] node1769;
	wire [14-1:0] node1772;
	wire [14-1:0] node1774;
	wire [14-1:0] node1777;
	wire [14-1:0] node1778;
	wire [14-1:0] node1779;
	wire [14-1:0] node1781;
	wire [14-1:0] node1784;
	wire [14-1:0] node1785;
	wire [14-1:0] node1788;
	wire [14-1:0] node1791;
	wire [14-1:0] node1793;
	wire [14-1:0] node1795;
	wire [14-1:0] node1798;
	wire [14-1:0] node1799;
	wire [14-1:0] node1800;
	wire [14-1:0] node1801;
	wire [14-1:0] node1802;
	wire [14-1:0] node1805;
	wire [14-1:0] node1809;
	wire [14-1:0] node1810;
	wire [14-1:0] node1811;
	wire [14-1:0] node1814;
	wire [14-1:0] node1817;
	wire [14-1:0] node1818;
	wire [14-1:0] node1821;
	wire [14-1:0] node1824;
	wire [14-1:0] node1825;
	wire [14-1:0] node1826;
	wire [14-1:0] node1827;
	wire [14-1:0] node1830;
	wire [14-1:0] node1833;
	wire [14-1:0] node1835;
	wire [14-1:0] node1838;
	wire [14-1:0] node1839;
	wire [14-1:0] node1841;
	wire [14-1:0] node1844;
	wire [14-1:0] node1846;
	wire [14-1:0] node1849;
	wire [14-1:0] node1850;
	wire [14-1:0] node1851;
	wire [14-1:0] node1852;
	wire [14-1:0] node1853;
	wire [14-1:0] node1854;
	wire [14-1:0] node1856;
	wire [14-1:0] node1859;
	wire [14-1:0] node1860;
	wire [14-1:0] node1863;
	wire [14-1:0] node1866;
	wire [14-1:0] node1867;
	wire [14-1:0] node1868;
	wire [14-1:0] node1871;
	wire [14-1:0] node1875;
	wire [14-1:0] node1876;
	wire [14-1:0] node1877;
	wire [14-1:0] node1878;
	wire [14-1:0] node1881;
	wire [14-1:0] node1884;
	wire [14-1:0] node1885;
	wire [14-1:0] node1888;
	wire [14-1:0] node1891;
	wire [14-1:0] node1892;
	wire [14-1:0] node1893;
	wire [14-1:0] node1897;
	wire [14-1:0] node1900;
	wire [14-1:0] node1901;
	wire [14-1:0] node1902;
	wire [14-1:0] node1903;
	wire [14-1:0] node1904;
	wire [14-1:0] node1908;
	wire [14-1:0] node1909;
	wire [14-1:0] node1912;
	wire [14-1:0] node1915;
	wire [14-1:0] node1916;
	wire [14-1:0] node1917;
	wire [14-1:0] node1920;
	wire [14-1:0] node1923;
	wire [14-1:0] node1926;
	wire [14-1:0] node1927;
	wire [14-1:0] node1928;
	wire [14-1:0] node1930;
	wire [14-1:0] node1933;
	wire [14-1:0] node1934;
	wire [14-1:0] node1938;
	wire [14-1:0] node1940;
	wire [14-1:0] node1941;
	wire [14-1:0] node1945;
	wire [14-1:0] node1946;
	wire [14-1:0] node1947;
	wire [14-1:0] node1948;
	wire [14-1:0] node1949;
	wire [14-1:0] node1951;
	wire [14-1:0] node1954;
	wire [14-1:0] node1955;
	wire [14-1:0] node1959;
	wire [14-1:0] node1960;
	wire [14-1:0] node1962;
	wire [14-1:0] node1966;
	wire [14-1:0] node1967;
	wire [14-1:0] node1968;
	wire [14-1:0] node1969;
	wire [14-1:0] node1972;
	wire [14-1:0] node1975;
	wire [14-1:0] node1976;
	wire [14-1:0] node1979;
	wire [14-1:0] node1982;
	wire [14-1:0] node1983;
	wire [14-1:0] node1985;
	wire [14-1:0] node1989;
	wire [14-1:0] node1990;
	wire [14-1:0] node1991;
	wire [14-1:0] node1992;
	wire [14-1:0] node1993;
	wire [14-1:0] node1996;
	wire [14-1:0] node1999;
	wire [14-1:0] node2000;
	wire [14-1:0] node2004;
	wire [14-1:0] node2005;
	wire [14-1:0] node2006;
	wire [14-1:0] node2010;
	wire [14-1:0] node2011;
	wire [14-1:0] node2014;
	wire [14-1:0] node2017;
	wire [14-1:0] node2018;
	wire [14-1:0] node2019;
	wire [14-1:0] node2020;
	wire [14-1:0] node2023;
	wire [14-1:0] node2027;
	wire [14-1:0] node2028;
	wire [14-1:0] node2030;
	wire [14-1:0] node2033;
	wire [14-1:0] node2034;
	wire [14-1:0] node2037;
	wire [14-1:0] node2040;
	wire [14-1:0] node2041;
	wire [14-1:0] node2042;
	wire [14-1:0] node2043;
	wire [14-1:0] node2044;
	wire [14-1:0] node2045;
	wire [14-1:0] node2046;
	wire [14-1:0] node2047;
	wire [14-1:0] node2051;
	wire [14-1:0] node2052;
	wire [14-1:0] node2055;
	wire [14-1:0] node2058;
	wire [14-1:0] node2059;
	wire [14-1:0] node2060;
	wire [14-1:0] node2063;
	wire [14-1:0] node2066;
	wire [14-1:0] node2069;
	wire [14-1:0] node2070;
	wire [14-1:0] node2071;
	wire [14-1:0] node2072;
	wire [14-1:0] node2077;
	wire [14-1:0] node2078;
	wire [14-1:0] node2079;
	wire [14-1:0] node2082;
	wire [14-1:0] node2085;
	wire [14-1:0] node2086;
	wire [14-1:0] node2089;
	wire [14-1:0] node2092;
	wire [14-1:0] node2093;
	wire [14-1:0] node2094;
	wire [14-1:0] node2095;
	wire [14-1:0] node2096;
	wire [14-1:0] node2099;
	wire [14-1:0] node2102;
	wire [14-1:0] node2103;
	wire [14-1:0] node2106;
	wire [14-1:0] node2109;
	wire [14-1:0] node2111;
	wire [14-1:0] node2112;
	wire [14-1:0] node2116;
	wire [14-1:0] node2117;
	wire [14-1:0] node2118;
	wire [14-1:0] node2119;
	wire [14-1:0] node2122;
	wire [14-1:0] node2125;
	wire [14-1:0] node2126;
	wire [14-1:0] node2130;
	wire [14-1:0] node2131;
	wire [14-1:0] node2132;
	wire [14-1:0] node2135;
	wire [14-1:0] node2138;
	wire [14-1:0] node2139;
	wire [14-1:0] node2143;
	wire [14-1:0] node2144;
	wire [14-1:0] node2145;
	wire [14-1:0] node2147;
	wire [14-1:0] node2148;
	wire [14-1:0] node2151;
	wire [14-1:0] node2152;
	wire [14-1:0] node2156;
	wire [14-1:0] node2157;
	wire [14-1:0] node2158;
	wire [14-1:0] node2159;
	wire [14-1:0] node2162;
	wire [14-1:0] node2166;
	wire [14-1:0] node2167;
	wire [14-1:0] node2168;
	wire [14-1:0] node2171;
	wire [14-1:0] node2174;
	wire [14-1:0] node2175;
	wire [14-1:0] node2179;
	wire [14-1:0] node2180;
	wire [14-1:0] node2181;
	wire [14-1:0] node2182;
	wire [14-1:0] node2183;
	wire [14-1:0] node2186;
	wire [14-1:0] node2189;
	wire [14-1:0] node2190;
	wire [14-1:0] node2193;
	wire [14-1:0] node2196;
	wire [14-1:0] node2197;
	wire [14-1:0] node2199;
	wire [14-1:0] node2202;
	wire [14-1:0] node2203;
	wire [14-1:0] node2206;
	wire [14-1:0] node2209;
	wire [14-1:0] node2210;
	wire [14-1:0] node2211;
	wire [14-1:0] node2212;
	wire [14-1:0] node2216;
	wire [14-1:0] node2217;
	wire [14-1:0] node2221;
	wire [14-1:0] node2222;
	wire [14-1:0] node2224;
	wire [14-1:0] node2227;
	wire [14-1:0] node2228;
	wire [14-1:0] node2232;
	wire [14-1:0] node2233;
	wire [14-1:0] node2234;
	wire [14-1:0] node2235;
	wire [14-1:0] node2236;
	wire [14-1:0] node2237;
	wire [14-1:0] node2240;
	wire [14-1:0] node2241;
	wire [14-1:0] node2245;
	wire [14-1:0] node2246;
	wire [14-1:0] node2247;
	wire [14-1:0] node2250;
	wire [14-1:0] node2253;
	wire [14-1:0] node2255;
	wire [14-1:0] node2258;
	wire [14-1:0] node2259;
	wire [14-1:0] node2260;
	wire [14-1:0] node2261;
	wire [14-1:0] node2264;
	wire [14-1:0] node2267;
	wire [14-1:0] node2268;
	wire [14-1:0] node2271;
	wire [14-1:0] node2274;
	wire [14-1:0] node2275;
	wire [14-1:0] node2276;
	wire [14-1:0] node2279;
	wire [14-1:0] node2282;
	wire [14-1:0] node2284;
	wire [14-1:0] node2287;
	wire [14-1:0] node2288;
	wire [14-1:0] node2289;
	wire [14-1:0] node2290;
	wire [14-1:0] node2291;
	wire [14-1:0] node2295;
	wire [14-1:0] node2296;
	wire [14-1:0] node2299;
	wire [14-1:0] node2302;
	wire [14-1:0] node2303;
	wire [14-1:0] node2304;
	wire [14-1:0] node2307;
	wire [14-1:0] node2310;
	wire [14-1:0] node2311;
	wire [14-1:0] node2314;
	wire [14-1:0] node2317;
	wire [14-1:0] node2318;
	wire [14-1:0] node2319;
	wire [14-1:0] node2320;
	wire [14-1:0] node2323;
	wire [14-1:0] node2326;
	wire [14-1:0] node2327;
	wire [14-1:0] node2330;
	wire [14-1:0] node2333;
	wire [14-1:0] node2334;
	wire [14-1:0] node2336;
	wire [14-1:0] node2339;
	wire [14-1:0] node2341;
	wire [14-1:0] node2344;
	wire [14-1:0] node2345;
	wire [14-1:0] node2346;
	wire [14-1:0] node2347;
	wire [14-1:0] node2348;
	wire [14-1:0] node2350;
	wire [14-1:0] node2353;
	wire [14-1:0] node2354;
	wire [14-1:0] node2358;
	wire [14-1:0] node2359;
	wire [14-1:0] node2363;
	wire [14-1:0] node2364;
	wire [14-1:0] node2365;
	wire [14-1:0] node2367;
	wire [14-1:0] node2370;
	wire [14-1:0] node2372;
	wire [14-1:0] node2375;
	wire [14-1:0] node2376;
	wire [14-1:0] node2378;
	wire [14-1:0] node2382;
	wire [14-1:0] node2383;
	wire [14-1:0] node2384;
	wire [14-1:0] node2385;
	wire [14-1:0] node2388;
	wire [14-1:0] node2389;
	wire [14-1:0] node2393;
	wire [14-1:0] node2394;
	wire [14-1:0] node2395;
	wire [14-1:0] node2398;
	wire [14-1:0] node2401;
	wire [14-1:0] node2403;
	wire [14-1:0] node2406;
	wire [14-1:0] node2407;
	wire [14-1:0] node2408;
	wire [14-1:0] node2410;
	wire [14-1:0] node2413;
	wire [14-1:0] node2414;
	wire [14-1:0] node2417;
	wire [14-1:0] node2420;
	wire [14-1:0] node2421;
	wire [14-1:0] node2423;
	wire [14-1:0] node2426;
	wire [14-1:0] node2427;
	wire [14-1:0] node2430;
	wire [14-1:0] node2433;
	wire [14-1:0] node2434;
	wire [14-1:0] node2435;
	wire [14-1:0] node2436;
	wire [14-1:0] node2437;
	wire [14-1:0] node2438;
	wire [14-1:0] node2439;
	wire [14-1:0] node2440;
	wire [14-1:0] node2443;
	wire [14-1:0] node2445;
	wire [14-1:0] node2448;
	wire [14-1:0] node2449;
	wire [14-1:0] node2450;
	wire [14-1:0] node2454;
	wire [14-1:0] node2455;
	wire [14-1:0] node2458;
	wire [14-1:0] node2461;
	wire [14-1:0] node2462;
	wire [14-1:0] node2464;
	wire [14-1:0] node2467;
	wire [14-1:0] node2468;
	wire [14-1:0] node2469;
	wire [14-1:0] node2472;
	wire [14-1:0] node2475;
	wire [14-1:0] node2476;
	wire [14-1:0] node2479;
	wire [14-1:0] node2482;
	wire [14-1:0] node2483;
	wire [14-1:0] node2484;
	wire [14-1:0] node2486;
	wire [14-1:0] node2487;
	wire [14-1:0] node2491;
	wire [14-1:0] node2492;
	wire [14-1:0] node2493;
	wire [14-1:0] node2497;
	wire [14-1:0] node2498;
	wire [14-1:0] node2501;
	wire [14-1:0] node2504;
	wire [14-1:0] node2505;
	wire [14-1:0] node2506;
	wire [14-1:0] node2508;
	wire [14-1:0] node2511;
	wire [14-1:0] node2512;
	wire [14-1:0] node2516;
	wire [14-1:0] node2517;
	wire [14-1:0] node2519;
	wire [14-1:0] node2522;
	wire [14-1:0] node2525;
	wire [14-1:0] node2526;
	wire [14-1:0] node2527;
	wire [14-1:0] node2528;
	wire [14-1:0] node2529;
	wire [14-1:0] node2530;
	wire [14-1:0] node2535;
	wire [14-1:0] node2536;
	wire [14-1:0] node2537;
	wire [14-1:0] node2541;
	wire [14-1:0] node2542;
	wire [14-1:0] node2546;
	wire [14-1:0] node2547;
	wire [14-1:0] node2548;
	wire [14-1:0] node2549;
	wire [14-1:0] node2552;
	wire [14-1:0] node2555;
	wire [14-1:0] node2558;
	wire [14-1:0] node2559;
	wire [14-1:0] node2560;
	wire [14-1:0] node2563;
	wire [14-1:0] node2566;
	wire [14-1:0] node2567;
	wire [14-1:0] node2571;
	wire [14-1:0] node2572;
	wire [14-1:0] node2573;
	wire [14-1:0] node2574;
	wire [14-1:0] node2576;
	wire [14-1:0] node2579;
	wire [14-1:0] node2580;
	wire [14-1:0] node2583;
	wire [14-1:0] node2586;
	wire [14-1:0] node2587;
	wire [14-1:0] node2588;
	wire [14-1:0] node2591;
	wire [14-1:0] node2594;
	wire [14-1:0] node2595;
	wire [14-1:0] node2598;
	wire [14-1:0] node2601;
	wire [14-1:0] node2602;
	wire [14-1:0] node2603;
	wire [14-1:0] node2605;
	wire [14-1:0] node2608;
	wire [14-1:0] node2609;
	wire [14-1:0] node2612;
	wire [14-1:0] node2615;
	wire [14-1:0] node2616;
	wire [14-1:0] node2620;
	wire [14-1:0] node2621;
	wire [14-1:0] node2622;
	wire [14-1:0] node2623;
	wire [14-1:0] node2624;
	wire [14-1:0] node2625;
	wire [14-1:0] node2627;
	wire [14-1:0] node2630;
	wire [14-1:0] node2631;
	wire [14-1:0] node2635;
	wire [14-1:0] node2636;
	wire [14-1:0] node2638;
	wire [14-1:0] node2641;
	wire [14-1:0] node2642;
	wire [14-1:0] node2646;
	wire [14-1:0] node2647;
	wire [14-1:0] node2648;
	wire [14-1:0] node2650;
	wire [14-1:0] node2653;
	wire [14-1:0] node2654;
	wire [14-1:0] node2657;
	wire [14-1:0] node2660;
	wire [14-1:0] node2661;
	wire [14-1:0] node2662;
	wire [14-1:0] node2665;
	wire [14-1:0] node2669;
	wire [14-1:0] node2670;
	wire [14-1:0] node2671;
	wire [14-1:0] node2672;
	wire [14-1:0] node2673;
	wire [14-1:0] node2676;
	wire [14-1:0] node2679;
	wire [14-1:0] node2680;
	wire [14-1:0] node2683;
	wire [14-1:0] node2686;
	wire [14-1:0] node2688;
	wire [14-1:0] node2689;
	wire [14-1:0] node2693;
	wire [14-1:0] node2694;
	wire [14-1:0] node2695;
	wire [14-1:0] node2696;
	wire [14-1:0] node2699;
	wire [14-1:0] node2702;
	wire [14-1:0] node2703;
	wire [14-1:0] node2707;
	wire [14-1:0] node2708;
	wire [14-1:0] node2710;
	wire [14-1:0] node2713;
	wire [14-1:0] node2715;
	wire [14-1:0] node2718;
	wire [14-1:0] node2719;
	wire [14-1:0] node2720;
	wire [14-1:0] node2721;
	wire [14-1:0] node2722;
	wire [14-1:0] node2723;
	wire [14-1:0] node2728;
	wire [14-1:0] node2729;
	wire [14-1:0] node2730;
	wire [14-1:0] node2734;
	wire [14-1:0] node2735;
	wire [14-1:0] node2739;
	wire [14-1:0] node2740;
	wire [14-1:0] node2741;
	wire [14-1:0] node2742;
	wire [14-1:0] node2745;
	wire [14-1:0] node2748;
	wire [14-1:0] node2750;
	wire [14-1:0] node2753;
	wire [14-1:0] node2754;
	wire [14-1:0] node2756;
	wire [14-1:0] node2759;
	wire [14-1:0] node2761;
	wire [14-1:0] node2764;
	wire [14-1:0] node2765;
	wire [14-1:0] node2766;
	wire [14-1:0] node2767;
	wire [14-1:0] node2769;
	wire [14-1:0] node2772;
	wire [14-1:0] node2773;
	wire [14-1:0] node2776;
	wire [14-1:0] node2779;
	wire [14-1:0] node2780;
	wire [14-1:0] node2781;
	wire [14-1:0] node2785;
	wire [14-1:0] node2786;
	wire [14-1:0] node2789;
	wire [14-1:0] node2792;
	wire [14-1:0] node2793;
	wire [14-1:0] node2794;
	wire [14-1:0] node2796;
	wire [14-1:0] node2800;
	wire [14-1:0] node2801;
	wire [14-1:0] node2803;
	wire [14-1:0] node2806;
	wire [14-1:0] node2807;
	wire [14-1:0] node2810;
	wire [14-1:0] node2813;
	wire [14-1:0] node2814;
	wire [14-1:0] node2815;
	wire [14-1:0] node2816;
	wire [14-1:0] node2817;
	wire [14-1:0] node2818;
	wire [14-1:0] node2819;
	wire [14-1:0] node2820;
	wire [14-1:0] node2823;
	wire [14-1:0] node2827;
	wire [14-1:0] node2828;
	wire [14-1:0] node2829;
	wire [14-1:0] node2832;
	wire [14-1:0] node2835;
	wire [14-1:0] node2836;
	wire [14-1:0] node2840;
	wire [14-1:0] node2841;
	wire [14-1:0] node2843;
	wire [14-1:0] node2844;
	wire [14-1:0] node2847;
	wire [14-1:0] node2850;
	wire [14-1:0] node2851;
	wire [14-1:0] node2853;
	wire [14-1:0] node2857;
	wire [14-1:0] node2858;
	wire [14-1:0] node2859;
	wire [14-1:0] node2860;
	wire [14-1:0] node2861;
	wire [14-1:0] node2865;
	wire [14-1:0] node2866;
	wire [14-1:0] node2869;
	wire [14-1:0] node2872;
	wire [14-1:0] node2873;
	wire [14-1:0] node2874;
	wire [14-1:0] node2877;
	wire [14-1:0] node2880;
	wire [14-1:0] node2883;
	wire [14-1:0] node2884;
	wire [14-1:0] node2885;
	wire [14-1:0] node2887;
	wire [14-1:0] node2890;
	wire [14-1:0] node2892;
	wire [14-1:0] node2895;
	wire [14-1:0] node2896;
	wire [14-1:0] node2897;
	wire [14-1:0] node2901;
	wire [14-1:0] node2902;
	wire [14-1:0] node2906;
	wire [14-1:0] node2907;
	wire [14-1:0] node2908;
	wire [14-1:0] node2909;
	wire [14-1:0] node2910;
	wire [14-1:0] node2911;
	wire [14-1:0] node2915;
	wire [14-1:0] node2917;
	wire [14-1:0] node2920;
	wire [14-1:0] node2921;
	wire [14-1:0] node2922;
	wire [14-1:0] node2925;
	wire [14-1:0] node2928;
	wire [14-1:0] node2929;
	wire [14-1:0] node2933;
	wire [14-1:0] node2934;
	wire [14-1:0] node2935;
	wire [14-1:0] node2936;
	wire [14-1:0] node2939;
	wire [14-1:0] node2942;
	wire [14-1:0] node2944;
	wire [14-1:0] node2947;
	wire [14-1:0] node2948;
	wire [14-1:0] node2949;
	wire [14-1:0] node2953;
	wire [14-1:0] node2955;
	wire [14-1:0] node2958;
	wire [14-1:0] node2959;
	wire [14-1:0] node2960;
	wire [14-1:0] node2961;
	wire [14-1:0] node2963;
	wire [14-1:0] node2966;
	wire [14-1:0] node2969;
	wire [14-1:0] node2970;
	wire [14-1:0] node2971;
	wire [14-1:0] node2974;
	wire [14-1:0] node2977;
	wire [14-1:0] node2978;
	wire [14-1:0] node2982;
	wire [14-1:0] node2983;
	wire [14-1:0] node2984;
	wire [14-1:0] node2986;
	wire [14-1:0] node2990;
	wire [14-1:0] node2991;
	wire [14-1:0] node2995;
	wire [14-1:0] node2996;
	wire [14-1:0] node2997;
	wire [14-1:0] node2998;
	wire [14-1:0] node2999;
	wire [14-1:0] node3000;
	wire [14-1:0] node3003;
	wire [14-1:0] node3004;
	wire [14-1:0] node3008;
	wire [14-1:0] node3010;
	wire [14-1:0] node3011;
	wire [14-1:0] node3015;
	wire [14-1:0] node3016;
	wire [14-1:0] node3017;
	wire [14-1:0] node3018;
	wire [14-1:0] node3022;
	wire [14-1:0] node3023;
	wire [14-1:0] node3026;
	wire [14-1:0] node3029;
	wire [14-1:0] node3030;
	wire [14-1:0] node3031;
	wire [14-1:0] node3034;
	wire [14-1:0] node3037;
	wire [14-1:0] node3038;
	wire [14-1:0] node3042;
	wire [14-1:0] node3043;
	wire [14-1:0] node3044;
	wire [14-1:0] node3045;
	wire [14-1:0] node3046;
	wire [14-1:0] node3049;
	wire [14-1:0] node3052;
	wire [14-1:0] node3054;
	wire [14-1:0] node3057;
	wire [14-1:0] node3058;
	wire [14-1:0] node3061;
	wire [14-1:0] node3062;
	wire [14-1:0] node3066;
	wire [14-1:0] node3067;
	wire [14-1:0] node3068;
	wire [14-1:0] node3069;
	wire [14-1:0] node3073;
	wire [14-1:0] node3074;
	wire [14-1:0] node3078;
	wire [14-1:0] node3079;
	wire [14-1:0] node3080;
	wire [14-1:0] node3083;
	wire [14-1:0] node3086;
	wire [14-1:0] node3087;
	wire [14-1:0] node3090;
	wire [14-1:0] node3093;
	wire [14-1:0] node3094;
	wire [14-1:0] node3095;
	wire [14-1:0] node3096;
	wire [14-1:0] node3097;
	wire [14-1:0] node3099;
	wire [14-1:0] node3102;
	wire [14-1:0] node3104;
	wire [14-1:0] node3107;
	wire [14-1:0] node3108;
	wire [14-1:0] node3110;
	wire [14-1:0] node3113;
	wire [14-1:0] node3114;
	wire [14-1:0] node3118;
	wire [14-1:0] node3119;
	wire [14-1:0] node3120;
	wire [14-1:0] node3121;
	wire [14-1:0] node3124;
	wire [14-1:0] node3127;
	wire [14-1:0] node3128;
	wire [14-1:0] node3131;
	wire [14-1:0] node3134;
	wire [14-1:0] node3135;
	wire [14-1:0] node3137;
	wire [14-1:0] node3140;
	wire [14-1:0] node3141;
	wire [14-1:0] node3144;
	wire [14-1:0] node3147;
	wire [14-1:0] node3148;
	wire [14-1:0] node3149;
	wire [14-1:0] node3150;
	wire [14-1:0] node3152;
	wire [14-1:0] node3155;
	wire [14-1:0] node3157;
	wire [14-1:0] node3160;
	wire [14-1:0] node3161;
	wire [14-1:0] node3162;
	wire [14-1:0] node3165;
	wire [14-1:0] node3168;
	wire [14-1:0] node3169;
	wire [14-1:0] node3173;
	wire [14-1:0] node3174;
	wire [14-1:0] node3175;
	wire [14-1:0] node3177;
	wire [14-1:0] node3180;
	wire [14-1:0] node3181;
	wire [14-1:0] node3184;
	wire [14-1:0] node3187;
	wire [14-1:0] node3188;
	wire [14-1:0] node3189;
	wire [14-1:0] node3192;
	wire [14-1:0] node3195;
	wire [14-1:0] node3196;
	wire [14-1:0] node3199;
	wire [14-1:0] node3202;
	wire [14-1:0] node3203;
	wire [14-1:0] node3204;
	wire [14-1:0] node3205;
	wire [14-1:0] node3206;
	wire [14-1:0] node3207;
	wire [14-1:0] node3208;
	wire [14-1:0] node3209;
	wire [14-1:0] node3210;
	wire [14-1:0] node3211;
	wire [14-1:0] node3212;
	wire [14-1:0] node3216;
	wire [14-1:0] node3217;
	wire [14-1:0] node3220;
	wire [14-1:0] node3223;
	wire [14-1:0] node3224;
	wire [14-1:0] node3225;
	wire [14-1:0] node3228;
	wire [14-1:0] node3231;
	wire [14-1:0] node3232;
	wire [14-1:0] node3235;
	wire [14-1:0] node3238;
	wire [14-1:0] node3239;
	wire [14-1:0] node3240;
	wire [14-1:0] node3241;
	wire [14-1:0] node3244;
	wire [14-1:0] node3247;
	wire [14-1:0] node3248;
	wire [14-1:0] node3251;
	wire [14-1:0] node3254;
	wire [14-1:0] node3255;
	wire [14-1:0] node3256;
	wire [14-1:0] node3260;
	wire [14-1:0] node3261;
	wire [14-1:0] node3265;
	wire [14-1:0] node3266;
	wire [14-1:0] node3267;
	wire [14-1:0] node3268;
	wire [14-1:0] node3270;
	wire [14-1:0] node3273;
	wire [14-1:0] node3274;
	wire [14-1:0] node3277;
	wire [14-1:0] node3280;
	wire [14-1:0] node3281;
	wire [14-1:0] node3282;
	wire [14-1:0] node3285;
	wire [14-1:0] node3288;
	wire [14-1:0] node3290;
	wire [14-1:0] node3293;
	wire [14-1:0] node3294;
	wire [14-1:0] node3295;
	wire [14-1:0] node3296;
	wire [14-1:0] node3299;
	wire [14-1:0] node3302;
	wire [14-1:0] node3303;
	wire [14-1:0] node3306;
	wire [14-1:0] node3309;
	wire [14-1:0] node3310;
	wire [14-1:0] node3312;
	wire [14-1:0] node3315;
	wire [14-1:0] node3316;
	wire [14-1:0] node3320;
	wire [14-1:0] node3321;
	wire [14-1:0] node3322;
	wire [14-1:0] node3323;
	wire [14-1:0] node3324;
	wire [14-1:0] node3325;
	wire [14-1:0] node3329;
	wire [14-1:0] node3330;
	wire [14-1:0] node3334;
	wire [14-1:0] node3335;
	wire [14-1:0] node3336;
	wire [14-1:0] node3339;
	wire [14-1:0] node3342;
	wire [14-1:0] node3343;
	wire [14-1:0] node3346;
	wire [14-1:0] node3349;
	wire [14-1:0] node3350;
	wire [14-1:0] node3351;
	wire [14-1:0] node3353;
	wire [14-1:0] node3356;
	wire [14-1:0] node3357;
	wire [14-1:0] node3360;
	wire [14-1:0] node3363;
	wire [14-1:0] node3364;
	wire [14-1:0] node3366;
	wire [14-1:0] node3369;
	wire [14-1:0] node3370;
	wire [14-1:0] node3373;
	wire [14-1:0] node3376;
	wire [14-1:0] node3377;
	wire [14-1:0] node3378;
	wire [14-1:0] node3379;
	wire [14-1:0] node3380;
	wire [14-1:0] node3383;
	wire [14-1:0] node3386;
	wire [14-1:0] node3387;
	wire [14-1:0] node3391;
	wire [14-1:0] node3392;
	wire [14-1:0] node3393;
	wire [14-1:0] node3396;
	wire [14-1:0] node3399;
	wire [14-1:0] node3400;
	wire [14-1:0] node3403;
	wire [14-1:0] node3406;
	wire [14-1:0] node3407;
	wire [14-1:0] node3408;
	wire [14-1:0] node3409;
	wire [14-1:0] node3412;
	wire [14-1:0] node3415;
	wire [14-1:0] node3418;
	wire [14-1:0] node3419;
	wire [14-1:0] node3421;
	wire [14-1:0] node3424;
	wire [14-1:0] node3425;
	wire [14-1:0] node3429;
	wire [14-1:0] node3430;
	wire [14-1:0] node3431;
	wire [14-1:0] node3432;
	wire [14-1:0] node3433;
	wire [14-1:0] node3434;
	wire [14-1:0] node3435;
	wire [14-1:0] node3438;
	wire [14-1:0] node3441;
	wire [14-1:0] node3442;
	wire [14-1:0] node3445;
	wire [14-1:0] node3448;
	wire [14-1:0] node3449;
	wire [14-1:0] node3450;
	wire [14-1:0] node3453;
	wire [14-1:0] node3456;
	wire [14-1:0] node3457;
	wire [14-1:0] node3460;
	wire [14-1:0] node3463;
	wire [14-1:0] node3464;
	wire [14-1:0] node3465;
	wire [14-1:0] node3466;
	wire [14-1:0] node3469;
	wire [14-1:0] node3473;
	wire [14-1:0] node3474;
	wire [14-1:0] node3475;
	wire [14-1:0] node3479;
	wire [14-1:0] node3480;
	wire [14-1:0] node3484;
	wire [14-1:0] node3485;
	wire [14-1:0] node3486;
	wire [14-1:0] node3487;
	wire [14-1:0] node3488;
	wire [14-1:0] node3491;
	wire [14-1:0] node3494;
	wire [14-1:0] node3495;
	wire [14-1:0] node3498;
	wire [14-1:0] node3501;
	wire [14-1:0] node3502;
	wire [14-1:0] node3503;
	wire [14-1:0] node3506;
	wire [14-1:0] node3509;
	wire [14-1:0] node3512;
	wire [14-1:0] node3513;
	wire [14-1:0] node3514;
	wire [14-1:0] node3515;
	wire [14-1:0] node3518;
	wire [14-1:0] node3521;
	wire [14-1:0] node3523;
	wire [14-1:0] node3526;
	wire [14-1:0] node3527;
	wire [14-1:0] node3528;
	wire [14-1:0] node3531;
	wire [14-1:0] node3534;
	wire [14-1:0] node3536;
	wire [14-1:0] node3539;
	wire [14-1:0] node3540;
	wire [14-1:0] node3541;
	wire [14-1:0] node3542;
	wire [14-1:0] node3543;
	wire [14-1:0] node3544;
	wire [14-1:0] node3547;
	wire [14-1:0] node3550;
	wire [14-1:0] node3551;
	wire [14-1:0] node3554;
	wire [14-1:0] node3557;
	wire [14-1:0] node3558;
	wire [14-1:0] node3560;
	wire [14-1:0] node3563;
	wire [14-1:0] node3566;
	wire [14-1:0] node3567;
	wire [14-1:0] node3568;
	wire [14-1:0] node3571;
	wire [14-1:0] node3574;
	wire [14-1:0] node3576;
	wire [14-1:0] node3577;
	wire [14-1:0] node3580;
	wire [14-1:0] node3583;
	wire [14-1:0] node3584;
	wire [14-1:0] node3585;
	wire [14-1:0] node3586;
	wire [14-1:0] node3590;
	wire [14-1:0] node3591;
	wire [14-1:0] node3592;
	wire [14-1:0] node3595;
	wire [14-1:0] node3599;
	wire [14-1:0] node3600;
	wire [14-1:0] node3601;
	wire [14-1:0] node3602;
	wire [14-1:0] node3605;
	wire [14-1:0] node3608;
	wire [14-1:0] node3610;
	wire [14-1:0] node3613;
	wire [14-1:0] node3614;
	wire [14-1:0] node3616;
	wire [14-1:0] node3619;
	wire [14-1:0] node3620;
	wire [14-1:0] node3623;
	wire [14-1:0] node3626;
	wire [14-1:0] node3627;
	wire [14-1:0] node3628;
	wire [14-1:0] node3629;
	wire [14-1:0] node3630;
	wire [14-1:0] node3631;
	wire [14-1:0] node3632;
	wire [14-1:0] node3633;
	wire [14-1:0] node3636;
	wire [14-1:0] node3639;
	wire [14-1:0] node3640;
	wire [14-1:0] node3644;
	wire [14-1:0] node3645;
	wire [14-1:0] node3648;
	wire [14-1:0] node3649;
	wire [14-1:0] node3653;
	wire [14-1:0] node3654;
	wire [14-1:0] node3655;
	wire [14-1:0] node3656;
	wire [14-1:0] node3659;
	wire [14-1:0] node3662;
	wire [14-1:0] node3663;
	wire [14-1:0] node3667;
	wire [14-1:0] node3668;
	wire [14-1:0] node3669;
	wire [14-1:0] node3672;
	wire [14-1:0] node3675;
	wire [14-1:0] node3678;
	wire [14-1:0] node3679;
	wire [14-1:0] node3680;
	wire [14-1:0] node3681;
	wire [14-1:0] node3682;
	wire [14-1:0] node3685;
	wire [14-1:0] node3688;
	wire [14-1:0] node3689;
	wire [14-1:0] node3693;
	wire [14-1:0] node3694;
	wire [14-1:0] node3697;
	wire [14-1:0] node3700;
	wire [14-1:0] node3701;
	wire [14-1:0] node3702;
	wire [14-1:0] node3703;
	wire [14-1:0] node3706;
	wire [14-1:0] node3709;
	wire [14-1:0] node3710;
	wire [14-1:0] node3713;
	wire [14-1:0] node3716;
	wire [14-1:0] node3717;
	wire [14-1:0] node3718;
	wire [14-1:0] node3723;
	wire [14-1:0] node3724;
	wire [14-1:0] node3725;
	wire [14-1:0] node3726;
	wire [14-1:0] node3727;
	wire [14-1:0] node3728;
	wire [14-1:0] node3731;
	wire [14-1:0] node3734;
	wire [14-1:0] node3735;
	wire [14-1:0] node3739;
	wire [14-1:0] node3740;
	wire [14-1:0] node3741;
	wire [14-1:0] node3744;
	wire [14-1:0] node3747;
	wire [14-1:0] node3750;
	wire [14-1:0] node3751;
	wire [14-1:0] node3752;
	wire [14-1:0] node3753;
	wire [14-1:0] node3757;
	wire [14-1:0] node3758;
	wire [14-1:0] node3762;
	wire [14-1:0] node3763;
	wire [14-1:0] node3764;
	wire [14-1:0] node3767;
	wire [14-1:0] node3770;
	wire [14-1:0] node3771;
	wire [14-1:0] node3774;
	wire [14-1:0] node3777;
	wire [14-1:0] node3778;
	wire [14-1:0] node3779;
	wire [14-1:0] node3780;
	wire [14-1:0] node3781;
	wire [14-1:0] node3785;
	wire [14-1:0] node3786;
	wire [14-1:0] node3789;
	wire [14-1:0] node3792;
	wire [14-1:0] node3794;
	wire [14-1:0] node3796;
	wire [14-1:0] node3799;
	wire [14-1:0] node3800;
	wire [14-1:0] node3801;
	wire [14-1:0] node3802;
	wire [14-1:0] node3805;
	wire [14-1:0] node3808;
	wire [14-1:0] node3810;
	wire [14-1:0] node3813;
	wire [14-1:0] node3815;
	wire [14-1:0] node3816;
	wire [14-1:0] node3819;
	wire [14-1:0] node3822;
	wire [14-1:0] node3823;
	wire [14-1:0] node3824;
	wire [14-1:0] node3825;
	wire [14-1:0] node3826;
	wire [14-1:0] node3827;
	wire [14-1:0] node3828;
	wire [14-1:0] node3832;
	wire [14-1:0] node3833;
	wire [14-1:0] node3836;
	wire [14-1:0] node3839;
	wire [14-1:0] node3840;
	wire [14-1:0] node3842;
	wire [14-1:0] node3845;
	wire [14-1:0] node3846;
	wire [14-1:0] node3849;
	wire [14-1:0] node3852;
	wire [14-1:0] node3853;
	wire [14-1:0] node3854;
	wire [14-1:0] node3855;
	wire [14-1:0] node3859;
	wire [14-1:0] node3860;
	wire [14-1:0] node3864;
	wire [14-1:0] node3866;
	wire [14-1:0] node3867;
	wire [14-1:0] node3870;
	wire [14-1:0] node3873;
	wire [14-1:0] node3874;
	wire [14-1:0] node3875;
	wire [14-1:0] node3876;
	wire [14-1:0] node3878;
	wire [14-1:0] node3881;
	wire [14-1:0] node3883;
	wire [14-1:0] node3886;
	wire [14-1:0] node3887;
	wire [14-1:0] node3889;
	wire [14-1:0] node3892;
	wire [14-1:0] node3893;
	wire [14-1:0] node3896;
	wire [14-1:0] node3899;
	wire [14-1:0] node3900;
	wire [14-1:0] node3901;
	wire [14-1:0] node3902;
	wire [14-1:0] node3906;
	wire [14-1:0] node3907;
	wire [14-1:0] node3911;
	wire [14-1:0] node3912;
	wire [14-1:0] node3913;
	wire [14-1:0] node3917;
	wire [14-1:0] node3918;
	wire [14-1:0] node3921;
	wire [14-1:0] node3924;
	wire [14-1:0] node3925;
	wire [14-1:0] node3926;
	wire [14-1:0] node3927;
	wire [14-1:0] node3928;
	wire [14-1:0] node3930;
	wire [14-1:0] node3933;
	wire [14-1:0] node3935;
	wire [14-1:0] node3938;
	wire [14-1:0] node3939;
	wire [14-1:0] node3941;
	wire [14-1:0] node3944;
	wire [14-1:0] node3945;
	wire [14-1:0] node3949;
	wire [14-1:0] node3950;
	wire [14-1:0] node3951;
	wire [14-1:0] node3952;
	wire [14-1:0] node3955;
	wire [14-1:0] node3958;
	wire [14-1:0] node3959;
	wire [14-1:0] node3963;
	wire [14-1:0] node3964;
	wire [14-1:0] node3965;
	wire [14-1:0] node3968;
	wire [14-1:0] node3971;
	wire [14-1:0] node3972;
	wire [14-1:0] node3975;
	wire [14-1:0] node3978;
	wire [14-1:0] node3979;
	wire [14-1:0] node3980;
	wire [14-1:0] node3981;
	wire [14-1:0] node3983;
	wire [14-1:0] node3986;
	wire [14-1:0] node3987;
	wire [14-1:0] node3990;
	wire [14-1:0] node3993;
	wire [14-1:0] node3994;
	wire [14-1:0] node3995;
	wire [14-1:0] node3999;
	wire [14-1:0] node4002;
	wire [14-1:0] node4003;
	wire [14-1:0] node4004;
	wire [14-1:0] node4006;
	wire [14-1:0] node4009;
	wire [14-1:0] node4010;
	wire [14-1:0] node4013;
	wire [14-1:0] node4016;
	wire [14-1:0] node4017;
	wire [14-1:0] node4018;
	wire [14-1:0] node4022;
	wire [14-1:0] node4023;
	wire [14-1:0] node4026;
	wire [14-1:0] node4029;
	wire [14-1:0] node4030;
	wire [14-1:0] node4031;
	wire [14-1:0] node4032;
	wire [14-1:0] node4033;
	wire [14-1:0] node4034;
	wire [14-1:0] node4035;
	wire [14-1:0] node4036;
	wire [14-1:0] node4037;
	wire [14-1:0] node4040;
	wire [14-1:0] node4043;
	wire [14-1:0] node4046;
	wire [14-1:0] node4047;
	wire [14-1:0] node4048;
	wire [14-1:0] node4051;
	wire [14-1:0] node4054;
	wire [14-1:0] node4055;
	wire [14-1:0] node4058;
	wire [14-1:0] node4061;
	wire [14-1:0] node4062;
	wire [14-1:0] node4063;
	wire [14-1:0] node4064;
	wire [14-1:0] node4068;
	wire [14-1:0] node4069;
	wire [14-1:0] node4072;
	wire [14-1:0] node4075;
	wire [14-1:0] node4076;
	wire [14-1:0] node4079;
	wire [14-1:0] node4080;
	wire [14-1:0] node4083;
	wire [14-1:0] node4086;
	wire [14-1:0] node4087;
	wire [14-1:0] node4088;
	wire [14-1:0] node4089;
	wire [14-1:0] node4090;
	wire [14-1:0] node4093;
	wire [14-1:0] node4096;
	wire [14-1:0] node4097;
	wire [14-1:0] node4100;
	wire [14-1:0] node4103;
	wire [14-1:0] node4104;
	wire [14-1:0] node4106;
	wire [14-1:0] node4109;
	wire [14-1:0] node4110;
	wire [14-1:0] node4114;
	wire [14-1:0] node4115;
	wire [14-1:0] node4116;
	wire [14-1:0] node4117;
	wire [14-1:0] node4121;
	wire [14-1:0] node4124;
	wire [14-1:0] node4125;
	wire [14-1:0] node4126;
	wire [14-1:0] node4129;
	wire [14-1:0] node4132;
	wire [14-1:0] node4134;
	wire [14-1:0] node4137;
	wire [14-1:0] node4138;
	wire [14-1:0] node4139;
	wire [14-1:0] node4140;
	wire [14-1:0] node4141;
	wire [14-1:0] node4142;
	wire [14-1:0] node4146;
	wire [14-1:0] node4147;
	wire [14-1:0] node4150;
	wire [14-1:0] node4153;
	wire [14-1:0] node4154;
	wire [14-1:0] node4155;
	wire [14-1:0] node4158;
	wire [14-1:0] node4161;
	wire [14-1:0] node4162;
	wire [14-1:0] node4165;
	wire [14-1:0] node4168;
	wire [14-1:0] node4169;
	wire [14-1:0] node4170;
	wire [14-1:0] node4171;
	wire [14-1:0] node4174;
	wire [14-1:0] node4177;
	wire [14-1:0] node4178;
	wire [14-1:0] node4181;
	wire [14-1:0] node4184;
	wire [14-1:0] node4185;
	wire [14-1:0] node4186;
	wire [14-1:0] node4189;
	wire [14-1:0] node4192;
	wire [14-1:0] node4193;
	wire [14-1:0] node4196;
	wire [14-1:0] node4199;
	wire [14-1:0] node4200;
	wire [14-1:0] node4201;
	wire [14-1:0] node4202;
	wire [14-1:0] node4203;
	wire [14-1:0] node4206;
	wire [14-1:0] node4209;
	wire [14-1:0] node4210;
	wire [14-1:0] node4213;
	wire [14-1:0] node4216;
	wire [14-1:0] node4217;
	wire [14-1:0] node4218;
	wire [14-1:0] node4221;
	wire [14-1:0] node4224;
	wire [14-1:0] node4225;
	wire [14-1:0] node4228;
	wire [14-1:0] node4231;
	wire [14-1:0] node4232;
	wire [14-1:0] node4233;
	wire [14-1:0] node4236;
	wire [14-1:0] node4238;
	wire [14-1:0] node4241;
	wire [14-1:0] node4242;
	wire [14-1:0] node4245;
	wire [14-1:0] node4246;
	wire [14-1:0] node4249;
	wire [14-1:0] node4252;
	wire [14-1:0] node4253;
	wire [14-1:0] node4254;
	wire [14-1:0] node4255;
	wire [14-1:0] node4256;
	wire [14-1:0] node4257;
	wire [14-1:0] node4258;
	wire [14-1:0] node4262;
	wire [14-1:0] node4263;
	wire [14-1:0] node4266;
	wire [14-1:0] node4269;
	wire [14-1:0] node4270;
	wire [14-1:0] node4272;
	wire [14-1:0] node4275;
	wire [14-1:0] node4278;
	wire [14-1:0] node4279;
	wire [14-1:0] node4280;
	wire [14-1:0] node4281;
	wire [14-1:0] node4284;
	wire [14-1:0] node4287;
	wire [14-1:0] node4288;
	wire [14-1:0] node4291;
	wire [14-1:0] node4294;
	wire [14-1:0] node4295;
	wire [14-1:0] node4297;
	wire [14-1:0] node4300;
	wire [14-1:0] node4302;
	wire [14-1:0] node4305;
	wire [14-1:0] node4306;
	wire [14-1:0] node4307;
	wire [14-1:0] node4309;
	wire [14-1:0] node4310;
	wire [14-1:0] node4314;
	wire [14-1:0] node4315;
	wire [14-1:0] node4318;
	wire [14-1:0] node4319;
	wire [14-1:0] node4322;
	wire [14-1:0] node4325;
	wire [14-1:0] node4326;
	wire [14-1:0] node4327;
	wire [14-1:0] node4328;
	wire [14-1:0] node4331;
	wire [14-1:0] node4334;
	wire [14-1:0] node4336;
	wire [14-1:0] node4339;
	wire [14-1:0] node4340;
	wire [14-1:0] node4341;
	wire [14-1:0] node4344;
	wire [14-1:0] node4347;
	wire [14-1:0] node4348;
	wire [14-1:0] node4351;
	wire [14-1:0] node4354;
	wire [14-1:0] node4355;
	wire [14-1:0] node4356;
	wire [14-1:0] node4357;
	wire [14-1:0] node4358;
	wire [14-1:0] node4361;
	wire [14-1:0] node4363;
	wire [14-1:0] node4366;
	wire [14-1:0] node4367;
	wire [14-1:0] node4369;
	wire [14-1:0] node4372;
	wire [14-1:0] node4373;
	wire [14-1:0] node4376;
	wire [14-1:0] node4379;
	wire [14-1:0] node4380;
	wire [14-1:0] node4381;
	wire [14-1:0] node4382;
	wire [14-1:0] node4385;
	wire [14-1:0] node4388;
	wire [14-1:0] node4389;
	wire [14-1:0] node4392;
	wire [14-1:0] node4395;
	wire [14-1:0] node4396;
	wire [14-1:0] node4397;
	wire [14-1:0] node4400;
	wire [14-1:0] node4403;
	wire [14-1:0] node4405;
	wire [14-1:0] node4408;
	wire [14-1:0] node4409;
	wire [14-1:0] node4410;
	wire [14-1:0] node4411;
	wire [14-1:0] node4413;
	wire [14-1:0] node4416;
	wire [14-1:0] node4417;
	wire [14-1:0] node4420;
	wire [14-1:0] node4423;
	wire [14-1:0] node4424;
	wire [14-1:0] node4426;
	wire [14-1:0] node4429;
	wire [14-1:0] node4432;
	wire [14-1:0] node4433;
	wire [14-1:0] node4434;
	wire [14-1:0] node4435;
	wire [14-1:0] node4440;
	wire [14-1:0] node4441;
	wire [14-1:0] node4442;
	wire [14-1:0] node4445;
	wire [14-1:0] node4448;
	wire [14-1:0] node4449;
	wire [14-1:0] node4452;
	wire [14-1:0] node4455;
	wire [14-1:0] node4456;
	wire [14-1:0] node4457;
	wire [14-1:0] node4458;
	wire [14-1:0] node4459;
	wire [14-1:0] node4460;
	wire [14-1:0] node4461;
	wire [14-1:0] node4462;
	wire [14-1:0] node4465;
	wire [14-1:0] node4468;
	wire [14-1:0] node4469;
	wire [14-1:0] node4473;
	wire [14-1:0] node4474;
	wire [14-1:0] node4475;
	wire [14-1:0] node4478;
	wire [14-1:0] node4482;
	wire [14-1:0] node4483;
	wire [14-1:0] node4484;
	wire [14-1:0] node4485;
	wire [14-1:0] node4488;
	wire [14-1:0] node4491;
	wire [14-1:0] node4492;
	wire [14-1:0] node4495;
	wire [14-1:0] node4498;
	wire [14-1:0] node4499;
	wire [14-1:0] node4501;
	wire [14-1:0] node4504;
	wire [14-1:0] node4505;
	wire [14-1:0] node4508;
	wire [14-1:0] node4511;
	wire [14-1:0] node4512;
	wire [14-1:0] node4513;
	wire [14-1:0] node4514;
	wire [14-1:0] node4515;
	wire [14-1:0] node4518;
	wire [14-1:0] node4522;
	wire [14-1:0] node4523;
	wire [14-1:0] node4524;
	wire [14-1:0] node4527;
	wire [14-1:0] node4530;
	wire [14-1:0] node4531;
	wire [14-1:0] node4534;
	wire [14-1:0] node4537;
	wire [14-1:0] node4538;
	wire [14-1:0] node4539;
	wire [14-1:0] node4540;
	wire [14-1:0] node4543;
	wire [14-1:0] node4546;
	wire [14-1:0] node4547;
	wire [14-1:0] node4550;
	wire [14-1:0] node4553;
	wire [14-1:0] node4554;
	wire [14-1:0] node4555;
	wire [14-1:0] node4558;
	wire [14-1:0] node4561;
	wire [14-1:0] node4563;
	wire [14-1:0] node4566;
	wire [14-1:0] node4567;
	wire [14-1:0] node4568;
	wire [14-1:0] node4569;
	wire [14-1:0] node4570;
	wire [14-1:0] node4572;
	wire [14-1:0] node4575;
	wire [14-1:0] node4576;
	wire [14-1:0] node4579;
	wire [14-1:0] node4582;
	wire [14-1:0] node4583;
	wire [14-1:0] node4586;
	wire [14-1:0] node4587;
	wire [14-1:0] node4591;
	wire [14-1:0] node4592;
	wire [14-1:0] node4593;
	wire [14-1:0] node4596;
	wire [14-1:0] node4597;
	wire [14-1:0] node4601;
	wire [14-1:0] node4602;
	wire [14-1:0] node4604;
	wire [14-1:0] node4607;
	wire [14-1:0] node4609;
	wire [14-1:0] node4612;
	wire [14-1:0] node4613;
	wire [14-1:0] node4614;
	wire [14-1:0] node4615;
	wire [14-1:0] node4616;
	wire [14-1:0] node4619;
	wire [14-1:0] node4622;
	wire [14-1:0] node4623;
	wire [14-1:0] node4626;
	wire [14-1:0] node4629;
	wire [14-1:0] node4630;
	wire [14-1:0] node4631;
	wire [14-1:0] node4634;
	wire [14-1:0] node4637;
	wire [14-1:0] node4638;
	wire [14-1:0] node4641;
	wire [14-1:0] node4644;
	wire [14-1:0] node4645;
	wire [14-1:0] node4646;
	wire [14-1:0] node4647;
	wire [14-1:0] node4650;
	wire [14-1:0] node4653;
	wire [14-1:0] node4654;
	wire [14-1:0] node4657;
	wire [14-1:0] node4660;
	wire [14-1:0] node4661;
	wire [14-1:0] node4663;
	wire [14-1:0] node4666;
	wire [14-1:0] node4667;
	wire [14-1:0] node4670;
	wire [14-1:0] node4673;
	wire [14-1:0] node4674;
	wire [14-1:0] node4675;
	wire [14-1:0] node4676;
	wire [14-1:0] node4677;
	wire [14-1:0] node4678;
	wire [14-1:0] node4681;
	wire [14-1:0] node4682;
	wire [14-1:0] node4685;
	wire [14-1:0] node4688;
	wire [14-1:0] node4689;
	wire [14-1:0] node4690;
	wire [14-1:0] node4693;
	wire [14-1:0] node4696;
	wire [14-1:0] node4697;
	wire [14-1:0] node4701;
	wire [14-1:0] node4702;
	wire [14-1:0] node4703;
	wire [14-1:0] node4704;
	wire [14-1:0] node4707;
	wire [14-1:0] node4710;
	wire [14-1:0] node4711;
	wire [14-1:0] node4714;
	wire [14-1:0] node4717;
	wire [14-1:0] node4719;
	wire [14-1:0] node4720;
	wire [14-1:0] node4723;
	wire [14-1:0] node4726;
	wire [14-1:0] node4727;
	wire [14-1:0] node4728;
	wire [14-1:0] node4729;
	wire [14-1:0] node4730;
	wire [14-1:0] node4734;
	wire [14-1:0] node4736;
	wire [14-1:0] node4739;
	wire [14-1:0] node4740;
	wire [14-1:0] node4741;
	wire [14-1:0] node4744;
	wire [14-1:0] node4747;
	wire [14-1:0] node4748;
	wire [14-1:0] node4751;
	wire [14-1:0] node4754;
	wire [14-1:0] node4755;
	wire [14-1:0] node4756;
	wire [14-1:0] node4757;
	wire [14-1:0] node4760;
	wire [14-1:0] node4763;
	wire [14-1:0] node4764;
	wire [14-1:0] node4767;
	wire [14-1:0] node4770;
	wire [14-1:0] node4771;
	wire [14-1:0] node4772;
	wire [14-1:0] node4775;
	wire [14-1:0] node4778;
	wire [14-1:0] node4781;
	wire [14-1:0] node4782;
	wire [14-1:0] node4783;
	wire [14-1:0] node4784;
	wire [14-1:0] node4785;
	wire [14-1:0] node4788;
	wire [14-1:0] node4790;
	wire [14-1:0] node4793;
	wire [14-1:0] node4794;
	wire [14-1:0] node4795;
	wire [14-1:0] node4798;
	wire [14-1:0] node4801;
	wire [14-1:0] node4803;
	wire [14-1:0] node4806;
	wire [14-1:0] node4807;
	wire [14-1:0] node4808;
	wire [14-1:0] node4810;
	wire [14-1:0] node4813;
	wire [14-1:0] node4816;
	wire [14-1:0] node4817;
	wire [14-1:0] node4819;
	wire [14-1:0] node4822;
	wire [14-1:0] node4823;
	wire [14-1:0] node4826;
	wire [14-1:0] node4829;
	wire [14-1:0] node4830;
	wire [14-1:0] node4831;
	wire [14-1:0] node4832;
	wire [14-1:0] node4833;
	wire [14-1:0] node4836;
	wire [14-1:0] node4839;
	wire [14-1:0] node4840;
	wire [14-1:0] node4843;
	wire [14-1:0] node4846;
	wire [14-1:0] node4847;
	wire [14-1:0] node4848;
	wire [14-1:0] node4852;
	wire [14-1:0] node4853;
	wire [14-1:0] node4856;
	wire [14-1:0] node4859;
	wire [14-1:0] node4860;
	wire [14-1:0] node4861;
	wire [14-1:0] node4863;
	wire [14-1:0] node4866;
	wire [14-1:0] node4867;
	wire [14-1:0] node4870;
	wire [14-1:0] node4873;
	wire [14-1:0] node4874;
	wire [14-1:0] node4876;
	wire [14-1:0] node4879;
	wire [14-1:0] node4880;
	wire [14-1:0] node4883;
	wire [14-1:0] node4886;
	wire [14-1:0] node4887;
	wire [14-1:0] node4888;
	wire [14-1:0] node4889;
	wire [14-1:0] node4890;
	wire [14-1:0] node4891;
	wire [14-1:0] node4892;
	wire [14-1:0] node4893;
	wire [14-1:0] node4894;
	wire [14-1:0] node4895;
	wire [14-1:0] node4899;
	wire [14-1:0] node4900;
	wire [14-1:0] node4903;
	wire [14-1:0] node4906;
	wire [14-1:0] node4907;
	wire [14-1:0] node4908;
	wire [14-1:0] node4911;
	wire [14-1:0] node4915;
	wire [14-1:0] node4916;
	wire [14-1:0] node4917;
	wire [14-1:0] node4918;
	wire [14-1:0] node4922;
	wire [14-1:0] node4923;
	wire [14-1:0] node4926;
	wire [14-1:0] node4929;
	wire [14-1:0] node4930;
	wire [14-1:0] node4933;
	wire [14-1:0] node4934;
	wire [14-1:0] node4937;
	wire [14-1:0] node4940;
	wire [14-1:0] node4941;
	wire [14-1:0] node4942;
	wire [14-1:0] node4943;
	wire [14-1:0] node4944;
	wire [14-1:0] node4948;
	wire [14-1:0] node4949;
	wire [14-1:0] node4953;
	wire [14-1:0] node4954;
	wire [14-1:0] node4956;
	wire [14-1:0] node4959;
	wire [14-1:0] node4960;
	wire [14-1:0] node4963;
	wire [14-1:0] node4966;
	wire [14-1:0] node4967;
	wire [14-1:0] node4968;
	wire [14-1:0] node4970;
	wire [14-1:0] node4973;
	wire [14-1:0] node4974;
	wire [14-1:0] node4977;
	wire [14-1:0] node4980;
	wire [14-1:0] node4981;
	wire [14-1:0] node4982;
	wire [14-1:0] node4985;
	wire [14-1:0] node4988;
	wire [14-1:0] node4989;
	wire [14-1:0] node4992;
	wire [14-1:0] node4995;
	wire [14-1:0] node4996;
	wire [14-1:0] node4997;
	wire [14-1:0] node4998;
	wire [14-1:0] node4999;
	wire [14-1:0] node5000;
	wire [14-1:0] node5003;
	wire [14-1:0] node5006;
	wire [14-1:0] node5007;
	wire [14-1:0] node5011;
	wire [14-1:0] node5012;
	wire [14-1:0] node5014;
	wire [14-1:0] node5017;
	wire [14-1:0] node5019;
	wire [14-1:0] node5022;
	wire [14-1:0] node5023;
	wire [14-1:0] node5024;
	wire [14-1:0] node5025;
	wire [14-1:0] node5028;
	wire [14-1:0] node5031;
	wire [14-1:0] node5032;
	wire [14-1:0] node5035;
	wire [14-1:0] node5038;
	wire [14-1:0] node5039;
	wire [14-1:0] node5040;
	wire [14-1:0] node5043;
	wire [14-1:0] node5046;
	wire [14-1:0] node5047;
	wire [14-1:0] node5051;
	wire [14-1:0] node5052;
	wire [14-1:0] node5053;
	wire [14-1:0] node5054;
	wire [14-1:0] node5055;
	wire [14-1:0] node5058;
	wire [14-1:0] node5061;
	wire [14-1:0] node5062;
	wire [14-1:0] node5066;
	wire [14-1:0] node5067;
	wire [14-1:0] node5069;
	wire [14-1:0] node5072;
	wire [14-1:0] node5074;
	wire [14-1:0] node5077;
	wire [14-1:0] node5078;
	wire [14-1:0] node5079;
	wire [14-1:0] node5081;
	wire [14-1:0] node5084;
	wire [14-1:0] node5085;
	wire [14-1:0] node5088;
	wire [14-1:0] node5091;
	wire [14-1:0] node5092;
	wire [14-1:0] node5093;
	wire [14-1:0] node5097;
	wire [14-1:0] node5098;
	wire [14-1:0] node5101;
	wire [14-1:0] node5104;
	wire [14-1:0] node5105;
	wire [14-1:0] node5106;
	wire [14-1:0] node5107;
	wire [14-1:0] node5108;
	wire [14-1:0] node5109;
	wire [14-1:0] node5112;
	wire [14-1:0] node5113;
	wire [14-1:0] node5116;
	wire [14-1:0] node5119;
	wire [14-1:0] node5120;
	wire [14-1:0] node5122;
	wire [14-1:0] node5125;
	wire [14-1:0] node5128;
	wire [14-1:0] node5129;
	wire [14-1:0] node5130;
	wire [14-1:0] node5132;
	wire [14-1:0] node5135;
	wire [14-1:0] node5136;
	wire [14-1:0] node5139;
	wire [14-1:0] node5142;
	wire [14-1:0] node5143;
	wire [14-1:0] node5145;
	wire [14-1:0] node5148;
	wire [14-1:0] node5149;
	wire [14-1:0] node5152;
	wire [14-1:0] node5155;
	wire [14-1:0] node5156;
	wire [14-1:0] node5157;
	wire [14-1:0] node5158;
	wire [14-1:0] node5159;
	wire [14-1:0] node5163;
	wire [14-1:0] node5165;
	wire [14-1:0] node5168;
	wire [14-1:0] node5169;
	wire [14-1:0] node5170;
	wire [14-1:0] node5174;
	wire [14-1:0] node5175;
	wire [14-1:0] node5178;
	wire [14-1:0] node5181;
	wire [14-1:0] node5182;
	wire [14-1:0] node5183;
	wire [14-1:0] node5184;
	wire [14-1:0] node5189;
	wire [14-1:0] node5190;
	wire [14-1:0] node5191;
	wire [14-1:0] node5194;
	wire [14-1:0] node5198;
	wire [14-1:0] node5199;
	wire [14-1:0] node5200;
	wire [14-1:0] node5201;
	wire [14-1:0] node5202;
	wire [14-1:0] node5203;
	wire [14-1:0] node5206;
	wire [14-1:0] node5209;
	wire [14-1:0] node5212;
	wire [14-1:0] node5215;
	wire [14-1:0] node5216;
	wire [14-1:0] node5218;
	wire [14-1:0] node5219;
	wire [14-1:0] node5222;
	wire [14-1:0] node5225;
	wire [14-1:0] node5226;
	wire [14-1:0] node5227;
	wire [14-1:0] node5230;
	wire [14-1:0] node5233;
	wire [14-1:0] node5234;
	wire [14-1:0] node5238;
	wire [14-1:0] node5239;
	wire [14-1:0] node5240;
	wire [14-1:0] node5241;
	wire [14-1:0] node5243;
	wire [14-1:0] node5246;
	wire [14-1:0] node5247;
	wire [14-1:0] node5251;
	wire [14-1:0] node5252;
	wire [14-1:0] node5253;
	wire [14-1:0] node5257;
	wire [14-1:0] node5258;
	wire [14-1:0] node5261;
	wire [14-1:0] node5264;
	wire [14-1:0] node5265;
	wire [14-1:0] node5266;
	wire [14-1:0] node5267;
	wire [14-1:0] node5271;
	wire [14-1:0] node5273;
	wire [14-1:0] node5276;
	wire [14-1:0] node5277;
	wire [14-1:0] node5281;
	wire [14-1:0] node5282;
	wire [14-1:0] node5283;
	wire [14-1:0] node5284;
	wire [14-1:0] node5285;
	wire [14-1:0] node5286;
	wire [14-1:0] node5287;
	wire [14-1:0] node5288;
	wire [14-1:0] node5291;
	wire [14-1:0] node5294;
	wire [14-1:0] node5295;
	wire [14-1:0] node5298;
	wire [14-1:0] node5301;
	wire [14-1:0] node5302;
	wire [14-1:0] node5303;
	wire [14-1:0] node5306;
	wire [14-1:0] node5309;
	wire [14-1:0] node5311;
	wire [14-1:0] node5314;
	wire [14-1:0] node5315;
	wire [14-1:0] node5316;
	wire [14-1:0] node5319;
	wire [14-1:0] node5320;
	wire [14-1:0] node5324;
	wire [14-1:0] node5325;
	wire [14-1:0] node5326;
	wire [14-1:0] node5330;
	wire [14-1:0] node5331;
	wire [14-1:0] node5334;
	wire [14-1:0] node5337;
	wire [14-1:0] node5338;
	wire [14-1:0] node5339;
	wire [14-1:0] node5340;
	wire [14-1:0] node5341;
	wire [14-1:0] node5344;
	wire [14-1:0] node5347;
	wire [14-1:0] node5348;
	wire [14-1:0] node5352;
	wire [14-1:0] node5354;
	wire [14-1:0] node5355;
	wire [14-1:0] node5358;
	wire [14-1:0] node5361;
	wire [14-1:0] node5362;
	wire [14-1:0] node5363;
	wire [14-1:0] node5364;
	wire [14-1:0] node5367;
	wire [14-1:0] node5370;
	wire [14-1:0] node5372;
	wire [14-1:0] node5375;
	wire [14-1:0] node5376;
	wire [14-1:0] node5377;
	wire [14-1:0] node5380;
	wire [14-1:0] node5383;
	wire [14-1:0] node5385;
	wire [14-1:0] node5388;
	wire [14-1:0] node5389;
	wire [14-1:0] node5390;
	wire [14-1:0] node5391;
	wire [14-1:0] node5392;
	wire [14-1:0] node5393;
	wire [14-1:0] node5396;
	wire [14-1:0] node5399;
	wire [14-1:0] node5402;
	wire [14-1:0] node5404;
	wire [14-1:0] node5405;
	wire [14-1:0] node5409;
	wire [14-1:0] node5410;
	wire [14-1:0] node5411;
	wire [14-1:0] node5413;
	wire [14-1:0] node5416;
	wire [14-1:0] node5418;
	wire [14-1:0] node5421;
	wire [14-1:0] node5422;
	wire [14-1:0] node5423;
	wire [14-1:0] node5427;
	wire [14-1:0] node5429;
	wire [14-1:0] node5432;
	wire [14-1:0] node5433;
	wire [14-1:0] node5434;
	wire [14-1:0] node5435;
	wire [14-1:0] node5438;
	wire [14-1:0] node5439;
	wire [14-1:0] node5442;
	wire [14-1:0] node5445;
	wire [14-1:0] node5446;
	wire [14-1:0] node5449;
	wire [14-1:0] node5451;
	wire [14-1:0] node5454;
	wire [14-1:0] node5455;
	wire [14-1:0] node5456;
	wire [14-1:0] node5458;
	wire [14-1:0] node5461;
	wire [14-1:0] node5462;
	wire [14-1:0] node5465;
	wire [14-1:0] node5468;
	wire [14-1:0] node5469;
	wire [14-1:0] node5471;
	wire [14-1:0] node5474;
	wire [14-1:0] node5475;
	wire [14-1:0] node5479;
	wire [14-1:0] node5480;
	wire [14-1:0] node5481;
	wire [14-1:0] node5482;
	wire [14-1:0] node5483;
	wire [14-1:0] node5484;
	wire [14-1:0] node5487;
	wire [14-1:0] node5488;
	wire [14-1:0] node5491;
	wire [14-1:0] node5494;
	wire [14-1:0] node5495;
	wire [14-1:0] node5496;
	wire [14-1:0] node5499;
	wire [14-1:0] node5502;
	wire [14-1:0] node5503;
	wire [14-1:0] node5507;
	wire [14-1:0] node5508;
	wire [14-1:0] node5509;
	wire [14-1:0] node5510;
	wire [14-1:0] node5513;
	wire [14-1:0] node5516;
	wire [14-1:0] node5517;
	wire [14-1:0] node5520;
	wire [14-1:0] node5523;
	wire [14-1:0] node5524;
	wire [14-1:0] node5525;
	wire [14-1:0] node5528;
	wire [14-1:0] node5531;
	wire [14-1:0] node5533;
	wire [14-1:0] node5536;
	wire [14-1:0] node5537;
	wire [14-1:0] node5538;
	wire [14-1:0] node5539;
	wire [14-1:0] node5541;
	wire [14-1:0] node5544;
	wire [14-1:0] node5547;
	wire [14-1:0] node5548;
	wire [14-1:0] node5549;
	wire [14-1:0] node5552;
	wire [14-1:0] node5556;
	wire [14-1:0] node5557;
	wire [14-1:0] node5558;
	wire [14-1:0] node5559;
	wire [14-1:0] node5562;
	wire [14-1:0] node5565;
	wire [14-1:0] node5566;
	wire [14-1:0] node5569;
	wire [14-1:0] node5572;
	wire [14-1:0] node5573;
	wire [14-1:0] node5574;
	wire [14-1:0] node5577;
	wire [14-1:0] node5580;
	wire [14-1:0] node5582;
	wire [14-1:0] node5585;
	wire [14-1:0] node5586;
	wire [14-1:0] node5587;
	wire [14-1:0] node5588;
	wire [14-1:0] node5589;
	wire [14-1:0] node5590;
	wire [14-1:0] node5593;
	wire [14-1:0] node5596;
	wire [14-1:0] node5597;
	wire [14-1:0] node5600;
	wire [14-1:0] node5603;
	wire [14-1:0] node5604;
	wire [14-1:0] node5606;
	wire [14-1:0] node5609;
	wire [14-1:0] node5611;
	wire [14-1:0] node5614;
	wire [14-1:0] node5615;
	wire [14-1:0] node5616;
	wire [14-1:0] node5618;
	wire [14-1:0] node5621;
	wire [14-1:0] node5622;
	wire [14-1:0] node5626;
	wire [14-1:0] node5627;
	wire [14-1:0] node5629;
	wire [14-1:0] node5632;
	wire [14-1:0] node5633;
	wire [14-1:0] node5637;
	wire [14-1:0] node5638;
	wire [14-1:0] node5639;
	wire [14-1:0] node5640;
	wire [14-1:0] node5641;
	wire [14-1:0] node5645;
	wire [14-1:0] node5647;
	wire [14-1:0] node5650;
	wire [14-1:0] node5651;
	wire [14-1:0] node5652;
	wire [14-1:0] node5655;
	wire [14-1:0] node5658;
	wire [14-1:0] node5659;
	wire [14-1:0] node5662;
	wire [14-1:0] node5665;
	wire [14-1:0] node5666;
	wire [14-1:0] node5667;
	wire [14-1:0] node5669;
	wire [14-1:0] node5672;
	wire [14-1:0] node5673;
	wire [14-1:0] node5676;
	wire [14-1:0] node5679;
	wire [14-1:0] node5680;
	wire [14-1:0] node5682;
	wire [14-1:0] node5685;
	wire [14-1:0] node5687;
	wire [14-1:0] node5690;
	wire [14-1:0] node5691;
	wire [14-1:0] node5692;
	wire [14-1:0] node5693;
	wire [14-1:0] node5694;
	wire [14-1:0] node5695;
	wire [14-1:0] node5696;
	wire [14-1:0] node5697;
	wire [14-1:0] node5699;
	wire [14-1:0] node5702;
	wire [14-1:0] node5703;
	wire [14-1:0] node5707;
	wire [14-1:0] node5708;
	wire [14-1:0] node5709;
	wire [14-1:0] node5712;
	wire [14-1:0] node5716;
	wire [14-1:0] node5717;
	wire [14-1:0] node5718;
	wire [14-1:0] node5720;
	wire [14-1:0] node5723;
	wire [14-1:0] node5724;
	wire [14-1:0] node5727;
	wire [14-1:0] node5730;
	wire [14-1:0] node5731;
	wire [14-1:0] node5732;
	wire [14-1:0] node5735;
	wire [14-1:0] node5738;
	wire [14-1:0] node5739;
	wire [14-1:0] node5743;
	wire [14-1:0] node5744;
	wire [14-1:0] node5745;
	wire [14-1:0] node5746;
	wire [14-1:0] node5747;
	wire [14-1:0] node5751;
	wire [14-1:0] node5752;
	wire [14-1:0] node5755;
	wire [14-1:0] node5758;
	wire [14-1:0] node5759;
	wire [14-1:0] node5760;
	wire [14-1:0] node5765;
	wire [14-1:0] node5766;
	wire [14-1:0] node5767;
	wire [14-1:0] node5768;
	wire [14-1:0] node5772;
	wire [14-1:0] node5773;
	wire [14-1:0] node5776;
	wire [14-1:0] node5779;
	wire [14-1:0] node5781;
	wire [14-1:0] node5782;
	wire [14-1:0] node5786;
	wire [14-1:0] node5787;
	wire [14-1:0] node5788;
	wire [14-1:0] node5789;
	wire [14-1:0] node5790;
	wire [14-1:0] node5792;
	wire [14-1:0] node5795;
	wire [14-1:0] node5796;
	wire [14-1:0] node5799;
	wire [14-1:0] node5802;
	wire [14-1:0] node5803;
	wire [14-1:0] node5804;
	wire [14-1:0] node5807;
	wire [14-1:0] node5810;
	wire [14-1:0] node5811;
	wire [14-1:0] node5815;
	wire [14-1:0] node5816;
	wire [14-1:0] node5817;
	wire [14-1:0] node5821;
	wire [14-1:0] node5822;
	wire [14-1:0] node5823;
	wire [14-1:0] node5826;
	wire [14-1:0] node5829;
	wire [14-1:0] node5830;
	wire [14-1:0] node5834;
	wire [14-1:0] node5835;
	wire [14-1:0] node5836;
	wire [14-1:0] node5837;
	wire [14-1:0] node5838;
	wire [14-1:0] node5842;
	wire [14-1:0] node5843;
	wire [14-1:0] node5846;
	wire [14-1:0] node5849;
	wire [14-1:0] node5851;
	wire [14-1:0] node5852;
	wire [14-1:0] node5855;
	wire [14-1:0] node5858;
	wire [14-1:0] node5859;
	wire [14-1:0] node5860;
	wire [14-1:0] node5862;
	wire [14-1:0] node5865;
	wire [14-1:0] node5868;
	wire [14-1:0] node5869;
	wire [14-1:0] node5871;
	wire [14-1:0] node5874;
	wire [14-1:0] node5876;
	wire [14-1:0] node5879;
	wire [14-1:0] node5880;
	wire [14-1:0] node5881;
	wire [14-1:0] node5882;
	wire [14-1:0] node5883;
	wire [14-1:0] node5885;
	wire [14-1:0] node5886;
	wire [14-1:0] node5889;
	wire [14-1:0] node5892;
	wire [14-1:0] node5893;
	wire [14-1:0] node5894;
	wire [14-1:0] node5897;
	wire [14-1:0] node5900;
	wire [14-1:0] node5901;
	wire [14-1:0] node5905;
	wire [14-1:0] node5906;
	wire [14-1:0] node5907;
	wire [14-1:0] node5908;
	wire [14-1:0] node5911;
	wire [14-1:0] node5914;
	wire [14-1:0] node5915;
	wire [14-1:0] node5918;
	wire [14-1:0] node5921;
	wire [14-1:0] node5922;
	wire [14-1:0] node5923;
	wire [14-1:0] node5926;
	wire [14-1:0] node5929;
	wire [14-1:0] node5930;
	wire [14-1:0] node5934;
	wire [14-1:0] node5935;
	wire [14-1:0] node5936;
	wire [14-1:0] node5937;
	wire [14-1:0] node5938;
	wire [14-1:0] node5941;
	wire [14-1:0] node5944;
	wire [14-1:0] node5945;
	wire [14-1:0] node5948;
	wire [14-1:0] node5951;
	wire [14-1:0] node5952;
	wire [14-1:0] node5953;
	wire [14-1:0] node5956;
	wire [14-1:0] node5959;
	wire [14-1:0] node5961;
	wire [14-1:0] node5964;
	wire [14-1:0] node5965;
	wire [14-1:0] node5966;
	wire [14-1:0] node5968;
	wire [14-1:0] node5971;
	wire [14-1:0] node5974;
	wire [14-1:0] node5975;
	wire [14-1:0] node5978;
	wire [14-1:0] node5979;
	wire [14-1:0] node5982;
	wire [14-1:0] node5985;
	wire [14-1:0] node5986;
	wire [14-1:0] node5987;
	wire [14-1:0] node5988;
	wire [14-1:0] node5989;
	wire [14-1:0] node5990;
	wire [14-1:0] node5994;
	wire [14-1:0] node5995;
	wire [14-1:0] node5998;
	wire [14-1:0] node6001;
	wire [14-1:0] node6002;
	wire [14-1:0] node6003;
	wire [14-1:0] node6006;
	wire [14-1:0] node6009;
	wire [14-1:0] node6011;
	wire [14-1:0] node6014;
	wire [14-1:0] node6015;
	wire [14-1:0] node6016;
	wire [14-1:0] node6018;
	wire [14-1:0] node6021;
	wire [14-1:0] node6023;
	wire [14-1:0] node6026;
	wire [14-1:0] node6027;
	wire [14-1:0] node6030;
	wire [14-1:0] node6032;
	wire [14-1:0] node6035;
	wire [14-1:0] node6036;
	wire [14-1:0] node6037;
	wire [14-1:0] node6039;
	wire [14-1:0] node6040;
	wire [14-1:0] node6043;
	wire [14-1:0] node6046;
	wire [14-1:0] node6047;
	wire [14-1:0] node6048;
	wire [14-1:0] node6051;
	wire [14-1:0] node6054;
	wire [14-1:0] node6056;
	wire [14-1:0] node6059;
	wire [14-1:0] node6060;
	wire [14-1:0] node6061;
	wire [14-1:0] node6063;
	wire [14-1:0] node6066;
	wire [14-1:0] node6067;
	wire [14-1:0] node6070;
	wire [14-1:0] node6073;
	wire [14-1:0] node6074;
	wire [14-1:0] node6076;
	wire [14-1:0] node6079;
	wire [14-1:0] node6080;
	wire [14-1:0] node6083;
	wire [14-1:0] node6086;
	wire [14-1:0] node6087;
	wire [14-1:0] node6088;
	wire [14-1:0] node6089;
	wire [14-1:0] node6090;
	wire [14-1:0] node6091;
	wire [14-1:0] node6092;
	wire [14-1:0] node6096;
	wire [14-1:0] node6097;
	wire [14-1:0] node6098;
	wire [14-1:0] node6101;
	wire [14-1:0] node6104;
	wire [14-1:0] node6105;
	wire [14-1:0] node6108;
	wire [14-1:0] node6111;
	wire [14-1:0] node6112;
	wire [14-1:0] node6113;
	wire [14-1:0] node6115;
	wire [14-1:0] node6119;
	wire [14-1:0] node6120;
	wire [14-1:0] node6121;
	wire [14-1:0] node6125;
	wire [14-1:0] node6126;
	wire [14-1:0] node6129;
	wire [14-1:0] node6132;
	wire [14-1:0] node6133;
	wire [14-1:0] node6134;
	wire [14-1:0] node6136;
	wire [14-1:0] node6137;
	wire [14-1:0] node6141;
	wire [14-1:0] node6142;
	wire [14-1:0] node6144;
	wire [14-1:0] node6147;
	wire [14-1:0] node6149;
	wire [14-1:0] node6152;
	wire [14-1:0] node6153;
	wire [14-1:0] node6154;
	wire [14-1:0] node6156;
	wire [14-1:0] node6159;
	wire [14-1:0] node6161;
	wire [14-1:0] node6164;
	wire [14-1:0] node6165;
	wire [14-1:0] node6167;
	wire [14-1:0] node6171;
	wire [14-1:0] node6172;
	wire [14-1:0] node6173;
	wire [14-1:0] node6174;
	wire [14-1:0] node6175;
	wire [14-1:0] node6177;
	wire [14-1:0] node6180;
	wire [14-1:0] node6182;
	wire [14-1:0] node6185;
	wire [14-1:0] node6186;
	wire [14-1:0] node6187;
	wire [14-1:0] node6191;
	wire [14-1:0] node6192;
	wire [14-1:0] node6195;
	wire [14-1:0] node6198;
	wire [14-1:0] node6199;
	wire [14-1:0] node6200;
	wire [14-1:0] node6202;
	wire [14-1:0] node6205;
	wire [14-1:0] node6206;
	wire [14-1:0] node6209;
	wire [14-1:0] node6212;
	wire [14-1:0] node6213;
	wire [14-1:0] node6214;
	wire [14-1:0] node6217;
	wire [14-1:0] node6220;
	wire [14-1:0] node6221;
	wire [14-1:0] node6224;
	wire [14-1:0] node6227;
	wire [14-1:0] node6228;
	wire [14-1:0] node6229;
	wire [14-1:0] node6231;
	wire [14-1:0] node6232;
	wire [14-1:0] node6236;
	wire [14-1:0] node6238;
	wire [14-1:0] node6239;
	wire [14-1:0] node6243;
	wire [14-1:0] node6244;
	wire [14-1:0] node6245;
	wire [14-1:0] node6246;
	wire [14-1:0] node6250;
	wire [14-1:0] node6251;
	wire [14-1:0] node6254;
	wire [14-1:0] node6257;
	wire [14-1:0] node6258;
	wire [14-1:0] node6259;
	wire [14-1:0] node6262;
	wire [14-1:0] node6265;
	wire [14-1:0] node6266;
	wire [14-1:0] node6269;
	wire [14-1:0] node6272;
	wire [14-1:0] node6273;
	wire [14-1:0] node6274;
	wire [14-1:0] node6275;
	wire [14-1:0] node6276;
	wire [14-1:0] node6277;
	wire [14-1:0] node6279;
	wire [14-1:0] node6282;
	wire [14-1:0] node6283;
	wire [14-1:0] node6286;
	wire [14-1:0] node6289;
	wire [14-1:0] node6290;
	wire [14-1:0] node6291;
	wire [14-1:0] node6294;
	wire [14-1:0] node6297;
	wire [14-1:0] node6298;
	wire [14-1:0] node6301;
	wire [14-1:0] node6304;
	wire [14-1:0] node6305;
	wire [14-1:0] node6306;
	wire [14-1:0] node6307;
	wire [14-1:0] node6310;
	wire [14-1:0] node6313;
	wire [14-1:0] node6315;
	wire [14-1:0] node6318;
	wire [14-1:0] node6320;
	wire [14-1:0] node6321;
	wire [14-1:0] node6325;
	wire [14-1:0] node6326;
	wire [14-1:0] node6327;
	wire [14-1:0] node6328;
	wire [14-1:0] node6330;
	wire [14-1:0] node6333;
	wire [14-1:0] node6334;
	wire [14-1:0] node6338;
	wire [14-1:0] node6339;
	wire [14-1:0] node6340;
	wire [14-1:0] node6344;
	wire [14-1:0] node6345;
	wire [14-1:0] node6348;
	wire [14-1:0] node6351;
	wire [14-1:0] node6352;
	wire [14-1:0] node6353;
	wire [14-1:0] node6356;
	wire [14-1:0] node6357;
	wire [14-1:0] node6361;
	wire [14-1:0] node6362;
	wire [14-1:0] node6364;
	wire [14-1:0] node6367;
	wire [14-1:0] node6369;
	wire [14-1:0] node6372;
	wire [14-1:0] node6373;
	wire [14-1:0] node6374;
	wire [14-1:0] node6375;
	wire [14-1:0] node6376;
	wire [14-1:0] node6377;
	wire [14-1:0] node6381;
	wire [14-1:0] node6382;
	wire [14-1:0] node6385;
	wire [14-1:0] node6388;
	wire [14-1:0] node6389;
	wire [14-1:0] node6390;
	wire [14-1:0] node6393;
	wire [14-1:0] node6396;
	wire [14-1:0] node6398;
	wire [14-1:0] node6401;
	wire [14-1:0] node6402;
	wire [14-1:0] node6403;
	wire [14-1:0] node6405;
	wire [14-1:0] node6408;
	wire [14-1:0] node6409;
	wire [14-1:0] node6412;
	wire [14-1:0] node6415;
	wire [14-1:0] node6416;
	wire [14-1:0] node6417;
	wire [14-1:0] node6420;
	wire [14-1:0] node6423;
	wire [14-1:0] node6424;
	wire [14-1:0] node6427;
	wire [14-1:0] node6430;
	wire [14-1:0] node6431;
	wire [14-1:0] node6432;
	wire [14-1:0] node6433;
	wire [14-1:0] node6434;
	wire [14-1:0] node6437;
	wire [14-1:0] node6440;
	wire [14-1:0] node6441;
	wire [14-1:0] node6444;
	wire [14-1:0] node6447;
	wire [14-1:0] node6448;
	wire [14-1:0] node6449;
	wire [14-1:0] node6453;
	wire [14-1:0] node6454;
	wire [14-1:0] node6458;
	wire [14-1:0] node6459;
	wire [14-1:0] node6460;
	wire [14-1:0] node6461;
	wire [14-1:0] node6465;
	wire [14-1:0] node6467;
	wire [14-1:0] node6470;
	wire [14-1:0] node6471;
	wire [14-1:0] node6472;
	wire [14-1:0] node6476;
	wire [14-1:0] node6478;

	assign outp = (inp[5]) ? node3202 : node1;
		assign node1 = (inp[1]) ? node1651 : node2;
			assign node2 = (inp[3]) ? node848 : node3;
				assign node3 = (inp[6]) ? node417 : node4;
					assign node4 = (inp[12]) ? node220 : node5;
						assign node5 = (inp[4]) ? node113 : node6;
							assign node6 = (inp[9]) ? node58 : node7;
								assign node7 = (inp[8]) ? node31 : node8;
									assign node8 = (inp[0]) ? node22 : node9;
										assign node9 = (inp[13]) ? node17 : node10;
											assign node10 = (inp[11]) ? node14 : node11;
												assign node11 = (inp[10]) ? 14'b00111111111111 : 14'b01111111111111;
												assign node14 = (inp[7]) ? 14'b00111111111111 : 14'b00111111111111;
											assign node17 = (inp[7]) ? node19 : 14'b00111111111111;
												assign node19 = (inp[11]) ? 14'b00011111111111 : 14'b00011111111111;
										assign node22 = (inp[11]) ? 14'b00001111111111 : node23;
											assign node23 = (inp[10]) ? node27 : node24;
												assign node24 = (inp[2]) ? 14'b00011111111111 : 14'b00111111111111;
												assign node27 = (inp[13]) ? 14'b00001111111111 : 14'b00011111111111;
									assign node31 = (inp[11]) ? node45 : node32;
										assign node32 = (inp[13]) ? node40 : node33;
											assign node33 = (inp[10]) ? node37 : node34;
												assign node34 = (inp[0]) ? 14'b00011111111111 : 14'b00111111111111;
												assign node37 = (inp[7]) ? 14'b00001111111111 : 14'b00011111111111;
											assign node40 = (inp[10]) ? 14'b00000111111111 : node41;
												assign node41 = (inp[0]) ? 14'b00001111111111 : 14'b00011111111111;
										assign node45 = (inp[2]) ? node53 : node46;
											assign node46 = (inp[7]) ? node50 : node47;
												assign node47 = (inp[10]) ? 14'b00001111111111 : 14'b00011111111111;
												assign node50 = (inp[0]) ? 14'b00000111111111 : 14'b00001111111111;
											assign node53 = (inp[0]) ? 14'b00000011111111 : node54;
												assign node54 = (inp[10]) ? 14'b00000111111111 : 14'b00001111111111;
								assign node58 = (inp[8]) ? node84 : node59;
									assign node59 = (inp[10]) ? node73 : node60;
										assign node60 = (inp[0]) ? node66 : node61;
											assign node61 = (inp[11]) ? 14'b00011111111111 : node62;
												assign node62 = (inp[13]) ? 14'b00011111111111 : 14'b00111111111111;
											assign node66 = (inp[11]) ? node70 : node67;
												assign node67 = (inp[13]) ? 14'b00000111111111 : 14'b00011111111111;
												assign node70 = (inp[2]) ? 14'b00000111111111 : 14'b00001111111111;
										assign node73 = (inp[11]) ? node81 : node74;
											assign node74 = (inp[2]) ? node78 : node75;
												assign node75 = (inp[7]) ? 14'b00001111111111 : 14'b00011111111111;
												assign node78 = (inp[13]) ? 14'b00000111111111 : 14'b00001111111111;
											assign node81 = (inp[2]) ? 14'b00000011111111 : 14'b00000111111111;
									assign node84 = (inp[7]) ? node98 : node85;
										assign node85 = (inp[10]) ? node93 : node86;
											assign node86 = (inp[2]) ? node90 : node87;
												assign node87 = (inp[11]) ? 14'b00001111111111 : 14'b00011111111111;
												assign node90 = (inp[11]) ? 14'b00000111111111 : 14'b00001111111111;
											assign node93 = (inp[11]) ? 14'b00000111111111 : node94;
												assign node94 = (inp[0]) ? 14'b00000111111111 : 14'b00001111111111;
										assign node98 = (inp[11]) ? node106 : node99;
											assign node99 = (inp[13]) ? node103 : node100;
												assign node100 = (inp[0]) ? 14'b00001111111111 : 14'b00011111111111;
												assign node103 = (inp[10]) ? 14'b00000011111111 : 14'b00000111111111;
											assign node106 = (inp[0]) ? node110 : node107;
												assign node107 = (inp[13]) ? 14'b00000011111111 : 14'b00000111111111;
												assign node110 = (inp[2]) ? 14'b00000000111111 : 14'b00000011111111;
							assign node113 = (inp[0]) ? node171 : node114;
								assign node114 = (inp[7]) ? node142 : node115;
									assign node115 = (inp[10]) ? node131 : node116;
										assign node116 = (inp[13]) ? node124 : node117;
											assign node117 = (inp[11]) ? node121 : node118;
												assign node118 = (inp[2]) ? 14'b00011111111111 : 14'b00111111111111;
												assign node121 = (inp[2]) ? 14'b00001111111111 : 14'b00011111111111;
											assign node124 = (inp[11]) ? node128 : node125;
												assign node125 = (inp[9]) ? 14'b00001111111111 : 14'b00001111111111;
												assign node128 = (inp[8]) ? 14'b00000011111111 : 14'b00001111111111;
										assign node131 = (inp[9]) ? node137 : node132;
											assign node132 = (inp[8]) ? node134 : 14'b00001111111111;
												assign node134 = (inp[2]) ? 14'b00000111111111 : 14'b00001111111111;
											assign node137 = (inp[11]) ? 14'b00000111111111 : node138;
												assign node138 = (inp[13]) ? 14'b00000111111111 : 14'b00001111111111;
									assign node142 = (inp[9]) ? node158 : node143;
										assign node143 = (inp[13]) ? node151 : node144;
											assign node144 = (inp[10]) ? node148 : node145;
												assign node145 = (inp[11]) ? 14'b00001111111111 : 14'b00011111111111;
												assign node148 = (inp[11]) ? 14'b00000111111111 : 14'b00001111111111;
											assign node151 = (inp[10]) ? node155 : node152;
												assign node152 = (inp[8]) ? 14'b00000111111111 : 14'b00001111111111;
												assign node155 = (inp[11]) ? 14'b00000011111111 : 14'b00000111111111;
										assign node158 = (inp[10]) ? node166 : node159;
											assign node159 = (inp[8]) ? node163 : node160;
												assign node160 = (inp[13]) ? 14'b00000111111111 : 14'b00001111111111;
												assign node163 = (inp[13]) ? 14'b00000011111111 : 14'b00000111111111;
											assign node166 = (inp[2]) ? 14'b00000011111111 : node167;
												assign node167 = (inp[13]) ? 14'b00000011111111 : 14'b00000111111111;
								assign node171 = (inp[11]) ? node195 : node172;
									assign node172 = (inp[8]) ? node184 : node173;
										assign node173 = (inp[10]) ? node179 : node174;
											assign node174 = (inp[9]) ? 14'b00001111111111 : node175;
												assign node175 = (inp[2]) ? 14'b00001111111111 : 14'b00011111111111;
											assign node179 = (inp[13]) ? 14'b00000011111111 : node180;
												assign node180 = (inp[2]) ? 14'b00000111111111 : 14'b00001111111111;
										assign node184 = (inp[9]) ? node190 : node185;
											assign node185 = (inp[10]) ? node187 : 14'b00001111111111;
												assign node187 = (inp[2]) ? 14'b00000011111111 : 14'b00000111111111;
											assign node190 = (inp[7]) ? node192 : 14'b00000011111111;
												assign node192 = (inp[10]) ? 14'b00000000111111 : 14'b00000001111111;
									assign node195 = (inp[2]) ? node209 : node196;
										assign node196 = (inp[9]) ? node202 : node197;
											assign node197 = (inp[10]) ? node199 : 14'b00000011111111;
												assign node199 = (inp[7]) ? 14'b00000111111111 : 14'b00000111111111;
											assign node202 = (inp[7]) ? node206 : node203;
												assign node203 = (inp[13]) ? 14'b00000011111111 : 14'b00000111111111;
												assign node206 = (inp[13]) ? 14'b00000000111111 : 14'b00000011111111;
										assign node209 = (inp[7]) ? node215 : node210;
											assign node210 = (inp[9]) ? node212 : 14'b00000011111111;
												assign node212 = (inp[8]) ? 14'b00000001111111 : 14'b00000011111111;
											assign node215 = (inp[9]) ? node217 : 14'b00000001111111;
												assign node217 = (inp[8]) ? 14'b00000000011111 : 14'b00000001111111;
						assign node220 = (inp[8]) ? node326 : node221;
							assign node221 = (inp[7]) ? node273 : node222;
								assign node222 = (inp[13]) ? node254 : node223;
									assign node223 = (inp[2]) ? node239 : node224;
										assign node224 = (inp[9]) ? node232 : node225;
											assign node225 = (inp[11]) ? node229 : node226;
												assign node226 = (inp[10]) ? 14'b00011111111111 : 14'b00111111111111;
												assign node229 = (inp[0]) ? 14'b00001111111111 : 14'b00011111111111;
											assign node232 = (inp[4]) ? node236 : node233;
												assign node233 = (inp[0]) ? 14'b00001111111111 : 14'b00011111111111;
												assign node236 = (inp[10]) ? 14'b00000111111111 : 14'b00001111111111;
										assign node239 = (inp[10]) ? node247 : node240;
											assign node240 = (inp[0]) ? node244 : node241;
												assign node241 = (inp[11]) ? 14'b00001111111111 : 14'b00011111111111;
												assign node244 = (inp[9]) ? 14'b00000111111111 : 14'b00001111111111;
											assign node247 = (inp[9]) ? node251 : node248;
												assign node248 = (inp[4]) ? 14'b00000111111111 : 14'b00000111111111;
												assign node251 = (inp[0]) ? 14'b00000011111111 : 14'b00000111111111;
									assign node254 = (inp[9]) ? node262 : node255;
										assign node255 = (inp[0]) ? 14'b00000111111111 : node256;
											assign node256 = (inp[11]) ? node258 : 14'b00001111111111;
												assign node258 = (inp[2]) ? 14'b00000111111111 : 14'b00000111111111;
										assign node262 = (inp[10]) ? node268 : node263;
											assign node263 = (inp[0]) ? node265 : 14'b00001111111111;
												assign node265 = (inp[4]) ? 14'b00000011111111 : 14'b00000111111111;
											assign node268 = (inp[11]) ? 14'b00000011111111 : node269;
												assign node269 = (inp[4]) ? 14'b00000011111111 : 14'b00000111111111;
								assign node273 = (inp[11]) ? node303 : node274;
									assign node274 = (inp[13]) ? node288 : node275;
										assign node275 = (inp[0]) ? node281 : node276;
											assign node276 = (inp[4]) ? 14'b00001111111111 : node277;
												assign node277 = (inp[10]) ? 14'b00001111111111 : 14'b00011111111111;
											assign node281 = (inp[2]) ? node285 : node282;
												assign node282 = (inp[10]) ? 14'b00000011111111 : 14'b00001111111111;
												assign node285 = (inp[9]) ? 14'b00000011111111 : 14'b00000111111111;
										assign node288 = (inp[9]) ? node296 : node289;
											assign node289 = (inp[4]) ? node293 : node290;
												assign node290 = (inp[10]) ? 14'b00000111111111 : 14'b00001111111111;
												assign node293 = (inp[10]) ? 14'b00000011111111 : 14'b00000111111111;
											assign node296 = (inp[0]) ? node300 : node297;
												assign node297 = (inp[2]) ? 14'b00000011111111 : 14'b00000111111111;
												assign node300 = (inp[10]) ? 14'b00000001111111 : 14'b00000011111111;
									assign node303 = (inp[4]) ? node317 : node304;
										assign node304 = (inp[0]) ? node312 : node305;
											assign node305 = (inp[10]) ? node309 : node306;
												assign node306 = (inp[2]) ? 14'b00000111111111 : 14'b00001111111111;
												assign node309 = (inp[9]) ? 14'b00000011111111 : 14'b00000111111111;
											assign node312 = (inp[13]) ? node314 : 14'b00000011111111;
												assign node314 = (inp[10]) ? 14'b00000000111111 : 14'b00000011111111;
										assign node317 = (inp[9]) ? node319 : 14'b00000011111111;
											assign node319 = (inp[10]) ? node323 : node320;
												assign node320 = (inp[13]) ? 14'b00000001111111 : 14'b00000011111111;
												assign node323 = (inp[0]) ? 14'b00000000111111 : 14'b00000001111111;
							assign node326 = (inp[4]) ? node376 : node327;
								assign node327 = (inp[7]) ? node347 : node328;
									assign node328 = (inp[0]) ? node340 : node329;
										assign node329 = (inp[2]) ? node335 : node330;
											assign node330 = (inp[9]) ? node332 : 14'b00011111111111;
												assign node332 = (inp[11]) ? 14'b00001111111111 : 14'b00001111111111;
											assign node335 = (inp[11]) ? node337 : 14'b00001111111111;
												assign node337 = (inp[13]) ? 14'b00000111111111 : 14'b00001111111111;
										assign node340 = (inp[10]) ? node342 : 14'b00000111111111;
											assign node342 = (inp[11]) ? 14'b00000011111111 : node343;
												assign node343 = (inp[13]) ? 14'b00000011111111 : 14'b00000111111111;
									assign node347 = (inp[13]) ? node361 : node348;
										assign node348 = (inp[10]) ? node354 : node349;
											assign node349 = (inp[11]) ? 14'b00000111111111 : node350;
												assign node350 = (inp[0]) ? 14'b00001111111111 : 14'b00011111111111;
											assign node354 = (inp[11]) ? node358 : node355;
												assign node355 = (inp[2]) ? 14'b00000011111111 : 14'b00000111111111;
												assign node358 = (inp[2]) ? 14'b00000001111111 : 14'b00000011111111;
										assign node361 = (inp[11]) ? node369 : node362;
											assign node362 = (inp[2]) ? node366 : node363;
												assign node363 = (inp[0]) ? 14'b00000011111111 : 14'b00000111111111;
												assign node366 = (inp[9]) ? 14'b00000001111111 : 14'b00000011111111;
											assign node369 = (inp[9]) ? node373 : node370;
												assign node370 = (inp[10]) ? 14'b00000001111111 : 14'b00000011111111;
												assign node373 = (inp[2]) ? 14'b00000000111111 : 14'b00000000111111;
								assign node376 = (inp[11]) ? node396 : node377;
									assign node377 = (inp[10]) ? node387 : node378;
										assign node378 = (inp[13]) ? node384 : node379;
											assign node379 = (inp[2]) ? 14'b00000111111111 : node380;
												assign node380 = (inp[7]) ? 14'b00000011111111 : 14'b00000111111111;
											assign node384 = (inp[7]) ? 14'b00000000111111 : 14'b00000011111111;
										assign node387 = (inp[7]) ? node393 : node388;
											assign node388 = (inp[13]) ? node390 : 14'b00000011111111;
												assign node390 = (inp[9]) ? 14'b00000001111111 : 14'b00000011111111;
											assign node393 = (inp[0]) ? 14'b00000001111111 : 14'b00000011111111;
									assign node396 = (inp[9]) ? node404 : node397;
										assign node397 = (inp[10]) ? 14'b00000001111111 : node398;
											assign node398 = (inp[13]) ? node400 : 14'b00000111111111;
												assign node400 = (inp[7]) ? 14'b00000001111111 : 14'b00000011111111;
										assign node404 = (inp[7]) ? node412 : node405;
											assign node405 = (inp[0]) ? node409 : node406;
												assign node406 = (inp[13]) ? 14'b00000001111111 : 14'b00000011111111;
												assign node409 = (inp[2]) ? 14'b00000000111111 : 14'b00000001111111;
											assign node412 = (inp[0]) ? node414 : 14'b00000000111111;
												assign node414 = (inp[13]) ? 14'b00000000011111 : 14'b00000000111111;
					assign node417 = (inp[10]) ? node631 : node418;
						assign node418 = (inp[0]) ? node528 : node419;
							assign node419 = (inp[9]) ? node477 : node420;
								assign node420 = (inp[2]) ? node450 : node421;
									assign node421 = (inp[13]) ? node437 : node422;
										assign node422 = (inp[7]) ? node430 : node423;
											assign node423 = (inp[12]) ? node427 : node424;
												assign node424 = (inp[4]) ? 14'b00011111111111 : 14'b00111111111111;
												assign node427 = (inp[4]) ? 14'b00001111111111 : 14'b00011111111111;
											assign node430 = (inp[8]) ? node434 : node431;
												assign node431 = (inp[4]) ? 14'b00001111111111 : 14'b00011111111111;
												assign node434 = (inp[12]) ? 14'b00000011111111 : 14'b00001111111111;
										assign node437 = (inp[11]) ? node443 : node438;
											assign node438 = (inp[8]) ? node440 : 14'b00001111111111;
												assign node440 = (inp[4]) ? 14'b00000111111111 : 14'b00001111111111;
											assign node443 = (inp[4]) ? node447 : node444;
												assign node444 = (inp[12]) ? 14'b00000111111111 : 14'b00001111111111;
												assign node447 = (inp[7]) ? 14'b00000011111111 : 14'b00000111111111;
									assign node450 = (inp[7]) ? node462 : node451;
										assign node451 = (inp[8]) ? node457 : node452;
											assign node452 = (inp[12]) ? node454 : 14'b00001111111111;
												assign node454 = (inp[11]) ? 14'b00000111111111 : 14'b00001111111111;
											assign node457 = (inp[4]) ? 14'b00000111111111 : node458;
												assign node458 = (inp[11]) ? 14'b00000111111111 : 14'b00001111111111;
										assign node462 = (inp[4]) ? node470 : node463;
											assign node463 = (inp[12]) ? node467 : node464;
												assign node464 = (inp[11]) ? 14'b00001111111111 : 14'b00001111111111;
												assign node467 = (inp[8]) ? 14'b00000011111111 : 14'b00000111111111;
											assign node470 = (inp[11]) ? node474 : node471;
												assign node471 = (inp[8]) ? 14'b00000011111111 : 14'b00000111111111;
												assign node474 = (inp[13]) ? 14'b00000001111111 : 14'b00000011111111;
								assign node477 = (inp[7]) ? node505 : node478;
									assign node478 = (inp[13]) ? node492 : node479;
										assign node479 = (inp[8]) ? node487 : node480;
											assign node480 = (inp[2]) ? node484 : node481;
												assign node481 = (inp[11]) ? 14'b00001111111111 : 14'b00111111111111;
												assign node484 = (inp[11]) ? 14'b00000111111111 : 14'b00001111111111;
											assign node487 = (inp[12]) ? 14'b00000011111111 : node488;
												assign node488 = (inp[2]) ? 14'b00000111111111 : 14'b00000111111111;
										assign node492 = (inp[2]) ? node500 : node493;
											assign node493 = (inp[11]) ? node497 : node494;
												assign node494 = (inp[4]) ? 14'b00000111111111 : 14'b00001111111111;
												assign node497 = (inp[8]) ? 14'b00000011111111 : 14'b00000111111111;
											assign node500 = (inp[4]) ? node502 : 14'b00000011111111;
												assign node502 = (inp[11]) ? 14'b00000001111111 : 14'b00000001111111;
									assign node505 = (inp[2]) ? node517 : node506;
										assign node506 = (inp[12]) ? node512 : node507;
											assign node507 = (inp[11]) ? node509 : 14'b00000111111111;
												assign node509 = (inp[8]) ? 14'b00000011111111 : 14'b00000111111111;
											assign node512 = (inp[4]) ? 14'b00000001111111 : node513;
												assign node513 = (inp[13]) ? 14'b00000111111111 : 14'b00000011111111;
										assign node517 = (inp[8]) ? node523 : node518;
											assign node518 = (inp[13]) ? 14'b00000001111111 : node519;
												assign node519 = (inp[11]) ? 14'b00000011111111 : 14'b00000111111111;
											assign node523 = (inp[13]) ? node525 : 14'b00000001111111;
												assign node525 = (inp[4]) ? 14'b00000000011111 : 14'b00000000111111;
							assign node528 = (inp[12]) ? node584 : node529;
								assign node529 = (inp[13]) ? node557 : node530;
									assign node530 = (inp[8]) ? node544 : node531;
										assign node531 = (inp[7]) ? node539 : node532;
											assign node532 = (inp[4]) ? node536 : node533;
												assign node533 = (inp[2]) ? 14'b00001111111111 : 14'b00011111111111;
												assign node536 = (inp[11]) ? 14'b00000111111111 : 14'b00001111111111;
											assign node539 = (inp[9]) ? 14'b00000011111111 : node540;
												assign node540 = (inp[11]) ? 14'b00000111111111 : 14'b00001111111111;
										assign node544 = (inp[2]) ? node550 : node545;
											assign node545 = (inp[11]) ? node547 : 14'b00000111111111;
												assign node547 = (inp[9]) ? 14'b00000011111111 : 14'b00000011111111;
											assign node550 = (inp[11]) ? node554 : node551;
												assign node551 = (inp[4]) ? 14'b00000011111111 : 14'b00000011111111;
												assign node554 = (inp[9]) ? 14'b00000001111111 : 14'b00000011111111;
									assign node557 = (inp[8]) ? node571 : node558;
										assign node558 = (inp[11]) ? node564 : node559;
											assign node559 = (inp[4]) ? node561 : 14'b00000111111111;
												assign node561 = (inp[9]) ? 14'b00000011111111 : 14'b00000111111111;
											assign node564 = (inp[2]) ? node568 : node565;
												assign node565 = (inp[9]) ? 14'b00000011111111 : 14'b00000111111111;
												assign node568 = (inp[7]) ? 14'b00000001111111 : 14'b00000011111111;
										assign node571 = (inp[11]) ? node579 : node572;
											assign node572 = (inp[4]) ? node576 : node573;
												assign node573 = (inp[9]) ? 14'b00000011111111 : 14'b00000111111111;
												assign node576 = (inp[9]) ? 14'b00000001111111 : 14'b00000011111111;
											assign node579 = (inp[4]) ? 14'b00000001111111 : node580;
												assign node580 = (inp[7]) ? 14'b00000001111111 : 14'b00000011111111;
								assign node584 = (inp[11]) ? node608 : node585;
									assign node585 = (inp[9]) ? node595 : node586;
										assign node586 = (inp[8]) ? node592 : node587;
											assign node587 = (inp[2]) ? 14'b00000111111111 : node588;
												assign node588 = (inp[13]) ? 14'b00000111111111 : 14'b00011111111111;
											assign node592 = (inp[13]) ? 14'b00000011111111 : 14'b00000111111111;
										assign node595 = (inp[13]) ? node603 : node596;
											assign node596 = (inp[2]) ? node600 : node597;
												assign node597 = (inp[7]) ? 14'b00000011111111 : 14'b00000111111111;
												assign node600 = (inp[7]) ? 14'b00000001111111 : 14'b00000011111111;
											assign node603 = (inp[2]) ? 14'b00000000111111 : node604;
												assign node604 = (inp[8]) ? 14'b00000000111111 : 14'b00000001111111;
									assign node608 = (inp[7]) ? node620 : node609;
										assign node609 = (inp[8]) ? node615 : node610;
											assign node610 = (inp[4]) ? node612 : 14'b00000011111111;
												assign node612 = (inp[2]) ? 14'b00000001111111 : 14'b00000011111111;
											assign node615 = (inp[13]) ? node617 : 14'b00000011111111;
												assign node617 = (inp[2]) ? 14'b00000000111111 : 14'b00000001111111;
										assign node620 = (inp[2]) ? node628 : node621;
											assign node621 = (inp[13]) ? node625 : node622;
												assign node622 = (inp[8]) ? 14'b00000000111111 : 14'b00000011111111;
												assign node625 = (inp[9]) ? 14'b00000000111111 : 14'b00000001111111;
											assign node628 = (inp[9]) ? 14'b00000000011111 : 14'b00000000111111;
						assign node631 = (inp[7]) ? node741 : node632;
							assign node632 = (inp[0]) ? node692 : node633;
								assign node633 = (inp[13]) ? node663 : node634;
									assign node634 = (inp[9]) ? node650 : node635;
										assign node635 = (inp[2]) ? node643 : node636;
											assign node636 = (inp[12]) ? node640 : node637;
												assign node637 = (inp[4]) ? 14'b00001111111111 : 14'b00011111111111;
												assign node640 = (inp[8]) ? 14'b00000111111111 : 14'b00001111111111;
											assign node643 = (inp[8]) ? node647 : node644;
												assign node644 = (inp[12]) ? 14'b00000111111111 : 14'b00001111111111;
												assign node647 = (inp[11]) ? 14'b00000011111111 : 14'b00000111111111;
										assign node650 = (inp[2]) ? node658 : node651;
											assign node651 = (inp[8]) ? node655 : node652;
												assign node652 = (inp[12]) ? 14'b00000111111111 : 14'b00001111111111;
												assign node655 = (inp[12]) ? 14'b00000011111111 : 14'b00000111111111;
											assign node658 = (inp[12]) ? 14'b00000011111111 : node659;
												assign node659 = (inp[11]) ? 14'b00000011111111 : 14'b00001111111111;
									assign node663 = (inp[4]) ? node677 : node664;
										assign node664 = (inp[2]) ? node672 : node665;
											assign node665 = (inp[8]) ? node669 : node666;
												assign node666 = (inp[11]) ? 14'b00000111111111 : 14'b00000111111111;
												assign node669 = (inp[12]) ? 14'b00000011111111 : 14'b00000111111111;
											assign node672 = (inp[12]) ? 14'b00000001111111 : node673;
												assign node673 = (inp[9]) ? 14'b00000011111111 : 14'b00000111111111;
										assign node677 = (inp[9]) ? node685 : node678;
											assign node678 = (inp[11]) ? node682 : node679;
												assign node679 = (inp[8]) ? 14'b00000011111111 : 14'b00000111111111;
												assign node682 = (inp[8]) ? 14'b00000001111111 : 14'b00000011111111;
											assign node685 = (inp[8]) ? node689 : node686;
												assign node686 = (inp[2]) ? 14'b00000001111111 : 14'b00000011111111;
												assign node689 = (inp[2]) ? 14'b00000000011111 : 14'b00000001111111;
								assign node692 = (inp[2]) ? node716 : node693;
									assign node693 = (inp[11]) ? node709 : node694;
										assign node694 = (inp[8]) ? node702 : node695;
											assign node695 = (inp[4]) ? node699 : node696;
												assign node696 = (inp[12]) ? 14'b00000111111111 : 14'b00011111111111;
												assign node699 = (inp[12]) ? 14'b00000011111111 : 14'b00000111111111;
											assign node702 = (inp[9]) ? node706 : node703;
												assign node703 = (inp[13]) ? 14'b00000011111111 : 14'b00000111111111;
												assign node706 = (inp[12]) ? 14'b00000001111111 : 14'b00000011111111;
										assign node709 = (inp[4]) ? 14'b00000001111111 : node710;
											assign node710 = (inp[12]) ? 14'b00000001111111 : node711;
												assign node711 = (inp[13]) ? 14'b00000011111111 : 14'b00000011111111;
									assign node716 = (inp[9]) ? node730 : node717;
										assign node717 = (inp[12]) ? node723 : node718;
											assign node718 = (inp[8]) ? 14'b00000011111111 : node719;
												assign node719 = (inp[4]) ? 14'b00000001111111 : 14'b00000011111111;
											assign node723 = (inp[4]) ? node727 : node724;
												assign node724 = (inp[8]) ? 14'b00000011111111 : 14'b00000001111111;
												assign node727 = (inp[11]) ? 14'b00000000111111 : 14'b00000001111111;
										assign node730 = (inp[13]) ? node736 : node731;
											assign node731 = (inp[11]) ? node733 : 14'b00000001111111;
												assign node733 = (inp[8]) ? 14'b00000000111111 : 14'b00000001111111;
											assign node736 = (inp[12]) ? node738 : 14'b00000000111111;
												assign node738 = (inp[11]) ? 14'b00000000011111 : 14'b00000000111111;
							assign node741 = (inp[11]) ? node789 : node742;
								assign node742 = (inp[9]) ? node760 : node743;
									assign node743 = (inp[4]) ? node753 : node744;
										assign node744 = (inp[2]) ? node748 : node745;
											assign node745 = (inp[12]) ? 14'b00000111111111 : 14'b00001111111111;
											assign node748 = (inp[0]) ? 14'b00000011111111 : node749;
												assign node749 = (inp[13]) ? 14'b00000011111111 : 14'b00000111111111;
										assign node753 = (inp[2]) ? node755 : 14'b00000011111111;
											assign node755 = (inp[13]) ? 14'b00000000111111 : node756;
												assign node756 = (inp[12]) ? 14'b00000001111111 : 14'b00000011111111;
									assign node760 = (inp[12]) ? node774 : node761;
										assign node761 = (inp[0]) ? node769 : node762;
											assign node762 = (inp[8]) ? node766 : node763;
												assign node763 = (inp[4]) ? 14'b00000011111111 : 14'b00000111111111;
												assign node766 = (inp[13]) ? 14'b00000001111111 : 14'b00000011111111;
											assign node769 = (inp[13]) ? node771 : 14'b00000011111111;
												assign node771 = (inp[2]) ? 14'b00000000111111 : 14'b00000001111111;
										assign node774 = (inp[8]) ? node782 : node775;
											assign node775 = (inp[2]) ? node779 : node776;
												assign node776 = (inp[13]) ? 14'b00000001111111 : 14'b00000011111111;
												assign node779 = (inp[13]) ? 14'b00000000111111 : 14'b00000001111111;
											assign node782 = (inp[2]) ? node786 : node783;
												assign node783 = (inp[0]) ? 14'b00000000111111 : 14'b00000000111111;
												assign node786 = (inp[0]) ? 14'b00000000011111 : 14'b00000000011111;
								assign node789 = (inp[9]) ? node819 : node790;
									assign node790 = (inp[4]) ? node804 : node791;
										assign node791 = (inp[0]) ? node799 : node792;
											assign node792 = (inp[2]) ? node796 : node793;
												assign node793 = (inp[12]) ? 14'b00000001111111 : 14'b00000011111111;
												assign node796 = (inp[12]) ? 14'b00000011111111 : 14'b00000011111111;
											assign node799 = (inp[2]) ? 14'b00000001111111 : node800;
												assign node800 = (inp[8]) ? 14'b00000001111111 : 14'b00000111111111;
										assign node804 = (inp[0]) ? node812 : node805;
											assign node805 = (inp[12]) ? node809 : node806;
												assign node806 = (inp[2]) ? 14'b00000001111111 : 14'b00000011111111;
												assign node809 = (inp[13]) ? 14'b00000000111111 : 14'b00000001111111;
											assign node812 = (inp[2]) ? node816 : node813;
												assign node813 = (inp[12]) ? 14'b00000000111111 : 14'b00000001111111;
												assign node816 = (inp[8]) ? 14'b00000000011111 : 14'b00000000111111;
									assign node819 = (inp[13]) ? node833 : node820;
										assign node820 = (inp[12]) ? node826 : node821;
											assign node821 = (inp[8]) ? node823 : 14'b00000001111111;
												assign node823 = (inp[0]) ? 14'b00000000111111 : 14'b00000001111111;
											assign node826 = (inp[4]) ? node830 : node827;
												assign node827 = (inp[8]) ? 14'b00000000111111 : 14'b00000001111111;
												assign node830 = (inp[8]) ? 14'b00000000001111 : 14'b00000000111111;
										assign node833 = (inp[0]) ? node841 : node834;
											assign node834 = (inp[8]) ? node838 : node835;
												assign node835 = (inp[12]) ? 14'b00000000111111 : 14'b00000000111111;
												assign node838 = (inp[4]) ? 14'b00000000011111 : 14'b00000000111111;
											assign node841 = (inp[2]) ? node845 : node842;
												assign node842 = (inp[4]) ? 14'b00000000011111 : 14'b00000000011111;
												assign node845 = (inp[12]) ? 14'b00000000001111 : 14'b00000000011111;
				assign node848 = (inp[2]) ? node1262 : node849;
					assign node849 = (inp[8]) ? node1059 : node850;
						assign node850 = (inp[6]) ? node950 : node851;
							assign node851 = (inp[10]) ? node897 : node852;
								assign node852 = (inp[12]) ? node874 : node853;
									assign node853 = (inp[4]) ? node865 : node854;
										assign node854 = (inp[7]) ? node860 : node855;
											assign node855 = (inp[11]) ? 14'b00001111111111 : node856;
												assign node856 = (inp[9]) ? 14'b00011111111111 : 14'b00111111111111;
											assign node860 = (inp[9]) ? node862 : 14'b00011111111111;
												assign node862 = (inp[13]) ? 14'b00001111111111 : 14'b00001111111111;
										assign node865 = (inp[9]) ? node867 : 14'b00001111111111;
											assign node867 = (inp[7]) ? node871 : node868;
												assign node868 = (inp[0]) ? 14'b00000111111111 : 14'b00011111111111;
												assign node871 = (inp[0]) ? 14'b00000011111111 : 14'b00000111111111;
									assign node874 = (inp[0]) ? node884 : node875;
										assign node875 = (inp[13]) ? node879 : node876;
											assign node876 = (inp[4]) ? 14'b00001111111111 : 14'b00011111111111;
											assign node879 = (inp[11]) ? 14'b00000111111111 : node880;
												assign node880 = (inp[7]) ? 14'b00000111111111 : 14'b00001111111111;
										assign node884 = (inp[11]) ? node892 : node885;
											assign node885 = (inp[7]) ? node889 : node886;
												assign node886 = (inp[13]) ? 14'b00000111111111 : 14'b00001111111111;
												assign node889 = (inp[13]) ? 14'b00000011111111 : 14'b00000111111111;
											assign node892 = (inp[9]) ? 14'b00000011111111 : node893;
												assign node893 = (inp[7]) ? 14'b00000001111111 : 14'b00000111111111;
								assign node897 = (inp[4]) ? node927 : node898;
									assign node898 = (inp[12]) ? node914 : node899;
										assign node899 = (inp[11]) ? node907 : node900;
											assign node900 = (inp[9]) ? node904 : node901;
												assign node901 = (inp[7]) ? 14'b00001111111111 : 14'b00011111111111;
												assign node904 = (inp[0]) ? 14'b00000111111111 : 14'b00001111111111;
											assign node907 = (inp[13]) ? node911 : node908;
												assign node908 = (inp[0]) ? 14'b00000111111111 : 14'b00001111111111;
												assign node911 = (inp[0]) ? 14'b00000011111111 : 14'b00000111111111;
										assign node914 = (inp[11]) ? node922 : node915;
											assign node915 = (inp[0]) ? node919 : node916;
												assign node916 = (inp[9]) ? 14'b00000111111111 : 14'b00001111111111;
												assign node919 = (inp[9]) ? 14'b00000011111111 : 14'b00000111111111;
											assign node922 = (inp[13]) ? 14'b00000011111111 : node923;
												assign node923 = (inp[9]) ? 14'b00000011111111 : 14'b00000011111111;
									assign node927 = (inp[11]) ? node939 : node928;
										assign node928 = (inp[12]) ? node934 : node929;
											assign node929 = (inp[9]) ? node931 : 14'b00000111111111;
												assign node931 = (inp[13]) ? 14'b00000011111111 : 14'b00001111111111;
											assign node934 = (inp[13]) ? 14'b00000001111111 : node935;
												assign node935 = (inp[7]) ? 14'b00000111111111 : 14'b00000011111111;
										assign node939 = (inp[13]) ? node945 : node940;
											assign node940 = (inp[7]) ? node942 : 14'b00000011111111;
												assign node942 = (inp[0]) ? 14'b00000011111111 : 14'b00000001111111;
											assign node945 = (inp[12]) ? 14'b00000000111111 : node946;
												assign node946 = (inp[9]) ? 14'b00000001111111 : 14'b00000011111111;
							assign node950 = (inp[0]) ? node1008 : node951;
								assign node951 = (inp[7]) ? node981 : node952;
									assign node952 = (inp[10]) ? node966 : node953;
										assign node953 = (inp[9]) ? node961 : node954;
											assign node954 = (inp[13]) ? node958 : node955;
												assign node955 = (inp[12]) ? 14'b00001111111111 : 14'b00011111111111;
												assign node958 = (inp[4]) ? 14'b00000111111111 : 14'b00001111111111;
											assign node961 = (inp[4]) ? 14'b00000011111111 : node962;
												assign node962 = (inp[11]) ? 14'b00000111111111 : 14'b00000111111111;
										assign node966 = (inp[13]) ? node974 : node967;
											assign node967 = (inp[11]) ? node971 : node968;
												assign node968 = (inp[4]) ? 14'b00000111111111 : 14'b00001111111111;
												assign node971 = (inp[9]) ? 14'b00000011111111 : 14'b00000111111111;
											assign node974 = (inp[4]) ? node978 : node975;
												assign node975 = (inp[12]) ? 14'b00000011111111 : 14'b00000111111111;
												assign node978 = (inp[11]) ? 14'b00000001111111 : 14'b00000011111111;
									assign node981 = (inp[11]) ? node995 : node982;
										assign node982 = (inp[9]) ? node990 : node983;
											assign node983 = (inp[13]) ? node987 : node984;
												assign node984 = (inp[12]) ? 14'b00000111111111 : 14'b00001111111111;
												assign node987 = (inp[4]) ? 14'b00000011111111 : 14'b00000111111111;
											assign node990 = (inp[12]) ? 14'b00000001111111 : node991;
												assign node991 = (inp[10]) ? 14'b00000011111111 : 14'b00000111111111;
										assign node995 = (inp[12]) ? node1003 : node996;
											assign node996 = (inp[9]) ? node1000 : node997;
												assign node997 = (inp[13]) ? 14'b00000011111111 : 14'b00000111111111;
												assign node1000 = (inp[13]) ? 14'b00000001111111 : 14'b00000011111111;
											assign node1003 = (inp[9]) ? 14'b00000000111111 : node1004;
												assign node1004 = (inp[4]) ? 14'b00000001111111 : 14'b00000011111111;
								assign node1008 = (inp[9]) ? node1036 : node1009;
									assign node1009 = (inp[4]) ? node1021 : node1010;
										assign node1010 = (inp[7]) ? node1016 : node1011;
											assign node1011 = (inp[11]) ? node1013 : 14'b00000111111111;
												assign node1013 = (inp[12]) ? 14'b00000011111111 : 14'b00000011111111;
											assign node1016 = (inp[13]) ? 14'b00000011111111 : node1017;
												assign node1017 = (inp[11]) ? 14'b00000011111111 : 14'b00000111111111;
										assign node1021 = (inp[13]) ? node1029 : node1022;
											assign node1022 = (inp[7]) ? node1026 : node1023;
												assign node1023 = (inp[12]) ? 14'b00000011111111 : 14'b00000111111111;
												assign node1026 = (inp[10]) ? 14'b00000001111111 : 14'b00000011111111;
											assign node1029 = (inp[11]) ? node1033 : node1030;
												assign node1030 = (inp[7]) ? 14'b00000000111111 : 14'b00000001111111;
												assign node1033 = (inp[10]) ? 14'b00000000111111 : 14'b00000000111111;
									assign node1036 = (inp[12]) ? node1050 : node1037;
										assign node1037 = (inp[4]) ? node1043 : node1038;
											assign node1038 = (inp[7]) ? node1040 : 14'b00000011111111;
												assign node1040 = (inp[13]) ? 14'b00000001111111 : 14'b00000011111111;
											assign node1043 = (inp[10]) ? node1047 : node1044;
												assign node1044 = (inp[13]) ? 14'b00000001111111 : 14'b00000011111111;
												assign node1047 = (inp[13]) ? 14'b00000000011111 : 14'b00000001111111;
										assign node1050 = (inp[10]) ? node1054 : node1051;
											assign node1051 = (inp[7]) ? 14'b00000000111111 : 14'b00000001111111;
											assign node1054 = (inp[13]) ? node1056 : 14'b00000001111111;
												assign node1056 = (inp[4]) ? 14'b00000000011111 : 14'b00000000111111;
						assign node1059 = (inp[11]) ? node1157 : node1060;
							assign node1060 = (inp[6]) ? node1104 : node1061;
								assign node1061 = (inp[12]) ? node1087 : node1062;
									assign node1062 = (inp[0]) ? node1076 : node1063;
										assign node1063 = (inp[10]) ? node1071 : node1064;
											assign node1064 = (inp[4]) ? node1068 : node1065;
												assign node1065 = (inp[13]) ? 14'b00001111111111 : 14'b00011111111111;
												assign node1068 = (inp[9]) ? 14'b00000111111111 : 14'b00001111111111;
											assign node1071 = (inp[9]) ? 14'b00000111111111 : node1072;
												assign node1072 = (inp[4]) ? 14'b00000111111111 : 14'b00001111111111;
										assign node1076 = (inp[9]) ? node1082 : node1077;
											assign node1077 = (inp[13]) ? node1079 : 14'b00001111111111;
												assign node1079 = (inp[4]) ? 14'b00000111111111 : 14'b00001111111111;
											assign node1082 = (inp[10]) ? 14'b00000001111111 : node1083;
												assign node1083 = (inp[4]) ? 14'b00000011111111 : 14'b00000111111111;
									assign node1087 = (inp[0]) ? node1095 : node1088;
										assign node1088 = (inp[13]) ? 14'b00000011111111 : node1089;
											assign node1089 = (inp[9]) ? node1091 : 14'b00000111111111;
												assign node1091 = (inp[7]) ? 14'b00000001111111 : 14'b00000011111111;
										assign node1095 = (inp[10]) ? node1101 : node1096;
											assign node1096 = (inp[4]) ? 14'b00000011111111 : node1097;
												assign node1097 = (inp[13]) ? 14'b00000011111111 : 14'b00000111111111;
											assign node1101 = (inp[9]) ? 14'b00000000111111 : 14'b00000001111111;
								assign node1104 = (inp[7]) ? node1130 : node1105;
									assign node1105 = (inp[0]) ? node1119 : node1106;
										assign node1106 = (inp[13]) ? node1112 : node1107;
											assign node1107 = (inp[4]) ? node1109 : 14'b00000111111111;
												assign node1109 = (inp[12]) ? 14'b00000011111111 : 14'b00000111111111;
											assign node1112 = (inp[9]) ? node1116 : node1113;
												assign node1113 = (inp[4]) ? 14'b00000011111111 : 14'b00000111111111;
												assign node1116 = (inp[12]) ? 14'b00000001111111 : 14'b00000001111111;
										assign node1119 = (inp[13]) ? node1127 : node1120;
											assign node1120 = (inp[12]) ? node1124 : node1121;
												assign node1121 = (inp[4]) ? 14'b00000011111111 : 14'b00000011111111;
												assign node1124 = (inp[4]) ? 14'b00000001111111 : 14'b00000011111111;
											assign node1127 = (inp[10]) ? 14'b00000000111111 : 14'b00000111111111;
									assign node1130 = (inp[4]) ? node1144 : node1131;
										assign node1131 = (inp[10]) ? node1139 : node1132;
											assign node1132 = (inp[9]) ? node1136 : node1133;
												assign node1133 = (inp[13]) ? 14'b00000011111111 : 14'b00000111111111;
												assign node1136 = (inp[0]) ? 14'b00000001111111 : 14'b00000011111111;
											assign node1139 = (inp[12]) ? node1141 : 14'b00000001111111;
												assign node1141 = (inp[9]) ? 14'b00000000111111 : 14'b00000001111111;
										assign node1144 = (inp[0]) ? node1150 : node1145;
											assign node1145 = (inp[13]) ? 14'b00000001111111 : node1146;
												assign node1146 = (inp[12]) ? 14'b00000001111111 : 14'b00000011111111;
											assign node1150 = (inp[13]) ? node1154 : node1151;
												assign node1151 = (inp[12]) ? 14'b00000000111111 : 14'b00000001111111;
												assign node1154 = (inp[10]) ? 14'b00000000001111 : 14'b00000000111111;
							assign node1157 = (inp[13]) ? node1215 : node1158;
								assign node1158 = (inp[4]) ? node1188 : node1159;
									assign node1159 = (inp[0]) ? node1175 : node1160;
										assign node1160 = (inp[7]) ? node1168 : node1161;
											assign node1161 = (inp[6]) ? node1165 : node1162;
												assign node1162 = (inp[9]) ? 14'b00000111111111 : 14'b00001111111111;
												assign node1165 = (inp[10]) ? 14'b00000011111111 : 14'b00000111111111;
											assign node1168 = (inp[10]) ? node1172 : node1169;
												assign node1169 = (inp[6]) ? 14'b00000011111111 : 14'b00000111111111;
												assign node1172 = (inp[12]) ? 14'b00000001111111 : 14'b00000011111111;
										assign node1175 = (inp[10]) ? node1183 : node1176;
											assign node1176 = (inp[12]) ? node1180 : node1177;
												assign node1177 = (inp[6]) ? 14'b00000011111111 : 14'b00000111111111;
												assign node1180 = (inp[9]) ? 14'b00000001111111 : 14'b00000011111111;
											assign node1183 = (inp[7]) ? node1185 : 14'b00000011111111;
												assign node1185 = (inp[9]) ? 14'b00000000111111 : 14'b00000001111111;
									assign node1188 = (inp[0]) ? node1204 : node1189;
										assign node1189 = (inp[6]) ? node1197 : node1190;
											assign node1190 = (inp[12]) ? node1194 : node1191;
												assign node1191 = (inp[10]) ? 14'b00000011111111 : 14'b00000111111111;
												assign node1194 = (inp[10]) ? 14'b00000001111111 : 14'b00000001111111;
											assign node1197 = (inp[10]) ? node1201 : node1198;
												assign node1198 = (inp[7]) ? 14'b00000001111111 : 14'b00000011111111;
												assign node1201 = (inp[7]) ? 14'b00000000011111 : 14'b00000000111111;
										assign node1204 = (inp[12]) ? node1210 : node1205;
											assign node1205 = (inp[7]) ? 14'b00000000111111 : node1206;
												assign node1206 = (inp[10]) ? 14'b00000001111111 : 14'b00000011111111;
											assign node1210 = (inp[6]) ? node1212 : 14'b00000000111111;
												assign node1212 = (inp[10]) ? 14'b00000000011111 : 14'b00000000111111;
								assign node1215 = (inp[7]) ? node1237 : node1216;
									assign node1216 = (inp[12]) ? node1226 : node1217;
										assign node1217 = (inp[6]) ? node1221 : node1218;
											assign node1218 = (inp[4]) ? 14'b00000000111111 : 14'b00000111111111;
											assign node1221 = (inp[9]) ? 14'b00000001111111 : node1222;
												assign node1222 = (inp[4]) ? 14'b00000001111111 : 14'b00000011111111;
										assign node1226 = (inp[10]) ? node1230 : node1227;
											assign node1227 = (inp[9]) ? 14'b00000001111111 : 14'b00000000111111;
											assign node1230 = (inp[9]) ? node1234 : node1231;
												assign node1231 = (inp[6]) ? 14'b00000000111111 : 14'b00000001111111;
												assign node1234 = (inp[4]) ? 14'b00000000011111 : 14'b00000000111111;
									assign node1237 = (inp[12]) ? node1251 : node1238;
										assign node1238 = (inp[6]) ? node1244 : node1239;
											assign node1239 = (inp[4]) ? node1241 : 14'b00000001111111;
												assign node1241 = (inp[9]) ? 14'b00000000011111 : 14'b00000001111111;
											assign node1244 = (inp[0]) ? node1248 : node1245;
												assign node1245 = (inp[9]) ? 14'b00000000111111 : 14'b00000000111111;
												assign node1248 = (inp[10]) ? 14'b00000000001111 : 14'b00000000111111;
										assign node1251 = (inp[9]) ? node1257 : node1252;
											assign node1252 = (inp[6]) ? 14'b00000000011111 : node1253;
												assign node1253 = (inp[0]) ? 14'b00000000011111 : 14'b00000001111111;
											assign node1257 = (inp[10]) ? node1259 : 14'b00000000011111;
												assign node1259 = (inp[4]) ? 14'b00000000001111 : 14'b00000000111111;
					assign node1262 = (inp[9]) ? node1448 : node1263;
						assign node1263 = (inp[0]) ? node1367 : node1264;
							assign node1264 = (inp[12]) ? node1310 : node1265;
								assign node1265 = (inp[4]) ? node1283 : node1266;
									assign node1266 = (inp[6]) ? node1276 : node1267;
										assign node1267 = (inp[8]) ? node1273 : node1268;
											assign node1268 = (inp[13]) ? node1270 : 14'b00001111111111;
												assign node1270 = (inp[10]) ? 14'b00000111111111 : 14'b00001111111111;
											assign node1273 = (inp[11]) ? 14'b00000011111111 : 14'b00000111111111;
										assign node1276 = (inp[10]) ? node1278 : 14'b00000111111111;
											assign node1278 = (inp[11]) ? 14'b00000011111111 : node1279;
												assign node1279 = (inp[7]) ? 14'b00000011111111 : 14'b00000111111111;
									assign node1283 = (inp[13]) ? node1295 : node1284;
										assign node1284 = (inp[6]) ? node1290 : node1285;
											assign node1285 = (inp[11]) ? node1287 : 14'b00001111111111;
												assign node1287 = (inp[7]) ? 14'b00000011111111 : 14'b00000111111111;
											assign node1290 = (inp[11]) ? 14'b00000011111111 : node1291;
												assign node1291 = (inp[7]) ? 14'b00000011111111 : 14'b00000111111111;
										assign node1295 = (inp[8]) ? node1303 : node1296;
											assign node1296 = (inp[11]) ? node1300 : node1297;
												assign node1297 = (inp[7]) ? 14'b00000011111111 : 14'b00000111111111;
												assign node1300 = (inp[7]) ? 14'b00000001111111 : 14'b00000011111111;
											assign node1303 = (inp[11]) ? node1307 : node1304;
												assign node1304 = (inp[7]) ? 14'b00000011111111 : 14'b00000001111111;
												assign node1307 = (inp[7]) ? 14'b00000000111111 : 14'b00000001111111;
								assign node1310 = (inp[6]) ? node1342 : node1311;
									assign node1311 = (inp[13]) ? node1327 : node1312;
										assign node1312 = (inp[7]) ? node1320 : node1313;
											assign node1313 = (inp[4]) ? node1317 : node1314;
												assign node1314 = (inp[10]) ? 14'b00000111111111 : 14'b00001111111111;
												assign node1317 = (inp[8]) ? 14'b00000111111111 : 14'b00000011111111;
											assign node1320 = (inp[11]) ? node1324 : node1321;
												assign node1321 = (inp[10]) ? 14'b00000011111111 : 14'b00000111111111;
												assign node1324 = (inp[8]) ? 14'b00000001111111 : 14'b00000011111111;
										assign node1327 = (inp[10]) ? node1335 : node1328;
											assign node1328 = (inp[11]) ? node1332 : node1329;
												assign node1329 = (inp[7]) ? 14'b00000011111111 : 14'b00000111111111;
												assign node1332 = (inp[7]) ? 14'b00000001111111 : 14'b00000011111111;
											assign node1335 = (inp[8]) ? node1339 : node1336;
												assign node1336 = (inp[4]) ? 14'b00000001111111 : 14'b00000011111111;
												assign node1339 = (inp[4]) ? 14'b00000000111111 : 14'b00000001111111;
									assign node1342 = (inp[11]) ? node1358 : node1343;
										assign node1343 = (inp[10]) ? node1351 : node1344;
											assign node1344 = (inp[8]) ? node1348 : node1345;
												assign node1345 = (inp[13]) ? 14'b00000011111111 : 14'b00000111111111;
												assign node1348 = (inp[7]) ? 14'b00000001111111 : 14'b00000011111111;
											assign node1351 = (inp[13]) ? node1355 : node1352;
												assign node1352 = (inp[8]) ? 14'b00000001111111 : 14'b00000011111111;
												assign node1355 = (inp[4]) ? 14'b00000000111111 : 14'b00000001111111;
										assign node1358 = (inp[7]) ? node1362 : node1359;
											assign node1359 = (inp[10]) ? 14'b00000011111111 : 14'b00000001111111;
											assign node1362 = (inp[13]) ? node1364 : 14'b00000000111111;
												assign node1364 = (inp[4]) ? 14'b00000000011111 : 14'b00000000111111;
							assign node1367 = (inp[4]) ? node1411 : node1368;
								assign node1368 = (inp[10]) ? node1386 : node1369;
									assign node1369 = (inp[8]) ? node1379 : node1370;
										assign node1370 = (inp[13]) ? node1376 : node1371;
											assign node1371 = (inp[6]) ? 14'b00000111111111 : node1372;
												assign node1372 = (inp[11]) ? 14'b00000111111111 : 14'b00001111111111;
											assign node1376 = (inp[11]) ? 14'b00000011111111 : 14'b00000111111111;
										assign node1379 = (inp[6]) ? node1381 : 14'b00000011111111;
											assign node1381 = (inp[12]) ? node1383 : 14'b00000001111111;
												assign node1383 = (inp[11]) ? 14'b00000001111111 : 14'b00000011111111;
									assign node1386 = (inp[12]) ? node1400 : node1387;
										assign node1387 = (inp[7]) ? node1393 : node1388;
											assign node1388 = (inp[13]) ? node1390 : 14'b00000011111111;
												assign node1390 = (inp[6]) ? 14'b00000001111111 : 14'b00000001111111;
											assign node1393 = (inp[11]) ? node1397 : node1394;
												assign node1394 = (inp[6]) ? 14'b00000011111111 : 14'b00000001111111;
												assign node1397 = (inp[8]) ? 14'b00000000111111 : 14'b00000001111111;
										assign node1400 = (inp[7]) ? node1406 : node1401;
											assign node1401 = (inp[8]) ? node1403 : 14'b00000001111111;
												assign node1403 = (inp[13]) ? 14'b00000000111111 : 14'b00000001111111;
											assign node1406 = (inp[11]) ? 14'b00000000111111 : node1407;
												assign node1407 = (inp[8]) ? 14'b00000000111111 : 14'b00000001111111;
								assign node1411 = (inp[13]) ? node1427 : node1412;
									assign node1412 = (inp[7]) ? 14'b00000000111111 : node1413;
										assign node1413 = (inp[12]) ? node1421 : node1414;
											assign node1414 = (inp[11]) ? node1418 : node1415;
												assign node1415 = (inp[8]) ? 14'b00000011111111 : 14'b00000011111111;
												assign node1418 = (inp[10]) ? 14'b00000001111111 : 14'b00000011111111;
											assign node1421 = (inp[6]) ? 14'b00000000111111 : node1422;
												assign node1422 = (inp[8]) ? 14'b00000001111111 : 14'b00000011111111;
									assign node1427 = (inp[6]) ? node1437 : node1428;
										assign node1428 = (inp[12]) ? node1434 : node1429;
											assign node1429 = (inp[10]) ? node1431 : 14'b00000011111111;
												assign node1431 = (inp[11]) ? 14'b00000000111111 : 14'b00000001111111;
											assign node1434 = (inp[10]) ? 14'b00000000111111 : 14'b00000000011111;
										assign node1437 = (inp[10]) ? node1441 : node1438;
											assign node1438 = (inp[11]) ? 14'b00000000111111 : 14'b00000000011111;
											assign node1441 = (inp[12]) ? node1445 : node1442;
												assign node1442 = (inp[7]) ? 14'b00000000011111 : 14'b00000000111111;
												assign node1445 = (inp[8]) ? 14'b00000000001111 : 14'b00000000011111;
						assign node1448 = (inp[6]) ? node1546 : node1449;
							assign node1449 = (inp[7]) ? node1499 : node1450;
								assign node1450 = (inp[12]) ? node1472 : node1451;
									assign node1451 = (inp[4]) ? node1465 : node1452;
										assign node1452 = (inp[10]) ? node1460 : node1453;
											assign node1453 = (inp[11]) ? node1457 : node1454;
												assign node1454 = (inp[8]) ? 14'b00000111111111 : 14'b00001111111111;
												assign node1457 = (inp[13]) ? 14'b00000011111111 : 14'b00000111111111;
											assign node1460 = (inp[0]) ? 14'b00000001111111 : node1461;
												assign node1461 = (inp[13]) ? 14'b00000011111111 : 14'b00000011111111;
										assign node1465 = (inp[13]) ? 14'b00000001111111 : node1466;
											assign node1466 = (inp[0]) ? 14'b00000001111111 : node1467;
												assign node1467 = (inp[11]) ? 14'b00000011111111 : 14'b00000111111111;
									assign node1472 = (inp[0]) ? node1488 : node1473;
										assign node1473 = (inp[11]) ? node1481 : node1474;
											assign node1474 = (inp[4]) ? node1478 : node1475;
												assign node1475 = (inp[13]) ? 14'b00000011111111 : 14'b00000011111111;
												assign node1478 = (inp[8]) ? 14'b00000001111111 : 14'b00000011111111;
											assign node1481 = (inp[13]) ? node1485 : node1482;
												assign node1482 = (inp[8]) ? 14'b00000001111111 : 14'b00000111111111;
												assign node1485 = (inp[10]) ? 14'b00000000011111 : 14'b00000001111111;
										assign node1488 = (inp[10]) ? node1494 : node1489;
											assign node1489 = (inp[4]) ? node1491 : 14'b00000001111111;
												assign node1491 = (inp[11]) ? 14'b00000000111111 : 14'b00000001111111;
											assign node1494 = (inp[4]) ? node1496 : 14'b00000000111111;
												assign node1496 = (inp[11]) ? 14'b00000000011111 : 14'b00000001111111;
								assign node1499 = (inp[11]) ? node1525 : node1500;
									assign node1500 = (inp[4]) ? node1510 : node1501;
										assign node1501 = (inp[8]) ? 14'b00000001111111 : node1502;
											assign node1502 = (inp[12]) ? node1506 : node1503;
												assign node1503 = (inp[10]) ? 14'b00000011111111 : 14'b00000111111111;
												assign node1506 = (inp[13]) ? 14'b00000001111111 : 14'b00000011111111;
										assign node1510 = (inp[12]) ? node1518 : node1511;
											assign node1511 = (inp[10]) ? node1515 : node1512;
												assign node1512 = (inp[0]) ? 14'b00000001111111 : 14'b00000011111111;
												assign node1515 = (inp[0]) ? 14'b00000000111111 : 14'b00000001111111;
											assign node1518 = (inp[13]) ? node1522 : node1519;
												assign node1519 = (inp[0]) ? 14'b00000000111111 : 14'b00000001111111;
												assign node1522 = (inp[10]) ? 14'b00000000011111 : 14'b00000000111111;
									assign node1525 = (inp[8]) ? node1537 : node1526;
										assign node1526 = (inp[10]) ? node1530 : node1527;
											assign node1527 = (inp[13]) ? 14'b00000001111111 : 14'b00000011111111;
											assign node1530 = (inp[0]) ? node1534 : node1531;
												assign node1531 = (inp[12]) ? 14'b00000000111111 : 14'b00000001111111;
												assign node1534 = (inp[12]) ? 14'b00000000011111 : 14'b00000000111111;
										assign node1537 = (inp[12]) ? node1543 : node1538;
											assign node1538 = (inp[13]) ? node1540 : 14'b00000000111111;
												assign node1540 = (inp[10]) ? 14'b00000000011111 : 14'b00000000111111;
											assign node1543 = (inp[13]) ? 14'b00000000011111 : 14'b00000000001111;
							assign node1546 = (inp[8]) ? node1602 : node1547;
								assign node1547 = (inp[12]) ? node1573 : node1548;
									assign node1548 = (inp[10]) ? node1562 : node1549;
										assign node1549 = (inp[4]) ? node1555 : node1550;
											assign node1550 = (inp[7]) ? 14'b00000011111111 : node1551;
												assign node1551 = (inp[11]) ? 14'b00000011111111 : 14'b00001111111111;
											assign node1555 = (inp[0]) ? node1559 : node1556;
												assign node1556 = (inp[13]) ? 14'b00000001111111 : 14'b00000011111111;
												assign node1559 = (inp[11]) ? 14'b00000000111111 : 14'b00000001111111;
										assign node1562 = (inp[13]) ? node1568 : node1563;
											assign node1563 = (inp[7]) ? node1565 : 14'b00000001111111;
												assign node1565 = (inp[0]) ? 14'b00000000111111 : 14'b00000001111111;
											assign node1568 = (inp[0]) ? node1570 : 14'b00000000111111;
												assign node1570 = (inp[11]) ? 14'b00000000111111 : 14'b00000001111111;
									assign node1573 = (inp[11]) ? node1589 : node1574;
										assign node1574 = (inp[13]) ? node1582 : node1575;
											assign node1575 = (inp[0]) ? node1579 : node1576;
												assign node1576 = (inp[7]) ? 14'b00000001111111 : 14'b00000011111111;
												assign node1579 = (inp[4]) ? 14'b00000000111111 : 14'b00000001111111;
											assign node1582 = (inp[4]) ? node1586 : node1583;
												assign node1583 = (inp[7]) ? 14'b00000000111111 : 14'b00000001111111;
												assign node1586 = (inp[0]) ? 14'b00000000011111 : 14'b00000000111111;
										assign node1589 = (inp[7]) ? node1595 : node1590;
											assign node1590 = (inp[4]) ? 14'b00000000111111 : node1591;
												assign node1591 = (inp[10]) ? 14'b00000000111111 : 14'b00000001111111;
											assign node1595 = (inp[4]) ? node1599 : node1596;
												assign node1596 = (inp[10]) ? 14'b00000000011111 : 14'b00000000111111;
												assign node1599 = (inp[13]) ? 14'b00000000001111 : 14'b00000000011111;
								assign node1602 = (inp[12]) ? node1624 : node1603;
									assign node1603 = (inp[0]) ? node1617 : node1604;
										assign node1604 = (inp[11]) ? node1610 : node1605;
											assign node1605 = (inp[7]) ? 14'b00000000111111 : node1606;
												assign node1606 = (inp[4]) ? 14'b00000011111111 : 14'b00000011111111;
											assign node1610 = (inp[13]) ? node1614 : node1611;
												assign node1611 = (inp[4]) ? 14'b00000000111111 : 14'b00000000111111;
												assign node1614 = (inp[10]) ? 14'b00000000011111 : 14'b00000000111111;
										assign node1617 = (inp[13]) ? node1619 : 14'b00000000111111;
											assign node1619 = (inp[10]) ? 14'b00000000001111 : node1620;
												assign node1620 = (inp[7]) ? 14'b00000000001111 : 14'b00000001111111;
									assign node1624 = (inp[13]) ? node1636 : node1625;
										assign node1625 = (inp[11]) ? node1631 : node1626;
											assign node1626 = (inp[7]) ? node1628 : 14'b00000000111111;
												assign node1628 = (inp[10]) ? 14'b00000000011111 : 14'b00000000111111;
											assign node1631 = (inp[10]) ? node1633 : 14'b00000000011111;
												assign node1633 = (inp[7]) ? 14'b00000000001111 : 14'b00000000011111;
										assign node1636 = (inp[10]) ? node1644 : node1637;
											assign node1637 = (inp[0]) ? node1641 : node1638;
												assign node1638 = (inp[11]) ? 14'b00000000011111 : 14'b00000000111111;
												assign node1641 = (inp[11]) ? 14'b00000000001111 : 14'b00000000011111;
											assign node1644 = (inp[0]) ? node1648 : node1645;
												assign node1645 = (inp[7]) ? 14'b00000000001111 : 14'b00000000001111;
												assign node1648 = (inp[7]) ? 14'b00000000000111 : 14'b00000000001111;
			assign node1651 = (inp[7]) ? node2433 : node1652;
				assign node1652 = (inp[9]) ? node2040 : node1653;
					assign node1653 = (inp[12]) ? node1849 : node1654;
						assign node1654 = (inp[2]) ? node1754 : node1655;
							assign node1655 = (inp[6]) ? node1703 : node1656;
								assign node1656 = (inp[13]) ? node1680 : node1657;
									assign node1657 = (inp[0]) ? node1669 : node1658;
										assign node1658 = (inp[3]) ? node1666 : node1659;
											assign node1659 = (inp[4]) ? node1663 : node1660;
												assign node1660 = (inp[10]) ? 14'b00011111111111 : 14'b00111111111111;
												assign node1663 = (inp[8]) ? 14'b00011111111111 : 14'b00011111111111;
											assign node1666 = (inp[4]) ? 14'b00011111111111 : 14'b00001111111111;
										assign node1669 = (inp[4]) ? node1675 : node1670;
											assign node1670 = (inp[3]) ? 14'b00001111111111 : node1671;
												assign node1671 = (inp[8]) ? 14'b00001111111111 : 14'b00011111111111;
											assign node1675 = (inp[10]) ? node1677 : 14'b00001111111111;
												assign node1677 = (inp[8]) ? 14'b00000011111111 : 14'b00000111111111;
									assign node1680 = (inp[4]) ? node1690 : node1681;
										assign node1681 = (inp[0]) ? node1687 : node1682;
											assign node1682 = (inp[3]) ? 14'b00001111111111 : node1683;
												assign node1683 = (inp[8]) ? 14'b00001111111111 : 14'b00011111111111;
											assign node1687 = (inp[11]) ? 14'b00000111111111 : 14'b00001111111111;
										assign node1690 = (inp[11]) ? node1696 : node1691;
											assign node1691 = (inp[0]) ? 14'b00000111111111 : node1692;
												assign node1692 = (inp[8]) ? 14'b00000111111111 : 14'b00001111111111;
											assign node1696 = (inp[10]) ? node1700 : node1697;
												assign node1697 = (inp[8]) ? 14'b00000011111111 : 14'b00000111111111;
												assign node1700 = (inp[8]) ? 14'b00000000111111 : 14'b00000011111111;
								assign node1703 = (inp[8]) ? node1733 : node1704;
									assign node1704 = (inp[0]) ? node1718 : node1705;
										assign node1705 = (inp[11]) ? node1713 : node1706;
											assign node1706 = (inp[13]) ? node1710 : node1707;
												assign node1707 = (inp[3]) ? 14'b00011111111111 : 14'b00011111111111;
												assign node1710 = (inp[3]) ? 14'b00000111111111 : 14'b00001111111111;
											assign node1713 = (inp[3]) ? node1715 : 14'b00000111111111;
												assign node1715 = (inp[13]) ? 14'b00000011111111 : 14'b00000111111111;
										assign node1718 = (inp[4]) ? node1726 : node1719;
											assign node1719 = (inp[10]) ? node1723 : node1720;
												assign node1720 = (inp[13]) ? 14'b00000111111111 : 14'b00001111111111;
												assign node1723 = (inp[13]) ? 14'b00000011111111 : 14'b00000111111111;
											assign node1726 = (inp[3]) ? node1730 : node1727;
												assign node1727 = (inp[13]) ? 14'b00000011111111 : 14'b00000111111111;
												assign node1730 = (inp[10]) ? 14'b00000001111111 : 14'b00000011111111;
									assign node1733 = (inp[10]) ? node1741 : node1734;
										assign node1734 = (inp[0]) ? node1736 : 14'b00000111111111;
											assign node1736 = (inp[4]) ? node1738 : 14'b00000111111111;
												assign node1738 = (inp[3]) ? 14'b00000011111111 : 14'b00000011111111;
										assign node1741 = (inp[4]) ? node1749 : node1742;
											assign node1742 = (inp[3]) ? node1746 : node1743;
												assign node1743 = (inp[13]) ? 14'b00000011111111 : 14'b00000111111111;
												assign node1746 = (inp[0]) ? 14'b00000001111111 : 14'b00000011111111;
											assign node1749 = (inp[11]) ? 14'b00000000111111 : node1750;
												assign node1750 = (inp[0]) ? 14'b00000001111111 : 14'b00000011111111;
							assign node1754 = (inp[11]) ? node1798 : node1755;
								assign node1755 = (inp[13]) ? node1777 : node1756;
									assign node1756 = (inp[0]) ? node1764 : node1757;
										assign node1757 = (inp[3]) ? 14'b00000111111111 : node1758;
											assign node1758 = (inp[4]) ? 14'b00000111111111 : node1759;
												assign node1759 = (inp[10]) ? 14'b00001111111111 : 14'b00011111111111;
										assign node1764 = (inp[4]) ? node1772 : node1765;
											assign node1765 = (inp[6]) ? node1769 : node1766;
												assign node1766 = (inp[10]) ? 14'b00000111111111 : 14'b00000111111111;
												assign node1769 = (inp[10]) ? 14'b00000011111111 : 14'b00000111111111;
											assign node1772 = (inp[6]) ? node1774 : 14'b00000111111111;
												assign node1774 = (inp[8]) ? 14'b00000001111111 : 14'b00000011111111;
									assign node1777 = (inp[8]) ? node1791 : node1778;
										assign node1778 = (inp[0]) ? node1784 : node1779;
											assign node1779 = (inp[4]) ? node1781 : 14'b00001111111111;
												assign node1781 = (inp[6]) ? 14'b00000011111111 : 14'b00000111111111;
											assign node1784 = (inp[6]) ? node1788 : node1785;
												assign node1785 = (inp[3]) ? 14'b00000011111111 : 14'b00000111111111;
												assign node1788 = (inp[4]) ? 14'b00000001111111 : 14'b00000011111111;
										assign node1791 = (inp[10]) ? node1793 : 14'b00000011111111;
											assign node1793 = (inp[3]) ? node1795 : 14'b00000001111111;
												assign node1795 = (inp[4]) ? 14'b00000000111111 : 14'b00000001111111;
								assign node1798 = (inp[13]) ? node1824 : node1799;
									assign node1799 = (inp[4]) ? node1809 : node1800;
										assign node1800 = (inp[6]) ? 14'b00000001111111 : node1801;
											assign node1801 = (inp[8]) ? node1805 : node1802;
												assign node1802 = (inp[0]) ? 14'b00000111111111 : 14'b00000111111111;
												assign node1805 = (inp[3]) ? 14'b00000011111111 : 14'b00000011111111;
										assign node1809 = (inp[10]) ? node1817 : node1810;
											assign node1810 = (inp[3]) ? node1814 : node1811;
												assign node1811 = (inp[8]) ? 14'b00000011111111 : 14'b00000111111111;
												assign node1814 = (inp[8]) ? 14'b00000001111111 : 14'b00000011111111;
											assign node1817 = (inp[0]) ? node1821 : node1818;
												assign node1818 = (inp[3]) ? 14'b00000001111111 : 14'b00000011111111;
												assign node1821 = (inp[6]) ? 14'b00000000111111 : 14'b00000001111111;
									assign node1824 = (inp[3]) ? node1838 : node1825;
										assign node1825 = (inp[10]) ? node1833 : node1826;
											assign node1826 = (inp[0]) ? node1830 : node1827;
												assign node1827 = (inp[8]) ? 14'b00000011111111 : 14'b00000111111111;
												assign node1830 = (inp[6]) ? 14'b00000011111111 : 14'b00000001111111;
											assign node1833 = (inp[4]) ? node1835 : 14'b00000001111111;
												assign node1835 = (inp[0]) ? 14'b00000000111111 : 14'b00000001111111;
										assign node1838 = (inp[6]) ? node1844 : node1839;
											assign node1839 = (inp[4]) ? node1841 : 14'b00000001111111;
												assign node1841 = (inp[8]) ? 14'b00000000111111 : 14'b00000001111111;
											assign node1844 = (inp[10]) ? node1846 : 14'b00000000111111;
												assign node1846 = (inp[0]) ? 14'b00000000011111 : 14'b00000000011111;
						assign node1849 = (inp[6]) ? node1945 : node1850;
							assign node1850 = (inp[3]) ? node1900 : node1851;
								assign node1851 = (inp[10]) ? node1875 : node1852;
									assign node1852 = (inp[0]) ? node1866 : node1853;
										assign node1853 = (inp[8]) ? node1859 : node1854;
											assign node1854 = (inp[13]) ? node1856 : 14'b00001111111111;
												assign node1856 = (inp[4]) ? 14'b00001111111111 : 14'b00011111111111;
											assign node1859 = (inp[11]) ? node1863 : node1860;
												assign node1860 = (inp[4]) ? 14'b00000111111111 : 14'b00001111111111;
												assign node1863 = (inp[4]) ? 14'b00000111111111 : 14'b00000011111111;
										assign node1866 = (inp[13]) ? 14'b00000011111111 : node1867;
											assign node1867 = (inp[11]) ? node1871 : node1868;
												assign node1868 = (inp[2]) ? 14'b00000111111111 : 14'b00001111111111;
												assign node1871 = (inp[8]) ? 14'b00000011111111 : 14'b00000111111111;
									assign node1875 = (inp[4]) ? node1891 : node1876;
										assign node1876 = (inp[0]) ? node1884 : node1877;
											assign node1877 = (inp[2]) ? node1881 : node1878;
												assign node1878 = (inp[11]) ? 14'b00000111111111 : 14'b00001111111111;
												assign node1881 = (inp[11]) ? 14'b00000011111111 : 14'b00000111111111;
											assign node1884 = (inp[13]) ? node1888 : node1885;
												assign node1885 = (inp[2]) ? 14'b00000011111111 : 14'b00000111111111;
												assign node1888 = (inp[11]) ? 14'b00000001111111 : 14'b00000011111111;
										assign node1891 = (inp[8]) ? node1897 : node1892;
											assign node1892 = (inp[11]) ? 14'b00000001111111 : node1893;
												assign node1893 = (inp[13]) ? 14'b00000011111111 : 14'b00000011111111;
											assign node1897 = (inp[2]) ? 14'b00000000111111 : 14'b00000001111111;
								assign node1900 = (inp[8]) ? node1926 : node1901;
									assign node1901 = (inp[2]) ? node1915 : node1902;
										assign node1902 = (inp[11]) ? node1908 : node1903;
											assign node1903 = (inp[13]) ? 14'b00000111111111 : node1904;
												assign node1904 = (inp[0]) ? 14'b00000111111111 : 14'b00001111111111;
											assign node1908 = (inp[0]) ? node1912 : node1909;
												assign node1909 = (inp[4]) ? 14'b00000011111111 : 14'b00000111111111;
												assign node1912 = (inp[10]) ? 14'b00000001111111 : 14'b00000011111111;
										assign node1915 = (inp[11]) ? node1923 : node1916;
											assign node1916 = (inp[0]) ? node1920 : node1917;
												assign node1917 = (inp[4]) ? 14'b00000011111111 : 14'b00000111111111;
												assign node1920 = (inp[10]) ? 14'b00000000111111 : 14'b00000011111111;
											assign node1923 = (inp[4]) ? 14'b00000000111111 : 14'b00000001111111;
									assign node1926 = (inp[4]) ? node1938 : node1927;
										assign node1927 = (inp[0]) ? node1933 : node1928;
											assign node1928 = (inp[2]) ? node1930 : 14'b00000011111111;
												assign node1930 = (inp[10]) ? 14'b00000001111111 : 14'b00000011111111;
											assign node1933 = (inp[2]) ? 14'b00000000011111 : node1934;
												assign node1934 = (inp[13]) ? 14'b00000001111111 : 14'b00000011111111;
										assign node1938 = (inp[10]) ? node1940 : 14'b00000001111111;
											assign node1940 = (inp[13]) ? 14'b00000000111111 : node1941;
												assign node1941 = (inp[11]) ? 14'b00000000111111 : 14'b00000001111111;
							assign node1945 = (inp[10]) ? node1989 : node1946;
								assign node1946 = (inp[13]) ? node1966 : node1947;
									assign node1947 = (inp[2]) ? node1959 : node1948;
										assign node1948 = (inp[8]) ? node1954 : node1949;
											assign node1949 = (inp[11]) ? node1951 : 14'b00000111111111;
												assign node1951 = (inp[0]) ? 14'b00000011111111 : 14'b00000111111111;
											assign node1954 = (inp[3]) ? 14'b00000001111111 : node1955;
												assign node1955 = (inp[0]) ? 14'b00000011111111 : 14'b00000111111111;
										assign node1959 = (inp[0]) ? 14'b00000001111111 : node1960;
											assign node1960 = (inp[8]) ? node1962 : 14'b00000011111111;
												assign node1962 = (inp[11]) ? 14'b00000001111111 : 14'b00000011111111;
									assign node1966 = (inp[3]) ? node1982 : node1967;
										assign node1967 = (inp[8]) ? node1975 : node1968;
											assign node1968 = (inp[11]) ? node1972 : node1969;
												assign node1969 = (inp[0]) ? 14'b00000111111111 : 14'b00001111111111;
												assign node1972 = (inp[4]) ? 14'b00000001111111 : 14'b00000011111111;
											assign node1975 = (inp[2]) ? node1979 : node1976;
												assign node1976 = (inp[11]) ? 14'b00000001111111 : 14'b00000011111111;
												assign node1979 = (inp[11]) ? 14'b00000000111111 : 14'b00000001111111;
										assign node1982 = (inp[4]) ? 14'b00000000111111 : node1983;
											assign node1983 = (inp[8]) ? node1985 : 14'b00000001111111;
												assign node1985 = (inp[2]) ? 14'b00000000111111 : 14'b00000001111111;
								assign node1989 = (inp[0]) ? node2017 : node1990;
									assign node1990 = (inp[3]) ? node2004 : node1991;
										assign node1991 = (inp[8]) ? node1999 : node1992;
											assign node1992 = (inp[4]) ? node1996 : node1993;
												assign node1993 = (inp[11]) ? 14'b00000011111111 : 14'b00000111111111;
												assign node1996 = (inp[11]) ? 14'b00000001111111 : 14'b00000011111111;
											assign node1999 = (inp[13]) ? 14'b00000001111111 : node2000;
												assign node2000 = (inp[11]) ? 14'b00000001111111 : 14'b00000011111111;
										assign node2004 = (inp[11]) ? node2010 : node2005;
											assign node2005 = (inp[13]) ? 14'b00000000111111 : node2006;
												assign node2006 = (inp[4]) ? 14'b00000001111111 : 14'b00000011111111;
											assign node2010 = (inp[4]) ? node2014 : node2011;
												assign node2011 = (inp[13]) ? 14'b00000000111111 : 14'b00000001111111;
												assign node2014 = (inp[2]) ? 14'b00000000011111 : 14'b00000000111111;
									assign node2017 = (inp[4]) ? node2027 : node2018;
										assign node2018 = (inp[11]) ? 14'b00000000111111 : node2019;
											assign node2019 = (inp[8]) ? node2023 : node2020;
												assign node2020 = (inp[2]) ? 14'b00000000111111 : 14'b00000011111111;
												assign node2023 = (inp[3]) ? 14'b00000000111111 : 14'b00000001111111;
										assign node2027 = (inp[8]) ? node2033 : node2028;
											assign node2028 = (inp[11]) ? node2030 : 14'b00000000111111;
												assign node2030 = (inp[2]) ? 14'b00000000011111 : 14'b00000000111111;
											assign node2033 = (inp[13]) ? node2037 : node2034;
												assign node2034 = (inp[3]) ? 14'b00000000011111 : 14'b00000000011111;
												assign node2037 = (inp[3]) ? 14'b00000000001111 : 14'b00000000011111;
					assign node2040 = (inp[13]) ? node2232 : node2041;
						assign node2041 = (inp[0]) ? node2143 : node2042;
							assign node2042 = (inp[6]) ? node2092 : node2043;
								assign node2043 = (inp[4]) ? node2069 : node2044;
									assign node2044 = (inp[10]) ? node2058 : node2045;
										assign node2045 = (inp[2]) ? node2051 : node2046;
											assign node2046 = (inp[11]) ? 14'b00001111111111 : node2047;
												assign node2047 = (inp[3]) ? 14'b00001111111111 : 14'b00011111111111;
											assign node2051 = (inp[11]) ? node2055 : node2052;
												assign node2052 = (inp[3]) ? 14'b00000111111111 : 14'b00001111111111;
												assign node2055 = (inp[3]) ? 14'b00000011111111 : 14'b00000111111111;
										assign node2058 = (inp[3]) ? node2066 : node2059;
											assign node2059 = (inp[2]) ? node2063 : node2060;
												assign node2060 = (inp[12]) ? 14'b00000111111111 : 14'b00001111111111;
												assign node2063 = (inp[11]) ? 14'b00000011111111 : 14'b00000111111111;
											assign node2066 = (inp[12]) ? 14'b00000001111111 : 14'b00000011111111;
									assign node2069 = (inp[2]) ? node2077 : node2070;
										assign node2070 = (inp[3]) ? 14'b00000111111111 : node2071;
											assign node2071 = (inp[10]) ? 14'b00000011111111 : node2072;
												assign node2072 = (inp[8]) ? 14'b00000011111111 : 14'b00000111111111;
										assign node2077 = (inp[12]) ? node2085 : node2078;
											assign node2078 = (inp[10]) ? node2082 : node2079;
												assign node2079 = (inp[8]) ? 14'b00000011111111 : 14'b00000011111111;
												assign node2082 = (inp[11]) ? 14'b00000001111111 : 14'b00000011111111;
											assign node2085 = (inp[11]) ? node2089 : node2086;
												assign node2086 = (inp[3]) ? 14'b00000001111111 : 14'b00000111111111;
												assign node2089 = (inp[3]) ? 14'b00000000111111 : 14'b00000001111111;
								assign node2092 = (inp[3]) ? node2116 : node2093;
									assign node2093 = (inp[8]) ? node2109 : node2094;
										assign node2094 = (inp[4]) ? node2102 : node2095;
											assign node2095 = (inp[10]) ? node2099 : node2096;
												assign node2096 = (inp[11]) ? 14'b00001111111111 : 14'b00011111111111;
												assign node2099 = (inp[2]) ? 14'b00000011111111 : 14'b00000111111111;
											assign node2102 = (inp[10]) ? node2106 : node2103;
												assign node2103 = (inp[2]) ? 14'b00000011111111 : 14'b00000111111111;
												assign node2106 = (inp[12]) ? 14'b00000001111111 : 14'b00000011111111;
										assign node2109 = (inp[11]) ? node2111 : 14'b00000011111111;
											assign node2111 = (inp[4]) ? 14'b00000001111111 : node2112;
												assign node2112 = (inp[12]) ? 14'b00000001111111 : 14'b00000011111111;
									assign node2116 = (inp[12]) ? node2130 : node2117;
										assign node2117 = (inp[10]) ? node2125 : node2118;
											assign node2118 = (inp[4]) ? node2122 : node2119;
												assign node2119 = (inp[2]) ? 14'b00000011111111 : 14'b00000111111111;
												assign node2122 = (inp[2]) ? 14'b00000001111111 : 14'b00000011111111;
											assign node2125 = (inp[8]) ? 14'b00000000111111 : node2126;
												assign node2126 = (inp[4]) ? 14'b00000001111111 : 14'b00000011111111;
										assign node2130 = (inp[10]) ? node2138 : node2131;
											assign node2131 = (inp[11]) ? node2135 : node2132;
												assign node2132 = (inp[4]) ? 14'b00000001111111 : 14'b00000011111111;
												assign node2135 = (inp[4]) ? 14'b00000000111111 : 14'b00000001111111;
											assign node2138 = (inp[4]) ? 14'b00000000011111 : node2139;
												assign node2139 = (inp[8]) ? 14'b00000000111111 : 14'b00000001111111;
							assign node2143 = (inp[8]) ? node2179 : node2144;
								assign node2144 = (inp[6]) ? node2156 : node2145;
									assign node2145 = (inp[2]) ? node2147 : 14'b00000011111111;
										assign node2147 = (inp[12]) ? node2151 : node2148;
											assign node2148 = (inp[11]) ? 14'b00000011111111 : 14'b00000111111111;
											assign node2151 = (inp[4]) ? 14'b00000001111111 : node2152;
												assign node2152 = (inp[11]) ? 14'b00000001111111 : 14'b00000011111111;
									assign node2156 = (inp[3]) ? node2166 : node2157;
										assign node2157 = (inp[10]) ? 14'b00000001111111 : node2158;
											assign node2158 = (inp[12]) ? node2162 : node2159;
												assign node2159 = (inp[11]) ? 14'b00000011111111 : 14'b00000111111111;
												assign node2162 = (inp[4]) ? 14'b00000001111111 : 14'b00000011111111;
										assign node2166 = (inp[12]) ? node2174 : node2167;
											assign node2167 = (inp[4]) ? node2171 : node2168;
												assign node2168 = (inp[10]) ? 14'b00000001111111 : 14'b00000011111111;
												assign node2171 = (inp[2]) ? 14'b00000000111111 : 14'b00000001111111;
											assign node2174 = (inp[11]) ? 14'b00000000011111 : node2175;
												assign node2175 = (inp[2]) ? 14'b00000000111111 : 14'b00000000111111;
								assign node2179 = (inp[2]) ? node2209 : node2180;
									assign node2180 = (inp[4]) ? node2196 : node2181;
										assign node2181 = (inp[12]) ? node2189 : node2182;
											assign node2182 = (inp[11]) ? node2186 : node2183;
												assign node2183 = (inp[6]) ? 14'b00000001111111 : 14'b00000111111111;
												assign node2186 = (inp[3]) ? 14'b00000001111111 : 14'b00000011111111;
											assign node2189 = (inp[11]) ? node2193 : node2190;
												assign node2190 = (inp[10]) ? 14'b00000001111111 : 14'b00000011111111;
												assign node2193 = (inp[3]) ? 14'b00000000111111 : 14'b00000001111111;
										assign node2196 = (inp[10]) ? node2202 : node2197;
											assign node2197 = (inp[3]) ? node2199 : 14'b00000001111111;
												assign node2199 = (inp[6]) ? 14'b00000000111111 : 14'b00000001111111;
											assign node2202 = (inp[11]) ? node2206 : node2203;
												assign node2203 = (inp[3]) ? 14'b00000000111111 : 14'b00000011111111;
												assign node2206 = (inp[6]) ? 14'b00000000011111 : 14'b00000000111111;
									assign node2209 = (inp[3]) ? node2221 : node2210;
										assign node2210 = (inp[4]) ? node2216 : node2211;
											assign node2211 = (inp[6]) ? 14'b00000000111111 : node2212;
												assign node2212 = (inp[10]) ? 14'b00000001111111 : 14'b00000011111111;
											assign node2216 = (inp[10]) ? 14'b00000000011111 : node2217;
												assign node2217 = (inp[12]) ? 14'b00000000111111 : 14'b00000000111111;
										assign node2221 = (inp[11]) ? node2227 : node2222;
											assign node2222 = (inp[6]) ? node2224 : 14'b00000001111111;
												assign node2224 = (inp[12]) ? 14'b00000000011111 : 14'b00000000111111;
											assign node2227 = (inp[12]) ? 14'b00000000011111 : node2228;
												assign node2228 = (inp[6]) ? 14'b00000000011111 : 14'b00000000111111;
						assign node2232 = (inp[4]) ? node2344 : node2233;
							assign node2233 = (inp[2]) ? node2287 : node2234;
								assign node2234 = (inp[10]) ? node2258 : node2235;
									assign node2235 = (inp[3]) ? node2245 : node2236;
										assign node2236 = (inp[6]) ? node2240 : node2237;
											assign node2237 = (inp[11]) ? 14'b00000111111111 : 14'b00001111111111;
											assign node2240 = (inp[8]) ? 14'b00000011111111 : node2241;
												assign node2241 = (inp[12]) ? 14'b00000011111111 : 14'b00000111111111;
										assign node2245 = (inp[12]) ? node2253 : node2246;
											assign node2246 = (inp[8]) ? node2250 : node2247;
												assign node2247 = (inp[0]) ? 14'b00000011111111 : 14'b00000111111111;
												assign node2250 = (inp[0]) ? 14'b00000001111111 : 14'b00000011111111;
											assign node2253 = (inp[8]) ? node2255 : 14'b00000001111111;
												assign node2255 = (inp[6]) ? 14'b00000001111111 : 14'b00000011111111;
									assign node2258 = (inp[0]) ? node2274 : node2259;
										assign node2259 = (inp[6]) ? node2267 : node2260;
											assign node2260 = (inp[11]) ? node2264 : node2261;
												assign node2261 = (inp[12]) ? 14'b00000001111111 : 14'b00000111111111;
												assign node2264 = (inp[8]) ? 14'b00000001111111 : 14'b00000011111111;
											assign node2267 = (inp[8]) ? node2271 : node2268;
												assign node2268 = (inp[3]) ? 14'b00000000111111 : 14'b00000011111111;
												assign node2271 = (inp[11]) ? 14'b00000000111111 : 14'b00000001111111;
										assign node2274 = (inp[12]) ? node2282 : node2275;
											assign node2275 = (inp[11]) ? node2279 : node2276;
												assign node2276 = (inp[6]) ? 14'b00000011111111 : 14'b00000001111111;
												assign node2279 = (inp[3]) ? 14'b00000000111111 : 14'b00000001111111;
											assign node2282 = (inp[8]) ? node2284 : 14'b00000001111111;
												assign node2284 = (inp[11]) ? 14'b00000000011111 : 14'b00000000111111;
								assign node2287 = (inp[3]) ? node2317 : node2288;
									assign node2288 = (inp[11]) ? node2302 : node2289;
										assign node2289 = (inp[6]) ? node2295 : node2290;
											assign node2290 = (inp[12]) ? 14'b00000011111111 : node2291;
												assign node2291 = (inp[0]) ? 14'b00000011111111 : 14'b00000111111111;
											assign node2295 = (inp[0]) ? node2299 : node2296;
												assign node2296 = (inp[8]) ? 14'b00000001111111 : 14'b00000011111111;
												assign node2299 = (inp[12]) ? 14'b00000000011111 : 14'b00000001111111;
										assign node2302 = (inp[10]) ? node2310 : node2303;
											assign node2303 = (inp[12]) ? node2307 : node2304;
												assign node2304 = (inp[0]) ? 14'b00000001111111 : 14'b00000001111111;
												assign node2307 = (inp[6]) ? 14'b00000001111111 : 14'b00000001111111;
											assign node2310 = (inp[0]) ? node2314 : node2311;
												assign node2311 = (inp[6]) ? 14'b00000000111111 : 14'b00000001111111;
												assign node2314 = (inp[6]) ? 14'b00000000011111 : 14'b00000000111111;
									assign node2317 = (inp[6]) ? node2333 : node2318;
										assign node2318 = (inp[8]) ? node2326 : node2319;
											assign node2319 = (inp[11]) ? node2323 : node2320;
												assign node2320 = (inp[10]) ? 14'b00000001111111 : 14'b00000011111111;
												assign node2323 = (inp[0]) ? 14'b00000000111111 : 14'b00000001111111;
											assign node2326 = (inp[10]) ? node2330 : node2327;
												assign node2327 = (inp[12]) ? 14'b00000000111111 : 14'b00000001111111;
												assign node2330 = (inp[12]) ? 14'b00000000011111 : 14'b00000000111111;
										assign node2333 = (inp[10]) ? node2339 : node2334;
											assign node2334 = (inp[0]) ? node2336 : 14'b00000000111111;
												assign node2336 = (inp[11]) ? 14'b00000000011111 : 14'b00000000111111;
											assign node2339 = (inp[11]) ? node2341 : 14'b00000000011111;
												assign node2341 = (inp[12]) ? 14'b00000000001111 : 14'b00000000011111;
							assign node2344 = (inp[2]) ? node2382 : node2345;
								assign node2345 = (inp[10]) ? node2363 : node2346;
									assign node2346 = (inp[6]) ? node2358 : node2347;
										assign node2347 = (inp[0]) ? node2353 : node2348;
											assign node2348 = (inp[11]) ? node2350 : 14'b00000111111111;
												assign node2350 = (inp[12]) ? 14'b00000001111111 : 14'b00000011111111;
											assign node2353 = (inp[11]) ? 14'b00000000111111 : node2354;
												assign node2354 = (inp[8]) ? 14'b00000001111111 : 14'b00000011111111;
										assign node2358 = (inp[0]) ? 14'b00000000111111 : node2359;
											assign node2359 = (inp[8]) ? 14'b00000000111111 : 14'b00000001111111;
									assign node2363 = (inp[3]) ? node2375 : node2364;
										assign node2364 = (inp[0]) ? node2370 : node2365;
											assign node2365 = (inp[11]) ? node2367 : 14'b00000011111111;
												assign node2367 = (inp[6]) ? 14'b00000000111111 : 14'b00000001111111;
											assign node2370 = (inp[11]) ? node2372 : 14'b00000000111111;
												assign node2372 = (inp[6]) ? 14'b00000000011111 : 14'b00000000111111;
										assign node2375 = (inp[11]) ? 14'b00000000011111 : node2376;
											assign node2376 = (inp[8]) ? node2378 : 14'b00000000111111;
												assign node2378 = (inp[6]) ? 14'b00000000001111 : 14'b00000000011111;
								assign node2382 = (inp[12]) ? node2406 : node2383;
									assign node2383 = (inp[8]) ? node2393 : node2384;
										assign node2384 = (inp[0]) ? node2388 : node2385;
											assign node2385 = (inp[11]) ? 14'b00000000111111 : 14'b00000001111111;
											assign node2388 = (inp[10]) ? 14'b00000000011111 : node2389;
												assign node2389 = (inp[3]) ? 14'b00000000111111 : 14'b00000000111111;
										assign node2393 = (inp[0]) ? node2401 : node2394;
											assign node2394 = (inp[10]) ? node2398 : node2395;
												assign node2395 = (inp[11]) ? 14'b00000000111111 : 14'b00000001111111;
												assign node2398 = (inp[11]) ? 14'b00000000011111 : 14'b00000000011111;
											assign node2401 = (inp[11]) ? node2403 : 14'b00000000011111;
												assign node2403 = (inp[3]) ? 14'b00000000001111 : 14'b00000000011111;
									assign node2406 = (inp[11]) ? node2420 : node2407;
										assign node2407 = (inp[6]) ? node2413 : node2408;
											assign node2408 = (inp[3]) ? node2410 : 14'b00000000111111;
												assign node2410 = (inp[10]) ? 14'b00000000011111 : 14'b00000000011111;
											assign node2413 = (inp[3]) ? node2417 : node2414;
												assign node2414 = (inp[10]) ? 14'b00000000011111 : 14'b00000000111111;
												assign node2417 = (inp[10]) ? 14'b00000000001111 : 14'b00000000011111;
										assign node2420 = (inp[3]) ? node2426 : node2421;
											assign node2421 = (inp[8]) ? node2423 : 14'b00000000011111;
												assign node2423 = (inp[0]) ? 14'b00000000001111 : 14'b00000000011111;
											assign node2426 = (inp[10]) ? node2430 : node2427;
												assign node2427 = (inp[0]) ? 14'b00000000001111 : 14'b00000000011111;
												assign node2430 = (inp[6]) ? 14'b00000000000111 : 14'b00000000001111;
				assign node2433 = (inp[0]) ? node2813 : node2434;
					assign node2434 = (inp[11]) ? node2620 : node2435;
						assign node2435 = (inp[13]) ? node2525 : node2436;
							assign node2436 = (inp[3]) ? node2482 : node2437;
								assign node2437 = (inp[4]) ? node2461 : node2438;
									assign node2438 = (inp[12]) ? node2448 : node2439;
										assign node2439 = (inp[10]) ? node2443 : node2440;
											assign node2440 = (inp[8]) ? 14'b00001111111111 : 14'b00011111111111;
											assign node2443 = (inp[9]) ? node2445 : 14'b00001111111111;
												assign node2445 = (inp[2]) ? 14'b00000111111111 : 14'b00001111111111;
										assign node2448 = (inp[6]) ? node2454 : node2449;
											assign node2449 = (inp[10]) ? 14'b00000111111111 : node2450;
												assign node2450 = (inp[8]) ? 14'b00001111111111 : 14'b00011111111111;
											assign node2454 = (inp[8]) ? node2458 : node2455;
												assign node2455 = (inp[2]) ? 14'b00000011111111 : 14'b00000111111111;
												assign node2458 = (inp[2]) ? 14'b00000001111111 : 14'b00000011111111;
									assign node2461 = (inp[10]) ? node2467 : node2462;
										assign node2462 = (inp[2]) ? node2464 : 14'b00000111111111;
											assign node2464 = (inp[9]) ? 14'b00000011111111 : 14'b00000111111111;
										assign node2467 = (inp[2]) ? node2475 : node2468;
											assign node2468 = (inp[9]) ? node2472 : node2469;
												assign node2469 = (inp[12]) ? 14'b00000011111111 : 14'b00000011111111;
												assign node2472 = (inp[6]) ? 14'b00000001111111 : 14'b00000011111111;
											assign node2475 = (inp[6]) ? node2479 : node2476;
												assign node2476 = (inp[8]) ? 14'b00000001111111 : 14'b00000011111111;
												assign node2479 = (inp[12]) ? 14'b00000000111111 : 14'b00000001111111;
								assign node2482 = (inp[6]) ? node2504 : node2483;
									assign node2483 = (inp[12]) ? node2491 : node2484;
										assign node2484 = (inp[9]) ? node2486 : 14'b00000111111111;
											assign node2486 = (inp[4]) ? 14'b00000011111111 : node2487;
												assign node2487 = (inp[2]) ? 14'b00000011111111 : 14'b00000111111111;
										assign node2491 = (inp[9]) ? node2497 : node2492;
											assign node2492 = (inp[8]) ? 14'b00000001111111 : node2493;
												assign node2493 = (inp[2]) ? 14'b00000011111111 : 14'b00000111111111;
											assign node2497 = (inp[10]) ? node2501 : node2498;
												assign node2498 = (inp[2]) ? 14'b00000001111111 : 14'b00000011111111;
												assign node2501 = (inp[8]) ? 14'b00000000111111 : 14'b00000001111111;
									assign node2504 = (inp[4]) ? node2516 : node2505;
										assign node2505 = (inp[10]) ? node2511 : node2506;
											assign node2506 = (inp[8]) ? node2508 : 14'b00000011111111;
												assign node2508 = (inp[9]) ? 14'b00000001111111 : 14'b00000011111111;
											assign node2511 = (inp[12]) ? 14'b00000001111111 : node2512;
												assign node2512 = (inp[8]) ? 14'b00000001111111 : 14'b00000011111111;
										assign node2516 = (inp[12]) ? node2522 : node2517;
											assign node2517 = (inp[10]) ? node2519 : 14'b00000011111111;
												assign node2519 = (inp[9]) ? 14'b00000000111111 : 14'b00000001111111;
											assign node2522 = (inp[2]) ? 14'b00000000111111 : 14'b00000001111111;
							assign node2525 = (inp[9]) ? node2571 : node2526;
								assign node2526 = (inp[10]) ? node2546 : node2527;
									assign node2527 = (inp[12]) ? node2535 : node2528;
										assign node2528 = (inp[3]) ? 14'b00000011111111 : node2529;
											assign node2529 = (inp[4]) ? 14'b00000111111111 : node2530;
												assign node2530 = (inp[8]) ? 14'b00000111111111 : 14'b00001111111111;
										assign node2535 = (inp[6]) ? node2541 : node2536;
											assign node2536 = (inp[2]) ? 14'b00000001111111 : node2537;
												assign node2537 = (inp[3]) ? 14'b00000011111111 : 14'b00000011111111;
											assign node2541 = (inp[4]) ? 14'b00000000111111 : node2542;
												assign node2542 = (inp[3]) ? 14'b00000001111111 : 14'b00000011111111;
									assign node2546 = (inp[6]) ? node2558 : node2547;
										assign node2547 = (inp[8]) ? node2555 : node2548;
											assign node2548 = (inp[2]) ? node2552 : node2549;
												assign node2549 = (inp[4]) ? 14'b00000011111111 : 14'b00000111111111;
												assign node2552 = (inp[12]) ? 14'b00000001111111 : 14'b00000011111111;
											assign node2555 = (inp[3]) ? 14'b00000001111111 : 14'b00000011111111;
										assign node2558 = (inp[8]) ? node2566 : node2559;
											assign node2559 = (inp[2]) ? node2563 : node2560;
												assign node2560 = (inp[4]) ? 14'b00000001111111 : 14'b00000011111111;
												assign node2563 = (inp[4]) ? 14'b00000000111111 : 14'b00000001111111;
											assign node2566 = (inp[2]) ? 14'b00000000011111 : node2567;
												assign node2567 = (inp[4]) ? 14'b00000000111111 : 14'b00000001111111;
								assign node2571 = (inp[4]) ? node2601 : node2572;
									assign node2572 = (inp[3]) ? node2586 : node2573;
										assign node2573 = (inp[6]) ? node2579 : node2574;
											assign node2574 = (inp[2]) ? node2576 : 14'b00000111111111;
												assign node2576 = (inp[8]) ? 14'b00000001111111 : 14'b00000111111111;
											assign node2579 = (inp[2]) ? node2583 : node2580;
												assign node2580 = (inp[12]) ? 14'b00000001111111 : 14'b00000011111111;
												assign node2583 = (inp[8]) ? 14'b00000000111111 : 14'b00000001111111;
										assign node2586 = (inp[6]) ? node2594 : node2587;
											assign node2587 = (inp[10]) ? node2591 : node2588;
												assign node2588 = (inp[8]) ? 14'b00000001111111 : 14'b00000001111111;
												assign node2591 = (inp[2]) ? 14'b00000000111111 : 14'b00000001111111;
											assign node2594 = (inp[12]) ? node2598 : node2595;
												assign node2595 = (inp[8]) ? 14'b00000000111111 : 14'b00000001111111;
												assign node2598 = (inp[8]) ? 14'b00000000011111 : 14'b00000000011111;
									assign node2601 = (inp[10]) ? node2615 : node2602;
										assign node2602 = (inp[2]) ? node2608 : node2603;
											assign node2603 = (inp[6]) ? node2605 : 14'b00000011111111;
												assign node2605 = (inp[3]) ? 14'b00000000111111 : 14'b00000001111111;
											assign node2608 = (inp[12]) ? node2612 : node2609;
												assign node2609 = (inp[6]) ? 14'b00000000111111 : 14'b00000001111111;
												assign node2612 = (inp[8]) ? 14'b00000000011111 : 14'b00000000111111;
										assign node2615 = (inp[12]) ? 14'b00000000011111 : node2616;
											assign node2616 = (inp[8]) ? 14'b00000000011111 : 14'b00000000111111;
						assign node2620 = (inp[12]) ? node2718 : node2621;
							assign node2621 = (inp[4]) ? node2669 : node2622;
								assign node2622 = (inp[9]) ? node2646 : node2623;
									assign node2623 = (inp[3]) ? node2635 : node2624;
										assign node2624 = (inp[13]) ? node2630 : node2625;
											assign node2625 = (inp[10]) ? node2627 : 14'b00000111111111;
												assign node2627 = (inp[8]) ? 14'b00000111111111 : 14'b00001111111111;
											assign node2630 = (inp[6]) ? 14'b00000011111111 : node2631;
												assign node2631 = (inp[10]) ? 14'b00000011111111 : 14'b00000111111111;
										assign node2635 = (inp[6]) ? node2641 : node2636;
											assign node2636 = (inp[10]) ? node2638 : 14'b00000111111111;
												assign node2638 = (inp[2]) ? 14'b00000000111111 : 14'b00000011111111;
											assign node2641 = (inp[2]) ? 14'b00000001111111 : node2642;
												assign node2642 = (inp[10]) ? 14'b00000001111111 : 14'b00000011111111;
									assign node2646 = (inp[10]) ? node2660 : node2647;
										assign node2647 = (inp[6]) ? node2653 : node2648;
											assign node2648 = (inp[3]) ? node2650 : 14'b00000011111111;
												assign node2650 = (inp[2]) ? 14'b00000001111111 : 14'b00000011111111;
											assign node2653 = (inp[2]) ? node2657 : node2654;
												assign node2654 = (inp[3]) ? 14'b00000001111111 : 14'b00000011111111;
												assign node2657 = (inp[8]) ? 14'b00000000111111 : 14'b00000001111111;
										assign node2660 = (inp[13]) ? 14'b00000000111111 : node2661;
											assign node2661 = (inp[3]) ? node2665 : node2662;
												assign node2662 = (inp[2]) ? 14'b00000000111111 : 14'b00000011111111;
												assign node2665 = (inp[6]) ? 14'b00000000111111 : 14'b00000001111111;
								assign node2669 = (inp[2]) ? node2693 : node2670;
									assign node2670 = (inp[6]) ? node2686 : node2671;
										assign node2671 = (inp[8]) ? node2679 : node2672;
											assign node2672 = (inp[9]) ? node2676 : node2673;
												assign node2673 = (inp[13]) ? 14'b00000011111111 : 14'b00001111111111;
												assign node2676 = (inp[13]) ? 14'b00000001111111 : 14'b00000001111111;
											assign node2679 = (inp[13]) ? node2683 : node2680;
												assign node2680 = (inp[10]) ? 14'b00000001111111 : 14'b00000011111111;
												assign node2683 = (inp[10]) ? 14'b00000000111111 : 14'b00000001111111;
										assign node2686 = (inp[13]) ? node2688 : 14'b00000001111111;
											assign node2688 = (inp[10]) ? 14'b00000000111111 : node2689;
												assign node2689 = (inp[3]) ? 14'b00000000111111 : 14'b00000001111111;
									assign node2693 = (inp[9]) ? node2707 : node2694;
										assign node2694 = (inp[6]) ? node2702 : node2695;
											assign node2695 = (inp[13]) ? node2699 : node2696;
												assign node2696 = (inp[10]) ? 14'b00000001111111 : 14'b00000111111111;
												assign node2699 = (inp[10]) ? 14'b00000000111111 : 14'b00000001111111;
											assign node2702 = (inp[8]) ? 14'b00000000111111 : node2703;
												assign node2703 = (inp[13]) ? 14'b00000001111111 : 14'b00000000111111;
										assign node2707 = (inp[10]) ? node2713 : node2708;
											assign node2708 = (inp[8]) ? node2710 : 14'b00000000111111;
												assign node2710 = (inp[6]) ? 14'b00000000011111 : 14'b00000000111111;
											assign node2713 = (inp[13]) ? node2715 : 14'b00000000011111;
												assign node2715 = (inp[8]) ? 14'b00000000000111 : 14'b00000000001111;
							assign node2718 = (inp[6]) ? node2764 : node2719;
								assign node2719 = (inp[10]) ? node2739 : node2720;
									assign node2720 = (inp[4]) ? node2728 : node2721;
										assign node2721 = (inp[13]) ? 14'b00000001111111 : node2722;
											assign node2722 = (inp[8]) ? 14'b00000011111111 : node2723;
												assign node2723 = (inp[9]) ? 14'b00000011111111 : 14'b00000111111111;
										assign node2728 = (inp[9]) ? node2734 : node2729;
											assign node2729 = (inp[2]) ? 14'b00000001111111 : node2730;
												assign node2730 = (inp[3]) ? 14'b00000001111111 : 14'b00000011111111;
											assign node2734 = (inp[13]) ? 14'b00000001111111 : node2735;
												assign node2735 = (inp[8]) ? 14'b00000000011111 : 14'b00000000111111;
									assign node2739 = (inp[8]) ? node2753 : node2740;
										assign node2740 = (inp[2]) ? node2748 : node2741;
											assign node2741 = (inp[3]) ? node2745 : node2742;
												assign node2742 = (inp[4]) ? 14'b00000001111111 : 14'b00000001111111;
												assign node2745 = (inp[9]) ? 14'b00000000111111 : 14'b00000000111111;
											assign node2748 = (inp[9]) ? node2750 : 14'b00000000111111;
												assign node2750 = (inp[4]) ? 14'b00000000011111 : 14'b00000000111111;
										assign node2753 = (inp[13]) ? node2759 : node2754;
											assign node2754 = (inp[2]) ? node2756 : 14'b00000011111111;
												assign node2756 = (inp[3]) ? 14'b00000000011111 : 14'b00000000111111;
											assign node2759 = (inp[2]) ? node2761 : 14'b00000000011111;
												assign node2761 = (inp[3]) ? 14'b00000000000111 : 14'b00000000011111;
								assign node2764 = (inp[9]) ? node2792 : node2765;
									assign node2765 = (inp[10]) ? node2779 : node2766;
										assign node2766 = (inp[8]) ? node2772 : node2767;
											assign node2767 = (inp[13]) ? node2769 : 14'b00000111111111;
												assign node2769 = (inp[3]) ? 14'b00000000111111 : 14'b00000001111111;
											assign node2772 = (inp[13]) ? node2776 : node2773;
												assign node2773 = (inp[3]) ? 14'b00000000111111 : 14'b00000001111111;
												assign node2776 = (inp[4]) ? 14'b00000000011111 : 14'b00000000111111;
										assign node2779 = (inp[2]) ? node2785 : node2780;
											assign node2780 = (inp[4]) ? 14'b00000000011111 : node2781;
												assign node2781 = (inp[13]) ? 14'b00000000111111 : 14'b00000000111111;
											assign node2785 = (inp[3]) ? node2789 : node2786;
												assign node2786 = (inp[13]) ? 14'b00000000011111 : 14'b00000000011111;
												assign node2789 = (inp[8]) ? 14'b00000000001111 : 14'b00000000001111;
									assign node2792 = (inp[4]) ? node2800 : node2793;
										assign node2793 = (inp[8]) ? 14'b00000000011111 : node2794;
											assign node2794 = (inp[3]) ? node2796 : 14'b00000001111111;
												assign node2796 = (inp[2]) ? 14'b00000000011111 : 14'b00000000111111;
										assign node2800 = (inp[8]) ? node2806 : node2801;
											assign node2801 = (inp[2]) ? node2803 : 14'b00000000011111;
												assign node2803 = (inp[3]) ? 14'b00000000001111 : 14'b00000000011111;
											assign node2806 = (inp[10]) ? node2810 : node2807;
												assign node2807 = (inp[2]) ? 14'b00000000001111 : 14'b00000000011111;
												assign node2810 = (inp[2]) ? 14'b00000000000011 : 14'b00000000000111;
					assign node2813 = (inp[4]) ? node2995 : node2814;
						assign node2814 = (inp[8]) ? node2906 : node2815;
							assign node2815 = (inp[9]) ? node2857 : node2816;
								assign node2816 = (inp[2]) ? node2840 : node2817;
									assign node2817 = (inp[11]) ? node2827 : node2818;
										assign node2818 = (inp[3]) ? 14'b00000011111111 : node2819;
											assign node2819 = (inp[12]) ? node2823 : node2820;
												assign node2820 = (inp[13]) ? 14'b00000111111111 : 14'b00001111111111;
												assign node2823 = (inp[13]) ? 14'b00000011111111 : 14'b00000111111111;
										assign node2827 = (inp[10]) ? node2835 : node2828;
											assign node2828 = (inp[6]) ? node2832 : node2829;
												assign node2829 = (inp[3]) ? 14'b00000011111111 : 14'b00000111111111;
												assign node2832 = (inp[13]) ? 14'b00000000111111 : 14'b00000011111111;
											assign node2835 = (inp[13]) ? 14'b00000001111111 : node2836;
												assign node2836 = (inp[3]) ? 14'b00000001111111 : 14'b00000011111111;
									assign node2840 = (inp[12]) ? node2850 : node2841;
										assign node2841 = (inp[3]) ? node2843 : 14'b00000011111111;
											assign node2843 = (inp[6]) ? node2847 : node2844;
												assign node2844 = (inp[10]) ? 14'b00000001111111 : 14'b00000011111111;
												assign node2847 = (inp[13]) ? 14'b00000001111111 : 14'b00000011111111;
										assign node2850 = (inp[13]) ? 14'b00000000111111 : node2851;
											assign node2851 = (inp[6]) ? node2853 : 14'b00000001111111;
												assign node2853 = (inp[11]) ? 14'b00000000111111 : 14'b00000001111111;
								assign node2857 = (inp[10]) ? node2883 : node2858;
									assign node2858 = (inp[3]) ? node2872 : node2859;
										assign node2859 = (inp[2]) ? node2865 : node2860;
											assign node2860 = (inp[12]) ? 14'b00000011111111 : node2861;
												assign node2861 = (inp[6]) ? 14'b00000011111111 : 14'b00000111111111;
											assign node2865 = (inp[13]) ? node2869 : node2866;
												assign node2866 = (inp[6]) ? 14'b00000001111111 : 14'b00000011111111;
												assign node2869 = (inp[11]) ? 14'b00000000111111 : 14'b00000001111111;
										assign node2872 = (inp[13]) ? node2880 : node2873;
											assign node2873 = (inp[2]) ? node2877 : node2874;
												assign node2874 = (inp[11]) ? 14'b00000001111111 : 14'b00000011111111;
												assign node2877 = (inp[11]) ? 14'b00000000111111 : 14'b00000001111111;
											assign node2880 = (inp[11]) ? 14'b00000000011111 : 14'b00000000111111;
									assign node2883 = (inp[3]) ? node2895 : node2884;
										assign node2884 = (inp[6]) ? node2890 : node2885;
											assign node2885 = (inp[13]) ? node2887 : 14'b00000001111111;
												assign node2887 = (inp[2]) ? 14'b00000000111111 : 14'b00000000111111;
											assign node2890 = (inp[11]) ? node2892 : 14'b00000000111111;
												assign node2892 = (inp[12]) ? 14'b00000000011111 : 14'b00000000111111;
										assign node2895 = (inp[11]) ? node2901 : node2896;
											assign node2896 = (inp[13]) ? 14'b00000000011111 : node2897;
												assign node2897 = (inp[6]) ? 14'b00000000111111 : 14'b00000001111111;
											assign node2901 = (inp[12]) ? 14'b00000000001111 : node2902;
												assign node2902 = (inp[13]) ? 14'b00000000011111 : 14'b00000000011111;
							assign node2906 = (inp[6]) ? node2958 : node2907;
								assign node2907 = (inp[3]) ? node2933 : node2908;
									assign node2908 = (inp[12]) ? node2920 : node2909;
										assign node2909 = (inp[2]) ? node2915 : node2910;
											assign node2910 = (inp[13]) ? 14'b00000011111111 : node2911;
												assign node2911 = (inp[9]) ? 14'b00000011111111 : 14'b00000111111111;
											assign node2915 = (inp[10]) ? node2917 : 14'b00000011111111;
												assign node2917 = (inp[9]) ? 14'b00000000111111 : 14'b00000001111111;
										assign node2920 = (inp[9]) ? node2928 : node2921;
											assign node2921 = (inp[10]) ? node2925 : node2922;
												assign node2922 = (inp[2]) ? 14'b00000001111111 : 14'b00000011111111;
												assign node2925 = (inp[13]) ? 14'b00000000111111 : 14'b00000001111111;
											assign node2928 = (inp[11]) ? 14'b00000000111111 : node2929;
												assign node2929 = (inp[10]) ? 14'b00000000111111 : 14'b00000000111111;
									assign node2933 = (inp[10]) ? node2947 : node2934;
										assign node2934 = (inp[9]) ? node2942 : node2935;
											assign node2935 = (inp[11]) ? node2939 : node2936;
												assign node2936 = (inp[12]) ? 14'b00000001111111 : 14'b00000011111111;
												assign node2939 = (inp[13]) ? 14'b00000000111111 : 14'b00000001111111;
											assign node2942 = (inp[13]) ? node2944 : 14'b00000000111111;
												assign node2944 = (inp[12]) ? 14'b00000000011111 : 14'b00000000111111;
										assign node2947 = (inp[13]) ? node2953 : node2948;
											assign node2948 = (inp[9]) ? 14'b00000000111111 : node2949;
												assign node2949 = (inp[11]) ? 14'b00000000111111 : 14'b00000000111111;
											assign node2953 = (inp[12]) ? node2955 : 14'b00000000011111;
												assign node2955 = (inp[11]) ? 14'b00000000000111 : 14'b00000000001111;
								assign node2958 = (inp[9]) ? node2982 : node2959;
									assign node2959 = (inp[13]) ? node2969 : node2960;
										assign node2960 = (inp[10]) ? node2966 : node2961;
											assign node2961 = (inp[11]) ? node2963 : 14'b00000001111111;
												assign node2963 = (inp[12]) ? 14'b00000000111111 : 14'b00000001111111;
											assign node2966 = (inp[12]) ? 14'b00000000011111 : 14'b00000001111111;
										assign node2969 = (inp[2]) ? node2977 : node2970;
											assign node2970 = (inp[12]) ? node2974 : node2971;
												assign node2971 = (inp[11]) ? 14'b00000000111111 : 14'b00000001111111;
												assign node2974 = (inp[11]) ? 14'b00000000001111 : 14'b00000000111111;
											assign node2977 = (inp[12]) ? 14'b00000000011111 : node2978;
												assign node2978 = (inp[10]) ? 14'b00000000001111 : 14'b00000000011111;
									assign node2982 = (inp[2]) ? node2990 : node2983;
										assign node2983 = (inp[11]) ? 14'b00000000011111 : node2984;
											assign node2984 = (inp[3]) ? node2986 : 14'b00000000111111;
												assign node2986 = (inp[12]) ? 14'b00000000011111 : 14'b00000000111111;
										assign node2990 = (inp[10]) ? 14'b00000000001111 : node2991;
											assign node2991 = (inp[3]) ? 14'b00000000001111 : 14'b00000000011111;
						assign node2995 = (inp[2]) ? node3093 : node2996;
							assign node2996 = (inp[6]) ? node3042 : node2997;
								assign node2997 = (inp[8]) ? node3015 : node2998;
									assign node2998 = (inp[9]) ? node3008 : node2999;
										assign node2999 = (inp[10]) ? node3003 : node3000;
											assign node3000 = (inp[13]) ? 14'b00000011111111 : 14'b00000111111111;
											assign node3003 = (inp[12]) ? 14'b00000001111111 : node3004;
												assign node3004 = (inp[3]) ? 14'b00000001111111 : 14'b00000011111111;
										assign node3008 = (inp[10]) ? node3010 : 14'b00000001111111;
											assign node3010 = (inp[11]) ? 14'b00000000111111 : node3011;
												assign node3011 = (inp[13]) ? 14'b00000000111111 : 14'b00000001111111;
									assign node3015 = (inp[11]) ? node3029 : node3016;
										assign node3016 = (inp[3]) ? node3022 : node3017;
											assign node3017 = (inp[9]) ? 14'b00000001111111 : node3018;
												assign node3018 = (inp[12]) ? 14'b00000011111111 : 14'b00000011111111;
											assign node3022 = (inp[13]) ? node3026 : node3023;
												assign node3023 = (inp[9]) ? 14'b00000000111111 : 14'b00000001111111;
												assign node3026 = (inp[12]) ? 14'b00000000011111 : 14'b00000000111111;
										assign node3029 = (inp[10]) ? node3037 : node3030;
											assign node3030 = (inp[9]) ? node3034 : node3031;
												assign node3031 = (inp[3]) ? 14'b00000001111111 : 14'b00000000111111;
												assign node3034 = (inp[13]) ? 14'b00000000011111 : 14'b00000000111111;
											assign node3037 = (inp[9]) ? 14'b00000000001111 : node3038;
												assign node3038 = (inp[13]) ? 14'b00000000011111 : 14'b00000000111111;
								assign node3042 = (inp[10]) ? node3066 : node3043;
									assign node3043 = (inp[3]) ? node3057 : node3044;
										assign node3044 = (inp[13]) ? node3052 : node3045;
											assign node3045 = (inp[9]) ? node3049 : node3046;
												assign node3046 = (inp[12]) ? 14'b00000001111111 : 14'b00000011111111;
												assign node3049 = (inp[12]) ? 14'b00000000111111 : 14'b00000001111111;
											assign node3052 = (inp[8]) ? node3054 : 14'b00000001111111;
												assign node3054 = (inp[9]) ? 14'b00000000011111 : 14'b00000000111111;
										assign node3057 = (inp[8]) ? node3061 : node3058;
											assign node3058 = (inp[12]) ? 14'b00000000111111 : 14'b00000001111111;
											assign node3061 = (inp[9]) ? 14'b00000000011111 : node3062;
												assign node3062 = (inp[11]) ? 14'b00000000011111 : 14'b00000000111111;
									assign node3066 = (inp[9]) ? node3078 : node3067;
										assign node3067 = (inp[11]) ? node3073 : node3068;
											assign node3068 = (inp[3]) ? 14'b00000001111111 : node3069;
												assign node3069 = (inp[12]) ? 14'b00000000011111 : 14'b00000000111111;
											assign node3073 = (inp[12]) ? 14'b00000000011111 : node3074;
												assign node3074 = (inp[8]) ? 14'b00000000011111 : 14'b00000000111111;
										assign node3078 = (inp[11]) ? node3086 : node3079;
											assign node3079 = (inp[8]) ? node3083 : node3080;
												assign node3080 = (inp[13]) ? 14'b00000000011111 : 14'b00000000111111;
												assign node3083 = (inp[13]) ? 14'b00000000001111 : 14'b00000000011111;
											assign node3086 = (inp[13]) ? node3090 : node3087;
												assign node3087 = (inp[3]) ? 14'b00000000001111 : 14'b00000000011111;
												assign node3090 = (inp[3]) ? 14'b00000000000111 : 14'b00000000000111;
							assign node3093 = (inp[8]) ? node3147 : node3094;
								assign node3094 = (inp[3]) ? node3118 : node3095;
									assign node3095 = (inp[9]) ? node3107 : node3096;
										assign node3096 = (inp[13]) ? node3102 : node3097;
											assign node3097 = (inp[10]) ? node3099 : 14'b00000001111111;
												assign node3099 = (inp[11]) ? 14'b00000000111111 : 14'b00000001111111;
											assign node3102 = (inp[10]) ? node3104 : 14'b00000000111111;
												assign node3104 = (inp[6]) ? 14'b00000000011111 : 14'b00000000011111;
										assign node3107 = (inp[12]) ? node3113 : node3108;
											assign node3108 = (inp[11]) ? node3110 : 14'b00000000111111;
												assign node3110 = (inp[13]) ? 14'b00000000011111 : 14'b00000000111111;
											assign node3113 = (inp[6]) ? 14'b00000000001111 : node3114;
												assign node3114 = (inp[10]) ? 14'b00000000111111 : 14'b00000000011111;
									assign node3118 = (inp[11]) ? node3134 : node3119;
										assign node3119 = (inp[12]) ? node3127 : node3120;
											assign node3120 = (inp[13]) ? node3124 : node3121;
												assign node3121 = (inp[6]) ? 14'b00000000111111 : 14'b00000001111111;
												assign node3124 = (inp[9]) ? 14'b00000000001111 : 14'b00000000111111;
											assign node3127 = (inp[9]) ? node3131 : node3128;
												assign node3128 = (inp[10]) ? 14'b00000000011111 : 14'b00000000111111;
												assign node3131 = (inp[13]) ? 14'b00000000001111 : 14'b00000000011111;
										assign node3134 = (inp[10]) ? node3140 : node3135;
											assign node3135 = (inp[12]) ? node3137 : 14'b00000000011111;
												assign node3137 = (inp[9]) ? 14'b00000000001111 : 14'b00000000011111;
											assign node3140 = (inp[6]) ? node3144 : node3141;
												assign node3141 = (inp[9]) ? 14'b00000000001111 : 14'b00000000001111;
												assign node3144 = (inp[12]) ? 14'b00000000000011 : 14'b00000000000111;
								assign node3147 = (inp[9]) ? node3173 : node3148;
									assign node3148 = (inp[3]) ? node3160 : node3149;
										assign node3149 = (inp[12]) ? node3155 : node3150;
											assign node3150 = (inp[11]) ? node3152 : 14'b00000000111111;
												assign node3152 = (inp[10]) ? 14'b00000000111111 : 14'b00000000011111;
											assign node3155 = (inp[10]) ? node3157 : 14'b00000000011111;
												assign node3157 = (inp[13]) ? 14'b00000000001111 : 14'b00000000011111;
										assign node3160 = (inp[11]) ? node3168 : node3161;
											assign node3161 = (inp[13]) ? node3165 : node3162;
												assign node3162 = (inp[12]) ? 14'b00000000011111 : 14'b00000000011111;
												assign node3165 = (inp[10]) ? 14'b00000000001111 : 14'b00000000011111;
											assign node3168 = (inp[6]) ? 14'b00000000001111 : node3169;
												assign node3169 = (inp[13]) ? 14'b00000000001111 : 14'b00000000011111;
									assign node3173 = (inp[12]) ? node3187 : node3174;
										assign node3174 = (inp[3]) ? node3180 : node3175;
											assign node3175 = (inp[11]) ? node3177 : 14'b00000000111111;
												assign node3177 = (inp[10]) ? 14'b00000000001111 : 14'b00000000011111;
											assign node3180 = (inp[6]) ? node3184 : node3181;
												assign node3181 = (inp[13]) ? 14'b00000000001111 : 14'b00000000011111;
												assign node3184 = (inp[10]) ? 14'b00000000000111 : 14'b00000000001111;
										assign node3187 = (inp[13]) ? node3195 : node3188;
											assign node3188 = (inp[6]) ? node3192 : node3189;
												assign node3189 = (inp[3]) ? 14'b00000000001111 : 14'b00000000011111;
												assign node3192 = (inp[11]) ? 14'b00000000000111 : 14'b00000000001111;
											assign node3195 = (inp[10]) ? node3199 : node3196;
												assign node3196 = (inp[3]) ? 14'b00000000000111 : 14'b00000000011111;
												assign node3199 = (inp[6]) ? 14'b00000000000011 : 14'b00000000000011;
		assign node3202 = (inp[4]) ? node4886 : node3203;
			assign node3203 = (inp[11]) ? node4029 : node3204;
				assign node3204 = (inp[10]) ? node3626 : node3205;
					assign node3205 = (inp[3]) ? node3429 : node3206;
						assign node3206 = (inp[6]) ? node3320 : node3207;
							assign node3207 = (inp[0]) ? node3265 : node3208;
								assign node3208 = (inp[8]) ? node3238 : node3209;
									assign node3209 = (inp[9]) ? node3223 : node3210;
										assign node3210 = (inp[7]) ? node3216 : node3211;
											assign node3211 = (inp[1]) ? 14'b00011111111111 : node3212;
												assign node3212 = (inp[12]) ? 14'b00011111111111 : 14'b00111111111111;
											assign node3216 = (inp[2]) ? node3220 : node3217;
												assign node3217 = (inp[13]) ? 14'b00001111111111 : 14'b00011111111111;
												assign node3220 = (inp[13]) ? 14'b00000111111111 : 14'b00001111111111;
										assign node3223 = (inp[13]) ? node3231 : node3224;
											assign node3224 = (inp[1]) ? node3228 : node3225;
												assign node3225 = (inp[12]) ? 14'b00001111111111 : 14'b00001111111111;
												assign node3228 = (inp[2]) ? 14'b00000011111111 : 14'b00001111111111;
											assign node3231 = (inp[12]) ? node3235 : node3232;
												assign node3232 = (inp[1]) ? 14'b00000111111111 : 14'b00011111111111;
												assign node3235 = (inp[1]) ? 14'b00000011111111 : 14'b00000111111111;
									assign node3238 = (inp[12]) ? node3254 : node3239;
										assign node3239 = (inp[7]) ? node3247 : node3240;
											assign node3240 = (inp[9]) ? node3244 : node3241;
												assign node3241 = (inp[13]) ? 14'b00001111111111 : 14'b00011111111111;
												assign node3244 = (inp[2]) ? 14'b00000111111111 : 14'b00001111111111;
											assign node3247 = (inp[9]) ? node3251 : node3248;
												assign node3248 = (inp[2]) ? 14'b00000111111111 : 14'b00001111111111;
												assign node3251 = (inp[2]) ? 14'b00000011111111 : 14'b00000111111111;
										assign node3254 = (inp[13]) ? node3260 : node3255;
											assign node3255 = (inp[9]) ? 14'b00000111111111 : node3256;
												assign node3256 = (inp[2]) ? 14'b00000111111111 : 14'b00000111111111;
											assign node3260 = (inp[7]) ? 14'b00000011111111 : node3261;
												assign node3261 = (inp[9]) ? 14'b00000011111111 : 14'b00000111111111;
								assign node3265 = (inp[12]) ? node3293 : node3266;
									assign node3266 = (inp[8]) ? node3280 : node3267;
										assign node3267 = (inp[1]) ? node3273 : node3268;
											assign node3268 = (inp[13]) ? node3270 : 14'b00011111111111;
												assign node3270 = (inp[2]) ? 14'b00000111111111 : 14'b00001111111111;
											assign node3273 = (inp[13]) ? node3277 : node3274;
												assign node3274 = (inp[7]) ? 14'b00000111111111 : 14'b00001111111111;
												assign node3277 = (inp[7]) ? 14'b00000011111111 : 14'b00000111111111;
										assign node3280 = (inp[13]) ? node3288 : node3281;
											assign node3281 = (inp[1]) ? node3285 : node3282;
												assign node3282 = (inp[9]) ? 14'b00000111111111 : 14'b00000111111111;
												assign node3285 = (inp[2]) ? 14'b00000011111111 : 14'b00000111111111;
											assign node3288 = (inp[7]) ? node3290 : 14'b00000111111111;
												assign node3290 = (inp[2]) ? 14'b00000001111111 : 14'b00000011111111;
									assign node3293 = (inp[8]) ? node3309 : node3294;
										assign node3294 = (inp[7]) ? node3302 : node3295;
											assign node3295 = (inp[1]) ? node3299 : node3296;
												assign node3296 = (inp[9]) ? 14'b00000111111111 : 14'b00001111111111;
												assign node3299 = (inp[2]) ? 14'b00000011111111 : 14'b00000111111111;
											assign node3302 = (inp[13]) ? node3306 : node3303;
												assign node3303 = (inp[9]) ? 14'b00000011111111 : 14'b00000111111111;
												assign node3306 = (inp[9]) ? 14'b00000001111111 : 14'b00000001111111;
										assign node3309 = (inp[2]) ? node3315 : node3310;
											assign node3310 = (inp[13]) ? node3312 : 14'b00000111111111;
												assign node3312 = (inp[9]) ? 14'b00000001111111 : 14'b00000001111111;
											assign node3315 = (inp[13]) ? 14'b00000001111111 : node3316;
												assign node3316 = (inp[7]) ? 14'b00000000111111 : 14'b00000001111111;
							assign node3320 = (inp[9]) ? node3376 : node3321;
								assign node3321 = (inp[12]) ? node3349 : node3322;
									assign node3322 = (inp[7]) ? node3334 : node3323;
										assign node3323 = (inp[8]) ? node3329 : node3324;
											assign node3324 = (inp[13]) ? 14'b00001111111111 : node3325;
												assign node3325 = (inp[0]) ? 14'b00001111111111 : 14'b00011111111111;
											assign node3329 = (inp[0]) ? 14'b00000111111111 : node3330;
												assign node3330 = (inp[13]) ? 14'b00000111111111 : 14'b00001111111111;
										assign node3334 = (inp[13]) ? node3342 : node3335;
											assign node3335 = (inp[0]) ? node3339 : node3336;
												assign node3336 = (inp[1]) ? 14'b00001111111111 : 14'b00001111111111;
												assign node3339 = (inp[1]) ? 14'b00000011111111 : 14'b00000011111111;
											assign node3342 = (inp[2]) ? node3346 : node3343;
												assign node3343 = (inp[1]) ? 14'b00000011111111 : 14'b00000111111111;
												assign node3346 = (inp[0]) ? 14'b00000001111111 : 14'b00000011111111;
									assign node3349 = (inp[8]) ? node3363 : node3350;
										assign node3350 = (inp[2]) ? node3356 : node3351;
											assign node3351 = (inp[0]) ? node3353 : 14'b00001111111111;
												assign node3353 = (inp[7]) ? 14'b00000011111111 : 14'b00000111111111;
											assign node3356 = (inp[7]) ? node3360 : node3357;
												assign node3357 = (inp[0]) ? 14'b00000011111111 : 14'b00000011111111;
												assign node3360 = (inp[13]) ? 14'b00000001111111 : 14'b00000011111111;
										assign node3363 = (inp[1]) ? node3369 : node3364;
											assign node3364 = (inp[7]) ? node3366 : 14'b00000011111111;
												assign node3366 = (inp[0]) ? 14'b00000001111111 : 14'b00000111111111;
											assign node3369 = (inp[0]) ? node3373 : node3370;
												assign node3370 = (inp[2]) ? 14'b00000001111111 : 14'b00000011111111;
												assign node3373 = (inp[13]) ? 14'b00000000011111 : 14'b00000000111111;
								assign node3376 = (inp[2]) ? node3406 : node3377;
									assign node3377 = (inp[13]) ? node3391 : node3378;
										assign node3378 = (inp[8]) ? node3386 : node3379;
											assign node3379 = (inp[0]) ? node3383 : node3380;
												assign node3380 = (inp[12]) ? 14'b00000111111111 : 14'b00001111111111;
												assign node3383 = (inp[1]) ? 14'b00000011111111 : 14'b00001111111111;
											assign node3386 = (inp[12]) ? 14'b00000001111111 : node3387;
												assign node3387 = (inp[7]) ? 14'b00000011111111 : 14'b00000011111111;
										assign node3391 = (inp[12]) ? node3399 : node3392;
											assign node3392 = (inp[0]) ? node3396 : node3393;
												assign node3393 = (inp[7]) ? 14'b00000011111111 : 14'b00000111111111;
												assign node3396 = (inp[7]) ? 14'b00000000111111 : 14'b00000011111111;
											assign node3399 = (inp[8]) ? node3403 : node3400;
												assign node3400 = (inp[7]) ? 14'b00000001111111 : 14'b00000011111111;
												assign node3403 = (inp[1]) ? 14'b00000000111111 : 14'b00000001111111;
									assign node3406 = (inp[1]) ? node3418 : node3407;
										assign node3407 = (inp[12]) ? node3415 : node3408;
											assign node3408 = (inp[8]) ? node3412 : node3409;
												assign node3409 = (inp[0]) ? 14'b00000001111111 : 14'b00000011111111;
												assign node3412 = (inp[13]) ? 14'b00000001111111 : 14'b00000001111111;
											assign node3415 = (inp[8]) ? 14'b00000000111111 : 14'b00000001111111;
										assign node3418 = (inp[0]) ? node3424 : node3419;
											assign node3419 = (inp[13]) ? node3421 : 14'b00000001111111;
												assign node3421 = (inp[12]) ? 14'b00000000111111 : 14'b00000001111111;
											assign node3424 = (inp[13]) ? 14'b00000000011111 : node3425;
												assign node3425 = (inp[7]) ? 14'b00000000111111 : 14'b00000001111111;
						assign node3429 = (inp[6]) ? node3539 : node3430;
							assign node3430 = (inp[9]) ? node3484 : node3431;
								assign node3431 = (inp[12]) ? node3463 : node3432;
									assign node3432 = (inp[7]) ? node3448 : node3433;
										assign node3433 = (inp[8]) ? node3441 : node3434;
											assign node3434 = (inp[2]) ? node3438 : node3435;
												assign node3435 = (inp[0]) ? 14'b00001111111111 : 14'b00011111111111;
												assign node3438 = (inp[0]) ? 14'b00000111111111 : 14'b00001111111111;
											assign node3441 = (inp[13]) ? node3445 : node3442;
												assign node3442 = (inp[1]) ? 14'b00000111111111 : 14'b00001111111111;
												assign node3445 = (inp[1]) ? 14'b00000011111111 : 14'b00000111111111;
										assign node3448 = (inp[8]) ? node3456 : node3449;
											assign node3449 = (inp[13]) ? node3453 : node3450;
												assign node3450 = (inp[2]) ? 14'b00000111111111 : 14'b00001111111111;
												assign node3453 = (inp[1]) ? 14'b00000011111111 : 14'b00000111111111;
											assign node3456 = (inp[1]) ? node3460 : node3457;
												assign node3457 = (inp[0]) ? 14'b00000011111111 : 14'b00000111111111;
												assign node3460 = (inp[13]) ? 14'b00000001111111 : 14'b00000011111111;
									assign node3463 = (inp[2]) ? node3473 : node3464;
										assign node3464 = (inp[0]) ? 14'b00000011111111 : node3465;
											assign node3465 = (inp[13]) ? node3469 : node3466;
												assign node3466 = (inp[1]) ? 14'b00000111111111 : 14'b00001111111111;
												assign node3469 = (inp[7]) ? 14'b00000011111111 : 14'b00000111111111;
										assign node3473 = (inp[13]) ? node3479 : node3474;
											assign node3474 = (inp[0]) ? 14'b00000001111111 : node3475;
												assign node3475 = (inp[7]) ? 14'b00000011111111 : 14'b00000111111111;
											assign node3479 = (inp[7]) ? 14'b00000000111111 : node3480;
												assign node3480 = (inp[8]) ? 14'b00000001111111 : 14'b00000011111111;
								assign node3484 = (inp[7]) ? node3512 : node3485;
									assign node3485 = (inp[12]) ? node3501 : node3486;
										assign node3486 = (inp[8]) ? node3494 : node3487;
											assign node3487 = (inp[1]) ? node3491 : node3488;
												assign node3488 = (inp[2]) ? 14'b00000011111111 : 14'b00000111111111;
												assign node3491 = (inp[13]) ? 14'b00000011111111 : 14'b00000011111111;
											assign node3494 = (inp[0]) ? node3498 : node3495;
												assign node3495 = (inp[1]) ? 14'b00000011111111 : 14'b00000011111111;
												assign node3498 = (inp[1]) ? 14'b00000001111111 : 14'b00000011111111;
										assign node3501 = (inp[13]) ? node3509 : node3502;
											assign node3502 = (inp[2]) ? node3506 : node3503;
												assign node3503 = (inp[1]) ? 14'b00000011111111 : 14'b00000111111111;
												assign node3506 = (inp[8]) ? 14'b00000001111111 : 14'b00000011111111;
											assign node3509 = (inp[0]) ? 14'b00000000011111 : 14'b00000001111111;
									assign node3512 = (inp[8]) ? node3526 : node3513;
										assign node3513 = (inp[13]) ? node3521 : node3514;
											assign node3514 = (inp[12]) ? node3518 : node3515;
												assign node3515 = (inp[2]) ? 14'b00000111111111 : 14'b00000111111111;
												assign node3518 = (inp[0]) ? 14'b00000001111111 : 14'b00000001111111;
											assign node3521 = (inp[1]) ? node3523 : 14'b00000001111111;
												assign node3523 = (inp[2]) ? 14'b00000000111111 : 14'b00000001111111;
										assign node3526 = (inp[2]) ? node3534 : node3527;
											assign node3527 = (inp[13]) ? node3531 : node3528;
												assign node3528 = (inp[0]) ? 14'b00000001111111 : 14'b00000011111111;
												assign node3531 = (inp[0]) ? 14'b00000000011111 : 14'b00000001111111;
											assign node3534 = (inp[12]) ? node3536 : 14'b00000000111111;
												assign node3536 = (inp[0]) ? 14'b00000000011111 : 14'b00000000111111;
							assign node3539 = (inp[0]) ? node3583 : node3540;
								assign node3540 = (inp[12]) ? node3566 : node3541;
									assign node3541 = (inp[13]) ? node3557 : node3542;
										assign node3542 = (inp[9]) ? node3550 : node3543;
											assign node3543 = (inp[7]) ? node3547 : node3544;
												assign node3544 = (inp[8]) ? 14'b00000111111111 : 14'b00001111111111;
												assign node3547 = (inp[1]) ? 14'b00000011111111 : 14'b00000111111111;
											assign node3550 = (inp[7]) ? node3554 : node3551;
												assign node3551 = (inp[2]) ? 14'b00000011111111 : 14'b00000111111111;
												assign node3554 = (inp[8]) ? 14'b00000001111111 : 14'b00000011111111;
										assign node3557 = (inp[8]) ? node3563 : node3558;
											assign node3558 = (inp[7]) ? node3560 : 14'b00000011111111;
												assign node3560 = (inp[2]) ? 14'b00000001111111 : 14'b00000011111111;
											assign node3563 = (inp[9]) ? 14'b00000000011111 : 14'b00000000111111;
									assign node3566 = (inp[7]) ? node3574 : node3567;
										assign node3567 = (inp[1]) ? node3571 : node3568;
											assign node3568 = (inp[9]) ? 14'b00000001111111 : 14'b00000111111111;
											assign node3571 = (inp[9]) ? 14'b00000011111111 : 14'b00000001111111;
										assign node3574 = (inp[1]) ? node3576 : 14'b00000001111111;
											assign node3576 = (inp[2]) ? node3580 : node3577;
												assign node3577 = (inp[9]) ? 14'b00000000111111 : 14'b00000001111111;
												assign node3580 = (inp[9]) ? 14'b00000000001111 : 14'b00000000011111;
								assign node3583 = (inp[2]) ? node3599 : node3584;
									assign node3584 = (inp[13]) ? node3590 : node3585;
										assign node3585 = (inp[12]) ? 14'b00000001111111 : node3586;
											assign node3586 = (inp[1]) ? 14'b00000001111111 : 14'b00000011111111;
										assign node3590 = (inp[12]) ? 14'b00000000111111 : node3591;
											assign node3591 = (inp[9]) ? node3595 : node3592;
												assign node3592 = (inp[1]) ? 14'b00000001111111 : 14'b00000001111111;
												assign node3595 = (inp[1]) ? 14'b00000000111111 : 14'b00000001111111;
									assign node3599 = (inp[7]) ? node3613 : node3600;
										assign node3600 = (inp[13]) ? node3608 : node3601;
											assign node3601 = (inp[12]) ? node3605 : node3602;
												assign node3602 = (inp[9]) ? 14'b00000001111111 : 14'b00000011111111;
												assign node3605 = (inp[9]) ? 14'b00000000111111 : 14'b00000001111111;
											assign node3608 = (inp[12]) ? node3610 : 14'b00000000111111;
												assign node3610 = (inp[8]) ? 14'b00000000011111 : 14'b00000000111111;
										assign node3613 = (inp[1]) ? node3619 : node3614;
											assign node3614 = (inp[8]) ? node3616 : 14'b00000001111111;
												assign node3616 = (inp[12]) ? 14'b00000000011111 : 14'b00000000111111;
											assign node3619 = (inp[12]) ? node3623 : node3620;
												assign node3620 = (inp[13]) ? 14'b00000000011111 : 14'b00000000111111;
												assign node3623 = (inp[13]) ? 14'b00000000001111 : 14'b00000000011111;
					assign node3626 = (inp[7]) ? node3822 : node3627;
						assign node3627 = (inp[9]) ? node3723 : node3628;
							assign node3628 = (inp[6]) ? node3678 : node3629;
								assign node3629 = (inp[12]) ? node3653 : node3630;
									assign node3630 = (inp[3]) ? node3644 : node3631;
										assign node3631 = (inp[1]) ? node3639 : node3632;
											assign node3632 = (inp[13]) ? node3636 : node3633;
												assign node3633 = (inp[2]) ? 14'b00001111111111 : 14'b00011111111111;
												assign node3636 = (inp[2]) ? 14'b00000111111111 : 14'b00001111111111;
											assign node3639 = (inp[0]) ? 14'b00000111111111 : node3640;
												assign node3640 = (inp[13]) ? 14'b00000111111111 : 14'b00001111111111;
										assign node3644 = (inp[8]) ? node3648 : node3645;
											assign node3645 = (inp[13]) ? 14'b00000111111111 : 14'b00001111111111;
											assign node3648 = (inp[2]) ? 14'b00000011111111 : node3649;
												assign node3649 = (inp[0]) ? 14'b00000011111111 : 14'b00000111111111;
									assign node3653 = (inp[13]) ? node3667 : node3654;
										assign node3654 = (inp[8]) ? node3662 : node3655;
											assign node3655 = (inp[3]) ? node3659 : node3656;
												assign node3656 = (inp[1]) ? 14'b00000111111111 : 14'b00001111111111;
												assign node3659 = (inp[1]) ? 14'b00000011111111 : 14'b00000111111111;
											assign node3662 = (inp[1]) ? 14'b00000011111111 : node3663;
												assign node3663 = (inp[3]) ? 14'b00000001111111 : 14'b00000111111111;
										assign node3667 = (inp[1]) ? node3675 : node3668;
											assign node3668 = (inp[2]) ? node3672 : node3669;
												assign node3669 = (inp[8]) ? 14'b00000011111111 : 14'b00000111111111;
												assign node3672 = (inp[3]) ? 14'b00000001111111 : 14'b00000011111111;
											assign node3675 = (inp[2]) ? 14'b00000000111111 : 14'b00000001111111;
								assign node3678 = (inp[13]) ? node3700 : node3679;
									assign node3679 = (inp[0]) ? node3693 : node3680;
										assign node3680 = (inp[2]) ? node3688 : node3681;
											assign node3681 = (inp[3]) ? node3685 : node3682;
												assign node3682 = (inp[1]) ? 14'b00000111111111 : 14'b00001111111111;
												assign node3685 = (inp[12]) ? 14'b00000011111111 : 14'b00000111111111;
											assign node3688 = (inp[3]) ? 14'b00000001111111 : node3689;
												assign node3689 = (inp[12]) ? 14'b00000011111111 : 14'b00000111111111;
										assign node3693 = (inp[1]) ? node3697 : node3694;
											assign node3694 = (inp[3]) ? 14'b00000001111111 : 14'b00000011111111;
											assign node3697 = (inp[2]) ? 14'b00000000011111 : 14'b00000001111111;
									assign node3700 = (inp[1]) ? node3716 : node3701;
										assign node3701 = (inp[12]) ? node3709 : node3702;
											assign node3702 = (inp[2]) ? node3706 : node3703;
												assign node3703 = (inp[0]) ? 14'b00000011111111 : 14'b00000011111111;
												assign node3706 = (inp[0]) ? 14'b00000001111111 : 14'b00000011111111;
											assign node3709 = (inp[0]) ? node3713 : node3710;
												assign node3710 = (inp[3]) ? 14'b00000001111111 : 14'b00000011111111;
												assign node3713 = (inp[3]) ? 14'b00000000111111 : 14'b00000001111111;
										assign node3716 = (inp[12]) ? 14'b00000001111111 : node3717;
											assign node3717 = (inp[0]) ? 14'b00000000111111 : node3718;
												assign node3718 = (inp[3]) ? 14'b00000000111111 : 14'b00000001111111;
							assign node3723 = (inp[12]) ? node3777 : node3724;
								assign node3724 = (inp[1]) ? node3750 : node3725;
									assign node3725 = (inp[6]) ? node3739 : node3726;
										assign node3726 = (inp[0]) ? node3734 : node3727;
											assign node3727 = (inp[13]) ? node3731 : node3728;
												assign node3728 = (inp[2]) ? 14'b00000111111111 : 14'b00001111111111;
												assign node3731 = (inp[3]) ? 14'b00000011111111 : 14'b00000111111111;
											assign node3734 = (inp[3]) ? 14'b00000001111111 : node3735;
												assign node3735 = (inp[13]) ? 14'b00000011111111 : 14'b00000011111111;
										assign node3739 = (inp[0]) ? node3747 : node3740;
											assign node3740 = (inp[3]) ? node3744 : node3741;
												assign node3741 = (inp[13]) ? 14'b00000011111111 : 14'b00000011111111;
												assign node3744 = (inp[13]) ? 14'b00000001111111 : 14'b00000011111111;
											assign node3747 = (inp[8]) ? 14'b00000001111111 : 14'b00000111111111;
									assign node3750 = (inp[0]) ? node3762 : node3751;
										assign node3751 = (inp[2]) ? node3757 : node3752;
											assign node3752 = (inp[6]) ? 14'b00000011111111 : node3753;
												assign node3753 = (inp[8]) ? 14'b00000011111111 : 14'b00000111111111;
											assign node3757 = (inp[8]) ? 14'b00000000111111 : node3758;
												assign node3758 = (inp[6]) ? 14'b00000001111111 : 14'b00000011111111;
										assign node3762 = (inp[6]) ? node3770 : node3763;
											assign node3763 = (inp[13]) ? node3767 : node3764;
												assign node3764 = (inp[2]) ? 14'b00000001111111 : 14'b00000111111111;
												assign node3767 = (inp[2]) ? 14'b00000000111111 : 14'b00000001111111;
											assign node3770 = (inp[13]) ? node3774 : node3771;
												assign node3771 = (inp[8]) ? 14'b00000000111111 : 14'b00000001111111;
												assign node3774 = (inp[2]) ? 14'b00000000011111 : 14'b00000000111111;
								assign node3777 = (inp[2]) ? node3799 : node3778;
									assign node3778 = (inp[6]) ? node3792 : node3779;
										assign node3779 = (inp[3]) ? node3785 : node3780;
											assign node3780 = (inp[8]) ? 14'b00000011111111 : node3781;
												assign node3781 = (inp[13]) ? 14'b00000011111111 : 14'b00000111111111;
											assign node3785 = (inp[8]) ? node3789 : node3786;
												assign node3786 = (inp[13]) ? 14'b00000001111111 : 14'b00000011111111;
												assign node3789 = (inp[0]) ? 14'b00000000111111 : 14'b00000001111111;
										assign node3792 = (inp[13]) ? node3794 : 14'b00000001111111;
											assign node3794 = (inp[3]) ? node3796 : 14'b00000001111111;
												assign node3796 = (inp[8]) ? 14'b00000000011111 : 14'b00000000111111;
									assign node3799 = (inp[0]) ? node3813 : node3800;
										assign node3800 = (inp[13]) ? node3808 : node3801;
											assign node3801 = (inp[1]) ? node3805 : node3802;
												assign node3802 = (inp[6]) ? 14'b00000001111111 : 14'b00000011111111;
												assign node3805 = (inp[3]) ? 14'b00000000111111 : 14'b00000001111111;
											assign node3808 = (inp[1]) ? node3810 : 14'b00000000111111;
												assign node3810 = (inp[8]) ? 14'b00000000011111 : 14'b00000000111111;
										assign node3813 = (inp[3]) ? node3815 : 14'b00000001111111;
											assign node3815 = (inp[1]) ? node3819 : node3816;
												assign node3816 = (inp[6]) ? 14'b00000000011111 : 14'b00000000111111;
												assign node3819 = (inp[8]) ? 14'b00000000001111 : 14'b00000000011111;
						assign node3822 = (inp[13]) ? node3924 : node3823;
							assign node3823 = (inp[12]) ? node3873 : node3824;
								assign node3824 = (inp[0]) ? node3852 : node3825;
									assign node3825 = (inp[1]) ? node3839 : node3826;
										assign node3826 = (inp[8]) ? node3832 : node3827;
											assign node3827 = (inp[6]) ? 14'b00000111111111 : node3828;
												assign node3828 = (inp[3]) ? 14'b00000111111111 : 14'b00001111111111;
											assign node3832 = (inp[9]) ? node3836 : node3833;
												assign node3833 = (inp[3]) ? 14'b00000011111111 : 14'b00000111111111;
												assign node3836 = (inp[3]) ? 14'b00000001111111 : 14'b00000011111111;
										assign node3839 = (inp[6]) ? node3845 : node3840;
											assign node3840 = (inp[8]) ? node3842 : 14'b00000011111111;
												assign node3842 = (inp[9]) ? 14'b00000001111111 : 14'b00000011111111;
											assign node3845 = (inp[9]) ? node3849 : node3846;
												assign node3846 = (inp[3]) ? 14'b00000001111111 : 14'b00000001111111;
												assign node3849 = (inp[8]) ? 14'b00000000011111 : 14'b00000001111111;
									assign node3852 = (inp[9]) ? node3864 : node3853;
										assign node3853 = (inp[6]) ? node3859 : node3854;
											assign node3854 = (inp[2]) ? 14'b00000011111111 : node3855;
												assign node3855 = (inp[1]) ? 14'b00000001111111 : 14'b00000011111111;
											assign node3859 = (inp[2]) ? 14'b00000001111111 : node3860;
												assign node3860 = (inp[1]) ? 14'b00000001111111 : 14'b00000011111111;
										assign node3864 = (inp[2]) ? node3866 : 14'b00000001111111;
											assign node3866 = (inp[1]) ? node3870 : node3867;
												assign node3867 = (inp[6]) ? 14'b00000000111111 : 14'b00000001111111;
												assign node3870 = (inp[3]) ? 14'b00000000011111 : 14'b00000000011111;
								assign node3873 = (inp[6]) ? node3899 : node3874;
									assign node3874 = (inp[3]) ? node3886 : node3875;
										assign node3875 = (inp[8]) ? node3881 : node3876;
											assign node3876 = (inp[0]) ? node3878 : 14'b00000011111111;
												assign node3878 = (inp[2]) ? 14'b00000001111111 : 14'b00000001111111;
											assign node3881 = (inp[1]) ? node3883 : 14'b00000001111111;
												assign node3883 = (inp[2]) ? 14'b00000000111111 : 14'b00000001111111;
										assign node3886 = (inp[2]) ? node3892 : node3887;
											assign node3887 = (inp[0]) ? node3889 : 14'b00000011111111;
												assign node3889 = (inp[1]) ? 14'b00000000111111 : 14'b00000001111111;
											assign node3892 = (inp[9]) ? node3896 : node3893;
												assign node3893 = (inp[1]) ? 14'b00000000011111 : 14'b00000000111111;
												assign node3896 = (inp[8]) ? 14'b00000000111111 : 14'b00000000111111;
									assign node3899 = (inp[9]) ? node3911 : node3900;
										assign node3900 = (inp[1]) ? node3906 : node3901;
											assign node3901 = (inp[8]) ? 14'b00000000111111 : node3902;
												assign node3902 = (inp[3]) ? 14'b00000000111111 : 14'b00000001111111;
											assign node3906 = (inp[3]) ? 14'b00000001111111 : node3907;
												assign node3907 = (inp[8]) ? 14'b00000001111111 : 14'b00000011111111;
										assign node3911 = (inp[1]) ? node3917 : node3912;
											assign node3912 = (inp[0]) ? 14'b00000000111111 : node3913;
												assign node3913 = (inp[2]) ? 14'b00000000111111 : 14'b00000001111111;
											assign node3917 = (inp[2]) ? node3921 : node3918;
												assign node3918 = (inp[8]) ? 14'b00000000011111 : 14'b00000000111111;
												assign node3921 = (inp[0]) ? 14'b00000000001111 : 14'b00000000011111;
							assign node3924 = (inp[3]) ? node3978 : node3925;
								assign node3925 = (inp[0]) ? node3949 : node3926;
									assign node3926 = (inp[2]) ? node3938 : node3927;
										assign node3927 = (inp[8]) ? node3933 : node3928;
											assign node3928 = (inp[1]) ? node3930 : 14'b00000011111111;
												assign node3930 = (inp[12]) ? 14'b00000000111111 : 14'b00000001111111;
											assign node3933 = (inp[6]) ? node3935 : 14'b00000001111111;
												assign node3935 = (inp[12]) ? 14'b00000001111111 : 14'b00000001111111;
										assign node3938 = (inp[8]) ? node3944 : node3939;
											assign node3939 = (inp[6]) ? node3941 : 14'b00000011111111;
												assign node3941 = (inp[1]) ? 14'b00000000111111 : 14'b00000001111111;
											assign node3944 = (inp[6]) ? 14'b00000000011111 : node3945;
												assign node3945 = (inp[12]) ? 14'b00000000111111 : 14'b00000001111111;
									assign node3949 = (inp[8]) ? node3963 : node3950;
										assign node3950 = (inp[9]) ? node3958 : node3951;
											assign node3951 = (inp[2]) ? node3955 : node3952;
												assign node3952 = (inp[6]) ? 14'b00000001111111 : 14'b00000011111111;
												assign node3955 = (inp[1]) ? 14'b00000000111111 : 14'b00000001111111;
											assign node3958 = (inp[1]) ? 14'b00000000011111 : node3959;
												assign node3959 = (inp[12]) ? 14'b00000000111111 : 14'b00000001111111;
										assign node3963 = (inp[2]) ? node3971 : node3964;
											assign node3964 = (inp[6]) ? node3968 : node3965;
												assign node3965 = (inp[12]) ? 14'b00000000111111 : 14'b00000001111111;
												assign node3968 = (inp[1]) ? 14'b00000000001111 : 14'b00000000111111;
											assign node3971 = (inp[12]) ? node3975 : node3972;
												assign node3972 = (inp[9]) ? 14'b00000000011111 : 14'b00000000111111;
												assign node3975 = (inp[6]) ? 14'b00000000001111 : 14'b00000000011111;
								assign node3978 = (inp[8]) ? node4002 : node3979;
									assign node3979 = (inp[6]) ? node3993 : node3980;
										assign node3980 = (inp[12]) ? node3986 : node3981;
											assign node3981 = (inp[1]) ? node3983 : 14'b00000001111111;
												assign node3983 = (inp[9]) ? 14'b00000000111111 : 14'b00000001111111;
											assign node3986 = (inp[2]) ? node3990 : node3987;
												assign node3987 = (inp[9]) ? 14'b00000000111111 : 14'b00000000111111;
												assign node3990 = (inp[1]) ? 14'b00000000011111 : 14'b00000000111111;
										assign node3993 = (inp[0]) ? node3999 : node3994;
											assign node3994 = (inp[1]) ? 14'b00000000011111 : node3995;
												assign node3995 = (inp[9]) ? 14'b00000000111111 : 14'b00000001111111;
											assign node3999 = (inp[9]) ? 14'b00000000001111 : 14'b00000000011111;
									assign node4002 = (inp[1]) ? node4016 : node4003;
										assign node4003 = (inp[0]) ? node4009 : node4004;
											assign node4004 = (inp[6]) ? node4006 : 14'b00000001111111;
												assign node4006 = (inp[9]) ? 14'b00000000011111 : 14'b00000000111111;
											assign node4009 = (inp[2]) ? node4013 : node4010;
												assign node4010 = (inp[9]) ? 14'b00000000011111 : 14'b00000000111111;
												assign node4013 = (inp[6]) ? 14'b00000000001111 : 14'b00000000011111;
										assign node4016 = (inp[2]) ? node4022 : node4017;
											assign node4017 = (inp[6]) ? 14'b00000000001111 : node4018;
												assign node4018 = (inp[9]) ? 14'b00000000001111 : 14'b00000000011111;
											assign node4022 = (inp[12]) ? node4026 : node4023;
												assign node4023 = (inp[6]) ? 14'b00000000001111 : 14'b00000000011111;
												assign node4026 = (inp[0]) ? 14'b00000000000111 : 14'b00000000000111;
				assign node4029 = (inp[6]) ? node4455 : node4030;
					assign node4030 = (inp[0]) ? node4252 : node4031;
						assign node4031 = (inp[12]) ? node4137 : node4032;
							assign node4032 = (inp[3]) ? node4086 : node4033;
								assign node4033 = (inp[10]) ? node4061 : node4034;
									assign node4034 = (inp[1]) ? node4046 : node4035;
										assign node4035 = (inp[7]) ? node4043 : node4036;
											assign node4036 = (inp[13]) ? node4040 : node4037;
												assign node4037 = (inp[9]) ? 14'b00011111111111 : 14'b00111111111111;
												assign node4040 = (inp[2]) ? 14'b00001111111111 : 14'b00001111111111;
											assign node4043 = (inp[13]) ? 14'b00000111111111 : 14'b00001111111111;
										assign node4046 = (inp[8]) ? node4054 : node4047;
											assign node4047 = (inp[9]) ? node4051 : node4048;
												assign node4048 = (inp[7]) ? 14'b00001111111111 : 14'b00001111111111;
												assign node4051 = (inp[13]) ? 14'b00000001111111 : 14'b00000111111111;
											assign node4054 = (inp[13]) ? node4058 : node4055;
												assign node4055 = (inp[9]) ? 14'b00000011111111 : 14'b00000111111111;
												assign node4058 = (inp[9]) ? 14'b00000001111111 : 14'b00000011111111;
									assign node4061 = (inp[13]) ? node4075 : node4062;
										assign node4062 = (inp[7]) ? node4068 : node4063;
											assign node4063 = (inp[2]) ? 14'b00000111111111 : node4064;
												assign node4064 = (inp[9]) ? 14'b00000111111111 : 14'b00001111111111;
											assign node4068 = (inp[1]) ? node4072 : node4069;
												assign node4069 = (inp[9]) ? 14'b00000011111111 : 14'b00001111111111;
												assign node4072 = (inp[2]) ? 14'b00000011111111 : 14'b00000011111111;
										assign node4075 = (inp[2]) ? node4079 : node4076;
											assign node4076 = (inp[1]) ? 14'b00000111111111 : 14'b00000011111111;
											assign node4079 = (inp[7]) ? node4083 : node4080;
												assign node4080 = (inp[9]) ? 14'b00000001111111 : 14'b00000011111111;
												assign node4083 = (inp[8]) ? 14'b00000000111111 : 14'b00000001111111;
								assign node4086 = (inp[1]) ? node4114 : node4087;
									assign node4087 = (inp[13]) ? node4103 : node4088;
										assign node4088 = (inp[7]) ? node4096 : node4089;
											assign node4089 = (inp[9]) ? node4093 : node4090;
												assign node4090 = (inp[2]) ? 14'b00000111111111 : 14'b00001111111111;
												assign node4093 = (inp[8]) ? 14'b00000011111111 : 14'b00000011111111;
											assign node4096 = (inp[10]) ? node4100 : node4097;
												assign node4097 = (inp[8]) ? 14'b00000011111111 : 14'b00000111111111;
												assign node4100 = (inp[9]) ? 14'b00000001111111 : 14'b00000011111111;
										assign node4103 = (inp[7]) ? node4109 : node4104;
											assign node4104 = (inp[8]) ? node4106 : 14'b00000011111111;
												assign node4106 = (inp[10]) ? 14'b00000011111111 : 14'b00000011111111;
											assign node4109 = (inp[9]) ? 14'b00000001111111 : node4110;
												assign node4110 = (inp[8]) ? 14'b00000001111111 : 14'b00000011111111;
									assign node4114 = (inp[9]) ? node4124 : node4115;
										assign node4115 = (inp[13]) ? node4121 : node4116;
											assign node4116 = (inp[10]) ? 14'b00000011111111 : node4117;
												assign node4117 = (inp[2]) ? 14'b00000011111111 : 14'b00000111111111;
											assign node4121 = (inp[7]) ? 14'b00000011111111 : 14'b00000001111111;
										assign node4124 = (inp[7]) ? node4132 : node4125;
											assign node4125 = (inp[8]) ? node4129 : node4126;
												assign node4126 = (inp[10]) ? 14'b00000001111111 : 14'b00000011111111;
												assign node4129 = (inp[13]) ? 14'b00000000111111 : 14'b00000001111111;
											assign node4132 = (inp[13]) ? node4134 : 14'b00000000011111;
												assign node4134 = (inp[2]) ? 14'b00000000001111 : 14'b00000000011111;
							assign node4137 = (inp[7]) ? node4199 : node4138;
								assign node4138 = (inp[3]) ? node4168 : node4139;
									assign node4139 = (inp[1]) ? node4153 : node4140;
										assign node4140 = (inp[8]) ? node4146 : node4141;
											assign node4141 = (inp[13]) ? 14'b00000111111111 : node4142;
												assign node4142 = (inp[10]) ? 14'b00000011111111 : 14'b00001111111111;
											assign node4146 = (inp[13]) ? node4150 : node4147;
												assign node4147 = (inp[9]) ? 14'b00000011111111 : 14'b00000111111111;
												assign node4150 = (inp[9]) ? 14'b00000001111111 : 14'b00000011111111;
										assign node4153 = (inp[8]) ? node4161 : node4154;
											assign node4154 = (inp[2]) ? node4158 : node4155;
												assign node4155 = (inp[13]) ? 14'b00000011111111 : 14'b00000111111111;
												assign node4158 = (inp[10]) ? 14'b00000001111111 : 14'b00000011111111;
											assign node4161 = (inp[13]) ? node4165 : node4162;
												assign node4162 = (inp[2]) ? 14'b00000001111111 : 14'b00000011111111;
												assign node4165 = (inp[9]) ? 14'b00000000111111 : 14'b00000001111111;
									assign node4168 = (inp[1]) ? node4184 : node4169;
										assign node4169 = (inp[13]) ? node4177 : node4170;
											assign node4170 = (inp[2]) ? node4174 : node4171;
												assign node4171 = (inp[10]) ? 14'b00000011111111 : 14'b00000111111111;
												assign node4174 = (inp[10]) ? 14'b00000001111111 : 14'b00000011111111;
											assign node4177 = (inp[8]) ? node4181 : node4178;
												assign node4178 = (inp[10]) ? 14'b00000001111111 : 14'b00000001111111;
												assign node4181 = (inp[10]) ? 14'b00000000111111 : 14'b00000001111111;
										assign node4184 = (inp[13]) ? node4192 : node4185;
											assign node4185 = (inp[9]) ? node4189 : node4186;
												assign node4186 = (inp[2]) ? 14'b00000000111111 : 14'b00000011111111;
												assign node4189 = (inp[10]) ? 14'b00000000111111 : 14'b00000001111111;
											assign node4192 = (inp[10]) ? node4196 : node4193;
												assign node4193 = (inp[8]) ? 14'b00000000111111 : 14'b00000000111111;
												assign node4196 = (inp[9]) ? 14'b00000000011111 : 14'b00000000111111;
								assign node4199 = (inp[13]) ? node4231 : node4200;
									assign node4200 = (inp[8]) ? node4216 : node4201;
										assign node4201 = (inp[10]) ? node4209 : node4202;
											assign node4202 = (inp[9]) ? node4206 : node4203;
												assign node4203 = (inp[3]) ? 14'b00000001111111 : 14'b00000011111111;
												assign node4206 = (inp[3]) ? 14'b00000011111111 : 14'b00000111111111;
											assign node4209 = (inp[2]) ? node4213 : node4210;
												assign node4210 = (inp[1]) ? 14'b00000011111111 : 14'b00000001111111;
												assign node4213 = (inp[3]) ? 14'b00000000111111 : 14'b00000001111111;
										assign node4216 = (inp[10]) ? node4224 : node4217;
											assign node4217 = (inp[3]) ? node4221 : node4218;
												assign node4218 = (inp[2]) ? 14'b00000001111111 : 14'b00000011111111;
												assign node4221 = (inp[1]) ? 14'b00000000111111 : 14'b00000001111111;
											assign node4224 = (inp[3]) ? node4228 : node4225;
												assign node4225 = (inp[2]) ? 14'b00000000111111 : 14'b00000001111111;
												assign node4228 = (inp[1]) ? 14'b00000000001111 : 14'b00000000111111;
									assign node4231 = (inp[8]) ? node4241 : node4232;
										assign node4232 = (inp[3]) ? node4236 : node4233;
											assign node4233 = (inp[9]) ? 14'b00000000111111 : 14'b00000001111111;
											assign node4236 = (inp[9]) ? node4238 : 14'b00000000111111;
												assign node4238 = (inp[2]) ? 14'b00000000011111 : 14'b00000000111111;
										assign node4241 = (inp[1]) ? node4245 : node4242;
											assign node4242 = (inp[9]) ? 14'b00000000011111 : 14'b00000001111111;
											assign node4245 = (inp[10]) ? node4249 : node4246;
												assign node4246 = (inp[3]) ? 14'b00000000001111 : 14'b00000000011111;
												assign node4249 = (inp[9]) ? 14'b00000000001111 : 14'b00000000011111;
						assign node4252 = (inp[13]) ? node4354 : node4253;
							assign node4253 = (inp[9]) ? node4305 : node4254;
								assign node4254 = (inp[1]) ? node4278 : node4255;
									assign node4255 = (inp[12]) ? node4269 : node4256;
										assign node4256 = (inp[2]) ? node4262 : node4257;
											assign node4257 = (inp[10]) ? 14'b00000111111111 : node4258;
												assign node4258 = (inp[8]) ? 14'b00001111111111 : 14'b00001111111111;
											assign node4262 = (inp[3]) ? node4266 : node4263;
												assign node4263 = (inp[8]) ? 14'b00000011111111 : 14'b00000111111111;
												assign node4266 = (inp[8]) ? 14'b00000001111111 : 14'b00000011111111;
										assign node4269 = (inp[8]) ? node4275 : node4270;
											assign node4270 = (inp[3]) ? node4272 : 14'b00000111111111;
												assign node4272 = (inp[10]) ? 14'b00000001111111 : 14'b00000011111111;
											assign node4275 = (inp[3]) ? 14'b00000001111111 : 14'b00000000111111;
									assign node4278 = (inp[7]) ? node4294 : node4279;
										assign node4279 = (inp[3]) ? node4287 : node4280;
											assign node4280 = (inp[12]) ? node4284 : node4281;
												assign node4281 = (inp[8]) ? 14'b00000011111111 : 14'b00000111111111;
												assign node4284 = (inp[2]) ? 14'b00000001111111 : 14'b00000011111111;
											assign node4287 = (inp[8]) ? node4291 : node4288;
												assign node4288 = (inp[2]) ? 14'b00000001111111 : 14'b00000011111111;
												assign node4291 = (inp[12]) ? 14'b00000000111111 : 14'b00000001111111;
										assign node4294 = (inp[12]) ? node4300 : node4295;
											assign node4295 = (inp[3]) ? node4297 : 14'b00000001111111;
												assign node4297 = (inp[2]) ? 14'b00000000111111 : 14'b00000001111111;
											assign node4300 = (inp[10]) ? node4302 : 14'b00000000111111;
												assign node4302 = (inp[8]) ? 14'b00000000001111 : 14'b00000000011111;
								assign node4305 = (inp[3]) ? node4325 : node4306;
									assign node4306 = (inp[1]) ? node4314 : node4307;
										assign node4307 = (inp[12]) ? node4309 : 14'b00000011111111;
											assign node4309 = (inp[2]) ? 14'b00000001111111 : node4310;
												assign node4310 = (inp[8]) ? 14'b00000001111111 : 14'b00000011111111;
										assign node4314 = (inp[8]) ? node4318 : node4315;
											assign node4315 = (inp[12]) ? 14'b00000001111111 : 14'b00000011111111;
											assign node4318 = (inp[7]) ? node4322 : node4319;
												assign node4319 = (inp[2]) ? 14'b00000000111111 : 14'b00000001111111;
												assign node4322 = (inp[10]) ? 14'b00000000011111 : 14'b00000000111111;
									assign node4325 = (inp[8]) ? node4339 : node4326;
										assign node4326 = (inp[10]) ? node4334 : node4327;
											assign node4327 = (inp[7]) ? node4331 : node4328;
												assign node4328 = (inp[12]) ? 14'b00000001111111 : 14'b00000011111111;
												assign node4331 = (inp[12]) ? 14'b00000000111111 : 14'b00000000111111;
											assign node4334 = (inp[1]) ? node4336 : 14'b00000000111111;
												assign node4336 = (inp[7]) ? 14'b00000000011111 : 14'b00000000111111;
										assign node4339 = (inp[12]) ? node4347 : node4340;
											assign node4340 = (inp[10]) ? node4344 : node4341;
												assign node4341 = (inp[2]) ? 14'b00000000111111 : 14'b00000001111111;
												assign node4344 = (inp[1]) ? 14'b00000000011111 : 14'b00000000111111;
											assign node4347 = (inp[1]) ? node4351 : node4348;
												assign node4348 = (inp[10]) ? 14'b00000000011111 : 14'b00000000111111;
												assign node4351 = (inp[7]) ? 14'b00000000001111 : 14'b00000000011111;
							assign node4354 = (inp[1]) ? node4408 : node4355;
								assign node4355 = (inp[7]) ? node4379 : node4356;
									assign node4356 = (inp[12]) ? node4366 : node4357;
										assign node4357 = (inp[8]) ? node4361 : node4358;
											assign node4358 = (inp[2]) ? 14'b00000011111111 : 14'b00000111111111;
											assign node4361 = (inp[9]) ? node4363 : 14'b00000011111111;
												assign node4363 = (inp[10]) ? 14'b00000000111111 : 14'b00000001111111;
										assign node4366 = (inp[10]) ? node4372 : node4367;
											assign node4367 = (inp[8]) ? node4369 : 14'b00000001111111;
												assign node4369 = (inp[9]) ? 14'b00000000111111 : 14'b00000001111111;
											assign node4372 = (inp[9]) ? node4376 : node4373;
												assign node4373 = (inp[8]) ? 14'b00000000111111 : 14'b00000000111111;
												assign node4376 = (inp[2]) ? 14'b00000000011111 : 14'b00000000111111;
									assign node4379 = (inp[3]) ? node4395 : node4380;
										assign node4380 = (inp[12]) ? node4388 : node4381;
											assign node4381 = (inp[10]) ? node4385 : node4382;
												assign node4382 = (inp[9]) ? 14'b00000001111111 : 14'b00000011111111;
												assign node4385 = (inp[9]) ? 14'b00000000111111 : 14'b00000001111111;
											assign node4388 = (inp[2]) ? node4392 : node4389;
												assign node4389 = (inp[9]) ? 14'b00000000011111 : 14'b00000001111111;
												assign node4392 = (inp[8]) ? 14'b00000000011111 : 14'b00000000111111;
										assign node4395 = (inp[9]) ? node4403 : node4396;
											assign node4396 = (inp[2]) ? node4400 : node4397;
												assign node4397 = (inp[8]) ? 14'b00000000111111 : 14'b00000001111111;
												assign node4400 = (inp[8]) ? 14'b00000000011111 : 14'b00000000111111;
											assign node4403 = (inp[8]) ? node4405 : 14'b00000000011111;
												assign node4405 = (inp[12]) ? 14'b00000000001111 : 14'b00000000001111;
								assign node4408 = (inp[8]) ? node4432 : node4409;
									assign node4409 = (inp[7]) ? node4423 : node4410;
										assign node4410 = (inp[2]) ? node4416 : node4411;
											assign node4411 = (inp[10]) ? node4413 : 14'b00000011111111;
												assign node4413 = (inp[3]) ? 14'b00000000111111 : 14'b00000001111111;
											assign node4416 = (inp[10]) ? node4420 : node4417;
												assign node4417 = (inp[9]) ? 14'b00000000111111 : 14'b00000001111111;
												assign node4420 = (inp[9]) ? 14'b00000000011111 : 14'b00000000111111;
										assign node4423 = (inp[12]) ? node4429 : node4424;
											assign node4424 = (inp[2]) ? node4426 : 14'b00000000111111;
												assign node4426 = (inp[3]) ? 14'b00000000011111 : 14'b00000000111111;
											assign node4429 = (inp[9]) ? 14'b00000000000111 : 14'b00000000011111;
									assign node4432 = (inp[2]) ? node4440 : node4433;
										assign node4433 = (inp[3]) ? 14'b00000000011111 : node4434;
											assign node4434 = (inp[7]) ? 14'b00000000011111 : node4435;
												assign node4435 = (inp[9]) ? 14'b00000000111111 : 14'b00000001111111;
										assign node4440 = (inp[10]) ? node4448 : node4441;
											assign node4441 = (inp[3]) ? node4445 : node4442;
												assign node4442 = (inp[9]) ? 14'b00000000011111 : 14'b00000000111111;
												assign node4445 = (inp[9]) ? 14'b00000000001111 : 14'b00000000011111;
											assign node4448 = (inp[9]) ? node4452 : node4449;
												assign node4449 = (inp[12]) ? 14'b00000000001111 : 14'b00000000011111;
												assign node4452 = (inp[3]) ? 14'b00000000000111 : 14'b00000000001111;
					assign node4455 = (inp[1]) ? node4673 : node4456;
						assign node4456 = (inp[12]) ? node4566 : node4457;
							assign node4457 = (inp[8]) ? node4511 : node4458;
								assign node4458 = (inp[2]) ? node4482 : node4459;
									assign node4459 = (inp[0]) ? node4473 : node4460;
										assign node4460 = (inp[13]) ? node4468 : node4461;
											assign node4461 = (inp[3]) ? node4465 : node4462;
												assign node4462 = (inp[10]) ? 14'b00000111111111 : 14'b00001111111111;
												assign node4465 = (inp[10]) ? 14'b00000011111111 : 14'b00000111111111;
											assign node4468 = (inp[3]) ? 14'b00000011111111 : node4469;
												assign node4469 = (inp[7]) ? 14'b00000011111111 : 14'b00000111111111;
										assign node4473 = (inp[7]) ? 14'b00000001111111 : node4474;
											assign node4474 = (inp[13]) ? node4478 : node4475;
												assign node4475 = (inp[3]) ? 14'b00000011111111 : 14'b00000011111111;
												assign node4478 = (inp[10]) ? 14'b00000001111111 : 14'b00000001111111;
									assign node4482 = (inp[3]) ? node4498 : node4483;
										assign node4483 = (inp[10]) ? node4491 : node4484;
											assign node4484 = (inp[13]) ? node4488 : node4485;
												assign node4485 = (inp[9]) ? 14'b00000011111111 : 14'b00000111111111;
												assign node4488 = (inp[7]) ? 14'b00000001111111 : 14'b00000011111111;
											assign node4491 = (inp[7]) ? node4495 : node4492;
												assign node4492 = (inp[9]) ? 14'b00000001111111 : 14'b00000011111111;
												assign node4495 = (inp[13]) ? 14'b00000000111111 : 14'b00000001111111;
										assign node4498 = (inp[13]) ? node4504 : node4499;
											assign node4499 = (inp[7]) ? node4501 : 14'b00000011111111;
												assign node4501 = (inp[10]) ? 14'b00000000111111 : 14'b00000001111111;
											assign node4504 = (inp[10]) ? node4508 : node4505;
												assign node4505 = (inp[9]) ? 14'b00000000111111 : 14'b00000000111111;
												assign node4508 = (inp[7]) ? 14'b00000000011111 : 14'b00000000111111;
								assign node4511 = (inp[3]) ? node4537 : node4512;
									assign node4512 = (inp[13]) ? node4522 : node4513;
										assign node4513 = (inp[10]) ? 14'b00000001111111 : node4514;
											assign node4514 = (inp[0]) ? node4518 : node4515;
												assign node4515 = (inp[2]) ? 14'b00000011111111 : 14'b00000111111111;
												assign node4518 = (inp[7]) ? 14'b00000001111111 : 14'b00000011111111;
										assign node4522 = (inp[9]) ? node4530 : node4523;
											assign node4523 = (inp[7]) ? node4527 : node4524;
												assign node4524 = (inp[0]) ? 14'b00000001111111 : 14'b00000001111111;
												assign node4527 = (inp[10]) ? 14'b00000000111111 : 14'b00000001111111;
											assign node4530 = (inp[10]) ? node4534 : node4531;
												assign node4531 = (inp[7]) ? 14'b00000000111111 : 14'b00000001111111;
												assign node4534 = (inp[0]) ? 14'b00000000011111 : 14'b00000000111111;
									assign node4537 = (inp[7]) ? node4553 : node4538;
										assign node4538 = (inp[13]) ? node4546 : node4539;
											assign node4539 = (inp[0]) ? node4543 : node4540;
												assign node4540 = (inp[9]) ? 14'b00000001111111 : 14'b00000011111111;
												assign node4543 = (inp[9]) ? 14'b00000000111111 : 14'b00000001111111;
											assign node4546 = (inp[10]) ? node4550 : node4547;
												assign node4547 = (inp[9]) ? 14'b00000000111111 : 14'b00000011111111;
												assign node4550 = (inp[0]) ? 14'b00000000011111 : 14'b00000000111111;
										assign node4553 = (inp[13]) ? node4561 : node4554;
											assign node4554 = (inp[2]) ? node4558 : node4555;
												assign node4555 = (inp[0]) ? 14'b00000000111111 : 14'b00000000111111;
												assign node4558 = (inp[9]) ? 14'b00000000001111 : 14'b00000000111111;
											assign node4561 = (inp[0]) ? node4563 : 14'b00000000111111;
												assign node4563 = (inp[9]) ? 14'b00000000001111 : 14'b00000000001111;
							assign node4566 = (inp[10]) ? node4612 : node4567;
								assign node4567 = (inp[9]) ? node4591 : node4568;
									assign node4568 = (inp[3]) ? node4582 : node4569;
										assign node4569 = (inp[0]) ? node4575 : node4570;
											assign node4570 = (inp[2]) ? node4572 : 14'b00000111111111;
												assign node4572 = (inp[8]) ? 14'b00000000111111 : 14'b00000011111111;
											assign node4575 = (inp[13]) ? node4579 : node4576;
												assign node4576 = (inp[7]) ? 14'b00000001111111 : 14'b00000011111111;
												assign node4579 = (inp[8]) ? 14'b00000000111111 : 14'b00000001111111;
										assign node4582 = (inp[13]) ? node4586 : node4583;
											assign node4583 = (inp[8]) ? 14'b00000001111111 : 14'b00000000111111;
											assign node4586 = (inp[8]) ? 14'b00000000111111 : node4587;
												assign node4587 = (inp[7]) ? 14'b00000000111111 : 14'b00000001111111;
									assign node4591 = (inp[13]) ? node4601 : node4592;
										assign node4592 = (inp[2]) ? node4596 : node4593;
											assign node4593 = (inp[3]) ? 14'b00000001111111 : 14'b00000011111111;
											assign node4596 = (inp[7]) ? 14'b00000000011111 : node4597;
												assign node4597 = (inp[0]) ? 14'b00000000111111 : 14'b00000001111111;
										assign node4601 = (inp[2]) ? node4607 : node4602;
											assign node4602 = (inp[7]) ? node4604 : 14'b00000000111111;
												assign node4604 = (inp[0]) ? 14'b00000000011111 : 14'b00000000111111;
											assign node4607 = (inp[3]) ? node4609 : 14'b00000000111111;
												assign node4609 = (inp[0]) ? 14'b00000000001111 : 14'b00000000001111;
								assign node4612 = (inp[0]) ? node4644 : node4613;
									assign node4613 = (inp[8]) ? node4629 : node4614;
										assign node4614 = (inp[7]) ? node4622 : node4615;
											assign node4615 = (inp[2]) ? node4619 : node4616;
												assign node4616 = (inp[13]) ? 14'b00000001111111 : 14'b00000011111111;
												assign node4619 = (inp[9]) ? 14'b00000000111111 : 14'b00000001111111;
											assign node4622 = (inp[3]) ? node4626 : node4623;
												assign node4623 = (inp[13]) ? 14'b00000000111111 : 14'b00000001111111;
												assign node4626 = (inp[2]) ? 14'b00000000011111 : 14'b00000000111111;
										assign node4629 = (inp[7]) ? node4637 : node4630;
											assign node4630 = (inp[13]) ? node4634 : node4631;
												assign node4631 = (inp[2]) ? 14'b00000000111111 : 14'b00000001111111;
												assign node4634 = (inp[3]) ? 14'b00000000011111 : 14'b00000000111111;
											assign node4637 = (inp[9]) ? node4641 : node4638;
												assign node4638 = (inp[3]) ? 14'b00000000001111 : 14'b00000000011111;
												assign node4641 = (inp[3]) ? 14'b00000000001111 : 14'b00000000001111;
									assign node4644 = (inp[2]) ? node4660 : node4645;
										assign node4645 = (inp[7]) ? node4653 : node4646;
											assign node4646 = (inp[8]) ? node4650 : node4647;
												assign node4647 = (inp[13]) ? 14'b00000000111111 : 14'b00000001111111;
												assign node4650 = (inp[13]) ? 14'b00000000011111 : 14'b00000000111111;
											assign node4653 = (inp[3]) ? node4657 : node4654;
												assign node4654 = (inp[13]) ? 14'b00000000011111 : 14'b00000000011111;
												assign node4657 = (inp[13]) ? 14'b00000000001111 : 14'b00000000011111;
										assign node4660 = (inp[8]) ? node4666 : node4661;
											assign node4661 = (inp[7]) ? node4663 : 14'b00000000011111;
												assign node4663 = (inp[9]) ? 14'b00000000001111 : 14'b00000000011111;
											assign node4666 = (inp[3]) ? node4670 : node4667;
												assign node4667 = (inp[7]) ? 14'b00000000001111 : 14'b00000000011111;
												assign node4670 = (inp[7]) ? 14'b00000000000111 : 14'b00000000001111;
						assign node4673 = (inp[2]) ? node4781 : node4674;
							assign node4674 = (inp[13]) ? node4726 : node4675;
								assign node4675 = (inp[8]) ? node4701 : node4676;
									assign node4676 = (inp[10]) ? node4688 : node4677;
										assign node4677 = (inp[7]) ? node4681 : node4678;
											assign node4678 = (inp[12]) ? 14'b00000011111111 : 14'b00000111111111;
											assign node4681 = (inp[0]) ? node4685 : node4682;
												assign node4682 = (inp[12]) ? 14'b00000001111111 : 14'b00000011111111;
												assign node4685 = (inp[12]) ? 14'b00000000111111 : 14'b00000001111111;
										assign node4688 = (inp[9]) ? node4696 : node4689;
											assign node4689 = (inp[12]) ? node4693 : node4690;
												assign node4690 = (inp[7]) ? 14'b00000001111111 : 14'b00000011111111;
												assign node4693 = (inp[7]) ? 14'b00000000111111 : 14'b00000001111111;
											assign node4696 = (inp[3]) ? 14'b00000000011111 : node4697;
												assign node4697 = (inp[7]) ? 14'b00000000111111 : 14'b00000000111111;
									assign node4701 = (inp[3]) ? node4717 : node4702;
										assign node4702 = (inp[0]) ? node4710 : node4703;
											assign node4703 = (inp[9]) ? node4707 : node4704;
												assign node4704 = (inp[12]) ? 14'b00000001111111 : 14'b00000011111111;
												assign node4707 = (inp[10]) ? 14'b00000000111111 : 14'b00000000111111;
											assign node4710 = (inp[9]) ? node4714 : node4711;
												assign node4711 = (inp[7]) ? 14'b00000000111111 : 14'b00000000111111;
												assign node4714 = (inp[10]) ? 14'b00000000011111 : 14'b00000000111111;
										assign node4717 = (inp[10]) ? node4719 : 14'b00000000111111;
											assign node4719 = (inp[0]) ? node4723 : node4720;
												assign node4720 = (inp[9]) ? 14'b00000000011111 : 14'b00000000111111;
												assign node4723 = (inp[9]) ? 14'b00000000001111 : 14'b00000000011111;
								assign node4726 = (inp[12]) ? node4754 : node4727;
									assign node4727 = (inp[8]) ? node4739 : node4728;
										assign node4728 = (inp[9]) ? node4734 : node4729;
											assign node4729 = (inp[7]) ? 14'b00000001111111 : node4730;
												assign node4730 = (inp[3]) ? 14'b00000001111111 : 14'b00000011111111;
											assign node4734 = (inp[0]) ? node4736 : 14'b00000001111111;
												assign node4736 = (inp[10]) ? 14'b00000000011111 : 14'b00000000111111;
										assign node4739 = (inp[0]) ? node4747 : node4740;
											assign node4740 = (inp[10]) ? node4744 : node4741;
												assign node4741 = (inp[3]) ? 14'b00000000111111 : 14'b00000000111111;
												assign node4744 = (inp[7]) ? 14'b00000000011111 : 14'b00000000111111;
											assign node4747 = (inp[9]) ? node4751 : node4748;
												assign node4748 = (inp[10]) ? 14'b00000000111111 : 14'b00000000011111;
												assign node4751 = (inp[7]) ? 14'b00000000000111 : 14'b00000000001111;
									assign node4754 = (inp[0]) ? node4770 : node4755;
										assign node4755 = (inp[10]) ? node4763 : node4756;
											assign node4756 = (inp[9]) ? node4760 : node4757;
												assign node4757 = (inp[8]) ? 14'b00000000111111 : 14'b00000001111111;
												assign node4760 = (inp[3]) ? 14'b00000000011111 : 14'b00000000111111;
											assign node4763 = (inp[3]) ? node4767 : node4764;
												assign node4764 = (inp[9]) ? 14'b00000000011111 : 14'b00000000111111;
												assign node4767 = (inp[8]) ? 14'b00000000001111 : 14'b00000000011111;
										assign node4770 = (inp[9]) ? node4778 : node4771;
											assign node4771 = (inp[3]) ? node4775 : node4772;
												assign node4772 = (inp[8]) ? 14'b00000000011111 : 14'b00000000111111;
												assign node4775 = (inp[7]) ? 14'b00000000001111 : 14'b00000000011111;
											assign node4778 = (inp[10]) ? 14'b00000000000111 : 14'b00000000001111;
							assign node4781 = (inp[7]) ? node4829 : node4782;
								assign node4782 = (inp[3]) ? node4806 : node4783;
									assign node4783 = (inp[8]) ? node4793 : node4784;
										assign node4784 = (inp[13]) ? node4788 : node4785;
											assign node4785 = (inp[10]) ? 14'b00000000111111 : 14'b00000001111111;
											assign node4788 = (inp[10]) ? node4790 : 14'b00000000111111;
												assign node4790 = (inp[0]) ? 14'b00000000011111 : 14'b00000000111111;
										assign node4793 = (inp[9]) ? node4801 : node4794;
											assign node4794 = (inp[12]) ? node4798 : node4795;
												assign node4795 = (inp[0]) ? 14'b00000000111111 : 14'b00000001111111;
												assign node4798 = (inp[10]) ? 14'b00000000011111 : 14'b00000000111111;
											assign node4801 = (inp[13]) ? node4803 : 14'b00000000011111;
												assign node4803 = (inp[10]) ? 14'b00000000001111 : 14'b00000000011111;
									assign node4806 = (inp[8]) ? node4816 : node4807;
										assign node4807 = (inp[10]) ? node4813 : node4808;
											assign node4808 = (inp[13]) ? node4810 : 14'b00000001111111;
												assign node4810 = (inp[12]) ? 14'b00000000011111 : 14'b00000000011111;
											assign node4813 = (inp[13]) ? 14'b00000000001111 : 14'b00000000011111;
										assign node4816 = (inp[0]) ? node4822 : node4817;
											assign node4817 = (inp[13]) ? node4819 : 14'b00000000011111;
												assign node4819 = (inp[12]) ? 14'b00000000001111 : 14'b00000000011111;
											assign node4822 = (inp[9]) ? node4826 : node4823;
												assign node4823 = (inp[10]) ? 14'b00000000001111 : 14'b00000000111111;
												assign node4826 = (inp[10]) ? 14'b00000000000011 : 14'b00000000001111;
								assign node4829 = (inp[0]) ? node4859 : node4830;
									assign node4830 = (inp[3]) ? node4846 : node4831;
										assign node4831 = (inp[10]) ? node4839 : node4832;
											assign node4832 = (inp[9]) ? node4836 : node4833;
												assign node4833 = (inp[13]) ? 14'b00000000111111 : 14'b00000011111111;
												assign node4836 = (inp[8]) ? 14'b00000000011111 : 14'b00000000111111;
											assign node4839 = (inp[12]) ? node4843 : node4840;
												assign node4840 = (inp[13]) ? 14'b00000000011111 : 14'b00000000111111;
												assign node4843 = (inp[8]) ? 14'b00000000001111 : 14'b00000000011111;
										assign node4846 = (inp[12]) ? node4852 : node4847;
											assign node4847 = (inp[10]) ? 14'b00000000001111 : node4848;
												assign node4848 = (inp[8]) ? 14'b00000000011111 : 14'b00000000011111;
											assign node4852 = (inp[13]) ? node4856 : node4853;
												assign node4853 = (inp[8]) ? 14'b00000000001111 : 14'b00000000011111;
												assign node4856 = (inp[10]) ? 14'b00000000000011 : 14'b00000000001111;
									assign node4859 = (inp[12]) ? node4873 : node4860;
										assign node4860 = (inp[9]) ? node4866 : node4861;
											assign node4861 = (inp[10]) ? node4863 : 14'b00000000011111;
												assign node4863 = (inp[8]) ? 14'b00000000001111 : 14'b00000000011111;
											assign node4866 = (inp[8]) ? node4870 : node4867;
												assign node4867 = (inp[13]) ? 14'b00000000001111 : 14'b00000000111111;
												assign node4870 = (inp[10]) ? 14'b00000000000111 : 14'b00000000001111;
										assign node4873 = (inp[13]) ? node4879 : node4874;
											assign node4874 = (inp[10]) ? node4876 : 14'b00000000001111;
												assign node4876 = (inp[3]) ? 14'b00000000000111 : 14'b00000000001111;
											assign node4879 = (inp[10]) ? node4883 : node4880;
												assign node4880 = (inp[3]) ? 14'b00000000000111 : 14'b00000000000111;
												assign node4883 = (inp[3]) ? 14'b00000000000001 : 14'b00000000000011;
			assign node4886 = (inp[1]) ? node5690 : node4887;
				assign node4887 = (inp[13]) ? node5281 : node4888;
					assign node4888 = (inp[10]) ? node5104 : node4889;
						assign node4889 = (inp[2]) ? node4995 : node4890;
							assign node4890 = (inp[9]) ? node4940 : node4891;
								assign node4891 = (inp[8]) ? node4915 : node4892;
									assign node4892 = (inp[6]) ? node4906 : node4893;
										assign node4893 = (inp[11]) ? node4899 : node4894;
											assign node4894 = (inp[7]) ? 14'b00000111111111 : node4895;
												assign node4895 = (inp[12]) ? 14'b00001111111111 : 14'b00011111111111;
											assign node4899 = (inp[0]) ? node4903 : node4900;
												assign node4900 = (inp[3]) ? 14'b00000111111111 : 14'b00001111111111;
												assign node4903 = (inp[3]) ? 14'b00000011111111 : 14'b00000111111111;
										assign node4906 = (inp[7]) ? 14'b00000011111111 : node4907;
											assign node4907 = (inp[0]) ? node4911 : node4908;
												assign node4908 = (inp[3]) ? 14'b00000111111111 : 14'b00000111111111;
												assign node4911 = (inp[12]) ? 14'b00000011111111 : 14'b00000111111111;
									assign node4915 = (inp[0]) ? node4929 : node4916;
										assign node4916 = (inp[11]) ? node4922 : node4917;
											assign node4917 = (inp[7]) ? 14'b00000111111111 : node4918;
												assign node4918 = (inp[3]) ? 14'b00000011111111 : 14'b00000111111111;
											assign node4922 = (inp[7]) ? node4926 : node4923;
												assign node4923 = (inp[3]) ? 14'b00000011111111 : 14'b00000111111111;
												assign node4926 = (inp[6]) ? 14'b00000001111111 : 14'b00000011111111;
										assign node4929 = (inp[11]) ? node4933 : node4930;
											assign node4930 = (inp[6]) ? 14'b00000001111111 : 14'b00000011111111;
											assign node4933 = (inp[12]) ? node4937 : node4934;
												assign node4934 = (inp[6]) ? 14'b00000001111111 : 14'b00000111111111;
												assign node4937 = (inp[3]) ? 14'b00000000111111 : 14'b00000001111111;
								assign node4940 = (inp[6]) ? node4966 : node4941;
									assign node4941 = (inp[0]) ? node4953 : node4942;
										assign node4942 = (inp[3]) ? node4948 : node4943;
											assign node4943 = (inp[8]) ? 14'b00000111111111 : node4944;
												assign node4944 = (inp[7]) ? 14'b00000111111111 : 14'b00001111111111;
											assign node4948 = (inp[12]) ? 14'b00000001111111 : node4949;
												assign node4949 = (inp[8]) ? 14'b00000011111111 : 14'b00000111111111;
										assign node4953 = (inp[3]) ? node4959 : node4954;
											assign node4954 = (inp[12]) ? node4956 : 14'b00000111111111;
												assign node4956 = (inp[11]) ? 14'b00000001111111 : 14'b00000011111111;
											assign node4959 = (inp[7]) ? node4963 : node4960;
												assign node4960 = (inp[8]) ? 14'b00000001111111 : 14'b00000011111111;
												assign node4963 = (inp[12]) ? 14'b00000000111111 : 14'b00000001111111;
									assign node4966 = (inp[8]) ? node4980 : node4967;
										assign node4967 = (inp[3]) ? node4973 : node4968;
											assign node4968 = (inp[0]) ? node4970 : 14'b00000111111111;
												assign node4970 = (inp[7]) ? 14'b00000001111111 : 14'b00000011111111;
											assign node4973 = (inp[12]) ? node4977 : node4974;
												assign node4974 = (inp[0]) ? 14'b00000001111111 : 14'b00000011111111;
												assign node4977 = (inp[7]) ? 14'b00000000111111 : 14'b00000001111111;
										assign node4980 = (inp[3]) ? node4988 : node4981;
											assign node4981 = (inp[11]) ? node4985 : node4982;
												assign node4982 = (inp[0]) ? 14'b00000001111111 : 14'b00000011111111;
												assign node4985 = (inp[7]) ? 14'b00000000111111 : 14'b00000001111111;
											assign node4988 = (inp[11]) ? node4992 : node4989;
												assign node4989 = (inp[0]) ? 14'b00000000011111 : 14'b00000000111111;
												assign node4992 = (inp[0]) ? 14'b00000000111111 : 14'b00000001111111;
							assign node4995 = (inp[3]) ? node5051 : node4996;
								assign node4996 = (inp[9]) ? node5022 : node4997;
									assign node4997 = (inp[12]) ? node5011 : node4998;
										assign node4998 = (inp[11]) ? node5006 : node4999;
											assign node4999 = (inp[8]) ? node5003 : node5000;
												assign node5000 = (inp[7]) ? 14'b00000111111111 : 14'b00001111111111;
												assign node5003 = (inp[6]) ? 14'b00000011111111 : 14'b00000111111111;
											assign node5006 = (inp[0]) ? 14'b00000011111111 : node5007;
												assign node5007 = (inp[7]) ? 14'b00000011111111 : 14'b00000111111111;
										assign node5011 = (inp[0]) ? node5017 : node5012;
											assign node5012 = (inp[8]) ? node5014 : 14'b00000111111111;
												assign node5014 = (inp[11]) ? 14'b00000001111111 : 14'b00000001111111;
											assign node5017 = (inp[7]) ? node5019 : 14'b00000011111111;
												assign node5019 = (inp[6]) ? 14'b00000000111111 : 14'b00000001111111;
									assign node5022 = (inp[8]) ? node5038 : node5023;
										assign node5023 = (inp[0]) ? node5031 : node5024;
											assign node5024 = (inp[12]) ? node5028 : node5025;
												assign node5025 = (inp[6]) ? 14'b00000011111111 : 14'b00000111111111;
												assign node5028 = (inp[6]) ? 14'b00000001111111 : 14'b00000011111111;
											assign node5031 = (inp[7]) ? node5035 : node5032;
												assign node5032 = (inp[12]) ? 14'b00000001111111 : 14'b00000011111111;
												assign node5035 = (inp[11]) ? 14'b00000000111111 : 14'b00000001111111;
										assign node5038 = (inp[6]) ? node5046 : node5039;
											assign node5039 = (inp[0]) ? node5043 : node5040;
												assign node5040 = (inp[7]) ? 14'b00000001111111 : 14'b00000011111111;
												assign node5043 = (inp[11]) ? 14'b00000000111111 : 14'b00000000111111;
											assign node5046 = (inp[7]) ? 14'b00000000111111 : node5047;
												assign node5047 = (inp[0]) ? 14'b00000000011111 : 14'b00000000111111;
								assign node5051 = (inp[6]) ? node5077 : node5052;
									assign node5052 = (inp[9]) ? node5066 : node5053;
										assign node5053 = (inp[7]) ? node5061 : node5054;
											assign node5054 = (inp[8]) ? node5058 : node5055;
												assign node5055 = (inp[11]) ? 14'b00000011111111 : 14'b00000111111111;
												assign node5058 = (inp[12]) ? 14'b00000001111111 : 14'b00000011111111;
											assign node5061 = (inp[12]) ? 14'b00000000111111 : node5062;
												assign node5062 = (inp[11]) ? 14'b00000001111111 : 14'b00000001111111;
										assign node5066 = (inp[0]) ? node5072 : node5067;
											assign node5067 = (inp[12]) ? node5069 : 14'b00000001111111;
												assign node5069 = (inp[7]) ? 14'b00000000111111 : 14'b00000001111111;
											assign node5072 = (inp[8]) ? node5074 : 14'b00000001111111;
												assign node5074 = (inp[11]) ? 14'b00000000011111 : 14'b00000000111111;
									assign node5077 = (inp[8]) ? node5091 : node5078;
										assign node5078 = (inp[11]) ? node5084 : node5079;
											assign node5079 = (inp[9]) ? node5081 : 14'b00000001111111;
												assign node5081 = (inp[12]) ? 14'b00000000111111 : 14'b00000001111111;
											assign node5084 = (inp[7]) ? node5088 : node5085;
												assign node5085 = (inp[0]) ? 14'b00000000111111 : 14'b00000001111111;
												assign node5088 = (inp[12]) ? 14'b00000000011111 : 14'b00000000111111;
										assign node5091 = (inp[12]) ? node5097 : node5092;
											assign node5092 = (inp[0]) ? 14'b00000000011111 : node5093;
												assign node5093 = (inp[7]) ? 14'b00000000111111 : 14'b00000001111111;
											assign node5097 = (inp[7]) ? node5101 : node5098;
												assign node5098 = (inp[11]) ? 14'b00000000011111 : 14'b00000000111111;
												assign node5101 = (inp[0]) ? 14'b00000000001111 : 14'b00000000011111;
						assign node5104 = (inp[7]) ? node5198 : node5105;
							assign node5105 = (inp[2]) ? node5155 : node5106;
								assign node5106 = (inp[8]) ? node5128 : node5107;
									assign node5107 = (inp[9]) ? node5119 : node5108;
										assign node5108 = (inp[6]) ? node5112 : node5109;
											assign node5109 = (inp[11]) ? 14'b00001111111111 : 14'b00000111111111;
											assign node5112 = (inp[12]) ? node5116 : node5113;
												assign node5113 = (inp[0]) ? 14'b00000011111111 : 14'b00000111111111;
												assign node5116 = (inp[3]) ? 14'b00000001111111 : 14'b00000011111111;
										assign node5119 = (inp[0]) ? node5125 : node5120;
											assign node5120 = (inp[12]) ? node5122 : 14'b00000011111111;
												assign node5122 = (inp[6]) ? 14'b00000001111111 : 14'b00000011111111;
											assign node5125 = (inp[6]) ? 14'b00000001111111 : 14'b00000000111111;
									assign node5128 = (inp[9]) ? node5142 : node5129;
										assign node5129 = (inp[0]) ? node5135 : node5130;
											assign node5130 = (inp[6]) ? node5132 : 14'b00001111111111;
												assign node5132 = (inp[11]) ? 14'b00000001111111 : 14'b00000011111111;
											assign node5135 = (inp[6]) ? node5139 : node5136;
												assign node5136 = (inp[3]) ? 14'b00000001111111 : 14'b00000011111111;
												assign node5139 = (inp[11]) ? 14'b00000000111111 : 14'b00000000111111;
										assign node5142 = (inp[0]) ? node5148 : node5143;
											assign node5143 = (inp[12]) ? node5145 : 14'b00000001111111;
												assign node5145 = (inp[3]) ? 14'b00000000111111 : 14'b00000001111111;
											assign node5148 = (inp[11]) ? node5152 : node5149;
												assign node5149 = (inp[3]) ? 14'b00000000111111 : 14'b00000001111111;
												assign node5152 = (inp[12]) ? 14'b00000000011111 : 14'b00000000111111;
								assign node5155 = (inp[3]) ? node5181 : node5156;
									assign node5156 = (inp[8]) ? node5168 : node5157;
										assign node5157 = (inp[6]) ? node5163 : node5158;
											assign node5158 = (inp[0]) ? 14'b00000011111111 : node5159;
												assign node5159 = (inp[9]) ? 14'b00000011111111 : 14'b00000111111111;
											assign node5163 = (inp[11]) ? node5165 : 14'b00000011111111;
												assign node5165 = (inp[9]) ? 14'b00000000111111 : 14'b00000001111111;
										assign node5168 = (inp[11]) ? node5174 : node5169;
											assign node5169 = (inp[6]) ? 14'b00000011111111 : node5170;
												assign node5170 = (inp[12]) ? 14'b00000001111111 : 14'b00000001111111;
											assign node5174 = (inp[9]) ? node5178 : node5175;
												assign node5175 = (inp[6]) ? 14'b00000000111111 : 14'b00000001111111;
												assign node5178 = (inp[12]) ? 14'b00000000001111 : 14'b00000000011111;
									assign node5181 = (inp[11]) ? node5189 : node5182;
										assign node5182 = (inp[6]) ? 14'b00000000111111 : node5183;
											assign node5183 = (inp[8]) ? 14'b00000000111111 : node5184;
												assign node5184 = (inp[9]) ? 14'b00000000111111 : 14'b00000001111111;
										assign node5189 = (inp[12]) ? 14'b00000000011111 : node5190;
											assign node5190 = (inp[9]) ? node5194 : node5191;
												assign node5191 = (inp[8]) ? 14'b00000000111111 : 14'b00000001111111;
												assign node5194 = (inp[6]) ? 14'b00000000001111 : 14'b00000000111111;
							assign node5198 = (inp[0]) ? node5238 : node5199;
								assign node5199 = (inp[6]) ? node5215 : node5200;
									assign node5200 = (inp[12]) ? node5212 : node5201;
										assign node5201 = (inp[8]) ? node5209 : node5202;
											assign node5202 = (inp[9]) ? node5206 : node5203;
												assign node5203 = (inp[3]) ? 14'b00000011111111 : 14'b00000111111111;
												assign node5206 = (inp[3]) ? 14'b00000001111111 : 14'b00000011111111;
											assign node5209 = (inp[2]) ? 14'b00000000111111 : 14'b00000001111111;
										assign node5212 = (inp[9]) ? 14'b00000000111111 : 14'b00000001111111;
									assign node5215 = (inp[9]) ? node5225 : node5216;
										assign node5216 = (inp[11]) ? node5218 : 14'b00000001111111;
											assign node5218 = (inp[8]) ? node5222 : node5219;
												assign node5219 = (inp[2]) ? 14'b00000000111111 : 14'b00000001111111;
												assign node5222 = (inp[3]) ? 14'b00000000011111 : 14'b00000000111111;
										assign node5225 = (inp[3]) ? node5233 : node5226;
											assign node5226 = (inp[2]) ? node5230 : node5227;
												assign node5227 = (inp[11]) ? 14'b00000000111111 : 14'b00000001111111;
												assign node5230 = (inp[11]) ? 14'b00000000011111 : 14'b00000000111111;
											assign node5233 = (inp[8]) ? 14'b00000000011111 : node5234;
												assign node5234 = (inp[11]) ? 14'b00000000001111 : 14'b00000000011111;
								assign node5238 = (inp[6]) ? node5264 : node5239;
									assign node5239 = (inp[2]) ? node5251 : node5240;
										assign node5240 = (inp[12]) ? node5246 : node5241;
											assign node5241 = (inp[9]) ? node5243 : 14'b00000001111111;
												assign node5243 = (inp[11]) ? 14'b00000000111111 : 14'b00000000111111;
											assign node5246 = (inp[3]) ? 14'b00000000111111 : node5247;
												assign node5247 = (inp[8]) ? 14'b00000000111111 : 14'b00000001111111;
										assign node5251 = (inp[12]) ? node5257 : node5252;
											assign node5252 = (inp[11]) ? 14'b00000000011111 : node5253;
												assign node5253 = (inp[8]) ? 14'b00000000111111 : 14'b00000001111111;
											assign node5257 = (inp[9]) ? node5261 : node5258;
												assign node5258 = (inp[8]) ? 14'b00000000011111 : 14'b00000000111111;
												assign node5261 = (inp[3]) ? 14'b00000000001111 : 14'b00000000001111;
									assign node5264 = (inp[11]) ? node5276 : node5265;
										assign node5265 = (inp[8]) ? node5271 : node5266;
											assign node5266 = (inp[2]) ? 14'b00000000011111 : node5267;
												assign node5267 = (inp[3]) ? 14'b00000000011111 : 14'b00000000111111;
											assign node5271 = (inp[12]) ? node5273 : 14'b00000000011111;
												assign node5273 = (inp[3]) ? 14'b00000000001111 : 14'b00000000011111;
										assign node5276 = (inp[9]) ? 14'b00000000001111 : node5277;
											assign node5277 = (inp[2]) ? 14'b00000000001111 : 14'b00000000011111;
					assign node5281 = (inp[2]) ? node5479 : node5282;
						assign node5282 = (inp[9]) ? node5388 : node5283;
							assign node5283 = (inp[7]) ? node5337 : node5284;
								assign node5284 = (inp[11]) ? node5314 : node5285;
									assign node5285 = (inp[10]) ? node5301 : node5286;
										assign node5286 = (inp[6]) ? node5294 : node5287;
											assign node5287 = (inp[3]) ? node5291 : node5288;
												assign node5288 = (inp[8]) ? 14'b00001111111111 : 14'b00000111111111;
												assign node5291 = (inp[8]) ? 14'b00000011111111 : 14'b00000111111111;
											assign node5294 = (inp[8]) ? node5298 : node5295;
												assign node5295 = (inp[0]) ? 14'b00000011111111 : 14'b00000111111111;
												assign node5298 = (inp[0]) ? 14'b00000001111111 : 14'b00000011111111;
										assign node5301 = (inp[6]) ? node5309 : node5302;
											assign node5302 = (inp[8]) ? node5306 : node5303;
												assign node5303 = (inp[0]) ? 14'b00000011111111 : 14'b00000111111111;
												assign node5306 = (inp[3]) ? 14'b00000001111111 : 14'b00000011111111;
											assign node5309 = (inp[12]) ? node5311 : 14'b00000011111111;
												assign node5311 = (inp[3]) ? 14'b00000000111111 : 14'b00000001111111;
									assign node5314 = (inp[8]) ? node5324 : node5315;
										assign node5315 = (inp[6]) ? node5319 : node5316;
											assign node5316 = (inp[0]) ? 14'b00000011111111 : 14'b00000111111111;
											assign node5319 = (inp[10]) ? 14'b00000001111111 : node5320;
												assign node5320 = (inp[3]) ? 14'b00000001111111 : 14'b00000011111111;
										assign node5324 = (inp[3]) ? node5330 : node5325;
											assign node5325 = (inp[0]) ? 14'b00000001111111 : node5326;
												assign node5326 = (inp[6]) ? 14'b00000001111111 : 14'b00000011111111;
											assign node5330 = (inp[12]) ? node5334 : node5331;
												assign node5331 = (inp[10]) ? 14'b00000000111111 : 14'b00000001111111;
												assign node5334 = (inp[6]) ? 14'b00000000011111 : 14'b00000000111111;
								assign node5337 = (inp[12]) ? node5361 : node5338;
									assign node5338 = (inp[11]) ? node5352 : node5339;
										assign node5339 = (inp[0]) ? node5347 : node5340;
											assign node5340 = (inp[8]) ? node5344 : node5341;
												assign node5341 = (inp[10]) ? 14'b00000011111111 : 14'b00000111111111;
												assign node5344 = (inp[10]) ? 14'b00000001111111 : 14'b00000011111111;
											assign node5347 = (inp[3]) ? 14'b00000000111111 : node5348;
												assign node5348 = (inp[8]) ? 14'b00000001111111 : 14'b00000001111111;
										assign node5352 = (inp[6]) ? node5354 : 14'b00000001111111;
											assign node5354 = (inp[10]) ? node5358 : node5355;
												assign node5355 = (inp[0]) ? 14'b00000000111111 : 14'b00000001111111;
												assign node5358 = (inp[0]) ? 14'b00000000001111 : 14'b00000000111111;
									assign node5361 = (inp[3]) ? node5375 : node5362;
										assign node5362 = (inp[11]) ? node5370 : node5363;
											assign node5363 = (inp[10]) ? node5367 : node5364;
												assign node5364 = (inp[0]) ? 14'b00000001111111 : 14'b00000001111111;
												assign node5367 = (inp[6]) ? 14'b00000000111111 : 14'b00000001111111;
											assign node5370 = (inp[6]) ? node5372 : 14'b00000001111111;
												assign node5372 = (inp[0]) ? 14'b00000000011111 : 14'b00000000111111;
										assign node5375 = (inp[10]) ? node5383 : node5376;
											assign node5376 = (inp[8]) ? node5380 : node5377;
												assign node5377 = (inp[11]) ? 14'b00000000011111 : 14'b00000001111111;
												assign node5380 = (inp[6]) ? 14'b00000000011111 : 14'b00000000111111;
											assign node5383 = (inp[6]) ? node5385 : 14'b00000000011111;
												assign node5385 = (inp[11]) ? 14'b00000000000111 : 14'b00000000011111;
							assign node5388 = (inp[12]) ? node5432 : node5389;
								assign node5389 = (inp[3]) ? node5409 : node5390;
									assign node5390 = (inp[8]) ? node5402 : node5391;
										assign node5391 = (inp[7]) ? node5399 : node5392;
											assign node5392 = (inp[0]) ? node5396 : node5393;
												assign node5393 = (inp[11]) ? 14'b00000011111111 : 14'b00000111111111;
												assign node5396 = (inp[11]) ? 14'b00000001111111 : 14'b00000011111111;
											assign node5399 = (inp[6]) ? 14'b00000000111111 : 14'b00000001111111;
										assign node5402 = (inp[11]) ? node5404 : 14'b00000011111111;
											assign node5404 = (inp[7]) ? 14'b00000000111111 : node5405;
												assign node5405 = (inp[0]) ? 14'b00000000111111 : 14'b00000001111111;
									assign node5409 = (inp[10]) ? node5421 : node5410;
										assign node5410 = (inp[7]) ? node5416 : node5411;
											assign node5411 = (inp[6]) ? node5413 : 14'b00000001111111;
												assign node5413 = (inp[8]) ? 14'b00000000111111 : 14'b00000001111111;
											assign node5416 = (inp[6]) ? node5418 : 14'b00000000111111;
												assign node5418 = (inp[8]) ? 14'b00000000111111 : 14'b00000001111111;
										assign node5421 = (inp[6]) ? node5427 : node5422;
											assign node5422 = (inp[7]) ? 14'b00000000111111 : node5423;
												assign node5423 = (inp[11]) ? 14'b00000000111111 : 14'b00000000111111;
											assign node5427 = (inp[7]) ? node5429 : 14'b00000000011111;
												assign node5429 = (inp[11]) ? 14'b00000000001111 : 14'b00000000111111;
								assign node5432 = (inp[8]) ? node5454 : node5433;
									assign node5433 = (inp[6]) ? node5445 : node5434;
										assign node5434 = (inp[0]) ? node5438 : node5435;
											assign node5435 = (inp[7]) ? 14'b00000000111111 : 14'b00000001111111;
											assign node5438 = (inp[11]) ? node5442 : node5439;
												assign node5439 = (inp[3]) ? 14'b00000000111111 : 14'b00000001111111;
												assign node5442 = (inp[10]) ? 14'b00000000011111 : 14'b00000000111111;
										assign node5445 = (inp[10]) ? node5449 : node5446;
											assign node5446 = (inp[3]) ? 14'b00000000011111 : 14'b00000001111111;
											assign node5449 = (inp[11]) ? node5451 : 14'b00000000011111;
												assign node5451 = (inp[3]) ? 14'b00000000001111 : 14'b00000000011111;
									assign node5454 = (inp[10]) ? node5468 : node5455;
										assign node5455 = (inp[6]) ? node5461 : node5456;
											assign node5456 = (inp[7]) ? node5458 : 14'b00000000111111;
												assign node5458 = (inp[3]) ? 14'b00000000011111 : 14'b00000000111111;
											assign node5461 = (inp[0]) ? node5465 : node5462;
												assign node5462 = (inp[3]) ? 14'b00000000011111 : 14'b00000000011111;
												assign node5465 = (inp[7]) ? 14'b00000000000111 : 14'b00000000001111;
										assign node5468 = (inp[6]) ? node5474 : node5469;
											assign node5469 = (inp[11]) ? node5471 : 14'b00000000011111;
												assign node5471 = (inp[3]) ? 14'b00000000001111 : 14'b00000000011111;
											assign node5474 = (inp[11]) ? 14'b00000000000111 : node5475;
												assign node5475 = (inp[3]) ? 14'b00000000001111 : 14'b00000000011111;
						assign node5479 = (inp[12]) ? node5585 : node5480;
							assign node5480 = (inp[0]) ? node5536 : node5481;
								assign node5481 = (inp[9]) ? node5507 : node5482;
									assign node5482 = (inp[8]) ? node5494 : node5483;
										assign node5483 = (inp[10]) ? node5487 : node5484;
											assign node5484 = (inp[3]) ? 14'b00000011111111 : 14'b00000111111111;
											assign node5487 = (inp[6]) ? node5491 : node5488;
												assign node5488 = (inp[7]) ? 14'b00000001111111 : 14'b00000011111111;
												assign node5491 = (inp[11]) ? 14'b00000000111111 : 14'b00000000111111;
										assign node5494 = (inp[10]) ? node5502 : node5495;
											assign node5495 = (inp[11]) ? node5499 : node5496;
												assign node5496 = (inp[6]) ? 14'b00000001111111 : 14'b00000001111111;
												assign node5499 = (inp[3]) ? 14'b00000000111111 : 14'b00000001111111;
											assign node5502 = (inp[3]) ? 14'b00000001111111 : node5503;
												assign node5503 = (inp[11]) ? 14'b00000000111111 : 14'b00000000111111;
									assign node5507 = (inp[6]) ? node5523 : node5508;
										assign node5508 = (inp[11]) ? node5516 : node5509;
											assign node5509 = (inp[7]) ? node5513 : node5510;
												assign node5510 = (inp[3]) ? 14'b00000001111111 : 14'b00000001111111;
												assign node5513 = (inp[10]) ? 14'b00000000011111 : 14'b00000001111111;
											assign node5516 = (inp[7]) ? node5520 : node5517;
												assign node5517 = (inp[8]) ? 14'b00000000111111 : 14'b00000001111111;
												assign node5520 = (inp[10]) ? 14'b00000000011111 : 14'b00000000111111;
										assign node5523 = (inp[10]) ? node5531 : node5524;
											assign node5524 = (inp[11]) ? node5528 : node5525;
												assign node5525 = (inp[7]) ? 14'b00000000111111 : 14'b00000001111111;
												assign node5528 = (inp[8]) ? 14'b00000000011111 : 14'b00000000011111;
											assign node5531 = (inp[11]) ? node5533 : 14'b00000000011111;
												assign node5533 = (inp[8]) ? 14'b00000000001111 : 14'b00000000011111;
								assign node5536 = (inp[10]) ? node5556 : node5537;
									assign node5537 = (inp[3]) ? node5547 : node5538;
										assign node5538 = (inp[7]) ? node5544 : node5539;
											assign node5539 = (inp[9]) ? node5541 : 14'b00000011111111;
												assign node5541 = (inp[8]) ? 14'b00000000111111 : 14'b00000001111111;
											assign node5544 = (inp[9]) ? 14'b00000000011111 : 14'b00000000111111;
										assign node5547 = (inp[6]) ? 14'b00000000011111 : node5548;
											assign node5548 = (inp[8]) ? node5552 : node5549;
												assign node5549 = (inp[7]) ? 14'b00000000111111 : 14'b00000001111111;
												assign node5552 = (inp[11]) ? 14'b00000000011111 : 14'b00000000111111;
									assign node5556 = (inp[8]) ? node5572 : node5557;
										assign node5557 = (inp[9]) ? node5565 : node5558;
											assign node5558 = (inp[3]) ? node5562 : node5559;
												assign node5559 = (inp[7]) ? 14'b00000000111111 : 14'b00000001111111;
												assign node5562 = (inp[6]) ? 14'b00000000011111 : 14'b00000000111111;
											assign node5565 = (inp[11]) ? node5569 : node5566;
												assign node5566 = (inp[3]) ? 14'b00000000011111 : 14'b00000000011111;
												assign node5569 = (inp[6]) ? 14'b00000000001111 : 14'b00000000011111;
										assign node5572 = (inp[7]) ? node5580 : node5573;
											assign node5573 = (inp[3]) ? node5577 : node5574;
												assign node5574 = (inp[6]) ? 14'b00000000011111 : 14'b00000000111111;
												assign node5577 = (inp[6]) ? 14'b00000000001111 : 14'b00000000011111;
											assign node5580 = (inp[9]) ? node5582 : 14'b00000000001111;
												assign node5582 = (inp[11]) ? 14'b00000000000111 : 14'b00000000000111;
							assign node5585 = (inp[9]) ? node5637 : node5586;
								assign node5586 = (inp[6]) ? node5614 : node5587;
									assign node5587 = (inp[0]) ? node5603 : node5588;
										assign node5588 = (inp[7]) ? node5596 : node5589;
											assign node5589 = (inp[10]) ? node5593 : node5590;
												assign node5590 = (inp[3]) ? 14'b00000001111111 : 14'b00000011111111;
												assign node5593 = (inp[11]) ? 14'b00000000111111 : 14'b00000001111111;
											assign node5596 = (inp[11]) ? node5600 : node5597;
												assign node5597 = (inp[8]) ? 14'b00000000111111 : 14'b00000001111111;
												assign node5600 = (inp[8]) ? 14'b00000000011111 : 14'b00000000111111;
										assign node5603 = (inp[3]) ? node5609 : node5604;
											assign node5604 = (inp[7]) ? node5606 : 14'b00000000111111;
												assign node5606 = (inp[11]) ? 14'b00000000011111 : 14'b00000000111111;
											assign node5609 = (inp[10]) ? node5611 : 14'b00000000111111;
												assign node5611 = (inp[11]) ? 14'b00000000001111 : 14'b00000000001111;
									assign node5614 = (inp[10]) ? node5626 : node5615;
										assign node5615 = (inp[3]) ? node5621 : node5616;
											assign node5616 = (inp[0]) ? node5618 : 14'b00000000111111;
												assign node5618 = (inp[8]) ? 14'b00000000011111 : 14'b00000000111111;
											assign node5621 = (inp[0]) ? 14'b00000000001111 : node5622;
												assign node5622 = (inp[11]) ? 14'b00000000001111 : 14'b00000000011111;
										assign node5626 = (inp[0]) ? node5632 : node5627;
											assign node5627 = (inp[8]) ? node5629 : 14'b00000000011111;
												assign node5629 = (inp[3]) ? 14'b00000000000111 : 14'b00000000011111;
											assign node5632 = (inp[7]) ? 14'b00000000001111 : node5633;
												assign node5633 = (inp[11]) ? 14'b00000000001111 : 14'b00000000011111;
								assign node5637 = (inp[11]) ? node5665 : node5638;
									assign node5638 = (inp[7]) ? node5650 : node5639;
										assign node5639 = (inp[8]) ? node5645 : node5640;
											assign node5640 = (inp[0]) ? 14'b00000000001111 : node5641;
												assign node5641 = (inp[10]) ? 14'b00000000111111 : 14'b00000001111111;
											assign node5645 = (inp[0]) ? node5647 : 14'b00000000011111;
												assign node5647 = (inp[3]) ? 14'b00000000001111 : 14'b00000000011111;
										assign node5650 = (inp[3]) ? node5658 : node5651;
											assign node5651 = (inp[10]) ? node5655 : node5652;
												assign node5652 = (inp[6]) ? 14'b00000000011111 : 14'b00000000111111;
												assign node5655 = (inp[8]) ? 14'b00000000001111 : 14'b00000000011111;
											assign node5658 = (inp[6]) ? node5662 : node5659;
												assign node5659 = (inp[10]) ? 14'b00000000001111 : 14'b00000000011111;
												assign node5662 = (inp[8]) ? 14'b00000000000111 : 14'b00000000001111;
									assign node5665 = (inp[8]) ? node5679 : node5666;
										assign node5666 = (inp[10]) ? node5672 : node5667;
											assign node5667 = (inp[6]) ? node5669 : 14'b00000000011111;
												assign node5669 = (inp[3]) ? 14'b00000000001111 : 14'b00000000011111;
											assign node5672 = (inp[6]) ? node5676 : node5673;
												assign node5673 = (inp[3]) ? 14'b00000000001111 : 14'b00000000001111;
												assign node5676 = (inp[3]) ? 14'b00000000000111 : 14'b00000000000111;
										assign node5679 = (inp[10]) ? node5685 : node5680;
											assign node5680 = (inp[7]) ? node5682 : 14'b00000000001111;
												assign node5682 = (inp[6]) ? 14'b00000000000111 : 14'b00000000000111;
											assign node5685 = (inp[6]) ? node5687 : 14'b00000000000111;
												assign node5687 = (inp[3]) ? 14'b00000000000011 : 14'b00000000000011;
				assign node5690 = (inp[3]) ? node6086 : node5691;
					assign node5691 = (inp[10]) ? node5879 : node5692;
						assign node5692 = (inp[13]) ? node5786 : node5693;
							assign node5693 = (inp[9]) ? node5743 : node5694;
								assign node5694 = (inp[7]) ? node5716 : node5695;
									assign node5695 = (inp[2]) ? node5707 : node5696;
										assign node5696 = (inp[0]) ? node5702 : node5697;
											assign node5697 = (inp[11]) ? node5699 : 14'b00000111111111;
												assign node5699 = (inp[6]) ? 14'b00000011111111 : 14'b00000111111111;
											assign node5702 = (inp[11]) ? 14'b00000011111111 : node5703;
												assign node5703 = (inp[8]) ? 14'b00000011111111 : 14'b00000111111111;
										assign node5707 = (inp[0]) ? 14'b00000001111111 : node5708;
											assign node5708 = (inp[6]) ? node5712 : node5709;
												assign node5709 = (inp[11]) ? 14'b00000011111111 : 14'b00000111111111;
												assign node5712 = (inp[11]) ? 14'b00000001111111 : 14'b00000011111111;
									assign node5716 = (inp[2]) ? node5730 : node5717;
										assign node5717 = (inp[0]) ? node5723 : node5718;
											assign node5718 = (inp[12]) ? node5720 : 14'b00000111111111;
												assign node5720 = (inp[11]) ? 14'b00000001111111 : 14'b00000111111111;
											assign node5723 = (inp[11]) ? node5727 : node5724;
												assign node5724 = (inp[12]) ? 14'b00000001111111 : 14'b00000011111111;
												assign node5727 = (inp[12]) ? 14'b00000000111111 : 14'b00000001111111;
										assign node5730 = (inp[0]) ? node5738 : node5731;
											assign node5731 = (inp[6]) ? node5735 : node5732;
												assign node5732 = (inp[8]) ? 14'b00000001111111 : 14'b00000011111111;
												assign node5735 = (inp[8]) ? 14'b00000000111111 : 14'b00000001111111;
											assign node5738 = (inp[11]) ? 14'b00000000111111 : node5739;
												assign node5739 = (inp[12]) ? 14'b00000000111111 : 14'b00000011111111;
								assign node5743 = (inp[12]) ? node5765 : node5744;
									assign node5744 = (inp[7]) ? node5758 : node5745;
										assign node5745 = (inp[8]) ? node5751 : node5746;
											assign node5746 = (inp[0]) ? 14'b00000011111111 : node5747;
												assign node5747 = (inp[11]) ? 14'b00000011111111 : 14'b00000111111111;
											assign node5751 = (inp[2]) ? node5755 : node5752;
												assign node5752 = (inp[11]) ? 14'b00000001111111 : 14'b00000011111111;
												assign node5755 = (inp[0]) ? 14'b00000000111111 : 14'b00000001111111;
										assign node5758 = (inp[0]) ? 14'b00000000011111 : node5759;
											assign node5759 = (inp[8]) ? 14'b00000000111111 : node5760;
												assign node5760 = (inp[2]) ? 14'b00000001111111 : 14'b00000001111111;
									assign node5765 = (inp[8]) ? node5779 : node5766;
										assign node5766 = (inp[0]) ? node5772 : node5767;
											assign node5767 = (inp[11]) ? 14'b00000001111111 : node5768;
												assign node5768 = (inp[6]) ? 14'b00000001111111 : 14'b00000011111111;
											assign node5772 = (inp[2]) ? node5776 : node5773;
												assign node5773 = (inp[7]) ? 14'b00000000111111 : 14'b00000011111111;
												assign node5776 = (inp[6]) ? 14'b00000000001111 : 14'b00000000111111;
										assign node5779 = (inp[6]) ? node5781 : 14'b00000000111111;
											assign node5781 = (inp[0]) ? 14'b00000000011111 : node5782;
												assign node5782 = (inp[2]) ? 14'b00000000011111 : 14'b00000000111111;
							assign node5786 = (inp[2]) ? node5834 : node5787;
								assign node5787 = (inp[6]) ? node5815 : node5788;
									assign node5788 = (inp[9]) ? node5802 : node5789;
										assign node5789 = (inp[0]) ? node5795 : node5790;
											assign node5790 = (inp[11]) ? node5792 : 14'b00000011111111;
												assign node5792 = (inp[7]) ? 14'b00000001111111 : 14'b00000011111111;
											assign node5795 = (inp[12]) ? node5799 : node5796;
												assign node5796 = (inp[8]) ? 14'b00000001111111 : 14'b00000011111111;
												assign node5799 = (inp[8]) ? 14'b00000000111111 : 14'b00000001111111;
										assign node5802 = (inp[8]) ? node5810 : node5803;
											assign node5803 = (inp[0]) ? node5807 : node5804;
												assign node5804 = (inp[12]) ? 14'b00000001111111 : 14'b00000011111111;
												assign node5807 = (inp[11]) ? 14'b00000000111111 : 14'b00000011111111;
											assign node5810 = (inp[0]) ? 14'b00000000111111 : node5811;
												assign node5811 = (inp[7]) ? 14'b00000000111111 : 14'b00000000111111;
									assign node5815 = (inp[7]) ? node5821 : node5816;
										assign node5816 = (inp[11]) ? 14'b00000001111111 : node5817;
											assign node5817 = (inp[0]) ? 14'b00000001111111 : 14'b00000011111111;
										assign node5821 = (inp[11]) ? node5829 : node5822;
											assign node5822 = (inp[12]) ? node5826 : node5823;
												assign node5823 = (inp[0]) ? 14'b00000000111111 : 14'b00000001111111;
												assign node5826 = (inp[8]) ? 14'b00000000001111 : 14'b00000000111111;
											assign node5829 = (inp[12]) ? 14'b00000000011111 : node5830;
												assign node5830 = (inp[9]) ? 14'b00000000011111 : 14'b00000000111111;
								assign node5834 = (inp[9]) ? node5858 : node5835;
									assign node5835 = (inp[6]) ? node5849 : node5836;
										assign node5836 = (inp[11]) ? node5842 : node5837;
											assign node5837 = (inp[8]) ? 14'b00000000111111 : node5838;
												assign node5838 = (inp[0]) ? 14'b00000001111111 : 14'b00000011111111;
											assign node5842 = (inp[0]) ? node5846 : node5843;
												assign node5843 = (inp[12]) ? 14'b00000000111111 : 14'b00000000111111;
												assign node5846 = (inp[12]) ? 14'b00000000011111 : 14'b00000000111111;
										assign node5849 = (inp[0]) ? node5851 : 14'b00000000111111;
											assign node5851 = (inp[11]) ? node5855 : node5852;
												assign node5852 = (inp[7]) ? 14'b00000000011111 : 14'b00000000111111;
												assign node5855 = (inp[8]) ? 14'b00000000000111 : 14'b00000000011111;
									assign node5858 = (inp[8]) ? node5868 : node5859;
										assign node5859 = (inp[12]) ? node5865 : node5860;
											assign node5860 = (inp[0]) ? node5862 : 14'b00000000111111;
												assign node5862 = (inp[7]) ? 14'b00000000011111 : 14'b00000000111111;
											assign node5865 = (inp[11]) ? 14'b00000000000111 : 14'b00000000011111;
										assign node5868 = (inp[12]) ? node5874 : node5869;
											assign node5869 = (inp[6]) ? node5871 : 14'b00000000011111;
												assign node5871 = (inp[11]) ? 14'b00000000000111 : 14'b00000000001111;
											assign node5874 = (inp[11]) ? node5876 : 14'b00000000001111;
												assign node5876 = (inp[0]) ? 14'b00000000000111 : 14'b00000000001111;
						assign node5879 = (inp[9]) ? node5985 : node5880;
							assign node5880 = (inp[8]) ? node5934 : node5881;
								assign node5881 = (inp[11]) ? node5905 : node5882;
									assign node5882 = (inp[6]) ? node5892 : node5883;
										assign node5883 = (inp[7]) ? node5885 : 14'b00000011111111;
											assign node5885 = (inp[0]) ? node5889 : node5886;
												assign node5886 = (inp[2]) ? 14'b00000001111111 : 14'b00000011111111;
												assign node5889 = (inp[12]) ? 14'b00000000111111 : 14'b00000001111111;
										assign node5892 = (inp[13]) ? node5900 : node5893;
											assign node5893 = (inp[0]) ? node5897 : node5894;
												assign node5894 = (inp[7]) ? 14'b00000001111111 : 14'b00000011111111;
												assign node5897 = (inp[7]) ? 14'b00000000111111 : 14'b00000001111111;
											assign node5900 = (inp[0]) ? 14'b00000000011111 : node5901;
												assign node5901 = (inp[2]) ? 14'b00000000111111 : 14'b00000001111111;
									assign node5905 = (inp[6]) ? node5921 : node5906;
										assign node5906 = (inp[12]) ? node5914 : node5907;
											assign node5907 = (inp[13]) ? node5911 : node5908;
												assign node5908 = (inp[2]) ? 14'b00000001111111 : 14'b00000011111111;
												assign node5911 = (inp[2]) ? 14'b00000000111111 : 14'b00000000111111;
											assign node5914 = (inp[7]) ? node5918 : node5915;
												assign node5915 = (inp[0]) ? 14'b00000000111111 : 14'b00000001111111;
												assign node5918 = (inp[13]) ? 14'b00000000011111 : 14'b00000000111111;
										assign node5921 = (inp[13]) ? node5929 : node5922;
											assign node5922 = (inp[7]) ? node5926 : node5923;
												assign node5923 = (inp[2]) ? 14'b00000000111111 : 14'b00000001111111;
												assign node5926 = (inp[0]) ? 14'b00000000011111 : 14'b00000000111111;
											assign node5929 = (inp[7]) ? 14'b00000000011111 : node5930;
												assign node5930 = (inp[0]) ? 14'b00000000011111 : 14'b00000000111111;
								assign node5934 = (inp[12]) ? node5964 : node5935;
									assign node5935 = (inp[11]) ? node5951 : node5936;
										assign node5936 = (inp[2]) ? node5944 : node5937;
											assign node5937 = (inp[0]) ? node5941 : node5938;
												assign node5938 = (inp[13]) ? 14'b00000001111111 : 14'b00000001111111;
												assign node5941 = (inp[7]) ? 14'b00000000111111 : 14'b00000001111111;
											assign node5944 = (inp[6]) ? node5948 : node5945;
												assign node5945 = (inp[0]) ? 14'b00000000111111 : 14'b00000001111111;
												assign node5948 = (inp[7]) ? 14'b00000000011111 : 14'b00000000111111;
										assign node5951 = (inp[6]) ? node5959 : node5952;
											assign node5952 = (inp[0]) ? node5956 : node5953;
												assign node5953 = (inp[7]) ? 14'b00000000111111 : 14'b00000000111111;
												assign node5956 = (inp[7]) ? 14'b00000000011111 : 14'b00000000111111;
											assign node5959 = (inp[2]) ? node5961 : 14'b00000000111111;
												assign node5961 = (inp[0]) ? 14'b00000000001111 : 14'b00000000011111;
									assign node5964 = (inp[2]) ? node5974 : node5965;
										assign node5965 = (inp[11]) ? node5971 : node5966;
											assign node5966 = (inp[7]) ? node5968 : 14'b00000000111111;
												assign node5968 = (inp[0]) ? 14'b00000000011111 : 14'b00000000111111;
											assign node5971 = (inp[13]) ? 14'b00000000011111 : 14'b00000000001111;
										assign node5974 = (inp[6]) ? node5978 : node5975;
											assign node5975 = (inp[0]) ? 14'b00000000001111 : 14'b00000000111111;
											assign node5978 = (inp[7]) ? node5982 : node5979;
												assign node5979 = (inp[11]) ? 14'b00000000001111 : 14'b00000000011111;
												assign node5982 = (inp[13]) ? 14'b00000000000111 : 14'b00000000000111;
							assign node5985 = (inp[7]) ? node6035 : node5986;
								assign node5986 = (inp[6]) ? node6014 : node5987;
									assign node5987 = (inp[11]) ? node6001 : node5988;
										assign node5988 = (inp[0]) ? node5994 : node5989;
											assign node5989 = (inp[13]) ? 14'b00000001111111 : node5990;
												assign node5990 = (inp[8]) ? 14'b00000001111111 : 14'b00000011111111;
											assign node5994 = (inp[13]) ? node5998 : node5995;
												assign node5995 = (inp[12]) ? 14'b00000000111111 : 14'b00000011111111;
												assign node5998 = (inp[8]) ? 14'b00000000011111 : 14'b00000000111111;
										assign node6001 = (inp[2]) ? node6009 : node6002;
											assign node6002 = (inp[13]) ? node6006 : node6003;
												assign node6003 = (inp[0]) ? 14'b00000000111111 : 14'b00000001111111;
												assign node6006 = (inp[8]) ? 14'b00000000011111 : 14'b00000000011111;
											assign node6009 = (inp[0]) ? node6011 : 14'b00000000011111;
												assign node6011 = (inp[8]) ? 14'b00000000001111 : 14'b00000000011111;
									assign node6014 = (inp[11]) ? node6026 : node6015;
										assign node6015 = (inp[12]) ? node6021 : node6016;
											assign node6016 = (inp[2]) ? node6018 : 14'b00000001111111;
												assign node6018 = (inp[0]) ? 14'b00000000011111 : 14'b00000000111111;
											assign node6021 = (inp[2]) ? node6023 : 14'b00000000011111;
												assign node6023 = (inp[13]) ? 14'b00000000001111 : 14'b00000000011111;
										assign node6026 = (inp[13]) ? node6030 : node6027;
											assign node6027 = (inp[2]) ? 14'b00000000001111 : 14'b00000000011111;
											assign node6030 = (inp[8]) ? node6032 : 14'b00000000001111;
												assign node6032 = (inp[12]) ? 14'b00000000000011 : 14'b00000000000111;
								assign node6035 = (inp[13]) ? node6059 : node6036;
									assign node6036 = (inp[2]) ? node6046 : node6037;
										assign node6037 = (inp[8]) ? node6039 : 14'b00000000111111;
											assign node6039 = (inp[6]) ? node6043 : node6040;
												assign node6040 = (inp[11]) ? 14'b00000000011111 : 14'b00000000111111;
												assign node6043 = (inp[0]) ? 14'b00000000001111 : 14'b00000000011111;
										assign node6046 = (inp[8]) ? node6054 : node6047;
											assign node6047 = (inp[6]) ? node6051 : node6048;
												assign node6048 = (inp[11]) ? 14'b00000000011111 : 14'b00000000111111;
												assign node6051 = (inp[11]) ? 14'b00000000001111 : 14'b00000000011111;
											assign node6054 = (inp[6]) ? node6056 : 14'b00000000001111;
												assign node6056 = (inp[0]) ? 14'b00000000000111 : 14'b00000000000111;
									assign node6059 = (inp[8]) ? node6073 : node6060;
										assign node6060 = (inp[6]) ? node6066 : node6061;
											assign node6061 = (inp[12]) ? node6063 : 14'b00000000011111;
												assign node6063 = (inp[11]) ? 14'b00000000000111 : 14'b00000000011111;
											assign node6066 = (inp[0]) ? node6070 : node6067;
												assign node6067 = (inp[2]) ? 14'b00000000001111 : 14'b00000000001111;
												assign node6070 = (inp[12]) ? 14'b00000000000111 : 14'b00000000001111;
										assign node6073 = (inp[2]) ? node6079 : node6074;
											assign node6074 = (inp[12]) ? node6076 : 14'b00000000001111;
												assign node6076 = (inp[11]) ? 14'b00000000000111 : 14'b00000000001111;
											assign node6079 = (inp[12]) ? node6083 : node6080;
												assign node6080 = (inp[6]) ? 14'b00000000000111 : 14'b00000000000111;
												assign node6083 = (inp[0]) ? 14'b00000000000001 : 14'b00000000000111;
					assign node6086 = (inp[9]) ? node6272 : node6087;
						assign node6087 = (inp[10]) ? node6171 : node6088;
							assign node6088 = (inp[12]) ? node6132 : node6089;
								assign node6089 = (inp[6]) ? node6111 : node6090;
									assign node6090 = (inp[0]) ? node6096 : node6091;
										assign node6091 = (inp[11]) ? 14'b00000001111111 : node6092;
											assign node6092 = (inp[8]) ? 14'b00000001111111 : 14'b00000111111111;
										assign node6096 = (inp[13]) ? node6104 : node6097;
											assign node6097 = (inp[8]) ? node6101 : node6098;
												assign node6098 = (inp[2]) ? 14'b00000001111111 : 14'b00000011111111;
												assign node6101 = (inp[7]) ? 14'b00000000111111 : 14'b00000001111111;
											assign node6104 = (inp[11]) ? node6108 : node6105;
												assign node6105 = (inp[2]) ? 14'b00000000111111 : 14'b00000001111111;
												assign node6108 = (inp[7]) ? 14'b00000000011111 : 14'b00000000111111;
									assign node6111 = (inp[7]) ? node6119 : node6112;
										assign node6112 = (inp[13]) ? 14'b00000000111111 : node6113;
											assign node6113 = (inp[11]) ? node6115 : 14'b00000011111111;
												assign node6115 = (inp[2]) ? 14'b00000000111111 : 14'b00000001111111;
										assign node6119 = (inp[0]) ? node6125 : node6120;
											assign node6120 = (inp[8]) ? 14'b00000000011111 : node6121;
												assign node6121 = (inp[11]) ? 14'b00000000011111 : 14'b00000001111111;
											assign node6125 = (inp[11]) ? node6129 : node6126;
												assign node6126 = (inp[2]) ? 14'b00000000011111 : 14'b00000000111111;
												assign node6129 = (inp[13]) ? 14'b00000000001111 : 14'b00000000011111;
								assign node6132 = (inp[11]) ? node6152 : node6133;
									assign node6133 = (inp[2]) ? node6141 : node6134;
										assign node6134 = (inp[7]) ? node6136 : 14'b00000001111111;
											assign node6136 = (inp[13]) ? 14'b00000000111111 : node6137;
												assign node6137 = (inp[8]) ? 14'b00000000111111 : 14'b00000001111111;
										assign node6141 = (inp[8]) ? node6147 : node6142;
											assign node6142 = (inp[6]) ? node6144 : 14'b00000000111111;
												assign node6144 = (inp[7]) ? 14'b00000000011111 : 14'b00000000111111;
											assign node6147 = (inp[6]) ? node6149 : 14'b00000000011111;
												assign node6149 = (inp[13]) ? 14'b00000000001111 : 14'b00000000011111;
									assign node6152 = (inp[2]) ? node6164 : node6153;
										assign node6153 = (inp[13]) ? node6159 : node6154;
											assign node6154 = (inp[6]) ? node6156 : 14'b00000000111111;
												assign node6156 = (inp[7]) ? 14'b00000000001111 : 14'b00000000011111;
											assign node6159 = (inp[7]) ? node6161 : 14'b00000000011111;
												assign node6161 = (inp[0]) ? 14'b00000000011111 : 14'b00000000001111;
										assign node6164 = (inp[0]) ? 14'b00000000001111 : node6165;
											assign node6165 = (inp[6]) ? node6167 : 14'b00000000011111;
												assign node6167 = (inp[7]) ? 14'b00000000001111 : 14'b00000000011111;
							assign node6171 = (inp[2]) ? node6227 : node6172;
								assign node6172 = (inp[7]) ? node6198 : node6173;
									assign node6173 = (inp[12]) ? node6185 : node6174;
										assign node6174 = (inp[6]) ? node6180 : node6175;
											assign node6175 = (inp[0]) ? node6177 : 14'b00000001111111;
												assign node6177 = (inp[8]) ? 14'b00000000111111 : 14'b00000000111111;
											assign node6180 = (inp[11]) ? node6182 : 14'b00000000111111;
												assign node6182 = (inp[0]) ? 14'b00000000001111 : 14'b00000000111111;
										assign node6185 = (inp[0]) ? node6191 : node6186;
											assign node6186 = (inp[8]) ? 14'b00000000111111 : node6187;
												assign node6187 = (inp[13]) ? 14'b00000000011111 : 14'b00000000111111;
											assign node6191 = (inp[8]) ? node6195 : node6192;
												assign node6192 = (inp[11]) ? 14'b00000000011111 : 14'b00000000111111;
												assign node6195 = (inp[13]) ? 14'b00000000001111 : 14'b00000000011111;
									assign node6198 = (inp[12]) ? node6212 : node6199;
										assign node6199 = (inp[13]) ? node6205 : node6200;
											assign node6200 = (inp[6]) ? node6202 : 14'b00000000111111;
												assign node6202 = (inp[8]) ? 14'b00000000011111 : 14'b00000000111111;
											assign node6205 = (inp[11]) ? node6209 : node6206;
												assign node6206 = (inp[8]) ? 14'b00000000011111 : 14'b00000000111111;
												assign node6209 = (inp[8]) ? 14'b00000000001111 : 14'b00000000011111;
										assign node6212 = (inp[8]) ? node6220 : node6213;
											assign node6213 = (inp[0]) ? node6217 : node6214;
												assign node6214 = (inp[13]) ? 14'b00000000011111 : 14'b00000000111111;
												assign node6217 = (inp[6]) ? 14'b00000000001111 : 14'b00000000011111;
											assign node6220 = (inp[13]) ? node6224 : node6221;
												assign node6221 = (inp[6]) ? 14'b00000000001111 : 14'b00000000001111;
												assign node6224 = (inp[11]) ? 14'b00000000000111 : 14'b00000000000111;
								assign node6227 = (inp[6]) ? node6243 : node6228;
									assign node6228 = (inp[11]) ? node6236 : node6229;
										assign node6229 = (inp[0]) ? node6231 : 14'b00000001111111;
											assign node6231 = (inp[8]) ? 14'b00000000011111 : node6232;
												assign node6232 = (inp[12]) ? 14'b00000000011111 : 14'b00000000111111;
										assign node6236 = (inp[12]) ? node6238 : 14'b00000000011111;
											assign node6238 = (inp[8]) ? 14'b00000000001111 : node6239;
												assign node6239 = (inp[13]) ? 14'b00000000001111 : 14'b00000000011111;
									assign node6243 = (inp[0]) ? node6257 : node6244;
										assign node6244 = (inp[7]) ? node6250 : node6245;
											assign node6245 = (inp[8]) ? 14'b00000000001111 : node6246;
												assign node6246 = (inp[12]) ? 14'b00000000111111 : 14'b00000000011111;
											assign node6250 = (inp[12]) ? node6254 : node6251;
												assign node6251 = (inp[8]) ? 14'b00000000001111 : 14'b00000000001111;
												assign node6254 = (inp[11]) ? 14'b00000000000111 : 14'b00000000001111;
										assign node6257 = (inp[13]) ? node6265 : node6258;
											assign node6258 = (inp[7]) ? node6262 : node6259;
												assign node6259 = (inp[8]) ? 14'b00000000001111 : 14'b00000000011111;
												assign node6262 = (inp[11]) ? 14'b00000000000111 : 14'b00000000001111;
											assign node6265 = (inp[12]) ? node6269 : node6266;
												assign node6266 = (inp[11]) ? 14'b00000000000111 : 14'b00000000001111;
												assign node6269 = (inp[8]) ? 14'b00000000000011 : 14'b00000000000111;
						assign node6272 = (inp[2]) ? node6372 : node6273;
							assign node6273 = (inp[6]) ? node6325 : node6274;
								assign node6274 = (inp[0]) ? node6304 : node6275;
									assign node6275 = (inp[11]) ? node6289 : node6276;
										assign node6276 = (inp[7]) ? node6282 : node6277;
											assign node6277 = (inp[10]) ? node6279 : 14'b00000011111111;
												assign node6279 = (inp[8]) ? 14'b00000001111111 : 14'b00000001111111;
											assign node6282 = (inp[12]) ? node6286 : node6283;
												assign node6283 = (inp[13]) ? 14'b00000000111111 : 14'b00000001111111;
												assign node6286 = (inp[10]) ? 14'b00000000011111 : 14'b00000000111111;
										assign node6289 = (inp[13]) ? node6297 : node6290;
											assign node6290 = (inp[7]) ? node6294 : node6291;
												assign node6291 = (inp[12]) ? 14'b00000000111111 : 14'b00000001111111;
												assign node6294 = (inp[8]) ? 14'b00000000011111 : 14'b00000000111111;
											assign node6297 = (inp[10]) ? node6301 : node6298;
												assign node6298 = (inp[12]) ? 14'b00000000011111 : 14'b00000000111111;
												assign node6301 = (inp[8]) ? 14'b00000000000111 : 14'b00000000011111;
									assign node6304 = (inp[8]) ? node6318 : node6305;
										assign node6305 = (inp[10]) ? node6313 : node6306;
											assign node6306 = (inp[11]) ? node6310 : node6307;
												assign node6307 = (inp[7]) ? 14'b00000000111111 : 14'b00000001111111;
												assign node6310 = (inp[7]) ? 14'b00000000011111 : 14'b00000000011111;
											assign node6313 = (inp[12]) ? node6315 : 14'b00000000011111;
												assign node6315 = (inp[13]) ? 14'b00000000001111 : 14'b00000000011111;
										assign node6318 = (inp[12]) ? node6320 : 14'b00000000011111;
											assign node6320 = (inp[10]) ? 14'b00000000001111 : node6321;
												assign node6321 = (inp[7]) ? 14'b00000000000111 : 14'b00000000001111;
								assign node6325 = (inp[10]) ? node6351 : node6326;
									assign node6326 = (inp[8]) ? node6338 : node6327;
										assign node6327 = (inp[0]) ? node6333 : node6328;
											assign node6328 = (inp[12]) ? node6330 : 14'b00000000111111;
												assign node6330 = (inp[11]) ? 14'b00000000011111 : 14'b00000000111111;
											assign node6333 = (inp[11]) ? 14'b00000000011111 : node6334;
												assign node6334 = (inp[13]) ? 14'b00000000011111 : 14'b00000000011111;
										assign node6338 = (inp[7]) ? node6344 : node6339;
											assign node6339 = (inp[12]) ? 14'b00000000011111 : node6340;
												assign node6340 = (inp[13]) ? 14'b00000000011111 : 14'b00000000111111;
											assign node6344 = (inp[11]) ? node6348 : node6345;
												assign node6345 = (inp[13]) ? 14'b00000000001111 : 14'b00000000011111;
												assign node6348 = (inp[12]) ? 14'b00000000000111 : 14'b00000000001111;
									assign node6351 = (inp[13]) ? node6361 : node6352;
										assign node6352 = (inp[11]) ? node6356 : node6353;
											assign node6353 = (inp[0]) ? 14'b00000000001111 : 14'b00000000011111;
											assign node6356 = (inp[8]) ? 14'b00000000000111 : node6357;
												assign node6357 = (inp[7]) ? 14'b00000000000111 : 14'b00000000001111;
										assign node6361 = (inp[0]) ? node6367 : node6362;
											assign node6362 = (inp[8]) ? node6364 : 14'b00000000001111;
												assign node6364 = (inp[7]) ? 14'b00000000000111 : 14'b00000000000111;
											assign node6367 = (inp[8]) ? node6369 : 14'b00000000000111;
												assign node6369 = (inp[7]) ? 14'b00000000000001 : 14'b00000000000011;
							assign node6372 = (inp[11]) ? node6430 : node6373;
								assign node6373 = (inp[7]) ? node6401 : node6374;
									assign node6374 = (inp[10]) ? node6388 : node6375;
										assign node6375 = (inp[12]) ? node6381 : node6376;
											assign node6376 = (inp[8]) ? 14'b00000000111111 : node6377;
												assign node6377 = (inp[6]) ? 14'b00000000011111 : 14'b00000001111111;
											assign node6381 = (inp[0]) ? node6385 : node6382;
												assign node6382 = (inp[13]) ? 14'b00000000011111 : 14'b00000000111111;
												assign node6385 = (inp[13]) ? 14'b00000000001111 : 14'b00000000011111;
										assign node6388 = (inp[8]) ? node6396 : node6389;
											assign node6389 = (inp[0]) ? node6393 : node6390;
												assign node6390 = (inp[6]) ? 14'b00000000011111 : 14'b00000000111111;
												assign node6393 = (inp[6]) ? 14'b00000000001111 : 14'b00000000011111;
											assign node6396 = (inp[12]) ? node6398 : 14'b00000000011111;
												assign node6398 = (inp[13]) ? 14'b00000000000111 : 14'b00000000000111;
									assign node6401 = (inp[8]) ? node6415 : node6402;
										assign node6402 = (inp[12]) ? node6408 : node6403;
											assign node6403 = (inp[13]) ? node6405 : 14'b00000000111111;
												assign node6405 = (inp[6]) ? 14'b00000000001111 : 14'b00000000011111;
											assign node6408 = (inp[6]) ? node6412 : node6409;
												assign node6409 = (inp[13]) ? 14'b00000000001111 : 14'b00000000011111;
												assign node6412 = (inp[0]) ? 14'b00000000000111 : 14'b00000000001111;
										assign node6415 = (inp[13]) ? node6423 : node6416;
											assign node6416 = (inp[12]) ? node6420 : node6417;
												assign node6417 = (inp[6]) ? 14'b00000000001111 : 14'b00000000011111;
												assign node6420 = (inp[6]) ? 14'b00000000000111 : 14'b00000000000111;
											assign node6423 = (inp[0]) ? node6427 : node6424;
												assign node6424 = (inp[10]) ? 14'b00000000000111 : 14'b00000000001111;
												assign node6427 = (inp[12]) ? 14'b00000000000011 : 14'b00000000000111;
								assign node6430 = (inp[12]) ? node6458 : node6431;
									assign node6431 = (inp[7]) ? node6447 : node6432;
										assign node6432 = (inp[13]) ? node6440 : node6433;
											assign node6433 = (inp[8]) ? node6437 : node6434;
												assign node6434 = (inp[0]) ? 14'b00000000011111 : 14'b00000000111111;
												assign node6437 = (inp[6]) ? 14'b00000000001111 : 14'b00000000011111;
											assign node6440 = (inp[0]) ? node6444 : node6441;
												assign node6441 = (inp[8]) ? 14'b00000000001111 : 14'b00000000001111;
												assign node6444 = (inp[10]) ? 14'b00000000000111 : 14'b00000000001111;
										assign node6447 = (inp[8]) ? node6453 : node6448;
											assign node6448 = (inp[10]) ? 14'b00000000000111 : node6449;
												assign node6449 = (inp[13]) ? 14'b00000000000111 : 14'b00000000011111;
											assign node6453 = (inp[6]) ? 14'b00000000000011 : node6454;
												assign node6454 = (inp[10]) ? 14'b00000000000011 : 14'b00000000001111;
									assign node6458 = (inp[10]) ? node6470 : node6459;
										assign node6459 = (inp[0]) ? node6465 : node6460;
											assign node6460 = (inp[6]) ? 14'b00000000000111 : node6461;
												assign node6461 = (inp[13]) ? 14'b00000000001111 : 14'b00000000011111;
											assign node6465 = (inp[13]) ? node6467 : 14'b00000000000111;
												assign node6467 = (inp[6]) ? 14'b00000000000001 : 14'b00000000000111;
										assign node6470 = (inp[8]) ? node6476 : node6471;
											assign node6471 = (inp[13]) ? 14'b00000000000011 : node6472;
												assign node6472 = (inp[6]) ? 14'b00000000000011 : 14'b00000000001111;
											assign node6476 = (inp[13]) ? node6478 : 14'b00000000000011;
												assign node6478 = (inp[0]) ? 14'b00000000000001 : 14'b00000000000011;

endmodule