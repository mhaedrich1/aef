module dtc_split33_bm58 (
	input  wire [12-1:0] inp,
	output wire [3-1:0] outp
);

	wire [3-1:0] node2;
	wire [3-1:0] node3;
	wire [3-1:0] node4;
	wire [3-1:0] node5;
	wire [3-1:0] node6;
	wire [3-1:0] node7;
	wire [3-1:0] node8;
	wire [3-1:0] node10;
	wire [3-1:0] node11;
	wire [3-1:0] node12;
	wire [3-1:0] node18;
	wire [3-1:0] node19;
	wire [3-1:0] node21;
	wire [3-1:0] node26;
	wire [3-1:0] node27;
	wire [3-1:0] node28;
	wire [3-1:0] node29;
	wire [3-1:0] node30;
	wire [3-1:0] node31;
	wire [3-1:0] node36;
	wire [3-1:0] node37;
	wire [3-1:0] node39;
	wire [3-1:0] node43;
	wire [3-1:0] node44;
	wire [3-1:0] node45;
	wire [3-1:0] node47;
	wire [3-1:0] node49;
	wire [3-1:0] node52;
	wire [3-1:0] node53;
	wire [3-1:0] node55;
	wire [3-1:0] node59;
	wire [3-1:0] node60;
	wire [3-1:0] node62;
	wire [3-1:0] node66;
	wire [3-1:0] node68;
	wire [3-1:0] node69;
	wire [3-1:0] node70;
	wire [3-1:0] node72;
	wire [3-1:0] node77;
	wire [3-1:0] node78;
	wire [3-1:0] node80;
	wire [3-1:0] node81;
	wire [3-1:0] node82;
	wire [3-1:0] node84;
	wire [3-1:0] node86;
	wire [3-1:0] node90;
	wire [3-1:0] node91;
	wire [3-1:0] node93;
	wire [3-1:0] node94;
	wire [3-1:0] node99;
	wire [3-1:0] node100;
	wire [3-1:0] node101;
	wire [3-1:0] node102;
	wire [3-1:0] node103;
	wire [3-1:0] node104;
	wire [3-1:0] node109;
	wire [3-1:0] node112;
	wire [3-1:0] node113;
	wire [3-1:0] node114;
	wire [3-1:0] node115;
	wire [3-1:0] node120;
	wire [3-1:0] node123;
	wire [3-1:0] node124;
	wire [3-1:0] node125;
	wire [3-1:0] node126;
	wire [3-1:0] node127;
	wire [3-1:0] node131;
	wire [3-1:0] node134;
	wire [3-1:0] node135;
	wire [3-1:0] node138;
	wire [3-1:0] node141;
	wire [3-1:0] node142;
	wire [3-1:0] node143;
	wire [3-1:0] node147;
	wire [3-1:0] node148;
	wire [3-1:0] node152;
	wire [3-1:0] node154;
	wire [3-1:0] node155;
	wire [3-1:0] node156;
	wire [3-1:0] node157;
	wire [3-1:0] node158;
	wire [3-1:0] node160;
	wire [3-1:0] node163;
	wire [3-1:0] node164;
	wire [3-1:0] node165;
	wire [3-1:0] node170;
	wire [3-1:0] node172;
	wire [3-1:0] node174;
	wire [3-1:0] node175;
	wire [3-1:0] node179;
	wire [3-1:0] node180;
	wire [3-1:0] node182;
	wire [3-1:0] node184;
	wire [3-1:0] node186;
	wire [3-1:0] node187;
	wire [3-1:0] node191;
	wire [3-1:0] node192;
	wire [3-1:0] node194;
	wire [3-1:0] node197;
	wire [3-1:0] node198;
	wire [3-1:0] node200;
	wire [3-1:0] node203;
	wire [3-1:0] node204;
	wire [3-1:0] node208;
	wire [3-1:0] node210;
	wire [3-1:0] node211;
	wire [3-1:0] node212;
	wire [3-1:0] node214;
	wire [3-1:0] node217;
	wire [3-1:0] node218;
	wire [3-1:0] node219;
	wire [3-1:0] node220;
	wire [3-1:0] node226;
	wire [3-1:0] node227;
	wire [3-1:0] node229;

	assign outp = (inp[6]) ? node2 : 3'b000;
		assign node2 = (inp[0]) ? node152 : node3;
			assign node3 = (inp[4]) ? node77 : node4;
				assign node4 = (inp[9]) ? node26 : node5;
					assign node5 = (inp[1]) ? 3'b000 : node6;
						assign node6 = (inp[8]) ? node18 : node7;
							assign node7 = (inp[11]) ? 3'b000 : node8;
								assign node8 = (inp[7]) ? node10 : 3'b100;
									assign node10 = (inp[3]) ? 3'b000 : node11;
										assign node11 = (inp[5]) ? 3'b100 : node12;
											assign node12 = (inp[2]) ? 3'b100 : 3'b000;
							assign node18 = (inp[10]) ? 3'b100 : node19;
								assign node19 = (inp[7]) ? node21 : 3'b100;
									assign node21 = (inp[11]) ? 3'b000 : 3'b100;
					assign node26 = (inp[1]) ? node66 : node27;
						assign node27 = (inp[11]) ? node43 : node28;
							assign node28 = (inp[8]) ? node36 : node29;
								assign node29 = (inp[10]) ? 3'b000 : node30;
									assign node30 = (inp[2]) ? 3'b000 : node31;
										assign node31 = (inp[3]) ? 3'b100 : 3'b000;
								assign node36 = (inp[10]) ? 3'b100 : node37;
									assign node37 = (inp[2]) ? node39 : 3'b000;
										assign node39 = (inp[3]) ? 3'b000 : 3'b100;
							assign node43 = (inp[5]) ? node59 : node44;
								assign node44 = (inp[7]) ? node52 : node45;
									assign node45 = (inp[8]) ? node47 : 3'b100;
										assign node47 = (inp[10]) ? node49 : 3'b000;
											assign node49 = (inp[2]) ? 3'b100 : 3'b000;
									assign node52 = (inp[8]) ? 3'b100 : node53;
										assign node53 = (inp[3]) ? node55 : 3'b000;
											assign node55 = (inp[2]) ? 3'b000 : 3'b100;
								assign node59 = (inp[8]) ? 3'b000 : node60;
									assign node60 = (inp[2]) ? node62 : 3'b100;
										assign node62 = (inp[10]) ? 3'b000 : 3'b100;
						assign node66 = (inp[8]) ? node68 : 3'b100;
							assign node68 = (inp[10]) ? 3'b000 : node69;
								assign node69 = (inp[11]) ? 3'b100 : node70;
									assign node70 = (inp[3]) ? node72 : 3'b000;
										assign node72 = (inp[7]) ? 3'b000 : 3'b100;
				assign node77 = (inp[9]) ? node99 : node78;
					assign node78 = (inp[1]) ? node80 : 3'b100;
						assign node80 = (inp[8]) ? node90 : node81;
							assign node81 = (inp[11]) ? 3'b000 : node82;
								assign node82 = (inp[3]) ? node84 : 3'b100;
									assign node84 = (inp[10]) ? node86 : 3'b000;
										assign node86 = (inp[7]) ? 3'b000 : 3'b100;
							assign node90 = (inp[10]) ? 3'b100 : node91;
								assign node91 = (inp[11]) ? node93 : 3'b100;
									assign node93 = (inp[5]) ? 3'b000 : node94;
										assign node94 = (inp[3]) ? 3'b000 : 3'b100;
					assign node99 = (inp[8]) ? node123 : node100;
						assign node100 = (inp[10]) ? node112 : node101;
							assign node101 = (inp[1]) ? node109 : node102;
								assign node102 = (inp[7]) ? 3'b001 : node103;
									assign node103 = (inp[11]) ? 3'b100 : node104;
										assign node104 = (inp[2]) ? 3'b101 : 3'b001;
								assign node109 = (inp[11]) ? 3'b000 : 3'b100;
							assign node112 = (inp[11]) ? node120 : node113;
								assign node113 = (inp[2]) ? 3'b101 : node114;
									assign node114 = (inp[1]) ? 3'b001 : node115;
										assign node115 = (inp[3]) ? 3'b101 : 3'b001;
								assign node120 = (inp[2]) ? 3'b001 : 3'b100;
						assign node123 = (inp[2]) ? node141 : node124;
							assign node124 = (inp[10]) ? node134 : node125;
								assign node125 = (inp[1]) ? node131 : node126;
									assign node126 = (inp[11]) ? 3'b000 : node127;
										assign node127 = (inp[3]) ? 3'b100 : 3'b000;
									assign node131 = (inp[3]) ? 3'b101 : 3'b001;
								assign node134 = (inp[11]) ? node138 : node135;
									assign node135 = (inp[7]) ? 3'b011 : 3'b111;
									assign node138 = (inp[7]) ? 3'b010 : 3'b110;
							assign node141 = (inp[1]) ? node147 : node142;
								assign node142 = (inp[10]) ? 3'b000 : node143;
									assign node143 = (inp[3]) ? 3'b001 : 3'b101;
								assign node147 = (inp[3]) ? 3'b000 : node148;
									assign node148 = (inp[10]) ? 3'b000 : 3'b100;
			assign node152 = (inp[9]) ? node154 : 3'b000;
				assign node154 = (inp[1]) ? node208 : node155;
					assign node155 = (inp[8]) ? node179 : node156;
						assign node156 = (inp[11]) ? node170 : node157;
							assign node157 = (inp[10]) ? node163 : node158;
								assign node158 = (inp[5]) ? node160 : 3'b000;
									assign node160 = (inp[3]) ? 3'b100 : 3'b000;
								assign node163 = (inp[2]) ? 3'b100 : node164;
									assign node164 = (inp[4]) ? 3'b000 : node165;
										assign node165 = (inp[3]) ? 3'b000 : 3'b100;
							assign node170 = (inp[4]) ? node172 : 3'b000;
								assign node172 = (inp[10]) ? node174 : 3'b100;
									assign node174 = (inp[2]) ? 3'b000 : node175;
										assign node175 = (inp[3]) ? 3'b100 : 3'b000;
						assign node179 = (inp[4]) ? node191 : node180;
							assign node180 = (inp[5]) ? node182 : 3'b100;
								assign node182 = (inp[11]) ? node184 : 3'b100;
									assign node184 = (inp[3]) ? node186 : 3'b100;
										assign node186 = (inp[7]) ? 3'b000 : node187;
											assign node187 = (inp[2]) ? 3'b000 : 3'b100;
							assign node191 = (inp[7]) ? node197 : node192;
								assign node192 = (inp[11]) ? node194 : 3'b101;
									assign node194 = (inp[2]) ? 3'b000 : 3'b100;
								assign node197 = (inp[11]) ? node203 : node198;
									assign node198 = (inp[10]) ? node200 : 3'b001;
										assign node200 = (inp[2]) ? 3'b000 : 3'b001;
									assign node203 = (inp[10]) ? 3'b000 : node204;
										assign node204 = (inp[2]) ? 3'b001 : 3'b000;
					assign node208 = (inp[4]) ? node210 : 3'b000;
						assign node210 = (inp[11]) ? node226 : node211;
							assign node211 = (inp[3]) ? node217 : node212;
								assign node212 = (inp[8]) ? node214 : 3'b100;
									assign node214 = (inp[2]) ? 3'b000 : 3'b101;
								assign node217 = (inp[2]) ? 3'b000 : node218;
									assign node218 = (inp[8]) ? 3'b101 : node219;
										assign node219 = (inp[7]) ? 3'b000 : node220;
											assign node220 = (inp[5]) ? 3'b100 : 3'b000;
							assign node226 = (inp[7]) ? 3'b000 : node227;
								assign node227 = (inp[8]) ? node229 : 3'b000;
									assign node229 = (inp[2]) ? 3'b000 : 3'b100;

endmodule