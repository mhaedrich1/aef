module dtc_split25_bm66 (
	input  wire [16-1:0] inp,
	output wire [4-1:0] outp
);

	wire [4-1:0] node1;
	wire [4-1:0] node2;
	wire [4-1:0] node3;
	wire [4-1:0] node4;
	wire [4-1:0] node6;
	wire [4-1:0] node7;
	wire [4-1:0] node9;
	wire [4-1:0] node11;
	wire [4-1:0] node13;
	wire [4-1:0] node14;
	wire [4-1:0] node15;
	wire [4-1:0] node17;
	wire [4-1:0] node21;
	wire [4-1:0] node24;
	wire [4-1:0] node25;
	wire [4-1:0] node26;
	wire [4-1:0] node28;
	wire [4-1:0] node29;
	wire [4-1:0] node31;
	wire [4-1:0] node33;
	wire [4-1:0] node35;
	wire [4-1:0] node39;
	wire [4-1:0] node40;
	wire [4-1:0] node41;
	wire [4-1:0] node42;
	wire [4-1:0] node44;
	wire [4-1:0] node51;
	wire [4-1:0] node52;
	wire [4-1:0] node54;
	wire [4-1:0] node56;
	wire [4-1:0] node58;
	wire [4-1:0] node60;
	wire [4-1:0] node63;
	wire [4-1:0] node64;
	wire [4-1:0] node66;
	wire [4-1:0] node68;
	wire [4-1:0] node70;
	wire [4-1:0] node71;
	wire [4-1:0] node73;
	wire [4-1:0] node77;
	wire [4-1:0] node78;
	wire [4-1:0] node79;
	wire [4-1:0] node80;
	wire [4-1:0] node82;
	wire [4-1:0] node84;
	wire [4-1:0] node90;
	wire [4-1:0] node91;
	wire [4-1:0] node92;
	wire [4-1:0] node93;
	wire [4-1:0] node95;
	wire [4-1:0] node97;
	wire [4-1:0] node99;
	wire [4-1:0] node100;
	wire [4-1:0] node104;
	wire [4-1:0] node105;
	wire [4-1:0] node107;
	wire [4-1:0] node108;
	wire [4-1:0] node110;
	wire [4-1:0] node111;
	wire [4-1:0] node113;
	wire [4-1:0] node119;
	wire [4-1:0] node120;
	wire [4-1:0] node122;
	wire [4-1:0] node124;
	wire [4-1:0] node125;
	wire [4-1:0] node127;
	wire [4-1:0] node129;
	wire [4-1:0] node133;
	wire [4-1:0] node134;
	wire [4-1:0] node135;
	wire [4-1:0] node137;
	wire [4-1:0] node139;
	wire [4-1:0] node141;
	wire [4-1:0] node146;
	wire [4-1:0] node147;
	wire [4-1:0] node148;
	wire [4-1:0] node150;
	wire [4-1:0] node152;
	wire [4-1:0] node153;
	wire [4-1:0] node154;
	wire [4-1:0] node156;
	wire [4-1:0] node157;
	wire [4-1:0] node163;
	wire [4-1:0] node164;
	wire [4-1:0] node165;
	wire [4-1:0] node166;
	wire [4-1:0] node168;
	wire [4-1:0] node170;
	wire [4-1:0] node176;
	wire [4-1:0] node177;
	wire [4-1:0] node179;
	wire [4-1:0] node182;
	wire [4-1:0] node184;
	wire [4-1:0] node186;
	wire [4-1:0] node187;
	wire [4-1:0] node189;
	wire [4-1:0] node193;
	wire [4-1:0] node194;
	wire [4-1:0] node195;
	wire [4-1:0] node196;
	wire [4-1:0] node197;
	wire [4-1:0] node198;
	wire [4-1:0] node200;
	wire [4-1:0] node201;
	wire [4-1:0] node203;
	wire [4-1:0] node205;
	wire [4-1:0] node209;
	wire [4-1:0] node211;
	wire [4-1:0] node213;
	wire [4-1:0] node216;
	wire [4-1:0] node217;
	wire [4-1:0] node218;
	wire [4-1:0] node220;
	wire [4-1:0] node221;
	wire [4-1:0] node227;
	wire [4-1:0] node228;
	wire [4-1:0] node230;
	wire [4-1:0] node232;
	wire [4-1:0] node234;
	wire [4-1:0] node236;
	wire [4-1:0] node238;
	wire [4-1:0] node241;
	wire [4-1:0] node243;
	wire [4-1:0] node246;
	wire [4-1:0] node247;
	wire [4-1:0] node248;
	wire [4-1:0] node249;
	wire [4-1:0] node251;
	wire [4-1:0] node252;
	wire [4-1:0] node254;
	wire [4-1:0] node256;
	wire [4-1:0] node258;
	wire [4-1:0] node261;
	wire [4-1:0] node265;
	wire [4-1:0] node266;
	wire [4-1:0] node268;
	wire [4-1:0] node272;
	wire [4-1:0] node273;
	wire [4-1:0] node274;
	wire [4-1:0] node275;
	wire [4-1:0] node276;
	wire [4-1:0] node278;
	wire [4-1:0] node280;
	wire [4-1:0] node285;
	wire [4-1:0] node287;
	wire [4-1:0] node288;
	wire [4-1:0] node289;
	wire [4-1:0] node294;
	wire [4-1:0] node296;
	wire [4-1:0] node297;
	wire [4-1:0] node301;
	wire [4-1:0] node302;
	wire [4-1:0] node303;
	wire [4-1:0] node304;
	wire [4-1:0] node305;
	wire [4-1:0] node306;
	wire [4-1:0] node309;
	wire [4-1:0] node311;
	wire [4-1:0] node312;
	wire [4-1:0] node314;
	wire [4-1:0] node316;
	wire [4-1:0] node319;
	wire [4-1:0] node322;
	wire [4-1:0] node323;
	wire [4-1:0] node324;
	wire [4-1:0] node325;
	wire [4-1:0] node326;
	wire [4-1:0] node327;
	wire [4-1:0] node330;
	wire [4-1:0] node333;
	wire [4-1:0] node334;
	wire [4-1:0] node335;
	wire [4-1:0] node340;
	wire [4-1:0] node341;
	wire [4-1:0] node342;
	wire [4-1:0] node345;
	wire [4-1:0] node346;
	wire [4-1:0] node351;
	wire [4-1:0] node352;
	wire [4-1:0] node353;
	wire [4-1:0] node354;
	wire [4-1:0] node357;
	wire [4-1:0] node360;
	wire [4-1:0] node362;
	wire [4-1:0] node365;
	wire [4-1:0] node366;
	wire [4-1:0] node367;
	wire [4-1:0] node370;
	wire [4-1:0] node373;
	wire [4-1:0] node374;
	wire [4-1:0] node377;
	wire [4-1:0] node380;
	wire [4-1:0] node381;
	wire [4-1:0] node382;
	wire [4-1:0] node385;
	wire [4-1:0] node388;
	wire [4-1:0] node389;
	wire [4-1:0] node390;
	wire [4-1:0] node394;
	wire [4-1:0] node397;
	wire [4-1:0] node398;
	wire [4-1:0] node400;
	wire [4-1:0] node401;
	wire [4-1:0] node402;
	wire [4-1:0] node404;
	wire [4-1:0] node406;
	wire [4-1:0] node411;
	wire [4-1:0] node413;
	wire [4-1:0] node414;
	wire [4-1:0] node416;
	wire [4-1:0] node418;
	wire [4-1:0] node422;
	wire [4-1:0] node423;
	wire [4-1:0] node424;
	wire [4-1:0] node426;
	wire [4-1:0] node428;
	wire [4-1:0] node431;
	wire [4-1:0] node433;
	wire [4-1:0] node435;
	wire [4-1:0] node436;
	wire [4-1:0] node440;
	wire [4-1:0] node442;
	wire [4-1:0] node444;
	wire [4-1:0] node446;
	wire [4-1:0] node449;
	wire [4-1:0] node450;
	wire [4-1:0] node451;
	wire [4-1:0] node452;
	wire [4-1:0] node453;
	wire [4-1:0] node454;
	wire [4-1:0] node455;
	wire [4-1:0] node456;
	wire [4-1:0] node458;
	wire [4-1:0] node464;
	wire [4-1:0] node466;
	wire [4-1:0] node470;
	wire [4-1:0] node472;
	wire [4-1:0] node474;
	wire [4-1:0] node475;
	wire [4-1:0] node477;
	wire [4-1:0] node479;
	wire [4-1:0] node480;
	wire [4-1:0] node484;
	wire [4-1:0] node485;
	wire [4-1:0] node488;
	wire [4-1:0] node490;
	wire [4-1:0] node493;
	wire [4-1:0] node494;
	wire [4-1:0] node495;
	wire [4-1:0] node496;
	wire [4-1:0] node497;
	wire [4-1:0] node499;
	wire [4-1:0] node501;
	wire [4-1:0] node506;
	wire [4-1:0] node509;
	wire [4-1:0] node511;
	wire [4-1:0] node513;
	wire [4-1:0] node515;
	wire [4-1:0] node516;
	wire [4-1:0] node518;
	wire [4-1:0] node522;
	wire [4-1:0] node523;
	wire [4-1:0] node524;
	wire [4-1:0] node525;
	wire [4-1:0] node526;
	wire [4-1:0] node527;
	wire [4-1:0] node528;
	wire [4-1:0] node530;
	wire [4-1:0] node532;
	wire [4-1:0] node533;
	wire [4-1:0] node534;
	wire [4-1:0] node535;
	wire [4-1:0] node542;
	wire [4-1:0] node543;
	wire [4-1:0] node545;
	wire [4-1:0] node546;
	wire [4-1:0] node548;
	wire [4-1:0] node550;
	wire [4-1:0] node554;
	wire [4-1:0] node556;
	wire [4-1:0] node558;
	wire [4-1:0] node561;
	wire [4-1:0] node562;
	wire [4-1:0] node564;
	wire [4-1:0] node565;
	wire [4-1:0] node566;
	wire [4-1:0] node567;
	wire [4-1:0] node569;
	wire [4-1:0] node571;
	wire [4-1:0] node574;
	wire [4-1:0] node579;
	wire [4-1:0] node581;
	wire [4-1:0] node582;
	wire [4-1:0] node584;
	wire [4-1:0] node586;
	wire [4-1:0] node587;
	wire [4-1:0] node589;
	wire [4-1:0] node594;
	wire [4-1:0] node595;
	wire [4-1:0] node596;
	wire [4-1:0] node597;
	wire [4-1:0] node599;
	wire [4-1:0] node601;
	wire [4-1:0] node604;
	wire [4-1:0] node606;
	wire [4-1:0] node608;
	wire [4-1:0] node610;
	wire [4-1:0] node612;
	wire [4-1:0] node614;
	wire [4-1:0] node618;
	wire [4-1:0] node619;
	wire [4-1:0] node620;
	wire [4-1:0] node622;
	wire [4-1:0] node624;
	wire [4-1:0] node626;
	wire [4-1:0] node628;
	wire [4-1:0] node630;
	wire [4-1:0] node632;
	wire [4-1:0] node635;
	wire [4-1:0] node636;
	wire [4-1:0] node637;
	wire [4-1:0] node638;
	wire [4-1:0] node639;
	wire [4-1:0] node641;
	wire [4-1:0] node649;
	wire [4-1:0] node650;
	wire [4-1:0] node651;
	wire [4-1:0] node652;
	wire [4-1:0] node653;
	wire [4-1:0] node654;
	wire [4-1:0] node655;
	wire [4-1:0] node659;
	wire [4-1:0] node661;
	wire [4-1:0] node663;
	wire [4-1:0] node665;
	wire [4-1:0] node667;
	wire [4-1:0] node670;
	wire [4-1:0] node671;
	wire [4-1:0] node672;
	wire [4-1:0] node673;
	wire [4-1:0] node675;
	wire [4-1:0] node680;
	wire [4-1:0] node682;
	wire [4-1:0] node685;
	wire [4-1:0] node687;
	wire [4-1:0] node690;
	wire [4-1:0] node691;
	wire [4-1:0] node693;
	wire [4-1:0] node694;
	wire [4-1:0] node695;
	wire [4-1:0] node700;
	wire [4-1:0] node701;
	wire [4-1:0] node703;
	wire [4-1:0] node704;
	wire [4-1:0] node706;
	wire [4-1:0] node708;
	wire [4-1:0] node713;
	wire [4-1:0] node714;
	wire [4-1:0] node715;
	wire [4-1:0] node717;
	wire [4-1:0] node718;
	wire [4-1:0] node720;
	wire [4-1:0] node722;
	wire [4-1:0] node724;
	wire [4-1:0] node726;
	wire [4-1:0] node730;
	wire [4-1:0] node731;
	wire [4-1:0] node733;
	wire [4-1:0] node735;
	wire [4-1:0] node736;
	wire [4-1:0] node738;
	wire [4-1:0] node739;
	wire [4-1:0] node745;
	wire [4-1:0] node746;
	wire [4-1:0] node747;
	wire [4-1:0] node748;
	wire [4-1:0] node750;
	wire [4-1:0] node752;
	wire [4-1:0] node753;
	wire [4-1:0] node755;
	wire [4-1:0] node760;
	wire [4-1:0] node762;
	wire [4-1:0] node764;
	wire [4-1:0] node767;
	wire [4-1:0] node769;
	wire [4-1:0] node770;
	wire [4-1:0] node772;
	wire [4-1:0] node773;
	wire [4-1:0] node774;
	wire [4-1:0] node776;
	wire [4-1:0] node778;
	wire [4-1:0] node784;
	wire [4-1:0] node785;
	wire [4-1:0] node786;
	wire [4-1:0] node787;
	wire [4-1:0] node788;
	wire [4-1:0] node790;
	wire [4-1:0] node792;
	wire [4-1:0] node794;
	wire [4-1:0] node796;
	wire [4-1:0] node799;
	wire [4-1:0] node800;
	wire [4-1:0] node801;
	wire [4-1:0] node803;
	wire [4-1:0] node806;
	wire [4-1:0] node807;
	wire [4-1:0] node808;
	wire [4-1:0] node809;
	wire [4-1:0] node811;
	wire [4-1:0] node813;
	wire [4-1:0] node819;
	wire [4-1:0] node821;
	wire [4-1:0] node823;
	wire [4-1:0] node826;
	wire [4-1:0] node827;
	wire [4-1:0] node829;
	wire [4-1:0] node831;
	wire [4-1:0] node833;
	wire [4-1:0] node834;
	wire [4-1:0] node836;
	wire [4-1:0] node840;
	wire [4-1:0] node841;
	wire [4-1:0] node842;
	wire [4-1:0] node843;
	wire [4-1:0] node845;
	wire [4-1:0] node847;
	wire [4-1:0] node852;
	wire [4-1:0] node854;
	wire [4-1:0] node855;
	wire [4-1:0] node857;
	wire [4-1:0] node858;
	wire [4-1:0] node859;
	wire [4-1:0] node861;
	wire [4-1:0] node867;
	wire [4-1:0] node868;
	wire [4-1:0] node869;
	wire [4-1:0] node870;
	wire [4-1:0] node872;
	wire [4-1:0] node874;
	wire [4-1:0] node875;
	wire [4-1:0] node879;
	wire [4-1:0] node880;
	wire [4-1:0] node882;
	wire [4-1:0] node884;
	wire [4-1:0] node886;
	wire [4-1:0] node890;
	wire [4-1:0] node891;
	wire [4-1:0] node892;
	wire [4-1:0] node894;
	wire [4-1:0] node897;
	wire [4-1:0] node899;
	wire [4-1:0] node902;
	wire [4-1:0] node903;
	wire [4-1:0] node904;
	wire [4-1:0] node906;
	wire [4-1:0] node908;
	wire [4-1:0] node910;
	wire [4-1:0] node914;
	wire [4-1:0] node915;
	wire [4-1:0] node916;
	wire [4-1:0] node918;
	wire [4-1:0] node923;
	wire [4-1:0] node924;
	wire [4-1:0] node925;
	wire [4-1:0] node928;
	wire [4-1:0] node929;
	wire [4-1:0] node930;
	wire [4-1:0] node931;
	wire [4-1:0] node933;
	wire [4-1:0] node935;
	wire [4-1:0] node941;
	wire [4-1:0] node942;
	wire [4-1:0] node944;
	wire [4-1:0] node946;
	wire [4-1:0] node948;
	wire [4-1:0] node950;
	wire [4-1:0] node953;
	wire [4-1:0] node954;
	wire [4-1:0] node955;
	wire [4-1:0] node957;
	wire [4-1:0] node959;
	wire [4-1:0] node961;
	wire [4-1:0] node963;
	wire [4-1:0] node967;
	wire [4-1:0] node970;
	wire [4-1:0] node971;
	wire [4-1:0] node972;
	wire [4-1:0] node973;
	wire [4-1:0] node974;
	wire [4-1:0] node975;
	wire [4-1:0] node976;
	wire [4-1:0] node978;
	wire [4-1:0] node980;
	wire [4-1:0] node982;
	wire [4-1:0] node985;
	wire [4-1:0] node986;
	wire [4-1:0] node987;
	wire [4-1:0] node989;
	wire [4-1:0] node991;
	wire [4-1:0] node997;
	wire [4-1:0] node998;
	wire [4-1:0] node1000;
	wire [4-1:0] node1002;
	wire [4-1:0] node1004;
	wire [4-1:0] node1007;
	wire [4-1:0] node1008;
	wire [4-1:0] node1012;
	wire [4-1:0] node1013;
	wire [4-1:0] node1015;
	wire [4-1:0] node1016;
	wire [4-1:0] node1017;
	wire [4-1:0] node1022;
	wire [4-1:0] node1023;
	wire [4-1:0] node1025;
	wire [4-1:0] node1026;
	wire [4-1:0] node1027;
	wire [4-1:0] node1029;
	wire [4-1:0] node1034;
	wire [4-1:0] node1036;
	wire [4-1:0] node1039;
	wire [4-1:0] node1040;
	wire [4-1:0] node1041;
	wire [4-1:0] node1042;
	wire [4-1:0] node1043;
	wire [4-1:0] node1045;
	wire [4-1:0] node1047;
	wire [4-1:0] node1051;
	wire [4-1:0] node1053;
	wire [4-1:0] node1054;
	wire [4-1:0] node1056;
	wire [4-1:0] node1058;
	wire [4-1:0] node1059;
	wire [4-1:0] node1063;
	wire [4-1:0] node1066;
	wire [4-1:0] node1067;
	wire [4-1:0] node1069;
	wire [4-1:0] node1070;
	wire [4-1:0] node1072;
	wire [4-1:0] node1074;
	wire [4-1:0] node1075;
	wire [4-1:0] node1080;
	wire [4-1:0] node1082;
	wire [4-1:0] node1084;
	wire [4-1:0] node1086;
	wire [4-1:0] node1089;
	wire [4-1:0] node1090;
	wire [4-1:0] node1092;
	wire [4-1:0] node1094;
	wire [4-1:0] node1096;
	wire [4-1:0] node1098;
	wire [4-1:0] node1101;
	wire [4-1:0] node1104;
	wire [4-1:0] node1105;
	wire [4-1:0] node1106;
	wire [4-1:0] node1107;
	wire [4-1:0] node1109;
	wire [4-1:0] node1111;
	wire [4-1:0] node1113;
	wire [4-1:0] node1116;
	wire [4-1:0] node1118;
	wire [4-1:0] node1120;
	wire [4-1:0] node1121;
	wire [4-1:0] node1123;
	wire [4-1:0] node1127;
	wire [4-1:0] node1128;
	wire [4-1:0] node1129;
	wire [4-1:0] node1130;
	wire [4-1:0] node1131;
	wire [4-1:0] node1133;
	wire [4-1:0] node1135;
	wire [4-1:0] node1138;
	wire [4-1:0] node1139;
	wire [4-1:0] node1143;
	wire [4-1:0] node1144;
	wire [4-1:0] node1145;
	wire [4-1:0] node1146;
	wire [4-1:0] node1147;
	wire [4-1:0] node1151;
	wire [4-1:0] node1155;
	wire [4-1:0] node1156;
	wire [4-1:0] node1157;
	wire [4-1:0] node1161;
	wire [4-1:0] node1164;
	wire [4-1:0] node1165;
	wire [4-1:0] node1168;
	wire [4-1:0] node1171;
	wire [4-1:0] node1172;
	wire [4-1:0] node1174;
	wire [4-1:0] node1176;
	wire [4-1:0] node1178;
	wire [4-1:0] node1179;
	wire [4-1:0] node1183;
	wire [4-1:0] node1185;
	wire [4-1:0] node1186;
	wire [4-1:0] node1188;
	wire [4-1:0] node1192;
	wire [4-1:0] node1193;
	wire [4-1:0] node1194;
	wire [4-1:0] node1195;
	wire [4-1:0] node1196;
	wire [4-1:0] node1197;
	wire [4-1:0] node1199;
	wire [4-1:0] node1201;
	wire [4-1:0] node1205;
	wire [4-1:0] node1208;
	wire [4-1:0] node1209;
	wire [4-1:0] node1210;
	wire [4-1:0] node1211;
	wire [4-1:0] node1213;
	wire [4-1:0] node1219;
	wire [4-1:0] node1220;
	wire [4-1:0] node1221;
	wire [4-1:0] node1223;
	wire [4-1:0] node1225;
	wire [4-1:0] node1229;
	wire [4-1:0] node1230;
	wire [4-1:0] node1232;
	wire [4-1:0] node1234;
	wire [4-1:0] node1236;
	wire [4-1:0] node1239;
	wire [4-1:0] node1242;
	wire [4-1:0] node1243;
	wire [4-1:0] node1244;
	wire [4-1:0] node1246;
	wire [4-1:0] node1247;
	wire [4-1:0] node1249;
	wire [4-1:0] node1251;
	wire [4-1:0] node1254;
	wire [4-1:0] node1255;
	wire [4-1:0] node1257;
	wire [4-1:0] node1261;
	wire [4-1:0] node1263;
	wire [4-1:0] node1264;
	wire [4-1:0] node1266;
	wire [4-1:0] node1270;
	wire [4-1:0] node1271;
	wire [4-1:0] node1272;
	wire [4-1:0] node1273;
	wire [4-1:0] node1276;
	wire [4-1:0] node1278;
	wire [4-1:0] node1280;
	wire [4-1:0] node1283;
	wire [4-1:0] node1284;
	wire [4-1:0] node1286;
	wire [4-1:0] node1290;
	wire [4-1:0] node1291;
	wire [4-1:0] node1292;
	wire [4-1:0] node1293;
	wire [4-1:0] node1295;
	wire [4-1:0] node1297;
	wire [4-1:0] node1301;
	wire [4-1:0] node1302;
	wire [4-1:0] node1304;
	wire [4-1:0] node1308;
	wire [4-1:0] node1309;
	wire [4-1:0] node1311;
	wire [4-1:0] node1314;
	wire [4-1:0] node1315;

	assign outp = (inp[10]) ? node522 : node1;
		assign node1 = (inp[5]) ? node193 : node2;
			assign node2 = (inp[4]) ? node90 : node3;
				assign node3 = (inp[14]) ? node51 : node4;
					assign node4 = (inp[13]) ? node6 : 4'b1111;
						assign node6 = (inp[12]) ? node24 : node7;
							assign node7 = (inp[9]) ? node9 : 4'b1111;
								assign node9 = (inp[2]) ? node11 : 4'b1111;
									assign node11 = (inp[8]) ? node13 : 4'b1111;
										assign node13 = (inp[6]) ? node21 : node14;
											assign node14 = (inp[3]) ? 4'b1111 : node15;
												assign node15 = (inp[0]) ? node17 : 4'b1111;
													assign node17 = (inp[1]) ? 4'b1101 : 4'b1111;
											assign node21 = (inp[7]) ? 4'b1101 : 4'b1111;
							assign node24 = (inp[2]) ? 4'b1101 : node25;
								assign node25 = (inp[6]) ? node39 : node26;
									assign node26 = (inp[9]) ? node28 : 4'b1111;
										assign node28 = (inp[8]) ? 4'b1101 : node29;
											assign node29 = (inp[7]) ? node31 : 4'b1111;
												assign node31 = (inp[0]) ? node33 : 4'b1111;
													assign node33 = (inp[15]) ? node35 : 4'b1111;
														assign node35 = (inp[11]) ? 4'b1101 : 4'b1111;
									assign node39 = (inp[9]) ? 4'b1101 : node40;
										assign node40 = (inp[8]) ? 4'b1101 : node41;
											assign node41 = (inp[7]) ? 4'b1101 : node42;
												assign node42 = (inp[11]) ? node44 : 4'b1111;
													assign node44 = (inp[1]) ? 4'b1101 : 4'b1111;
					assign node51 = (inp[13]) ? node63 : node52;
						assign node52 = (inp[6]) ? node54 : 4'b1101;
							assign node54 = (inp[2]) ? node56 : 4'b1101;
								assign node56 = (inp[12]) ? node58 : 4'b1101;
									assign node58 = (inp[9]) ? node60 : 4'b1101;
										assign node60 = (inp[8]) ? 4'b1011 : 4'b1101;
						assign node63 = (inp[12]) ? node77 : node64;
							assign node64 = (inp[2]) ? node66 : 4'b1101;
								assign node66 = (inp[8]) ? node68 : 4'b1101;
									assign node68 = (inp[9]) ? node70 : 4'b1101;
										assign node70 = (inp[6]) ? 4'b1011 : node71;
											assign node71 = (inp[7]) ? node73 : 4'b1101;
												assign node73 = (inp[15]) ? 4'b1111 : 4'b1101;
							assign node77 = (inp[6]) ? 4'b1011 : node78;
								assign node78 = (inp[9]) ? 4'b1111 : node79;
									assign node79 = (inp[2]) ? 4'b1111 : node80;
										assign node80 = (inp[7]) ? node82 : 4'b1101;
											assign node82 = (inp[15]) ? node84 : 4'b1101;
												assign node84 = (inp[1]) ? 4'b1111 : 4'b1101;
				assign node90 = (inp[6]) ? node146 : node91;
					assign node91 = (inp[14]) ? node119 : node92;
						assign node92 = (inp[12]) ? node104 : node93;
							assign node93 = (inp[2]) ? node95 : 4'b1011;
								assign node95 = (inp[9]) ? node97 : 4'b1011;
									assign node97 = (inp[13]) ? node99 : 4'b1011;
										assign node99 = (inp[7]) ? 4'b1001 : node100;
											assign node100 = (inp[8]) ? 4'b1001 : 4'b1011;
							assign node104 = (inp[13]) ? 4'b1001 : node105;
								assign node105 = (inp[2]) ? node107 : 4'b1011;
									assign node107 = (inp[9]) ? 4'b1001 : node108;
										assign node108 = (inp[8]) ? node110 : 4'b1011;
											assign node110 = (inp[7]) ? 4'b1001 : node111;
												assign node111 = (inp[1]) ? node113 : 4'b1011;
													assign node113 = (inp[0]) ? 4'b1011 : 4'b1001;
						assign node119 = (inp[12]) ? node133 : node120;
							assign node120 = (inp[13]) ? node122 : 4'b1001;
								assign node122 = (inp[2]) ? node124 : 4'b1001;
									assign node124 = (inp[9]) ? 4'b1011 : node125;
										assign node125 = (inp[8]) ? node127 : 4'b1001;
											assign node127 = (inp[7]) ? node129 : 4'b1001;
												assign node129 = (inp[15]) ? 4'b1011 : 4'b1001;
							assign node133 = (inp[13]) ? 4'b1011 : node134;
								assign node134 = (inp[2]) ? 4'b1011 : node135;
									assign node135 = (inp[8]) ? node137 : 4'b1001;
										assign node137 = (inp[7]) ? node139 : 4'b1001;
											assign node139 = (inp[9]) ? node141 : 4'b1001;
												assign node141 = (inp[15]) ? 4'b1011 : 4'b1001;
					assign node146 = (inp[14]) ? node176 : node147;
						assign node147 = (inp[12]) ? node163 : node148;
							assign node148 = (inp[2]) ? node150 : 4'b1011;
								assign node150 = (inp[13]) ? node152 : 4'b1011;
									assign node152 = (inp[9]) ? 4'b1001 : node153;
										assign node153 = (inp[8]) ? 4'b1001 : node154;
											assign node154 = (inp[11]) ? node156 : 4'b1011;
												assign node156 = (inp[0]) ? 4'b1011 : node157;
													assign node157 = (inp[15]) ? 4'b1001 : 4'b1011;
							assign node163 = (inp[13]) ? 4'b1001 : node164;
								assign node164 = (inp[9]) ? 4'b1001 : node165;
									assign node165 = (inp[2]) ? 4'b1001 : node166;
										assign node166 = (inp[7]) ? node168 : 4'b1011;
											assign node168 = (inp[15]) ? node170 : 4'b1011;
												assign node170 = (inp[11]) ? 4'b1001 : 4'b1011;
						assign node176 = (inp[12]) ? node182 : node177;
							assign node177 = (inp[13]) ? node179 : 4'b1001;
								assign node179 = (inp[2]) ? 4'b1111 : 4'b1001;
							assign node182 = (inp[13]) ? node184 : 4'b1110;
								assign node184 = (inp[2]) ? node186 : 4'b1110;
									assign node186 = (inp[9]) ? 4'b1100 : node187;
										assign node187 = (inp[1]) ? node189 : 4'b1110;
											assign node189 = (inp[0]) ? 4'b1100 : 4'b1110;
			assign node193 = (inp[12]) ? node301 : node194;
				assign node194 = (inp[6]) ? node246 : node195;
					assign node195 = (inp[13]) ? node227 : node196;
						assign node196 = (inp[14]) ? node216 : node197;
							assign node197 = (inp[4]) ? node209 : node198;
								assign node198 = (inp[2]) ? node200 : 4'b1001;
									assign node200 = (inp[9]) ? 4'b1011 : node201;
										assign node201 = (inp[8]) ? node203 : 4'b1001;
											assign node203 = (inp[15]) ? node205 : 4'b1001;
												assign node205 = (inp[7]) ? 4'b1011 : 4'b1001;
								assign node209 = (inp[8]) ? node211 : 4'b1101;
									assign node211 = (inp[9]) ? node213 : 4'b1101;
										assign node213 = (inp[2]) ? 4'b1011 : 4'b1101;
							assign node216 = (inp[2]) ? 4'b1001 : node217;
								assign node217 = (inp[9]) ? 4'b1001 : node218;
									assign node218 = (inp[8]) ? node220 : 4'b1011;
										assign node220 = (inp[7]) ? 4'b1001 : node221;
											assign node221 = (inp[4]) ? 4'b1011 : 4'b1001;
						assign node227 = (inp[2]) ? node241 : node228;
							assign node228 = (inp[14]) ? node230 : 4'b1011;
								assign node230 = (inp[0]) ? node232 : 4'b1001;
									assign node232 = (inp[8]) ? node234 : 4'b1001;
										assign node234 = (inp[7]) ? node236 : 4'b1001;
											assign node236 = (inp[4]) ? node238 : 4'b1001;
												assign node238 = (inp[9]) ? 4'b1011 : 4'b1001;
							assign node241 = (inp[14]) ? node243 : 4'b1011;
								assign node243 = (inp[4]) ? 4'b1011 : 4'b1111;
					assign node246 = (inp[14]) ? node272 : node247;
						assign node247 = (inp[4]) ? node265 : node248;
							assign node248 = (inp[13]) ? 4'b1101 : node249;
								assign node249 = (inp[2]) ? node251 : 4'b1111;
									assign node251 = (inp[8]) ? node261 : node252;
										assign node252 = (inp[1]) ? node254 : 4'b1111;
											assign node254 = (inp[15]) ? node256 : 4'b1111;
												assign node256 = (inp[9]) ? node258 : 4'b1111;
													assign node258 = (inp[0]) ? 4'b1111 : 4'b1101;
										assign node261 = (inp[9]) ? 4'b1101 : 4'b1111;
							assign node265 = (inp[13]) ? 4'b1001 : node266;
								assign node266 = (inp[2]) ? node268 : 4'b1011;
									assign node268 = (inp[9]) ? 4'b1001 : 4'b1011;
						assign node272 = (inp[4]) ? node294 : node273;
							assign node273 = (inp[13]) ? node285 : node274;
								assign node274 = (inp[2]) ? 4'b1111 : node275;
									assign node275 = (inp[9]) ? 4'b1111 : node276;
										assign node276 = (inp[8]) ? node278 : 4'b1101;
											assign node278 = (inp[7]) ? node280 : 4'b1101;
												assign node280 = (inp[15]) ? 4'b1111 : 4'b1101;
								assign node285 = (inp[2]) ? node287 : 4'b1111;
									assign node287 = (inp[8]) ? 4'b1101 : node288;
										assign node288 = (inp[9]) ? 4'b1101 : node289;
											assign node289 = (inp[7]) ? 4'b1101 : 4'b1111;
							assign node294 = (inp[13]) ? node296 : 4'b1110;
								assign node296 = (inp[2]) ? 4'b1100 : node297;
									assign node297 = (inp[9]) ? 4'b1100 : 4'b1110;
				assign node301 = (inp[6]) ? node449 : node302;
					assign node302 = (inp[14]) ? node422 : node303;
						assign node303 = (inp[4]) ? node397 : node304;
							assign node304 = (inp[9]) ? node322 : node305;
								assign node305 = (inp[2]) ? node309 : node306;
									assign node306 = (inp[13]) ? 4'b1110 : 4'b1100;
									assign node309 = (inp[13]) ? node311 : 4'b1110;
										assign node311 = (inp[7]) ? node319 : node312;
											assign node312 = (inp[15]) ? node314 : 4'b1110;
												assign node314 = (inp[11]) ? node316 : 4'b1110;
													assign node316 = (inp[8]) ? 4'b1100 : 4'b1110;
											assign node319 = (inp[8]) ? 4'b1100 : 4'b1110;
								assign node322 = (inp[8]) ? node380 : node323;
									assign node323 = (inp[3]) ? node351 : node324;
										assign node324 = (inp[15]) ? node340 : node325;
											assign node325 = (inp[11]) ? node333 : node326;
												assign node326 = (inp[2]) ? node330 : node327;
													assign node327 = (inp[13]) ? 4'b1110 : 4'b1100;
													assign node330 = (inp[13]) ? 4'b1100 : 4'b1110;
												assign node333 = (inp[7]) ? 4'b1100 : node334;
													assign node334 = (inp[13]) ? 4'b1100 : node335;
														assign node335 = (inp[2]) ? 4'b1110 : 4'b1100;
											assign node340 = (inp[0]) ? 4'b1100 : node341;
												assign node341 = (inp[1]) ? node345 : node342;
													assign node342 = (inp[11]) ? 4'b1100 : 4'b1110;
													assign node345 = (inp[13]) ? 4'b1100 : node346;
														assign node346 = (inp[2]) ? 4'b1110 : 4'b1100;
										assign node351 = (inp[0]) ? node365 : node352;
											assign node352 = (inp[11]) ? node360 : node353;
												assign node353 = (inp[2]) ? node357 : node354;
													assign node354 = (inp[13]) ? 4'b1110 : 4'b1100;
													assign node357 = (inp[13]) ? 4'b1100 : 4'b1110;
												assign node360 = (inp[13]) ? node362 : 4'b1100;
													assign node362 = (inp[2]) ? 4'b1100 : 4'b1110;
											assign node365 = (inp[1]) ? node373 : node366;
												assign node366 = (inp[15]) ? node370 : node367;
													assign node367 = (inp[2]) ? 4'b1110 : 4'b1100;
													assign node370 = (inp[7]) ? 4'b1110 : 4'b1100;
												assign node373 = (inp[2]) ? node377 : node374;
													assign node374 = (inp[13]) ? 4'b1110 : 4'b1100;
													assign node377 = (inp[7]) ? 4'b1110 : 4'b1100;
									assign node380 = (inp[7]) ? node388 : node381;
										assign node381 = (inp[13]) ? node385 : node382;
											assign node382 = (inp[2]) ? 4'b1110 : 4'b1100;
											assign node385 = (inp[2]) ? 4'b1100 : 4'b1110;
										assign node388 = (inp[13]) ? node394 : node389;
											assign node389 = (inp[15]) ? 4'b1110 : node390;
												assign node390 = (inp[2]) ? 4'b1110 : 4'b1100;
											assign node394 = (inp[2]) ? 4'b1100 : 4'b1110;
							assign node397 = (inp[13]) ? node411 : node398;
								assign node398 = (inp[2]) ? node400 : 4'b1110;
									assign node400 = (inp[9]) ? 4'b1100 : node401;
										assign node401 = (inp[8]) ? 4'b1100 : node402;
											assign node402 = (inp[3]) ? node404 : 4'b1110;
												assign node404 = (inp[15]) ? node406 : 4'b1110;
													assign node406 = (inp[11]) ? 4'b1100 : 4'b1110;
								assign node411 = (inp[2]) ? node413 : 4'b1100;
									assign node413 = (inp[9]) ? 4'b1110 : node414;
										assign node414 = (inp[8]) ? node416 : 4'b1100;
											assign node416 = (inp[15]) ? node418 : 4'b1100;
												assign node418 = (inp[7]) ? 4'b1110 : 4'b1100;
						assign node422 = (inp[13]) ? node440 : node423;
							assign node423 = (inp[4]) ? node431 : node424;
								assign node424 = (inp[8]) ? node426 : 4'b1100;
									assign node426 = (inp[9]) ? node428 : 4'b1100;
										assign node428 = (inp[2]) ? 4'b1010 : 4'b1100;
								assign node431 = (inp[9]) ? node433 : 4'b1110;
									assign node433 = (inp[2]) ? node435 : 4'b1110;
										assign node435 = (inp[8]) ? 4'b1100 : node436;
											assign node436 = (inp[7]) ? 4'b1100 : 4'b1110;
							assign node440 = (inp[4]) ? node442 : 4'b1010;
								assign node442 = (inp[9]) ? node444 : 4'b1100;
									assign node444 = (inp[8]) ? node446 : 4'b1100;
										assign node446 = (inp[2]) ? 4'b1010 : 4'b1100;
					assign node449 = (inp[13]) ? node493 : node450;
						assign node450 = (inp[4]) ? node470 : node451;
							assign node451 = (inp[2]) ? 4'b1000 : node452;
								assign node452 = (inp[14]) ? node464 : node453;
									assign node453 = (inp[7]) ? 4'b1000 : node454;
										assign node454 = (inp[8]) ? 4'b1000 : node455;
											assign node455 = (inp[9]) ? 4'b1000 : node456;
												assign node456 = (inp[1]) ? node458 : 4'b1010;
													assign node458 = (inp[11]) ? 4'b1000 : 4'b1010;
									assign node464 = (inp[8]) ? node466 : 4'b1010;
										assign node466 = (inp[9]) ? 4'b1000 : 4'b1010;
							assign node470 = (inp[2]) ? node472 : 4'b1010;
								assign node472 = (inp[8]) ? node474 : 4'b1010;
									assign node474 = (inp[7]) ? node484 : node475;
										assign node475 = (inp[15]) ? node477 : 4'b1010;
											assign node477 = (inp[11]) ? node479 : 4'b1010;
												assign node479 = (inp[14]) ? 4'b1010 : node480;
													assign node480 = (inp[0]) ? 4'b1000 : 4'b1010;
										assign node484 = (inp[14]) ? node488 : node485;
											assign node485 = (inp[9]) ? 4'b1000 : 4'b1010;
											assign node488 = (inp[1]) ? node490 : 4'b1010;
												assign node490 = (inp[9]) ? 4'b1000 : 4'b1010;
						assign node493 = (inp[4]) ? node509 : node494;
							assign node494 = (inp[2]) ? node506 : node495;
								assign node495 = (inp[14]) ? 4'b1000 : node496;
									assign node496 = (inp[9]) ? 4'b1010 : node497;
										assign node497 = (inp[7]) ? node499 : 4'b1000;
											assign node499 = (inp[8]) ? node501 : 4'b1000;
												assign node501 = (inp[15]) ? 4'b1010 : 4'b1000;
								assign node506 = (inp[14]) ? 4'b1110 : 4'b1010;
							assign node509 = (inp[15]) ? node511 : 4'b1000;
								assign node511 = (inp[8]) ? node513 : 4'b1000;
									assign node513 = (inp[9]) ? node515 : 4'b1000;
										assign node515 = (inp[14]) ? 4'b1000 : node516;
											assign node516 = (inp[2]) ? node518 : 4'b1000;
												assign node518 = (inp[7]) ? 4'b1010 : 4'b1000;
		assign node522 = (inp[5]) ? node784 : node523;
			assign node523 = (inp[4]) ? node649 : node524;
				assign node524 = (inp[6]) ? node594 : node525;
					assign node525 = (inp[14]) ? node561 : node526;
						assign node526 = (inp[13]) ? node542 : node527;
							assign node527 = (inp[2]) ? 4'b1100 : node528;
								assign node528 = (inp[12]) ? node530 : 4'b1100;
									assign node530 = (inp[9]) ? node532 : 4'b1110;
										assign node532 = (inp[8]) ? 4'b1100 : node533;
											assign node533 = (inp[7]) ? 4'b1100 : node534;
												assign node534 = (inp[0]) ? 4'b1110 : node535;
													assign node535 = (inp[11]) ? 4'b1100 : 4'b1110;
							assign node542 = (inp[2]) ? node554 : node543;
								assign node543 = (inp[8]) ? node545 : 4'b1100;
									assign node545 = (inp[12]) ? 4'b1100 : node546;
										assign node546 = (inp[7]) ? node548 : 4'b1100;
											assign node548 = (inp[15]) ? node550 : 4'b1100;
												assign node550 = (inp[9]) ? 4'b1110 : 4'b1100;
								assign node554 = (inp[12]) ? node556 : 4'b1110;
									assign node556 = (inp[8]) ? node558 : 4'b1100;
										assign node558 = (inp[9]) ? 4'b1010 : 4'b1100;
						assign node561 = (inp[12]) ? node579 : node562;
							assign node562 = (inp[13]) ? node564 : 4'b1110;
								assign node564 = (inp[2]) ? 4'b1100 : node565;
									assign node565 = (inp[9]) ? 4'b1100 : node566;
										assign node566 = (inp[7]) ? node574 : node567;
											assign node567 = (inp[3]) ? node569 : 4'b1110;
												assign node569 = (inp[1]) ? node571 : 4'b1110;
													assign node571 = (inp[0]) ? 4'b1110 : 4'b1100;
											assign node574 = (inp[8]) ? 4'b1100 : 4'b1110;
							assign node579 = (inp[13]) ? node581 : 4'b1010;
								assign node581 = (inp[2]) ? 4'b1000 : node582;
									assign node582 = (inp[8]) ? node584 : 4'b1010;
										assign node584 = (inp[9]) ? node586 : 4'b1010;
											assign node586 = (inp[7]) ? 4'b1000 : node587;
												assign node587 = (inp[11]) ? node589 : 4'b1010;
													assign node589 = (inp[1]) ? 4'b1000 : 4'b1010;
					assign node594 = (inp[14]) ? node618 : node595;
						assign node595 = (inp[13]) ? 4'b1010 : node596;
							assign node596 = (inp[12]) ? node604 : node597;
								assign node597 = (inp[2]) ? node599 : 4'b1100;
									assign node599 = (inp[8]) ? node601 : 4'b1100;
										assign node601 = (inp[9]) ? 4'b1010 : 4'b1100;
								assign node604 = (inp[9]) ? node606 : 4'b1000;
									assign node606 = (inp[1]) ? node608 : 4'b1000;
										assign node608 = (inp[7]) ? node610 : 4'b1000;
											assign node610 = (inp[8]) ? node612 : 4'b1000;
												assign node612 = (inp[15]) ? node614 : 4'b1000;
													assign node614 = (inp[2]) ? 4'b1010 : 4'b1000;
						assign node618 = (inp[13]) ? 4'b1000 : node619;
							assign node619 = (inp[2]) ? node635 : node620;
								assign node620 = (inp[12]) ? node622 : 4'b1010;
									assign node622 = (inp[1]) ? node624 : 4'b1010;
										assign node624 = (inp[8]) ? node626 : 4'b1010;
											assign node626 = (inp[15]) ? node628 : 4'b1010;
												assign node628 = (inp[7]) ? node630 : 4'b1010;
													assign node630 = (inp[11]) ? node632 : 4'b1010;
														assign node632 = (inp[9]) ? 4'b1000 : 4'b1010;
								assign node635 = (inp[8]) ? 4'b1000 : node636;
									assign node636 = (inp[12]) ? 4'b1000 : node637;
										assign node637 = (inp[9]) ? 4'b1000 : node638;
											assign node638 = (inp[7]) ? 4'b1000 : node639;
												assign node639 = (inp[11]) ? node641 : 4'b1010;
													assign node641 = (inp[1]) ? 4'b1000 : 4'b1010;
				assign node649 = (inp[12]) ? node713 : node650;
					assign node650 = (inp[6]) ? node690 : node651;
						assign node651 = (inp[14]) ? node685 : node652;
							assign node652 = (inp[8]) ? node670 : node653;
								assign node653 = (inp[2]) ? node659 : node654;
									assign node654 = (inp[9]) ? 4'b1010 : node655;
										assign node655 = (inp[13]) ? 4'b1010 : 4'b1000;
									assign node659 = (inp[7]) ? node661 : 4'b1010;
										assign node661 = (inp[11]) ? node663 : 4'b1010;
											assign node663 = (inp[9]) ? node665 : 4'b1010;
												assign node665 = (inp[1]) ? node667 : 4'b1010;
													assign node667 = (inp[13]) ? 4'b1000 : 4'b1010;
								assign node670 = (inp[13]) ? node680 : node671;
									assign node671 = (inp[2]) ? 4'b1010 : node672;
										assign node672 = (inp[9]) ? 4'b1010 : node673;
											assign node673 = (inp[7]) ? node675 : 4'b1000;
												assign node675 = (inp[15]) ? 4'b1010 : 4'b1000;
									assign node680 = (inp[2]) ? node682 : 4'b1010;
										assign node682 = (inp[9]) ? 4'b1000 : 4'b1010;
							assign node685 = (inp[2]) ? node687 : 4'b1000;
								assign node687 = (inp[13]) ? 4'b1110 : 4'b1000;
						assign node690 = (inp[14]) ? node700 : node691;
							assign node691 = (inp[13]) ? node693 : 4'b1110;
								assign node693 = (inp[8]) ? 4'b1100 : node694;
									assign node694 = (inp[2]) ? 4'b1100 : node695;
										assign node695 = (inp[9]) ? 4'b1100 : 4'b1110;
							assign node700 = (inp[13]) ? 4'b1110 : node701;
								assign node701 = (inp[2]) ? node703 : 4'b1100;
									assign node703 = (inp[9]) ? 4'b1110 : node704;
										assign node704 = (inp[1]) ? node706 : 4'b1100;
											assign node706 = (inp[7]) ? node708 : 4'b1100;
												assign node708 = (inp[15]) ? 4'b1110 : 4'b1100;
					assign node713 = (inp[6]) ? node745 : node714;
						assign node714 = (inp[14]) ? node730 : node715;
							assign node715 = (inp[13]) ? node717 : 4'b1111;
								assign node717 = (inp[2]) ? 4'b1101 : node718;
									assign node718 = (inp[0]) ? node720 : 4'b1111;
										assign node720 = (inp[11]) ? node722 : 4'b1111;
											assign node722 = (inp[15]) ? node724 : 4'b1111;
												assign node724 = (inp[3]) ? node726 : 4'b1111;
													assign node726 = (inp[9]) ? 4'b1101 : 4'b1111;
							assign node730 = (inp[13]) ? 4'b1111 : node731;
								assign node731 = (inp[8]) ? node733 : 4'b1101;
									assign node733 = (inp[15]) ? node735 : 4'b1101;
										assign node735 = (inp[0]) ? 4'b1101 : node736;
											assign node736 = (inp[1]) ? node738 : 4'b1101;
												assign node738 = (inp[3]) ? 4'b1101 : node739;
													assign node739 = (inp[9]) ? 4'b1111 : 4'b1101;
						assign node745 = (inp[14]) ? node767 : node746;
							assign node746 = (inp[2]) ? node760 : node747;
								assign node747 = (inp[13]) ? 4'b1101 : node748;
									assign node748 = (inp[8]) ? node750 : 4'b1111;
										assign node750 = (inp[9]) ? node752 : 4'b1111;
											assign node752 = (inp[7]) ? 4'b1101 : node753;
												assign node753 = (inp[11]) ? node755 : 4'b1111;
													assign node755 = (inp[15]) ? 4'b1101 : 4'b1111;
								assign node760 = (inp[8]) ? node762 : 4'b1101;
									assign node762 = (inp[13]) ? node764 : 4'b1101;
										assign node764 = (inp[9]) ? 4'b1011 : 4'b1101;
							assign node767 = (inp[13]) ? node769 : 4'b1011;
								assign node769 = (inp[2]) ? 4'b1001 : node770;
									assign node770 = (inp[9]) ? node772 : 4'b1011;
										assign node772 = (inp[8]) ? 4'b1001 : node773;
											assign node773 = (inp[7]) ? 4'b1001 : node774;
												assign node774 = (inp[15]) ? node776 : 4'b1011;
													assign node776 = (inp[1]) ? node778 : 4'b1011;
														assign node778 = (inp[11]) ? 4'b1001 : 4'b1011;
			assign node784 = (inp[12]) ? node970 : node785;
				assign node785 = (inp[6]) ? node867 : node786;
					assign node786 = (inp[13]) ? node826 : node787;
						assign node787 = (inp[4]) ? node799 : node788;
							assign node788 = (inp[8]) ? node790 : 4'b0111;
								assign node790 = (inp[14]) ? node792 : 4'b0111;
									assign node792 = (inp[9]) ? node794 : 4'b0111;
										assign node794 = (inp[2]) ? node796 : 4'b0111;
											assign node796 = (inp[7]) ? 4'b0101 : 4'b0111;
							assign node799 = (inp[2]) ? node819 : node800;
								assign node800 = (inp[14]) ? node806 : node801;
									assign node801 = (inp[9]) ? node803 : 4'b0111;
										assign node803 = (inp[8]) ? 4'b0101 : 4'b0111;
									assign node806 = (inp[7]) ? 4'b0101 : node807;
										assign node807 = (inp[9]) ? 4'b0101 : node808;
											assign node808 = (inp[8]) ? 4'b0101 : node809;
												assign node809 = (inp[11]) ? node811 : 4'b0111;
													assign node811 = (inp[1]) ? node813 : 4'b0111;
														assign node813 = (inp[15]) ? 4'b0101 : 4'b0111;
								assign node819 = (inp[14]) ? node821 : 4'b0101;
									assign node821 = (inp[8]) ? node823 : 4'b0101;
										assign node823 = (inp[9]) ? 4'b0011 : 4'b0101;
						assign node826 = (inp[4]) ? node840 : node827;
							assign node827 = (inp[9]) ? node829 : 4'b0101;
								assign node829 = (inp[2]) ? node831 : 4'b0101;
									assign node831 = (inp[8]) ? node833 : 4'b0101;
										assign node833 = (inp[14]) ? 4'b0011 : node834;
											assign node834 = (inp[15]) ? node836 : 4'b0101;
												assign node836 = (inp[7]) ? 4'b0111 : 4'b0101;
							assign node840 = (inp[14]) ? node852 : node841;
								assign node841 = (inp[2]) ? 4'b0111 : node842;
									assign node842 = (inp[9]) ? 4'b0111 : node843;
										assign node843 = (inp[8]) ? node845 : 4'b0101;
											assign node845 = (inp[7]) ? node847 : 4'b0101;
												assign node847 = (inp[15]) ? 4'b0111 : 4'b0101;
								assign node852 = (inp[2]) ? node854 : 4'b0011;
									assign node854 = (inp[9]) ? 4'b0001 : node855;
										assign node855 = (inp[8]) ? node857 : 4'b0011;
											assign node857 = (inp[7]) ? 4'b0001 : node858;
												assign node858 = (inp[3]) ? 4'b0011 : node859;
													assign node859 = (inp[11]) ? node861 : 4'b0011;
														assign node861 = (inp[0]) ? 4'b0011 : 4'b0001;
					assign node867 = (inp[14]) ? node923 : node868;
						assign node868 = (inp[13]) ? node890 : node869;
							assign node869 = (inp[4]) ? node879 : node870;
								assign node870 = (inp[2]) ? node872 : 4'b0011;
									assign node872 = (inp[9]) ? node874 : 4'b0011;
										assign node874 = (inp[7]) ? 4'b0001 : node875;
											assign node875 = (inp[8]) ? 4'b0001 : 4'b0011;
								assign node879 = (inp[2]) ? 4'b0011 : node880;
									assign node880 = (inp[8]) ? node882 : 4'b0001;
										assign node882 = (inp[15]) ? node884 : 4'b0001;
											assign node884 = (inp[7]) ? node886 : 4'b0001;
												assign node886 = (inp[9]) ? 4'b0011 : 4'b0001;
							assign node890 = (inp[7]) ? node902 : node891;
								assign node891 = (inp[9]) ? node897 : node892;
									assign node892 = (inp[4]) ? node894 : 4'b0001;
										assign node894 = (inp[2]) ? 4'b0001 : 4'b0011;
									assign node897 = (inp[2]) ? node899 : 4'b0001;
										assign node899 = (inp[4]) ? 4'b0001 : 4'b0011;
								assign node902 = (inp[2]) ? node914 : node903;
									assign node903 = (inp[9]) ? 4'b0001 : node904;
										assign node904 = (inp[4]) ? node906 : 4'b0001;
											assign node906 = (inp[8]) ? node908 : 4'b0011;
												assign node908 = (inp[15]) ? node910 : 4'b0011;
													assign node910 = (inp[1]) ? 4'b0001 : 4'b0011;
									assign node914 = (inp[4]) ? 4'b0001 : node915;
										assign node915 = (inp[9]) ? 4'b0011 : node916;
											assign node916 = (inp[15]) ? node918 : 4'b0001;
												assign node918 = (inp[8]) ? 4'b0011 : 4'b0001;
						assign node923 = (inp[4]) ? node941 : node924;
							assign node924 = (inp[2]) ? node928 : node925;
								assign node925 = (inp[13]) ? 4'b0001 : 4'b0011;
								assign node928 = (inp[13]) ? 4'b0111 : node929;
									assign node929 = (inp[9]) ? 4'b0001 : node930;
										assign node930 = (inp[8]) ? 4'b0001 : node931;
											assign node931 = (inp[1]) ? node933 : 4'b0011;
												assign node933 = (inp[15]) ? node935 : 4'b0011;
													assign node935 = (inp[11]) ? 4'b0001 : 4'b0011;
							assign node941 = (inp[2]) ? node953 : node942;
								assign node942 = (inp[13]) ? node944 : 4'b0110;
									assign node944 = (inp[9]) ? node946 : 4'b0100;
										assign node946 = (inp[7]) ? node948 : 4'b0100;
											assign node948 = (inp[8]) ? node950 : 4'b0100;
												assign node950 = (inp[15]) ? 4'b0110 : 4'b0100;
								assign node953 = (inp[9]) ? node967 : node954;
									assign node954 = (inp[0]) ? 4'b0110 : node955;
										assign node955 = (inp[1]) ? node957 : 4'b0110;
											assign node957 = (inp[11]) ? node959 : 4'b0110;
												assign node959 = (inp[7]) ? node961 : 4'b0110;
													assign node961 = (inp[8]) ? node963 : 4'b0110;
														assign node963 = (inp[3]) ? 4'b0100 : 4'b0110;
									assign node967 = (inp[13]) ? 4'b0110 : 4'b0100;
				assign node970 = (inp[4]) ? node1104 : node971;
					assign node971 = (inp[14]) ? node1039 : node972;
						assign node972 = (inp[13]) ? node1012 : node973;
							assign node973 = (inp[2]) ? node997 : node974;
								assign node974 = (inp[9]) ? 4'b0100 : node975;
									assign node975 = (inp[8]) ? node985 : node976;
										assign node976 = (inp[6]) ? node978 : 4'b0110;
											assign node978 = (inp[11]) ? node980 : 4'b0110;
												assign node980 = (inp[1]) ? node982 : 4'b0110;
													assign node982 = (inp[15]) ? 4'b0100 : 4'b0110;
										assign node985 = (inp[6]) ? 4'b0100 : node986;
											assign node986 = (inp[7]) ? 4'b0100 : node987;
												assign node987 = (inp[1]) ? node989 : 4'b0110;
													assign node989 = (inp[15]) ? node991 : 4'b0110;
														assign node991 = (inp[11]) ? 4'b0100 : 4'b0110;
								assign node997 = (inp[9]) ? node1007 : node998;
									assign node998 = (inp[0]) ? node1000 : 4'b0100;
										assign node1000 = (inp[1]) ? node1002 : 4'b0100;
											assign node1002 = (inp[7]) ? node1004 : 4'b0100;
												assign node1004 = (inp[8]) ? 4'b0110 : 4'b0100;
									assign node1007 = (inp[6]) ? 4'b0110 : node1008;
										assign node1008 = (inp[8]) ? 4'b0010 : 4'b0100;
							assign node1012 = (inp[6]) ? node1022 : node1013;
								assign node1013 = (inp[2]) ? node1015 : 4'b0010;
									assign node1015 = (inp[8]) ? 4'b0000 : node1016;
										assign node1016 = (inp[9]) ? 4'b0000 : node1017;
											assign node1017 = (inp[7]) ? 4'b0000 : 4'b0010;
								assign node1022 = (inp[2]) ? node1034 : node1023;
									assign node1023 = (inp[9]) ? node1025 : 4'b0110;
										assign node1025 = (inp[7]) ? 4'b0100 : node1026;
											assign node1026 = (inp[8]) ? 4'b0100 : node1027;
												assign node1027 = (inp[15]) ? node1029 : 4'b0110;
													assign node1029 = (inp[11]) ? 4'b0100 : 4'b0110;
									assign node1034 = (inp[9]) ? node1036 : 4'b0100;
										assign node1036 = (inp[8]) ? 4'b0010 : 4'b0100;
						assign node1039 = (inp[13]) ? node1089 : node1040;
							assign node1040 = (inp[2]) ? node1066 : node1041;
								assign node1041 = (inp[6]) ? node1051 : node1042;
									assign node1042 = (inp[9]) ? 4'b0010 : node1043;
										assign node1043 = (inp[8]) ? node1045 : 4'b0000;
											assign node1045 = (inp[15]) ? node1047 : 4'b0000;
												assign node1047 = (inp[7]) ? 4'b0010 : 4'b0000;
									assign node1051 = (inp[8]) ? node1053 : 4'b0010;
										assign node1053 = (inp[7]) ? node1063 : node1054;
											assign node1054 = (inp[1]) ? node1056 : 4'b0010;
												assign node1056 = (inp[11]) ? node1058 : 4'b0010;
													assign node1058 = (inp[0]) ? 4'b0010 : node1059;
														assign node1059 = (inp[9]) ? 4'b0000 : 4'b0010;
											assign node1063 = (inp[9]) ? 4'b0000 : 4'b0010;
								assign node1066 = (inp[6]) ? node1080 : node1067;
									assign node1067 = (inp[9]) ? node1069 : 4'b0010;
										assign node1069 = (inp[8]) ? 4'b0000 : node1070;
											assign node1070 = (inp[1]) ? node1072 : 4'b0010;
												assign node1072 = (inp[15]) ? node1074 : 4'b0010;
													assign node1074 = (inp[0]) ? 4'b0010 : node1075;
														assign node1075 = (inp[11]) ? 4'b0000 : 4'b0010;
									assign node1080 = (inp[15]) ? node1082 : 4'b0000;
										assign node1082 = (inp[8]) ? node1084 : 4'b0000;
											assign node1084 = (inp[9]) ? node1086 : 4'b0000;
												assign node1086 = (inp[7]) ? 4'b0010 : 4'b0000;
							assign node1089 = (inp[2]) ? node1101 : node1090;
								assign node1090 = (inp[6]) ? node1092 : 4'b0000;
									assign node1092 = (inp[9]) ? node1094 : 4'b0010;
										assign node1094 = (inp[1]) ? node1096 : 4'b0010;
											assign node1096 = (inp[3]) ? node1098 : 4'b0010;
												assign node1098 = (inp[15]) ? 4'b0000 : 4'b0010;
								assign node1101 = (inp[6]) ? 4'b0000 : 4'b0110;
					assign node1104 = (inp[14]) ? node1192 : node1105;
						assign node1105 = (inp[6]) ? node1127 : node1106;
							assign node1106 = (inp[2]) ? node1116 : node1107;
								assign node1107 = (inp[8]) ? node1109 : 4'b0111;
									assign node1109 = (inp[9]) ? node1111 : 4'b0111;
										assign node1111 = (inp[13]) ? node1113 : 4'b0111;
											assign node1113 = (inp[7]) ? 4'b0101 : 4'b0111;
								assign node1116 = (inp[8]) ? node1118 : 4'b0101;
									assign node1118 = (inp[9]) ? node1120 : 4'b0101;
										assign node1120 = (inp[13]) ? 4'b0011 : node1121;
											assign node1121 = (inp[7]) ? node1123 : 4'b0101;
												assign node1123 = (inp[15]) ? 4'b0111 : 4'b0101;
							assign node1127 = (inp[13]) ? node1171 : node1128;
								assign node1128 = (inp[9]) ? node1164 : node1129;
									assign node1129 = (inp[1]) ? node1143 : node1130;
										assign node1130 = (inp[2]) ? node1138 : node1131;
											assign node1131 = (inp[15]) ? node1133 : 4'b0101;
												assign node1133 = (inp[3]) ? node1135 : 4'b0101;
													assign node1135 = (inp[7]) ? 4'b0111 : 4'b0101;
											assign node1138 = (inp[8]) ? 4'b0101 : node1139;
												assign node1139 = (inp[7]) ? 4'b0101 : 4'b0111;
										assign node1143 = (inp[11]) ? node1155 : node1144;
											assign node1144 = (inp[0]) ? 4'b0101 : node1145;
												assign node1145 = (inp[7]) ? node1151 : node1146;
													assign node1146 = (inp[8]) ? 4'b0101 : node1147;
														assign node1147 = (inp[2]) ? 4'b0111 : 4'b0101;
													assign node1151 = (inp[8]) ? 4'b0111 : 4'b0101;
											assign node1155 = (inp[8]) ? node1161 : node1156;
												assign node1156 = (inp[7]) ? 4'b0101 : node1157;
													assign node1157 = (inp[2]) ? 4'b0111 : 4'b0101;
												assign node1161 = (inp[7]) ? 4'b0111 : 4'b0101;
									assign node1164 = (inp[8]) ? node1168 : node1165;
										assign node1165 = (inp[2]) ? 4'b0101 : 4'b0111;
										assign node1168 = (inp[2]) ? 4'b0011 : 4'b0111;
								assign node1171 = (inp[9]) ? node1183 : node1172;
									assign node1172 = (inp[7]) ? node1174 : 4'b0011;
										assign node1174 = (inp[8]) ? node1176 : 4'b0011;
											assign node1176 = (inp[2]) ? node1178 : 4'b0001;
												assign node1178 = (inp[3]) ? 4'b0011 : node1179;
													assign node1179 = (inp[1]) ? 4'b0001 : 4'b0011;
									assign node1183 = (inp[15]) ? node1185 : 4'b0001;
										assign node1185 = (inp[2]) ? 4'b0001 : node1186;
											assign node1186 = (inp[7]) ? node1188 : 4'b0001;
												assign node1188 = (inp[1]) ? 4'b0011 : 4'b0001;
						assign node1192 = (inp[6]) ? node1242 : node1193;
							assign node1193 = (inp[2]) ? node1219 : node1194;
								assign node1194 = (inp[9]) ? node1208 : node1195;
									assign node1195 = (inp[8]) ? node1205 : node1196;
										assign node1196 = (inp[0]) ? 4'b0011 : node1197;
											assign node1197 = (inp[15]) ? node1199 : 4'b0011;
												assign node1199 = (inp[3]) ? node1201 : 4'b0011;
													assign node1201 = (inp[13]) ? 4'b0001 : 4'b0011;
										assign node1205 = (inp[13]) ? 4'b0001 : 4'b0011;
									assign node1208 = (inp[13]) ? 4'b0001 : node1209;
										assign node1209 = (inp[8]) ? 4'b0001 : node1210;
											assign node1210 = (inp[7]) ? 4'b0001 : node1211;
												assign node1211 = (inp[15]) ? node1213 : 4'b0011;
													assign node1213 = (inp[11]) ? 4'b0001 : 4'b0011;
								assign node1219 = (inp[13]) ? node1229 : node1220;
									assign node1220 = (inp[9]) ? 4'b0011 : node1221;
										assign node1221 = (inp[8]) ? node1223 : 4'b0001;
											assign node1223 = (inp[15]) ? node1225 : 4'b0001;
												assign node1225 = (inp[7]) ? 4'b0011 : 4'b0001;
									assign node1229 = (inp[8]) ? node1239 : node1230;
										assign node1230 = (inp[1]) ? node1232 : 4'b0111;
											assign node1232 = (inp[9]) ? node1234 : 4'b0111;
												assign node1234 = (inp[3]) ? node1236 : 4'b0111;
													assign node1236 = (inp[7]) ? 4'b0101 : 4'b0111;
										assign node1239 = (inp[9]) ? 4'b0101 : 4'b0111;
							assign node1242 = (inp[13]) ? node1270 : node1243;
								assign node1243 = (inp[9]) ? node1261 : node1244;
									assign node1244 = (inp[8]) ? node1246 : 4'b0110;
										assign node1246 = (inp[2]) ? node1254 : node1247;
											assign node1247 = (inp[15]) ? node1249 : 4'b0110;
												assign node1249 = (inp[11]) ? node1251 : 4'b0110;
													assign node1251 = (inp[1]) ? 4'b0100 : 4'b0110;
											assign node1254 = (inp[7]) ? 4'b0100 : node1255;
												assign node1255 = (inp[1]) ? node1257 : 4'b0110;
													assign node1257 = (inp[15]) ? 4'b0100 : 4'b0110;
									assign node1261 = (inp[8]) ? node1263 : 4'b0100;
										assign node1263 = (inp[2]) ? 4'b0010 : node1264;
											assign node1264 = (inp[7]) ? node1266 : 4'b0100;
												assign node1266 = (inp[15]) ? 4'b0110 : 4'b0100;
								assign node1270 = (inp[2]) ? node1290 : node1271;
									assign node1271 = (inp[8]) ? node1283 : node1272;
										assign node1272 = (inp[9]) ? node1276 : node1273;
											assign node1273 = (inp[7]) ? 4'b0000 : 4'b0010;
											assign node1276 = (inp[15]) ? node1278 : 4'b0010;
												assign node1278 = (inp[1]) ? node1280 : 4'b0010;
													assign node1280 = (inp[11]) ? 4'b0000 : 4'b0010;
										assign node1283 = (inp[9]) ? 4'b0000 : node1284;
											assign node1284 = (inp[7]) ? node1286 : 4'b0000;
												assign node1286 = (inp[15]) ? 4'b0010 : 4'b0000;
									assign node1290 = (inp[8]) ? node1308 : node1291;
										assign node1291 = (inp[9]) ? node1301 : node1292;
											assign node1292 = (inp[0]) ? 4'b0110 : node1293;
												assign node1293 = (inp[7]) ? node1295 : 4'b0110;
													assign node1295 = (inp[15]) ? node1297 : 4'b0110;
														assign node1297 = (inp[1]) ? 4'b0100 : 4'b0110;
											assign node1301 = (inp[7]) ? 4'b0100 : node1302;
												assign node1302 = (inp[11]) ? node1304 : 4'b0110;
													assign node1304 = (inp[15]) ? 4'b0100 : 4'b0110;
										assign node1308 = (inp[9]) ? node1314 : node1309;
											assign node1309 = (inp[15]) ? node1311 : 4'b0100;
												assign node1311 = (inp[7]) ? 4'b0110 : 4'b0100;
											assign node1314 = (inp[15]) ? 4'b0010 : node1315;
												assign node1315 = (inp[7]) ? 4'b0000 : 4'b0010;

endmodule