module dtc_split5_bm89 (
	input  wire [12-1:0] inp,
	output wire [3-1:0] outp
);

	wire [3-1:0] node1;
	wire [3-1:0] node2;
	wire [3-1:0] node3;
	wire [3-1:0] node4;
	wire [3-1:0] node5;
	wire [3-1:0] node6;
	wire [3-1:0] node7;
	wire [3-1:0] node8;
	wire [3-1:0] node10;
	wire [3-1:0] node14;
	wire [3-1:0] node15;
	wire [3-1:0] node16;
	wire [3-1:0] node17;
	wire [3-1:0] node18;
	wire [3-1:0] node22;
	wire [3-1:0] node25;
	wire [3-1:0] node28;
	wire [3-1:0] node29;
	wire [3-1:0] node30;
	wire [3-1:0] node36;
	wire [3-1:0] node37;
	wire [3-1:0] node38;
	wire [3-1:0] node41;
	wire [3-1:0] node42;
	wire [3-1:0] node43;
	wire [3-1:0] node47;
	wire [3-1:0] node50;
	wire [3-1:0] node51;
	wire [3-1:0] node52;
	wire [3-1:0] node53;
	wire [3-1:0] node57;
	wire [3-1:0] node58;
	wire [3-1:0] node60;
	wire [3-1:0] node64;
	wire [3-1:0] node65;
	wire [3-1:0] node66;
	wire [3-1:0] node67;
	wire [3-1:0] node71;
	wire [3-1:0] node73;
	wire [3-1:0] node76;
	wire [3-1:0] node78;
	wire [3-1:0] node82;
	wire [3-1:0] node83;
	wire [3-1:0] node84;
	wire [3-1:0] node85;
	wire [3-1:0] node86;
	wire [3-1:0] node87;
	wire [3-1:0] node88;
	wire [3-1:0] node91;
	wire [3-1:0] node93;
	wire [3-1:0] node96;
	wire [3-1:0] node99;
	wire [3-1:0] node100;
	wire [3-1:0] node101;
	wire [3-1:0] node104;
	wire [3-1:0] node107;
	wire [3-1:0] node108;
	wire [3-1:0] node112;
	wire [3-1:0] node113;
	wire [3-1:0] node114;
	wire [3-1:0] node115;
	wire [3-1:0] node117;
	wire [3-1:0] node121;
	wire [3-1:0] node122;
	wire [3-1:0] node126;
	wire [3-1:0] node128;
	wire [3-1:0] node129;
	wire [3-1:0] node133;
	wire [3-1:0] node134;
	wire [3-1:0] node135;
	wire [3-1:0] node136;
	wire [3-1:0] node138;
	wire [3-1:0] node141;
	wire [3-1:0] node142;
	wire [3-1:0] node144;
	wire [3-1:0] node148;
	wire [3-1:0] node150;
	wire [3-1:0] node152;
	wire [3-1:0] node155;
	wire [3-1:0] node156;
	wire [3-1:0] node158;
	wire [3-1:0] node160;
	wire [3-1:0] node162;
	wire [3-1:0] node165;
	wire [3-1:0] node166;
	wire [3-1:0] node169;
	wire [3-1:0] node170;
	wire [3-1:0] node174;
	wire [3-1:0] node175;
	wire [3-1:0] node176;
	wire [3-1:0] node177;
	wire [3-1:0] node178;
	wire [3-1:0] node179;
	wire [3-1:0] node181;
	wire [3-1:0] node183;
	wire [3-1:0] node186;
	wire [3-1:0] node189;
	wire [3-1:0] node190;
	wire [3-1:0] node192;
	wire [3-1:0] node195;
	wire [3-1:0] node198;
	wire [3-1:0] node199;
	wire [3-1:0] node200;
	wire [3-1:0] node203;
	wire [3-1:0] node205;
	wire [3-1:0] node208;
	wire [3-1:0] node209;
	wire [3-1:0] node211;
	wire [3-1:0] node213;
	wire [3-1:0] node216;
	wire [3-1:0] node218;
	wire [3-1:0] node222;
	wire [3-1:0] node223;
	wire [3-1:0] node224;
	wire [3-1:0] node226;
	wire [3-1:0] node228;
	wire [3-1:0] node231;
	wire [3-1:0] node232;
	wire [3-1:0] node233;
	wire [3-1:0] node235;
	wire [3-1:0] node238;
	wire [3-1:0] node240;
	wire [3-1:0] node243;
	wire [3-1:0] node245;
	wire [3-1:0] node248;
	wire [3-1:0] node249;
	wire [3-1:0] node250;
	wire [3-1:0] node252;
	wire [3-1:0] node255;
	wire [3-1:0] node257;
	wire [3-1:0] node260;
	wire [3-1:0] node261;
	wire [3-1:0] node264;
	wire [3-1:0] node266;
	wire [3-1:0] node269;
	wire [3-1:0] node270;
	wire [3-1:0] node271;
	wire [3-1:0] node272;
	wire [3-1:0] node273;
	wire [3-1:0] node274;
	wire [3-1:0] node275;
	wire [3-1:0] node277;
	wire [3-1:0] node279;
	wire [3-1:0] node283;
	wire [3-1:0] node284;
	wire [3-1:0] node285;
	wire [3-1:0] node288;
	wire [3-1:0] node291;
	wire [3-1:0] node292;
	wire [3-1:0] node294;
	wire [3-1:0] node297;
	wire [3-1:0] node302;
	wire [3-1:0] node303;
	wire [3-1:0] node304;
	wire [3-1:0] node305;
	wire [3-1:0] node306;
	wire [3-1:0] node307;
	wire [3-1:0] node310;
	wire [3-1:0] node312;
	wire [3-1:0] node315;
	wire [3-1:0] node316;
	wire [3-1:0] node320;
	wire [3-1:0] node321;
	wire [3-1:0] node322;
	wire [3-1:0] node325;
	wire [3-1:0] node326;
	wire [3-1:0] node330;
	wire [3-1:0] node331;
	wire [3-1:0] node332;
	wire [3-1:0] node335;
	wire [3-1:0] node339;
	wire [3-1:0] node340;
	wire [3-1:0] node343;
	wire [3-1:0] node344;
	wire [3-1:0] node345;
	wire [3-1:0] node346;
	wire [3-1:0] node351;
	wire [3-1:0] node352;
	wire [3-1:0] node354;
	wire [3-1:0] node357;
	wire [3-1:0] node360;
	wire [3-1:0] node361;
	wire [3-1:0] node362;
	wire [3-1:0] node363;
	wire [3-1:0] node365;
	wire [3-1:0] node369;
	wire [3-1:0] node370;
	wire [3-1:0] node371;
	wire [3-1:0] node375;
	wire [3-1:0] node376;
	wire [3-1:0] node381;
	wire [3-1:0] node382;
	wire [3-1:0] node383;
	wire [3-1:0] node384;
	wire [3-1:0] node385;
	wire [3-1:0] node387;
	wire [3-1:0] node388;
	wire [3-1:0] node391;
	wire [3-1:0] node393;
	wire [3-1:0] node396;
	wire [3-1:0] node398;
	wire [3-1:0] node402;
	wire [3-1:0] node403;
	wire [3-1:0] node404;
	wire [3-1:0] node405;
	wire [3-1:0] node407;
	wire [3-1:0] node410;
	wire [3-1:0] node413;
	wire [3-1:0] node414;
	wire [3-1:0] node415;
	wire [3-1:0] node418;
	wire [3-1:0] node419;
	wire [3-1:0] node422;
	wire [3-1:0] node424;
	wire [3-1:0] node427;
	wire [3-1:0] node428;
	wire [3-1:0] node429;
	wire [3-1:0] node432;
	wire [3-1:0] node434;
	wire [3-1:0] node437;
	wire [3-1:0] node440;
	wire [3-1:0] node441;
	wire [3-1:0] node443;
	wire [3-1:0] node445;
	wire [3-1:0] node448;
	wire [3-1:0] node449;
	wire [3-1:0] node452;
	wire [3-1:0] node454;
	wire [3-1:0] node457;
	wire [3-1:0] node458;
	wire [3-1:0] node459;
	wire [3-1:0] node460;
	wire [3-1:0] node463;
	wire [3-1:0] node465;
	wire [3-1:0] node466;
	wire [3-1:0] node468;
	wire [3-1:0] node469;
	wire [3-1:0] node474;
	wire [3-1:0] node475;
	wire [3-1:0] node477;
	wire [3-1:0] node479;
	wire [3-1:0] node482;
	wire [3-1:0] node484;
	wire [3-1:0] node486;
	wire [3-1:0] node487;
	wire [3-1:0] node490;
	wire [3-1:0] node493;
	wire [3-1:0] node494;
	wire [3-1:0] node495;
	wire [3-1:0] node496;
	wire [3-1:0] node498;
	wire [3-1:0] node499;
	wire [3-1:0] node503;
	wire [3-1:0] node505;
	wire [3-1:0] node508;
	wire [3-1:0] node509;
	wire [3-1:0] node510;
	wire [3-1:0] node512;
	wire [3-1:0] node516;
	wire [3-1:0] node518;
	wire [3-1:0] node521;
	wire [3-1:0] node522;
	wire [3-1:0] node523;
	wire [3-1:0] node525;
	wire [3-1:0] node528;
	wire [3-1:0] node530;
	wire [3-1:0] node531;
	wire [3-1:0] node534;
	wire [3-1:0] node536;
	wire [3-1:0] node539;
	wire [3-1:0] node540;
	wire [3-1:0] node542;
	wire [3-1:0] node545;
	wire [3-1:0] node546;
	wire [3-1:0] node550;
	wire [3-1:0] node551;
	wire [3-1:0] node552;
	wire [3-1:0] node553;
	wire [3-1:0] node554;
	wire [3-1:0] node555;
	wire [3-1:0] node556;
	wire [3-1:0] node559;
	wire [3-1:0] node560;
	wire [3-1:0] node562;
	wire [3-1:0] node563;
	wire [3-1:0] node566;
	wire [3-1:0] node569;
	wire [3-1:0] node570;
	wire [3-1:0] node572;
	wire [3-1:0] node576;
	wire [3-1:0] node577;
	wire [3-1:0] node578;
	wire [3-1:0] node579;
	wire [3-1:0] node582;
	wire [3-1:0] node584;
	wire [3-1:0] node587;
	wire [3-1:0] node588;
	wire [3-1:0] node590;
	wire [3-1:0] node593;
	wire [3-1:0] node596;
	wire [3-1:0] node597;
	wire [3-1:0] node598;
	wire [3-1:0] node601;
	wire [3-1:0] node602;
	wire [3-1:0] node603;
	wire [3-1:0] node608;
	wire [3-1:0] node609;
	wire [3-1:0] node610;
	wire [3-1:0] node615;
	wire [3-1:0] node617;
	wire [3-1:0] node618;
	wire [3-1:0] node619;
	wire [3-1:0] node621;
	wire [3-1:0] node624;
	wire [3-1:0] node625;
	wire [3-1:0] node627;
	wire [3-1:0] node630;
	wire [3-1:0] node632;
	wire [3-1:0] node633;
	wire [3-1:0] node636;
	wire [3-1:0] node639;
	wire [3-1:0] node640;
	wire [3-1:0] node642;
	wire [3-1:0] node645;
	wire [3-1:0] node646;
	wire [3-1:0] node649;
	wire [3-1:0] node650;
	wire [3-1:0] node653;
	wire [3-1:0] node656;
	wire [3-1:0] node658;
	wire [3-1:0] node660;
	wire [3-1:0] node661;
	wire [3-1:0] node663;
	wire [3-1:0] node668;
	wire [3-1:0] node669;
	wire [3-1:0] node670;
	wire [3-1:0] node671;
	wire [3-1:0] node672;
	wire [3-1:0] node673;
	wire [3-1:0] node674;
	wire [3-1:0] node677;
	wire [3-1:0] node679;
	wire [3-1:0] node682;
	wire [3-1:0] node683;
	wire [3-1:0] node686;
	wire [3-1:0] node687;
	wire [3-1:0] node689;
	wire [3-1:0] node694;
	wire [3-1:0] node695;
	wire [3-1:0] node696;
	wire [3-1:0] node697;
	wire [3-1:0] node698;
	wire [3-1:0] node699;
	wire [3-1:0] node704;
	wire [3-1:0] node705;
	wire [3-1:0] node708;
	wire [3-1:0] node711;
	wire [3-1:0] node712;
	wire [3-1:0] node713;
	wire [3-1:0] node715;
	wire [3-1:0] node718;
	wire [3-1:0] node721;
	wire [3-1:0] node722;
	wire [3-1:0] node725;
	wire [3-1:0] node728;
	wire [3-1:0] node729;
	wire [3-1:0] node730;
	wire [3-1:0] node731;
	wire [3-1:0] node732;
	wire [3-1:0] node736;
	wire [3-1:0] node739;
	wire [3-1:0] node740;
	wire [3-1:0] node741;
	wire [3-1:0] node743;
	wire [3-1:0] node746;
	wire [3-1:0] node748;
	wire [3-1:0] node751;
	wire [3-1:0] node752;
	wire [3-1:0] node755;
	wire [3-1:0] node758;
	wire [3-1:0] node759;
	wire [3-1:0] node760;
	wire [3-1:0] node764;
	wire [3-1:0] node765;
	wire [3-1:0] node767;
	wire [3-1:0] node769;
	wire [3-1:0] node772;
	wire [3-1:0] node774;
	wire [3-1:0] node777;
	wire [3-1:0] node778;
	wire [3-1:0] node779;
	wire [3-1:0] node780;
	wire [3-1:0] node782;
	wire [3-1:0] node783;
	wire [3-1:0] node784;
	wire [3-1:0] node789;
	wire [3-1:0] node791;
	wire [3-1:0] node792;
	wire [3-1:0] node796;
	wire [3-1:0] node797;
	wire [3-1:0] node798;
	wire [3-1:0] node800;
	wire [3-1:0] node802;
	wire [3-1:0] node806;
	wire [3-1:0] node807;
	wire [3-1:0] node809;
	wire [3-1:0] node810;
	wire [3-1:0] node814;
	wire [3-1:0] node815;
	wire [3-1:0] node819;
	wire [3-1:0] node820;
	wire [3-1:0] node821;
	wire [3-1:0] node822;
	wire [3-1:0] node824;
	wire [3-1:0] node827;
	wire [3-1:0] node829;
	wire [3-1:0] node832;
	wire [3-1:0] node833;
	wire [3-1:0] node834;
	wire [3-1:0] node836;
	wire [3-1:0] node839;
	wire [3-1:0] node842;
	wire [3-1:0] node844;
	wire [3-1:0] node847;
	wire [3-1:0] node848;
	wire [3-1:0] node849;
	wire [3-1:0] node851;
	wire [3-1:0] node855;
	wire [3-1:0] node856;
	wire [3-1:0] node858;
	wire [3-1:0] node859;
	wire [3-1:0] node863;
	wire [3-1:0] node866;
	wire [3-1:0] node867;
	wire [3-1:0] node868;
	wire [3-1:0] node869;
	wire [3-1:0] node870;
	wire [3-1:0] node871;
	wire [3-1:0] node873;
	wire [3-1:0] node874;
	wire [3-1:0] node878;
	wire [3-1:0] node880;
	wire [3-1:0] node881;
	wire [3-1:0] node884;
	wire [3-1:0] node887;
	wire [3-1:0] node889;
	wire [3-1:0] node891;
	wire [3-1:0] node894;
	wire [3-1:0] node895;
	wire [3-1:0] node897;
	wire [3-1:0] node901;
	wire [3-1:0] node902;
	wire [3-1:0] node903;
	wire [3-1:0] node904;
	wire [3-1:0] node905;
	wire [3-1:0] node909;
	wire [3-1:0] node910;
	wire [3-1:0] node912;
	wire [3-1:0] node916;
	wire [3-1:0] node917;
	wire [3-1:0] node919;
	wire [3-1:0] node922;
	wire [3-1:0] node924;
	wire [3-1:0] node926;
	wire [3-1:0] node929;
	wire [3-1:0] node931;
	wire [3-1:0] node932;
	wire [3-1:0] node933;
	wire [3-1:0] node935;
	wire [3-1:0] node939;
	wire [3-1:0] node940;
	wire [3-1:0] node942;
	wire [3-1:0] node945;
	wire [3-1:0] node946;
	wire [3-1:0] node950;
	wire [3-1:0] node952;
	wire [3-1:0] node953;
	wire [3-1:0] node954;
	wire [3-1:0] node955;
	wire [3-1:0] node957;
	wire [3-1:0] node961;
	wire [3-1:0] node962;
	wire [3-1:0] node964;
	wire [3-1:0] node965;
	wire [3-1:0] node968;
	wire [3-1:0] node970;
	wire [3-1:0] node973;
	wire [3-1:0] node974;
	wire [3-1:0] node978;
	wire [3-1:0] node979;
	wire [3-1:0] node980;
	wire [3-1:0] node982;

	assign outp = (inp[3]) ? node550 : node1;
		assign node1 = (inp[6]) ? node269 : node2;
			assign node2 = (inp[7]) ? node82 : node3;
				assign node3 = (inp[9]) ? 3'b111 : node4;
					assign node4 = (inp[4]) ? node36 : node5;
						assign node5 = (inp[10]) ? 3'b111 : node6;
							assign node6 = (inp[8]) ? node14 : node7;
								assign node7 = (inp[5]) ? 3'b011 : node8;
									assign node8 = (inp[0]) ? node10 : 3'b101;
										assign node10 = (inp[2]) ? 3'b011 : 3'b101;
								assign node14 = (inp[2]) ? node28 : node15;
									assign node15 = (inp[0]) ? node25 : node16;
										assign node16 = (inp[1]) ? node22 : node17;
											assign node17 = (inp[11]) ? 3'b101 : node18;
												assign node18 = (inp[5]) ? 3'b011 : 3'b101;
											assign node22 = (inp[11]) ? 3'b011 : 3'b101;
										assign node25 = (inp[11]) ? 3'b101 : 3'b011;
									assign node28 = (inp[1]) ? 3'b101 : node29;
										assign node29 = (inp[5]) ? 3'b101 : node30;
											assign node30 = (inp[11]) ? 3'b011 : 3'b101;
						assign node36 = (inp[10]) ? node50 : node37;
							assign node37 = (inp[11]) ? node41 : node38;
								assign node38 = (inp[8]) ? 3'b100 : 3'b010;
								assign node41 = (inp[1]) ? node47 : node42;
									assign node42 = (inp[0]) ? 3'b110 : node43;
										assign node43 = (inp[2]) ? 3'b110 : 3'b001;
									assign node47 = (inp[8]) ? 3'b010 : 3'b110;
							assign node50 = (inp[5]) ? node64 : node51;
								assign node51 = (inp[8]) ? node57 : node52;
									assign node52 = (inp[11]) ? 3'b011 : node53;
										assign node53 = (inp[1]) ? 3'b001 : 3'b101;
									assign node57 = (inp[11]) ? 3'b101 : node58;
										assign node58 = (inp[1]) ? node60 : 3'b001;
											assign node60 = (inp[2]) ? 3'b110 : 3'b001;
								assign node64 = (inp[11]) ? node76 : node65;
									assign node65 = (inp[8]) ? node71 : node66;
										assign node66 = (inp[2]) ? 3'b101 : node67;
											assign node67 = (inp[0]) ? 3'b001 : 3'b101;
										assign node71 = (inp[1]) ? node73 : 3'b001;
											assign node73 = (inp[0]) ? 3'b110 : 3'b001;
									assign node76 = (inp[0]) ? node78 : 3'b101;
										assign node78 = (inp[8]) ? 3'b001 : 3'b101;
				assign node82 = (inp[10]) ? node174 : node83;
					assign node83 = (inp[4]) ? node133 : node84;
						assign node84 = (inp[9]) ? node112 : node85;
							assign node85 = (inp[11]) ? node99 : node86;
								assign node86 = (inp[8]) ? node96 : node87;
									assign node87 = (inp[0]) ? node91 : node88;
										assign node88 = (inp[5]) ? 3'b110 : 3'b010;
										assign node91 = (inp[1]) ? node93 : 3'b110;
											assign node93 = (inp[2]) ? 3'b110 : 3'b010;
									assign node96 = (inp[5]) ? 3'b000 : 3'b010;
								assign node99 = (inp[8]) ? node107 : node100;
									assign node100 = (inp[2]) ? node104 : node101;
										assign node101 = (inp[5]) ? 3'b001 : 3'b011;
										assign node104 = (inp[5]) ? 3'b011 : 3'b001;
									assign node107 = (inp[2]) ? 3'b110 : node108;
										assign node108 = (inp[5]) ? 3'b110 : 3'b001;
							assign node112 = (inp[5]) ? node126 : node113;
								assign node113 = (inp[11]) ? node121 : node114;
									assign node114 = (inp[2]) ? 3'b110 : node115;
										assign node115 = (inp[8]) ? node117 : 3'b110;
											assign node117 = (inp[0]) ? 3'b000 : 3'b110;
									assign node121 = (inp[8]) ? 3'b000 : node122;
										assign node122 = (inp[2]) ? 3'b000 : 3'b110;
								assign node126 = (inp[11]) ? node128 : 3'b000;
									assign node128 = (inp[2]) ? 3'b110 : node129;
										assign node129 = (inp[1]) ? 3'b000 : 3'b110;
						assign node133 = (inp[9]) ? node155 : node134;
							assign node134 = (inp[5]) ? node148 : node135;
								assign node135 = (inp[8]) ? node141 : node136;
									assign node136 = (inp[11]) ? node138 : 3'b100;
										assign node138 = (inp[1]) ? 3'b010 : 3'b100;
									assign node141 = (inp[2]) ? 3'b100 : node142;
										assign node142 = (inp[1]) ? node144 : 3'b000;
											assign node144 = (inp[11]) ? 3'b100 : 3'b000;
								assign node148 = (inp[11]) ? node150 : 3'b000;
									assign node150 = (inp[2]) ? node152 : 3'b100;
										assign node152 = (inp[1]) ? 3'b100 : 3'b010;
							assign node155 = (inp[8]) ? node165 : node156;
								assign node156 = (inp[11]) ? node158 : 3'b001;
									assign node158 = (inp[2]) ? node160 : 3'b010;
										assign node160 = (inp[0]) ? node162 : 3'b101;
											assign node162 = (inp[5]) ? 3'b101 : 3'b100;
								assign node165 = (inp[11]) ? node169 : node166;
									assign node166 = (inp[5]) ? 3'b110 : 3'b111;
									assign node169 = (inp[1]) ? 3'b001 : node170;
										assign node170 = (inp[5]) ? 3'b101 : 3'b110;
					assign node174 = (inp[4]) ? node222 : node175;
						assign node175 = (inp[9]) ? 3'b100 : node176;
							assign node176 = (inp[8]) ? node198 : node177;
								assign node177 = (inp[11]) ? node189 : node178;
									assign node178 = (inp[2]) ? node186 : node179;
										assign node179 = (inp[0]) ? node181 : 3'b101;
											assign node181 = (inp[1]) ? node183 : 3'b101;
												assign node183 = (inp[5]) ? 3'b001 : 3'b101;
										assign node186 = (inp[0]) ? 3'b101 : 3'b001;
									assign node189 = (inp[5]) ? node195 : node190;
										assign node190 = (inp[0]) ? node192 : 3'b101;
											assign node192 = (inp[2]) ? 3'b011 : 3'b001;
										assign node195 = (inp[2]) ? 3'b001 : 3'b011;
								assign node198 = (inp[11]) ? node208 : node199;
									assign node199 = (inp[5]) ? node203 : node200;
										assign node200 = (inp[2]) ? 3'b001 : 3'b101;
										assign node203 = (inp[0]) ? node205 : 3'b010;
											assign node205 = (inp[2]) ? 3'b110 : 3'b010;
									assign node208 = (inp[5]) ? node216 : node209;
										assign node209 = (inp[2]) ? node211 : 3'b011;
											assign node211 = (inp[1]) ? node213 : 3'b111;
												assign node213 = (inp[0]) ? 3'b101 : 3'b111;
										assign node216 = (inp[1]) ? node218 : 3'b101;
											assign node218 = (inp[2]) ? 3'b001 : 3'b101;
						assign node222 = (inp[9]) ? node248 : node223;
							assign node223 = (inp[11]) ? node231 : node224;
								assign node224 = (inp[8]) ? node226 : 3'b110;
									assign node226 = (inp[0]) ? node228 : 3'b010;
										assign node228 = (inp[5]) ? 3'b100 : 3'b010;
								assign node231 = (inp[5]) ? node243 : node232;
									assign node232 = (inp[2]) ? node238 : node233;
										assign node233 = (inp[0]) ? node235 : 3'b001;
											assign node235 = (inp[8]) ? 3'b101 : 3'b001;
										assign node238 = (inp[8]) ? node240 : 3'b001;
											assign node240 = (inp[1]) ? 3'b110 : 3'b010;
									assign node243 = (inp[0]) ? node245 : 3'b110;
										assign node245 = (inp[8]) ? 3'b010 : 3'b110;
							assign node248 = (inp[8]) ? node260 : node249;
								assign node249 = (inp[11]) ? node255 : node250;
									assign node250 = (inp[2]) ? node252 : 3'b111;
										assign node252 = (inp[1]) ? 3'b011 : 3'b111;
									assign node255 = (inp[0]) ? node257 : 3'b001;
										assign node257 = (inp[5]) ? 3'b111 : 3'b001;
								assign node260 = (inp[11]) ? node264 : node261;
									assign node261 = (inp[2]) ? 3'b101 : 3'b011;
									assign node264 = (inp[0]) ? node266 : 3'b111;
										assign node266 = (inp[5]) ? 3'b011 : 3'b111;
			assign node269 = (inp[9]) ? node381 : node270;
				assign node270 = (inp[10]) ? node302 : node271;
					assign node271 = (inp[7]) ? 3'b000 : node272;
						assign node272 = (inp[4]) ? 3'b000 : node273;
							assign node273 = (inp[11]) ? node283 : node274;
								assign node274 = (inp[8]) ? 3'b000 : node275;
									assign node275 = (inp[5]) ? node277 : 3'b100;
										assign node277 = (inp[2]) ? node279 : 3'b100;
											assign node279 = (inp[0]) ? 3'b000 : 3'b100;
								assign node283 = (inp[5]) ? node291 : node284;
									assign node284 = (inp[0]) ? node288 : node285;
										assign node285 = (inp[8]) ? 3'b010 : 3'b110;
										assign node288 = (inp[8]) ? 3'b110 : 3'b010;
									assign node291 = (inp[8]) ? node297 : node292;
										assign node292 = (inp[0]) ? node294 : 3'b010;
											assign node294 = (inp[1]) ? 3'b100 : 3'b010;
										assign node297 = (inp[1]) ? 3'b000 : 3'b100;
					assign node302 = (inp[4]) ? node360 : node303;
						assign node303 = (inp[7]) ? node339 : node304;
							assign node304 = (inp[11]) ? node320 : node305;
								assign node305 = (inp[8]) ? node315 : node306;
									assign node306 = (inp[0]) ? node310 : node307;
										assign node307 = (inp[5]) ? 3'b110 : 3'b010;
										assign node310 = (inp[5]) ? node312 : 3'b110;
											assign node312 = (inp[1]) ? 3'b010 : 3'b110;
									assign node315 = (inp[5]) ? 3'b000 : node316;
										assign node316 = (inp[2]) ? 3'b010 : 3'b110;
								assign node320 = (inp[2]) ? node330 : node321;
									assign node321 = (inp[5]) ? node325 : node322;
										assign node322 = (inp[0]) ? 3'b011 : 3'b001;
										assign node325 = (inp[8]) ? 3'b110 : node326;
											assign node326 = (inp[1]) ? 3'b100 : 3'b001;
									assign node330 = (inp[1]) ? 3'b110 : node331;
										assign node331 = (inp[8]) ? node335 : node332;
											assign node332 = (inp[5]) ? 3'b011 : 3'b111;
											assign node335 = (inp[0]) ? 3'b110 : 3'b101;
							assign node339 = (inp[11]) ? node343 : node340;
								assign node340 = (inp[8]) ? 3'b000 : 3'b100;
								assign node343 = (inp[5]) ? node351 : node344;
									assign node344 = (inp[2]) ? 3'b110 : node345;
										assign node345 = (inp[0]) ? 3'b010 : node346;
											assign node346 = (inp[8]) ? 3'b010 : 3'b110;
									assign node351 = (inp[8]) ? node357 : node352;
										assign node352 = (inp[1]) ? node354 : 3'b010;
											assign node354 = (inp[0]) ? 3'b100 : 3'b010;
										assign node357 = (inp[1]) ? 3'b000 : 3'b100;
						assign node360 = (inp[7]) ? 3'b000 : node361;
							assign node361 = (inp[11]) ? node369 : node362;
								assign node362 = (inp[8]) ? 3'b000 : node363;
									assign node363 = (inp[1]) ? node365 : 3'b100;
										assign node365 = (inp[5]) ? 3'b000 : 3'b100;
								assign node369 = (inp[8]) ? node375 : node370;
									assign node370 = (inp[5]) ? 3'b010 : node371;
										assign node371 = (inp[0]) ? 3'b010 : 3'b110;
									assign node375 = (inp[5]) ? 3'b100 : node376;
										assign node376 = (inp[2]) ? 3'b110 : 3'b010;
				assign node381 = (inp[4]) ? node457 : node382;
					assign node382 = (inp[7]) ? node402 : node383;
						assign node383 = (inp[10]) ? 3'b011 : node384;
							assign node384 = (inp[5]) ? node396 : node385;
								assign node385 = (inp[11]) ? node387 : 3'b001;
									assign node387 = (inp[8]) ? node391 : node388;
										assign node388 = (inp[2]) ? 3'b011 : 3'b001;
										assign node391 = (inp[0]) ? node393 : 3'b011;
											assign node393 = (inp[2]) ? 3'b001 : 3'b011;
								assign node396 = (inp[11]) ? node398 : 3'b011;
									assign node398 = (inp[2]) ? 3'b001 : 3'b011;
						assign node402 = (inp[10]) ? node440 : node403;
							assign node403 = (inp[11]) ? node413 : node404;
								assign node404 = (inp[5]) ? node410 : node405;
									assign node405 = (inp[2]) ? node407 : 3'b110;
										assign node407 = (inp[8]) ? 3'b010 : 3'b110;
									assign node410 = (inp[8]) ? 3'b000 : 3'b110;
								assign node413 = (inp[5]) ? node427 : node414;
									assign node414 = (inp[0]) ? node418 : node415;
										assign node415 = (inp[8]) ? 3'b001 : 3'b111;
										assign node418 = (inp[8]) ? node422 : node419;
											assign node419 = (inp[2]) ? 3'b001 : 3'b011;
											assign node422 = (inp[2]) ? node424 : 3'b001;
												assign node424 = (inp[1]) ? 3'b110 : 3'b101;
									assign node427 = (inp[8]) ? node437 : node428;
										assign node428 = (inp[2]) ? node432 : node429;
											assign node429 = (inp[1]) ? 3'b100 : 3'b001;
											assign node432 = (inp[0]) ? node434 : 3'b011;
												assign node434 = (inp[1]) ? 3'b110 : 3'b011;
										assign node437 = (inp[1]) ? 3'b010 : 3'b110;
							assign node440 = (inp[5]) ? node448 : node441;
								assign node441 = (inp[11]) ? node443 : 3'b001;
									assign node443 = (inp[1]) ? node445 : 3'b011;
										assign node445 = (inp[8]) ? 3'b101 : 3'b011;
								assign node448 = (inp[11]) ? node452 : node449;
									assign node449 = (inp[8]) ? 3'b110 : 3'b111;
									assign node452 = (inp[8]) ? node454 : 3'b101;
										assign node454 = (inp[1]) ? 3'b001 : 3'b101;
					assign node457 = (inp[10]) ? node493 : node458;
						assign node458 = (inp[7]) ? node474 : node459;
							assign node459 = (inp[8]) ? node463 : node460;
								assign node460 = (inp[11]) ? 3'b110 : 3'b010;
								assign node463 = (inp[11]) ? node465 : 3'b100;
									assign node465 = (inp[1]) ? 3'b010 : node466;
										assign node466 = (inp[5]) ? node468 : 3'b110;
											assign node468 = (inp[0]) ? 3'b110 : node469;
												assign node469 = (inp[2]) ? 3'b110 : 3'b101;
							assign node474 = (inp[5]) ? node482 : node475;
								assign node475 = (inp[8]) ? node477 : 3'b010;
									assign node477 = (inp[11]) ? node479 : 3'b010;
										assign node479 = (inp[0]) ? 3'b100 : 3'b110;
								assign node482 = (inp[11]) ? node484 : 3'b000;
									assign node484 = (inp[1]) ? node486 : 3'b000;
										assign node486 = (inp[0]) ? node490 : node487;
											assign node487 = (inp[8]) ? 3'b100 : 3'b000;
											assign node490 = (inp[8]) ? 3'b000 : 3'b100;
						assign node493 = (inp[7]) ? node521 : node494;
							assign node494 = (inp[8]) ? node508 : node495;
								assign node495 = (inp[11]) ? node503 : node496;
									assign node496 = (inp[1]) ? node498 : 3'b101;
										assign node498 = (inp[2]) ? 3'b001 : node499;
											assign node499 = (inp[5]) ? 3'b001 : 3'b101;
									assign node503 = (inp[0]) ? node505 : 3'b011;
										assign node505 = (inp[5]) ? 3'b101 : 3'b011;
								assign node508 = (inp[11]) ? node516 : node509;
									assign node509 = (inp[1]) ? 3'b110 : node510;
										assign node510 = (inp[0]) ? node512 : 3'b001;
											assign node512 = (inp[2]) ? 3'b001 : 3'b110;
									assign node516 = (inp[5]) ? node518 : 3'b101;
										assign node518 = (inp[0]) ? 3'b001 : 3'b101;
							assign node521 = (inp[11]) ? node539 : node522;
								assign node522 = (inp[8]) ? node528 : node523;
									assign node523 = (inp[0]) ? node525 : 3'b110;
										assign node525 = (inp[5]) ? 3'b010 : 3'b110;
									assign node528 = (inp[2]) ? node530 : 3'b010;
										assign node530 = (inp[0]) ? node534 : node531;
											assign node531 = (inp[5]) ? 3'b010 : 3'b110;
											assign node534 = (inp[1]) ? node536 : 3'b010;
												assign node536 = (inp[5]) ? 3'b100 : 3'b010;
								assign node539 = (inp[5]) ? node545 : node540;
									assign node540 = (inp[0]) ? node542 : 3'b001;
										assign node542 = (inp[8]) ? 3'b110 : 3'b001;
									assign node545 = (inp[8]) ? 3'b110 : node546;
										assign node546 = (inp[1]) ? 3'b110 : 3'b101;
		assign node550 = (inp[9]) ? node668 : node551;
			assign node551 = (inp[6]) ? 3'b000 : node552;
				assign node552 = (inp[4]) ? node656 : node553;
					assign node553 = (inp[7]) ? node615 : node554;
						assign node554 = (inp[10]) ? node576 : node555;
							assign node555 = (inp[11]) ? node559 : node556;
								assign node556 = (inp[8]) ? 3'b000 : 3'b100;
								assign node559 = (inp[8]) ? node569 : node560;
									assign node560 = (inp[1]) ? node562 : 3'b010;
										assign node562 = (inp[5]) ? node566 : node563;
											assign node563 = (inp[0]) ? 3'b010 : 3'b110;
											assign node566 = (inp[0]) ? 3'b100 : 3'b010;
									assign node569 = (inp[5]) ? 3'b100 : node570;
										assign node570 = (inp[2]) ? node572 : 3'b010;
											assign node572 = (inp[1]) ? 3'b100 : 3'b110;
							assign node576 = (inp[11]) ? node596 : node577;
								assign node577 = (inp[5]) ? node587 : node578;
									assign node578 = (inp[0]) ? node582 : node579;
										assign node579 = (inp[8]) ? 3'b110 : 3'b010;
										assign node582 = (inp[8]) ? node584 : 3'b110;
											assign node584 = (inp[2]) ? 3'b010 : 3'b110;
									assign node587 = (inp[8]) ? node593 : node588;
										assign node588 = (inp[0]) ? node590 : 3'b110;
											assign node590 = (inp[2]) ? 3'b010 : 3'b110;
										assign node593 = (inp[2]) ? 3'b100 : 3'b000;
								assign node596 = (inp[5]) ? node608 : node597;
									assign node597 = (inp[0]) ? node601 : node598;
										assign node598 = (inp[2]) ? 3'b101 : 3'b111;
										assign node601 = (inp[1]) ? 3'b011 : node602;
											assign node602 = (inp[8]) ? 3'b001 : node603;
												assign node603 = (inp[2]) ? 3'b001 : 3'b011;
									assign node608 = (inp[8]) ? 3'b110 : node609;
										assign node609 = (inp[1]) ? 3'b100 : node610;
											assign node610 = (inp[0]) ? 3'b001 : 3'b011;
						assign node615 = (inp[10]) ? node617 : 3'b000;
							assign node617 = (inp[8]) ? node639 : node618;
								assign node618 = (inp[11]) ? node624 : node619;
									assign node619 = (inp[0]) ? node621 : 3'b100;
										assign node621 = (inp[5]) ? 3'b000 : 3'b100;
									assign node624 = (inp[0]) ? node630 : node625;
										assign node625 = (inp[2]) ? node627 : 3'b000;
											assign node627 = (inp[1]) ? 3'b000 : 3'b010;
										assign node630 = (inp[5]) ? node632 : 3'b000;
											assign node632 = (inp[2]) ? node636 : node633;
												assign node633 = (inp[1]) ? 3'b110 : 3'b000;
												assign node636 = (inp[1]) ? 3'b100 : 3'b110;
								assign node639 = (inp[0]) ? node645 : node640;
									assign node640 = (inp[11]) ? node642 : 3'b000;
										assign node642 = (inp[5]) ? 3'b100 : 3'b000;
									assign node645 = (inp[1]) ? node649 : node646;
										assign node646 = (inp[11]) ? 3'b100 : 3'b000;
										assign node649 = (inp[11]) ? node653 : node650;
											assign node650 = (inp[5]) ? 3'b100 : 3'b000;
											assign node653 = (inp[5]) ? 3'b000 : 3'b100;
					assign node656 = (inp[10]) ? node658 : 3'b000;
						assign node658 = (inp[11]) ? node660 : 3'b000;
							assign node660 = (inp[7]) ? 3'b000 : node661;
								assign node661 = (inp[5]) ? node663 : 3'b100;
									assign node663 = (inp[8]) ? 3'b000 : 3'b100;
			assign node668 = (inp[6]) ? node866 : node669;
				assign node669 = (inp[4]) ? node777 : node670;
					assign node670 = (inp[7]) ? node694 : node671;
						assign node671 = (inp[10]) ? 3'b111 : node672;
							assign node672 = (inp[2]) ? node682 : node673;
								assign node673 = (inp[5]) ? node677 : node674;
									assign node674 = (inp[8]) ? 3'b011 : 3'b101;
									assign node677 = (inp[8]) ? node679 : 3'b011;
										assign node679 = (inp[11]) ? 3'b101 : 3'b011;
								assign node682 = (inp[11]) ? node686 : node683;
									assign node683 = (inp[5]) ? 3'b011 : 3'b101;
									assign node686 = (inp[5]) ? 3'b101 : node687;
										assign node687 = (inp[0]) ? node689 : 3'b011;
											assign node689 = (inp[8]) ? 3'b101 : 3'b011;
						assign node694 = (inp[10]) ? node728 : node695;
							assign node695 = (inp[11]) ? node711 : node696;
								assign node696 = (inp[5]) ? node704 : node697;
									assign node697 = (inp[0]) ? 3'b110 : node698;
										assign node698 = (inp[2]) ? 3'b010 : node699;
											assign node699 = (inp[8]) ? 3'b110 : 3'b010;
									assign node704 = (inp[8]) ? node708 : node705;
										assign node705 = (inp[1]) ? 3'b010 : 3'b110;
										assign node708 = (inp[1]) ? 3'b100 : 3'b000;
								assign node711 = (inp[5]) ? node721 : node712;
									assign node712 = (inp[8]) ? node718 : node713;
										assign node713 = (inp[0]) ? node715 : 3'b111;
											assign node715 = (inp[2]) ? 3'b001 : 3'b011;
										assign node718 = (inp[2]) ? 3'b101 : 3'b001;
									assign node721 = (inp[8]) ? node725 : node722;
										assign node722 = (inp[2]) ? 3'b011 : 3'b001;
										assign node725 = (inp[2]) ? 3'b010 : 3'b110;
							assign node728 = (inp[8]) ? node758 : node729;
								assign node729 = (inp[1]) ? node739 : node730;
									assign node730 = (inp[0]) ? node736 : node731;
										assign node731 = (inp[11]) ? 3'b101 : node732;
											assign node732 = (inp[5]) ? 3'b101 : 3'b001;
										assign node736 = (inp[11]) ? 3'b001 : 3'b101;
									assign node739 = (inp[11]) ? node751 : node740;
										assign node740 = (inp[2]) ? node746 : node741;
											assign node741 = (inp[5]) ? node743 : 3'b001;
												assign node743 = (inp[0]) ? 3'b001 : 3'b101;
											assign node746 = (inp[0]) ? node748 : 3'b001;
												assign node748 = (inp[5]) ? 3'b001 : 3'b101;
										assign node751 = (inp[5]) ? node755 : node752;
											assign node752 = (inp[0]) ? 3'b001 : 3'b101;
											assign node755 = (inp[0]) ? 3'b111 : 3'b011;
								assign node758 = (inp[11]) ? node764 : node759;
									assign node759 = (inp[5]) ? 3'b010 : node760;
										assign node760 = (inp[2]) ? 3'b001 : 3'b101;
									assign node764 = (inp[5]) ? node772 : node765;
										assign node765 = (inp[2]) ? node767 : 3'b011;
											assign node767 = (inp[0]) ? node769 : 3'b111;
												assign node769 = (inp[1]) ? 3'b101 : 3'b111;
										assign node772 = (inp[0]) ? node774 : 3'b101;
											assign node774 = (inp[1]) ? 3'b001 : 3'b101;
					assign node777 = (inp[10]) ? node819 : node778;
						assign node778 = (inp[7]) ? node796 : node779;
							assign node779 = (inp[8]) ? node789 : node780;
								assign node780 = (inp[11]) ? node782 : 3'b010;
									assign node782 = (inp[1]) ? 3'b110 : node783;
										assign node783 = (inp[2]) ? 3'b110 : node784;
											assign node784 = (inp[0]) ? 3'b110 : 3'b001;
								assign node789 = (inp[11]) ? node791 : 3'b100;
									assign node791 = (inp[1]) ? 3'b010 : node792;
										assign node792 = (inp[0]) ? 3'b110 : 3'b101;
							assign node796 = (inp[11]) ? node806 : node797;
								assign node797 = (inp[5]) ? 3'b000 : node798;
									assign node798 = (inp[0]) ? node800 : 3'b100;
										assign node800 = (inp[1]) ? node802 : 3'b100;
											assign node802 = (inp[8]) ? 3'b000 : 3'b100;
								assign node806 = (inp[8]) ? node814 : node807;
									assign node807 = (inp[5]) ? node809 : 3'b010;
										assign node809 = (inp[1]) ? 3'b100 : node810;
											assign node810 = (inp[2]) ? 3'b010 : 3'b100;
									assign node814 = (inp[1]) ? 3'b100 : node815;
										assign node815 = (inp[2]) ? 3'b100 : 3'b000;
						assign node819 = (inp[7]) ? node847 : node820;
							assign node820 = (inp[8]) ? node832 : node821;
								assign node821 = (inp[11]) ? node827 : node822;
									assign node822 = (inp[0]) ? node824 : 3'b101;
										assign node824 = (inp[1]) ? 3'b001 : 3'b101;
									assign node827 = (inp[0]) ? node829 : 3'b011;
										assign node829 = (inp[5]) ? 3'b101 : 3'b011;
								assign node832 = (inp[11]) ? node842 : node833;
									assign node833 = (inp[1]) ? node839 : node834;
										assign node834 = (inp[0]) ? node836 : 3'b001;
											assign node836 = (inp[2]) ? 3'b001 : 3'b110;
										assign node839 = (inp[2]) ? 3'b110 : 3'b001;
									assign node842 = (inp[5]) ? node844 : 3'b101;
										assign node844 = (inp[0]) ? 3'b001 : 3'b101;
							assign node847 = (inp[11]) ? node855 : node848;
								assign node848 = (inp[8]) ? 3'b010 : node849;
									assign node849 = (inp[0]) ? node851 : 3'b110;
										assign node851 = (inp[5]) ? 3'b010 : 3'b110;
								assign node855 = (inp[8]) ? node863 : node856;
									assign node856 = (inp[0]) ? node858 : 3'b001;
										assign node858 = (inp[2]) ? 3'b001 : node859;
											assign node859 = (inp[1]) ? 3'b110 : 3'b001;
									assign node863 = (inp[5]) ? 3'b110 : 3'b101;
				assign node866 = (inp[7]) ? node950 : node867;
					assign node867 = (inp[11]) ? node901 : node868;
						assign node868 = (inp[8]) ? node894 : node869;
							assign node869 = (inp[4]) ? node887 : node870;
								assign node870 = (inp[10]) ? node878 : node871;
									assign node871 = (inp[0]) ? node873 : 3'b100;
										assign node873 = (inp[1]) ? 3'b000 : node874;
											assign node874 = (inp[2]) ? 3'b000 : 3'b100;
									assign node878 = (inp[1]) ? node880 : 3'b110;
										assign node880 = (inp[0]) ? node884 : node881;
											assign node881 = (inp[5]) ? 3'b110 : 3'b010;
											assign node884 = (inp[5]) ? 3'b010 : 3'b110;
								assign node887 = (inp[10]) ? node889 : 3'b000;
									assign node889 = (inp[5]) ? node891 : 3'b100;
										assign node891 = (inp[0]) ? 3'b000 : 3'b100;
							assign node894 = (inp[5]) ? 3'b000 : node895;
								assign node895 = (inp[10]) ? node897 : 3'b000;
									assign node897 = (inp[4]) ? 3'b000 : 3'b110;
						assign node901 = (inp[4]) ? node929 : node902;
							assign node902 = (inp[10]) ? node916 : node903;
								assign node903 = (inp[5]) ? node909 : node904;
									assign node904 = (inp[2]) ? 3'b110 : node905;
										assign node905 = (inp[8]) ? 3'b010 : 3'b110;
									assign node909 = (inp[8]) ? 3'b100 : node910;
										assign node910 = (inp[0]) ? node912 : 3'b010;
											assign node912 = (inp[1]) ? 3'b100 : 3'b010;
								assign node916 = (inp[5]) ? node922 : node917;
									assign node917 = (inp[2]) ? node919 : 3'b001;
										assign node919 = (inp[8]) ? 3'b101 : 3'b111;
									assign node922 = (inp[8]) ? node924 : 3'b011;
										assign node924 = (inp[2]) ? node926 : 3'b110;
											assign node926 = (inp[0]) ? 3'b010 : 3'b110;
							assign node929 = (inp[10]) ? node931 : 3'b000;
								assign node931 = (inp[0]) ? node939 : node932;
									assign node932 = (inp[5]) ? 3'b010 : node933;
										assign node933 = (inp[8]) ? node935 : 3'b110;
											assign node935 = (inp[2]) ? 3'b110 : 3'b010;
									assign node939 = (inp[8]) ? node945 : node940;
										assign node940 = (inp[1]) ? node942 : 3'b010;
											assign node942 = (inp[5]) ? 3'b100 : 3'b010;
										assign node945 = (inp[1]) ? 3'b100 : node946;
											assign node946 = (inp[2]) ? 3'b100 : 3'b010;
					assign node950 = (inp[10]) ? node952 : 3'b000;
						assign node952 = (inp[4]) ? node978 : node953;
							assign node953 = (inp[11]) ? node961 : node954;
								assign node954 = (inp[5]) ? 3'b000 : node955;
									assign node955 = (inp[0]) ? node957 : 3'b100;
										assign node957 = (inp[2]) ? 3'b100 : 3'b000;
								assign node961 = (inp[5]) ? node973 : node962;
									assign node962 = (inp[0]) ? node964 : 3'b010;
										assign node964 = (inp[1]) ? node968 : node965;
											assign node965 = (inp[2]) ? 3'b010 : 3'b110;
											assign node968 = (inp[8]) ? node970 : 3'b010;
												assign node970 = (inp[2]) ? 3'b100 : 3'b010;
									assign node973 = (inp[8]) ? 3'b100 : node974;
										assign node974 = (inp[2]) ? 3'b110 : 3'b010;
							assign node978 = (inp[8]) ? 3'b000 : node979;
								assign node979 = (inp[5]) ? 3'b000 : node980;
									assign node980 = (inp[11]) ? node982 : 3'b000;
										assign node982 = (inp[2]) ? 3'b000 : 3'b100;

endmodule