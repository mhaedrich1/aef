module dtc_split75_bm70 (
	input  wire [12-1:0] inp,
	output wire [3-1:0] outp
);

	wire [3-1:0] node1;
	wire [3-1:0] node2;
	wire [3-1:0] node3;
	wire [3-1:0] node4;
	wire [3-1:0] node5;
	wire [3-1:0] node8;
	wire [3-1:0] node11;
	wire [3-1:0] node12;
	wire [3-1:0] node15;
	wire [3-1:0] node18;
	wire [3-1:0] node19;
	wire [3-1:0] node20;
	wire [3-1:0] node23;
	wire [3-1:0] node26;
	wire [3-1:0] node27;
	wire [3-1:0] node30;
	wire [3-1:0] node33;
	wire [3-1:0] node34;
	wire [3-1:0] node35;
	wire [3-1:0] node36;
	wire [3-1:0] node39;
	wire [3-1:0] node42;
	wire [3-1:0] node43;
	wire [3-1:0] node46;
	wire [3-1:0] node49;
	wire [3-1:0] node50;
	wire [3-1:0] node51;
	wire [3-1:0] node54;
	wire [3-1:0] node57;
	wire [3-1:0] node58;
	wire [3-1:0] node61;
	wire [3-1:0] node64;
	wire [3-1:0] node65;
	wire [3-1:0] node66;
	wire [3-1:0] node68;
	wire [3-1:0] node69;
	wire [3-1:0] node72;
	wire [3-1:0] node76;
	wire [3-1:0] node77;
	wire [3-1:0] node78;
	wire [3-1:0] node79;
	wire [3-1:0] node82;
	wire [3-1:0] node85;
	wire [3-1:0] node86;
	wire [3-1:0] node89;
	wire [3-1:0] node92;
	wire [3-1:0] node93;
	wire [3-1:0] node95;
	wire [3-1:0] node98;
	wire [3-1:0] node99;
	wire [3-1:0] node102;

	assign outp = (inp[3]) ? node64 : node1;
		assign node1 = (inp[0]) ? node33 : node2;
			assign node2 = (inp[4]) ? node18 : node3;
				assign node3 = (inp[1]) ? node11 : node4;
					assign node4 = (inp[9]) ? node8 : node5;
						assign node5 = (inp[6]) ? 3'b010 : 3'b000;
						assign node8 = (inp[6]) ? 3'b111 : 3'b010;
					assign node11 = (inp[9]) ? node15 : node12;
						assign node12 = (inp[6]) ? 3'b001 : 3'b110;
						assign node15 = (inp[6]) ? 3'b111 : 3'b111;
				assign node18 = (inp[1]) ? node26 : node19;
					assign node19 = (inp[9]) ? node23 : node20;
						assign node20 = (inp[8]) ? 3'b000 : 3'b000;
						assign node23 = (inp[6]) ? 3'b000 : 3'b000;
					assign node26 = (inp[9]) ? node30 : node27;
						assign node27 = (inp[6]) ? 3'b000 : 3'b000;
						assign node30 = (inp[6]) ? 3'b010 : 3'b000;
			assign node33 = (inp[4]) ? node49 : node34;
				assign node34 = (inp[6]) ? node42 : node35;
					assign node35 = (inp[9]) ? node39 : node36;
						assign node36 = (inp[1]) ? 3'b111 : 3'b011;
						assign node39 = (inp[1]) ? 3'b111 : 3'b111;
					assign node42 = (inp[9]) ? node46 : node43;
						assign node43 = (inp[1]) ? 3'b111 : 3'b111;
						assign node46 = (inp[5]) ? 3'b111 : 3'b111;
				assign node49 = (inp[9]) ? node57 : node50;
					assign node50 = (inp[6]) ? node54 : node51;
						assign node51 = (inp[1]) ? 3'b110 : 3'b000;
						assign node54 = (inp[1]) ? 3'b011 : 3'b010;
					assign node57 = (inp[6]) ? node61 : node58;
						assign node58 = (inp[1]) ? 3'b111 : 3'b110;
						assign node61 = (inp[1]) ? 3'b111 : 3'b111;
		assign node64 = (inp[0]) ? node76 : node65;
			assign node65 = (inp[4]) ? 3'b000 : node66;
				assign node66 = (inp[9]) ? node68 : 3'b000;
					assign node68 = (inp[6]) ? node72 : node69;
						assign node69 = (inp[11]) ? 3'b000 : 3'b000;
						assign node72 = (inp[5]) ? 3'b000 : 3'b000;
			assign node76 = (inp[4]) ? node92 : node77;
				assign node77 = (inp[9]) ? node85 : node78;
					assign node78 = (inp[1]) ? node82 : node79;
						assign node79 = (inp[6]) ? 3'b000 : 3'b000;
						assign node82 = (inp[6]) ? 3'b010 : 3'b000;
					assign node85 = (inp[1]) ? node89 : node86;
						assign node86 = (inp[6]) ? 3'b010 : 3'b000;
						assign node89 = (inp[6]) ? 3'b011 : 3'b010;
				assign node92 = (inp[9]) ? node98 : node93;
					assign node93 = (inp[1]) ? node95 : 3'b000;
						assign node95 = (inp[8]) ? 3'b000 : 3'b000;
					assign node98 = (inp[1]) ? node102 : node99;
						assign node99 = (inp[6]) ? 3'b000 : 3'b000;
						assign node102 = (inp[6]) ? 3'b000 : 3'b000;

endmodule