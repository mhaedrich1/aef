module dtc_split25_bm78 (
	input  wire [12-1:0] inp,
	output wire [3-1:0] outp
);

	wire [3-1:0] node1;
	wire [3-1:0] node2;
	wire [3-1:0] node3;
	wire [3-1:0] node4;
	wire [3-1:0] node5;
	wire [3-1:0] node6;
	wire [3-1:0] node7;
	wire [3-1:0] node8;
	wire [3-1:0] node10;
	wire [3-1:0] node13;
	wire [3-1:0] node15;
	wire [3-1:0] node18;
	wire [3-1:0] node19;
	wire [3-1:0] node22;
	wire [3-1:0] node25;
	wire [3-1:0] node26;
	wire [3-1:0] node27;
	wire [3-1:0] node28;
	wire [3-1:0] node32;
	wire [3-1:0] node35;
	wire [3-1:0] node36;
	wire [3-1:0] node37;
	wire [3-1:0] node40;
	wire [3-1:0] node43;
	wire [3-1:0] node44;
	wire [3-1:0] node48;
	wire [3-1:0] node49;
	wire [3-1:0] node50;
	wire [3-1:0] node51;
	wire [3-1:0] node53;
	wire [3-1:0] node56;
	wire [3-1:0] node58;
	wire [3-1:0] node61;
	wire [3-1:0] node62;
	wire [3-1:0] node63;
	wire [3-1:0] node67;
	wire [3-1:0] node68;
	wire [3-1:0] node72;
	wire [3-1:0] node73;
	wire [3-1:0] node75;
	wire [3-1:0] node76;
	wire [3-1:0] node80;
	wire [3-1:0] node82;
	wire [3-1:0] node83;
	wire [3-1:0] node86;
	wire [3-1:0] node89;
	wire [3-1:0] node90;
	wire [3-1:0] node92;
	wire [3-1:0] node93;
	wire [3-1:0] node94;
	wire [3-1:0] node95;
	wire [3-1:0] node99;
	wire [3-1:0] node102;
	wire [3-1:0] node104;
	wire [3-1:0] node105;
	wire [3-1:0] node109;
	wire [3-1:0] node110;
	wire [3-1:0] node111;
	wire [3-1:0] node112;
	wire [3-1:0] node117;
	wire [3-1:0] node118;
	wire [3-1:0] node119;
	wire [3-1:0] node120;
	wire [3-1:0] node123;
	wire [3-1:0] node126;
	wire [3-1:0] node127;
	wire [3-1:0] node131;
	wire [3-1:0] node132;
	wire [3-1:0] node135;
	wire [3-1:0] node136;
	wire [3-1:0] node140;
	wire [3-1:0] node141;
	wire [3-1:0] node142;
	wire [3-1:0] node143;
	wire [3-1:0] node144;
	wire [3-1:0] node145;
	wire [3-1:0] node146;
	wire [3-1:0] node149;
	wire [3-1:0] node152;
	wire [3-1:0] node154;
	wire [3-1:0] node157;
	wire [3-1:0] node159;
	wire [3-1:0] node160;
	wire [3-1:0] node164;
	wire [3-1:0] node165;
	wire [3-1:0] node166;
	wire [3-1:0] node168;
	wire [3-1:0] node171;
	wire [3-1:0] node173;
	wire [3-1:0] node176;
	wire [3-1:0] node177;
	wire [3-1:0] node180;
	wire [3-1:0] node182;
	wire [3-1:0] node185;
	wire [3-1:0] node186;
	wire [3-1:0] node187;
	wire [3-1:0] node188;
	wire [3-1:0] node192;
	wire [3-1:0] node194;
	wire [3-1:0] node199;
	wire [3-1:0] node200;
	wire [3-1:0] node202;
	wire [3-1:0] node203;
	wire [3-1:0] node204;
	wire [3-1:0] node206;
	wire [3-1:0] node207;
	wire [3-1:0] node211;
	wire [3-1:0] node212;
	wire [3-1:0] node214;
	wire [3-1:0] node217;
	wire [3-1:0] node218;
	wire [3-1:0] node220;
	wire [3-1:0] node224;
	wire [3-1:0] node225;
	wire [3-1:0] node227;
	wire [3-1:0] node228;
	wire [3-1:0] node232;
	wire [3-1:0] node234;
	wire [3-1:0] node236;
	wire [3-1:0] node238;
	wire [3-1:0] node241;
	wire [3-1:0] node242;
	wire [3-1:0] node243;
	wire [3-1:0] node244;
	wire [3-1:0] node245;
	wire [3-1:0] node246;
	wire [3-1:0] node247;
	wire [3-1:0] node251;
	wire [3-1:0] node252;
	wire [3-1:0] node256;
	wire [3-1:0] node257;
	wire [3-1:0] node259;
	wire [3-1:0] node262;
	wire [3-1:0] node263;
	wire [3-1:0] node267;
	wire [3-1:0] node269;
	wire [3-1:0] node273;
	wire [3-1:0] node274;
	wire [3-1:0] node275;
	wire [3-1:0] node276;
	wire [3-1:0] node277;
	wire [3-1:0] node278;
	wire [3-1:0] node281;
	wire [3-1:0] node286;
	wire [3-1:0] node287;
	wire [3-1:0] node288;
	wire [3-1:0] node289;
	wire [3-1:0] node293;
	wire [3-1:0] node295;
	wire [3-1:0] node298;
	wire [3-1:0] node299;
	wire [3-1:0] node300;
	wire [3-1:0] node303;
	wire [3-1:0] node307;
	wire [3-1:0] node308;
	wire [3-1:0] node312;
	wire [3-1:0] node313;
	wire [3-1:0] node315;
	wire [3-1:0] node316;
	wire [3-1:0] node317;
	wire [3-1:0] node319;
	wire [3-1:0] node321;
	wire [3-1:0] node326;
	wire [3-1:0] node327;
	wire [3-1:0] node328;
	wire [3-1:0] node329;
	wire [3-1:0] node330;
	wire [3-1:0] node332;
	wire [3-1:0] node334;
	wire [3-1:0] node339;
	wire [3-1:0] node340;
	wire [3-1:0] node341;
	wire [3-1:0] node342;
	wire [3-1:0] node343;
	wire [3-1:0] node345;
	wire [3-1:0] node348;
	wire [3-1:0] node351;
	wire [3-1:0] node352;
	wire [3-1:0] node355;
	wire [3-1:0] node356;
	wire [3-1:0] node359;
	wire [3-1:0] node362;
	wire [3-1:0] node363;
	wire [3-1:0] node365;
	wire [3-1:0] node367;
	wire [3-1:0] node370;
	wire [3-1:0] node371;
	wire [3-1:0] node373;
	wire [3-1:0] node376;
	wire [3-1:0] node379;
	wire [3-1:0] node380;
	wire [3-1:0] node381;
	wire [3-1:0] node382;
	wire [3-1:0] node383;
	wire [3-1:0] node387;
	wire [3-1:0] node388;
	wire [3-1:0] node392;
	wire [3-1:0] node393;
	wire [3-1:0] node395;
	wire [3-1:0] node399;
	wire [3-1:0] node401;
	wire [3-1:0] node402;
	wire [3-1:0] node404;
	wire [3-1:0] node408;
	wire [3-1:0] node410;
	wire [3-1:0] node412;
	wire [3-1:0] node413;
	wire [3-1:0] node414;
	wire [3-1:0] node415;
	wire [3-1:0] node417;
	wire [3-1:0] node420;
	wire [3-1:0] node421;
	wire [3-1:0] node425;
	wire [3-1:0] node428;
	wire [3-1:0] node429;
	wire [3-1:0] node431;
	wire [3-1:0] node433;
	wire [3-1:0] node436;

	assign outp = (inp[3]) ? node312 : node1;
		assign node1 = (inp[4]) ? node199 : node2;
			assign node2 = (inp[0]) ? node140 : node3;
				assign node3 = (inp[6]) ? node89 : node4;
					assign node4 = (inp[5]) ? node48 : node5;
						assign node5 = (inp[9]) ? node25 : node6;
							assign node6 = (inp[1]) ? node18 : node7;
								assign node7 = (inp[7]) ? node13 : node8;
									assign node8 = (inp[11]) ? node10 : 3'b000;
										assign node10 = (inp[10]) ? 3'b100 : 3'b000;
									assign node13 = (inp[2]) ? node15 : 3'b100;
										assign node15 = (inp[11]) ? 3'b010 : 3'b100;
								assign node18 = (inp[2]) ? node22 : node19;
									assign node19 = (inp[8]) ? 3'b011 : 3'b010;
									assign node22 = (inp[7]) ? 3'b101 : 3'b110;
							assign node25 = (inp[1]) ? node35 : node26;
								assign node26 = (inp[2]) ? node32 : node27;
									assign node27 = (inp[8]) ? 3'b011 : node28;
										assign node28 = (inp[10]) ? 3'b110 : 3'b010;
									assign node32 = (inp[10]) ? 3'b001 : 3'b111;
								assign node35 = (inp[10]) ? node43 : node36;
									assign node36 = (inp[8]) ? node40 : node37;
										assign node37 = (inp[2]) ? 3'b001 : 3'b001;
										assign node40 = (inp[11]) ? 3'b001 : 3'b110;
									assign node43 = (inp[2]) ? 3'b011 : node44;
										assign node44 = (inp[8]) ? 3'b011 : 3'b001;
						assign node48 = (inp[1]) ? node72 : node49;
							assign node49 = (inp[10]) ? node61 : node50;
								assign node50 = (inp[7]) ? node56 : node51;
									assign node51 = (inp[11]) ? node53 : 3'b000;
										assign node53 = (inp[2]) ? 3'b100 : 3'b000;
									assign node56 = (inp[8]) ? node58 : 3'b100;
										assign node58 = (inp[9]) ? 3'b000 : 3'b000;
								assign node61 = (inp[9]) ? node67 : node62;
									assign node62 = (inp[7]) ? 3'b000 : node63;
										assign node63 = (inp[11]) ? 3'b100 : 3'b000;
									assign node67 = (inp[2]) ? 3'b010 : node68;
										assign node68 = (inp[7]) ? 3'b110 : 3'b100;
							assign node72 = (inp[10]) ? node80 : node73;
								assign node73 = (inp[9]) ? node75 : 3'b100;
									assign node75 = (inp[8]) ? 3'b100 : node76;
										assign node76 = (inp[11]) ? 3'b010 : 3'b000;
								assign node80 = (inp[9]) ? node82 : 3'b110;
									assign node82 = (inp[2]) ? node86 : node83;
										assign node83 = (inp[8]) ? 3'b001 : 3'b100;
										assign node86 = (inp[8]) ? 3'b011 : 3'b001;
					assign node89 = (inp[9]) ? node109 : node90;
						assign node90 = (inp[5]) ? node92 : 3'b011;
							assign node92 = (inp[8]) ? node102 : node93;
								assign node93 = (inp[1]) ? node99 : node94;
									assign node94 = (inp[7]) ? 3'b010 : node95;
										assign node95 = (inp[10]) ? 3'b010 : 3'b011;
									assign node99 = (inp[7]) ? 3'b011 : 3'b010;
								assign node102 = (inp[11]) ? node104 : 3'b011;
									assign node104 = (inp[2]) ? 3'b011 : node105;
										assign node105 = (inp[1]) ? 3'b011 : 3'b010;
						assign node109 = (inp[2]) ? node117 : node110;
							assign node110 = (inp[7]) ? 3'b011 : node111;
								assign node111 = (inp[10]) ? 3'b101 : node112;
									assign node112 = (inp[11]) ? 3'b011 : 3'b111;
							assign node117 = (inp[1]) ? node131 : node118;
								assign node118 = (inp[11]) ? node126 : node119;
									assign node119 = (inp[5]) ? node123 : node120;
										assign node120 = (inp[10]) ? 3'b111 : 3'b011;
										assign node123 = (inp[7]) ? 3'b111 : 3'b101;
									assign node126 = (inp[8]) ? 3'b011 : node127;
										assign node127 = (inp[7]) ? 3'b111 : 3'b011;
								assign node131 = (inp[7]) ? node135 : node132;
									assign node132 = (inp[5]) ? 3'b101 : 3'b111;
									assign node135 = (inp[11]) ? 3'b111 : node136;
										assign node136 = (inp[10]) ? 3'b011 : 3'b111;
				assign node140 = (inp[6]) ? 3'b111 : node141;
					assign node141 = (inp[1]) ? node185 : node142;
						assign node142 = (inp[9]) ? node164 : node143;
							assign node143 = (inp[10]) ? node157 : node144;
								assign node144 = (inp[7]) ? node152 : node145;
									assign node145 = (inp[11]) ? node149 : node146;
										assign node146 = (inp[8]) ? 3'b110 : 3'b010;
										assign node149 = (inp[8]) ? 3'b110 : 3'b101;
									assign node152 = (inp[11]) ? node154 : 3'b101;
										assign node154 = (inp[8]) ? 3'b011 : 3'b001;
								assign node157 = (inp[2]) ? node159 : 3'b001;
									assign node159 = (inp[5]) ? 3'b101 : node160;
										assign node160 = (inp[7]) ? 3'b111 : 3'b101;
							assign node164 = (inp[11]) ? node176 : node165;
								assign node165 = (inp[7]) ? node171 : node166;
									assign node166 = (inp[2]) ? node168 : 3'b101;
										assign node168 = (inp[8]) ? 3'b101 : 3'b011;
									assign node171 = (inp[5]) ? node173 : 3'b111;
										assign node173 = (inp[10]) ? 3'b011 : 3'b001;
								assign node176 = (inp[10]) ? node180 : node177;
									assign node177 = (inp[7]) ? 3'b101 : 3'b011;
									assign node180 = (inp[5]) ? node182 : 3'b111;
										assign node182 = (inp[8]) ? 3'b111 : 3'b011;
						assign node185 = (inp[9]) ? 3'b111 : node186;
							assign node186 = (inp[7]) ? node192 : node187;
								assign node187 = (inp[5]) ? 3'b101 : node188;
									assign node188 = (inp[10]) ? 3'b111 : 3'b011;
								assign node192 = (inp[2]) ? node194 : 3'b111;
									assign node194 = (inp[11]) ? 3'b111 : 3'b011;
			assign node199 = (inp[0]) ? node241 : node200;
				assign node200 = (inp[9]) ? node202 : 3'b000;
					assign node202 = (inp[6]) ? node224 : node203;
						assign node203 = (inp[1]) ? node211 : node204;
							assign node204 = (inp[7]) ? node206 : 3'b000;
								assign node206 = (inp[8]) ? 3'b100 : node207;
									assign node207 = (inp[2]) ? 3'b000 : 3'b100;
							assign node211 = (inp[8]) ? node217 : node212;
								assign node212 = (inp[7]) ? node214 : 3'b100;
									assign node214 = (inp[2]) ? 3'b010 : 3'b100;
								assign node217 = (inp[5]) ? 3'b000 : node218;
									assign node218 = (inp[7]) ? node220 : 3'b010;
										assign node220 = (inp[11]) ? 3'b001 : 3'b010;
						assign node224 = (inp[5]) ? node232 : node225;
							assign node225 = (inp[1]) ? node227 : 3'b000;
								assign node227 = (inp[2]) ? 3'b001 : node228;
									assign node228 = (inp[7]) ? 3'b001 : 3'b000;
							assign node232 = (inp[8]) ? node234 : 3'b000;
								assign node234 = (inp[11]) ? node236 : 3'b000;
									assign node236 = (inp[2]) ? node238 : 3'b000;
										assign node238 = (inp[1]) ? 3'b001 : 3'b000;
				assign node241 = (inp[9]) ? node273 : node242;
					assign node242 = (inp[6]) ? 3'b000 : node243;
						assign node243 = (inp[7]) ? node267 : node244;
							assign node244 = (inp[2]) ? node256 : node245;
								assign node245 = (inp[1]) ? node251 : node246;
									assign node246 = (inp[5]) ? 3'b000 : node247;
										assign node247 = (inp[11]) ? 3'b000 : 3'b100;
									assign node251 = (inp[11]) ? 3'b010 : node252;
										assign node252 = (inp[5]) ? 3'b000 : 3'b010;
								assign node256 = (inp[5]) ? node262 : node257;
									assign node257 = (inp[1]) ? node259 : 3'b010;
										assign node259 = (inp[8]) ? 3'b101 : 3'b001;
									assign node262 = (inp[8]) ? 3'b000 : node263;
										assign node263 = (inp[10]) ? 3'b000 : 3'b100;
							assign node267 = (inp[1]) ? node269 : 3'b110;
								assign node269 = (inp[8]) ? 3'b110 : 3'b111;
					assign node273 = (inp[6]) ? node307 : node274;
						assign node274 = (inp[1]) ? node286 : node275;
							assign node275 = (inp[5]) ? 3'b110 : node276;
								assign node276 = (inp[7]) ? 3'b101 : node277;
									assign node277 = (inp[10]) ? node281 : node278;
										assign node278 = (inp[2]) ? 3'b110 : 3'b010;
										assign node281 = (inp[11]) ? 3'b001 : 3'b001;
							assign node286 = (inp[5]) ? node298 : node287;
								assign node287 = (inp[10]) ? node293 : node288;
									assign node288 = (inp[2]) ? 3'b011 : node289;
										assign node289 = (inp[7]) ? 3'b111 : 3'b101;
									assign node293 = (inp[2]) ? node295 : 3'b011;
										assign node295 = (inp[11]) ? 3'b111 : 3'b011;
								assign node298 = (inp[7]) ? 3'b011 : node299;
									assign node299 = (inp[10]) ? node303 : node300;
										assign node300 = (inp[2]) ? 3'b001 : 3'b010;
										assign node303 = (inp[2]) ? 3'b101 : 3'b001;
						assign node307 = (inp[7]) ? 3'b111 : node308;
							assign node308 = (inp[10]) ? 3'b111 : 3'b011;
		assign node312 = (inp[0]) ? node326 : node313;
			assign node313 = (inp[11]) ? node315 : 3'b000;
				assign node315 = (inp[6]) ? 3'b000 : node316;
					assign node316 = (inp[4]) ? 3'b000 : node317;
						assign node317 = (inp[8]) ? node319 : 3'b000;
							assign node319 = (inp[9]) ? node321 : 3'b000;
								assign node321 = (inp[7]) ? 3'b100 : 3'b000;
			assign node326 = (inp[4]) ? node408 : node327;
				assign node327 = (inp[9]) ? node339 : node328;
					assign node328 = (inp[6]) ? 3'b000 : node329;
						assign node329 = (inp[7]) ? 3'b100 : node330;
							assign node330 = (inp[1]) ? node332 : 3'b000;
								assign node332 = (inp[10]) ? node334 : 3'b000;
									assign node334 = (inp[5]) ? 3'b000 : 3'b100;
					assign node339 = (inp[6]) ? node379 : node340;
						assign node340 = (inp[5]) ? node362 : node341;
							assign node341 = (inp[10]) ? node351 : node342;
								assign node342 = (inp[2]) ? node348 : node343;
									assign node343 = (inp[8]) ? node345 : 3'b100;
										assign node345 = (inp[7]) ? 3'b000 : 3'b000;
									assign node348 = (inp[8]) ? 3'b001 : 3'b010;
								assign node351 = (inp[11]) ? node355 : node352;
									assign node352 = (inp[2]) ? 3'b101 : 3'b011;
									assign node355 = (inp[2]) ? node359 : node356;
										assign node356 = (inp[1]) ? 3'b010 : 3'b100;
										assign node359 = (inp[1]) ? 3'b100 : 3'b010;
							assign node362 = (inp[1]) ? node370 : node363;
								assign node363 = (inp[8]) ? node365 : 3'b000;
									assign node365 = (inp[7]) ? node367 : 3'b000;
										assign node367 = (inp[10]) ? 3'b100 : 3'b000;
								assign node370 = (inp[11]) ? node376 : node371;
									assign node371 = (inp[8]) ? node373 : 3'b000;
										assign node373 = (inp[2]) ? 3'b000 : 3'b100;
									assign node376 = (inp[7]) ? 3'b110 : 3'b100;
						assign node379 = (inp[7]) ? node399 : node380;
							assign node380 = (inp[1]) ? node392 : node381;
								assign node381 = (inp[10]) ? node387 : node382;
									assign node382 = (inp[2]) ? 3'b011 : node383;
										assign node383 = (inp[5]) ? 3'b011 : 3'b010;
									assign node387 = (inp[8]) ? 3'b010 : node388;
										assign node388 = (inp[5]) ? 3'b011 : 3'b010;
								assign node392 = (inp[2]) ? 3'b011 : node393;
									assign node393 = (inp[5]) ? node395 : 3'b001;
										assign node395 = (inp[10]) ? 3'b011 : 3'b010;
							assign node399 = (inp[5]) ? node401 : 3'b101;
								assign node401 = (inp[1]) ? 3'b101 : node402;
									assign node402 = (inp[10]) ? node404 : 3'b100;
										assign node404 = (inp[8]) ? 3'b101 : 3'b100;
				assign node408 = (inp[1]) ? node410 : 3'b000;
					assign node410 = (inp[9]) ? node412 : 3'b000;
						assign node412 = (inp[5]) ? node428 : node413;
							assign node413 = (inp[6]) ? node425 : node414;
								assign node414 = (inp[7]) ? node420 : node415;
									assign node415 = (inp[10]) ? node417 : 3'b000;
										assign node417 = (inp[8]) ? 3'b100 : 3'b000;
									assign node420 = (inp[2]) ? 3'b100 : node421;
										assign node421 = (inp[10]) ? 3'b000 : 3'b000;
								assign node425 = (inp[7]) ? 3'b110 : 3'b010;
							assign node428 = (inp[2]) ? node436 : node429;
								assign node429 = (inp[8]) ? node431 : 3'b000;
									assign node431 = (inp[7]) ? node433 : 3'b000;
										assign node433 = (inp[11]) ? 3'b100 : 3'b000;
								assign node436 = (inp[6]) ? 3'b010 : 3'b000;

endmodule