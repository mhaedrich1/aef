module dtc_split66_bm85 (
	input  wire [12-1:0] inp,
	output wire [3-1:0] outp
);

	wire [3-1:0] node1;
	wire [3-1:0] node2;
	wire [3-1:0] node4;
	wire [3-1:0] node6;
	wire [3-1:0] node7;
	wire [3-1:0] node9;
	wire [3-1:0] node10;
	wire [3-1:0] node12;
	wire [3-1:0] node13;
	wire [3-1:0] node14;
	wire [3-1:0] node20;
	wire [3-1:0] node21;
	wire [3-1:0] node22;
	wire [3-1:0] node23;
	wire [3-1:0] node24;
	wire [3-1:0] node25;
	wire [3-1:0] node29;
	wire [3-1:0] node32;
	wire [3-1:0] node33;
	wire [3-1:0] node35;
	wire [3-1:0] node38;
	wire [3-1:0] node40;
	wire [3-1:0] node44;
	wire [3-1:0] node45;
	wire [3-1:0] node46;
	wire [3-1:0] node47;
	wire [3-1:0] node49;
	wire [3-1:0] node51;
	wire [3-1:0] node54;
	wire [3-1:0] node56;
	wire [3-1:0] node59;
	wire [3-1:0] node60;
	wire [3-1:0] node61;
	wire [3-1:0] node65;
	wire [3-1:0] node67;
	wire [3-1:0] node70;
	wire [3-1:0] node71;
	wire [3-1:0] node72;
	wire [3-1:0] node75;
	wire [3-1:0] node76;
	wire [3-1:0] node78;
	wire [3-1:0] node81;
	wire [3-1:0] node84;
	wire [3-1:0] node85;
	wire [3-1:0] node87;
	wire [3-1:0] node89;
	wire [3-1:0] node92;
	wire [3-1:0] node93;
	wire [3-1:0] node96;
	wire [3-1:0] node97;
	wire [3-1:0] node102;
	wire [3-1:0] node103;
	wire [3-1:0] node104;
	wire [3-1:0] node105;
	wire [3-1:0] node107;
	wire [3-1:0] node108;
	wire [3-1:0] node110;
	wire [3-1:0] node112;
	wire [3-1:0] node114;
	wire [3-1:0] node115;
	wire [3-1:0] node118;
	wire [3-1:0] node122;
	wire [3-1:0] node123;
	wire [3-1:0] node124;
	wire [3-1:0] node125;
	wire [3-1:0] node127;
	wire [3-1:0] node128;
	wire [3-1:0] node131;
	wire [3-1:0] node134;
	wire [3-1:0] node135;
	wire [3-1:0] node136;
	wire [3-1:0] node138;
	wire [3-1:0] node141;
	wire [3-1:0] node142;
	wire [3-1:0] node145;
	wire [3-1:0] node146;
	wire [3-1:0] node150;
	wire [3-1:0] node151;
	wire [3-1:0] node154;
	wire [3-1:0] node158;
	wire [3-1:0] node159;
	wire [3-1:0] node160;
	wire [3-1:0] node161;
	wire [3-1:0] node162;
	wire [3-1:0] node166;
	wire [3-1:0] node167;
	wire [3-1:0] node168;
	wire [3-1:0] node173;
	wire [3-1:0] node174;
	wire [3-1:0] node175;
	wire [3-1:0] node176;
	wire [3-1:0] node177;
	wire [3-1:0] node181;
	wire [3-1:0] node183;
	wire [3-1:0] node187;
	wire [3-1:0] node190;
	wire [3-1:0] node191;
	wire [3-1:0] node193;
	wire [3-1:0] node194;
	wire [3-1:0] node195;
	wire [3-1:0] node196;
	wire [3-1:0] node200;
	wire [3-1:0] node203;
	wire [3-1:0] node204;
	wire [3-1:0] node207;
	wire [3-1:0] node209;
	wire [3-1:0] node212;
	wire [3-1:0] node213;
	wire [3-1:0] node214;
	wire [3-1:0] node215;
	wire [3-1:0] node216;
	wire [3-1:0] node219;
	wire [3-1:0] node222;
	wire [3-1:0] node225;
	wire [3-1:0] node226;
	wire [3-1:0] node230;
	wire [3-1:0] node231;
	wire [3-1:0] node234;
	wire [3-1:0] node237;
	wire [3-1:0] node238;
	wire [3-1:0] node239;
	wire [3-1:0] node240;
	wire [3-1:0] node241;
	wire [3-1:0] node243;
	wire [3-1:0] node244;
	wire [3-1:0] node245;
	wire [3-1:0] node246;
	wire [3-1:0] node249;
	wire [3-1:0] node252;
	wire [3-1:0] node253;
	wire [3-1:0] node258;
	wire [3-1:0] node259;
	wire [3-1:0] node262;
	wire [3-1:0] node267;
	wire [3-1:0] node268;
	wire [3-1:0] node269;
	wire [3-1:0] node270;
	wire [3-1:0] node271;
	wire [3-1:0] node272;
	wire [3-1:0] node273;
	wire [3-1:0] node276;
	wire [3-1:0] node280;
	wire [3-1:0] node281;
	wire [3-1:0] node285;
	wire [3-1:0] node286;
	wire [3-1:0] node288;
	wire [3-1:0] node291;
	wire [3-1:0] node294;
	wire [3-1:0] node295;
	wire [3-1:0] node296;
	wire [3-1:0] node298;
	wire [3-1:0] node299;
	wire [3-1:0] node303;
	wire [3-1:0] node304;
	wire [3-1:0] node305;
	wire [3-1:0] node308;
	wire [3-1:0] node311;
	wire [3-1:0] node312;
	wire [3-1:0] node315;
	wire [3-1:0] node318;
	wire [3-1:0] node319;
	wire [3-1:0] node320;
	wire [3-1:0] node322;
	wire [3-1:0] node325;
	wire [3-1:0] node326;
	wire [3-1:0] node328;
	wire [3-1:0] node331;
	wire [3-1:0] node332;
	wire [3-1:0] node336;
	wire [3-1:0] node337;
	wire [3-1:0] node339;
	wire [3-1:0] node342;
	wire [3-1:0] node343;
	wire [3-1:0] node345;
	wire [3-1:0] node348;
	wire [3-1:0] node351;
	wire [3-1:0] node352;
	wire [3-1:0] node353;
	wire [3-1:0] node354;
	wire [3-1:0] node355;
	wire [3-1:0] node358;
	wire [3-1:0] node360;
	wire [3-1:0] node363;
	wire [3-1:0] node364;
	wire [3-1:0] node365;
	wire [3-1:0] node366;
	wire [3-1:0] node369;
	wire [3-1:0] node373;
	wire [3-1:0] node374;
	wire [3-1:0] node378;
	wire [3-1:0] node379;
	wire [3-1:0] node380;
	wire [3-1:0] node381;
	wire [3-1:0] node384;
	wire [3-1:0] node387;
	wire [3-1:0] node388;
	wire [3-1:0] node389;
	wire [3-1:0] node393;
	wire [3-1:0] node394;
	wire [3-1:0] node397;
	wire [3-1:0] node400;
	wire [3-1:0] node401;
	wire [3-1:0] node402;
	wire [3-1:0] node403;
	wire [3-1:0] node406;
	wire [3-1:0] node409;
	wire [3-1:0] node411;
	wire [3-1:0] node414;
	wire [3-1:0] node417;
	wire [3-1:0] node418;
	wire [3-1:0] node419;
	wire [3-1:0] node421;
	wire [3-1:0] node422;
	wire [3-1:0] node427;
	wire [3-1:0] node428;
	wire [3-1:0] node429;
	wire [3-1:0] node433;
	wire [3-1:0] node434;
	wire [3-1:0] node435;
	wire [3-1:0] node437;
	wire [3-1:0] node440;
	wire [3-1:0] node442;
	wire [3-1:0] node446;
	wire [3-1:0] node448;
	wire [3-1:0] node450;
	wire [3-1:0] node451;
	wire [3-1:0] node452;
	wire [3-1:0] node453;
	wire [3-1:0] node454;
	wire [3-1:0] node456;
	wire [3-1:0] node460;
	wire [3-1:0] node462;
	wire [3-1:0] node463;
	wire [3-1:0] node464;
	wire [3-1:0] node467;
	wire [3-1:0] node470;
	wire [3-1:0] node471;
	wire [3-1:0] node472;
	wire [3-1:0] node475;
	wire [3-1:0] node478;
	wire [3-1:0] node479;
	wire [3-1:0] node482;
	wire [3-1:0] node485;
	wire [3-1:0] node486;
	wire [3-1:0] node487;
	wire [3-1:0] node490;
	wire [3-1:0] node493;
	wire [3-1:0] node494;
	wire [3-1:0] node495;
	wire [3-1:0] node498;
	wire [3-1:0] node499;
	wire [3-1:0] node503;
	wire [3-1:0] node504;
	wire [3-1:0] node507;
	wire [3-1:0] node508;
	wire [3-1:0] node510;
	wire [3-1:0] node514;
	wire [3-1:0] node516;
	wire [3-1:0] node518;
	wire [3-1:0] node519;
	wire [3-1:0] node520;
	wire [3-1:0] node522;
	wire [3-1:0] node526;
	wire [3-1:0] node527;
	wire [3-1:0] node528;
	wire [3-1:0] node530;
	wire [3-1:0] node533;
	wire [3-1:0] node536;
	wire [3-1:0] node537;
	wire [3-1:0] node540;
	wire [3-1:0] node541;

	assign outp = (inp[0]) ? node102 : node1;
		assign node1 = (inp[6]) ? 3'b000 : node2;
			assign node2 = (inp[3]) ? node4 : 3'b000;
				assign node4 = (inp[9]) ? node6 : 3'b000;
					assign node6 = (inp[4]) ? node20 : node7;
						assign node7 = (inp[2]) ? node9 : 3'b000;
							assign node9 = (inp[7]) ? 3'b000 : node10;
								assign node10 = (inp[1]) ? node12 : 3'b000;
									assign node12 = (inp[10]) ? 3'b100 : node13;
										assign node13 = (inp[5]) ? 3'b000 : node14;
											assign node14 = (inp[8]) ? 3'b100 : 3'b000;
						assign node20 = (inp[1]) ? node44 : node21;
							assign node21 = (inp[7]) ? 3'b000 : node22;
								assign node22 = (inp[2]) ? node32 : node23;
									assign node23 = (inp[10]) ? node29 : node24;
										assign node24 = (inp[8]) ? 3'b000 : node25;
											assign node25 = (inp[5]) ? 3'b100 : 3'b000;
										assign node29 = (inp[5]) ? 3'b010 : 3'b000;
									assign node32 = (inp[10]) ? node38 : node33;
										assign node33 = (inp[5]) ? node35 : 3'b010;
											assign node35 = (inp[8]) ? 3'b011 : 3'b010;
										assign node38 = (inp[5]) ? node40 : 3'b000;
											assign node40 = (inp[8]) ? 3'b000 : 3'b001;
							assign node44 = (inp[7]) ? node70 : node45;
								assign node45 = (inp[11]) ? node59 : node46;
									assign node46 = (inp[10]) ? node54 : node47;
										assign node47 = (inp[2]) ? node49 : 3'b110;
											assign node49 = (inp[8]) ? node51 : 3'b001;
												assign node51 = (inp[5]) ? 3'b110 : 3'b101;
										assign node54 = (inp[8]) ? node56 : 3'b001;
											assign node56 = (inp[5]) ? 3'b110 : 3'b010;
									assign node59 = (inp[10]) ? node65 : node60;
										assign node60 = (inp[2]) ? 3'b001 : node61;
											assign node61 = (inp[8]) ? 3'b010 : 3'b001;
										assign node65 = (inp[2]) ? node67 : 3'b101;
											assign node67 = (inp[8]) ? 3'b101 : 3'b001;
								assign node70 = (inp[2]) ? node84 : node71;
									assign node71 = (inp[8]) ? node75 : node72;
										assign node72 = (inp[10]) ? 3'b110 : 3'b100;
										assign node75 = (inp[5]) ? node81 : node76;
											assign node76 = (inp[10]) ? node78 : 3'b100;
												assign node78 = (inp[11]) ? 3'b000 : 3'b100;
											assign node81 = (inp[11]) ? 3'b100 : 3'b000;
									assign node84 = (inp[10]) ? node92 : node85;
										assign node85 = (inp[8]) ? node87 : 3'b010;
											assign node87 = (inp[11]) ? node89 : 3'b100;
												assign node89 = (inp[5]) ? 3'b100 : 3'b000;
										assign node92 = (inp[8]) ? node96 : node93;
											assign node93 = (inp[11]) ? 3'b010 : 3'b110;
											assign node96 = (inp[5]) ? 3'b010 : node97;
												assign node97 = (inp[11]) ? 3'b110 : 3'b010;
		assign node102 = (inp[6]) ? node446 : node103;
			assign node103 = (inp[3]) ? node237 : node104;
				assign node104 = (inp[4]) ? node122 : node105;
					assign node105 = (inp[5]) ? node107 : 3'b000;
						assign node107 = (inp[7]) ? 3'b000 : node108;
							assign node108 = (inp[9]) ? node110 : 3'b000;
								assign node110 = (inp[1]) ? node112 : 3'b000;
									assign node112 = (inp[2]) ? node114 : 3'b000;
										assign node114 = (inp[8]) ? node118 : node115;
											assign node115 = (inp[10]) ? 3'b100 : 3'b000;
											assign node118 = (inp[10]) ? 3'b000 : 3'b100;
					assign node122 = (inp[9]) ? node158 : node123;
						assign node123 = (inp[7]) ? 3'b100 : node124;
							assign node124 = (inp[11]) ? node134 : node125;
								assign node125 = (inp[5]) ? node127 : 3'b100;
									assign node127 = (inp[8]) ? node131 : node128;
										assign node128 = (inp[10]) ? 3'b000 : 3'b100;
										assign node131 = (inp[10]) ? 3'b100 : 3'b000;
								assign node134 = (inp[5]) ? node150 : node135;
									assign node135 = (inp[2]) ? node141 : node136;
										assign node136 = (inp[10]) ? node138 : 3'b000;
											assign node138 = (inp[8]) ? 3'b000 : 3'b100;
										assign node141 = (inp[1]) ? node145 : node142;
											assign node142 = (inp[8]) ? 3'b000 : 3'b100;
											assign node145 = (inp[10]) ? 3'b100 : node146;
												assign node146 = (inp[8]) ? 3'b100 : 3'b000;
									assign node150 = (inp[8]) ? node154 : node151;
										assign node151 = (inp[10]) ? 3'b000 : 3'b100;
										assign node154 = (inp[10]) ? 3'b100 : 3'b000;
						assign node158 = (inp[2]) ? node190 : node159;
							assign node159 = (inp[8]) ? node173 : node160;
								assign node160 = (inp[10]) ? node166 : node161;
									assign node161 = (inp[7]) ? 3'b100 : node162;
										assign node162 = (inp[5]) ? 3'b000 : 3'b100;
									assign node166 = (inp[7]) ? 3'b000 : node167;
										assign node167 = (inp[5]) ? 3'b100 : node168;
											assign node168 = (inp[1]) ? 3'b000 : 3'b100;
								assign node173 = (inp[10]) ? node187 : node174;
									assign node174 = (inp[7]) ? 3'b000 : node175;
										assign node175 = (inp[11]) ? node181 : node176;
											assign node176 = (inp[5]) ? 3'b000 : node177;
												assign node177 = (inp[1]) ? 3'b000 : 3'b100;
											assign node181 = (inp[1]) ? node183 : 3'b000;
												assign node183 = (inp[5]) ? 3'b100 : 3'b000;
									assign node187 = (inp[7]) ? 3'b100 : 3'b000;
							assign node190 = (inp[1]) ? node212 : node191;
								assign node191 = (inp[7]) ? node193 : 3'b100;
									assign node193 = (inp[11]) ? node203 : node194;
										assign node194 = (inp[5]) ? node200 : node195;
											assign node195 = (inp[8]) ? 3'b000 : node196;
												assign node196 = (inp[10]) ? 3'b000 : 3'b100;
											assign node200 = (inp[8]) ? 3'b100 : 3'b000;
										assign node203 = (inp[5]) ? node207 : node204;
											assign node204 = (inp[10]) ? 3'b100 : 3'b000;
											assign node207 = (inp[10]) ? node209 : 3'b100;
												assign node209 = (inp[8]) ? 3'b100 : 3'b000;
								assign node212 = (inp[7]) ? node230 : node213;
									assign node213 = (inp[5]) ? node225 : node214;
										assign node214 = (inp[10]) ? node222 : node215;
											assign node215 = (inp[11]) ? node219 : node216;
												assign node216 = (inp[8]) ? 3'b010 : 3'b100;
												assign node219 = (inp[8]) ? 3'b100 : 3'b010;
											assign node222 = (inp[8]) ? 3'b010 : 3'b110;
										assign node225 = (inp[10]) ? 3'b001 : node226;
											assign node226 = (inp[8]) ? 3'b011 : 3'b110;
									assign node230 = (inp[10]) ? node234 : node231;
										assign node231 = (inp[8]) ? 3'b000 : 3'b100;
										assign node234 = (inp[8]) ? 3'b100 : 3'b000;
				assign node237 = (inp[9]) ? node267 : node238;
					assign node238 = (inp[7]) ? 3'b001 : node239;
						assign node239 = (inp[4]) ? 3'b111 : node240;
							assign node240 = (inp[5]) ? node258 : node241;
								assign node241 = (inp[11]) ? node243 : 3'b001;
									assign node243 = (inp[1]) ? 3'b001 : node244;
										assign node244 = (inp[2]) ? node252 : node245;
											assign node245 = (inp[8]) ? node249 : node246;
												assign node246 = (inp[10]) ? 3'b001 : 3'b101;
												assign node249 = (inp[10]) ? 3'b101 : 3'b001;
											assign node252 = (inp[8]) ? 3'b001 : node253;
												assign node253 = (inp[10]) ? 3'b001 : 3'b101;
								assign node258 = (inp[10]) ? node262 : node259;
									assign node259 = (inp[8]) ? 3'b101 : 3'b001;
									assign node262 = (inp[8]) ? 3'b001 : 3'b101;
					assign node267 = (inp[4]) ? node351 : node268;
						assign node268 = (inp[1]) ? node294 : node269;
							assign node269 = (inp[8]) ? node285 : node270;
								assign node270 = (inp[10]) ? node280 : node271;
									assign node271 = (inp[7]) ? 3'b010 : node272;
										assign node272 = (inp[5]) ? node276 : node273;
											assign node273 = (inp[11]) ? 3'b110 : 3'b010;
											assign node276 = (inp[11]) ? 3'b001 : 3'b110;
									assign node280 = (inp[7]) ? 3'b110 : node281;
										assign node281 = (inp[5]) ? 3'b110 : 3'b010;
								assign node285 = (inp[7]) ? node291 : node286;
									assign node286 = (inp[5]) ? node288 : 3'b010;
										assign node288 = (inp[2]) ? 3'b010 : 3'b110;
									assign node291 = (inp[10]) ? 3'b001 : 3'b101;
							assign node294 = (inp[7]) ? node318 : node295;
								assign node295 = (inp[5]) ? node303 : node296;
									assign node296 = (inp[11]) ? node298 : 3'b101;
										assign node298 = (inp[10]) ? 3'b101 : node299;
											assign node299 = (inp[8]) ? 3'b001 : 3'b011;
									assign node303 = (inp[2]) ? node311 : node304;
										assign node304 = (inp[10]) ? node308 : node305;
											assign node305 = (inp[8]) ? 3'b011 : 3'b101;
											assign node308 = (inp[8]) ? 3'b101 : 3'b011;
										assign node311 = (inp[8]) ? node315 : node312;
											assign node312 = (inp[10]) ? 3'b111 : 3'b011;
											assign node315 = (inp[10]) ? 3'b011 : 3'b111;
								assign node318 = (inp[5]) ? node336 : node319;
									assign node319 = (inp[2]) ? node325 : node320;
										assign node320 = (inp[8]) ? node322 : 3'b101;
											assign node322 = (inp[10]) ? 3'b010 : 3'b101;
										assign node325 = (inp[11]) ? node331 : node326;
											assign node326 = (inp[8]) ? node328 : 3'b110;
												assign node328 = (inp[10]) ? 3'b010 : 3'b110;
											assign node331 = (inp[10]) ? 3'b010 : node332;
												assign node332 = (inp[8]) ? 3'b110 : 3'b010;
									assign node336 = (inp[10]) ? node342 : node337;
										assign node337 = (inp[8]) ? node339 : 3'b010;
											assign node339 = (inp[2]) ? 3'b110 : 3'b101;
										assign node342 = (inp[8]) ? node348 : node343;
											assign node343 = (inp[2]) ? node345 : 3'b101;
												assign node345 = (inp[11]) ? 3'b101 : 3'b110;
											assign node348 = (inp[2]) ? 3'b001 : 3'b010;
						assign node351 = (inp[1]) ? node417 : node352;
							assign node352 = (inp[7]) ? node378 : node353;
								assign node353 = (inp[5]) ? node363 : node354;
									assign node354 = (inp[10]) ? node358 : node355;
										assign node355 = (inp[8]) ? 3'b110 : 3'b001;
										assign node358 = (inp[8]) ? node360 : 3'b101;
											assign node360 = (inp[2]) ? 3'b101 : 3'b001;
									assign node363 = (inp[2]) ? node373 : node364;
										assign node364 = (inp[8]) ? 3'b101 : node365;
											assign node365 = (inp[11]) ? node369 : node366;
												assign node366 = (inp[10]) ? 3'b011 : 3'b101;
												assign node369 = (inp[10]) ? 3'b111 : 3'b011;
										assign node373 = (inp[10]) ? 3'b111 : node374;
											assign node374 = (inp[8]) ? 3'b011 : 3'b111;
								assign node378 = (inp[10]) ? node400 : node379;
									assign node379 = (inp[11]) ? node387 : node380;
										assign node380 = (inp[8]) ? node384 : node381;
											assign node381 = (inp[2]) ? 3'b111 : 3'b110;
											assign node384 = (inp[5]) ? 3'b100 : 3'b101;
										assign node387 = (inp[5]) ? node393 : node388;
											assign node388 = (inp[8]) ? 3'b101 : node389;
												assign node389 = (inp[2]) ? 3'b100 : 3'b000;
											assign node393 = (inp[8]) ? node397 : node394;
												assign node394 = (inp[2]) ? 3'b101 : 3'b001;
												assign node397 = (inp[2]) ? 3'b001 : 3'b100;
									assign node400 = (inp[5]) ? node414 : node401;
										assign node401 = (inp[8]) ? node409 : node402;
											assign node402 = (inp[2]) ? node406 : node403;
												assign node403 = (inp[11]) ? 3'b110 : 3'b100;
												assign node406 = (inp[11]) ? 3'b011 : 3'b001;
											assign node409 = (inp[11]) ? node411 : 3'b110;
												assign node411 = (inp[2]) ? 3'b110 : 3'b010;
										assign node414 = (inp[8]) ? 3'b011 : 3'b001;
							assign node417 = (inp[7]) ? node427 : node418;
								assign node418 = (inp[2]) ? 3'b111 : node419;
									assign node419 = (inp[5]) ? node421 : 3'b111;
										assign node421 = (inp[11]) ? 3'b111 : node422;
											assign node422 = (inp[10]) ? 3'b111 : 3'b011;
								assign node427 = (inp[2]) ? node433 : node428;
									assign node428 = (inp[8]) ? 3'b001 : node429;
										assign node429 = (inp[10]) ? 3'b111 : 3'b011;
									assign node433 = (inp[11]) ? 3'b111 : node434;
										assign node434 = (inp[8]) ? node440 : node435;
											assign node435 = (inp[5]) ? node437 : 3'b111;
												assign node437 = (inp[10]) ? 3'b111 : 3'b011;
											assign node440 = (inp[10]) ? node442 : 3'b101;
												assign node442 = (inp[5]) ? 3'b011 : 3'b111;
			assign node446 = (inp[3]) ? node448 : 3'b000;
				assign node448 = (inp[9]) ? node450 : 3'b000;
					assign node450 = (inp[7]) ? node514 : node451;
						assign node451 = (inp[4]) ? node485 : node452;
							assign node452 = (inp[2]) ? node460 : node453;
								assign node453 = (inp[8]) ? 3'b000 : node454;
									assign node454 = (inp[11]) ? node456 : 3'b000;
										assign node456 = (inp[5]) ? 3'b010 : 3'b000;
								assign node460 = (inp[1]) ? node462 : 3'b000;
									assign node462 = (inp[8]) ? node470 : node463;
										assign node463 = (inp[10]) ? node467 : node464;
											assign node464 = (inp[11]) ? 3'b010 : 3'b000;
											assign node467 = (inp[11]) ? 3'b110 : 3'b100;
										assign node470 = (inp[11]) ? node478 : node471;
											assign node471 = (inp[5]) ? node475 : node472;
												assign node472 = (inp[10]) ? 3'b000 : 3'b100;
												assign node475 = (inp[10]) ? 3'b100 : 3'b000;
											assign node478 = (inp[5]) ? node482 : node479;
												assign node479 = (inp[10]) ? 3'b000 : 3'b100;
												assign node482 = (inp[10]) ? 3'b100 : 3'b000;
							assign node485 = (inp[1]) ? node493 : node486;
								assign node486 = (inp[10]) ? node490 : node487;
									assign node487 = (inp[8]) ? 3'b000 : 3'b100;
									assign node490 = (inp[8]) ? 3'b010 : 3'b110;
								assign node493 = (inp[10]) ? node503 : node494;
									assign node494 = (inp[2]) ? node498 : node495;
										assign node495 = (inp[8]) ? 3'b010 : 3'b110;
										assign node498 = (inp[8]) ? 3'b110 : node499;
											assign node499 = (inp[5]) ? 3'b001 : 3'b110;
									assign node503 = (inp[2]) ? node507 : node504;
										assign node504 = (inp[8]) ? 3'b101 : 3'b001;
										assign node507 = (inp[8]) ? 3'b110 : node508;
											assign node508 = (inp[11]) ? node510 : 3'b101;
												assign node510 = (inp[5]) ? 3'b011 : 3'b111;
						assign node514 = (inp[4]) ? node516 : 3'b000;
							assign node516 = (inp[2]) ? node518 : 3'b000;
								assign node518 = (inp[1]) ? node526 : node519;
									assign node519 = (inp[10]) ? 3'b000 : node520;
										assign node520 = (inp[11]) ? node522 : 3'b000;
											assign node522 = (inp[5]) ? 3'b100 : 3'b000;
									assign node526 = (inp[10]) ? node536 : node527;
										assign node527 = (inp[5]) ? node533 : node528;
											assign node528 = (inp[11]) ? node530 : 3'b000;
												assign node530 = (inp[8]) ? 3'b000 : 3'b100;
											assign node533 = (inp[8]) ? 3'b100 : 3'b010;
										assign node536 = (inp[8]) ? node540 : node537;
											assign node537 = (inp[5]) ? 3'b110 : 3'b010;
											assign node540 = (inp[5]) ? 3'b010 : node541;
												assign node541 = (inp[11]) ? 3'b100 : 3'b000;

endmodule