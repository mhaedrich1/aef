module dtc_split125_bm76 (
	input  wire [12-1:0] inp,
	output wire [3-1:0] outp
);

	wire [3-1:0] node1;
	wire [3-1:0] node2;
	wire [3-1:0] node3;
	wire [3-1:0] node4;
	wire [3-1:0] node6;
	wire [3-1:0] node8;
	wire [3-1:0] node10;
	wire [3-1:0] node11;
	wire [3-1:0] node15;
	wire [3-1:0] node16;
	wire [3-1:0] node17;
	wire [3-1:0] node19;
	wire [3-1:0] node22;
	wire [3-1:0] node24;
	wire [3-1:0] node25;
	wire [3-1:0] node28;
	wire [3-1:0] node31;
	wire [3-1:0] node32;
	wire [3-1:0] node33;
	wire [3-1:0] node37;
	wire [3-1:0] node40;
	wire [3-1:0] node41;
	wire [3-1:0] node42;
	wire [3-1:0] node43;
	wire [3-1:0] node46;
	wire [3-1:0] node47;
	wire [3-1:0] node48;
	wire [3-1:0] node52;
	wire [3-1:0] node55;
	wire [3-1:0] node56;
	wire [3-1:0] node58;
	wire [3-1:0] node60;
	wire [3-1:0] node63;
	wire [3-1:0] node65;
	wire [3-1:0] node68;
	wire [3-1:0] node69;
	wire [3-1:0] node70;
	wire [3-1:0] node72;
	wire [3-1:0] node76;
	wire [3-1:0] node77;
	wire [3-1:0] node78;
	wire [3-1:0] node79;
	wire [3-1:0] node83;
	wire [3-1:0] node86;
	wire [3-1:0] node87;
	wire [3-1:0] node91;
	wire [3-1:0] node92;
	wire [3-1:0] node93;
	wire [3-1:0] node94;
	wire [3-1:0] node95;
	wire [3-1:0] node96;
	wire [3-1:0] node100;
	wire [3-1:0] node102;
	wire [3-1:0] node103;
	wire [3-1:0] node104;
	wire [3-1:0] node107;
	wire [3-1:0] node108;
	wire [3-1:0] node113;
	wire [3-1:0] node114;
	wire [3-1:0] node116;
	wire [3-1:0] node119;
	wire [3-1:0] node120;
	wire [3-1:0] node123;
	wire [3-1:0] node126;
	wire [3-1:0] node127;
	wire [3-1:0] node129;
	wire [3-1:0] node130;
	wire [3-1:0] node134;
	wire [3-1:0] node135;
	wire [3-1:0] node137;
	wire [3-1:0] node138;
	wire [3-1:0] node142;
	wire [3-1:0] node143;
	wire [3-1:0] node145;
	wire [3-1:0] node148;
	wire [3-1:0] node151;
	wire [3-1:0] node152;
	wire [3-1:0] node153;
	wire [3-1:0] node154;
	wire [3-1:0] node157;
	wire [3-1:0] node160;
	wire [3-1:0] node161;
	wire [3-1:0] node164;
	wire [3-1:0] node166;
	wire [3-1:0] node169;
	wire [3-1:0] node170;
	wire [3-1:0] node171;
	wire [3-1:0] node173;
	wire [3-1:0] node176;
	wire [3-1:0] node177;
	wire [3-1:0] node181;
	wire [3-1:0] node182;
	wire [3-1:0] node184;
	wire [3-1:0] node186;
	wire [3-1:0] node189;
	wire [3-1:0] node190;
	wire [3-1:0] node194;
	wire [3-1:0] node195;
	wire [3-1:0] node196;
	wire [3-1:0] node197;
	wire [3-1:0] node198;
	wire [3-1:0] node199;
	wire [3-1:0] node200;
	wire [3-1:0] node202;
	wire [3-1:0] node206;
	wire [3-1:0] node209;
	wire [3-1:0] node212;
	wire [3-1:0] node213;
	wire [3-1:0] node215;
	wire [3-1:0] node218;
	wire [3-1:0] node219;
	wire [3-1:0] node220;
	wire [3-1:0] node221;
	wire [3-1:0] node225;
	wire [3-1:0] node226;
	wire [3-1:0] node230;
	wire [3-1:0] node232;
	wire [3-1:0] node234;
	wire [3-1:0] node236;
	wire [3-1:0] node239;
	wire [3-1:0] node240;
	wire [3-1:0] node241;
	wire [3-1:0] node242;
	wire [3-1:0] node243;
	wire [3-1:0] node245;
	wire [3-1:0] node249;
	wire [3-1:0] node250;
	wire [3-1:0] node252;
	wire [3-1:0] node254;
	wire [3-1:0] node256;
	wire [3-1:0] node260;
	wire [3-1:0] node261;
	wire [3-1:0] node262;
	wire [3-1:0] node265;
	wire [3-1:0] node267;
	wire [3-1:0] node270;
	wire [3-1:0] node272;
	wire [3-1:0] node275;
	wire [3-1:0] node276;
	wire [3-1:0] node277;
	wire [3-1:0] node279;
	wire [3-1:0] node284;
	wire [3-1:0] node285;
	wire [3-1:0] node286;
	wire [3-1:0] node287;
	wire [3-1:0] node288;
	wire [3-1:0] node289;
	wire [3-1:0] node293;
	wire [3-1:0] node294;
	wire [3-1:0] node296;
	wire [3-1:0] node300;
	wire [3-1:0] node301;
	wire [3-1:0] node302;

	assign outp = (inp[9]) ? node194 : node1;
		assign node1 = (inp[6]) ? node91 : node2;
			assign node2 = (inp[10]) ? node40 : node3;
				assign node3 = (inp[7]) ? node15 : node4;
					assign node4 = (inp[8]) ? node6 : 3'b111;
						assign node6 = (inp[11]) ? node8 : 3'b111;
							assign node8 = (inp[3]) ? node10 : 3'b111;
								assign node10 = (inp[4]) ? 3'b011 : node11;
									assign node11 = (inp[0]) ? 3'b011 : 3'b111;
					assign node15 = (inp[8]) ? node31 : node16;
						assign node16 = (inp[11]) ? node22 : node17;
							assign node17 = (inp[1]) ? node19 : 3'b111;
								assign node19 = (inp[0]) ? 3'b011 : 3'b111;
							assign node22 = (inp[5]) ? node24 : 3'b011;
								assign node24 = (inp[3]) ? node28 : node25;
									assign node25 = (inp[2]) ? 3'b111 : 3'b011;
									assign node28 = (inp[4]) ? 3'b101 : 3'b011;
						assign node31 = (inp[4]) ? node37 : node32;
							assign node32 = (inp[11]) ? 3'b011 : node33;
								assign node33 = (inp[3]) ? 3'b011 : 3'b111;
							assign node37 = (inp[11]) ? 3'b101 : 3'b011;
				assign node40 = (inp[7]) ? node68 : node41;
					assign node41 = (inp[11]) ? node55 : node42;
						assign node42 = (inp[3]) ? node46 : node43;
							assign node43 = (inp[8]) ? 3'b011 : 3'b111;
							assign node46 = (inp[0]) ? node52 : node47;
								assign node47 = (inp[8]) ? 3'b011 : node48;
									assign node48 = (inp[1]) ? 3'b011 : 3'b111;
								assign node52 = (inp[8]) ? 3'b101 : 3'b011;
						assign node55 = (inp[1]) ? node63 : node56;
							assign node56 = (inp[0]) ? node58 : 3'b101;
								assign node58 = (inp[4]) ? node60 : 3'b011;
									assign node60 = (inp[8]) ? 3'b001 : 3'b101;
							assign node63 = (inp[3]) ? node65 : 3'b011;
								assign node65 = (inp[8]) ? 3'b001 : 3'b101;
					assign node68 = (inp[11]) ? node76 : node69;
						assign node69 = (inp[8]) ? 3'b001 : node70;
							assign node70 = (inp[5]) ? node72 : 3'b101;
								assign node72 = (inp[2]) ? 3'b001 : 3'b101;
						assign node76 = (inp[3]) ? node86 : node77;
							assign node77 = (inp[8]) ? node83 : node78;
								assign node78 = (inp[5]) ? 3'b001 : node79;
									assign node79 = (inp[0]) ? 3'b001 : 3'b101;
								assign node83 = (inp[2]) ? 3'b001 : 3'b110;
							assign node86 = (inp[1]) ? 3'b110 : node87;
								assign node87 = (inp[8]) ? 3'b110 : 3'b001;
			assign node91 = (inp[10]) ? node151 : node92;
				assign node92 = (inp[7]) ? node126 : node93;
					assign node93 = (inp[0]) ? node113 : node94;
						assign node94 = (inp[1]) ? node100 : node95;
							assign node95 = (inp[3]) ? 3'b001 : node96;
								assign node96 = (inp[8]) ? 3'b001 : 3'b101;
							assign node100 = (inp[8]) ? node102 : 3'b011;
								assign node102 = (inp[4]) ? 3'b001 : node103;
									assign node103 = (inp[5]) ? node107 : node104;
										assign node104 = (inp[2]) ? 3'b011 : 3'b001;
										assign node107 = (inp[3]) ? 3'b110 : node108;
											assign node108 = (inp[11]) ? 3'b001 : 3'b101;
						assign node113 = (inp[11]) ? node119 : node114;
							assign node114 = (inp[8]) ? node116 : 3'b101;
								assign node116 = (inp[4]) ? 3'b001 : 3'b101;
							assign node119 = (inp[8]) ? node123 : node120;
								assign node120 = (inp[3]) ? 3'b001 : 3'b101;
								assign node123 = (inp[3]) ? 3'b110 : 3'b001;
					assign node126 = (inp[11]) ? node134 : node127;
						assign node127 = (inp[8]) ? node129 : 3'b001;
							assign node129 = (inp[3]) ? 3'b110 : node130;
								assign node130 = (inp[4]) ? 3'b110 : 3'b001;
						assign node134 = (inp[5]) ? node142 : node135;
							assign node135 = (inp[0]) ? node137 : 3'b110;
								assign node137 = (inp[1]) ? 3'b110 : node138;
									assign node138 = (inp[3]) ? 3'b110 : 3'b001;
							assign node142 = (inp[4]) ? node148 : node143;
								assign node143 = (inp[8]) ? node145 : 3'b001;
									assign node145 = (inp[2]) ? 3'b010 : 3'b100;
								assign node148 = (inp[0]) ? 3'b010 : 3'b110;
				assign node151 = (inp[7]) ? node169 : node152;
					assign node152 = (inp[3]) ? node160 : node153;
						assign node153 = (inp[8]) ? node157 : node154;
							assign node154 = (inp[11]) ? 3'b110 : 3'b001;
							assign node157 = (inp[11]) ? 3'b010 : 3'b110;
						assign node160 = (inp[11]) ? node164 : node161;
							assign node161 = (inp[8]) ? 3'b010 : 3'b110;
							assign node164 = (inp[8]) ? node166 : 3'b010;
								assign node166 = (inp[4]) ? 3'b100 : 3'b010;
					assign node169 = (inp[11]) ? node181 : node170;
						assign node170 = (inp[8]) ? node176 : node171;
							assign node171 = (inp[5]) ? node173 : 3'b010;
								assign node173 = (inp[3]) ? 3'b100 : 3'b010;
							assign node176 = (inp[1]) ? 3'b100 : node177;
								assign node177 = (inp[2]) ? 3'b100 : 3'b000;
						assign node181 = (inp[8]) ? node189 : node182;
							assign node182 = (inp[2]) ? node184 : 3'b100;
								assign node184 = (inp[4]) ? node186 : 3'b100;
									assign node186 = (inp[3]) ? 3'b000 : 3'b100;
							assign node189 = (inp[0]) ? 3'b000 : node190;
								assign node190 = (inp[1]) ? 3'b000 : 3'b100;
		assign node194 = (inp[6]) ? node284 : node195;
			assign node195 = (inp[10]) ? node239 : node196;
				assign node196 = (inp[8]) ? node212 : node197;
					assign node197 = (inp[7]) ? node209 : node198;
						assign node198 = (inp[11]) ? node206 : node199;
							assign node199 = (inp[3]) ? 3'b001 : node200;
								assign node200 = (inp[4]) ? node202 : 3'b101;
									assign node202 = (inp[2]) ? 3'b001 : 3'b101;
							assign node206 = (inp[0]) ? 3'b110 : 3'b001;
						assign node209 = (inp[4]) ? 3'b010 : 3'b110;
					assign node212 = (inp[7]) ? node218 : node213;
						assign node213 = (inp[11]) ? node215 : 3'b110;
							assign node215 = (inp[3]) ? 3'b010 : 3'b110;
						assign node218 = (inp[11]) ? node230 : node219;
							assign node219 = (inp[5]) ? node225 : node220;
								assign node220 = (inp[3]) ? 3'b010 : node221;
									assign node221 = (inp[4]) ? 3'b010 : 3'b110;
								assign node225 = (inp[3]) ? 3'b100 : node226;
									assign node226 = (inp[0]) ? 3'b010 : 3'b110;
							assign node230 = (inp[3]) ? node232 : 3'b010;
								assign node232 = (inp[1]) ? node234 : 3'b100;
									assign node234 = (inp[0]) ? node236 : 3'b100;
										assign node236 = (inp[4]) ? 3'b000 : 3'b100;
				assign node239 = (inp[7]) ? node275 : node240;
					assign node240 = (inp[11]) ? node260 : node241;
						assign node241 = (inp[8]) ? node249 : node242;
							assign node242 = (inp[3]) ? 3'b010 : node243;
								assign node243 = (inp[5]) ? node245 : 3'b110;
									assign node245 = (inp[1]) ? 3'b010 : 3'b110;
							assign node249 = (inp[3]) ? 3'b100 : node250;
								assign node250 = (inp[1]) ? node252 : 3'b100;
									assign node252 = (inp[0]) ? node254 : 3'b010;
										assign node254 = (inp[2]) ? node256 : 3'b010;
											assign node256 = (inp[5]) ? 3'b100 : 3'b010;
						assign node260 = (inp[0]) ? node270 : node261;
							assign node261 = (inp[1]) ? node265 : node262;
								assign node262 = (inp[8]) ? 3'b000 : 3'b100;
								assign node265 = (inp[8]) ? node267 : 3'b000;
									assign node267 = (inp[4]) ? 3'b000 : 3'b100;
							assign node270 = (inp[1]) ? node272 : 3'b000;
								assign node272 = (inp[4]) ? 3'b000 : 3'b100;
					assign node275 = (inp[11]) ? 3'b000 : node276;
						assign node276 = (inp[8]) ? 3'b000 : node277;
							assign node277 = (inp[3]) ? node279 : 3'b100;
								assign node279 = (inp[4]) ? 3'b000 : 3'b100;
			assign node284 = (inp[7]) ? 3'b000 : node285;
				assign node285 = (inp[10]) ? 3'b000 : node286;
					assign node286 = (inp[11]) ? node300 : node287;
						assign node287 = (inp[8]) ? node293 : node288;
							assign node288 = (inp[4]) ? 3'b100 : node289;
								assign node289 = (inp[3]) ? 3'b100 : 3'b010;
							assign node293 = (inp[3]) ? 3'b000 : node294;
								assign node294 = (inp[2]) ? node296 : 3'b100;
									assign node296 = (inp[1]) ? 3'b100 : 3'b000;
						assign node300 = (inp[8]) ? 3'b000 : node301;
							assign node301 = (inp[2]) ? 3'b000 : node302;
								assign node302 = (inp[5]) ? 3'b100 : 3'b000;

endmodule