module dtc_split25_bm34 (
	input  wire [9-1:0] inp,
	output wire [5-1:0] outp
);

	wire [5-1:0] node1;
	wire [5-1:0] node2;
	wire [5-1:0] node3;
	wire [5-1:0] node4;
	wire [5-1:0] node6;
	wire [5-1:0] node7;
	wire [5-1:0] node8;
	wire [5-1:0] node12;
	wire [5-1:0] node14;
	wire [5-1:0] node17;
	wire [5-1:0] node18;
	wire [5-1:0] node19;
	wire [5-1:0] node23;
	wire [5-1:0] node24;
	wire [5-1:0] node27;
	wire [5-1:0] node29;
	wire [5-1:0] node32;
	wire [5-1:0] node33;
	wire [5-1:0] node34;
	wire [5-1:0] node35;
	wire [5-1:0] node38;
	wire [5-1:0] node40;
	wire [5-1:0] node42;
	wire [5-1:0] node45;
	wire [5-1:0] node47;
	wire [5-1:0] node50;
	wire [5-1:0] node51;
	wire [5-1:0] node52;
	wire [5-1:0] node53;
	wire [5-1:0] node56;
	wire [5-1:0] node60;
	wire [5-1:0] node61;
	wire [5-1:0] node65;
	wire [5-1:0] node66;
	wire [5-1:0] node67;
	wire [5-1:0] node68;
	wire [5-1:0] node70;
	wire [5-1:0] node74;
	wire [5-1:0] node75;
	wire [5-1:0] node76;
	wire [5-1:0] node79;
	wire [5-1:0] node80;
	wire [5-1:0] node84;
	wire [5-1:0] node85;
	wire [5-1:0] node88;
	wire [5-1:0] node90;
	wire [5-1:0] node93;
	wire [5-1:0] node94;
	wire [5-1:0] node95;
	wire [5-1:0] node96;
	wire [5-1:0] node100;
	wire [5-1:0] node103;
	wire [5-1:0] node104;
	wire [5-1:0] node105;
	wire [5-1:0] node106;
	wire [5-1:0] node109;
	wire [5-1:0] node112;
	wire [5-1:0] node115;
	wire [5-1:0] node116;
	wire [5-1:0] node120;
	wire [5-1:0] node121;
	wire [5-1:0] node122;
	wire [5-1:0] node123;
	wire [5-1:0] node124;
	wire [5-1:0] node126;
	wire [5-1:0] node129;
	wire [5-1:0] node130;
	wire [5-1:0] node133;
	wire [5-1:0] node136;
	wire [5-1:0] node137;
	wire [5-1:0] node138;
	wire [5-1:0] node139;
	wire [5-1:0] node142;
	wire [5-1:0] node144;
	wire [5-1:0] node149;
	wire [5-1:0] node150;
	wire [5-1:0] node152;
	wire [5-1:0] node154;
	wire [5-1:0] node157;
	wire [5-1:0] node158;
	wire [5-1:0] node160;
	wire [5-1:0] node163;
	wire [5-1:0] node166;
	wire [5-1:0] node167;
	wire [5-1:0] node168;
	wire [5-1:0] node169;
	wire [5-1:0] node171;
	wire [5-1:0] node174;
	wire [5-1:0] node175;
	wire [5-1:0] node176;
	wire [5-1:0] node180;
	wire [5-1:0] node183;
	wire [5-1:0] node184;
	wire [5-1:0] node185;
	wire [5-1:0] node186;
	wire [5-1:0] node190;
	wire [5-1:0] node193;
	wire [5-1:0] node196;
	wire [5-1:0] node197;
	wire [5-1:0] node198;
	wire [5-1:0] node199;
	wire [5-1:0] node202;
	wire [5-1:0] node205;
	wire [5-1:0] node208;
	wire [5-1:0] node209;
	wire [5-1:0] node210;
	wire [5-1:0] node211;
	wire [5-1:0] node216;
	wire [5-1:0] node217;

	assign outp = (inp[2]) ? node120 : node1;
		assign node1 = (inp[0]) ? node65 : node2;
			assign node2 = (inp[7]) ? node32 : node3;
				assign node3 = (inp[5]) ? node17 : node4;
					assign node4 = (inp[8]) ? node6 : 5'b11011;
						assign node6 = (inp[3]) ? node12 : node7;
							assign node7 = (inp[1]) ? 5'b11000 : node8;
								assign node8 = (inp[4]) ? 5'b10001 : 5'b01001;
							assign node12 = (inp[6]) ? node14 : 5'b10001;
								assign node14 = (inp[1]) ? 5'b00001 : 5'b10001;
					assign node17 = (inp[3]) ? node23 : node18;
						assign node18 = (inp[8]) ? 5'b10000 : node19;
							assign node19 = (inp[6]) ? 5'b01010 : 5'b10010;
						assign node23 = (inp[8]) ? node27 : node24;
							assign node24 = (inp[4]) ? 5'b11010 : 5'b01011;
							assign node27 = (inp[1]) ? node29 : 5'b01111;
								assign node29 = (inp[6]) ? 5'b01110 : 5'b11110;
				assign node32 = (inp[5]) ? node50 : node33;
					assign node33 = (inp[3]) ? node45 : node34;
						assign node34 = (inp[8]) ? node38 : node35;
							assign node35 = (inp[1]) ? 5'b10111 : 5'b01110;
							assign node38 = (inp[6]) ? node40 : 5'b00000;
								assign node40 = (inp[4]) ? node42 : 5'b00000;
									assign node42 = (inp[1]) ? 5'b01111 : 5'b11111;
						assign node45 = (inp[6]) ? node47 : 5'b01111;
							assign node47 = (inp[1]) ? 5'b01110 : 5'b11110;
					assign node50 = (inp[8]) ? node60 : node51;
						assign node51 = (inp[4]) ? 5'b00110 : node52;
							assign node52 = (inp[6]) ? node56 : node53;
								assign node53 = (inp[3]) ? 5'b10110 : 5'b11011;
								assign node56 = (inp[1]) ? 5'b00110 : 5'b10110;
						assign node60 = (inp[1]) ? 5'b10111 : node61;
							assign node61 = (inp[6]) ? 5'b11110 : 5'b01111;
			assign node65 = (inp[7]) ? node93 : node66;
				assign node66 = (inp[8]) ? node74 : node67;
					assign node67 = (inp[5]) ? 5'b00010 : node68;
						assign node68 = (inp[1]) ? node70 : 5'b00011;
							assign node70 = (inp[3]) ? 5'b10010 : 5'b00010;
					assign node74 = (inp[6]) ? node84 : node75;
						assign node75 = (inp[1]) ? node79 : node76;
							assign node76 = (inp[5]) ? 5'b00110 : 5'b01110;
							assign node79 = (inp[4]) ? 5'b11011 : node80;
								assign node80 = (inp[5]) ? 5'b10110 : 5'b11110;
						assign node84 = (inp[1]) ? node88 : node85;
							assign node85 = (inp[5]) ? 5'b10110 : 5'b10111;
							assign node88 = (inp[3]) ? node90 : 5'b00110;
								assign node90 = (inp[5]) ? 5'b01011 : 5'b00110;
				assign node93 = (inp[5]) ? node103 : node94;
					assign node94 = (inp[3]) ? node100 : node95;
						assign node95 = (inp[4]) ? 5'b10011 : node96;
							assign node96 = (inp[1]) ? 5'b10011 : 5'b11010;
						assign node100 = (inp[1]) ? 5'b01010 : 5'b11011;
					assign node103 = (inp[3]) ? node115 : node104;
						assign node104 = (inp[1]) ? node112 : node105;
							assign node105 = (inp[6]) ? node109 : node106;
								assign node106 = (inp[8]) ? 5'b01010 : 5'b00010;
								assign node109 = (inp[4]) ? 5'b10011 : 5'b10010;
							assign node112 = (inp[6]) ? 5'b00011 : 5'b10011;
						assign node115 = (inp[8]) ? 5'b10010 : node116;
							assign node116 = (inp[6]) ? 5'b10011 : 5'b10010;
		assign node120 = (inp[0]) ? node166 : node121;
			assign node121 = (inp[8]) ? node149 : node122;
				assign node122 = (inp[7]) ? node136 : node123;
					assign node123 = (inp[3]) ? node129 : node124;
						assign node124 = (inp[1]) ? node126 : 5'b01000;
							assign node126 = (inp[4]) ? 5'b11000 : 5'b11001;
						assign node129 = (inp[5]) ? node133 : node130;
							assign node130 = (inp[1]) ? 5'b00100 : 5'b00101;
							assign node133 = (inp[4]) ? 5'b01000 : 5'b01001;
					assign node136 = (inp[4]) ? 5'b11001 : node137;
						assign node137 = (inp[5]) ? 5'b10100 : node138;
							assign node138 = (inp[3]) ? node142 : node139;
								assign node139 = (inp[6]) ? 5'b01100 : 5'b10101;
								assign node142 = (inp[6]) ? node144 : 5'b01101;
									assign node144 = (inp[1]) ? 5'b01101 : 5'b11101;
				assign node149 = (inp[7]) ? node157 : node150;
					assign node150 = (inp[5]) ? node152 : 5'b11101;
						assign node152 = (inp[3]) ? node154 : 5'b11101;
							assign node154 = (inp[4]) ? 5'b11100 : 5'b11101;
					assign node157 = (inp[3]) ? node163 : node158;
						assign node158 = (inp[4]) ? node160 : 5'b11100;
							assign node160 = (inp[1]) ? 5'b00101 : 5'b10101;
						assign node163 = (inp[5]) ? 5'b10100 : 5'b11100;
			assign node166 = (inp[3]) ? node196 : node167;
				assign node167 = (inp[6]) ? node183 : node168;
					assign node168 = (inp[8]) ? node174 : node169;
						assign node169 = (inp[4]) ? node171 : 5'b11111;
							assign node171 = (inp[1]) ? 5'b10110 : 5'b00111;
						assign node174 = (inp[4]) ? node180 : node175;
							assign node175 = (inp[5]) ? 5'b00101 : node176;
								assign node176 = (inp[7]) ? 5'b00101 : 5'b01101;
							assign node180 = (inp[7]) ? 5'b00100 : 5'b01100;
					assign node183 = (inp[1]) ? node193 : node184;
						assign node184 = (inp[4]) ? node190 : node185;
							assign node185 = (inp[5]) ? 5'b11000 : node186;
								assign node186 = (inp[7]) ? 5'b10100 : 5'b11100;
							assign node190 = (inp[5]) ? 5'b10001 : 5'b10101;
						assign node193 = (inp[8]) ? 5'b00100 : 5'b00000;
				assign node196 = (inp[1]) ? node208 : node197;
					assign node197 = (inp[6]) ? node205 : node198;
						assign node198 = (inp[8]) ? node202 : node199;
							assign node199 = (inp[4]) ? 5'b01110 : 5'b01111;
							assign node202 = (inp[4]) ? 5'b01001 : 5'b01100;
						assign node205 = (inp[7]) ? 5'b11001 : 5'b11000;
					assign node208 = (inp[6]) ? node216 : node209;
						assign node209 = (inp[7]) ? 5'b11000 : node210;
							assign node210 = (inp[5]) ? 5'b11000 : node211;
								assign node211 = (inp[4]) ? 5'b10100 : 5'b10000;
						assign node216 = (inp[5]) ? 5'b00001 : node217;
							assign node217 = (inp[7]) ? 5'b01000 : 5'b00000;

endmodule