module dtc_split25_bm88 (
	input  wire [12-1:0] inp,
	output wire [3-1:0] outp
);

	wire [3-1:0] node1;
	wire [3-1:0] node2;
	wire [3-1:0] node3;
	wire [3-1:0] node4;
	wire [3-1:0] node5;
	wire [3-1:0] node6;
	wire [3-1:0] node8;
	wire [3-1:0] node11;
	wire [3-1:0] node12;
	wire [3-1:0] node14;
	wire [3-1:0] node17;
	wire [3-1:0] node20;
	wire [3-1:0] node21;
	wire [3-1:0] node22;
	wire [3-1:0] node25;
	wire [3-1:0] node27;
	wire [3-1:0] node28;
	wire [3-1:0] node33;
	wire [3-1:0] node34;
	wire [3-1:0] node36;
	wire [3-1:0] node38;
	wire [3-1:0] node42;
	wire [3-1:0] node43;
	wire [3-1:0] node44;
	wire [3-1:0] node45;
	wire [3-1:0] node46;
	wire [3-1:0] node47;
	wire [3-1:0] node48;
	wire [3-1:0] node52;
	wire [3-1:0] node53;
	wire [3-1:0] node57;
	wire [3-1:0] node58;
	wire [3-1:0] node59;
	wire [3-1:0] node63;
	wire [3-1:0] node64;
	wire [3-1:0] node68;
	wire [3-1:0] node69;
	wire [3-1:0] node72;
	wire [3-1:0] node73;
	wire [3-1:0] node75;
	wire [3-1:0] node79;
	wire [3-1:0] node80;
	wire [3-1:0] node81;
	wire [3-1:0] node82;
	wire [3-1:0] node83;
	wire [3-1:0] node87;
	wire [3-1:0] node88;
	wire [3-1:0] node92;
	wire [3-1:0] node93;
	wire [3-1:0] node94;
	wire [3-1:0] node98;
	wire [3-1:0] node99;
	wire [3-1:0] node103;
	wire [3-1:0] node104;
	wire [3-1:0] node105;
	wire [3-1:0] node107;
	wire [3-1:0] node110;
	wire [3-1:0] node113;
	wire [3-1:0] node114;
	wire [3-1:0] node115;
	wire [3-1:0] node118;
	wire [3-1:0] node121;
	wire [3-1:0] node124;
	wire [3-1:0] node126;
	wire [3-1:0] node127;
	wire [3-1:0] node128;
	wire [3-1:0] node129;
	wire [3-1:0] node132;
	wire [3-1:0] node135;
	wire [3-1:0] node137;
	wire [3-1:0] node138;
	wire [3-1:0] node142;
	wire [3-1:0] node144;
	wire [3-1:0] node146;
	wire [3-1:0] node149;
	wire [3-1:0] node150;
	wire [3-1:0] node151;
	wire [3-1:0] node152;
	wire [3-1:0] node153;
	wire [3-1:0] node155;
	wire [3-1:0] node161;
	wire [3-1:0] node162;
	wire [3-1:0] node163;
	wire [3-1:0] node165;
	wire [3-1:0] node166;
	wire [3-1:0] node167;
	wire [3-1:0] node171;
	wire [3-1:0] node172;
	wire [3-1:0] node173;
	wire [3-1:0] node178;
	wire [3-1:0] node179;
	wire [3-1:0] node181;
	wire [3-1:0] node183;
	wire [3-1:0] node185;
	wire [3-1:0] node188;
	wire [3-1:0] node189;
	wire [3-1:0] node190;
	wire [3-1:0] node191;
	wire [3-1:0] node196;
	wire [3-1:0] node197;
	wire [3-1:0] node200;
	wire [3-1:0] node203;
	wire [3-1:0] node204;
	wire [3-1:0] node205;
	wire [3-1:0] node206;
	wire [3-1:0] node207;
	wire [3-1:0] node208;
	wire [3-1:0] node215;
	wire [3-1:0] node217;
	wire [3-1:0] node218;
	wire [3-1:0] node222;
	wire [3-1:0] node223;
	wire [3-1:0] node224;
	wire [3-1:0] node225;
	wire [3-1:0] node226;
	wire [3-1:0] node228;
	wire [3-1:0] node230;
	wire [3-1:0] node231;
	wire [3-1:0] node236;
	wire [3-1:0] node237;
	wire [3-1:0] node238;
	wire [3-1:0] node239;
	wire [3-1:0] node241;
	wire [3-1:0] node242;
	wire [3-1:0] node245;
	wire [3-1:0] node248;
	wire [3-1:0] node249;
	wire [3-1:0] node251;
	wire [3-1:0] node254;
	wire [3-1:0] node256;
	wire [3-1:0] node259;
	wire [3-1:0] node260;
	wire [3-1:0] node261;
	wire [3-1:0] node265;
	wire [3-1:0] node266;
	wire [3-1:0] node269;
	wire [3-1:0] node272;
	wire [3-1:0] node273;
	wire [3-1:0] node274;
	wire [3-1:0] node277;
	wire [3-1:0] node279;
	wire [3-1:0] node282;
	wire [3-1:0] node284;
	wire [3-1:0] node285;
	wire [3-1:0] node289;
	wire [3-1:0] node290;
	wire [3-1:0] node291;
	wire [3-1:0] node293;
	wire [3-1:0] node294;
	wire [3-1:0] node297;
	wire [3-1:0] node299;
	wire [3-1:0] node301;
	wire [3-1:0] node304;
	wire [3-1:0] node305;
	wire [3-1:0] node306;
	wire [3-1:0] node307;
	wire [3-1:0] node309;
	wire [3-1:0] node313;
	wire [3-1:0] node314;
	wire [3-1:0] node317;
	wire [3-1:0] node318;
	wire [3-1:0] node322;
	wire [3-1:0] node323;
	wire [3-1:0] node324;
	wire [3-1:0] node326;
	wire [3-1:0] node329;
	wire [3-1:0] node330;
	wire [3-1:0] node334;
	wire [3-1:0] node335;
	wire [3-1:0] node337;
	wire [3-1:0] node340;
	wire [3-1:0] node341;
	wire [3-1:0] node344;
	wire [3-1:0] node347;
	wire [3-1:0] node348;
	wire [3-1:0] node349;
	wire [3-1:0] node350;
	wire [3-1:0] node351;
	wire [3-1:0] node353;
	wire [3-1:0] node357;
	wire [3-1:0] node358;
	wire [3-1:0] node359;
	wire [3-1:0] node362;
	wire [3-1:0] node365;
	wire [3-1:0] node367;
	wire [3-1:0] node370;
	wire [3-1:0] node371;
	wire [3-1:0] node374;
	wire [3-1:0] node375;
	wire [3-1:0] node377;
	wire [3-1:0] node381;
	wire [3-1:0] node382;
	wire [3-1:0] node383;
	wire [3-1:0] node385;
	wire [3-1:0] node386;
	wire [3-1:0] node390;
	wire [3-1:0] node391;
	wire [3-1:0] node392;
	wire [3-1:0] node397;
	wire [3-1:0] node398;
	wire [3-1:0] node400;
	wire [3-1:0] node401;
	wire [3-1:0] node405;
	wire [3-1:0] node406;
	wire [3-1:0] node407;
	wire [3-1:0] node410;
	wire [3-1:0] node413;
	wire [3-1:0] node415;
	wire [3-1:0] node418;
	wire [3-1:0] node419;
	wire [3-1:0] node420;
	wire [3-1:0] node421;
	wire [3-1:0] node422;
	wire [3-1:0] node423;
	wire [3-1:0] node424;
	wire [3-1:0] node428;
	wire [3-1:0] node429;
	wire [3-1:0] node432;
	wire [3-1:0] node434;
	wire [3-1:0] node437;
	wire [3-1:0] node439;
	wire [3-1:0] node440;
	wire [3-1:0] node443;
	wire [3-1:0] node445;
	wire [3-1:0] node448;
	wire [3-1:0] node449;
	wire [3-1:0] node450;
	wire [3-1:0] node451;
	wire [3-1:0] node453;
	wire [3-1:0] node456;
	wire [3-1:0] node458;
	wire [3-1:0] node461;
	wire [3-1:0] node464;
	wire [3-1:0] node465;
	wire [3-1:0] node466;
	wire [3-1:0] node467;
	wire [3-1:0] node471;
	wire [3-1:0] node472;
	wire [3-1:0] node475;
	wire [3-1:0] node478;
	wire [3-1:0] node481;
	wire [3-1:0] node482;
	wire [3-1:0] node483;
	wire [3-1:0] node484;
	wire [3-1:0] node485;
	wire [3-1:0] node488;
	wire [3-1:0] node491;
	wire [3-1:0] node492;
	wire [3-1:0] node495;
	wire [3-1:0] node498;
	wire [3-1:0] node499;
	wire [3-1:0] node502;
	wire [3-1:0] node504;
	wire [3-1:0] node507;
	wire [3-1:0] node508;
	wire [3-1:0] node509;
	wire [3-1:0] node514;
	wire [3-1:0] node515;
	wire [3-1:0] node516;
	wire [3-1:0] node517;
	wire [3-1:0] node518;
	wire [3-1:0] node519;
	wire [3-1:0] node521;
	wire [3-1:0] node524;
	wire [3-1:0] node525;
	wire [3-1:0] node529;
	wire [3-1:0] node530;
	wire [3-1:0] node532;
	wire [3-1:0] node535;
	wire [3-1:0] node536;
	wire [3-1:0] node540;
	wire [3-1:0] node541;
	wire [3-1:0] node542;
	wire [3-1:0] node544;
	wire [3-1:0] node547;
	wire [3-1:0] node549;
	wire [3-1:0] node552;
	wire [3-1:0] node553;
	wire [3-1:0] node554;
	wire [3-1:0] node557;
	wire [3-1:0] node561;
	wire [3-1:0] node562;
	wire [3-1:0] node563;
	wire [3-1:0] node564;
	wire [3-1:0] node567;
	wire [3-1:0] node568;
	wire [3-1:0] node572;
	wire [3-1:0] node573;
	wire [3-1:0] node574;
	wire [3-1:0] node578;
	wire [3-1:0] node580;
	wire [3-1:0] node583;
	wire [3-1:0] node584;
	wire [3-1:0] node585;
	wire [3-1:0] node586;
	wire [3-1:0] node590;
	wire [3-1:0] node594;
	wire [3-1:0] node595;
	wire [3-1:0] node596;
	wire [3-1:0] node597;
	wire [3-1:0] node598;
	wire [3-1:0] node599;
	wire [3-1:0] node602;
	wire [3-1:0] node605;
	wire [3-1:0] node608;
	wire [3-1:0] node609;
	wire [3-1:0] node610;
	wire [3-1:0] node613;
	wire [3-1:0] node616;
	wire [3-1:0] node619;
	wire [3-1:0] node620;
	wire [3-1:0] node621;
	wire [3-1:0] node623;
	wire [3-1:0] node626;
	wire [3-1:0] node629;
	wire [3-1:0] node630;
	wire [3-1:0] node631;
	wire [3-1:0] node635;
	wire [3-1:0] node637;
	wire [3-1:0] node640;
	wire [3-1:0] node641;
	wire [3-1:0] node642;
	wire [3-1:0] node643;
	wire [3-1:0] node645;
	wire [3-1:0] node648;
	wire [3-1:0] node649;
	wire [3-1:0] node654;
	wire [3-1:0] node655;
	wire [3-1:0] node656;
	wire [3-1:0] node659;
	wire [3-1:0] node662;
	wire [3-1:0] node663;
	wire [3-1:0] node665;
	wire [3-1:0] node668;
	wire [3-1:0] node669;

	assign outp = (inp[6]) ? node222 : node1;
		assign node1 = (inp[3]) ? node149 : node2;
			assign node2 = (inp[0]) ? node42 : node3;
				assign node3 = (inp[9]) ? node33 : node4;
					assign node4 = (inp[7]) ? node20 : node5;
						assign node5 = (inp[5]) ? node11 : node6;
							assign node6 = (inp[10]) ? node8 : 3'b000;
								assign node8 = (inp[8]) ? 3'b000 : 3'b010;
							assign node11 = (inp[8]) ? node17 : node12;
								assign node12 = (inp[10]) ? node14 : 3'b010;
									assign node14 = (inp[11]) ? 3'b110 : 3'b100;
								assign node17 = (inp[10]) ? 3'b010 : 3'b000;
						assign node20 = (inp[8]) ? 3'b000 : node21;
							assign node21 = (inp[4]) ? node25 : node22;
								assign node22 = (inp[5]) ? 3'b010 : 3'b000;
								assign node25 = (inp[5]) ? node27 : 3'b000;
									assign node27 = (inp[11]) ? 3'b000 : node28;
										assign node28 = (inp[10]) ? 3'b000 : 3'b010;
					assign node33 = (inp[8]) ? 3'b000 : node34;
						assign node34 = (inp[10]) ? node36 : 3'b000;
							assign node36 = (inp[7]) ? node38 : 3'b000;
								assign node38 = (inp[5]) ? 3'b010 : 3'b000;
				assign node42 = (inp[9]) ? node124 : node43;
					assign node43 = (inp[8]) ? node79 : node44;
						assign node44 = (inp[5]) ? node68 : node45;
							assign node45 = (inp[7]) ? node57 : node46;
								assign node46 = (inp[10]) ? node52 : node47;
									assign node47 = (inp[11]) ? 3'b010 : node48;
										assign node48 = (inp[4]) ? 3'b100 : 3'b110;
									assign node52 = (inp[2]) ? 3'b000 : node53;
										assign node53 = (inp[1]) ? 3'b010 : 3'b000;
								assign node57 = (inp[4]) ? node63 : node58;
									assign node58 = (inp[1]) ? 3'b001 : node59;
										assign node59 = (inp[2]) ? 3'b100 : 3'b000;
									assign node63 = (inp[11]) ? 3'b010 : node64;
										assign node64 = (inp[2]) ? 3'b010 : 3'b001;
							assign node68 = (inp[10]) ? node72 : node69;
								assign node69 = (inp[2]) ? 3'b100 : 3'b000;
								assign node72 = (inp[11]) ? 3'b000 : node73;
									assign node73 = (inp[1]) ? node75 : 3'b000;
										assign node75 = (inp[4]) ? 3'b000 : 3'b010;
						assign node79 = (inp[1]) ? node103 : node80;
							assign node80 = (inp[5]) ? node92 : node81;
								assign node81 = (inp[11]) ? node87 : node82;
									assign node82 = (inp[10]) ? 3'b000 : node83;
										assign node83 = (inp[2]) ? 3'b000 : 3'b100;
									assign node87 = (inp[10]) ? 3'b110 : node88;
										assign node88 = (inp[4]) ? 3'b000 : 3'b010;
								assign node92 = (inp[2]) ? node98 : node93;
									assign node93 = (inp[4]) ? 3'b010 : node94;
										assign node94 = (inp[10]) ? 3'b100 : 3'b000;
									assign node98 = (inp[4]) ? 3'b111 : node99;
										assign node99 = (inp[10]) ? 3'b100 : 3'b110;
							assign node103 = (inp[4]) ? node113 : node104;
								assign node104 = (inp[7]) ? node110 : node105;
									assign node105 = (inp[2]) ? node107 : 3'b010;
										assign node107 = (inp[5]) ? 3'b010 : 3'b010;
									assign node110 = (inp[10]) ? 3'b110 : 3'b100;
								assign node113 = (inp[7]) ? node121 : node114;
									assign node114 = (inp[11]) ? node118 : node115;
										assign node115 = (inp[10]) ? 3'b000 : 3'b010;
										assign node118 = (inp[10]) ? 3'b000 : 3'b100;
									assign node121 = (inp[10]) ? 3'b010 : 3'b110;
					assign node124 = (inp[7]) ? node126 : 3'b000;
						assign node126 = (inp[4]) ? node142 : node127;
							assign node127 = (inp[10]) ? node135 : node128;
								assign node128 = (inp[8]) ? node132 : node129;
									assign node129 = (inp[5]) ? 3'b100 : 3'b010;
									assign node132 = (inp[5]) ? 3'b010 : 3'b110;
								assign node135 = (inp[1]) ? node137 : 3'b110;
									assign node137 = (inp[11]) ? 3'b100 : node138;
										assign node138 = (inp[8]) ? 3'b100 : 3'b000;
							assign node142 = (inp[8]) ? node144 : 3'b000;
								assign node144 = (inp[5]) ? node146 : 3'b010;
									assign node146 = (inp[11]) ? 3'b000 : 3'b100;
			assign node149 = (inp[7]) ? node161 : node150;
				assign node150 = (inp[4]) ? 3'b000 : node151;
					assign node151 = (inp[8]) ? 3'b000 : node152;
						assign node152 = (inp[9]) ? 3'b000 : node153;
							assign node153 = (inp[1]) ? node155 : 3'b000;
								assign node155 = (inp[5]) ? 3'b000 : 3'b100;
				assign node161 = (inp[0]) ? node203 : node162;
					assign node162 = (inp[8]) ? node178 : node163;
						assign node163 = (inp[1]) ? node165 : 3'b000;
							assign node165 = (inp[5]) ? node171 : node166;
								assign node166 = (inp[9]) ? 3'b000 : node167;
									assign node167 = (inp[10]) ? 3'b010 : 3'b000;
								assign node171 = (inp[9]) ? 3'b000 : node172;
									assign node172 = (inp[2]) ? 3'b100 : node173;
										assign node173 = (inp[11]) ? 3'b000 : 3'b100;
						assign node178 = (inp[5]) ? node188 : node179;
							assign node179 = (inp[4]) ? node181 : 3'b100;
								assign node181 = (inp[11]) ? node183 : 3'b100;
									assign node183 = (inp[10]) ? node185 : 3'b000;
										assign node185 = (inp[1]) ? 3'b100 : 3'b000;
							assign node188 = (inp[1]) ? node196 : node189;
								assign node189 = (inp[4]) ? 3'b000 : node190;
									assign node190 = (inp[10]) ? 3'b000 : node191;
										assign node191 = (inp[11]) ? 3'b100 : 3'b000;
								assign node196 = (inp[4]) ? node200 : node197;
									assign node197 = (inp[10]) ? 3'b110 : 3'b010;
									assign node200 = (inp[11]) ? 3'b000 : 3'b100;
					assign node203 = (inp[9]) ? node215 : node204;
						assign node204 = (inp[4]) ? 3'b000 : node205;
							assign node205 = (inp[10]) ? 3'b000 : node206;
								assign node206 = (inp[8]) ? 3'b100 : node207;
									assign node207 = (inp[5]) ? 3'b000 : node208;
										assign node208 = (inp[1]) ? 3'b100 : 3'b000;
						assign node215 = (inp[8]) ? node217 : 3'b000;
							assign node217 = (inp[10]) ? 3'b000 : node218;
								assign node218 = (inp[11]) ? 3'b000 : 3'b010;
		assign node222 = (inp[3]) ? node418 : node223;
			assign node223 = (inp[7]) ? node289 : node224;
				assign node224 = (inp[0]) ? node236 : node225;
					assign node225 = (inp[8]) ? 3'b001 : node226;
						assign node226 = (inp[5]) ? node228 : 3'b001;
							assign node228 = (inp[2]) ? node230 : 3'b000;
								assign node230 = (inp[9]) ? 3'b000 : node231;
									assign node231 = (inp[10]) ? 3'b001 : 3'b000;
					assign node236 = (inp[10]) ? node272 : node237;
						assign node237 = (inp[11]) ? node259 : node238;
							assign node238 = (inp[9]) ? node248 : node239;
								assign node239 = (inp[4]) ? node241 : 3'b011;
									assign node241 = (inp[8]) ? node245 : node242;
										assign node242 = (inp[5]) ? 3'b010 : 3'b001;
										assign node245 = (inp[5]) ? 3'b001 : 3'b101;
								assign node248 = (inp[8]) ? node254 : node249;
									assign node249 = (inp[4]) ? node251 : 3'b101;
										assign node251 = (inp[5]) ? 3'b110 : 3'b001;
									assign node254 = (inp[4]) ? node256 : 3'b011;
										assign node256 = (inp[2]) ? 3'b101 : 3'b001;
							assign node259 = (inp[4]) ? node265 : node260;
								assign node260 = (inp[8]) ? 3'b111 : node261;
									assign node261 = (inp[5]) ? 3'b001 : 3'b111;
								assign node265 = (inp[8]) ? node269 : node266;
									assign node266 = (inp[5]) ? 3'b010 : 3'b011;
									assign node269 = (inp[5]) ? 3'b011 : 3'b111;
						assign node272 = (inp[4]) ? node282 : node273;
							assign node273 = (inp[11]) ? node277 : node274;
								assign node274 = (inp[5]) ? 3'b100 : 3'b110;
								assign node277 = (inp[1]) ? node279 : 3'b010;
									assign node279 = (inp[5]) ? 3'b010 : 3'b110;
							assign node282 = (inp[11]) ? node284 : 3'b110;
								assign node284 = (inp[8]) ? 3'b100 : node285;
									assign node285 = (inp[5]) ? 3'b110 : 3'b100;
				assign node289 = (inp[9]) ? node347 : node290;
					assign node290 = (inp[0]) ? node304 : node291;
						assign node291 = (inp[10]) ? node293 : 3'b111;
							assign node293 = (inp[8]) ? node297 : node294;
								assign node294 = (inp[2]) ? 3'b011 : 3'b000;
								assign node297 = (inp[11]) ? node299 : 3'b111;
									assign node299 = (inp[5]) ? node301 : 3'b111;
										assign node301 = (inp[1]) ? 3'b011 : 3'b111;
						assign node304 = (inp[1]) ? node322 : node305;
							assign node305 = (inp[5]) ? node313 : node306;
								assign node306 = (inp[8]) ? 3'b111 : node307;
									assign node307 = (inp[4]) ? node309 : 3'b111;
										assign node309 = (inp[2]) ? 3'b111 : 3'b011;
								assign node313 = (inp[2]) ? node317 : node314;
									assign node314 = (inp[11]) ? 3'b101 : 3'b100;
									assign node317 = (inp[10]) ? 3'b111 : node318;
										assign node318 = (inp[11]) ? 3'b001 : 3'b011;
							assign node322 = (inp[10]) ? node334 : node323;
								assign node323 = (inp[4]) ? node329 : node324;
									assign node324 = (inp[2]) ? node326 : 3'b011;
										assign node326 = (inp[11]) ? 3'b011 : 3'b011;
									assign node329 = (inp[5]) ? 3'b101 : node330;
										assign node330 = (inp[8]) ? 3'b011 : 3'b101;
								assign node334 = (inp[5]) ? node340 : node335;
									assign node335 = (inp[4]) ? node337 : 3'b101;
										assign node337 = (inp[8]) ? 3'b101 : 3'b001;
									assign node340 = (inp[11]) ? node344 : node341;
										assign node341 = (inp[8]) ? 3'b011 : 3'b010;
										assign node344 = (inp[4]) ? 3'b001 : 3'b101;
					assign node347 = (inp[4]) ? node381 : node348;
						assign node348 = (inp[5]) ? node370 : node349;
							assign node349 = (inp[10]) ? node357 : node350;
								assign node350 = (inp[11]) ? 3'b111 : node351;
									assign node351 = (inp[0]) ? node353 : 3'b011;
										assign node353 = (inp[1]) ? 3'b011 : 3'b111;
								assign node357 = (inp[8]) ? node365 : node358;
									assign node358 = (inp[1]) ? node362 : node359;
										assign node359 = (inp[0]) ? 3'b101 : 3'b111;
										assign node362 = (inp[0]) ? 3'b110 : 3'b011;
									assign node365 = (inp[11]) ? node367 : 3'b101;
										assign node367 = (inp[0]) ? 3'b001 : 3'b011;
							assign node370 = (inp[0]) ? node374 : node371;
								assign node371 = (inp[8]) ? 3'b111 : 3'b000;
								assign node374 = (inp[10]) ? 3'b110 : node375;
									assign node375 = (inp[8]) ? node377 : 3'b111;
										assign node377 = (inp[1]) ? 3'b110 : 3'b011;
						assign node381 = (inp[5]) ? node397 : node382;
							assign node382 = (inp[0]) ? node390 : node383;
								assign node383 = (inp[1]) ? node385 : 3'b111;
									assign node385 = (inp[10]) ? 3'b101 : node386;
										assign node386 = (inp[11]) ? 3'b101 : 3'b011;
								assign node390 = (inp[2]) ? 3'b001 : node391;
									assign node391 = (inp[10]) ? 3'b101 : node392;
										assign node392 = (inp[8]) ? 3'b001 : 3'b101;
							assign node397 = (inp[8]) ? node405 : node398;
								assign node398 = (inp[0]) ? node400 : 3'b000;
									assign node400 = (inp[11]) ? 3'b100 : node401;
										assign node401 = (inp[2]) ? 3'b101 : 3'b111;
								assign node405 = (inp[0]) ? node413 : node406;
									assign node406 = (inp[1]) ? node410 : node407;
										assign node407 = (inp[2]) ? 3'b011 : 3'b111;
										assign node410 = (inp[2]) ? 3'b101 : 3'b001;
									assign node413 = (inp[11]) ? node415 : 3'b001;
										assign node415 = (inp[2]) ? 3'b110 : 3'b010;
			assign node418 = (inp[7]) ? node514 : node419;
				assign node419 = (inp[9]) ? node481 : node420;
					assign node420 = (inp[5]) ? node448 : node421;
						assign node421 = (inp[8]) ? node437 : node422;
							assign node422 = (inp[0]) ? node428 : node423;
								assign node423 = (inp[11]) ? 3'b100 : node424;
									assign node424 = (inp[10]) ? 3'b010 : 3'b110;
								assign node428 = (inp[1]) ? node432 : node429;
									assign node429 = (inp[10]) ? 3'b100 : 3'b010;
									assign node432 = (inp[10]) ? node434 : 3'b100;
										assign node434 = (inp[2]) ? 3'b000 : 3'b100;
							assign node437 = (inp[0]) ? node439 : 3'b000;
								assign node439 = (inp[4]) ? node443 : node440;
									assign node440 = (inp[10]) ? 3'b010 : 3'b110;
									assign node443 = (inp[11]) ? node445 : 3'b000;
										assign node445 = (inp[1]) ? 3'b100 : 3'b000;
						assign node448 = (inp[10]) ? node464 : node449;
							assign node449 = (inp[8]) ? node461 : node450;
								assign node450 = (inp[0]) ? node456 : node451;
									assign node451 = (inp[1]) ? node453 : 3'b000;
										assign node453 = (inp[2]) ? 3'b000 : 3'b010;
									assign node456 = (inp[1]) ? node458 : 3'b100;
										assign node458 = (inp[4]) ? 3'b000 : 3'b100;
								assign node461 = (inp[11]) ? 3'b010 : 3'b110;
							assign node464 = (inp[0]) ? node478 : node465;
								assign node465 = (inp[4]) ? node471 : node466;
									assign node466 = (inp[1]) ? 3'b100 : node467;
										assign node467 = (inp[8]) ? 3'b100 : 3'b110;
									assign node471 = (inp[8]) ? node475 : node472;
										assign node472 = (inp[11]) ? 3'b110 : 3'b100;
										assign node475 = (inp[11]) ? 3'b100 : 3'b010;
								assign node478 = (inp[4]) ? 3'b000 : 3'b100;
					assign node481 = (inp[0]) ? node507 : node482;
						assign node482 = (inp[10]) ? node498 : node483;
							assign node483 = (inp[11]) ? node491 : node484;
								assign node484 = (inp[5]) ? node488 : node485;
									assign node485 = (inp[8]) ? 3'b000 : 3'b110;
									assign node488 = (inp[8]) ? 3'b110 : 3'b000;
								assign node491 = (inp[8]) ? node495 : node492;
									assign node492 = (inp[5]) ? 3'b000 : 3'b010;
									assign node495 = (inp[5]) ? 3'b010 : 3'b000;
							assign node498 = (inp[5]) ? node502 : node499;
								assign node499 = (inp[8]) ? 3'b000 : 3'b010;
								assign node502 = (inp[8]) ? node504 : 3'b100;
									assign node504 = (inp[11]) ? 3'b100 : 3'b010;
						assign node507 = (inp[4]) ? 3'b000 : node508;
							assign node508 = (inp[10]) ? 3'b000 : node509;
								assign node509 = (inp[8]) ? 3'b000 : 3'b010;
				assign node514 = (inp[0]) ? node594 : node515;
					assign node515 = (inp[10]) ? node561 : node516;
						assign node516 = (inp[9]) ? node540 : node517;
							assign node517 = (inp[4]) ? node529 : node518;
								assign node518 = (inp[5]) ? node524 : node519;
									assign node519 = (inp[1]) ? node521 : 3'b111;
										assign node521 = (inp[8]) ? 3'b111 : 3'b011;
									assign node524 = (inp[11]) ? 3'b111 : node525;
										assign node525 = (inp[8]) ? 3'b011 : 3'b000;
								assign node529 = (inp[5]) ? node535 : node530;
									assign node530 = (inp[11]) ? node532 : 3'b011;
										assign node532 = (inp[2]) ? 3'b001 : 3'b001;
									assign node535 = (inp[11]) ? 3'b110 : node536;
										assign node536 = (inp[2]) ? 3'b101 : 3'b000;
							assign node540 = (inp[5]) ? node552 : node541;
								assign node541 = (inp[11]) ? node547 : node542;
									assign node542 = (inp[8]) ? node544 : 3'b001;
										assign node544 = (inp[4]) ? 3'b001 : 3'b011;
									assign node547 = (inp[2]) ? node549 : 3'b001;
										assign node549 = (inp[1]) ? 3'b001 : 3'b000;
								assign node552 = (inp[4]) ? 3'b110 : node553;
									assign node553 = (inp[8]) ? node557 : node554;
										assign node554 = (inp[11]) ? 3'b110 : 3'b000;
										assign node557 = (inp[1]) ? 3'b001 : 3'b101;
						assign node561 = (inp[5]) ? node583 : node562;
							assign node562 = (inp[9]) ? node572 : node563;
								assign node563 = (inp[8]) ? node567 : node564;
									assign node564 = (inp[1]) ? 3'b001 : 3'b011;
									assign node567 = (inp[11]) ? 3'b101 : node568;
										assign node568 = (inp[4]) ? 3'b101 : 3'b011;
								assign node572 = (inp[4]) ? node578 : node573;
									assign node573 = (inp[11]) ? 3'b001 : node574;
										assign node574 = (inp[8]) ? 3'b101 : 3'b110;
									assign node578 = (inp[1]) ? node580 : 3'b110;
										assign node580 = (inp[2]) ? 3'b100 : 3'b010;
							assign node583 = (inp[9]) ? 3'b110 : node584;
								assign node584 = (inp[8]) ? node590 : node585;
									assign node585 = (inp[2]) ? 3'b110 : node586;
										assign node586 = (inp[4]) ? 3'b110 : 3'b111;
									assign node590 = (inp[11]) ? 3'b001 : 3'b101;
					assign node594 = (inp[9]) ? node640 : node595;
						assign node595 = (inp[5]) ? node619 : node596;
							assign node596 = (inp[10]) ? node608 : node597;
								assign node597 = (inp[4]) ? node605 : node598;
									assign node598 = (inp[1]) ? node602 : node599;
										assign node599 = (inp[8]) ? 3'b011 : 3'b101;
										assign node602 = (inp[8]) ? 3'b001 : 3'b001;
									assign node605 = (inp[1]) ? 3'b110 : 3'b001;
								assign node608 = (inp[11]) ? node616 : node609;
									assign node609 = (inp[4]) ? node613 : node610;
										assign node610 = (inp[1]) ? 3'b001 : 3'b101;
										assign node613 = (inp[8]) ? 3'b010 : 3'b110;
									assign node616 = (inp[8]) ? 3'b110 : 3'b100;
							assign node619 = (inp[11]) ? node629 : node620;
								assign node620 = (inp[10]) ? node626 : node621;
									assign node621 = (inp[1]) ? node623 : 3'b110;
										assign node623 = (inp[4]) ? 3'b010 : 3'b110;
									assign node626 = (inp[4]) ? 3'b100 : 3'b110;
								assign node629 = (inp[2]) ? node635 : node630;
									assign node630 = (inp[8]) ? 3'b110 : node631;
										assign node631 = (inp[1]) ? 3'b010 : 3'b010;
									assign node635 = (inp[4]) ? node637 : 3'b001;
										assign node637 = (inp[8]) ? 3'b010 : 3'b000;
						assign node640 = (inp[8]) ? node654 : node641;
							assign node641 = (inp[5]) ? 3'b000 : node642;
								assign node642 = (inp[4]) ? node648 : node643;
									assign node643 = (inp[1]) ? node645 : 3'b010;
										assign node645 = (inp[10]) ? 3'b100 : 3'b010;
									assign node648 = (inp[11]) ? 3'b000 : node649;
										assign node649 = (inp[2]) ? 3'b100 : 3'b000;
							assign node654 = (inp[4]) ? node662 : node655;
								assign node655 = (inp[11]) ? node659 : node656;
									assign node656 = (inp[10]) ? 3'b010 : 3'b110;
									assign node659 = (inp[1]) ? 3'b100 : 3'b001;
								assign node662 = (inp[11]) ? node668 : node663;
									assign node663 = (inp[10]) ? node665 : 3'b100;
										assign node665 = (inp[5]) ? 3'b100 : 3'b000;
									assign node668 = (inp[1]) ? 3'b100 : node669;
										assign node669 = (inp[10]) ? 3'b100 : 3'b010;

endmodule