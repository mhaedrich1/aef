module dtc_split66_bm95 (
	input  wire [11-1:0] inp,
	output wire [3-1:0] outp
);

	wire [3-1:0] node2;
	wire [3-1:0] node3;
	wire [3-1:0] node4;
	wire [3-1:0] node5;
	wire [3-1:0] node7;
	wire [3-1:0] node8;
	wire [3-1:0] node9;
	wire [3-1:0] node10;
	wire [3-1:0] node11;
	wire [3-1:0] node14;
	wire [3-1:0] node17;
	wire [3-1:0] node18;
	wire [3-1:0] node21;
	wire [3-1:0] node24;
	wire [3-1:0] node25;
	wire [3-1:0] node28;
	wire [3-1:0] node31;
	wire [3-1:0] node33;
	wire [3-1:0] node34;
	wire [3-1:0] node35;
	wire [3-1:0] node38;
	wire [3-1:0] node41;
	wire [3-1:0] node42;
	wire [3-1:0] node44;
	wire [3-1:0] node47;
	wire [3-1:0] node48;
	wire [3-1:0] node53;
	wire [3-1:0] node55;
	wire [3-1:0] node57;
	wire [3-1:0] node58;
	wire [3-1:0] node59;
	wire [3-1:0] node60;
	wire [3-1:0] node63;
	wire [3-1:0] node66;
	wire [3-1:0] node67;
	wire [3-1:0] node68;
	wire [3-1:0] node69;
	wire [3-1:0] node73;
	wire [3-1:0] node74;
	wire [3-1:0] node77;
	wire [3-1:0] node80;
	wire [3-1:0] node82;
	wire [3-1:0] node85;
	wire [3-1:0] node87;
	wire [3-1:0] node88;
	wire [3-1:0] node89;
	wire [3-1:0] node92;
	wire [3-1:0] node95;
	wire [3-1:0] node97;
	wire [3-1:0] node100;
	wire [3-1:0] node101;
	wire [3-1:0] node102;
	wire [3-1:0] node104;
	wire [3-1:0] node105;
	wire [3-1:0] node106;
	wire [3-1:0] node107;
	wire [3-1:0] node108;
	wire [3-1:0] node109;
	wire [3-1:0] node113;
	wire [3-1:0] node116;
	wire [3-1:0] node117;
	wire [3-1:0] node121;
	wire [3-1:0] node122;
	wire [3-1:0] node123;
	wire [3-1:0] node124;
	wire [3-1:0] node127;
	wire [3-1:0] node130;
	wire [3-1:0] node132;
	wire [3-1:0] node135;
	wire [3-1:0] node136;
	wire [3-1:0] node140;
	wire [3-1:0] node141;
	wire [3-1:0] node142;
	wire [3-1:0] node143;
	wire [3-1:0] node147;
	wire [3-1:0] node150;
	wire [3-1:0] node153;
	wire [3-1:0] node154;
	wire [3-1:0] node155;
	wire [3-1:0] node156;
	wire [3-1:0] node157;
	wire [3-1:0] node160;
	wire [3-1:0] node163;
	wire [3-1:0] node164;
	wire [3-1:0] node165;
	wire [3-1:0] node166;
	wire [3-1:0] node170;
	wire [3-1:0] node171;
	wire [3-1:0] node175;
	wire [3-1:0] node176;
	wire [3-1:0] node180;
	wire [3-1:0] node182;
	wire [3-1:0] node183;
	wire [3-1:0] node185;
	wire [3-1:0] node188;
	wire [3-1:0] node190;
	wire [3-1:0] node193;
	wire [3-1:0] node194;
	wire [3-1:0] node195;
	wire [3-1:0] node196;
	wire [3-1:0] node199;
	wire [3-1:0] node202;
	wire [3-1:0] node203;
	wire [3-1:0] node207;
	wire [3-1:0] node208;
	wire [3-1:0] node209;
	wire [3-1:0] node212;
	wire [3-1:0] node215;
	wire [3-1:0] node216;
	wire [3-1:0] node220;
	wire [3-1:0] node222;
	wire [3-1:0] node223;
	wire [3-1:0] node224;
	wire [3-1:0] node225;
	wire [3-1:0] node228;
	wire [3-1:0] node231;
	wire [3-1:0] node232;
	wire [3-1:0] node234;
	wire [3-1:0] node238;
	wire [3-1:0] node240;
	wire [3-1:0] node241;
	wire [3-1:0] node243;
	wire [3-1:0] node245;
	wire [3-1:0] node248;
	wire [3-1:0] node249;
	wire [3-1:0] node250;

	assign outp = (inp[5]) ? node2 : 3'b000;
		assign node2 = (inp[8]) ? node100 : node3;
			assign node3 = (inp[6]) ? node53 : node4;
				assign node4 = (inp[0]) ? 3'b001 : node5;
					assign node5 = (inp[9]) ? node7 : 3'b011;
						assign node7 = (inp[1]) ? node31 : node8;
							assign node8 = (inp[7]) ? node24 : node9;
								assign node9 = (inp[4]) ? node17 : node10;
									assign node10 = (inp[2]) ? node14 : node11;
										assign node11 = (inp[10]) ? 3'b001 : 3'b101;
										assign node14 = (inp[10]) ? 3'b101 : 3'b001;
									assign node17 = (inp[10]) ? node21 : node18;
										assign node18 = (inp[2]) ? 3'b001 : 3'b101;
										assign node21 = (inp[2]) ? 3'b101 : 3'b001;
								assign node24 = (inp[2]) ? node28 : node25;
									assign node25 = (inp[10]) ? 3'b101 : 3'b011;
									assign node28 = (inp[10]) ? 3'b011 : 3'b101;
							assign node31 = (inp[7]) ? node33 : 3'b001;
								assign node33 = (inp[4]) ? node41 : node34;
									assign node34 = (inp[10]) ? node38 : node35;
										assign node35 = (inp[2]) ? 3'b001 : 3'b101;
										assign node38 = (inp[2]) ? 3'b101 : 3'b001;
									assign node41 = (inp[3]) ? node47 : node42;
										assign node42 = (inp[2]) ? node44 : 3'b001;
											assign node44 = (inp[10]) ? 3'b101 : 3'b001;
										assign node47 = (inp[10]) ? 3'b001 : node48;
											assign node48 = (inp[2]) ? 3'b001 : 3'b101;
				assign node53 = (inp[0]) ? node55 : 3'b111;
					assign node55 = (inp[9]) ? node57 : 3'b110;
						assign node57 = (inp[1]) ? node85 : node58;
							assign node58 = (inp[2]) ? node66 : node59;
								assign node59 = (inp[7]) ? node63 : node60;
									assign node60 = (inp[10]) ? 3'b110 : 3'b001;
									assign node63 = (inp[10]) ? 3'b001 : 3'b110;
								assign node66 = (inp[3]) ? node80 : node67;
									assign node67 = (inp[4]) ? node73 : node68;
										assign node68 = (inp[10]) ? 3'b001 : node69;
											assign node69 = (inp[7]) ? 3'b001 : 3'b110;
										assign node73 = (inp[10]) ? node77 : node74;
											assign node74 = (inp[7]) ? 3'b001 : 3'b110;
											assign node77 = (inp[7]) ? 3'b110 : 3'b001;
									assign node80 = (inp[10]) ? node82 : 3'b110;
										assign node82 = (inp[7]) ? 3'b110 : 3'b001;
							assign node85 = (inp[7]) ? node87 : 3'b110;
								assign node87 = (inp[3]) ? node95 : node88;
									assign node88 = (inp[2]) ? node92 : node89;
										assign node89 = (inp[10]) ? 3'b110 : 3'b001;
										assign node92 = (inp[10]) ? 3'b001 : 3'b110;
									assign node95 = (inp[4]) ? node97 : 3'b110;
										assign node97 = (inp[10]) ? 3'b110 : 3'b001;
			assign node100 = (inp[0]) ? node220 : node101;
				assign node101 = (inp[9]) ? node153 : node102;
					assign node102 = (inp[6]) ? node104 : 3'b010;
						assign node104 = (inp[10]) ? node140 : node105;
							assign node105 = (inp[3]) ? node121 : node106;
								assign node106 = (inp[7]) ? node116 : node107;
									assign node107 = (inp[2]) ? node113 : node108;
										assign node108 = (inp[1]) ? 3'b001 : node109;
											assign node109 = (inp[4]) ? 3'b101 : 3'b111;
										assign node113 = (inp[1]) ? 3'b111 : 3'b011;
									assign node116 = (inp[1]) ? 3'b101 : node117;
										assign node117 = (inp[2]) ? 3'b101 : 3'b011;
								assign node121 = (inp[1]) ? node135 : node122;
									assign node122 = (inp[4]) ? node130 : node123;
										assign node123 = (inp[2]) ? node127 : node124;
											assign node124 = (inp[7]) ? 3'b011 : 3'b111;
											assign node127 = (inp[7]) ? 3'b101 : 3'b011;
										assign node130 = (inp[7]) ? node132 : 3'b101;
											assign node132 = (inp[2]) ? 3'b101 : 3'b011;
									assign node135 = (inp[7]) ? 3'b001 : node136;
										assign node136 = (inp[2]) ? 3'b011 : 3'b001;
							assign node140 = (inp[1]) ? node150 : node141;
								assign node141 = (inp[7]) ? node147 : node142;
									assign node142 = (inp[2]) ? 3'b111 : node143;
										assign node143 = (inp[4]) ? 3'b001 : 3'b011;
									assign node147 = (inp[2]) ? 3'b001 : 3'b101;
								assign node150 = (inp[7]) ? 3'b110 : 3'b010;
					assign node153 = (inp[7]) ? node193 : node154;
						assign node154 = (inp[1]) ? node180 : node155;
							assign node155 = (inp[6]) ? node163 : node156;
								assign node156 = (inp[2]) ? node160 : node157;
									assign node157 = (inp[10]) ? 3'b000 : 3'b100;
									assign node160 = (inp[10]) ? 3'b100 : 3'b000;
								assign node163 = (inp[4]) ? node175 : node164;
									assign node164 = (inp[3]) ? node170 : node165;
										assign node165 = (inp[2]) ? 3'b100 : node166;
											assign node166 = (inp[10]) ? 3'b000 : 3'b100;
										assign node170 = (inp[2]) ? 3'b000 : node171;
											assign node171 = (inp[10]) ? 3'b000 : 3'b100;
									assign node175 = (inp[10]) ? 3'b100 : node176;
										assign node176 = (inp[2]) ? 3'b010 : 3'b110;
							assign node180 = (inp[6]) ? node182 : 3'b000;
								assign node182 = (inp[10]) ? node188 : node183;
									assign node183 = (inp[2]) ? node185 : 3'b010;
										assign node185 = (inp[3]) ? 3'b000 : 3'b100;
									assign node188 = (inp[4]) ? node190 : 3'b000;
										assign node190 = (inp[2]) ? 3'b000 : 3'b100;
						assign node193 = (inp[1]) ? node207 : node194;
							assign node194 = (inp[2]) ? node202 : node195;
								assign node195 = (inp[10]) ? node199 : node196;
									assign node196 = (inp[6]) ? 3'b001 : 3'b010;
									assign node199 = (inp[3]) ? 3'b110 : 3'b100;
								assign node202 = (inp[10]) ? 3'b010 : node203;
									assign node203 = (inp[6]) ? 3'b110 : 3'b100;
							assign node207 = (inp[10]) ? node215 : node208;
								assign node208 = (inp[6]) ? node212 : node209;
									assign node209 = (inp[2]) ? 3'b000 : 3'b100;
									assign node212 = (inp[3]) ? 3'b010 : 3'b110;
								assign node215 = (inp[6]) ? 3'b100 : node216;
									assign node216 = (inp[4]) ? 3'b000 : 3'b100;
				assign node220 = (inp[6]) ? node222 : 3'b000;
					assign node222 = (inp[1]) ? node238 : node223;
						assign node223 = (inp[9]) ? node231 : node224;
							assign node224 = (inp[10]) ? node228 : node225;
								assign node225 = (inp[2]) ? 3'b010 : 3'b110;
								assign node228 = (inp[2]) ? 3'b100 : 3'b000;
							assign node231 = (inp[10]) ? 3'b000 : node232;
								assign node232 = (inp[3]) ? node234 : 3'b000;
									assign node234 = (inp[7]) ? 3'b100 : 3'b000;
						assign node238 = (inp[4]) ? node240 : 3'b000;
							assign node240 = (inp[10]) ? node248 : node241;
								assign node241 = (inp[7]) ? node243 : 3'b000;
									assign node243 = (inp[3]) ? node245 : 3'b000;
										assign node245 = (inp[9]) ? 3'b000 : 3'b010;
								assign node248 = (inp[2]) ? 3'b000 : node249;
									assign node249 = (inp[9]) ? 3'b000 : node250;
										assign node250 = (inp[3]) ? 3'b100 : 3'b000;

endmodule