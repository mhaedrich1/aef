module dtc_split5_bm99 (
	input  wire [12-1:0] inp,
	output wire [3-1:0] outp
);

	wire [3-1:0] node1;
	wire [3-1:0] node2;
	wire [3-1:0] node3;
	wire [3-1:0] node4;
	wire [3-1:0] node5;
	wire [3-1:0] node6;
	wire [3-1:0] node11;
	wire [3-1:0] node12;
	wire [3-1:0] node13;
	wire [3-1:0] node14;
	wire [3-1:0] node16;
	wire [3-1:0] node17;
	wire [3-1:0] node20;
	wire [3-1:0] node21;
	wire [3-1:0] node26;
	wire [3-1:0] node27;
	wire [3-1:0] node28;
	wire [3-1:0] node29;
	wire [3-1:0] node30;
	wire [3-1:0] node34;
	wire [3-1:0] node37;
	wire [3-1:0] node38;
	wire [3-1:0] node39;
	wire [3-1:0] node46;
	wire [3-1:0] node48;
	wire [3-1:0] node49;
	wire [3-1:0] node50;
	wire [3-1:0] node51;
	wire [3-1:0] node53;
	wire [3-1:0] node55;
	wire [3-1:0] node59;
	wire [3-1:0] node60;
	wire [3-1:0] node62;
	wire [3-1:0] node66;
	wire [3-1:0] node67;
	wire [3-1:0] node71;
	wire [3-1:0] node72;
	wire [3-1:0] node73;
	wire [3-1:0] node74;
	wire [3-1:0] node75;
	wire [3-1:0] node76;
	wire [3-1:0] node80;
	wire [3-1:0] node83;
	wire [3-1:0] node84;
	wire [3-1:0] node85;
	wire [3-1:0] node86;
	wire [3-1:0] node87;
	wire [3-1:0] node89;
	wire [3-1:0] node92;
	wire [3-1:0] node93;
	wire [3-1:0] node98;
	wire [3-1:0] node99;
	wire [3-1:0] node100;
	wire [3-1:0] node102;
	wire [3-1:0] node107;
	wire [3-1:0] node108;
	wire [3-1:0] node109;
	wire [3-1:0] node110;
	wire [3-1:0] node112;
	wire [3-1:0] node116;
	wire [3-1:0] node117;
	wire [3-1:0] node119;
	wire [3-1:0] node122;
	wire [3-1:0] node126;
	wire [3-1:0] node127;
	wire [3-1:0] node128;
	wire [3-1:0] node130;
	wire [3-1:0] node132;
	wire [3-1:0] node133;
	wire [3-1:0] node138;
	wire [3-1:0] node139;
	wire [3-1:0] node140;
	wire [3-1:0] node142;
	wire [3-1:0] node144;
	wire [3-1:0] node148;
	wire [3-1:0] node149;
	wire [3-1:0] node151;
	wire [3-1:0] node155;
	wire [3-1:0] node156;
	wire [3-1:0] node158;
	wire [3-1:0] node160;
	wire [3-1:0] node161;
	wire [3-1:0] node162;
	wire [3-1:0] node164;
	wire [3-1:0] node169;
	wire [3-1:0] node170;
	wire [3-1:0] node171;
	wire [3-1:0] node173;
	wire [3-1:0] node175;
	wire [3-1:0] node178;
	wire [3-1:0] node181;
	wire [3-1:0] node182;
	wire [3-1:0] node183;
	wire [3-1:0] node185;
	wire [3-1:0] node187;
	wire [3-1:0] node191;
	wire [3-1:0] node192;
	wire [3-1:0] node194;
	wire [3-1:0] node198;
	wire [3-1:0] node200;
	wire [3-1:0] node201;
	wire [3-1:0] node202;
	wire [3-1:0] node205;
	wire [3-1:0] node206;
	wire [3-1:0] node208;
	wire [3-1:0] node210;
	wire [3-1:0] node211;
	wire [3-1:0] node216;
	wire [3-1:0] node217;
	wire [3-1:0] node220;
	wire [3-1:0] node221;
	wire [3-1:0] node222;
	wire [3-1:0] node223;
	wire [3-1:0] node225;
	wire [3-1:0] node227;
	wire [3-1:0] node231;
	wire [3-1:0] node233;
	wire [3-1:0] node234;
	wire [3-1:0] node236;
	wire [3-1:0] node239;
	wire [3-1:0] node241;
	wire [3-1:0] node244;
	wire [3-1:0] node246;
	wire [3-1:0] node247;
	wire [3-1:0] node249;
	wire [3-1:0] node251;
	wire [3-1:0] node252;

	assign outp = (inp[3]) ? node198 : node1;
		assign node1 = (inp[9]) ? node71 : node2;
			assign node2 = (inp[4]) ? node46 : node3;
				assign node3 = (inp[0]) ? node11 : node4;
					assign node4 = (inp[6]) ? 3'b000 : node5;
						assign node5 = (inp[1]) ? 3'b001 : node6;
							assign node6 = (inp[5]) ? 3'b000 : 3'b001;
					assign node11 = (inp[6]) ? 3'b001 : node12;
						assign node12 = (inp[5]) ? node26 : node13;
							assign node13 = (inp[1]) ? 3'b000 : node14;
								assign node14 = (inp[7]) ? node16 : 3'b000;
									assign node16 = (inp[10]) ? node20 : node17;
										assign node17 = (inp[11]) ? 3'b000 : 3'b001;
										assign node20 = (inp[8]) ? 3'b000 : node21;
											assign node21 = (inp[11]) ? 3'b001 : 3'b000;
							assign node26 = (inp[1]) ? 3'b001 : node27;
								assign node27 = (inp[7]) ? node37 : node28;
									assign node28 = (inp[2]) ? node34 : node29;
										assign node29 = (inp[8]) ? 3'b000 : node30;
											assign node30 = (inp[11]) ? 3'b001 : 3'b000;
										assign node34 = (inp[11]) ? 3'b000 : 3'b001;
									assign node37 = (inp[8]) ? 3'b000 : node38;
										assign node38 = (inp[2]) ? 3'b000 : node39;
											assign node39 = (inp[11]) ? 3'b001 : 3'b000;
				assign node46 = (inp[0]) ? node48 : 3'b000;
					assign node48 = (inp[6]) ? node66 : node49;
						assign node49 = (inp[5]) ? node59 : node50;
							assign node50 = (inp[1]) ? 3'b001 : node51;
								assign node51 = (inp[7]) ? node53 : 3'b000;
									assign node53 = (inp[2]) ? node55 : 3'b000;
										assign node55 = (inp[10]) ? 3'b001 : 3'b000;
							assign node59 = (inp[1]) ? 3'b000 : node60;
								assign node60 = (inp[7]) ? node62 : 3'b000;
									assign node62 = (inp[10]) ? 3'b001 : 3'b000;
						assign node66 = (inp[1]) ? 3'b000 : node67;
							assign node67 = (inp[5]) ? 3'b001 : 3'b000;
			assign node71 = (inp[6]) ? node155 : node72;
				assign node72 = (inp[4]) ? node126 : node73;
					assign node73 = (inp[0]) ? node83 : node74;
						assign node74 = (inp[5]) ? node80 : node75;
							assign node75 = (inp[1]) ? 3'b110 : node76;
								assign node76 = (inp[7]) ? 3'b110 : 3'b010;
							assign node80 = (inp[1]) ? 3'b010 : 3'b100;
						assign node83 = (inp[5]) ? node107 : node84;
							assign node84 = (inp[7]) ? node98 : node85;
								assign node85 = (inp[1]) ? 3'b001 : node86;
									assign node86 = (inp[11]) ? node92 : node87;
										assign node87 = (inp[2]) ? node89 : 3'b001;
											assign node89 = (inp[8]) ? 3'b110 : 3'b001;
										assign node92 = (inp[2]) ? 3'b001 : node93;
											assign node93 = (inp[10]) ? 3'b110 : 3'b001;
								assign node98 = (inp[1]) ? 3'b101 : node99;
									assign node99 = (inp[2]) ? 3'b110 : node100;
										assign node100 = (inp[11]) ? node102 : 3'b001;
											assign node102 = (inp[8]) ? 3'b001 : 3'b110;
							assign node107 = (inp[1]) ? 3'b110 : node108;
								assign node108 = (inp[7]) ? node116 : node109;
									assign node109 = (inp[11]) ? 3'b001 : node110;
										assign node110 = (inp[2]) ? node112 : 3'b001;
											assign node112 = (inp[8]) ? 3'b110 : 3'b001;
									assign node116 = (inp[11]) ? node122 : node117;
										assign node117 = (inp[2]) ? node119 : 3'b001;
											assign node119 = (inp[8]) ? 3'b110 : 3'b001;
										assign node122 = (inp[2]) ? 3'b001 : 3'b110;
					assign node126 = (inp[0]) ? node138 : node127;
						assign node127 = (inp[7]) ? 3'b000 : node128;
							assign node128 = (inp[2]) ? node130 : 3'b000;
								assign node130 = (inp[11]) ? node132 : 3'b000;
									assign node132 = (inp[5]) ? 3'b000 : node133;
										assign node133 = (inp[10]) ? 3'b100 : 3'b000;
						assign node138 = (inp[5]) ? node148 : node139;
							assign node139 = (inp[1]) ? 3'b010 : node140;
								assign node140 = (inp[2]) ? node142 : 3'b100;
									assign node142 = (inp[10]) ? node144 : 3'b100;
										assign node144 = (inp[7]) ? 3'b010 : 3'b100;
							assign node148 = (inp[1]) ? 3'b100 : node149;
								assign node149 = (inp[7]) ? node151 : 3'b100;
									assign node151 = (inp[10]) ? 3'b010 : 3'b100;
				assign node155 = (inp[0]) ? node169 : node156;
					assign node156 = (inp[8]) ? node158 : 3'b001;
						assign node158 = (inp[2]) ? node160 : 3'b001;
							assign node160 = (inp[5]) ? 3'b001 : node161;
								assign node161 = (inp[4]) ? 3'b001 : node162;
									assign node162 = (inp[10]) ? node164 : 3'b001;
										assign node164 = (inp[7]) ? 3'b011 : 3'b001;
					assign node169 = (inp[4]) ? node181 : node170;
						assign node170 = (inp[1]) ? node178 : node171;
							assign node171 = (inp[10]) ? node173 : 3'b011;
								assign node173 = (inp[7]) ? node175 : 3'b011;
									assign node175 = (inp[5]) ? 3'b111 : 3'b011;
							assign node178 = (inp[5]) ? 3'b011 : 3'b111;
						assign node181 = (inp[5]) ? node191 : node182;
							assign node182 = (inp[1]) ? 3'b101 : node183;
								assign node183 = (inp[7]) ? node185 : 3'b001;
									assign node185 = (inp[10]) ? node187 : 3'b001;
										assign node187 = (inp[2]) ? 3'b101 : 3'b001;
							assign node191 = (inp[1]) ? 3'b001 : node192;
								assign node192 = (inp[7]) ? node194 : 3'b010;
									assign node194 = (inp[10]) ? 3'b110 : 3'b010;
		assign node198 = (inp[6]) ? node200 : 3'b000;
			assign node200 = (inp[0]) ? node216 : node201;
				assign node201 = (inp[4]) ? node205 : node202;
					assign node202 = (inp[9]) ? 3'b100 : 3'b000;
					assign node205 = (inp[9]) ? 3'b000 : node206;
						assign node206 = (inp[10]) ? node208 : 3'b010;
							assign node208 = (inp[1]) ? node210 : 3'b010;
								assign node210 = (inp[5]) ? 3'b100 : node211;
									assign node211 = (inp[2]) ? 3'b100 : 3'b010;
				assign node216 = (inp[4]) ? node220 : node217;
					assign node217 = (inp[9]) ? 3'b010 : 3'b001;
					assign node220 = (inp[9]) ? node244 : node221;
						assign node221 = (inp[1]) ? node231 : node222;
							assign node222 = (inp[10]) ? 3'b010 : node223;
								assign node223 = (inp[7]) ? node225 : 3'b010;
									assign node225 = (inp[11]) ? node227 : 3'b110;
										assign node227 = (inp[2]) ? 3'b110 : 3'b010;
							assign node231 = (inp[7]) ? node233 : 3'b110;
								assign node233 = (inp[10]) ? node239 : node234;
									assign node234 = (inp[2]) ? node236 : 3'b110;
										assign node236 = (inp[11]) ? 3'b110 : 3'b001;
									assign node239 = (inp[2]) ? node241 : 3'b010;
										assign node241 = (inp[8]) ? 3'b110 : 3'b010;
						assign node244 = (inp[7]) ? node246 : 3'b000;
							assign node246 = (inp[10]) ? 3'b000 : node247;
								assign node247 = (inp[11]) ? node249 : 3'b100;
									assign node249 = (inp[1]) ? node251 : 3'b000;
										assign node251 = (inp[8]) ? 3'b100 : node252;
											assign node252 = (inp[2]) ? 3'b100 : 3'b000;

endmodule