module dtc_split75_bm62 (
	input  wire [16-1:0] inp,
	output wire [4-1:0] outp
);

	wire [4-1:0] node1;
	wire [4-1:0] node2;
	wire [4-1:0] node3;
	wire [4-1:0] node4;
	wire [4-1:0] node5;
	wire [4-1:0] node6;
	wire [4-1:0] node7;
	wire [4-1:0] node8;
	wire [4-1:0] node9;
	wire [4-1:0] node10;
	wire [4-1:0] node11;
	wire [4-1:0] node12;
	wire [4-1:0] node13;
	wire [4-1:0] node15;
	wire [4-1:0] node18;
	wire [4-1:0] node19;
	wire [4-1:0] node21;
	wire [4-1:0] node24;
	wire [4-1:0] node25;
	wire [4-1:0] node28;
	wire [4-1:0] node31;
	wire [4-1:0] node32;
	wire [4-1:0] node34;
	wire [4-1:0] node36;
	wire [4-1:0] node39;
	wire [4-1:0] node40;
	wire [4-1:0] node41;
	wire [4-1:0] node44;
	wire [4-1:0] node47;
	wire [4-1:0] node48;
	wire [4-1:0] node52;
	wire [4-1:0] node53;
	wire [4-1:0] node54;
	wire [4-1:0] node55;
	wire [4-1:0] node56;
	wire [4-1:0] node59;
	wire [4-1:0] node63;
	wire [4-1:0] node64;
	wire [4-1:0] node66;
	wire [4-1:0] node69;
	wire [4-1:0] node71;
	wire [4-1:0] node74;
	wire [4-1:0] node75;
	wire [4-1:0] node76;
	wire [4-1:0] node79;
	wire [4-1:0] node80;
	wire [4-1:0] node83;
	wire [4-1:0] node86;
	wire [4-1:0] node87;
	wire [4-1:0] node88;
	wire [4-1:0] node91;
	wire [4-1:0] node94;
	wire [4-1:0] node95;
	wire [4-1:0] node99;
	wire [4-1:0] node100;
	wire [4-1:0] node101;
	wire [4-1:0] node102;
	wire [4-1:0] node105;
	wire [4-1:0] node108;
	wire [4-1:0] node109;
	wire [4-1:0] node112;
	wire [4-1:0] node115;
	wire [4-1:0] node116;
	wire [4-1:0] node117;
	wire [4-1:0] node120;
	wire [4-1:0] node123;
	wire [4-1:0] node124;
	wire [4-1:0] node125;
	wire [4-1:0] node128;
	wire [4-1:0] node131;
	wire [4-1:0] node132;
	wire [4-1:0] node135;
	wire [4-1:0] node138;
	wire [4-1:0] node139;
	wire [4-1:0] node140;
	wire [4-1:0] node141;
	wire [4-1:0] node142;
	wire [4-1:0] node143;
	wire [4-1:0] node144;
	wire [4-1:0] node148;
	wire [4-1:0] node150;
	wire [4-1:0] node153;
	wire [4-1:0] node154;
	wire [4-1:0] node155;
	wire [4-1:0] node158;
	wire [4-1:0] node161;
	wire [4-1:0] node163;
	wire [4-1:0] node166;
	wire [4-1:0] node167;
	wire [4-1:0] node168;
	wire [4-1:0] node170;
	wire [4-1:0] node173;
	wire [4-1:0] node174;
	wire [4-1:0] node178;
	wire [4-1:0] node179;
	wire [4-1:0] node180;
	wire [4-1:0] node183;
	wire [4-1:0] node186;
	wire [4-1:0] node187;
	wire [4-1:0] node190;
	wire [4-1:0] node193;
	wire [4-1:0] node194;
	wire [4-1:0] node195;
	wire [4-1:0] node196;
	wire [4-1:0] node197;
	wire [4-1:0] node201;
	wire [4-1:0] node203;
	wire [4-1:0] node206;
	wire [4-1:0] node208;
	wire [4-1:0] node209;
	wire [4-1:0] node213;
	wire [4-1:0] node214;
	wire [4-1:0] node215;
	wire [4-1:0] node216;
	wire [4-1:0] node219;
	wire [4-1:0] node222;
	wire [4-1:0] node223;
	wire [4-1:0] node226;
	wire [4-1:0] node229;
	wire [4-1:0] node230;
	wire [4-1:0] node231;
	wire [4-1:0] node236;
	wire [4-1:0] node237;
	wire [4-1:0] node238;
	wire [4-1:0] node239;
	wire [4-1:0] node240;
	wire [4-1:0] node243;
	wire [4-1:0] node246;
	wire [4-1:0] node247;
	wire [4-1:0] node248;
	wire [4-1:0] node251;
	wire [4-1:0] node255;
	wire [4-1:0] node256;
	wire [4-1:0] node257;
	wire [4-1:0] node260;
	wire [4-1:0] node263;
	wire [4-1:0] node264;
	wire [4-1:0] node265;
	wire [4-1:0] node268;
	wire [4-1:0] node271;
	wire [4-1:0] node273;
	wire [4-1:0] node276;
	wire [4-1:0] node277;
	wire [4-1:0] node278;
	wire [4-1:0] node279;
	wire [4-1:0] node282;
	wire [4-1:0] node286;
	wire [4-1:0] node287;
	wire [4-1:0] node288;
	wire [4-1:0] node292;
	wire [4-1:0] node294;
	wire [4-1:0] node295;
	wire [4-1:0] node299;
	wire [4-1:0] node300;
	wire [4-1:0] node301;
	wire [4-1:0] node302;
	wire [4-1:0] node303;
	wire [4-1:0] node304;
	wire [4-1:0] node305;
	wire [4-1:0] node308;
	wire [4-1:0] node311;
	wire [4-1:0] node312;
	wire [4-1:0] node315;
	wire [4-1:0] node318;
	wire [4-1:0] node319;
	wire [4-1:0] node320;
	wire [4-1:0] node323;
	wire [4-1:0] node326;
	wire [4-1:0] node327;
	wire [4-1:0] node330;
	wire [4-1:0] node333;
	wire [4-1:0] node334;
	wire [4-1:0] node335;
	wire [4-1:0] node336;
	wire [4-1:0] node339;
	wire [4-1:0] node342;
	wire [4-1:0] node344;
	wire [4-1:0] node347;
	wire [4-1:0] node348;
	wire [4-1:0] node349;
	wire [4-1:0] node352;
	wire [4-1:0] node355;
	wire [4-1:0] node356;
	wire [4-1:0] node359;
	wire [4-1:0] node362;
	wire [4-1:0] node363;
	wire [4-1:0] node364;
	wire [4-1:0] node365;
	wire [4-1:0] node366;
	wire [4-1:0] node367;
	wire [4-1:0] node371;
	wire [4-1:0] node372;
	wire [4-1:0] node376;
	wire [4-1:0] node377;
	wire [4-1:0] node379;
	wire [4-1:0] node382;
	wire [4-1:0] node383;
	wire [4-1:0] node386;
	wire [4-1:0] node389;
	wire [4-1:0] node390;
	wire [4-1:0] node391;
	wire [4-1:0] node392;
	wire [4-1:0] node396;
	wire [4-1:0] node397;
	wire [4-1:0] node401;
	wire [4-1:0] node402;
	wire [4-1:0] node403;
	wire [4-1:0] node406;
	wire [4-1:0] node409;
	wire [4-1:0] node412;
	wire [4-1:0] node413;
	wire [4-1:0] node414;
	wire [4-1:0] node416;
	wire [4-1:0] node417;
	wire [4-1:0] node421;
	wire [4-1:0] node422;
	wire [4-1:0] node425;
	wire [4-1:0] node426;
	wire [4-1:0] node429;
	wire [4-1:0] node432;
	wire [4-1:0] node433;
	wire [4-1:0] node434;
	wire [4-1:0] node435;
	wire [4-1:0] node439;
	wire [4-1:0] node441;
	wire [4-1:0] node444;
	wire [4-1:0] node446;
	wire [4-1:0] node447;
	wire [4-1:0] node450;
	wire [4-1:0] node453;
	wire [4-1:0] node454;
	wire [4-1:0] node455;
	wire [4-1:0] node456;
	wire [4-1:0] node457;
	wire [4-1:0] node458;
	wire [4-1:0] node462;
	wire [4-1:0] node463;
	wire [4-1:0] node466;
	wire [4-1:0] node469;
	wire [4-1:0] node470;
	wire [4-1:0] node473;
	wire [4-1:0] node474;
	wire [4-1:0] node478;
	wire [4-1:0] node479;
	wire [4-1:0] node480;
	wire [4-1:0] node481;
	wire [4-1:0] node484;
	wire [4-1:0] node487;
	wire [4-1:0] node488;
	wire [4-1:0] node491;
	wire [4-1:0] node494;
	wire [4-1:0] node495;
	wire [4-1:0] node497;
	wire [4-1:0] node500;
	wire [4-1:0] node501;
	wire [4-1:0] node504;
	wire [4-1:0] node507;
	wire [4-1:0] node508;
	wire [4-1:0] node509;
	wire [4-1:0] node510;
	wire [4-1:0] node511;
	wire [4-1:0] node514;
	wire [4-1:0] node517;
	wire [4-1:0] node518;
	wire [4-1:0] node520;
	wire [4-1:0] node523;
	wire [4-1:0] node524;
	wire [4-1:0] node527;
	wire [4-1:0] node530;
	wire [4-1:0] node531;
	wire [4-1:0] node532;
	wire [4-1:0] node536;
	wire [4-1:0] node537;
	wire [4-1:0] node538;
	wire [4-1:0] node541;
	wire [4-1:0] node544;
	wire [4-1:0] node545;
	wire [4-1:0] node548;
	wire [4-1:0] node551;
	wire [4-1:0] node552;
	wire [4-1:0] node553;
	wire [4-1:0] node554;
	wire [4-1:0] node555;
	wire [4-1:0] node559;
	wire [4-1:0] node561;
	wire [4-1:0] node564;
	wire [4-1:0] node565;
	wire [4-1:0] node566;
	wire [4-1:0] node569;
	wire [4-1:0] node572;
	wire [4-1:0] node573;
	wire [4-1:0] node576;
	wire [4-1:0] node579;
	wire [4-1:0] node580;
	wire [4-1:0] node581;
	wire [4-1:0] node582;
	wire [4-1:0] node585;
	wire [4-1:0] node588;
	wire [4-1:0] node589;
	wire [4-1:0] node592;
	wire [4-1:0] node595;
	wire [4-1:0] node596;
	wire [4-1:0] node597;
	wire [4-1:0] node601;
	wire [4-1:0] node602;
	wire [4-1:0] node605;
	wire [4-1:0] node608;
	wire [4-1:0] node609;
	wire [4-1:0] node610;
	wire [4-1:0] node611;
	wire [4-1:0] node612;
	wire [4-1:0] node613;
	wire [4-1:0] node614;
	wire [4-1:0] node615;
	wire [4-1:0] node617;
	wire [4-1:0] node620;
	wire [4-1:0] node621;
	wire [4-1:0] node624;
	wire [4-1:0] node627;
	wire [4-1:0] node628;
	wire [4-1:0] node629;
	wire [4-1:0] node633;
	wire [4-1:0] node635;
	wire [4-1:0] node638;
	wire [4-1:0] node639;
	wire [4-1:0] node640;
	wire [4-1:0] node641;
	wire [4-1:0] node644;
	wire [4-1:0] node647;
	wire [4-1:0] node648;
	wire [4-1:0] node651;
	wire [4-1:0] node654;
	wire [4-1:0] node656;
	wire [4-1:0] node657;
	wire [4-1:0] node660;
	wire [4-1:0] node663;
	wire [4-1:0] node664;
	wire [4-1:0] node665;
	wire [4-1:0] node666;
	wire [4-1:0] node667;
	wire [4-1:0] node670;
	wire [4-1:0] node673;
	wire [4-1:0] node674;
	wire [4-1:0] node677;
	wire [4-1:0] node680;
	wire [4-1:0] node681;
	wire [4-1:0] node682;
	wire [4-1:0] node686;
	wire [4-1:0] node687;
	wire [4-1:0] node691;
	wire [4-1:0] node692;
	wire [4-1:0] node694;
	wire [4-1:0] node695;
	wire [4-1:0] node698;
	wire [4-1:0] node701;
	wire [4-1:0] node702;
	wire [4-1:0] node703;
	wire [4-1:0] node706;
	wire [4-1:0] node710;
	wire [4-1:0] node711;
	wire [4-1:0] node712;
	wire [4-1:0] node713;
	wire [4-1:0] node714;
	wire [4-1:0] node715;
	wire [4-1:0] node719;
	wire [4-1:0] node720;
	wire [4-1:0] node723;
	wire [4-1:0] node726;
	wire [4-1:0] node728;
	wire [4-1:0] node729;
	wire [4-1:0] node732;
	wire [4-1:0] node735;
	wire [4-1:0] node736;
	wire [4-1:0] node737;
	wire [4-1:0] node738;
	wire [4-1:0] node741;
	wire [4-1:0] node744;
	wire [4-1:0] node745;
	wire [4-1:0] node748;
	wire [4-1:0] node751;
	wire [4-1:0] node753;
	wire [4-1:0] node754;
	wire [4-1:0] node757;
	wire [4-1:0] node760;
	wire [4-1:0] node761;
	wire [4-1:0] node762;
	wire [4-1:0] node763;
	wire [4-1:0] node764;
	wire [4-1:0] node767;
	wire [4-1:0] node771;
	wire [4-1:0] node772;
	wire [4-1:0] node773;
	wire [4-1:0] node776;
	wire [4-1:0] node779;
	wire [4-1:0] node781;
	wire [4-1:0] node784;
	wire [4-1:0] node785;
	wire [4-1:0] node786;
	wire [4-1:0] node787;
	wire [4-1:0] node791;
	wire [4-1:0] node793;
	wire [4-1:0] node796;
	wire [4-1:0] node799;
	wire [4-1:0] node800;
	wire [4-1:0] node801;
	wire [4-1:0] node802;
	wire [4-1:0] node803;
	wire [4-1:0] node804;
	wire [4-1:0] node807;
	wire [4-1:0] node810;
	wire [4-1:0] node811;
	wire [4-1:0] node814;
	wire [4-1:0] node815;
	wire [4-1:0] node819;
	wire [4-1:0] node820;
	wire [4-1:0] node823;
	wire [4-1:0] node824;
	wire [4-1:0] node826;
	wire [4-1:0] node829;
	wire [4-1:0] node830;
	wire [4-1:0] node834;
	wire [4-1:0] node835;
	wire [4-1:0] node836;
	wire [4-1:0] node837;
	wire [4-1:0] node838;
	wire [4-1:0] node841;
	wire [4-1:0] node844;
	wire [4-1:0] node845;
	wire [4-1:0] node849;
	wire [4-1:0] node850;
	wire [4-1:0] node851;
	wire [4-1:0] node854;
	wire [4-1:0] node858;
	wire [4-1:0] node859;
	wire [4-1:0] node861;
	wire [4-1:0] node863;
	wire [4-1:0] node866;
	wire [4-1:0] node867;
	wire [4-1:0] node870;
	wire [4-1:0] node873;
	wire [4-1:0] node874;
	wire [4-1:0] node875;
	wire [4-1:0] node876;
	wire [4-1:0] node877;
	wire [4-1:0] node878;
	wire [4-1:0] node881;
	wire [4-1:0] node884;
	wire [4-1:0] node886;
	wire [4-1:0] node889;
	wire [4-1:0] node891;
	wire [4-1:0] node894;
	wire [4-1:0] node895;
	wire [4-1:0] node896;
	wire [4-1:0] node897;
	wire [4-1:0] node901;
	wire [4-1:0] node902;
	wire [4-1:0] node905;
	wire [4-1:0] node908;
	wire [4-1:0] node910;
	wire [4-1:0] node912;
	wire [4-1:0] node915;
	wire [4-1:0] node916;
	wire [4-1:0] node917;
	wire [4-1:0] node918;
	wire [4-1:0] node919;
	wire [4-1:0] node922;
	wire [4-1:0] node925;
	wire [4-1:0] node926;
	wire [4-1:0] node929;
	wire [4-1:0] node932;
	wire [4-1:0] node933;
	wire [4-1:0] node934;
	wire [4-1:0] node938;
	wire [4-1:0] node939;
	wire [4-1:0] node942;
	wire [4-1:0] node945;
	wire [4-1:0] node946;
	wire [4-1:0] node948;
	wire [4-1:0] node949;
	wire [4-1:0] node953;
	wire [4-1:0] node954;
	wire [4-1:0] node956;
	wire [4-1:0] node959;
	wire [4-1:0] node961;
	wire [4-1:0] node964;
	wire [4-1:0] node965;
	wire [4-1:0] node966;
	wire [4-1:0] node967;
	wire [4-1:0] node968;
	wire [4-1:0] node969;
	wire [4-1:0] node970;
	wire [4-1:0] node971;
	wire [4-1:0] node974;
	wire [4-1:0] node977;
	wire [4-1:0] node979;
	wire [4-1:0] node982;
	wire [4-1:0] node983;
	wire [4-1:0] node985;
	wire [4-1:0] node988;
	wire [4-1:0] node991;
	wire [4-1:0] node992;
	wire [4-1:0] node993;
	wire [4-1:0] node996;
	wire [4-1:0] node998;
	wire [4-1:0] node1001;
	wire [4-1:0] node1002;
	wire [4-1:0] node1003;
	wire [4-1:0] node1007;
	wire [4-1:0] node1008;
	wire [4-1:0] node1012;
	wire [4-1:0] node1013;
	wire [4-1:0] node1014;
	wire [4-1:0] node1016;
	wire [4-1:0] node1019;
	wire [4-1:0] node1020;
	wire [4-1:0] node1022;
	wire [4-1:0] node1025;
	wire [4-1:0] node1026;
	wire [4-1:0] node1030;
	wire [4-1:0] node1031;
	wire [4-1:0] node1032;
	wire [4-1:0] node1035;
	wire [4-1:0] node1038;
	wire [4-1:0] node1039;
	wire [4-1:0] node1040;
	wire [4-1:0] node1045;
	wire [4-1:0] node1046;
	wire [4-1:0] node1047;
	wire [4-1:0] node1049;
	wire [4-1:0] node1050;
	wire [4-1:0] node1052;
	wire [4-1:0] node1055;
	wire [4-1:0] node1057;
	wire [4-1:0] node1060;
	wire [4-1:0] node1061;
	wire [4-1:0] node1063;
	wire [4-1:0] node1064;
	wire [4-1:0] node1068;
	wire [4-1:0] node1069;
	wire [4-1:0] node1073;
	wire [4-1:0] node1074;
	wire [4-1:0] node1075;
	wire [4-1:0] node1077;
	wire [4-1:0] node1080;
	wire [4-1:0] node1081;
	wire [4-1:0] node1082;
	wire [4-1:0] node1086;
	wire [4-1:0] node1089;
	wire [4-1:0] node1090;
	wire [4-1:0] node1091;
	wire [4-1:0] node1092;
	wire [4-1:0] node1096;
	wire [4-1:0] node1097;
	wire [4-1:0] node1101;
	wire [4-1:0] node1103;
	wire [4-1:0] node1106;
	wire [4-1:0] node1107;
	wire [4-1:0] node1108;
	wire [4-1:0] node1109;
	wire [4-1:0] node1110;
	wire [4-1:0] node1112;
	wire [4-1:0] node1115;
	wire [4-1:0] node1116;
	wire [4-1:0] node1118;
	wire [4-1:0] node1121;
	wire [4-1:0] node1122;
	wire [4-1:0] node1125;
	wire [4-1:0] node1128;
	wire [4-1:0] node1129;
	wire [4-1:0] node1130;
	wire [4-1:0] node1132;
	wire [4-1:0] node1135;
	wire [4-1:0] node1136;
	wire [4-1:0] node1140;
	wire [4-1:0] node1141;
	wire [4-1:0] node1143;
	wire [4-1:0] node1146;
	wire [4-1:0] node1149;
	wire [4-1:0] node1150;
	wire [4-1:0] node1151;
	wire [4-1:0] node1152;
	wire [4-1:0] node1153;
	wire [4-1:0] node1156;
	wire [4-1:0] node1159;
	wire [4-1:0] node1161;
	wire [4-1:0] node1164;
	wire [4-1:0] node1165;
	wire [4-1:0] node1168;
	wire [4-1:0] node1171;
	wire [4-1:0] node1172;
	wire [4-1:0] node1173;
	wire [4-1:0] node1174;
	wire [4-1:0] node1177;
	wire [4-1:0] node1180;
	wire [4-1:0] node1181;
	wire [4-1:0] node1184;
	wire [4-1:0] node1187;
	wire [4-1:0] node1188;
	wire [4-1:0] node1191;
	wire [4-1:0] node1194;
	wire [4-1:0] node1195;
	wire [4-1:0] node1196;
	wire [4-1:0] node1197;
	wire [4-1:0] node1198;
	wire [4-1:0] node1199;
	wire [4-1:0] node1202;
	wire [4-1:0] node1205;
	wire [4-1:0] node1206;
	wire [4-1:0] node1210;
	wire [4-1:0] node1211;
	wire [4-1:0] node1212;
	wire [4-1:0] node1215;
	wire [4-1:0] node1219;
	wire [4-1:0] node1220;
	wire [4-1:0] node1221;
	wire [4-1:0] node1223;
	wire [4-1:0] node1226;
	wire [4-1:0] node1227;
	wire [4-1:0] node1231;
	wire [4-1:0] node1233;
	wire [4-1:0] node1234;
	wire [4-1:0] node1238;
	wire [4-1:0] node1239;
	wire [4-1:0] node1240;
	wire [4-1:0] node1241;
	wire [4-1:0] node1242;
	wire [4-1:0] node1245;
	wire [4-1:0] node1248;
	wire [4-1:0] node1250;
	wire [4-1:0] node1253;
	wire [4-1:0] node1254;
	wire [4-1:0] node1255;
	wire [4-1:0] node1258;
	wire [4-1:0] node1262;
	wire [4-1:0] node1263;
	wire [4-1:0] node1265;
	wire [4-1:0] node1267;
	wire [4-1:0] node1270;
	wire [4-1:0] node1271;
	wire [4-1:0] node1272;
	wire [4-1:0] node1276;
	wire [4-1:0] node1279;
	wire [4-1:0] node1280;
	wire [4-1:0] node1281;
	wire [4-1:0] node1282;
	wire [4-1:0] node1283;
	wire [4-1:0] node1284;
	wire [4-1:0] node1285;
	wire [4-1:0] node1286;
	wire [4-1:0] node1288;
	wire [4-1:0] node1291;
	wire [4-1:0] node1293;
	wire [4-1:0] node1296;
	wire [4-1:0] node1297;
	wire [4-1:0] node1298;
	wire [4-1:0] node1301;
	wire [4-1:0] node1304;
	wire [4-1:0] node1305;
	wire [4-1:0] node1308;
	wire [4-1:0] node1311;
	wire [4-1:0] node1312;
	wire [4-1:0] node1313;
	wire [4-1:0] node1316;
	wire [4-1:0] node1319;
	wire [4-1:0] node1320;
	wire [4-1:0] node1321;
	wire [4-1:0] node1324;
	wire [4-1:0] node1326;
	wire [4-1:0] node1329;
	wire [4-1:0] node1330;
	wire [4-1:0] node1332;
	wire [4-1:0] node1336;
	wire [4-1:0] node1337;
	wire [4-1:0] node1338;
	wire [4-1:0] node1339;
	wire [4-1:0] node1341;
	wire [4-1:0] node1344;
	wire [4-1:0] node1346;
	wire [4-1:0] node1349;
	wire [4-1:0] node1350;
	wire [4-1:0] node1353;
	wire [4-1:0] node1355;
	wire [4-1:0] node1358;
	wire [4-1:0] node1359;
	wire [4-1:0] node1360;
	wire [4-1:0] node1362;
	wire [4-1:0] node1365;
	wire [4-1:0] node1367;
	wire [4-1:0] node1368;
	wire [4-1:0] node1371;
	wire [4-1:0] node1374;
	wire [4-1:0] node1375;
	wire [4-1:0] node1376;
	wire [4-1:0] node1377;
	wire [4-1:0] node1380;
	wire [4-1:0] node1383;
	wire [4-1:0] node1385;
	wire [4-1:0] node1388;
	wire [4-1:0] node1389;
	wire [4-1:0] node1390;
	wire [4-1:0] node1393;
	wire [4-1:0] node1396;
	wire [4-1:0] node1397;
	wire [4-1:0] node1400;
	wire [4-1:0] node1403;
	wire [4-1:0] node1404;
	wire [4-1:0] node1405;
	wire [4-1:0] node1406;
	wire [4-1:0] node1407;
	wire [4-1:0] node1408;
	wire [4-1:0] node1409;
	wire [4-1:0] node1412;
	wire [4-1:0] node1416;
	wire [4-1:0] node1418;
	wire [4-1:0] node1419;
	wire [4-1:0] node1422;
	wire [4-1:0] node1425;
	wire [4-1:0] node1426;
	wire [4-1:0] node1428;
	wire [4-1:0] node1429;
	wire [4-1:0] node1432;
	wire [4-1:0] node1435;
	wire [4-1:0] node1437;
	wire [4-1:0] node1440;
	wire [4-1:0] node1441;
	wire [4-1:0] node1442;
	wire [4-1:0] node1444;
	wire [4-1:0] node1447;
	wire [4-1:0] node1449;
	wire [4-1:0] node1450;
	wire [4-1:0] node1453;
	wire [4-1:0] node1456;
	wire [4-1:0] node1457;
	wire [4-1:0] node1458;
	wire [4-1:0] node1459;
	wire [4-1:0] node1463;
	wire [4-1:0] node1464;
	wire [4-1:0] node1468;
	wire [4-1:0] node1471;
	wire [4-1:0] node1472;
	wire [4-1:0] node1473;
	wire [4-1:0] node1474;
	wire [4-1:0] node1475;
	wire [4-1:0] node1479;
	wire [4-1:0] node1480;
	wire [4-1:0] node1483;
	wire [4-1:0] node1486;
	wire [4-1:0] node1487;
	wire [4-1:0] node1488;
	wire [4-1:0] node1491;
	wire [4-1:0] node1494;
	wire [4-1:0] node1495;
	wire [4-1:0] node1496;
	wire [4-1:0] node1499;
	wire [4-1:0] node1502;
	wire [4-1:0] node1504;
	wire [4-1:0] node1507;
	wire [4-1:0] node1508;
	wire [4-1:0] node1509;
	wire [4-1:0] node1510;
	wire [4-1:0] node1511;
	wire [4-1:0] node1514;
	wire [4-1:0] node1518;
	wire [4-1:0] node1519;
	wire [4-1:0] node1520;
	wire [4-1:0] node1523;
	wire [4-1:0] node1526;
	wire [4-1:0] node1528;
	wire [4-1:0] node1531;
	wire [4-1:0] node1532;
	wire [4-1:0] node1533;
	wire [4-1:0] node1535;
	wire [4-1:0] node1538;
	wire [4-1:0] node1540;
	wire [4-1:0] node1543;
	wire [4-1:0] node1545;
	wire [4-1:0] node1548;
	wire [4-1:0] node1549;
	wire [4-1:0] node1550;
	wire [4-1:0] node1551;
	wire [4-1:0] node1552;
	wire [4-1:0] node1553;
	wire [4-1:0] node1555;
	wire [4-1:0] node1558;
	wire [4-1:0] node1559;
	wire [4-1:0] node1562;
	wire [4-1:0] node1565;
	wire [4-1:0] node1566;
	wire [4-1:0] node1567;
	wire [4-1:0] node1570;
	wire [4-1:0] node1573;
	wire [4-1:0] node1574;
	wire [4-1:0] node1577;
	wire [4-1:0] node1580;
	wire [4-1:0] node1581;
	wire [4-1:0] node1582;
	wire [4-1:0] node1583;
	wire [4-1:0] node1586;
	wire [4-1:0] node1589;
	wire [4-1:0] node1590;
	wire [4-1:0] node1593;
	wire [4-1:0] node1596;
	wire [4-1:0] node1597;
	wire [4-1:0] node1598;
	wire [4-1:0] node1599;
	wire [4-1:0] node1602;
	wire [4-1:0] node1605;
	wire [4-1:0] node1606;
	wire [4-1:0] node1610;
	wire [4-1:0] node1612;
	wire [4-1:0] node1615;
	wire [4-1:0] node1616;
	wire [4-1:0] node1617;
	wire [4-1:0] node1618;
	wire [4-1:0] node1619;
	wire [4-1:0] node1623;
	wire [4-1:0] node1624;
	wire [4-1:0] node1627;
	wire [4-1:0] node1630;
	wire [4-1:0] node1631;
	wire [4-1:0] node1632;
	wire [4-1:0] node1635;
	wire [4-1:0] node1638;
	wire [4-1:0] node1640;
	wire [4-1:0] node1643;
	wire [4-1:0] node1644;
	wire [4-1:0] node1646;
	wire [4-1:0] node1647;
	wire [4-1:0] node1648;
	wire [4-1:0] node1651;
	wire [4-1:0] node1654;
	wire [4-1:0] node1656;
	wire [4-1:0] node1659;
	wire [4-1:0] node1660;
	wire [4-1:0] node1662;
	wire [4-1:0] node1664;
	wire [4-1:0] node1667;
	wire [4-1:0] node1668;
	wire [4-1:0] node1669;
	wire [4-1:0] node1674;
	wire [4-1:0] node1675;
	wire [4-1:0] node1676;
	wire [4-1:0] node1677;
	wire [4-1:0] node1678;
	wire [4-1:0] node1679;
	wire [4-1:0] node1682;
	wire [4-1:0] node1685;
	wire [4-1:0] node1686;
	wire [4-1:0] node1687;
	wire [4-1:0] node1690;
	wire [4-1:0] node1693;
	wire [4-1:0] node1696;
	wire [4-1:0] node1697;
	wire [4-1:0] node1698;
	wire [4-1:0] node1699;
	wire [4-1:0] node1703;
	wire [4-1:0] node1704;
	wire [4-1:0] node1707;
	wire [4-1:0] node1710;
	wire [4-1:0] node1711;
	wire [4-1:0] node1712;
	wire [4-1:0] node1716;
	wire [4-1:0] node1717;
	wire [4-1:0] node1720;
	wire [4-1:0] node1723;
	wire [4-1:0] node1724;
	wire [4-1:0] node1725;
	wire [4-1:0] node1726;
	wire [4-1:0] node1729;
	wire [4-1:0] node1731;
	wire [4-1:0] node1734;
	wire [4-1:0] node1735;
	wire [4-1:0] node1738;
	wire [4-1:0] node1741;
	wire [4-1:0] node1742;
	wire [4-1:0] node1743;
	wire [4-1:0] node1745;
	wire [4-1:0] node1748;
	wire [4-1:0] node1750;
	wire [4-1:0] node1753;
	wire [4-1:0] node1754;
	wire [4-1:0] node1755;
	wire [4-1:0] node1759;
	wire [4-1:0] node1762;
	wire [4-1:0] node1763;
	wire [4-1:0] node1764;
	wire [4-1:0] node1765;
	wire [4-1:0] node1766;
	wire [4-1:0] node1767;
	wire [4-1:0] node1770;
	wire [4-1:0] node1774;
	wire [4-1:0] node1775;
	wire [4-1:0] node1776;
	wire [4-1:0] node1780;
	wire [4-1:0] node1782;
	wire [4-1:0] node1785;
	wire [4-1:0] node1786;
	wire [4-1:0] node1787;
	wire [4-1:0] node1789;
	wire [4-1:0] node1792;
	wire [4-1:0] node1795;
	wire [4-1:0] node1797;
	wire [4-1:0] node1800;
	wire [4-1:0] node1801;
	wire [4-1:0] node1802;
	wire [4-1:0] node1803;
	wire [4-1:0] node1804;
	wire [4-1:0] node1807;
	wire [4-1:0] node1810;
	wire [4-1:0] node1811;
	wire [4-1:0] node1814;
	wire [4-1:0] node1817;
	wire [4-1:0] node1818;
	wire [4-1:0] node1819;
	wire [4-1:0] node1822;
	wire [4-1:0] node1825;
	wire [4-1:0] node1827;
	wire [4-1:0] node1830;
	wire [4-1:0] node1831;
	wire [4-1:0] node1832;
	wire [4-1:0] node1833;
	wire [4-1:0] node1836;
	wire [4-1:0] node1840;
	wire [4-1:0] node1841;
	wire [4-1:0] node1843;
	wire [4-1:0] node1846;
	wire [4-1:0] node1847;
	wire [4-1:0] node1850;
	wire [4-1:0] node1853;
	wire [4-1:0] node1854;
	wire [4-1:0] node1855;
	wire [4-1:0] node1856;
	wire [4-1:0] node1857;
	wire [4-1:0] node1858;
	wire [4-1:0] node1859;
	wire [4-1:0] node1862;
	wire [4-1:0] node1865;
	wire [4-1:0] node1866;
	wire [4-1:0] node1867;
	wire [4-1:0] node1871;
	wire [4-1:0] node1873;
	wire [4-1:0] node1876;
	wire [4-1:0] node1877;
	wire [4-1:0] node1878;
	wire [4-1:0] node1881;
	wire [4-1:0] node1884;
	wire [4-1:0] node1885;
	wire [4-1:0] node1886;
	wire [4-1:0] node1889;
	wire [4-1:0] node1890;
	wire [4-1:0] node1894;
	wire [4-1:0] node1895;
	wire [4-1:0] node1896;
	wire [4-1:0] node1899;
	wire [4-1:0] node1902;
	wire [4-1:0] node1903;
	wire [4-1:0] node1906;
	wire [4-1:0] node1909;
	wire [4-1:0] node1910;
	wire [4-1:0] node1911;
	wire [4-1:0] node1912;
	wire [4-1:0] node1915;
	wire [4-1:0] node1918;
	wire [4-1:0] node1919;
	wire [4-1:0] node1920;
	wire [4-1:0] node1924;
	wire [4-1:0] node1926;
	wire [4-1:0] node1927;
	wire [4-1:0] node1930;
	wire [4-1:0] node1933;
	wire [4-1:0] node1934;
	wire [4-1:0] node1935;
	wire [4-1:0] node1936;
	wire [4-1:0] node1937;
	wire [4-1:0] node1940;
	wire [4-1:0] node1943;
	wire [4-1:0] node1944;
	wire [4-1:0] node1947;
	wire [4-1:0] node1951;
	wire [4-1:0] node1952;
	wire [4-1:0] node1954;
	wire [4-1:0] node1955;
	wire [4-1:0] node1959;
	wire [4-1:0] node1960;
	wire [4-1:0] node1961;
	wire [4-1:0] node1966;
	wire [4-1:0] node1967;
	wire [4-1:0] node1968;
	wire [4-1:0] node1969;
	wire [4-1:0] node1970;
	wire [4-1:0] node1971;
	wire [4-1:0] node1974;
	wire [4-1:0] node1975;
	wire [4-1:0] node1979;
	wire [4-1:0] node1981;
	wire [4-1:0] node1984;
	wire [4-1:0] node1985;
	wire [4-1:0] node1987;
	wire [4-1:0] node1988;
	wire [4-1:0] node1992;
	wire [4-1:0] node1993;
	wire [4-1:0] node1996;
	wire [4-1:0] node1999;
	wire [4-1:0] node2000;
	wire [4-1:0] node2001;
	wire [4-1:0] node2002;
	wire [4-1:0] node2005;
	wire [4-1:0] node2008;
	wire [4-1:0] node2009;
	wire [4-1:0] node2010;
	wire [4-1:0] node2013;
	wire [4-1:0] node2017;
	wire [4-1:0] node2018;
	wire [4-1:0] node2019;
	wire [4-1:0] node2022;
	wire [4-1:0] node2025;
	wire [4-1:0] node2026;
	wire [4-1:0] node2027;
	wire [4-1:0] node2030;
	wire [4-1:0] node2033;
	wire [4-1:0] node2034;
	wire [4-1:0] node2037;
	wire [4-1:0] node2040;
	wire [4-1:0] node2041;
	wire [4-1:0] node2042;
	wire [4-1:0] node2043;
	wire [4-1:0] node2044;
	wire [4-1:0] node2045;
	wire [4-1:0] node2048;
	wire [4-1:0] node2051;
	wire [4-1:0] node2052;
	wire [4-1:0] node2055;
	wire [4-1:0] node2058;
	wire [4-1:0] node2059;
	wire [4-1:0] node2061;
	wire [4-1:0] node2064;
	wire [4-1:0] node2066;
	wire [4-1:0] node2069;
	wire [4-1:0] node2070;
	wire [4-1:0] node2071;
	wire [4-1:0] node2072;
	wire [4-1:0] node2076;
	wire [4-1:0] node2078;
	wire [4-1:0] node2081;
	wire [4-1:0] node2083;
	wire [4-1:0] node2084;
	wire [4-1:0] node2087;
	wire [4-1:0] node2090;
	wire [4-1:0] node2091;
	wire [4-1:0] node2092;
	wire [4-1:0] node2093;
	wire [4-1:0] node2097;
	wire [4-1:0] node2098;
	wire [4-1:0] node2099;
	wire [4-1:0] node2103;
	wire [4-1:0] node2106;
	wire [4-1:0] node2107;
	wire [4-1:0] node2108;
	wire [4-1:0] node2111;
	wire [4-1:0] node2114;
	wire [4-1:0] node2116;
	wire [4-1:0] node2119;
	wire [4-1:0] node2120;
	wire [4-1:0] node2121;
	wire [4-1:0] node2122;
	wire [4-1:0] node2123;
	wire [4-1:0] node2124;
	wire [4-1:0] node2126;
	wire [4-1:0] node2129;
	wire [4-1:0] node2131;
	wire [4-1:0] node2134;
	wire [4-1:0] node2135;
	wire [4-1:0] node2137;
	wire [4-1:0] node2140;
	wire [4-1:0] node2143;
	wire [4-1:0] node2144;
	wire [4-1:0] node2145;
	wire [4-1:0] node2148;
	wire [4-1:0] node2151;
	wire [4-1:0] node2152;
	wire [4-1:0] node2153;
	wire [4-1:0] node2157;
	wire [4-1:0] node2158;
	wire [4-1:0] node2162;
	wire [4-1:0] node2163;
	wire [4-1:0] node2164;
	wire [4-1:0] node2165;
	wire [4-1:0] node2166;
	wire [4-1:0] node2170;
	wire [4-1:0] node2171;
	wire [4-1:0] node2174;
	wire [4-1:0] node2177;
	wire [4-1:0] node2178;
	wire [4-1:0] node2179;
	wire [4-1:0] node2183;
	wire [4-1:0] node2184;
	wire [4-1:0] node2185;
	wire [4-1:0] node2188;
	wire [4-1:0] node2191;
	wire [4-1:0] node2193;
	wire [4-1:0] node2196;
	wire [4-1:0] node2197;
	wire [4-1:0] node2198;
	wire [4-1:0] node2199;
	wire [4-1:0] node2202;
	wire [4-1:0] node2203;
	wire [4-1:0] node2207;
	wire [4-1:0] node2208;
	wire [4-1:0] node2211;
	wire [4-1:0] node2214;
	wire [4-1:0] node2215;
	wire [4-1:0] node2216;
	wire [4-1:0] node2217;
	wire [4-1:0] node2220;
	wire [4-1:0] node2223;
	wire [4-1:0] node2224;
	wire [4-1:0] node2227;
	wire [4-1:0] node2230;
	wire [4-1:0] node2232;
	wire [4-1:0] node2235;
	wire [4-1:0] node2236;
	wire [4-1:0] node2237;
	wire [4-1:0] node2238;
	wire [4-1:0] node2239;
	wire [4-1:0] node2240;
	wire [4-1:0] node2241;
	wire [4-1:0] node2244;
	wire [4-1:0] node2247;
	wire [4-1:0] node2248;
	wire [4-1:0] node2251;
	wire [4-1:0] node2254;
	wire [4-1:0] node2255;
	wire [4-1:0] node2256;
	wire [4-1:0] node2260;
	wire [4-1:0] node2261;
	wire [4-1:0] node2264;
	wire [4-1:0] node2267;
	wire [4-1:0] node2268;
	wire [4-1:0] node2269;
	wire [4-1:0] node2270;
	wire [4-1:0] node2273;
	wire [4-1:0] node2276;
	wire [4-1:0] node2278;
	wire [4-1:0] node2281;
	wire [4-1:0] node2282;
	wire [4-1:0] node2284;
	wire [4-1:0] node2287;
	wire [4-1:0] node2288;
	wire [4-1:0] node2291;
	wire [4-1:0] node2294;
	wire [4-1:0] node2295;
	wire [4-1:0] node2296;
	wire [4-1:0] node2297;
	wire [4-1:0] node2298;
	wire [4-1:0] node2302;
	wire [4-1:0] node2303;
	wire [4-1:0] node2307;
	wire [4-1:0] node2308;
	wire [4-1:0] node2312;
	wire [4-1:0] node2313;
	wire [4-1:0] node2314;
	wire [4-1:0] node2315;
	wire [4-1:0] node2319;
	wire [4-1:0] node2320;
	wire [4-1:0] node2324;
	wire [4-1:0] node2325;
	wire [4-1:0] node2327;
	wire [4-1:0] node2330;
	wire [4-1:0] node2331;
	wire [4-1:0] node2335;
	wire [4-1:0] node2336;
	wire [4-1:0] node2337;
	wire [4-1:0] node2338;
	wire [4-1:0] node2339;
	wire [4-1:0] node2341;
	wire [4-1:0] node2344;
	wire [4-1:0] node2345;
	wire [4-1:0] node2349;
	wire [4-1:0] node2350;
	wire [4-1:0] node2351;
	wire [4-1:0] node2354;
	wire [4-1:0] node2357;
	wire [4-1:0] node2358;
	wire [4-1:0] node2361;
	wire [4-1:0] node2364;
	wire [4-1:0] node2365;
	wire [4-1:0] node2366;
	wire [4-1:0] node2368;
	wire [4-1:0] node2371;
	wire [4-1:0] node2372;
	wire [4-1:0] node2375;
	wire [4-1:0] node2378;
	wire [4-1:0] node2379;
	wire [4-1:0] node2380;
	wire [4-1:0] node2383;
	wire [4-1:0] node2387;
	wire [4-1:0] node2388;
	wire [4-1:0] node2389;
	wire [4-1:0] node2390;
	wire [4-1:0] node2391;
	wire [4-1:0] node2395;
	wire [4-1:0] node2396;
	wire [4-1:0] node2400;
	wire [4-1:0] node2403;
	wire [4-1:0] node2404;
	wire [4-1:0] node2405;
	wire [4-1:0] node2406;
	wire [4-1:0] node2409;
	wire [4-1:0] node2412;
	wire [4-1:0] node2414;
	wire [4-1:0] node2417;
	wire [4-1:0] node2418;
	wire [4-1:0] node2420;
	wire [4-1:0] node2423;
	wire [4-1:0] node2424;
	wire [4-1:0] node2427;
	wire [4-1:0] node2430;
	wire [4-1:0] node2431;
	wire [4-1:0] node2432;
	wire [4-1:0] node2433;
	wire [4-1:0] node2434;
	wire [4-1:0] node2435;
	wire [4-1:0] node2436;
	wire [4-1:0] node2437;
	wire [4-1:0] node2438;
	wire [4-1:0] node2439;
	wire [4-1:0] node2440;
	wire [4-1:0] node2444;
	wire [4-1:0] node2445;
	wire [4-1:0] node2449;
	wire [4-1:0] node2450;
	wire [4-1:0] node2451;
	wire [4-1:0] node2454;
	wire [4-1:0] node2457;
	wire [4-1:0] node2458;
	wire [4-1:0] node2461;
	wire [4-1:0] node2464;
	wire [4-1:0] node2465;
	wire [4-1:0] node2466;
	wire [4-1:0] node2468;
	wire [4-1:0] node2471;
	wire [4-1:0] node2473;
	wire [4-1:0] node2476;
	wire [4-1:0] node2477;
	wire [4-1:0] node2478;
	wire [4-1:0] node2481;
	wire [4-1:0] node2485;
	wire [4-1:0] node2486;
	wire [4-1:0] node2487;
	wire [4-1:0] node2489;
	wire [4-1:0] node2490;
	wire [4-1:0] node2494;
	wire [4-1:0] node2495;
	wire [4-1:0] node2496;
	wire [4-1:0] node2499;
	wire [4-1:0] node2502;
	wire [4-1:0] node2503;
	wire [4-1:0] node2506;
	wire [4-1:0] node2509;
	wire [4-1:0] node2510;
	wire [4-1:0] node2512;
	wire [4-1:0] node2513;
	wire [4-1:0] node2517;
	wire [4-1:0] node2518;
	wire [4-1:0] node2522;
	wire [4-1:0] node2523;
	wire [4-1:0] node2524;
	wire [4-1:0] node2525;
	wire [4-1:0] node2528;
	wire [4-1:0] node2531;
	wire [4-1:0] node2532;
	wire [4-1:0] node2533;
	wire [4-1:0] node2536;
	wire [4-1:0] node2539;
	wire [4-1:0] node2541;
	wire [4-1:0] node2542;
	wire [4-1:0] node2545;
	wire [4-1:0] node2548;
	wire [4-1:0] node2549;
	wire [4-1:0] node2551;
	wire [4-1:0] node2552;
	wire [4-1:0] node2556;
	wire [4-1:0] node2557;
	wire [4-1:0] node2559;
	wire [4-1:0] node2560;
	wire [4-1:0] node2563;
	wire [4-1:0] node2566;
	wire [4-1:0] node2567;
	wire [4-1:0] node2570;
	wire [4-1:0] node2573;
	wire [4-1:0] node2574;
	wire [4-1:0] node2575;
	wire [4-1:0] node2576;
	wire [4-1:0] node2577;
	wire [4-1:0] node2578;
	wire [4-1:0] node2581;
	wire [4-1:0] node2584;
	wire [4-1:0] node2585;
	wire [4-1:0] node2588;
	wire [4-1:0] node2591;
	wire [4-1:0] node2592;
	wire [4-1:0] node2593;
	wire [4-1:0] node2596;
	wire [4-1:0] node2599;
	wire [4-1:0] node2600;
	wire [4-1:0] node2602;
	wire [4-1:0] node2605;
	wire [4-1:0] node2606;
	wire [4-1:0] node2610;
	wire [4-1:0] node2611;
	wire [4-1:0] node2612;
	wire [4-1:0] node2613;
	wire [4-1:0] node2616;
	wire [4-1:0] node2619;
	wire [4-1:0] node2621;
	wire [4-1:0] node2624;
	wire [4-1:0] node2625;
	wire [4-1:0] node2626;
	wire [4-1:0] node2629;
	wire [4-1:0] node2632;
	wire [4-1:0] node2633;
	wire [4-1:0] node2634;
	wire [4-1:0] node2639;
	wire [4-1:0] node2640;
	wire [4-1:0] node2641;
	wire [4-1:0] node2642;
	wire [4-1:0] node2645;
	wire [4-1:0] node2648;
	wire [4-1:0] node2649;
	wire [4-1:0] node2650;
	wire [4-1:0] node2653;
	wire [4-1:0] node2656;
	wire [4-1:0] node2657;
	wire [4-1:0] node2660;
	wire [4-1:0] node2663;
	wire [4-1:0] node2664;
	wire [4-1:0] node2665;
	wire [4-1:0] node2666;
	wire [4-1:0] node2669;
	wire [4-1:0] node2672;
	wire [4-1:0] node2673;
	wire [4-1:0] node2676;
	wire [4-1:0] node2679;
	wire [4-1:0] node2680;
	wire [4-1:0] node2683;
	wire [4-1:0] node2686;
	wire [4-1:0] node2687;
	wire [4-1:0] node2688;
	wire [4-1:0] node2689;
	wire [4-1:0] node2690;
	wire [4-1:0] node2691;
	wire [4-1:0] node2694;
	wire [4-1:0] node2697;
	wire [4-1:0] node2698;
	wire [4-1:0] node2699;
	wire [4-1:0] node2700;
	wire [4-1:0] node2703;
	wire [4-1:0] node2706;
	wire [4-1:0] node2707;
	wire [4-1:0] node2711;
	wire [4-1:0] node2712;
	wire [4-1:0] node2715;
	wire [4-1:0] node2718;
	wire [4-1:0] node2719;
	wire [4-1:0] node2720;
	wire [4-1:0] node2721;
	wire [4-1:0] node2723;
	wire [4-1:0] node2727;
	wire [4-1:0] node2728;
	wire [4-1:0] node2729;
	wire [4-1:0] node2733;
	wire [4-1:0] node2734;
	wire [4-1:0] node2737;
	wire [4-1:0] node2740;
	wire [4-1:0] node2741;
	wire [4-1:0] node2742;
	wire [4-1:0] node2744;
	wire [4-1:0] node2747;
	wire [4-1:0] node2749;
	wire [4-1:0] node2752;
	wire [4-1:0] node2753;
	wire [4-1:0] node2756;
	wire [4-1:0] node2759;
	wire [4-1:0] node2760;
	wire [4-1:0] node2761;
	wire [4-1:0] node2764;
	wire [4-1:0] node2767;
	wire [4-1:0] node2768;
	wire [4-1:0] node2769;
	wire [4-1:0] node2770;
	wire [4-1:0] node2774;
	wire [4-1:0] node2775;
	wire [4-1:0] node2778;
	wire [4-1:0] node2781;
	wire [4-1:0] node2782;
	wire [4-1:0] node2785;
	wire [4-1:0] node2788;
	wire [4-1:0] node2789;
	wire [4-1:0] node2790;
	wire [4-1:0] node2791;
	wire [4-1:0] node2792;
	wire [4-1:0] node2793;
	wire [4-1:0] node2794;
	wire [4-1:0] node2798;
	wire [4-1:0] node2799;
	wire [4-1:0] node2802;
	wire [4-1:0] node2805;
	wire [4-1:0] node2806;
	wire [4-1:0] node2809;
	wire [4-1:0] node2812;
	wire [4-1:0] node2813;
	wire [4-1:0] node2814;
	wire [4-1:0] node2817;
	wire [4-1:0] node2820;
	wire [4-1:0] node2822;
	wire [4-1:0] node2825;
	wire [4-1:0] node2826;
	wire [4-1:0] node2827;
	wire [4-1:0] node2828;
	wire [4-1:0] node2831;
	wire [4-1:0] node2834;
	wire [4-1:0] node2835;
	wire [4-1:0] node2838;
	wire [4-1:0] node2841;
	wire [4-1:0] node2842;
	wire [4-1:0] node2844;
	wire [4-1:0] node2845;
	wire [4-1:0] node2848;
	wire [4-1:0] node2851;
	wire [4-1:0] node2853;
	wire [4-1:0] node2856;
	wire [4-1:0] node2857;
	wire [4-1:0] node2858;
	wire [4-1:0] node2859;
	wire [4-1:0] node2860;
	wire [4-1:0] node2861;
	wire [4-1:0] node2864;
	wire [4-1:0] node2867;
	wire [4-1:0] node2869;
	wire [4-1:0] node2872;
	wire [4-1:0] node2873;
	wire [4-1:0] node2876;
	wire [4-1:0] node2879;
	wire [4-1:0] node2880;
	wire [4-1:0] node2882;
	wire [4-1:0] node2884;
	wire [4-1:0] node2887;
	wire [4-1:0] node2889;
	wire [4-1:0] node2892;
	wire [4-1:0] node2893;
	wire [4-1:0] node2894;
	wire [4-1:0] node2895;
	wire [4-1:0] node2898;
	wire [4-1:0] node2901;
	wire [4-1:0] node2902;
	wire [4-1:0] node2905;
	wire [4-1:0] node2908;
	wire [4-1:0] node2909;
	wire [4-1:0] node2911;
	wire [4-1:0] node2914;
	wire [4-1:0] node2915;
	wire [4-1:0] node2918;
	wire [4-1:0] node2921;
	wire [4-1:0] node2922;
	wire [4-1:0] node2923;
	wire [4-1:0] node2924;
	wire [4-1:0] node2925;
	wire [4-1:0] node2926;
	wire [4-1:0] node2927;
	wire [4-1:0] node2928;
	wire [4-1:0] node2931;
	wire [4-1:0] node2934;
	wire [4-1:0] node2936;
	wire [4-1:0] node2937;
	wire [4-1:0] node2940;
	wire [4-1:0] node2943;
	wire [4-1:0] node2944;
	wire [4-1:0] node2945;
	wire [4-1:0] node2948;
	wire [4-1:0] node2951;
	wire [4-1:0] node2952;
	wire [4-1:0] node2954;
	wire [4-1:0] node2958;
	wire [4-1:0] node2959;
	wire [4-1:0] node2960;
	wire [4-1:0] node2961;
	wire [4-1:0] node2964;
	wire [4-1:0] node2967;
	wire [4-1:0] node2968;
	wire [4-1:0] node2970;
	wire [4-1:0] node2973;
	wire [4-1:0] node2975;
	wire [4-1:0] node2978;
	wire [4-1:0] node2979;
	wire [4-1:0] node2980;
	wire [4-1:0] node2983;
	wire [4-1:0] node2986;
	wire [4-1:0] node2987;
	wire [4-1:0] node2988;
	wire [4-1:0] node2991;
	wire [4-1:0] node2994;
	wire [4-1:0] node2995;
	wire [4-1:0] node2999;
	wire [4-1:0] node3000;
	wire [4-1:0] node3001;
	wire [4-1:0] node3002;
	wire [4-1:0] node3003;
	wire [4-1:0] node3006;
	wire [4-1:0] node3009;
	wire [4-1:0] node3010;
	wire [4-1:0] node3013;
	wire [4-1:0] node3016;
	wire [4-1:0] node3017;
	wire [4-1:0] node3018;
	wire [4-1:0] node3021;
	wire [4-1:0] node3024;
	wire [4-1:0] node3025;
	wire [4-1:0] node3026;
	wire [4-1:0] node3029;
	wire [4-1:0] node3032;
	wire [4-1:0] node3033;
	wire [4-1:0] node3036;
	wire [4-1:0] node3039;
	wire [4-1:0] node3040;
	wire [4-1:0] node3041;
	wire [4-1:0] node3042;
	wire [4-1:0] node3045;
	wire [4-1:0] node3048;
	wire [4-1:0] node3049;
	wire [4-1:0] node3053;
	wire [4-1:0] node3055;
	wire [4-1:0] node3057;
	wire [4-1:0] node3058;
	wire [4-1:0] node3061;
	wire [4-1:0] node3064;
	wire [4-1:0] node3065;
	wire [4-1:0] node3066;
	wire [4-1:0] node3067;
	wire [4-1:0] node3068;
	wire [4-1:0] node3071;
	wire [4-1:0] node3074;
	wire [4-1:0] node3075;
	wire [4-1:0] node3076;
	wire [4-1:0] node3077;
	wire [4-1:0] node3080;
	wire [4-1:0] node3083;
	wire [4-1:0] node3084;
	wire [4-1:0] node3087;
	wire [4-1:0] node3090;
	wire [4-1:0] node3091;
	wire [4-1:0] node3092;
	wire [4-1:0] node3095;
	wire [4-1:0] node3099;
	wire [4-1:0] node3100;
	wire [4-1:0] node3101;
	wire [4-1:0] node3102;
	wire [4-1:0] node3106;
	wire [4-1:0] node3107;
	wire [4-1:0] node3109;
	wire [4-1:0] node3112;
	wire [4-1:0] node3114;
	wire [4-1:0] node3117;
	wire [4-1:0] node3118;
	wire [4-1:0] node3119;
	wire [4-1:0] node3122;
	wire [4-1:0] node3125;
	wire [4-1:0] node3126;
	wire [4-1:0] node3129;
	wire [4-1:0] node3132;
	wire [4-1:0] node3133;
	wire [4-1:0] node3134;
	wire [4-1:0] node3135;
	wire [4-1:0] node3136;
	wire [4-1:0] node3140;
	wire [4-1:0] node3141;
	wire [4-1:0] node3143;
	wire [4-1:0] node3146;
	wire [4-1:0] node3147;
	wire [4-1:0] node3150;
	wire [4-1:0] node3153;
	wire [4-1:0] node3154;
	wire [4-1:0] node3155;
	wire [4-1:0] node3158;
	wire [4-1:0] node3161;
	wire [4-1:0] node3162;
	wire [4-1:0] node3165;
	wire [4-1:0] node3168;
	wire [4-1:0] node3169;
	wire [4-1:0] node3170;
	wire [4-1:0] node3171;
	wire [4-1:0] node3172;
	wire [4-1:0] node3175;
	wire [4-1:0] node3178;
	wire [4-1:0] node3179;
	wire [4-1:0] node3183;
	wire [4-1:0] node3185;
	wire [4-1:0] node3186;
	wire [4-1:0] node3189;
	wire [4-1:0] node3192;
	wire [4-1:0] node3193;
	wire [4-1:0] node3194;
	wire [4-1:0] node3197;
	wire [4-1:0] node3200;
	wire [4-1:0] node3201;
	wire [4-1:0] node3204;
	wire [4-1:0] node3207;
	wire [4-1:0] node3208;
	wire [4-1:0] node3209;
	wire [4-1:0] node3210;
	wire [4-1:0] node3211;
	wire [4-1:0] node3212;
	wire [4-1:0] node3213;
	wire [4-1:0] node3216;
	wire [4-1:0] node3219;
	wire [4-1:0] node3220;
	wire [4-1:0] node3224;
	wire [4-1:0] node3225;
	wire [4-1:0] node3226;
	wire [4-1:0] node3229;
	wire [4-1:0] node3232;
	wire [4-1:0] node3234;
	wire [4-1:0] node3237;
	wire [4-1:0] node3238;
	wire [4-1:0] node3239;
	wire [4-1:0] node3242;
	wire [4-1:0] node3245;
	wire [4-1:0] node3246;
	wire [4-1:0] node3247;
	wire [4-1:0] node3249;
	wire [4-1:0] node3252;
	wire [4-1:0] node3253;
	wire [4-1:0] node3256;
	wire [4-1:0] node3260;
	wire [4-1:0] node3261;
	wire [4-1:0] node3262;
	wire [4-1:0] node3263;
	wire [4-1:0] node3265;
	wire [4-1:0] node3268;
	wire [4-1:0] node3269;
	wire [4-1:0] node3272;
	wire [4-1:0] node3275;
	wire [4-1:0] node3276;
	wire [4-1:0] node3277;
	wire [4-1:0] node3278;
	wire [4-1:0] node3281;
	wire [4-1:0] node3285;
	wire [4-1:0] node3286;
	wire [4-1:0] node3289;
	wire [4-1:0] node3292;
	wire [4-1:0] node3293;
	wire [4-1:0] node3294;
	wire [4-1:0] node3295;
	wire [4-1:0] node3298;
	wire [4-1:0] node3301;
	wire [4-1:0] node3302;
	wire [4-1:0] node3305;
	wire [4-1:0] node3308;
	wire [4-1:0] node3309;
	wire [4-1:0] node3312;
	wire [4-1:0] node3315;
	wire [4-1:0] node3316;
	wire [4-1:0] node3317;
	wire [4-1:0] node3318;
	wire [4-1:0] node3319;
	wire [4-1:0] node3320;
	wire [4-1:0] node3321;
	wire [4-1:0] node3325;
	wire [4-1:0] node3327;
	wire [4-1:0] node3330;
	wire [4-1:0] node3332;
	wire [4-1:0] node3335;
	wire [4-1:0] node3336;
	wire [4-1:0] node3339;
	wire [4-1:0] node3340;
	wire [4-1:0] node3342;
	wire [4-1:0] node3345;
	wire [4-1:0] node3346;
	wire [4-1:0] node3349;
	wire [4-1:0] node3352;
	wire [4-1:0] node3353;
	wire [4-1:0] node3354;
	wire [4-1:0] node3355;
	wire [4-1:0] node3356;
	wire [4-1:0] node3360;
	wire [4-1:0] node3362;
	wire [4-1:0] node3365;
	wire [4-1:0] node3366;
	wire [4-1:0] node3367;
	wire [4-1:0] node3372;
	wire [4-1:0] node3373;
	wire [4-1:0] node3374;
	wire [4-1:0] node3375;
	wire [4-1:0] node3378;
	wire [4-1:0] node3381;
	wire [4-1:0] node3382;
	wire [4-1:0] node3385;
	wire [4-1:0] node3388;
	wire [4-1:0] node3389;
	wire [4-1:0] node3390;
	wire [4-1:0] node3393;
	wire [4-1:0] node3396;
	wire [4-1:0] node3398;
	wire [4-1:0] node3401;
	wire [4-1:0] node3402;
	wire [4-1:0] node3403;
	wire [4-1:0] node3404;
	wire [4-1:0] node3405;
	wire [4-1:0] node3408;
	wire [4-1:0] node3411;
	wire [4-1:0] node3412;
	wire [4-1:0] node3415;
	wire [4-1:0] node3418;
	wire [4-1:0] node3419;
	wire [4-1:0] node3420;
	wire [4-1:0] node3421;
	wire [4-1:0] node3424;
	wire [4-1:0] node3427;
	wire [4-1:0] node3429;
	wire [4-1:0] node3432;
	wire [4-1:0] node3433;
	wire [4-1:0] node3436;
	wire [4-1:0] node3439;
	wire [4-1:0] node3440;
	wire [4-1:0] node3441;
	wire [4-1:0] node3442;
	wire [4-1:0] node3444;
	wire [4-1:0] node3447;
	wire [4-1:0] node3448;
	wire [4-1:0] node3451;
	wire [4-1:0] node3454;
	wire [4-1:0] node3455;
	wire [4-1:0] node3457;
	wire [4-1:0] node3460;
	wire [4-1:0] node3463;
	wire [4-1:0] node3464;
	wire [4-1:0] node3465;
	wire [4-1:0] node3467;
	wire [4-1:0] node3470;
	wire [4-1:0] node3471;
	wire [4-1:0] node3475;
	wire [4-1:0] node3476;
	wire [4-1:0] node3477;
	wire [4-1:0] node3480;
	wire [4-1:0] node3483;
	wire [4-1:0] node3484;
	wire [4-1:0] node3487;
	wire [4-1:0] node3490;
	wire [4-1:0] node3491;
	wire [4-1:0] node3492;
	wire [4-1:0] node3493;
	wire [4-1:0] node3494;
	wire [4-1:0] node3495;
	wire [4-1:0] node3496;
	wire [4-1:0] node3497;
	wire [4-1:0] node3498;
	wire [4-1:0] node3500;
	wire [4-1:0] node3503;
	wire [4-1:0] node3504;
	wire [4-1:0] node3507;
	wire [4-1:0] node3510;
	wire [4-1:0] node3511;
	wire [4-1:0] node3514;
	wire [4-1:0] node3517;
	wire [4-1:0] node3518;
	wire [4-1:0] node3521;
	wire [4-1:0] node3524;
	wire [4-1:0] node3525;
	wire [4-1:0] node3526;
	wire [4-1:0] node3527;
	wire [4-1:0] node3528;
	wire [4-1:0] node3532;
	wire [4-1:0] node3535;
	wire [4-1:0] node3536;
	wire [4-1:0] node3537;
	wire [4-1:0] node3540;
	wire [4-1:0] node3543;
	wire [4-1:0] node3545;
	wire [4-1:0] node3548;
	wire [4-1:0] node3549;
	wire [4-1:0] node3550;
	wire [4-1:0] node3554;
	wire [4-1:0] node3555;
	wire [4-1:0] node3558;
	wire [4-1:0] node3561;
	wire [4-1:0] node3562;
	wire [4-1:0] node3563;
	wire [4-1:0] node3564;
	wire [4-1:0] node3565;
	wire [4-1:0] node3566;
	wire [4-1:0] node3569;
	wire [4-1:0] node3572;
	wire [4-1:0] node3573;
	wire [4-1:0] node3576;
	wire [4-1:0] node3579;
	wire [4-1:0] node3580;
	wire [4-1:0] node3581;
	wire [4-1:0] node3584;
	wire [4-1:0] node3587;
	wire [4-1:0] node3589;
	wire [4-1:0] node3592;
	wire [4-1:0] node3593;
	wire [4-1:0] node3594;
	wire [4-1:0] node3595;
	wire [4-1:0] node3598;
	wire [4-1:0] node3601;
	wire [4-1:0] node3602;
	wire [4-1:0] node3605;
	wire [4-1:0] node3608;
	wire [4-1:0] node3609;
	wire [4-1:0] node3612;
	wire [4-1:0] node3615;
	wire [4-1:0] node3616;
	wire [4-1:0] node3617;
	wire [4-1:0] node3618;
	wire [4-1:0] node3619;
	wire [4-1:0] node3622;
	wire [4-1:0] node3625;
	wire [4-1:0] node3627;
	wire [4-1:0] node3630;
	wire [4-1:0] node3631;
	wire [4-1:0] node3632;
	wire [4-1:0] node3637;
	wire [4-1:0] node3638;
	wire [4-1:0] node3641;
	wire [4-1:0] node3644;
	wire [4-1:0] node3645;
	wire [4-1:0] node3646;
	wire [4-1:0] node3647;
	wire [4-1:0] node3648;
	wire [4-1:0] node3651;
	wire [4-1:0] node3654;
	wire [4-1:0] node3655;
	wire [4-1:0] node3658;
	wire [4-1:0] node3661;
	wire [4-1:0] node3662;
	wire [4-1:0] node3663;
	wire [4-1:0] node3665;
	wire [4-1:0] node3668;
	wire [4-1:0] node3669;
	wire [4-1:0] node3672;
	wire [4-1:0] node3675;
	wire [4-1:0] node3676;
	wire [4-1:0] node3679;
	wire [4-1:0] node3682;
	wire [4-1:0] node3683;
	wire [4-1:0] node3684;
	wire [4-1:0] node3685;
	wire [4-1:0] node3688;
	wire [4-1:0] node3691;
	wire [4-1:0] node3692;
	wire [4-1:0] node3695;
	wire [4-1:0] node3698;
	wire [4-1:0] node3699;
	wire [4-1:0] node3700;
	wire [4-1:0] node3703;
	wire [4-1:0] node3706;
	wire [4-1:0] node3707;
	wire [4-1:0] node3710;
	wire [4-1:0] node3713;
	wire [4-1:0] node3714;
	wire [4-1:0] node3715;
	wire [4-1:0] node3716;
	wire [4-1:0] node3717;
	wire [4-1:0] node3718;
	wire [4-1:0] node3721;
	wire [4-1:0] node3723;
	wire [4-1:0] node3724;
	wire [4-1:0] node3727;
	wire [4-1:0] node3730;
	wire [4-1:0] node3731;
	wire [4-1:0] node3732;
	wire [4-1:0] node3736;
	wire [4-1:0] node3737;
	wire [4-1:0] node3739;
	wire [4-1:0] node3742;
	wire [4-1:0] node3744;
	wire [4-1:0] node3747;
	wire [4-1:0] node3748;
	wire [4-1:0] node3749;
	wire [4-1:0] node3750;
	wire [4-1:0] node3752;
	wire [4-1:0] node3755;
	wire [4-1:0] node3757;
	wire [4-1:0] node3760;
	wire [4-1:0] node3762;
	wire [4-1:0] node3765;
	wire [4-1:0] node3766;
	wire [4-1:0] node3769;
	wire [4-1:0] node3770;
	wire [4-1:0] node3771;
	wire [4-1:0] node3774;
	wire [4-1:0] node3777;
	wire [4-1:0] node3778;
	wire [4-1:0] node3782;
	wire [4-1:0] node3783;
	wire [4-1:0] node3784;
	wire [4-1:0] node3785;
	wire [4-1:0] node3786;
	wire [4-1:0] node3789;
	wire [4-1:0] node3791;
	wire [4-1:0] node3794;
	wire [4-1:0] node3796;
	wire [4-1:0] node3798;
	wire [4-1:0] node3801;
	wire [4-1:0] node3802;
	wire [4-1:0] node3803;
	wire [4-1:0] node3805;
	wire [4-1:0] node3808;
	wire [4-1:0] node3810;
	wire [4-1:0] node3814;
	wire [4-1:0] node3815;
	wire [4-1:0] node3816;
	wire [4-1:0] node3817;
	wire [4-1:0] node3821;
	wire [4-1:0] node3822;
	wire [4-1:0] node3823;
	wire [4-1:0] node3826;
	wire [4-1:0] node3829;
	wire [4-1:0] node3830;
	wire [4-1:0] node3834;
	wire [4-1:0] node3835;
	wire [4-1:0] node3836;
	wire [4-1:0] node3840;
	wire [4-1:0] node3841;
	wire [4-1:0] node3843;
	wire [4-1:0] node3846;
	wire [4-1:0] node3848;
	wire [4-1:0] node3851;
	wire [4-1:0] node3852;
	wire [4-1:0] node3853;
	wire [4-1:0] node3854;
	wire [4-1:0] node3855;
	wire [4-1:0] node3856;
	wire [4-1:0] node3858;
	wire [4-1:0] node3861;
	wire [4-1:0] node3863;
	wire [4-1:0] node3866;
	wire [4-1:0] node3867;
	wire [4-1:0] node3869;
	wire [4-1:0] node3873;
	wire [4-1:0] node3874;
	wire [4-1:0] node3875;
	wire [4-1:0] node3877;
	wire [4-1:0] node3880;
	wire [4-1:0] node3882;
	wire [4-1:0] node3885;
	wire [4-1:0] node3886;
	wire [4-1:0] node3888;
	wire [4-1:0] node3891;
	wire [4-1:0] node3893;
	wire [4-1:0] node3896;
	wire [4-1:0] node3897;
	wire [4-1:0] node3898;
	wire [4-1:0] node3899;
	wire [4-1:0] node3903;
	wire [4-1:0] node3905;
	wire [4-1:0] node3908;
	wire [4-1:0] node3909;
	wire [4-1:0] node3910;
	wire [4-1:0] node3912;
	wire [4-1:0] node3915;
	wire [4-1:0] node3917;
	wire [4-1:0] node3920;
	wire [4-1:0] node3921;
	wire [4-1:0] node3925;
	wire [4-1:0] node3926;
	wire [4-1:0] node3927;
	wire [4-1:0] node3928;
	wire [4-1:0] node3929;
	wire [4-1:0] node3930;
	wire [4-1:0] node3933;
	wire [4-1:0] node3936;
	wire [4-1:0] node3937;
	wire [4-1:0] node3940;
	wire [4-1:0] node3943;
	wire [4-1:0] node3944;
	wire [4-1:0] node3945;
	wire [4-1:0] node3948;
	wire [4-1:0] node3952;
	wire [4-1:0] node3953;
	wire [4-1:0] node3954;
	wire [4-1:0] node3955;
	wire [4-1:0] node3959;
	wire [4-1:0] node3961;
	wire [4-1:0] node3964;
	wire [4-1:0] node3965;
	wire [4-1:0] node3968;
	wire [4-1:0] node3970;
	wire [4-1:0] node3973;
	wire [4-1:0] node3974;
	wire [4-1:0] node3975;
	wire [4-1:0] node3976;
	wire [4-1:0] node3979;
	wire [4-1:0] node3982;
	wire [4-1:0] node3983;
	wire [4-1:0] node3984;
	wire [4-1:0] node3988;
	wire [4-1:0] node3989;
	wire [4-1:0] node3993;
	wire [4-1:0] node3994;
	wire [4-1:0] node3995;
	wire [4-1:0] node3998;
	wire [4-1:0] node4001;
	wire [4-1:0] node4003;
	wire [4-1:0] node4004;
	wire [4-1:0] node4008;
	wire [4-1:0] node4009;
	wire [4-1:0] node4010;
	wire [4-1:0] node4011;
	wire [4-1:0] node4012;
	wire [4-1:0] node4013;
	wire [4-1:0] node4014;
	wire [4-1:0] node4017;
	wire [4-1:0] node4020;
	wire [4-1:0] node4021;
	wire [4-1:0] node4023;
	wire [4-1:0] node4026;
	wire [4-1:0] node4027;
	wire [4-1:0] node4031;
	wire [4-1:0] node4032;
	wire [4-1:0] node4033;
	wire [4-1:0] node4036;
	wire [4-1:0] node4039;
	wire [4-1:0] node4040;
	wire [4-1:0] node4041;
	wire [4-1:0] node4044;
	wire [4-1:0] node4045;
	wire [4-1:0] node4049;
	wire [4-1:0] node4050;
	wire [4-1:0] node4054;
	wire [4-1:0] node4055;
	wire [4-1:0] node4056;
	wire [4-1:0] node4057;
	wire [4-1:0] node4060;
	wire [4-1:0] node4063;
	wire [4-1:0] node4064;
	wire [4-1:0] node4065;
	wire [4-1:0] node4068;
	wire [4-1:0] node4072;
	wire [4-1:0] node4073;
	wire [4-1:0] node4074;
	wire [4-1:0] node4077;
	wire [4-1:0] node4080;
	wire [4-1:0] node4081;
	wire [4-1:0] node4082;
	wire [4-1:0] node4086;
	wire [4-1:0] node4087;
	wire [4-1:0] node4088;
	wire [4-1:0] node4091;
	wire [4-1:0] node4095;
	wire [4-1:0] node4096;
	wire [4-1:0] node4097;
	wire [4-1:0] node4098;
	wire [4-1:0] node4099;
	wire [4-1:0] node4100;
	wire [4-1:0] node4104;
	wire [4-1:0] node4105;
	wire [4-1:0] node4108;
	wire [4-1:0] node4110;
	wire [4-1:0] node4113;
	wire [4-1:0] node4114;
	wire [4-1:0] node4115;
	wire [4-1:0] node4116;
	wire [4-1:0] node4120;
	wire [4-1:0] node4122;
	wire [4-1:0] node4125;
	wire [4-1:0] node4126;
	wire [4-1:0] node4129;
	wire [4-1:0] node4130;
	wire [4-1:0] node4133;
	wire [4-1:0] node4136;
	wire [4-1:0] node4137;
	wire [4-1:0] node4138;
	wire [4-1:0] node4139;
	wire [4-1:0] node4140;
	wire [4-1:0] node4145;
	wire [4-1:0] node4146;
	wire [4-1:0] node4148;
	wire [4-1:0] node4151;
	wire [4-1:0] node4152;
	wire [4-1:0] node4155;
	wire [4-1:0] node4158;
	wire [4-1:0] node4159;
	wire [4-1:0] node4160;
	wire [4-1:0] node4161;
	wire [4-1:0] node4164;
	wire [4-1:0] node4167;
	wire [4-1:0] node4169;
	wire [4-1:0] node4172;
	wire [4-1:0] node4173;
	wire [4-1:0] node4175;
	wire [4-1:0] node4178;
	wire [4-1:0] node4179;
	wire [4-1:0] node4182;
	wire [4-1:0] node4185;
	wire [4-1:0] node4186;
	wire [4-1:0] node4187;
	wire [4-1:0] node4188;
	wire [4-1:0] node4189;
	wire [4-1:0] node4190;
	wire [4-1:0] node4193;
	wire [4-1:0] node4197;
	wire [4-1:0] node4198;
	wire [4-1:0] node4200;
	wire [4-1:0] node4203;
	wire [4-1:0] node4204;
	wire [4-1:0] node4208;
	wire [4-1:0] node4209;
	wire [4-1:0] node4211;
	wire [4-1:0] node4212;
	wire [4-1:0] node4215;
	wire [4-1:0] node4218;
	wire [4-1:0] node4219;
	wire [4-1:0] node4222;
	wire [4-1:0] node4225;
	wire [4-1:0] node4226;
	wire [4-1:0] node4227;
	wire [4-1:0] node4228;
	wire [4-1:0] node4231;
	wire [4-1:0] node4234;
	wire [4-1:0] node4235;
	wire [4-1:0] node4238;
	wire [4-1:0] node4241;
	wire [4-1:0] node4242;
	wire [4-1:0] node4243;
	wire [4-1:0] node4246;
	wire [4-1:0] node4248;
	wire [4-1:0] node4251;
	wire [4-1:0] node4253;
	wire [4-1:0] node4256;
	wire [4-1:0] node4257;
	wire [4-1:0] node4258;
	wire [4-1:0] node4259;
	wire [4-1:0] node4260;
	wire [4-1:0] node4261;
	wire [4-1:0] node4262;
	wire [4-1:0] node4264;
	wire [4-1:0] node4268;
	wire [4-1:0] node4270;
	wire [4-1:0] node4273;
	wire [4-1:0] node4274;
	wire [4-1:0] node4276;
	wire [4-1:0] node4279;
	wire [4-1:0] node4281;
	wire [4-1:0] node4284;
	wire [4-1:0] node4285;
	wire [4-1:0] node4286;
	wire [4-1:0] node4287;
	wire [4-1:0] node4289;
	wire [4-1:0] node4292;
	wire [4-1:0] node4293;
	wire [4-1:0] node4296;
	wire [4-1:0] node4299;
	wire [4-1:0] node4300;
	wire [4-1:0] node4303;
	wire [4-1:0] node4306;
	wire [4-1:0] node4307;
	wire [4-1:0] node4308;
	wire [4-1:0] node4311;
	wire [4-1:0] node4314;
	wire [4-1:0] node4315;
	wire [4-1:0] node4318;
	wire [4-1:0] node4321;
	wire [4-1:0] node4322;
	wire [4-1:0] node4323;
	wire [4-1:0] node4324;
	wire [4-1:0] node4326;
	wire [4-1:0] node4329;
	wire [4-1:0] node4331;
	wire [4-1:0] node4334;
	wire [4-1:0] node4335;
	wire [4-1:0] node4339;
	wire [4-1:0] node4340;
	wire [4-1:0] node4341;
	wire [4-1:0] node4343;
	wire [4-1:0] node4346;
	wire [4-1:0] node4348;
	wire [4-1:0] node4351;
	wire [4-1:0] node4352;
	wire [4-1:0] node4354;
	wire [4-1:0] node4357;
	wire [4-1:0] node4359;
	wire [4-1:0] node4362;
	wire [4-1:0] node4363;
	wire [4-1:0] node4364;
	wire [4-1:0] node4365;
	wire [4-1:0] node4366;
	wire [4-1:0] node4368;
	wire [4-1:0] node4371;
	wire [4-1:0] node4373;
	wire [4-1:0] node4376;
	wire [4-1:0] node4377;
	wire [4-1:0] node4379;
	wire [4-1:0] node4382;
	wire [4-1:0] node4384;
	wire [4-1:0] node4387;
	wire [4-1:0] node4388;
	wire [4-1:0] node4389;
	wire [4-1:0] node4390;
	wire [4-1:0] node4393;
	wire [4-1:0] node4396;
	wire [4-1:0] node4397;
	wire [4-1:0] node4400;
	wire [4-1:0] node4403;
	wire [4-1:0] node4404;
	wire [4-1:0] node4405;
	wire [4-1:0] node4406;
	wire [4-1:0] node4411;
	wire [4-1:0] node4412;
	wire [4-1:0] node4413;
	wire [4-1:0] node4416;
	wire [4-1:0] node4419;
	wire [4-1:0] node4420;
	wire [4-1:0] node4423;
	wire [4-1:0] node4426;
	wire [4-1:0] node4427;
	wire [4-1:0] node4428;
	wire [4-1:0] node4429;
	wire [4-1:0] node4432;
	wire [4-1:0] node4434;
	wire [4-1:0] node4437;
	wire [4-1:0] node4438;
	wire [4-1:0] node4440;
	wire [4-1:0] node4443;
	wire [4-1:0] node4445;
	wire [4-1:0] node4448;
	wire [4-1:0] node4449;
	wire [4-1:0] node4450;
	wire [4-1:0] node4451;
	wire [4-1:0] node4454;
	wire [4-1:0] node4457;
	wire [4-1:0] node4459;
	wire [4-1:0] node4462;
	wire [4-1:0] node4463;
	wire [4-1:0] node4464;
	wire [4-1:0] node4467;
	wire [4-1:0] node4470;
	wire [4-1:0] node4471;
	wire [4-1:0] node4475;
	wire [4-1:0] node4476;
	wire [4-1:0] node4477;
	wire [4-1:0] node4478;
	wire [4-1:0] node4479;
	wire [4-1:0] node4480;
	wire [4-1:0] node4481;
	wire [4-1:0] node4482;
	wire [4-1:0] node4483;
	wire [4-1:0] node4484;
	wire [4-1:0] node4486;
	wire [4-1:0] node4489;
	wire [4-1:0] node4491;
	wire [4-1:0] node4494;
	wire [4-1:0] node4495;
	wire [4-1:0] node4496;
	wire [4-1:0] node4498;
	wire [4-1:0] node4502;
	wire [4-1:0] node4503;
	wire [4-1:0] node4506;
	wire [4-1:0] node4509;
	wire [4-1:0] node4510;
	wire [4-1:0] node4511;
	wire [4-1:0] node4513;
	wire [4-1:0] node4515;
	wire [4-1:0] node4518;
	wire [4-1:0] node4519;
	wire [4-1:0] node4523;
	wire [4-1:0] node4524;
	wire [4-1:0] node4525;
	wire [4-1:0] node4527;
	wire [4-1:0] node4530;
	wire [4-1:0] node4533;
	wire [4-1:0] node4534;
	wire [4-1:0] node4538;
	wire [4-1:0] node4539;
	wire [4-1:0] node4540;
	wire [4-1:0] node4541;
	wire [4-1:0] node4542;
	wire [4-1:0] node4543;
	wire [4-1:0] node4546;
	wire [4-1:0] node4549;
	wire [4-1:0] node4550;
	wire [4-1:0] node4553;
	wire [4-1:0] node4556;
	wire [4-1:0] node4557;
	wire [4-1:0] node4558;
	wire [4-1:0] node4561;
	wire [4-1:0] node4564;
	wire [4-1:0] node4565;
	wire [4-1:0] node4568;
	wire [4-1:0] node4571;
	wire [4-1:0] node4572;
	wire [4-1:0] node4573;
	wire [4-1:0] node4575;
	wire [4-1:0] node4578;
	wire [4-1:0] node4580;
	wire [4-1:0] node4583;
	wire [4-1:0] node4584;
	wire [4-1:0] node4588;
	wire [4-1:0] node4589;
	wire [4-1:0] node4590;
	wire [4-1:0] node4591;
	wire [4-1:0] node4593;
	wire [4-1:0] node4596;
	wire [4-1:0] node4599;
	wire [4-1:0] node4600;
	wire [4-1:0] node4603;
	wire [4-1:0] node4605;
	wire [4-1:0] node4608;
	wire [4-1:0] node4609;
	wire [4-1:0] node4610;
	wire [4-1:0] node4614;
	wire [4-1:0] node4615;
	wire [4-1:0] node4619;
	wire [4-1:0] node4620;
	wire [4-1:0] node4621;
	wire [4-1:0] node4622;
	wire [4-1:0] node4623;
	wire [4-1:0] node4624;
	wire [4-1:0] node4626;
	wire [4-1:0] node4629;
	wire [4-1:0] node4631;
	wire [4-1:0] node4634;
	wire [4-1:0] node4635;
	wire [4-1:0] node4639;
	wire [4-1:0] node4640;
	wire [4-1:0] node4643;
	wire [4-1:0] node4644;
	wire [4-1:0] node4646;
	wire [4-1:0] node4649;
	wire [4-1:0] node4651;
	wire [4-1:0] node4654;
	wire [4-1:0] node4655;
	wire [4-1:0] node4656;
	wire [4-1:0] node4658;
	wire [4-1:0] node4659;
	wire [4-1:0] node4662;
	wire [4-1:0] node4665;
	wire [4-1:0] node4666;
	wire [4-1:0] node4668;
	wire [4-1:0] node4671;
	wire [4-1:0] node4674;
	wire [4-1:0] node4675;
	wire [4-1:0] node4677;
	wire [4-1:0] node4679;
	wire [4-1:0] node4682;
	wire [4-1:0] node4684;
	wire [4-1:0] node4686;
	wire [4-1:0] node4689;
	wire [4-1:0] node4690;
	wire [4-1:0] node4691;
	wire [4-1:0] node4692;
	wire [4-1:0] node4693;
	wire [4-1:0] node4696;
	wire [4-1:0] node4698;
	wire [4-1:0] node4701;
	wire [4-1:0] node4702;
	wire [4-1:0] node4704;
	wire [4-1:0] node4707;
	wire [4-1:0] node4710;
	wire [4-1:0] node4711;
	wire [4-1:0] node4712;
	wire [4-1:0] node4714;
	wire [4-1:0] node4717;
	wire [4-1:0] node4719;
	wire [4-1:0] node4722;
	wire [4-1:0] node4723;
	wire [4-1:0] node4725;
	wire [4-1:0] node4728;
	wire [4-1:0] node4730;
	wire [4-1:0] node4733;
	wire [4-1:0] node4734;
	wire [4-1:0] node4735;
	wire [4-1:0] node4736;
	wire [4-1:0] node4740;
	wire [4-1:0] node4741;
	wire [4-1:0] node4744;
	wire [4-1:0] node4746;
	wire [4-1:0] node4749;
	wire [4-1:0] node4750;
	wire [4-1:0] node4752;
	wire [4-1:0] node4754;
	wire [4-1:0] node4757;
	wire [4-1:0] node4759;
	wire [4-1:0] node4761;
	wire [4-1:0] node4764;
	wire [4-1:0] node4765;
	wire [4-1:0] node4766;
	wire [4-1:0] node4767;
	wire [4-1:0] node4768;
	wire [4-1:0] node4769;
	wire [4-1:0] node4770;
	wire [4-1:0] node4773;
	wire [4-1:0] node4775;
	wire [4-1:0] node4778;
	wire [4-1:0] node4779;
	wire [4-1:0] node4781;
	wire [4-1:0] node4785;
	wire [4-1:0] node4786;
	wire [4-1:0] node4787;
	wire [4-1:0] node4791;
	wire [4-1:0] node4792;
	wire [4-1:0] node4793;
	wire [4-1:0] node4796;
	wire [4-1:0] node4799;
	wire [4-1:0] node4801;
	wire [4-1:0] node4804;
	wire [4-1:0] node4805;
	wire [4-1:0] node4806;
	wire [4-1:0] node4808;
	wire [4-1:0] node4811;
	wire [4-1:0] node4812;
	wire [4-1:0] node4813;
	wire [4-1:0] node4817;
	wire [4-1:0] node4818;
	wire [4-1:0] node4822;
	wire [4-1:0] node4823;
	wire [4-1:0] node4824;
	wire [4-1:0] node4827;
	wire [4-1:0] node4830;
	wire [4-1:0] node4833;
	wire [4-1:0] node4834;
	wire [4-1:0] node4835;
	wire [4-1:0] node4836;
	wire [4-1:0] node4839;
	wire [4-1:0] node4842;
	wire [4-1:0] node4843;
	wire [4-1:0] node4844;
	wire [4-1:0] node4846;
	wire [4-1:0] node4849;
	wire [4-1:0] node4850;
	wire [4-1:0] node4854;
	wire [4-1:0] node4855;
	wire [4-1:0] node4858;
	wire [4-1:0] node4861;
	wire [4-1:0] node4862;
	wire [4-1:0] node4863;
	wire [4-1:0] node4865;
	wire [4-1:0] node4868;
	wire [4-1:0] node4869;
	wire [4-1:0] node4870;
	wire [4-1:0] node4873;
	wire [4-1:0] node4877;
	wire [4-1:0] node4878;
	wire [4-1:0] node4880;
	wire [4-1:0] node4883;
	wire [4-1:0] node4885;
	wire [4-1:0] node4888;
	wire [4-1:0] node4889;
	wire [4-1:0] node4890;
	wire [4-1:0] node4891;
	wire [4-1:0] node4892;
	wire [4-1:0] node4894;
	wire [4-1:0] node4897;
	wire [4-1:0] node4899;
	wire [4-1:0] node4902;
	wire [4-1:0] node4903;
	wire [4-1:0] node4905;
	wire [4-1:0] node4908;
	wire [4-1:0] node4910;
	wire [4-1:0] node4913;
	wire [4-1:0] node4914;
	wire [4-1:0] node4915;
	wire [4-1:0] node4917;
	wire [4-1:0] node4920;
	wire [4-1:0] node4921;
	wire [4-1:0] node4924;
	wire [4-1:0] node4926;
	wire [4-1:0] node4929;
	wire [4-1:0] node4930;
	wire [4-1:0] node4931;
	wire [4-1:0] node4932;
	wire [4-1:0] node4935;
	wire [4-1:0] node4938;
	wire [4-1:0] node4939;
	wire [4-1:0] node4943;
	wire [4-1:0] node4944;
	wire [4-1:0] node4947;
	wire [4-1:0] node4950;
	wire [4-1:0] node4951;
	wire [4-1:0] node4952;
	wire [4-1:0] node4953;
	wire [4-1:0] node4954;
	wire [4-1:0] node4958;
	wire [4-1:0] node4959;
	wire [4-1:0] node4963;
	wire [4-1:0] node4964;
	wire [4-1:0] node4967;
	wire [4-1:0] node4968;
	wire [4-1:0] node4972;
	wire [4-1:0] node4973;
	wire [4-1:0] node4974;
	wire [4-1:0] node4977;
	wire [4-1:0] node4978;
	wire [4-1:0] node4979;
	wire [4-1:0] node4982;
	wire [4-1:0] node4985;
	wire [4-1:0] node4986;
	wire [4-1:0] node4990;
	wire [4-1:0] node4991;
	wire [4-1:0] node4993;
	wire [4-1:0] node4996;
	wire [4-1:0] node4998;
	wire [4-1:0] node5001;
	wire [4-1:0] node5002;
	wire [4-1:0] node5003;
	wire [4-1:0] node5004;
	wire [4-1:0] node5005;
	wire [4-1:0] node5006;
	wire [4-1:0] node5007;
	wire [4-1:0] node5010;
	wire [4-1:0] node5012;
	wire [4-1:0] node5015;
	wire [4-1:0] node5017;
	wire [4-1:0] node5019;
	wire [4-1:0] node5022;
	wire [4-1:0] node5023;
	wire [4-1:0] node5025;
	wire [4-1:0] node5028;
	wire [4-1:0] node5029;
	wire [4-1:0] node5031;
	wire [4-1:0] node5034;
	wire [4-1:0] node5036;
	wire [4-1:0] node5039;
	wire [4-1:0] node5040;
	wire [4-1:0] node5041;
	wire [4-1:0] node5042;
	wire [4-1:0] node5043;
	wire [4-1:0] node5045;
	wire [4-1:0] node5048;
	wire [4-1:0] node5049;
	wire [4-1:0] node5052;
	wire [4-1:0] node5055;
	wire [4-1:0] node5056;
	wire [4-1:0] node5059;
	wire [4-1:0] node5062;
	wire [4-1:0] node5063;
	wire [4-1:0] node5064;
	wire [4-1:0] node5067;
	wire [4-1:0] node5070;
	wire [4-1:0] node5071;
	wire [4-1:0] node5074;
	wire [4-1:0] node5075;
	wire [4-1:0] node5079;
	wire [4-1:0] node5080;
	wire [4-1:0] node5082;
	wire [4-1:0] node5083;
	wire [4-1:0] node5086;
	wire [4-1:0] node5089;
	wire [4-1:0] node5090;
	wire [4-1:0] node5092;
	wire [4-1:0] node5093;
	wire [4-1:0] node5096;
	wire [4-1:0] node5099;
	wire [4-1:0] node5101;
	wire [4-1:0] node5102;
	wire [4-1:0] node5105;
	wire [4-1:0] node5108;
	wire [4-1:0] node5109;
	wire [4-1:0] node5110;
	wire [4-1:0] node5111;
	wire [4-1:0] node5112;
	wire [4-1:0] node5113;
	wire [4-1:0] node5114;
	wire [4-1:0] node5117;
	wire [4-1:0] node5120;
	wire [4-1:0] node5122;
	wire [4-1:0] node5125;
	wire [4-1:0] node5126;
	wire [4-1:0] node5130;
	wire [4-1:0] node5131;
	wire [4-1:0] node5132;
	wire [4-1:0] node5133;
	wire [4-1:0] node5136;
	wire [4-1:0] node5139;
	wire [4-1:0] node5141;
	wire [4-1:0] node5144;
	wire [4-1:0] node5145;
	wire [4-1:0] node5147;
	wire [4-1:0] node5151;
	wire [4-1:0] node5152;
	wire [4-1:0] node5153;
	wire [4-1:0] node5154;
	wire [4-1:0] node5155;
	wire [4-1:0] node5158;
	wire [4-1:0] node5161;
	wire [4-1:0] node5162;
	wire [4-1:0] node5166;
	wire [4-1:0] node5167;
	wire [4-1:0] node5170;
	wire [4-1:0] node5173;
	wire [4-1:0] node5174;
	wire [4-1:0] node5175;
	wire [4-1:0] node5176;
	wire [4-1:0] node5180;
	wire [4-1:0] node5182;
	wire [4-1:0] node5185;
	wire [4-1:0] node5186;
	wire [4-1:0] node5189;
	wire [4-1:0] node5192;
	wire [4-1:0] node5193;
	wire [4-1:0] node5194;
	wire [4-1:0] node5195;
	wire [4-1:0] node5196;
	wire [4-1:0] node5197;
	wire [4-1:0] node5201;
	wire [4-1:0] node5203;
	wire [4-1:0] node5206;
	wire [4-1:0] node5207;
	wire [4-1:0] node5211;
	wire [4-1:0] node5212;
	wire [4-1:0] node5213;
	wire [4-1:0] node5216;
	wire [4-1:0] node5219;
	wire [4-1:0] node5220;
	wire [4-1:0] node5223;
	wire [4-1:0] node5226;
	wire [4-1:0] node5227;
	wire [4-1:0] node5228;
	wire [4-1:0] node5229;
	wire [4-1:0] node5232;
	wire [4-1:0] node5235;
	wire [4-1:0] node5236;
	wire [4-1:0] node5240;
	wire [4-1:0] node5241;
	wire [4-1:0] node5242;
	wire [4-1:0] node5245;
	wire [4-1:0] node5248;
	wire [4-1:0] node5250;
	wire [4-1:0] node5253;
	wire [4-1:0] node5254;
	wire [4-1:0] node5255;
	wire [4-1:0] node5256;
	wire [4-1:0] node5257;
	wire [4-1:0] node5258;
	wire [4-1:0] node5259;
	wire [4-1:0] node5262;
	wire [4-1:0] node5265;
	wire [4-1:0] node5266;
	wire [4-1:0] node5269;
	wire [4-1:0] node5272;
	wire [4-1:0] node5273;
	wire [4-1:0] node5274;
	wire [4-1:0] node5277;
	wire [4-1:0] node5280;
	wire [4-1:0] node5281;
	wire [4-1:0] node5283;
	wire [4-1:0] node5287;
	wire [4-1:0] node5288;
	wire [4-1:0] node5290;
	wire [4-1:0] node5291;
	wire [4-1:0] node5294;
	wire [4-1:0] node5297;
	wire [4-1:0] node5298;
	wire [4-1:0] node5299;
	wire [4-1:0] node5302;
	wire [4-1:0] node5305;
	wire [4-1:0] node5306;
	wire [4-1:0] node5310;
	wire [4-1:0] node5311;
	wire [4-1:0] node5312;
	wire [4-1:0] node5313;
	wire [4-1:0] node5314;
	wire [4-1:0] node5317;
	wire [4-1:0] node5320;
	wire [4-1:0] node5322;
	wire [4-1:0] node5325;
	wire [4-1:0] node5326;
	wire [4-1:0] node5327;
	wire [4-1:0] node5328;
	wire [4-1:0] node5331;
	wire [4-1:0] node5334;
	wire [4-1:0] node5336;
	wire [4-1:0] node5339;
	wire [4-1:0] node5340;
	wire [4-1:0] node5344;
	wire [4-1:0] node5345;
	wire [4-1:0] node5346;
	wire [4-1:0] node5347;
	wire [4-1:0] node5350;
	wire [4-1:0] node5353;
	wire [4-1:0] node5355;
	wire [4-1:0] node5357;
	wire [4-1:0] node5360;
	wire [4-1:0] node5361;
	wire [4-1:0] node5362;
	wire [4-1:0] node5363;
	wire [4-1:0] node5367;
	wire [4-1:0] node5368;
	wire [4-1:0] node5371;
	wire [4-1:0] node5374;
	wire [4-1:0] node5376;
	wire [4-1:0] node5377;
	wire [4-1:0] node5380;
	wire [4-1:0] node5383;
	wire [4-1:0] node5384;
	wire [4-1:0] node5385;
	wire [4-1:0] node5386;
	wire [4-1:0] node5387;
	wire [4-1:0] node5390;
	wire [4-1:0] node5392;
	wire [4-1:0] node5395;
	wire [4-1:0] node5396;
	wire [4-1:0] node5397;
	wire [4-1:0] node5400;
	wire [4-1:0] node5403;
	wire [4-1:0] node5404;
	wire [4-1:0] node5405;
	wire [4-1:0] node5408;
	wire [4-1:0] node5411;
	wire [4-1:0] node5413;
	wire [4-1:0] node5416;
	wire [4-1:0] node5417;
	wire [4-1:0] node5418;
	wire [4-1:0] node5419;
	wire [4-1:0] node5422;
	wire [4-1:0] node5425;
	wire [4-1:0] node5426;
	wire [4-1:0] node5428;
	wire [4-1:0] node5431;
	wire [4-1:0] node5432;
	wire [4-1:0] node5436;
	wire [4-1:0] node5437;
	wire [4-1:0] node5438;
	wire [4-1:0] node5441;
	wire [4-1:0] node5444;
	wire [4-1:0] node5445;
	wire [4-1:0] node5448;
	wire [4-1:0] node5451;
	wire [4-1:0] node5452;
	wire [4-1:0] node5453;
	wire [4-1:0] node5454;
	wire [4-1:0] node5455;
	wire [4-1:0] node5456;
	wire [4-1:0] node5459;
	wire [4-1:0] node5462;
	wire [4-1:0] node5463;
	wire [4-1:0] node5467;
	wire [4-1:0] node5468;
	wire [4-1:0] node5471;
	wire [4-1:0] node5474;
	wire [4-1:0] node5475;
	wire [4-1:0] node5478;
	wire [4-1:0] node5481;
	wire [4-1:0] node5482;
	wire [4-1:0] node5483;
	wire [4-1:0] node5484;
	wire [4-1:0] node5487;
	wire [4-1:0] node5490;
	wire [4-1:0] node5491;
	wire [4-1:0] node5495;
	wire [4-1:0] node5496;
	wire [4-1:0] node5497;
	wire [4-1:0] node5501;
	wire [4-1:0] node5504;
	wire [4-1:0] node5505;
	wire [4-1:0] node5506;
	wire [4-1:0] node5507;
	wire [4-1:0] node5508;
	wire [4-1:0] node5509;
	wire [4-1:0] node5510;
	wire [4-1:0] node5511;
	wire [4-1:0] node5512;
	wire [4-1:0] node5515;
	wire [4-1:0] node5518;
	wire [4-1:0] node5519;
	wire [4-1:0] node5522;
	wire [4-1:0] node5525;
	wire [4-1:0] node5526;
	wire [4-1:0] node5527;
	wire [4-1:0] node5529;
	wire [4-1:0] node5532;
	wire [4-1:0] node5534;
	wire [4-1:0] node5537;
	wire [4-1:0] node5538;
	wire [4-1:0] node5539;
	wire [4-1:0] node5544;
	wire [4-1:0] node5545;
	wire [4-1:0] node5546;
	wire [4-1:0] node5547;
	wire [4-1:0] node5551;
	wire [4-1:0] node5552;
	wire [4-1:0] node5556;
	wire [4-1:0] node5557;
	wire [4-1:0] node5558;
	wire [4-1:0] node5561;
	wire [4-1:0] node5564;
	wire [4-1:0] node5565;
	wire [4-1:0] node5566;
	wire [4-1:0] node5569;
	wire [4-1:0] node5572;
	wire [4-1:0] node5573;
	wire [4-1:0] node5576;
	wire [4-1:0] node5579;
	wire [4-1:0] node5580;
	wire [4-1:0] node5581;
	wire [4-1:0] node5582;
	wire [4-1:0] node5584;
	wire [4-1:0] node5587;
	wire [4-1:0] node5589;
	wire [4-1:0] node5592;
	wire [4-1:0] node5593;
	wire [4-1:0] node5595;
	wire [4-1:0] node5598;
	wire [4-1:0] node5600;
	wire [4-1:0] node5603;
	wire [4-1:0] node5604;
	wire [4-1:0] node5605;
	wire [4-1:0] node5607;
	wire [4-1:0] node5608;
	wire [4-1:0] node5611;
	wire [4-1:0] node5614;
	wire [4-1:0] node5615;
	wire [4-1:0] node5618;
	wire [4-1:0] node5621;
	wire [4-1:0] node5622;
	wire [4-1:0] node5623;
	wire [4-1:0] node5624;
	wire [4-1:0] node5629;
	wire [4-1:0] node5632;
	wire [4-1:0] node5633;
	wire [4-1:0] node5634;
	wire [4-1:0] node5635;
	wire [4-1:0] node5636;
	wire [4-1:0] node5637;
	wire [4-1:0] node5640;
	wire [4-1:0] node5643;
	wire [4-1:0] node5644;
	wire [4-1:0] node5647;
	wire [4-1:0] node5650;
	wire [4-1:0] node5652;
	wire [4-1:0] node5653;
	wire [4-1:0] node5654;
	wire [4-1:0] node5657;
	wire [4-1:0] node5660;
	wire [4-1:0] node5661;
	wire [4-1:0] node5665;
	wire [4-1:0] node5666;
	wire [4-1:0] node5667;
	wire [4-1:0] node5668;
	wire [4-1:0] node5671;
	wire [4-1:0] node5674;
	wire [4-1:0] node5676;
	wire [4-1:0] node5677;
	wire [4-1:0] node5681;
	wire [4-1:0] node5682;
	wire [4-1:0] node5683;
	wire [4-1:0] node5684;
	wire [4-1:0] node5687;
	wire [4-1:0] node5691;
	wire [4-1:0] node5692;
	wire [4-1:0] node5695;
	wire [4-1:0] node5698;
	wire [4-1:0] node5699;
	wire [4-1:0] node5700;
	wire [4-1:0] node5701;
	wire [4-1:0] node5702;
	wire [4-1:0] node5706;
	wire [4-1:0] node5707;
	wire [4-1:0] node5711;
	wire [4-1:0] node5712;
	wire [4-1:0] node5713;
	wire [4-1:0] node5717;
	wire [4-1:0] node5718;
	wire [4-1:0] node5722;
	wire [4-1:0] node5723;
	wire [4-1:0] node5724;
	wire [4-1:0] node5725;
	wire [4-1:0] node5726;
	wire [4-1:0] node5730;
	wire [4-1:0] node5731;
	wire [4-1:0] node5735;
	wire [4-1:0] node5736;
	wire [4-1:0] node5737;
	wire [4-1:0] node5742;
	wire [4-1:0] node5743;
	wire [4-1:0] node5745;
	wire [4-1:0] node5748;
	wire [4-1:0] node5750;
	wire [4-1:0] node5753;
	wire [4-1:0] node5754;
	wire [4-1:0] node5755;
	wire [4-1:0] node5756;
	wire [4-1:0] node5757;
	wire [4-1:0] node5758;
	wire [4-1:0] node5761;
	wire [4-1:0] node5764;
	wire [4-1:0] node5765;
	wire [4-1:0] node5768;
	wire [4-1:0] node5771;
	wire [4-1:0] node5772;
	wire [4-1:0] node5773;
	wire [4-1:0] node5775;
	wire [4-1:0] node5778;
	wire [4-1:0] node5779;
	wire [4-1:0] node5782;
	wire [4-1:0] node5785;
	wire [4-1:0] node5786;
	wire [4-1:0] node5787;
	wire [4-1:0] node5788;
	wire [4-1:0] node5791;
	wire [4-1:0] node5794;
	wire [4-1:0] node5795;
	wire [4-1:0] node5798;
	wire [4-1:0] node5801;
	wire [4-1:0] node5802;
	wire [4-1:0] node5805;
	wire [4-1:0] node5808;
	wire [4-1:0] node5809;
	wire [4-1:0] node5810;
	wire [4-1:0] node5811;
	wire [4-1:0] node5812;
	wire [4-1:0] node5815;
	wire [4-1:0] node5818;
	wire [4-1:0] node5819;
	wire [4-1:0] node5822;
	wire [4-1:0] node5825;
	wire [4-1:0] node5826;
	wire [4-1:0] node5827;
	wire [4-1:0] node5830;
	wire [4-1:0] node5833;
	wire [4-1:0] node5834;
	wire [4-1:0] node5835;
	wire [4-1:0] node5838;
	wire [4-1:0] node5842;
	wire [4-1:0] node5843;
	wire [4-1:0] node5844;
	wire [4-1:0] node5845;
	wire [4-1:0] node5846;
	wire [4-1:0] node5849;
	wire [4-1:0] node5852;
	wire [4-1:0] node5853;
	wire [4-1:0] node5857;
	wire [4-1:0] node5860;
	wire [4-1:0] node5861;
	wire [4-1:0] node5862;
	wire [4-1:0] node5864;
	wire [4-1:0] node5867;
	wire [4-1:0] node5868;
	wire [4-1:0] node5871;
	wire [4-1:0] node5874;
	wire [4-1:0] node5875;
	wire [4-1:0] node5878;
	wire [4-1:0] node5881;
	wire [4-1:0] node5882;
	wire [4-1:0] node5883;
	wire [4-1:0] node5884;
	wire [4-1:0] node5885;
	wire [4-1:0] node5886;
	wire [4-1:0] node5890;
	wire [4-1:0] node5892;
	wire [4-1:0] node5893;
	wire [4-1:0] node5897;
	wire [4-1:0] node5898;
	wire [4-1:0] node5899;
	wire [4-1:0] node5903;
	wire [4-1:0] node5904;
	wire [4-1:0] node5905;
	wire [4-1:0] node5909;
	wire [4-1:0] node5911;
	wire [4-1:0] node5914;
	wire [4-1:0] node5915;
	wire [4-1:0] node5916;
	wire [4-1:0] node5917;
	wire [4-1:0] node5920;
	wire [4-1:0] node5923;
	wire [4-1:0] node5924;
	wire [4-1:0] node5926;
	wire [4-1:0] node5929;
	wire [4-1:0] node5930;
	wire [4-1:0] node5934;
	wire [4-1:0] node5935;
	wire [4-1:0] node5936;
	wire [4-1:0] node5939;
	wire [4-1:0] node5942;
	wire [4-1:0] node5944;
	wire [4-1:0] node5947;
	wire [4-1:0] node5948;
	wire [4-1:0] node5949;
	wire [4-1:0] node5950;
	wire [4-1:0] node5952;
	wire [4-1:0] node5955;
	wire [4-1:0] node5956;
	wire [4-1:0] node5958;
	wire [4-1:0] node5961;
	wire [4-1:0] node5962;
	wire [4-1:0] node5965;
	wire [4-1:0] node5968;
	wire [4-1:0] node5969;
	wire [4-1:0] node5970;
	wire [4-1:0] node5971;
	wire [4-1:0] node5974;
	wire [4-1:0] node5977;
	wire [4-1:0] node5978;
	wire [4-1:0] node5981;
	wire [4-1:0] node5984;
	wire [4-1:0] node5985;
	wire [4-1:0] node5986;
	wire [4-1:0] node5989;
	wire [4-1:0] node5992;
	wire [4-1:0] node5993;
	wire [4-1:0] node5996;
	wire [4-1:0] node5999;
	wire [4-1:0] node6000;
	wire [4-1:0] node6001;
	wire [4-1:0] node6002;
	wire [4-1:0] node6005;
	wire [4-1:0] node6008;
	wire [4-1:0] node6009;
	wire [4-1:0] node6010;
	wire [4-1:0] node6014;
	wire [4-1:0] node6015;
	wire [4-1:0] node6018;
	wire [4-1:0] node6021;
	wire [4-1:0] node6022;
	wire [4-1:0] node6023;
	wire [4-1:0] node6026;
	wire [4-1:0] node6029;
	wire [4-1:0] node6030;
	wire [4-1:0] node6032;
	wire [4-1:0] node6035;
	wire [4-1:0] node6038;
	wire [4-1:0] node6039;
	wire [4-1:0] node6040;
	wire [4-1:0] node6041;
	wire [4-1:0] node6042;
	wire [4-1:0] node6043;
	wire [4-1:0] node6044;
	wire [4-1:0] node6045;
	wire [4-1:0] node6047;
	wire [4-1:0] node6050;
	wire [4-1:0] node6051;
	wire [4-1:0] node6054;
	wire [4-1:0] node6057;
	wire [4-1:0] node6058;
	wire [4-1:0] node6062;
	wire [4-1:0] node6063;
	wire [4-1:0] node6064;
	wire [4-1:0] node6068;
	wire [4-1:0] node6070;
	wire [4-1:0] node6071;
	wire [4-1:0] node6074;
	wire [4-1:0] node6077;
	wire [4-1:0] node6078;
	wire [4-1:0] node6079;
	wire [4-1:0] node6081;
	wire [4-1:0] node6084;
	wire [4-1:0] node6086;
	wire [4-1:0] node6089;
	wire [4-1:0] node6090;
	wire [4-1:0] node6092;
	wire [4-1:0] node6095;
	wire [4-1:0] node6097;
	wire [4-1:0] node6100;
	wire [4-1:0] node6101;
	wire [4-1:0] node6102;
	wire [4-1:0] node6103;
	wire [4-1:0] node6105;
	wire [4-1:0] node6108;
	wire [4-1:0] node6110;
	wire [4-1:0] node6113;
	wire [4-1:0] node6114;
	wire [4-1:0] node6116;
	wire [4-1:0] node6119;
	wire [4-1:0] node6121;
	wire [4-1:0] node6124;
	wire [4-1:0] node6125;
	wire [4-1:0] node6126;
	wire [4-1:0] node6128;
	wire [4-1:0] node6130;
	wire [4-1:0] node6133;
	wire [4-1:0] node6136;
	wire [4-1:0] node6137;
	wire [4-1:0] node6139;
	wire [4-1:0] node6142;
	wire [4-1:0] node6144;
	wire [4-1:0] node6147;
	wire [4-1:0] node6148;
	wire [4-1:0] node6149;
	wire [4-1:0] node6150;
	wire [4-1:0] node6151;
	wire [4-1:0] node6153;
	wire [4-1:0] node6156;
	wire [4-1:0] node6157;
	wire [4-1:0] node6160;
	wire [4-1:0] node6163;
	wire [4-1:0] node6164;
	wire [4-1:0] node6166;
	wire [4-1:0] node6169;
	wire [4-1:0] node6170;
	wire [4-1:0] node6171;
	wire [4-1:0] node6174;
	wire [4-1:0] node6177;
	wire [4-1:0] node6178;
	wire [4-1:0] node6181;
	wire [4-1:0] node6184;
	wire [4-1:0] node6185;
	wire [4-1:0] node6186;
	wire [4-1:0] node6188;
	wire [4-1:0] node6191;
	wire [4-1:0] node6193;
	wire [4-1:0] node6196;
	wire [4-1:0] node6197;
	wire [4-1:0] node6199;
	wire [4-1:0] node6202;
	wire [4-1:0] node6204;
	wire [4-1:0] node6207;
	wire [4-1:0] node6208;
	wire [4-1:0] node6209;
	wire [4-1:0] node6210;
	wire [4-1:0] node6212;
	wire [4-1:0] node6215;
	wire [4-1:0] node6216;
	wire [4-1:0] node6218;
	wire [4-1:0] node6222;
	wire [4-1:0] node6223;
	wire [4-1:0] node6225;
	wire [4-1:0] node6228;
	wire [4-1:0] node6230;
	wire [4-1:0] node6233;
	wire [4-1:0] node6234;
	wire [4-1:0] node6235;
	wire [4-1:0] node6238;
	wire [4-1:0] node6241;
	wire [4-1:0] node6242;
	wire [4-1:0] node6243;
	wire [4-1:0] node6246;
	wire [4-1:0] node6250;
	wire [4-1:0] node6251;
	wire [4-1:0] node6252;
	wire [4-1:0] node6253;
	wire [4-1:0] node6254;
	wire [4-1:0] node6255;
	wire [4-1:0] node6258;
	wire [4-1:0] node6261;
	wire [4-1:0] node6262;
	wire [4-1:0] node6263;
	wire [4-1:0] node6266;
	wire [4-1:0] node6269;
	wire [4-1:0] node6270;
	wire [4-1:0] node6271;
	wire [4-1:0] node6275;
	wire [4-1:0] node6277;
	wire [4-1:0] node6280;
	wire [4-1:0] node6281;
	wire [4-1:0] node6282;
	wire [4-1:0] node6285;
	wire [4-1:0] node6287;
	wire [4-1:0] node6290;
	wire [4-1:0] node6291;
	wire [4-1:0] node6293;
	wire [4-1:0] node6296;
	wire [4-1:0] node6298;
	wire [4-1:0] node6301;
	wire [4-1:0] node6302;
	wire [4-1:0] node6303;
	wire [4-1:0] node6304;
	wire [4-1:0] node6306;
	wire [4-1:0] node6309;
	wire [4-1:0] node6311;
	wire [4-1:0] node6314;
	wire [4-1:0] node6315;
	wire [4-1:0] node6316;
	wire [4-1:0] node6319;
	wire [4-1:0] node6322;
	wire [4-1:0] node6324;
	wire [4-1:0] node6326;
	wire [4-1:0] node6329;
	wire [4-1:0] node6330;
	wire [4-1:0] node6331;
	wire [4-1:0] node6332;
	wire [4-1:0] node6335;
	wire [4-1:0] node6338;
	wire [4-1:0] node6339;
	wire [4-1:0] node6340;
	wire [4-1:0] node6343;
	wire [4-1:0] node6346;
	wire [4-1:0] node6347;
	wire [4-1:0] node6350;
	wire [4-1:0] node6353;
	wire [4-1:0] node6354;
	wire [4-1:0] node6355;
	wire [4-1:0] node6358;
	wire [4-1:0] node6360;
	wire [4-1:0] node6363;
	wire [4-1:0] node6365;
	wire [4-1:0] node6366;
	wire [4-1:0] node6369;
	wire [4-1:0] node6372;
	wire [4-1:0] node6373;
	wire [4-1:0] node6374;
	wire [4-1:0] node6375;
	wire [4-1:0] node6376;
	wire [4-1:0] node6379;
	wire [4-1:0] node6382;
	wire [4-1:0] node6383;
	wire [4-1:0] node6384;
	wire [4-1:0] node6385;
	wire [4-1:0] node6388;
	wire [4-1:0] node6392;
	wire [4-1:0] node6393;
	wire [4-1:0] node6397;
	wire [4-1:0] node6398;
	wire [4-1:0] node6399;
	wire [4-1:0] node6401;
	wire [4-1:0] node6404;
	wire [4-1:0] node6406;
	wire [4-1:0] node6409;
	wire [4-1:0] node6410;
	wire [4-1:0] node6412;
	wire [4-1:0] node6415;
	wire [4-1:0] node6416;
	wire [4-1:0] node6418;
	wire [4-1:0] node6422;
	wire [4-1:0] node6423;
	wire [4-1:0] node6424;
	wire [4-1:0] node6425;
	wire [4-1:0] node6427;
	wire [4-1:0] node6430;
	wire [4-1:0] node6432;
	wire [4-1:0] node6435;
	wire [4-1:0] node6437;
	wire [4-1:0] node6439;
	wire [4-1:0] node6442;
	wire [4-1:0] node6443;
	wire [4-1:0] node6444;
	wire [4-1:0] node6445;
	wire [4-1:0] node6448;
	wire [4-1:0] node6451;
	wire [4-1:0] node6452;
	wire [4-1:0] node6455;
	wire [4-1:0] node6456;
	wire [4-1:0] node6460;
	wire [4-1:0] node6461;
	wire [4-1:0] node6462;
	wire [4-1:0] node6466;
	wire [4-1:0] node6467;
	wire [4-1:0] node6468;
	wire [4-1:0] node6471;
	wire [4-1:0] node6474;
	wire [4-1:0] node6475;
	wire [4-1:0] node6478;
	wire [4-1:0] node6481;
	wire [4-1:0] node6482;
	wire [4-1:0] node6483;
	wire [4-1:0] node6484;
	wire [4-1:0] node6485;
	wire [4-1:0] node6486;
	wire [4-1:0] node6487;
	wire [4-1:0] node6488;
	wire [4-1:0] node6489;
	wire [4-1:0] node6492;
	wire [4-1:0] node6495;
	wire [4-1:0] node6496;
	wire [4-1:0] node6497;
	wire [4-1:0] node6500;
	wire [4-1:0] node6501;
	wire [4-1:0] node6505;
	wire [4-1:0] node6506;
	wire [4-1:0] node6509;
	wire [4-1:0] node6512;
	wire [4-1:0] node6513;
	wire [4-1:0] node6514;
	wire [4-1:0] node6515;
	wire [4-1:0] node6519;
	wire [4-1:0] node6520;
	wire [4-1:0] node6523;
	wire [4-1:0] node6524;
	wire [4-1:0] node6528;
	wire [4-1:0] node6529;
	wire [4-1:0] node6531;
	wire [4-1:0] node6534;
	wire [4-1:0] node6535;
	wire [4-1:0] node6536;
	wire [4-1:0] node6539;
	wire [4-1:0] node6542;
	wire [4-1:0] node6543;
	wire [4-1:0] node6546;
	wire [4-1:0] node6549;
	wire [4-1:0] node6550;
	wire [4-1:0] node6551;
	wire [4-1:0] node6552;
	wire [4-1:0] node6553;
	wire [4-1:0] node6556;
	wire [4-1:0] node6559;
	wire [4-1:0] node6560;
	wire [4-1:0] node6561;
	wire [4-1:0] node6564;
	wire [4-1:0] node6567;
	wire [4-1:0] node6568;
	wire [4-1:0] node6571;
	wire [4-1:0] node6574;
	wire [4-1:0] node6575;
	wire [4-1:0] node6576;
	wire [4-1:0] node6580;
	wire [4-1:0] node6581;
	wire [4-1:0] node6583;
	wire [4-1:0] node6586;
	wire [4-1:0] node6588;
	wire [4-1:0] node6591;
	wire [4-1:0] node6592;
	wire [4-1:0] node6593;
	wire [4-1:0] node6594;
	wire [4-1:0] node6597;
	wire [4-1:0] node6600;
	wire [4-1:0] node6601;
	wire [4-1:0] node6604;
	wire [4-1:0] node6607;
	wire [4-1:0] node6608;
	wire [4-1:0] node6611;
	wire [4-1:0] node6614;
	wire [4-1:0] node6615;
	wire [4-1:0] node6616;
	wire [4-1:0] node6617;
	wire [4-1:0] node6619;
	wire [4-1:0] node6620;
	wire [4-1:0] node6623;
	wire [4-1:0] node6626;
	wire [4-1:0] node6627;
	wire [4-1:0] node6628;
	wire [4-1:0] node6629;
	wire [4-1:0] node6632;
	wire [4-1:0] node6635;
	wire [4-1:0] node6636;
	wire [4-1:0] node6639;
	wire [4-1:0] node6642;
	wire [4-1:0] node6643;
	wire [4-1:0] node6644;
	wire [4-1:0] node6647;
	wire [4-1:0] node6650;
	wire [4-1:0] node6651;
	wire [4-1:0] node6654;
	wire [4-1:0] node6657;
	wire [4-1:0] node6658;
	wire [4-1:0] node6659;
	wire [4-1:0] node6660;
	wire [4-1:0] node6661;
	wire [4-1:0] node6665;
	wire [4-1:0] node6667;
	wire [4-1:0] node6670;
	wire [4-1:0] node6671;
	wire [4-1:0] node6675;
	wire [4-1:0] node6676;
	wire [4-1:0] node6677;
	wire [4-1:0] node6679;
	wire [4-1:0] node6682;
	wire [4-1:0] node6683;
	wire [4-1:0] node6687;
	wire [4-1:0] node6688;
	wire [4-1:0] node6690;
	wire [4-1:0] node6693;
	wire [4-1:0] node6694;
	wire [4-1:0] node6697;
	wire [4-1:0] node6700;
	wire [4-1:0] node6701;
	wire [4-1:0] node6702;
	wire [4-1:0] node6703;
	wire [4-1:0] node6704;
	wire [4-1:0] node6706;
	wire [4-1:0] node6709;
	wire [4-1:0] node6710;
	wire [4-1:0] node6713;
	wire [4-1:0] node6716;
	wire [4-1:0] node6717;
	wire [4-1:0] node6718;
	wire [4-1:0] node6721;
	wire [4-1:0] node6724;
	wire [4-1:0] node6726;
	wire [4-1:0] node6729;
	wire [4-1:0] node6730;
	wire [4-1:0] node6731;
	wire [4-1:0] node6734;
	wire [4-1:0] node6737;
	wire [4-1:0] node6739;
	wire [4-1:0] node6741;
	wire [4-1:0] node6744;
	wire [4-1:0] node6745;
	wire [4-1:0] node6746;
	wire [4-1:0] node6747;
	wire [4-1:0] node6749;
	wire [4-1:0] node6752;
	wire [4-1:0] node6753;
	wire [4-1:0] node6757;
	wire [4-1:0] node6758;
	wire [4-1:0] node6759;
	wire [4-1:0] node6762;
	wire [4-1:0] node6765;
	wire [4-1:0] node6766;
	wire [4-1:0] node6769;
	wire [4-1:0] node6772;
	wire [4-1:0] node6773;
	wire [4-1:0] node6774;
	wire [4-1:0] node6775;
	wire [4-1:0] node6778;
	wire [4-1:0] node6782;
	wire [4-1:0] node6783;
	wire [4-1:0] node6784;
	wire [4-1:0] node6788;
	wire [4-1:0] node6789;
	wire [4-1:0] node6793;
	wire [4-1:0] node6794;
	wire [4-1:0] node6795;
	wire [4-1:0] node6796;
	wire [4-1:0] node6797;
	wire [4-1:0] node6798;
	wire [4-1:0] node6801;
	wire [4-1:0] node6803;
	wire [4-1:0] node6806;
	wire [4-1:0] node6807;
	wire [4-1:0] node6809;
	wire [4-1:0] node6812;
	wire [4-1:0] node6814;
	wire [4-1:0] node6817;
	wire [4-1:0] node6818;
	wire [4-1:0] node6819;
	wire [4-1:0] node6820;
	wire [4-1:0] node6822;
	wire [4-1:0] node6825;
	wire [4-1:0] node6828;
	wire [4-1:0] node6830;
	wire [4-1:0] node6831;
	wire [4-1:0] node6834;
	wire [4-1:0] node6837;
	wire [4-1:0] node6838;
	wire [4-1:0] node6839;
	wire [4-1:0] node6842;
	wire [4-1:0] node6845;
	wire [4-1:0] node6846;
	wire [4-1:0] node6847;
	wire [4-1:0] node6851;
	wire [4-1:0] node6852;
	wire [4-1:0] node6855;
	wire [4-1:0] node6858;
	wire [4-1:0] node6859;
	wire [4-1:0] node6860;
	wire [4-1:0] node6861;
	wire [4-1:0] node6863;
	wire [4-1:0] node6866;
	wire [4-1:0] node6867;
	wire [4-1:0] node6870;
	wire [4-1:0] node6873;
	wire [4-1:0] node6874;
	wire [4-1:0] node6875;
	wire [4-1:0] node6876;
	wire [4-1:0] node6880;
	wire [4-1:0] node6881;
	wire [4-1:0] node6884;
	wire [4-1:0] node6887;
	wire [4-1:0] node6889;
	wire [4-1:0] node6890;
	wire [4-1:0] node6893;
	wire [4-1:0] node6896;
	wire [4-1:0] node6897;
	wire [4-1:0] node6898;
	wire [4-1:0] node6899;
	wire [4-1:0] node6903;
	wire [4-1:0] node6904;
	wire [4-1:0] node6907;
	wire [4-1:0] node6910;
	wire [4-1:0] node6911;
	wire [4-1:0] node6913;
	wire [4-1:0] node6914;
	wire [4-1:0] node6918;
	wire [4-1:0] node6919;
	wire [4-1:0] node6922;
	wire [4-1:0] node6925;
	wire [4-1:0] node6926;
	wire [4-1:0] node6927;
	wire [4-1:0] node6928;
	wire [4-1:0] node6929;
	wire [4-1:0] node6931;
	wire [4-1:0] node6934;
	wire [4-1:0] node6936;
	wire [4-1:0] node6939;
	wire [4-1:0] node6940;
	wire [4-1:0] node6942;
	wire [4-1:0] node6945;
	wire [4-1:0] node6948;
	wire [4-1:0] node6949;
	wire [4-1:0] node6950;
	wire [4-1:0] node6951;
	wire [4-1:0] node6954;
	wire [4-1:0] node6957;
	wire [4-1:0] node6959;
	wire [4-1:0] node6961;
	wire [4-1:0] node6964;
	wire [4-1:0] node6965;
	wire [4-1:0] node6966;
	wire [4-1:0] node6967;
	wire [4-1:0] node6970;
	wire [4-1:0] node6973;
	wire [4-1:0] node6974;
	wire [4-1:0] node6977;
	wire [4-1:0] node6980;
	wire [4-1:0] node6982;
	wire [4-1:0] node6985;
	wire [4-1:0] node6986;
	wire [4-1:0] node6987;
	wire [4-1:0] node6988;
	wire [4-1:0] node6989;
	wire [4-1:0] node6992;
	wire [4-1:0] node6995;
	wire [4-1:0] node6996;
	wire [4-1:0] node6998;
	wire [4-1:0] node7001;
	wire [4-1:0] node7003;
	wire [4-1:0] node7006;
	wire [4-1:0] node7007;
	wire [4-1:0] node7010;
	wire [4-1:0] node7013;
	wire [4-1:0] node7014;
	wire [4-1:0] node7015;
	wire [4-1:0] node7016;
	wire [4-1:0] node7019;
	wire [4-1:0] node7022;
	wire [4-1:0] node7025;
	wire [4-1:0] node7026;
	wire [4-1:0] node7027;
	wire [4-1:0] node7028;
	wire [4-1:0] node7031;
	wire [4-1:0] node7035;
	wire [4-1:0] node7036;
	wire [4-1:0] node7040;
	wire [4-1:0] node7041;
	wire [4-1:0] node7042;
	wire [4-1:0] node7043;
	wire [4-1:0] node7044;
	wire [4-1:0] node7045;
	wire [4-1:0] node7046;
	wire [4-1:0] node7048;
	wire [4-1:0] node7052;
	wire [4-1:0] node7053;
	wire [4-1:0] node7055;
	wire [4-1:0] node7059;
	wire [4-1:0] node7060;
	wire [4-1:0] node7061;
	wire [4-1:0] node7062;
	wire [4-1:0] node7064;
	wire [4-1:0] node7067;
	wire [4-1:0] node7069;
	wire [4-1:0] node7072;
	wire [4-1:0] node7073;
	wire [4-1:0] node7077;
	wire [4-1:0] node7078;
	wire [4-1:0] node7079;
	wire [4-1:0] node7083;
	wire [4-1:0] node7084;
	wire [4-1:0] node7087;
	wire [4-1:0] node7089;
	wire [4-1:0] node7092;
	wire [4-1:0] node7093;
	wire [4-1:0] node7094;
	wire [4-1:0] node7095;
	wire [4-1:0] node7097;
	wire [4-1:0] node7100;
	wire [4-1:0] node7102;
	wire [4-1:0] node7105;
	wire [4-1:0] node7106;
	wire [4-1:0] node7108;
	wire [4-1:0] node7111;
	wire [4-1:0] node7113;
	wire [4-1:0] node7116;
	wire [4-1:0] node7117;
	wire [4-1:0] node7118;
	wire [4-1:0] node7120;
	wire [4-1:0] node7123;
	wire [4-1:0] node7124;
	wire [4-1:0] node7125;
	wire [4-1:0] node7130;
	wire [4-1:0] node7131;
	wire [4-1:0] node7132;
	wire [4-1:0] node7135;
	wire [4-1:0] node7136;
	wire [4-1:0] node7140;
	wire [4-1:0] node7141;
	wire [4-1:0] node7142;
	wire [4-1:0] node7145;
	wire [4-1:0] node7149;
	wire [4-1:0] node7150;
	wire [4-1:0] node7151;
	wire [4-1:0] node7152;
	wire [4-1:0] node7153;
	wire [4-1:0] node7156;
	wire [4-1:0] node7159;
	wire [4-1:0] node7160;
	wire [4-1:0] node7162;
	wire [4-1:0] node7165;
	wire [4-1:0] node7166;
	wire [4-1:0] node7169;
	wire [4-1:0] node7172;
	wire [4-1:0] node7173;
	wire [4-1:0] node7174;
	wire [4-1:0] node7178;
	wire [4-1:0] node7179;
	wire [4-1:0] node7180;
	wire [4-1:0] node7183;
	wire [4-1:0] node7186;
	wire [4-1:0] node7187;
	wire [4-1:0] node7190;
	wire [4-1:0] node7193;
	wire [4-1:0] node7194;
	wire [4-1:0] node7195;
	wire [4-1:0] node7196;
	wire [4-1:0] node7199;
	wire [4-1:0] node7201;
	wire [4-1:0] node7204;
	wire [4-1:0] node7205;
	wire [4-1:0] node7206;
	wire [4-1:0] node7209;
	wire [4-1:0] node7212;
	wire [4-1:0] node7214;
	wire [4-1:0] node7217;
	wire [4-1:0] node7218;
	wire [4-1:0] node7219;
	wire [4-1:0] node7220;
	wire [4-1:0] node7223;
	wire [4-1:0] node7226;
	wire [4-1:0] node7227;
	wire [4-1:0] node7230;
	wire [4-1:0] node7233;
	wire [4-1:0] node7234;
	wire [4-1:0] node7235;
	wire [4-1:0] node7238;
	wire [4-1:0] node7241;
	wire [4-1:0] node7243;
	wire [4-1:0] node7245;
	wire [4-1:0] node7248;
	wire [4-1:0] node7249;
	wire [4-1:0] node7250;
	wire [4-1:0] node7251;
	wire [4-1:0] node7252;
	wire [4-1:0] node7253;
	wire [4-1:0] node7254;
	wire [4-1:0] node7257;
	wire [4-1:0] node7260;
	wire [4-1:0] node7261;
	wire [4-1:0] node7262;
	wire [4-1:0] node7266;
	wire [4-1:0] node7268;
	wire [4-1:0] node7271;
	wire [4-1:0] node7272;
	wire [4-1:0] node7273;
	wire [4-1:0] node7276;
	wire [4-1:0] node7279;
	wire [4-1:0] node7280;
	wire [4-1:0] node7282;
	wire [4-1:0] node7285;
	wire [4-1:0] node7287;
	wire [4-1:0] node7290;
	wire [4-1:0] node7291;
	wire [4-1:0] node7292;
	wire [4-1:0] node7294;
	wire [4-1:0] node7297;
	wire [4-1:0] node7298;
	wire [4-1:0] node7299;
	wire [4-1:0] node7303;
	wire [4-1:0] node7306;
	wire [4-1:0] node7307;
	wire [4-1:0] node7308;
	wire [4-1:0] node7309;
	wire [4-1:0] node7313;
	wire [4-1:0] node7314;
	wire [4-1:0] node7318;
	wire [4-1:0] node7319;
	wire [4-1:0] node7320;
	wire [4-1:0] node7323;
	wire [4-1:0] node7326;
	wire [4-1:0] node7327;
	wire [4-1:0] node7330;
	wire [4-1:0] node7333;
	wire [4-1:0] node7334;
	wire [4-1:0] node7335;
	wire [4-1:0] node7336;
	wire [4-1:0] node7337;
	wire [4-1:0] node7340;
	wire [4-1:0] node7342;
	wire [4-1:0] node7345;
	wire [4-1:0] node7346;
	wire [4-1:0] node7347;
	wire [4-1:0] node7350;
	wire [4-1:0] node7353;
	wire [4-1:0] node7354;
	wire [4-1:0] node7358;
	wire [4-1:0] node7359;
	wire [4-1:0] node7360;
	wire [4-1:0] node7363;
	wire [4-1:0] node7366;
	wire [4-1:0] node7367;
	wire [4-1:0] node7368;
	wire [4-1:0] node7371;
	wire [4-1:0] node7374;
	wire [4-1:0] node7375;
	wire [4-1:0] node7378;
	wire [4-1:0] node7381;
	wire [4-1:0] node7382;
	wire [4-1:0] node7383;
	wire [4-1:0] node7385;
	wire [4-1:0] node7386;
	wire [4-1:0] node7389;
	wire [4-1:0] node7392;
	wire [4-1:0] node7393;
	wire [4-1:0] node7394;
	wire [4-1:0] node7398;
	wire [4-1:0] node7399;
	wire [4-1:0] node7402;
	wire [4-1:0] node7405;
	wire [4-1:0] node7406;
	wire [4-1:0] node7409;
	wire [4-1:0] node7410;
	wire [4-1:0] node7412;
	wire [4-1:0] node7415;
	wire [4-1:0] node7416;
	wire [4-1:0] node7420;
	wire [4-1:0] node7421;
	wire [4-1:0] node7422;
	wire [4-1:0] node7423;
	wire [4-1:0] node7424;
	wire [4-1:0] node7425;
	wire [4-1:0] node7428;
	wire [4-1:0] node7431;
	wire [4-1:0] node7432;
	wire [4-1:0] node7433;
	wire [4-1:0] node7438;
	wire [4-1:0] node7439;
	wire [4-1:0] node7440;
	wire [4-1:0] node7441;
	wire [4-1:0] node7444;
	wire [4-1:0] node7447;
	wire [4-1:0] node7448;
	wire [4-1:0] node7451;
	wire [4-1:0] node7454;
	wire [4-1:0] node7455;
	wire [4-1:0] node7456;
	wire [4-1:0] node7459;
	wire [4-1:0] node7462;
	wire [4-1:0] node7463;
	wire [4-1:0] node7466;
	wire [4-1:0] node7469;
	wire [4-1:0] node7470;
	wire [4-1:0] node7471;
	wire [4-1:0] node7472;
	wire [4-1:0] node7473;
	wire [4-1:0] node7476;
	wire [4-1:0] node7479;
	wire [4-1:0] node7480;
	wire [4-1:0] node7483;
	wire [4-1:0] node7486;
	wire [4-1:0] node7487;
	wire [4-1:0] node7491;
	wire [4-1:0] node7492;
	wire [4-1:0] node7494;
	wire [4-1:0] node7497;
	wire [4-1:0] node7498;
	wire [4-1:0] node7499;
	wire [4-1:0] node7503;
	wire [4-1:0] node7505;
	wire [4-1:0] node7508;
	wire [4-1:0] node7509;
	wire [4-1:0] node7510;
	wire [4-1:0] node7511;
	wire [4-1:0] node7513;
	wire [4-1:0] node7514;
	wire [4-1:0] node7518;
	wire [4-1:0] node7519;
	wire [4-1:0] node7520;
	wire [4-1:0] node7524;
	wire [4-1:0] node7527;
	wire [4-1:0] node7528;
	wire [4-1:0] node7529;
	wire [4-1:0] node7530;
	wire [4-1:0] node7533;
	wire [4-1:0] node7536;
	wire [4-1:0] node7537;
	wire [4-1:0] node7540;
	wire [4-1:0] node7543;
	wire [4-1:0] node7545;
	wire [4-1:0] node7546;
	wire [4-1:0] node7549;
	wire [4-1:0] node7552;
	wire [4-1:0] node7553;
	wire [4-1:0] node7554;
	wire [4-1:0] node7555;
	wire [4-1:0] node7558;
	wire [4-1:0] node7559;
	wire [4-1:0] node7562;
	wire [4-1:0] node7565;
	wire [4-1:0] node7566;
	wire [4-1:0] node7567;
	wire [4-1:0] node7571;
	wire [4-1:0] node7574;
	wire [4-1:0] node7575;
	wire [4-1:0] node7576;
	wire [4-1:0] node7577;
	wire [4-1:0] node7580;
	wire [4-1:0] node7583;
	wire [4-1:0] node7586;
	wire [4-1:0] node7587;
	wire [4-1:0] node7588;
	wire [4-1:0] node7592;
	wire [4-1:0] node7595;
	wire [4-1:0] node7596;
	wire [4-1:0] node7597;
	wire [4-1:0] node7598;
	wire [4-1:0] node7599;
	wire [4-1:0] node7600;
	wire [4-1:0] node7601;
	wire [4-1:0] node7602;
	wire [4-1:0] node7603;
	wire [4-1:0] node7605;
	wire [4-1:0] node7608;
	wire [4-1:0] node7610;
	wire [4-1:0] node7613;
	wire [4-1:0] node7614;
	wire [4-1:0] node7616;
	wire [4-1:0] node7619;
	wire [4-1:0] node7621;
	wire [4-1:0] node7624;
	wire [4-1:0] node7625;
	wire [4-1:0] node7626;
	wire [4-1:0] node7628;
	wire [4-1:0] node7632;
	wire [4-1:0] node7633;
	wire [4-1:0] node7635;
	wire [4-1:0] node7638;
	wire [4-1:0] node7641;
	wire [4-1:0] node7642;
	wire [4-1:0] node7643;
	wire [4-1:0] node7644;
	wire [4-1:0] node7646;
	wire [4-1:0] node7650;
	wire [4-1:0] node7651;
	wire [4-1:0] node7653;
	wire [4-1:0] node7656;
	wire [4-1:0] node7659;
	wire [4-1:0] node7660;
	wire [4-1:0] node7662;
	wire [4-1:0] node7665;
	wire [4-1:0] node7666;
	wire [4-1:0] node7667;
	wire [4-1:0] node7670;
	wire [4-1:0] node7674;
	wire [4-1:0] node7675;
	wire [4-1:0] node7676;
	wire [4-1:0] node7677;
	wire [4-1:0] node7679;
	wire [4-1:0] node7682;
	wire [4-1:0] node7684;
	wire [4-1:0] node7686;
	wire [4-1:0] node7689;
	wire [4-1:0] node7691;
	wire [4-1:0] node7692;
	wire [4-1:0] node7694;
	wire [4-1:0] node7697;
	wire [4-1:0] node7700;
	wire [4-1:0] node7701;
	wire [4-1:0] node7702;
	wire [4-1:0] node7704;
	wire [4-1:0] node7705;
	wire [4-1:0] node7709;
	wire [4-1:0] node7710;
	wire [4-1:0] node7712;
	wire [4-1:0] node7716;
	wire [4-1:0] node7717;
	wire [4-1:0] node7719;
	wire [4-1:0] node7722;
	wire [4-1:0] node7723;
	wire [4-1:0] node7724;
	wire [4-1:0] node7727;
	wire [4-1:0] node7730;
	wire [4-1:0] node7731;
	wire [4-1:0] node7734;
	wire [4-1:0] node7737;
	wire [4-1:0] node7738;
	wire [4-1:0] node7739;
	wire [4-1:0] node7740;
	wire [4-1:0] node7741;
	wire [4-1:0] node7743;
	wire [4-1:0] node7744;
	wire [4-1:0] node7748;
	wire [4-1:0] node7749;
	wire [4-1:0] node7751;
	wire [4-1:0] node7754;
	wire [4-1:0] node7755;
	wire [4-1:0] node7759;
	wire [4-1:0] node7760;
	wire [4-1:0] node7761;
	wire [4-1:0] node7765;
	wire [4-1:0] node7766;
	wire [4-1:0] node7767;
	wire [4-1:0] node7771;
	wire [4-1:0] node7773;
	wire [4-1:0] node7776;
	wire [4-1:0] node7777;
	wire [4-1:0] node7778;
	wire [4-1:0] node7779;
	wire [4-1:0] node7780;
	wire [4-1:0] node7783;
	wire [4-1:0] node7787;
	wire [4-1:0] node7788;
	wire [4-1:0] node7789;
	wire [4-1:0] node7792;
	wire [4-1:0] node7795;
	wire [4-1:0] node7796;
	wire [4-1:0] node7799;
	wire [4-1:0] node7802;
	wire [4-1:0] node7803;
	wire [4-1:0] node7804;
	wire [4-1:0] node7807;
	wire [4-1:0] node7809;
	wire [4-1:0] node7812;
	wire [4-1:0] node7813;
	wire [4-1:0] node7815;
	wire [4-1:0] node7819;
	wire [4-1:0] node7820;
	wire [4-1:0] node7821;
	wire [4-1:0] node7822;
	wire [4-1:0] node7823;
	wire [4-1:0] node7827;
	wire [4-1:0] node7828;
	wire [4-1:0] node7831;
	wire [4-1:0] node7833;
	wire [4-1:0] node7836;
	wire [4-1:0] node7837;
	wire [4-1:0] node7839;
	wire [4-1:0] node7840;
	wire [4-1:0] node7843;
	wire [4-1:0] node7846;
	wire [4-1:0] node7847;
	wire [4-1:0] node7849;
	wire [4-1:0] node7852;
	wire [4-1:0] node7855;
	wire [4-1:0] node7856;
	wire [4-1:0] node7857;
	wire [4-1:0] node7858;
	wire [4-1:0] node7860;
	wire [4-1:0] node7863;
	wire [4-1:0] node7866;
	wire [4-1:0] node7867;
	wire [4-1:0] node7870;
	wire [4-1:0] node7873;
	wire [4-1:0] node7874;
	wire [4-1:0] node7875;
	wire [4-1:0] node7877;
	wire [4-1:0] node7880;
	wire [4-1:0] node7882;
	wire [4-1:0] node7885;
	wire [4-1:0] node7887;
	wire [4-1:0] node7889;
	wire [4-1:0] node7892;
	wire [4-1:0] node7893;
	wire [4-1:0] node7894;
	wire [4-1:0] node7895;
	wire [4-1:0] node7896;
	wire [4-1:0] node7897;
	wire [4-1:0] node7899;
	wire [4-1:0] node7902;
	wire [4-1:0] node7904;
	wire [4-1:0] node7907;
	wire [4-1:0] node7908;
	wire [4-1:0] node7911;
	wire [4-1:0] node7913;
	wire [4-1:0] node7916;
	wire [4-1:0] node7917;
	wire [4-1:0] node7918;
	wire [4-1:0] node7919;
	wire [4-1:0] node7923;
	wire [4-1:0] node7924;
	wire [4-1:0] node7928;
	wire [4-1:0] node7929;
	wire [4-1:0] node7931;
	wire [4-1:0] node7934;
	wire [4-1:0] node7935;
	wire [4-1:0] node7936;
	wire [4-1:0] node7940;
	wire [4-1:0] node7941;
	wire [4-1:0] node7944;
	wire [4-1:0] node7947;
	wire [4-1:0] node7948;
	wire [4-1:0] node7949;
	wire [4-1:0] node7950;
	wire [4-1:0] node7952;
	wire [4-1:0] node7955;
	wire [4-1:0] node7957;
	wire [4-1:0] node7960;
	wire [4-1:0] node7961;
	wire [4-1:0] node7963;
	wire [4-1:0] node7966;
	wire [4-1:0] node7968;
	wire [4-1:0] node7971;
	wire [4-1:0] node7972;
	wire [4-1:0] node7973;
	wire [4-1:0] node7974;
	wire [4-1:0] node7977;
	wire [4-1:0] node7980;
	wire [4-1:0] node7981;
	wire [4-1:0] node7983;
	wire [4-1:0] node7986;
	wire [4-1:0] node7987;
	wire [4-1:0] node7990;
	wire [4-1:0] node7993;
	wire [4-1:0] node7994;
	wire [4-1:0] node7995;
	wire [4-1:0] node7996;
	wire [4-1:0] node8000;
	wire [4-1:0] node8001;
	wire [4-1:0] node8005;
	wire [4-1:0] node8006;
	wire [4-1:0] node8010;
	wire [4-1:0] node8011;
	wire [4-1:0] node8012;
	wire [4-1:0] node8013;
	wire [4-1:0] node8014;
	wire [4-1:0] node8017;
	wire [4-1:0] node8020;
	wire [4-1:0] node8021;
	wire [4-1:0] node8022;
	wire [4-1:0] node8025;
	wire [4-1:0] node8028;
	wire [4-1:0] node8029;
	wire [4-1:0] node8032;
	wire [4-1:0] node8035;
	wire [4-1:0] node8036;
	wire [4-1:0] node8037;
	wire [4-1:0] node8038;
	wire [4-1:0] node8041;
	wire [4-1:0] node8044;
	wire [4-1:0] node8046;
	wire [4-1:0] node8048;
	wire [4-1:0] node8051;
	wire [4-1:0] node8052;
	wire [4-1:0] node8053;
	wire [4-1:0] node8054;
	wire [4-1:0] node8059;
	wire [4-1:0] node8060;
	wire [4-1:0] node8064;
	wire [4-1:0] node8065;
	wire [4-1:0] node8066;
	wire [4-1:0] node8067;
	wire [4-1:0] node8069;
	wire [4-1:0] node8072;
	wire [4-1:0] node8073;
	wire [4-1:0] node8074;
	wire [4-1:0] node8078;
	wire [4-1:0] node8079;
	wire [4-1:0] node8083;
	wire [4-1:0] node8084;
	wire [4-1:0] node8085;
	wire [4-1:0] node8088;
	wire [4-1:0] node8091;
	wire [4-1:0] node8092;
	wire [4-1:0] node8095;
	wire [4-1:0] node8098;
	wire [4-1:0] node8099;
	wire [4-1:0] node8100;
	wire [4-1:0] node8101;
	wire [4-1:0] node8102;
	wire [4-1:0] node8106;
	wire [4-1:0] node8107;
	wire [4-1:0] node8111;
	wire [4-1:0] node8112;
	wire [4-1:0] node8113;
	wire [4-1:0] node8117;
	wire [4-1:0] node8120;
	wire [4-1:0] node8121;
	wire [4-1:0] node8122;
	wire [4-1:0] node8125;
	wire [4-1:0] node8128;
	wire [4-1:0] node8129;
	wire [4-1:0] node8130;
	wire [4-1:0] node8135;
	wire [4-1:0] node8136;
	wire [4-1:0] node8137;
	wire [4-1:0] node8138;
	wire [4-1:0] node8139;
	wire [4-1:0] node8140;
	wire [4-1:0] node8141;
	wire [4-1:0] node8144;
	wire [4-1:0] node8146;
	wire [4-1:0] node8149;
	wire [4-1:0] node8150;
	wire [4-1:0] node8153;
	wire [4-1:0] node8154;
	wire [4-1:0] node8158;
	wire [4-1:0] node8159;
	wire [4-1:0] node8160;
	wire [4-1:0] node8162;
	wire [4-1:0] node8165;
	wire [4-1:0] node8166;
	wire [4-1:0] node8169;
	wire [4-1:0] node8172;
	wire [4-1:0] node8173;
	wire [4-1:0] node8176;
	wire [4-1:0] node8179;
	wire [4-1:0] node8180;
	wire [4-1:0] node8181;
	wire [4-1:0] node8182;
	wire [4-1:0] node8183;
	wire [4-1:0] node8186;
	wire [4-1:0] node8189;
	wire [4-1:0] node8190;
	wire [4-1:0] node8193;
	wire [4-1:0] node8195;
	wire [4-1:0] node8198;
	wire [4-1:0] node8199;
	wire [4-1:0] node8200;
	wire [4-1:0] node8201;
	wire [4-1:0] node8204;
	wire [4-1:0] node8207;
	wire [4-1:0] node8208;
	wire [4-1:0] node8211;
	wire [4-1:0] node8214;
	wire [4-1:0] node8215;
	wire [4-1:0] node8218;
	wire [4-1:0] node8221;
	wire [4-1:0] node8222;
	wire [4-1:0] node8223;
	wire [4-1:0] node8224;
	wire [4-1:0] node8227;
	wire [4-1:0] node8229;
	wire [4-1:0] node8232;
	wire [4-1:0] node8233;
	wire [4-1:0] node8234;
	wire [4-1:0] node8237;
	wire [4-1:0] node8240;
	wire [4-1:0] node8242;
	wire [4-1:0] node8245;
	wire [4-1:0] node8246;
	wire [4-1:0] node8247;
	wire [4-1:0] node8250;
	wire [4-1:0] node8253;
	wire [4-1:0] node8254;
	wire [4-1:0] node8256;
	wire [4-1:0] node8259;
	wire [4-1:0] node8262;
	wire [4-1:0] node8263;
	wire [4-1:0] node8264;
	wire [4-1:0] node8265;
	wire [4-1:0] node8266;
	wire [4-1:0] node8267;
	wire [4-1:0] node8268;
	wire [4-1:0] node8272;
	wire [4-1:0] node8273;
	wire [4-1:0] node8277;
	wire [4-1:0] node8278;
	wire [4-1:0] node8281;
	wire [4-1:0] node8284;
	wire [4-1:0] node8285;
	wire [4-1:0] node8286;
	wire [4-1:0] node8287;
	wire [4-1:0] node8290;
	wire [4-1:0] node8293;
	wire [4-1:0] node8295;
	wire [4-1:0] node8298;
	wire [4-1:0] node8299;
	wire [4-1:0] node8302;
	wire [4-1:0] node8305;
	wire [4-1:0] node8306;
	wire [4-1:0] node8307;
	wire [4-1:0] node8308;
	wire [4-1:0] node8311;
	wire [4-1:0] node8314;
	wire [4-1:0] node8315;
	wire [4-1:0] node8318;
	wire [4-1:0] node8321;
	wire [4-1:0] node8322;
	wire [4-1:0] node8323;
	wire [4-1:0] node8326;
	wire [4-1:0] node8329;
	wire [4-1:0] node8330;
	wire [4-1:0] node8333;
	wire [4-1:0] node8336;
	wire [4-1:0] node8337;
	wire [4-1:0] node8338;
	wire [4-1:0] node8339;
	wire [4-1:0] node8340;
	wire [4-1:0] node8343;
	wire [4-1:0] node8346;
	wire [4-1:0] node8347;
	wire [4-1:0] node8348;
	wire [4-1:0] node8352;
	wire [4-1:0] node8355;
	wire [4-1:0] node8356;
	wire [4-1:0] node8357;
	wire [4-1:0] node8359;
	wire [4-1:0] node8363;
	wire [4-1:0] node8364;
	wire [4-1:0] node8365;
	wire [4-1:0] node8368;
	wire [4-1:0] node8371;
	wire [4-1:0] node8373;
	wire [4-1:0] node8376;
	wire [4-1:0] node8377;
	wire [4-1:0] node8378;
	wire [4-1:0] node8379;
	wire [4-1:0] node8381;
	wire [4-1:0] node8384;
	wire [4-1:0] node8385;
	wire [4-1:0] node8388;
	wire [4-1:0] node8391;
	wire [4-1:0] node8392;
	wire [4-1:0] node8393;
	wire [4-1:0] node8396;
	wire [4-1:0] node8399;
	wire [4-1:0] node8400;
	wire [4-1:0] node8404;
	wire [4-1:0] node8405;
	wire [4-1:0] node8406;
	wire [4-1:0] node8407;
	wire [4-1:0] node8410;
	wire [4-1:0] node8414;
	wire [4-1:0] node8415;
	wire [4-1:0] node8418;
	wire [4-1:0] node8421;
	wire [4-1:0] node8422;
	wire [4-1:0] node8423;
	wire [4-1:0] node8424;
	wire [4-1:0] node8425;
	wire [4-1:0] node8426;
	wire [4-1:0] node8427;
	wire [4-1:0] node8430;
	wire [4-1:0] node8433;
	wire [4-1:0] node8435;
	wire [4-1:0] node8436;
	wire [4-1:0] node8440;
	wire [4-1:0] node8441;
	wire [4-1:0] node8444;
	wire [4-1:0] node8447;
	wire [4-1:0] node8448;
	wire [4-1:0] node8449;
	wire [4-1:0] node8452;
	wire [4-1:0] node8455;
	wire [4-1:0] node8456;
	wire [4-1:0] node8459;
	wire [4-1:0] node8462;
	wire [4-1:0] node8463;
	wire [4-1:0] node8464;
	wire [4-1:0] node8465;
	wire [4-1:0] node8468;
	wire [4-1:0] node8471;
	wire [4-1:0] node8472;
	wire [4-1:0] node8473;
	wire [4-1:0] node8476;
	wire [4-1:0] node8479;
	wire [4-1:0] node8480;
	wire [4-1:0] node8484;
	wire [4-1:0] node8485;
	wire [4-1:0] node8486;
	wire [4-1:0] node8489;
	wire [4-1:0] node8492;
	wire [4-1:0] node8493;
	wire [4-1:0] node8494;
	wire [4-1:0] node8498;
	wire [4-1:0] node8500;
	wire [4-1:0] node8501;
	wire [4-1:0] node8504;
	wire [4-1:0] node8507;
	wire [4-1:0] node8508;
	wire [4-1:0] node8509;
	wire [4-1:0] node8510;
	wire [4-1:0] node8511;
	wire [4-1:0] node8512;
	wire [4-1:0] node8515;
	wire [4-1:0] node8518;
	wire [4-1:0] node8519;
	wire [4-1:0] node8522;
	wire [4-1:0] node8525;
	wire [4-1:0] node8526;
	wire [4-1:0] node8527;
	wire [4-1:0] node8530;
	wire [4-1:0] node8533;
	wire [4-1:0] node8534;
	wire [4-1:0] node8537;
	wire [4-1:0] node8540;
	wire [4-1:0] node8541;
	wire [4-1:0] node8542;
	wire [4-1:0] node8543;
	wire [4-1:0] node8546;
	wire [4-1:0] node8549;
	wire [4-1:0] node8550;
	wire [4-1:0] node8553;
	wire [4-1:0] node8556;
	wire [4-1:0] node8557;
	wire [4-1:0] node8559;
	wire [4-1:0] node8560;
	wire [4-1:0] node8563;
	wire [4-1:0] node8566;
	wire [4-1:0] node8567;
	wire [4-1:0] node8570;
	wire [4-1:0] node8573;
	wire [4-1:0] node8574;
	wire [4-1:0] node8575;
	wire [4-1:0] node8576;
	wire [4-1:0] node8577;
	wire [4-1:0] node8580;
	wire [4-1:0] node8583;
	wire [4-1:0] node8584;
	wire [4-1:0] node8588;
	wire [4-1:0] node8589;
	wire [4-1:0] node8592;
	wire [4-1:0] node8595;
	wire [4-1:0] node8596;
	wire [4-1:0] node8597;
	wire [4-1:0] node8598;
	wire [4-1:0] node8602;
	wire [4-1:0] node8603;
	wire [4-1:0] node8604;
	wire [4-1:0] node8607;
	wire [4-1:0] node8611;
	wire [4-1:0] node8612;
	wire [4-1:0] node8613;
	wire [4-1:0] node8616;
	wire [4-1:0] node8619;
	wire [4-1:0] node8620;
	wire [4-1:0] node8621;
	wire [4-1:0] node8625;
	wire [4-1:0] node8626;
	wire [4-1:0] node8630;
	wire [4-1:0] node8631;
	wire [4-1:0] node8632;
	wire [4-1:0] node8633;
	wire [4-1:0] node8634;
	wire [4-1:0] node8635;
	wire [4-1:0] node8636;
	wire [4-1:0] node8637;
	wire [4-1:0] node8638;
	wire [4-1:0] node8639;
	wire [4-1:0] node8640;
	wire [4-1:0] node8641;
	wire [4-1:0] node8645;
	wire [4-1:0] node8647;
	wire [4-1:0] node8650;
	wire [4-1:0] node8651;
	wire [4-1:0] node8653;
	wire [4-1:0] node8656;
	wire [4-1:0] node8657;
	wire [4-1:0] node8659;
	wire [4-1:0] node8662;
	wire [4-1:0] node8663;
	wire [4-1:0] node8666;
	wire [4-1:0] node8669;
	wire [4-1:0] node8670;
	wire [4-1:0] node8671;
	wire [4-1:0] node8672;
	wire [4-1:0] node8673;
	wire [4-1:0] node8678;
	wire [4-1:0] node8679;
	wire [4-1:0] node8681;
	wire [4-1:0] node8684;
	wire [4-1:0] node8685;
	wire [4-1:0] node8688;
	wire [4-1:0] node8691;
	wire [4-1:0] node8692;
	wire [4-1:0] node8693;
	wire [4-1:0] node8694;
	wire [4-1:0] node8698;
	wire [4-1:0] node8699;
	wire [4-1:0] node8702;
	wire [4-1:0] node8705;
	wire [4-1:0] node8706;
	wire [4-1:0] node8707;
	wire [4-1:0] node8712;
	wire [4-1:0] node8713;
	wire [4-1:0] node8714;
	wire [4-1:0] node8715;
	wire [4-1:0] node8717;
	wire [4-1:0] node8719;
	wire [4-1:0] node8722;
	wire [4-1:0] node8724;
	wire [4-1:0] node8726;
	wire [4-1:0] node8729;
	wire [4-1:0] node8730;
	wire [4-1:0] node8731;
	wire [4-1:0] node8734;
	wire [4-1:0] node8737;
	wire [4-1:0] node8739;
	wire [4-1:0] node8741;
	wire [4-1:0] node8744;
	wire [4-1:0] node8745;
	wire [4-1:0] node8747;
	wire [4-1:0] node8748;
	wire [4-1:0] node8751;
	wire [4-1:0] node8753;
	wire [4-1:0] node8756;
	wire [4-1:0] node8757;
	wire [4-1:0] node8758;
	wire [4-1:0] node8759;
	wire [4-1:0] node8762;
	wire [4-1:0] node8766;
	wire [4-1:0] node8767;
	wire [4-1:0] node8768;
	wire [4-1:0] node8771;
	wire [4-1:0] node8774;
	wire [4-1:0] node8775;
	wire [4-1:0] node8778;
	wire [4-1:0] node8781;
	wire [4-1:0] node8782;
	wire [4-1:0] node8783;
	wire [4-1:0] node8784;
	wire [4-1:0] node8785;
	wire [4-1:0] node8787;
	wire [4-1:0] node8790;
	wire [4-1:0] node8791;
	wire [4-1:0] node8793;
	wire [4-1:0] node8796;
	wire [4-1:0] node8798;
	wire [4-1:0] node8801;
	wire [4-1:0] node8802;
	wire [4-1:0] node8803;
	wire [4-1:0] node8806;
	wire [4-1:0] node8809;
	wire [4-1:0] node8811;
	wire [4-1:0] node8814;
	wire [4-1:0] node8815;
	wire [4-1:0] node8816;
	wire [4-1:0] node8817;
	wire [4-1:0] node8821;
	wire [4-1:0] node8822;
	wire [4-1:0] node8824;
	wire [4-1:0] node8828;
	wire [4-1:0] node8829;
	wire [4-1:0] node8831;
	wire [4-1:0] node8832;
	wire [4-1:0] node8836;
	wire [4-1:0] node8838;
	wire [4-1:0] node8839;
	wire [4-1:0] node8843;
	wire [4-1:0] node8844;
	wire [4-1:0] node8845;
	wire [4-1:0] node8847;
	wire [4-1:0] node8848;
	wire [4-1:0] node8849;
	wire [4-1:0] node8853;
	wire [4-1:0] node8856;
	wire [4-1:0] node8857;
	wire [4-1:0] node8858;
	wire [4-1:0] node8859;
	wire [4-1:0] node8862;
	wire [4-1:0] node8865;
	wire [4-1:0] node8868;
	wire [4-1:0] node8869;
	wire [4-1:0] node8872;
	wire [4-1:0] node8875;
	wire [4-1:0] node8876;
	wire [4-1:0] node8877;
	wire [4-1:0] node8878;
	wire [4-1:0] node8879;
	wire [4-1:0] node8883;
	wire [4-1:0] node8885;
	wire [4-1:0] node8888;
	wire [4-1:0] node8889;
	wire [4-1:0] node8890;
	wire [4-1:0] node8893;
	wire [4-1:0] node8897;
	wire [4-1:0] node8898;
	wire [4-1:0] node8899;
	wire [4-1:0] node8901;
	wire [4-1:0] node8904;
	wire [4-1:0] node8905;
	wire [4-1:0] node8909;
	wire [4-1:0] node8910;
	wire [4-1:0] node8911;
	wire [4-1:0] node8914;
	wire [4-1:0] node8917;
	wire [4-1:0] node8918;
	wire [4-1:0] node8921;
	wire [4-1:0] node8924;
	wire [4-1:0] node8925;
	wire [4-1:0] node8926;
	wire [4-1:0] node8927;
	wire [4-1:0] node8928;
	wire [4-1:0] node8929;
	wire [4-1:0] node8930;
	wire [4-1:0] node8931;
	wire [4-1:0] node8934;
	wire [4-1:0] node8937;
	wire [4-1:0] node8938;
	wire [4-1:0] node8942;
	wire [4-1:0] node8943;
	wire [4-1:0] node8946;
	wire [4-1:0] node8948;
	wire [4-1:0] node8951;
	wire [4-1:0] node8952;
	wire [4-1:0] node8953;
	wire [4-1:0] node8956;
	wire [4-1:0] node8959;
	wire [4-1:0] node8960;
	wire [4-1:0] node8962;
	wire [4-1:0] node8965;
	wire [4-1:0] node8966;
	wire [4-1:0] node8969;
	wire [4-1:0] node8972;
	wire [4-1:0] node8973;
	wire [4-1:0] node8974;
	wire [4-1:0] node8975;
	wire [4-1:0] node8976;
	wire [4-1:0] node8979;
	wire [4-1:0] node8982;
	wire [4-1:0] node8983;
	wire [4-1:0] node8986;
	wire [4-1:0] node8989;
	wire [4-1:0] node8990;
	wire [4-1:0] node8993;
	wire [4-1:0] node8996;
	wire [4-1:0] node8997;
	wire [4-1:0] node8998;
	wire [4-1:0] node9001;
	wire [4-1:0] node9004;
	wire [4-1:0] node9005;
	wire [4-1:0] node9007;
	wire [4-1:0] node9010;
	wire [4-1:0] node9011;
	wire [4-1:0] node9014;
	wire [4-1:0] node9017;
	wire [4-1:0] node9018;
	wire [4-1:0] node9019;
	wire [4-1:0] node9020;
	wire [4-1:0] node9024;
	wire [4-1:0] node9025;
	wire [4-1:0] node9026;
	wire [4-1:0] node9030;
	wire [4-1:0] node9031;
	wire [4-1:0] node9034;
	wire [4-1:0] node9037;
	wire [4-1:0] node9038;
	wire [4-1:0] node9039;
	wire [4-1:0] node9041;
	wire [4-1:0] node9045;
	wire [4-1:0] node9046;
	wire [4-1:0] node9048;
	wire [4-1:0] node9051;
	wire [4-1:0] node9052;
	wire [4-1:0] node9056;
	wire [4-1:0] node9057;
	wire [4-1:0] node9058;
	wire [4-1:0] node9059;
	wire [4-1:0] node9060;
	wire [4-1:0] node9061;
	wire [4-1:0] node9065;
	wire [4-1:0] node9066;
	wire [4-1:0] node9067;
	wire [4-1:0] node9070;
	wire [4-1:0] node9074;
	wire [4-1:0] node9075;
	wire [4-1:0] node9076;
	wire [4-1:0] node9078;
	wire [4-1:0] node9081;
	wire [4-1:0] node9083;
	wire [4-1:0] node9086;
	wire [4-1:0] node9087;
	wire [4-1:0] node9089;
	wire [4-1:0] node9092;
	wire [4-1:0] node9094;
	wire [4-1:0] node9097;
	wire [4-1:0] node9098;
	wire [4-1:0] node9099;
	wire [4-1:0] node9101;
	wire [4-1:0] node9102;
	wire [4-1:0] node9105;
	wire [4-1:0] node9108;
	wire [4-1:0] node9109;
	wire [4-1:0] node9111;
	wire [4-1:0] node9114;
	wire [4-1:0] node9116;
	wire [4-1:0] node9119;
	wire [4-1:0] node9120;
	wire [4-1:0] node9121;
	wire [4-1:0] node9124;
	wire [4-1:0] node9127;
	wire [4-1:0] node9128;
	wire [4-1:0] node9129;
	wire [4-1:0] node9133;
	wire [4-1:0] node9136;
	wire [4-1:0] node9137;
	wire [4-1:0] node9138;
	wire [4-1:0] node9139;
	wire [4-1:0] node9140;
	wire [4-1:0] node9144;
	wire [4-1:0] node9145;
	wire [4-1:0] node9146;
	wire [4-1:0] node9150;
	wire [4-1:0] node9152;
	wire [4-1:0] node9155;
	wire [4-1:0] node9156;
	wire [4-1:0] node9158;
	wire [4-1:0] node9159;
	wire [4-1:0] node9163;
	wire [4-1:0] node9164;
	wire [4-1:0] node9167;
	wire [4-1:0] node9169;
	wire [4-1:0] node9172;
	wire [4-1:0] node9173;
	wire [4-1:0] node9174;
	wire [4-1:0] node9175;
	wire [4-1:0] node9177;
	wire [4-1:0] node9180;
	wire [4-1:0] node9181;
	wire [4-1:0] node9185;
	wire [4-1:0] node9186;
	wire [4-1:0] node9189;
	wire [4-1:0] node9192;
	wire [4-1:0] node9194;
	wire [4-1:0] node9195;
	wire [4-1:0] node9196;
	wire [4-1:0] node9200;
	wire [4-1:0] node9203;
	wire [4-1:0] node9204;
	wire [4-1:0] node9205;
	wire [4-1:0] node9206;
	wire [4-1:0] node9207;
	wire [4-1:0] node9208;
	wire [4-1:0] node9210;
	wire [4-1:0] node9213;
	wire [4-1:0] node9215;
	wire [4-1:0] node9218;
	wire [4-1:0] node9219;
	wire [4-1:0] node9221;
	wire [4-1:0] node9224;
	wire [4-1:0] node9226;
	wire [4-1:0] node9229;
	wire [4-1:0] node9230;
	wire [4-1:0] node9231;
	wire [4-1:0] node9232;
	wire [4-1:0] node9235;
	wire [4-1:0] node9238;
	wire [4-1:0] node9239;
	wire [4-1:0] node9240;
	wire [4-1:0] node9242;
	wire [4-1:0] node9245;
	wire [4-1:0] node9248;
	wire [4-1:0] node9249;
	wire [4-1:0] node9250;
	wire [4-1:0] node9253;
	wire [4-1:0] node9256;
	wire [4-1:0] node9257;
	wire [4-1:0] node9260;
	wire [4-1:0] node9263;
	wire [4-1:0] node9264;
	wire [4-1:0] node9265;
	wire [4-1:0] node9266;
	wire [4-1:0] node9269;
	wire [4-1:0] node9273;
	wire [4-1:0] node9274;
	wire [4-1:0] node9276;
	wire [4-1:0] node9277;
	wire [4-1:0] node9280;
	wire [4-1:0] node9283;
	wire [4-1:0] node9286;
	wire [4-1:0] node9287;
	wire [4-1:0] node9288;
	wire [4-1:0] node9289;
	wire [4-1:0] node9292;
	wire [4-1:0] node9295;
	wire [4-1:0] node9296;
	wire [4-1:0] node9297;
	wire [4-1:0] node9299;
	wire [4-1:0] node9302;
	wire [4-1:0] node9303;
	wire [4-1:0] node9307;
	wire [4-1:0] node9308;
	wire [4-1:0] node9309;
	wire [4-1:0] node9310;
	wire [4-1:0] node9313;
	wire [4-1:0] node9316;
	wire [4-1:0] node9318;
	wire [4-1:0] node9321;
	wire [4-1:0] node9322;
	wire [4-1:0] node9326;
	wire [4-1:0] node9327;
	wire [4-1:0] node9328;
	wire [4-1:0] node9329;
	wire [4-1:0] node9332;
	wire [4-1:0] node9335;
	wire [4-1:0] node9336;
	wire [4-1:0] node9337;
	wire [4-1:0] node9339;
	wire [4-1:0] node9343;
	wire [4-1:0] node9344;
	wire [4-1:0] node9345;
	wire [4-1:0] node9348;
	wire [4-1:0] node9352;
	wire [4-1:0] node9353;
	wire [4-1:0] node9354;
	wire [4-1:0] node9355;
	wire [4-1:0] node9358;
	wire [4-1:0] node9361;
	wire [4-1:0] node9362;
	wire [4-1:0] node9363;
	wire [4-1:0] node9366;
	wire [4-1:0] node9369;
	wire [4-1:0] node9370;
	wire [4-1:0] node9373;
	wire [4-1:0] node9376;
	wire [4-1:0] node9377;
	wire [4-1:0] node9380;
	wire [4-1:0] node9383;
	wire [4-1:0] node9384;
	wire [4-1:0] node9385;
	wire [4-1:0] node9386;
	wire [4-1:0] node9387;
	wire [4-1:0] node9390;
	wire [4-1:0] node9393;
	wire [4-1:0] node9394;
	wire [4-1:0] node9395;
	wire [4-1:0] node9396;
	wire [4-1:0] node9399;
	wire [4-1:0] node9402;
	wire [4-1:0] node9403;
	wire [4-1:0] node9406;
	wire [4-1:0] node9409;
	wire [4-1:0] node9411;
	wire [4-1:0] node9412;
	wire [4-1:0] node9415;
	wire [4-1:0] node9418;
	wire [4-1:0] node9419;
	wire [4-1:0] node9420;
	wire [4-1:0] node9421;
	wire [4-1:0] node9422;
	wire [4-1:0] node9424;
	wire [4-1:0] node9427;
	wire [4-1:0] node9429;
	wire [4-1:0] node9432;
	wire [4-1:0] node9435;
	wire [4-1:0] node9437;
	wire [4-1:0] node9438;
	wire [4-1:0] node9441;
	wire [4-1:0] node9443;
	wire [4-1:0] node9446;
	wire [4-1:0] node9447;
	wire [4-1:0] node9448;
	wire [4-1:0] node9449;
	wire [4-1:0] node9452;
	wire [4-1:0] node9455;
	wire [4-1:0] node9456;
	wire [4-1:0] node9459;
	wire [4-1:0] node9462;
	wire [4-1:0] node9463;
	wire [4-1:0] node9464;
	wire [4-1:0] node9467;
	wire [4-1:0] node9470;
	wire [4-1:0] node9471;
	wire [4-1:0] node9475;
	wire [4-1:0] node9476;
	wire [4-1:0] node9477;
	wire [4-1:0] node9478;
	wire [4-1:0] node9479;
	wire [4-1:0] node9480;
	wire [4-1:0] node9483;
	wire [4-1:0] node9486;
	wire [4-1:0] node9487;
	wire [4-1:0] node9490;
	wire [4-1:0] node9493;
	wire [4-1:0] node9494;
	wire [4-1:0] node9497;
	wire [4-1:0] node9500;
	wire [4-1:0] node9501;
	wire [4-1:0] node9503;
	wire [4-1:0] node9504;
	wire [4-1:0] node9506;
	wire [4-1:0] node9509;
	wire [4-1:0] node9510;
	wire [4-1:0] node9513;
	wire [4-1:0] node9516;
	wire [4-1:0] node9517;
	wire [4-1:0] node9520;
	wire [4-1:0] node9523;
	wire [4-1:0] node9524;
	wire [4-1:0] node9525;
	wire [4-1:0] node9526;
	wire [4-1:0] node9527;
	wire [4-1:0] node9530;
	wire [4-1:0] node9534;
	wire [4-1:0] node9535;
	wire [4-1:0] node9536;
	wire [4-1:0] node9540;
	wire [4-1:0] node9541;
	wire [4-1:0] node9545;
	wire [4-1:0] node9546;
	wire [4-1:0] node9547;
	wire [4-1:0] node9548;
	wire [4-1:0] node9552;
	wire [4-1:0] node9553;
	wire [4-1:0] node9557;
	wire [4-1:0] node9559;
	wire [4-1:0] node9560;
	wire [4-1:0] node9564;
	wire [4-1:0] node9565;
	wire [4-1:0] node9566;
	wire [4-1:0] node9567;
	wire [4-1:0] node9568;
	wire [4-1:0] node9569;
	wire [4-1:0] node9570;
	wire [4-1:0] node9571;
	wire [4-1:0] node9574;
	wire [4-1:0] node9576;
	wire [4-1:0] node9579;
	wire [4-1:0] node9580;
	wire [4-1:0] node9581;
	wire [4-1:0] node9584;
	wire [4-1:0] node9587;
	wire [4-1:0] node9588;
	wire [4-1:0] node9591;
	wire [4-1:0] node9594;
	wire [4-1:0] node9595;
	wire [4-1:0] node9596;
	wire [4-1:0] node9599;
	wire [4-1:0] node9601;
	wire [4-1:0] node9604;
	wire [4-1:0] node9605;
	wire [4-1:0] node9606;
	wire [4-1:0] node9609;
	wire [4-1:0] node9612;
	wire [4-1:0] node9613;
	wire [4-1:0] node9616;
	wire [4-1:0] node9619;
	wire [4-1:0] node9620;
	wire [4-1:0] node9621;
	wire [4-1:0] node9622;
	wire [4-1:0] node9625;
	wire [4-1:0] node9627;
	wire [4-1:0] node9630;
	wire [4-1:0] node9631;
	wire [4-1:0] node9632;
	wire [4-1:0] node9635;
	wire [4-1:0] node9638;
	wire [4-1:0] node9640;
	wire [4-1:0] node9641;
	wire [4-1:0] node9644;
	wire [4-1:0] node9647;
	wire [4-1:0] node9648;
	wire [4-1:0] node9649;
	wire [4-1:0] node9652;
	wire [4-1:0] node9654;
	wire [4-1:0] node9657;
	wire [4-1:0] node9658;
	wire [4-1:0] node9659;
	wire [4-1:0] node9662;
	wire [4-1:0] node9665;
	wire [4-1:0] node9666;
	wire [4-1:0] node9669;
	wire [4-1:0] node9672;
	wire [4-1:0] node9673;
	wire [4-1:0] node9674;
	wire [4-1:0] node9675;
	wire [4-1:0] node9676;
	wire [4-1:0] node9677;
	wire [4-1:0] node9678;
	wire [4-1:0] node9682;
	wire [4-1:0] node9684;
	wire [4-1:0] node9687;
	wire [4-1:0] node9689;
	wire [4-1:0] node9692;
	wire [4-1:0] node9693;
	wire [4-1:0] node9695;
	wire [4-1:0] node9698;
	wire [4-1:0] node9700;
	wire [4-1:0] node9701;
	wire [4-1:0] node9705;
	wire [4-1:0] node9706;
	wire [4-1:0] node9707;
	wire [4-1:0] node9708;
	wire [4-1:0] node9709;
	wire [4-1:0] node9712;
	wire [4-1:0] node9715;
	wire [4-1:0] node9717;
	wire [4-1:0] node9720;
	wire [4-1:0] node9723;
	wire [4-1:0] node9724;
	wire [4-1:0] node9725;
	wire [4-1:0] node9728;
	wire [4-1:0] node9729;
	wire [4-1:0] node9732;
	wire [4-1:0] node9735;
	wire [4-1:0] node9736;
	wire [4-1:0] node9737;
	wire [4-1:0] node9740;
	wire [4-1:0] node9743;
	wire [4-1:0] node9744;
	wire [4-1:0] node9747;
	wire [4-1:0] node9750;
	wire [4-1:0] node9751;
	wire [4-1:0] node9752;
	wire [4-1:0] node9753;
	wire [4-1:0] node9754;
	wire [4-1:0] node9755;
	wire [4-1:0] node9760;
	wire [4-1:0] node9761;
	wire [4-1:0] node9762;
	wire [4-1:0] node9765;
	wire [4-1:0] node9768;
	wire [4-1:0] node9770;
	wire [4-1:0] node9773;
	wire [4-1:0] node9774;
	wire [4-1:0] node9775;
	wire [4-1:0] node9776;
	wire [4-1:0] node9779;
	wire [4-1:0] node9782;
	wire [4-1:0] node9784;
	wire [4-1:0] node9787;
	wire [4-1:0] node9788;
	wire [4-1:0] node9790;
	wire [4-1:0] node9793;
	wire [4-1:0] node9794;
	wire [4-1:0] node9797;
	wire [4-1:0] node9800;
	wire [4-1:0] node9801;
	wire [4-1:0] node9802;
	wire [4-1:0] node9804;
	wire [4-1:0] node9806;
	wire [4-1:0] node9809;
	wire [4-1:0] node9810;
	wire [4-1:0] node9811;
	wire [4-1:0] node9815;
	wire [4-1:0] node9816;
	wire [4-1:0] node9819;
	wire [4-1:0] node9822;
	wire [4-1:0] node9823;
	wire [4-1:0] node9827;
	wire [4-1:0] node9828;
	wire [4-1:0] node9829;
	wire [4-1:0] node9830;
	wire [4-1:0] node9831;
	wire [4-1:0] node9832;
	wire [4-1:0] node9833;
	wire [4-1:0] node9835;
	wire [4-1:0] node9838;
	wire [4-1:0] node9840;
	wire [4-1:0] node9843;
	wire [4-1:0] node9844;
	wire [4-1:0] node9846;
	wire [4-1:0] node9849;
	wire [4-1:0] node9851;
	wire [4-1:0] node9854;
	wire [4-1:0] node9855;
	wire [4-1:0] node9856;
	wire [4-1:0] node9858;
	wire [4-1:0] node9861;
	wire [4-1:0] node9863;
	wire [4-1:0] node9866;
	wire [4-1:0] node9868;
	wire [4-1:0] node9869;
	wire [4-1:0] node9872;
	wire [4-1:0] node9875;
	wire [4-1:0] node9876;
	wire [4-1:0] node9877;
	wire [4-1:0] node9878;
	wire [4-1:0] node9880;
	wire [4-1:0] node9884;
	wire [4-1:0] node9885;
	wire [4-1:0] node9888;
	wire [4-1:0] node9891;
	wire [4-1:0] node9892;
	wire [4-1:0] node9893;
	wire [4-1:0] node9896;
	wire [4-1:0] node9899;
	wire [4-1:0] node9901;
	wire [4-1:0] node9904;
	wire [4-1:0] node9905;
	wire [4-1:0] node9906;
	wire [4-1:0] node9907;
	wire [4-1:0] node9908;
	wire [4-1:0] node9911;
	wire [4-1:0] node9913;
	wire [4-1:0] node9916;
	wire [4-1:0] node9917;
	wire [4-1:0] node9921;
	wire [4-1:0] node9922;
	wire [4-1:0] node9924;
	wire [4-1:0] node9925;
	wire [4-1:0] node9929;
	wire [4-1:0] node9931;
	wire [4-1:0] node9933;
	wire [4-1:0] node9936;
	wire [4-1:0] node9937;
	wire [4-1:0] node9938;
	wire [4-1:0] node9939;
	wire [4-1:0] node9942;
	wire [4-1:0] node9946;
	wire [4-1:0] node9947;
	wire [4-1:0] node9948;
	wire [4-1:0] node9950;
	wire [4-1:0] node9953;
	wire [4-1:0] node9956;
	wire [4-1:0] node9958;
	wire [4-1:0] node9960;
	wire [4-1:0] node9963;
	wire [4-1:0] node9964;
	wire [4-1:0] node9965;
	wire [4-1:0] node9966;
	wire [4-1:0] node9967;
	wire [4-1:0] node9968;
	wire [4-1:0] node9972;
	wire [4-1:0] node9973;
	wire [4-1:0] node9974;
	wire [4-1:0] node9977;
	wire [4-1:0] node9980;
	wire [4-1:0] node9982;
	wire [4-1:0] node9985;
	wire [4-1:0] node9986;
	wire [4-1:0] node9987;
	wire [4-1:0] node9988;
	wire [4-1:0] node9992;
	wire [4-1:0] node9993;
	wire [4-1:0] node9996;
	wire [4-1:0] node9999;
	wire [4-1:0] node10000;
	wire [4-1:0] node10001;
	wire [4-1:0] node10004;
	wire [4-1:0] node10007;
	wire [4-1:0] node10008;
	wire [4-1:0] node10012;
	wire [4-1:0] node10013;
	wire [4-1:0] node10014;
	wire [4-1:0] node10015;
	wire [4-1:0] node10019;
	wire [4-1:0] node10020;
	wire [4-1:0] node10021;
	wire [4-1:0] node10024;
	wire [4-1:0] node10027;
	wire [4-1:0] node10030;
	wire [4-1:0] node10031;
	wire [4-1:0] node10032;
	wire [4-1:0] node10033;
	wire [4-1:0] node10036;
	wire [4-1:0] node10040;
	wire [4-1:0] node10041;
	wire [4-1:0] node10042;
	wire [4-1:0] node10045;
	wire [4-1:0] node10048;
	wire [4-1:0] node10049;
	wire [4-1:0] node10052;
	wire [4-1:0] node10055;
	wire [4-1:0] node10056;
	wire [4-1:0] node10057;
	wire [4-1:0] node10058;
	wire [4-1:0] node10059;
	wire [4-1:0] node10061;
	wire [4-1:0] node10064;
	wire [4-1:0] node10066;
	wire [4-1:0] node10069;
	wire [4-1:0] node10070;
	wire [4-1:0] node10074;
	wire [4-1:0] node10075;
	wire [4-1:0] node10077;
	wire [4-1:0] node10079;
	wire [4-1:0] node10082;
	wire [4-1:0] node10083;
	wire [4-1:0] node10087;
	wire [4-1:0] node10088;
	wire [4-1:0] node10089;
	wire [4-1:0] node10090;
	wire [4-1:0] node10094;
	wire [4-1:0] node10095;
	wire [4-1:0] node10097;
	wire [4-1:0] node10101;
	wire [4-1:0] node10102;
	wire [4-1:0] node10103;
	wire [4-1:0] node10106;
	wire [4-1:0] node10109;
	wire [4-1:0] node10110;
	wire [4-1:0] node10111;
	wire [4-1:0] node10114;
	wire [4-1:0] node10117;
	wire [4-1:0] node10118;
	wire [4-1:0] node10121;
	wire [4-1:0] node10124;
	wire [4-1:0] node10125;
	wire [4-1:0] node10126;
	wire [4-1:0] node10127;
	wire [4-1:0] node10128;
	wire [4-1:0] node10129;
	wire [4-1:0] node10130;
	wire [4-1:0] node10131;
	wire [4-1:0] node10134;
	wire [4-1:0] node10137;
	wire [4-1:0] node10138;
	wire [4-1:0] node10139;
	wire [4-1:0] node10142;
	wire [4-1:0] node10145;
	wire [4-1:0] node10147;
	wire [4-1:0] node10150;
	wire [4-1:0] node10151;
	wire [4-1:0] node10152;
	wire [4-1:0] node10154;
	wire [4-1:0] node10157;
	wire [4-1:0] node10159;
	wire [4-1:0] node10162;
	wire [4-1:0] node10163;
	wire [4-1:0] node10165;
	wire [4-1:0] node10168;
	wire [4-1:0] node10171;
	wire [4-1:0] node10172;
	wire [4-1:0] node10173;
	wire [4-1:0] node10175;
	wire [4-1:0] node10178;
	wire [4-1:0] node10180;
	wire [4-1:0] node10183;
	wire [4-1:0] node10184;
	wire [4-1:0] node10186;
	wire [4-1:0] node10189;
	wire [4-1:0] node10191;
	wire [4-1:0] node10194;
	wire [4-1:0] node10195;
	wire [4-1:0] node10196;
	wire [4-1:0] node10198;
	wire [4-1:0] node10199;
	wire [4-1:0] node10201;
	wire [4-1:0] node10204;
	wire [4-1:0] node10205;
	wire [4-1:0] node10208;
	wire [4-1:0] node10211;
	wire [4-1:0] node10212;
	wire [4-1:0] node10213;
	wire [4-1:0] node10216;
	wire [4-1:0] node10219;
	wire [4-1:0] node10220;
	wire [4-1:0] node10221;
	wire [4-1:0] node10224;
	wire [4-1:0] node10227;
	wire [4-1:0] node10228;
	wire [4-1:0] node10231;
	wire [4-1:0] node10234;
	wire [4-1:0] node10235;
	wire [4-1:0] node10236;
	wire [4-1:0] node10239;
	wire [4-1:0] node10242;
	wire [4-1:0] node10243;
	wire [4-1:0] node10245;
	wire [4-1:0] node10248;
	wire [4-1:0] node10249;
	wire [4-1:0] node10250;
	wire [4-1:0] node10253;
	wire [4-1:0] node10256;
	wire [4-1:0] node10257;
	wire [4-1:0] node10260;
	wire [4-1:0] node10263;
	wire [4-1:0] node10264;
	wire [4-1:0] node10265;
	wire [4-1:0] node10266;
	wire [4-1:0] node10268;
	wire [4-1:0] node10271;
	wire [4-1:0] node10273;
	wire [4-1:0] node10276;
	wire [4-1:0] node10277;
	wire [4-1:0] node10279;
	wire [4-1:0] node10282;
	wire [4-1:0] node10284;
	wire [4-1:0] node10287;
	wire [4-1:0] node10288;
	wire [4-1:0] node10289;
	wire [4-1:0] node10290;
	wire [4-1:0] node10292;
	wire [4-1:0] node10295;
	wire [4-1:0] node10297;
	wire [4-1:0] node10300;
	wire [4-1:0] node10301;
	wire [4-1:0] node10303;
	wire [4-1:0] node10306;
	wire [4-1:0] node10309;
	wire [4-1:0] node10310;
	wire [4-1:0] node10311;
	wire [4-1:0] node10312;
	wire [4-1:0] node10316;
	wire [4-1:0] node10317;
	wire [4-1:0] node10321;
	wire [4-1:0] node10322;
	wire [4-1:0] node10323;
	wire [4-1:0] node10327;
	wire [4-1:0] node10329;
	wire [4-1:0] node10332;
	wire [4-1:0] node10333;
	wire [4-1:0] node10334;
	wire [4-1:0] node10335;
	wire [4-1:0] node10336;
	wire [4-1:0] node10337;
	wire [4-1:0] node10340;
	wire [4-1:0] node10343;
	wire [4-1:0] node10344;
	wire [4-1:0] node10347;
	wire [4-1:0] node10350;
	wire [4-1:0] node10351;
	wire [4-1:0] node10352;
	wire [4-1:0] node10353;
	wire [4-1:0] node10357;
	wire [4-1:0] node10358;
	wire [4-1:0] node10362;
	wire [4-1:0] node10363;
	wire [4-1:0] node10366;
	wire [4-1:0] node10369;
	wire [4-1:0] node10370;
	wire [4-1:0] node10371;
	wire [4-1:0] node10372;
	wire [4-1:0] node10373;
	wire [4-1:0] node10375;
	wire [4-1:0] node10379;
	wire [4-1:0] node10381;
	wire [4-1:0] node10383;
	wire [4-1:0] node10386;
	wire [4-1:0] node10387;
	wire [4-1:0] node10388;
	wire [4-1:0] node10390;
	wire [4-1:0] node10393;
	wire [4-1:0] node10395;
	wire [4-1:0] node10398;
	wire [4-1:0] node10399;
	wire [4-1:0] node10403;
	wire [4-1:0] node10404;
	wire [4-1:0] node10405;
	wire [4-1:0] node10406;
	wire [4-1:0] node10410;
	wire [4-1:0] node10411;
	wire [4-1:0] node10415;
	wire [4-1:0] node10416;
	wire [4-1:0] node10419;
	wire [4-1:0] node10420;
	wire [4-1:0] node10424;
	wire [4-1:0] node10425;
	wire [4-1:0] node10426;
	wire [4-1:0] node10427;
	wire [4-1:0] node10428;
	wire [4-1:0] node10429;
	wire [4-1:0] node10433;
	wire [4-1:0] node10434;
	wire [4-1:0] node10438;
	wire [4-1:0] node10439;
	wire [4-1:0] node10440;
	wire [4-1:0] node10444;
	wire [4-1:0] node10445;
	wire [4-1:0] node10446;
	wire [4-1:0] node10450;
	wire [4-1:0] node10452;
	wire [4-1:0] node10455;
	wire [4-1:0] node10456;
	wire [4-1:0] node10457;
	wire [4-1:0] node10460;
	wire [4-1:0] node10461;
	wire [4-1:0] node10465;
	wire [4-1:0] node10466;
	wire [4-1:0] node10467;
	wire [4-1:0] node10471;
	wire [4-1:0] node10474;
	wire [4-1:0] node10475;
	wire [4-1:0] node10476;
	wire [4-1:0] node10477;
	wire [4-1:0] node10478;
	wire [4-1:0] node10482;
	wire [4-1:0] node10483;
	wire [4-1:0] node10487;
	wire [4-1:0] node10488;
	wire [4-1:0] node10489;
	wire [4-1:0] node10493;
	wire [4-1:0] node10494;
	wire [4-1:0] node10498;
	wire [4-1:0] node10499;
	wire [4-1:0] node10500;
	wire [4-1:0] node10501;
	wire [4-1:0] node10502;
	wire [4-1:0] node10505;
	wire [4-1:0] node10509;
	wire [4-1:0] node10510;
	wire [4-1:0] node10513;
	wire [4-1:0] node10516;
	wire [4-1:0] node10518;
	wire [4-1:0] node10519;
	wire [4-1:0] node10521;
	wire [4-1:0] node10524;
	wire [4-1:0] node10527;
	wire [4-1:0] node10528;
	wire [4-1:0] node10529;
	wire [4-1:0] node10530;
	wire [4-1:0] node10531;
	wire [4-1:0] node10532;
	wire [4-1:0] node10533;
	wire [4-1:0] node10534;
	wire [4-1:0] node10535;
	wire [4-1:0] node10536;
	wire [4-1:0] node10539;
	wire [4-1:0] node10542;
	wire [4-1:0] node10543;
	wire [4-1:0] node10547;
	wire [4-1:0] node10548;
	wire [4-1:0] node10549;
	wire [4-1:0] node10552;
	wire [4-1:0] node10555;
	wire [4-1:0] node10557;
	wire [4-1:0] node10560;
	wire [4-1:0] node10561;
	wire [4-1:0] node10563;
	wire [4-1:0] node10564;
	wire [4-1:0] node10565;
	wire [4-1:0] node10569;
	wire [4-1:0] node10570;
	wire [4-1:0] node10574;
	wire [4-1:0] node10575;
	wire [4-1:0] node10576;
	wire [4-1:0] node10579;
	wire [4-1:0] node10582;
	wire [4-1:0] node10583;
	wire [4-1:0] node10584;
	wire [4-1:0] node10587;
	wire [4-1:0] node10590;
	wire [4-1:0] node10591;
	wire [4-1:0] node10595;
	wire [4-1:0] node10596;
	wire [4-1:0] node10597;
	wire [4-1:0] node10598;
	wire [4-1:0] node10600;
	wire [4-1:0] node10603;
	wire [4-1:0] node10605;
	wire [4-1:0] node10608;
	wire [4-1:0] node10609;
	wire [4-1:0] node10611;
	wire [4-1:0] node10614;
	wire [4-1:0] node10616;
	wire [4-1:0] node10619;
	wire [4-1:0] node10620;
	wire [4-1:0] node10621;
	wire [4-1:0] node10623;
	wire [4-1:0] node10624;
	wire [4-1:0] node10627;
	wire [4-1:0] node10630;
	wire [4-1:0] node10632;
	wire [4-1:0] node10633;
	wire [4-1:0] node10636;
	wire [4-1:0] node10639;
	wire [4-1:0] node10640;
	wire [4-1:0] node10641;
	wire [4-1:0] node10642;
	wire [4-1:0] node10647;
	wire [4-1:0] node10648;
	wire [4-1:0] node10652;
	wire [4-1:0] node10653;
	wire [4-1:0] node10654;
	wire [4-1:0] node10655;
	wire [4-1:0] node10656;
	wire [4-1:0] node10657;
	wire [4-1:0] node10659;
	wire [4-1:0] node10662;
	wire [4-1:0] node10663;
	wire [4-1:0] node10667;
	wire [4-1:0] node10668;
	wire [4-1:0] node10671;
	wire [4-1:0] node10673;
	wire [4-1:0] node10676;
	wire [4-1:0] node10677;
	wire [4-1:0] node10678;
	wire [4-1:0] node10681;
	wire [4-1:0] node10684;
	wire [4-1:0] node10685;
	wire [4-1:0] node10688;
	wire [4-1:0] node10690;
	wire [4-1:0] node10693;
	wire [4-1:0] node10694;
	wire [4-1:0] node10695;
	wire [4-1:0] node10696;
	wire [4-1:0] node10699;
	wire [4-1:0] node10702;
	wire [4-1:0] node10704;
	wire [4-1:0] node10705;
	wire [4-1:0] node10708;
	wire [4-1:0] node10711;
	wire [4-1:0] node10712;
	wire [4-1:0] node10713;
	wire [4-1:0] node10715;
	wire [4-1:0] node10718;
	wire [4-1:0] node10719;
	wire [4-1:0] node10722;
	wire [4-1:0] node10725;
	wire [4-1:0] node10726;
	wire [4-1:0] node10729;
	wire [4-1:0] node10732;
	wire [4-1:0] node10733;
	wire [4-1:0] node10734;
	wire [4-1:0] node10735;
	wire [4-1:0] node10738;
	wire [4-1:0] node10739;
	wire [4-1:0] node10743;
	wire [4-1:0] node10744;
	wire [4-1:0] node10745;
	wire [4-1:0] node10749;
	wire [4-1:0] node10750;
	wire [4-1:0] node10754;
	wire [4-1:0] node10755;
	wire [4-1:0] node10756;
	wire [4-1:0] node10757;
	wire [4-1:0] node10758;
	wire [4-1:0] node10762;
	wire [4-1:0] node10765;
	wire [4-1:0] node10766;
	wire [4-1:0] node10767;
	wire [4-1:0] node10771;
	wire [4-1:0] node10774;
	wire [4-1:0] node10775;
	wire [4-1:0] node10776;
	wire [4-1:0] node10777;
	wire [4-1:0] node10781;
	wire [4-1:0] node10782;
	wire [4-1:0] node10786;
	wire [4-1:0] node10788;
	wire [4-1:0] node10789;
	wire [4-1:0] node10793;
	wire [4-1:0] node10794;
	wire [4-1:0] node10795;
	wire [4-1:0] node10796;
	wire [4-1:0] node10797;
	wire [4-1:0] node10798;
	wire [4-1:0] node10799;
	wire [4-1:0] node10803;
	wire [4-1:0] node10804;
	wire [4-1:0] node10805;
	wire [4-1:0] node10808;
	wire [4-1:0] node10812;
	wire [4-1:0] node10813;
	wire [4-1:0] node10816;
	wire [4-1:0] node10819;
	wire [4-1:0] node10820;
	wire [4-1:0] node10821;
	wire [4-1:0] node10822;
	wire [4-1:0] node10825;
	wire [4-1:0] node10828;
	wire [4-1:0] node10830;
	wire [4-1:0] node10833;
	wire [4-1:0] node10834;
	wire [4-1:0] node10835;
	wire [4-1:0] node10836;
	wire [4-1:0] node10839;
	wire [4-1:0] node10842;
	wire [4-1:0] node10843;
	wire [4-1:0] node10847;
	wire [4-1:0] node10848;
	wire [4-1:0] node10849;
	wire [4-1:0] node10852;
	wire [4-1:0] node10855;
	wire [4-1:0] node10856;
	wire [4-1:0] node10860;
	wire [4-1:0] node10861;
	wire [4-1:0] node10862;
	wire [4-1:0] node10863;
	wire [4-1:0] node10864;
	wire [4-1:0] node10867;
	wire [4-1:0] node10870;
	wire [4-1:0] node10871;
	wire [4-1:0] node10874;
	wire [4-1:0] node10877;
	wire [4-1:0] node10878;
	wire [4-1:0] node10879;
	wire [4-1:0] node10882;
	wire [4-1:0] node10885;
	wire [4-1:0] node10886;
	wire [4-1:0] node10887;
	wire [4-1:0] node10891;
	wire [4-1:0] node10892;
	wire [4-1:0] node10896;
	wire [4-1:0] node10897;
	wire [4-1:0] node10898;
	wire [4-1:0] node10899;
	wire [4-1:0] node10902;
	wire [4-1:0] node10905;
	wire [4-1:0] node10906;
	wire [4-1:0] node10907;
	wire [4-1:0] node10910;
	wire [4-1:0] node10913;
	wire [4-1:0] node10914;
	wire [4-1:0] node10917;
	wire [4-1:0] node10920;
	wire [4-1:0] node10921;
	wire [4-1:0] node10922;
	wire [4-1:0] node10925;
	wire [4-1:0] node10928;
	wire [4-1:0] node10930;
	wire [4-1:0] node10933;
	wire [4-1:0] node10934;
	wire [4-1:0] node10935;
	wire [4-1:0] node10936;
	wire [4-1:0] node10937;
	wire [4-1:0] node10939;
	wire [4-1:0] node10942;
	wire [4-1:0] node10943;
	wire [4-1:0] node10944;
	wire [4-1:0] node10947;
	wire [4-1:0] node10950;
	wire [4-1:0] node10951;
	wire [4-1:0] node10955;
	wire [4-1:0] node10956;
	wire [4-1:0] node10957;
	wire [4-1:0] node10961;
	wire [4-1:0] node10962;
	wire [4-1:0] node10964;
	wire [4-1:0] node10968;
	wire [4-1:0] node10969;
	wire [4-1:0] node10970;
	wire [4-1:0] node10971;
	wire [4-1:0] node10972;
	wire [4-1:0] node10976;
	wire [4-1:0] node10977;
	wire [4-1:0] node10981;
	wire [4-1:0] node10982;
	wire [4-1:0] node10983;
	wire [4-1:0] node10986;
	wire [4-1:0] node10990;
	wire [4-1:0] node10991;
	wire [4-1:0] node10992;
	wire [4-1:0] node10993;
	wire [4-1:0] node10996;
	wire [4-1:0] node10999;
	wire [4-1:0] node11000;
	wire [4-1:0] node11003;
	wire [4-1:0] node11006;
	wire [4-1:0] node11008;
	wire [4-1:0] node11010;
	wire [4-1:0] node11013;
	wire [4-1:0] node11014;
	wire [4-1:0] node11015;
	wire [4-1:0] node11016;
	wire [4-1:0] node11017;
	wire [4-1:0] node11018;
	wire [4-1:0] node11021;
	wire [4-1:0] node11025;
	wire [4-1:0] node11026;
	wire [4-1:0] node11027;
	wire [4-1:0] node11030;
	wire [4-1:0] node11033;
	wire [4-1:0] node11034;
	wire [4-1:0] node11037;
	wire [4-1:0] node11040;
	wire [4-1:0] node11041;
	wire [4-1:0] node11042;
	wire [4-1:0] node11043;
	wire [4-1:0] node11046;
	wire [4-1:0] node11049;
	wire [4-1:0] node11050;
	wire [4-1:0] node11054;
	wire [4-1:0] node11055;
	wire [4-1:0] node11057;
	wire [4-1:0] node11060;
	wire [4-1:0] node11061;
	wire [4-1:0] node11064;
	wire [4-1:0] node11067;
	wire [4-1:0] node11068;
	wire [4-1:0] node11069;
	wire [4-1:0] node11071;
	wire [4-1:0] node11072;
	wire [4-1:0] node11076;
	wire [4-1:0] node11078;
	wire [4-1:0] node11079;
	wire [4-1:0] node11083;
	wire [4-1:0] node11084;
	wire [4-1:0] node11087;
	wire [4-1:0] node11088;
	wire [4-1:0] node11091;
	wire [4-1:0] node11092;
	wire [4-1:0] node11096;
	wire [4-1:0] node11097;
	wire [4-1:0] node11098;
	wire [4-1:0] node11099;
	wire [4-1:0] node11100;
	wire [4-1:0] node11101;
	wire [4-1:0] node11102;
	wire [4-1:0] node11105;
	wire [4-1:0] node11107;
	wire [4-1:0] node11110;
	wire [4-1:0] node11111;
	wire [4-1:0] node11112;
	wire [4-1:0] node11115;
	wire [4-1:0] node11118;
	wire [4-1:0] node11119;
	wire [4-1:0] node11122;
	wire [4-1:0] node11125;
	wire [4-1:0] node11126;
	wire [4-1:0] node11127;
	wire [4-1:0] node11130;
	wire [4-1:0] node11132;
	wire [4-1:0] node11135;
	wire [4-1:0] node11136;
	wire [4-1:0] node11137;
	wire [4-1:0] node11140;
	wire [4-1:0] node11143;
	wire [4-1:0] node11144;
	wire [4-1:0] node11147;
	wire [4-1:0] node11150;
	wire [4-1:0] node11151;
	wire [4-1:0] node11152;
	wire [4-1:0] node11153;
	wire [4-1:0] node11156;
	wire [4-1:0] node11158;
	wire [4-1:0] node11161;
	wire [4-1:0] node11162;
	wire [4-1:0] node11163;
	wire [4-1:0] node11166;
	wire [4-1:0] node11169;
	wire [4-1:0] node11170;
	wire [4-1:0] node11173;
	wire [4-1:0] node11176;
	wire [4-1:0] node11177;
	wire [4-1:0] node11178;
	wire [4-1:0] node11181;
	wire [4-1:0] node11183;
	wire [4-1:0] node11186;
	wire [4-1:0] node11187;
	wire [4-1:0] node11188;
	wire [4-1:0] node11191;
	wire [4-1:0] node11194;
	wire [4-1:0] node11195;
	wire [4-1:0] node11196;
	wire [4-1:0] node11199;
	wire [4-1:0] node11203;
	wire [4-1:0] node11204;
	wire [4-1:0] node11205;
	wire [4-1:0] node11206;
	wire [4-1:0] node11207;
	wire [4-1:0] node11210;
	wire [4-1:0] node11211;
	wire [4-1:0] node11215;
	wire [4-1:0] node11216;
	wire [4-1:0] node11217;
	wire [4-1:0] node11220;
	wire [4-1:0] node11223;
	wire [4-1:0] node11224;
	wire [4-1:0] node11225;
	wire [4-1:0] node11229;
	wire [4-1:0] node11230;
	wire [4-1:0] node11233;
	wire [4-1:0] node11236;
	wire [4-1:0] node11237;
	wire [4-1:0] node11238;
	wire [4-1:0] node11239;
	wire [4-1:0] node11242;
	wire [4-1:0] node11244;
	wire [4-1:0] node11247;
	wire [4-1:0] node11249;
	wire [4-1:0] node11252;
	wire [4-1:0] node11253;
	wire [4-1:0] node11254;
	wire [4-1:0] node11257;
	wire [4-1:0] node11260;
	wire [4-1:0] node11261;
	wire [4-1:0] node11262;
	wire [4-1:0] node11267;
	wire [4-1:0] node11268;
	wire [4-1:0] node11269;
	wire [4-1:0] node11270;
	wire [4-1:0] node11271;
	wire [4-1:0] node11274;
	wire [4-1:0] node11277;
	wire [4-1:0] node11278;
	wire [4-1:0] node11281;
	wire [4-1:0] node11284;
	wire [4-1:0] node11285;
	wire [4-1:0] node11286;
	wire [4-1:0] node11290;
	wire [4-1:0] node11291;
	wire [4-1:0] node11294;
	wire [4-1:0] node11297;
	wire [4-1:0] node11298;
	wire [4-1:0] node11299;
	wire [4-1:0] node11301;
	wire [4-1:0] node11305;
	wire [4-1:0] node11306;
	wire [4-1:0] node11308;
	wire [4-1:0] node11311;
	wire [4-1:0] node11312;
	wire [4-1:0] node11316;
	wire [4-1:0] node11317;
	wire [4-1:0] node11318;
	wire [4-1:0] node11319;
	wire [4-1:0] node11320;
	wire [4-1:0] node11321;
	wire [4-1:0] node11322;
	wire [4-1:0] node11323;
	wire [4-1:0] node11326;
	wire [4-1:0] node11329;
	wire [4-1:0] node11330;
	wire [4-1:0] node11333;
	wire [4-1:0] node11336;
	wire [4-1:0] node11337;
	wire [4-1:0] node11339;
	wire [4-1:0] node11342;
	wire [4-1:0] node11343;
	wire [4-1:0] node11347;
	wire [4-1:0] node11348;
	wire [4-1:0] node11349;
	wire [4-1:0] node11352;
	wire [4-1:0] node11353;
	wire [4-1:0] node11356;
	wire [4-1:0] node11359;
	wire [4-1:0] node11360;
	wire [4-1:0] node11361;
	wire [4-1:0] node11365;
	wire [4-1:0] node11368;
	wire [4-1:0] node11369;
	wire [4-1:0] node11370;
	wire [4-1:0] node11371;
	wire [4-1:0] node11372;
	wire [4-1:0] node11377;
	wire [4-1:0] node11378;
	wire [4-1:0] node11379;
	wire [4-1:0] node11382;
	wire [4-1:0] node11385;
	wire [4-1:0] node11387;
	wire [4-1:0] node11390;
	wire [4-1:0] node11391;
	wire [4-1:0] node11394;
	wire [4-1:0] node11395;
	wire [4-1:0] node11399;
	wire [4-1:0] node11400;
	wire [4-1:0] node11401;
	wire [4-1:0] node11402;
	wire [4-1:0] node11403;
	wire [4-1:0] node11406;
	wire [4-1:0] node11409;
	wire [4-1:0] node11410;
	wire [4-1:0] node11412;
	wire [4-1:0] node11415;
	wire [4-1:0] node11416;
	wire [4-1:0] node11419;
	wire [4-1:0] node11422;
	wire [4-1:0] node11423;
	wire [4-1:0] node11424;
	wire [4-1:0] node11425;
	wire [4-1:0] node11428;
	wire [4-1:0] node11431;
	wire [4-1:0] node11432;
	wire [4-1:0] node11436;
	wire [4-1:0] node11437;
	wire [4-1:0] node11438;
	wire [4-1:0] node11441;
	wire [4-1:0] node11444;
	wire [4-1:0] node11447;
	wire [4-1:0] node11448;
	wire [4-1:0] node11449;
	wire [4-1:0] node11450;
	wire [4-1:0] node11453;
	wire [4-1:0] node11455;
	wire [4-1:0] node11458;
	wire [4-1:0] node11459;
	wire [4-1:0] node11460;
	wire [4-1:0] node11463;
	wire [4-1:0] node11466;
	wire [4-1:0] node11467;
	wire [4-1:0] node11470;
	wire [4-1:0] node11473;
	wire [4-1:0] node11474;
	wire [4-1:0] node11475;
	wire [4-1:0] node11478;
	wire [4-1:0] node11481;
	wire [4-1:0] node11482;
	wire [4-1:0] node11483;
	wire [4-1:0] node11487;
	wire [4-1:0] node11488;
	wire [4-1:0] node11491;
	wire [4-1:0] node11494;
	wire [4-1:0] node11495;
	wire [4-1:0] node11496;
	wire [4-1:0] node11497;
	wire [4-1:0] node11498;
	wire [4-1:0] node11499;
	wire [4-1:0] node11503;
	wire [4-1:0] node11504;
	wire [4-1:0] node11507;
	wire [4-1:0] node11510;
	wire [4-1:0] node11511;
	wire [4-1:0] node11512;
	wire [4-1:0] node11515;
	wire [4-1:0] node11518;
	wire [4-1:0] node11519;
	wire [4-1:0] node11522;
	wire [4-1:0] node11525;
	wire [4-1:0] node11526;
	wire [4-1:0] node11527;
	wire [4-1:0] node11528;
	wire [4-1:0] node11532;
	wire [4-1:0] node11533;
	wire [4-1:0] node11537;
	wire [4-1:0] node11538;
	wire [4-1:0] node11539;
	wire [4-1:0] node11543;
	wire [4-1:0] node11544;
	wire [4-1:0] node11548;
	wire [4-1:0] node11549;
	wire [4-1:0] node11550;
	wire [4-1:0] node11551;
	wire [4-1:0] node11552;
	wire [4-1:0] node11555;
	wire [4-1:0] node11558;
	wire [4-1:0] node11561;
	wire [4-1:0] node11562;
	wire [4-1:0] node11563;
	wire [4-1:0] node11567;
	wire [4-1:0] node11568;
	wire [4-1:0] node11572;
	wire [4-1:0] node11573;
	wire [4-1:0] node11574;
	wire [4-1:0] node11575;
	wire [4-1:0] node11578;
	wire [4-1:0] node11581;
	wire [4-1:0] node11582;
	wire [4-1:0] node11585;
	wire [4-1:0] node11588;
	wire [4-1:0] node11589;
	wire [4-1:0] node11590;
	wire [4-1:0] node11593;
	wire [4-1:0] node11596;
	wire [4-1:0] node11597;
	wire [4-1:0] node11599;
	wire [4-1:0] node11602;
	wire [4-1:0] node11603;
	wire [4-1:0] node11607;
	wire [4-1:0] node11608;
	wire [4-1:0] node11609;
	wire [4-1:0] node11610;
	wire [4-1:0] node11611;
	wire [4-1:0] node11612;
	wire [4-1:0] node11613;
	wire [4-1:0] node11614;
	wire [4-1:0] node11616;
	wire [4-1:0] node11619;
	wire [4-1:0] node11621;
	wire [4-1:0] node11624;
	wire [4-1:0] node11625;
	wire [4-1:0] node11627;
	wire [4-1:0] node11630;
	wire [4-1:0] node11633;
	wire [4-1:0] node11634;
	wire [4-1:0] node11635;
	wire [4-1:0] node11636;
	wire [4-1:0] node11638;
	wire [4-1:0] node11641;
	wire [4-1:0] node11643;
	wire [4-1:0] node11646;
	wire [4-1:0] node11647;
	wire [4-1:0] node11651;
	wire [4-1:0] node11652;
	wire [4-1:0] node11653;
	wire [4-1:0] node11656;
	wire [4-1:0] node11659;
	wire [4-1:0] node11661;
	wire [4-1:0] node11664;
	wire [4-1:0] node11665;
	wire [4-1:0] node11666;
	wire [4-1:0] node11667;
	wire [4-1:0] node11669;
	wire [4-1:0] node11672;
	wire [4-1:0] node11674;
	wire [4-1:0] node11677;
	wire [4-1:0] node11678;
	wire [4-1:0] node11680;
	wire [4-1:0] node11683;
	wire [4-1:0] node11685;
	wire [4-1:0] node11688;
	wire [4-1:0] node11689;
	wire [4-1:0] node11690;
	wire [4-1:0] node11691;
	wire [4-1:0] node11693;
	wire [4-1:0] node11697;
	wire [4-1:0] node11699;
	wire [4-1:0] node11702;
	wire [4-1:0] node11703;
	wire [4-1:0] node11706;
	wire [4-1:0] node11708;
	wire [4-1:0] node11711;
	wire [4-1:0] node11712;
	wire [4-1:0] node11713;
	wire [4-1:0] node11714;
	wire [4-1:0] node11715;
	wire [4-1:0] node11717;
	wire [4-1:0] node11720;
	wire [4-1:0] node11722;
	wire [4-1:0] node11725;
	wire [4-1:0] node11726;
	wire [4-1:0] node11730;
	wire [4-1:0] node11731;
	wire [4-1:0] node11733;
	wire [4-1:0] node11734;
	wire [4-1:0] node11736;
	wire [4-1:0] node11739;
	wire [4-1:0] node11742;
	wire [4-1:0] node11743;
	wire [4-1:0] node11744;
	wire [4-1:0] node11745;
	wire [4-1:0] node11750;
	wire [4-1:0] node11751;
	wire [4-1:0] node11752;
	wire [4-1:0] node11756;
	wire [4-1:0] node11757;
	wire [4-1:0] node11761;
	wire [4-1:0] node11762;
	wire [4-1:0] node11763;
	wire [4-1:0] node11764;
	wire [4-1:0] node11765;
	wire [4-1:0] node11769;
	wire [4-1:0] node11770;
	wire [4-1:0] node11774;
	wire [4-1:0] node11775;
	wire [4-1:0] node11776;
	wire [4-1:0] node11780;
	wire [4-1:0] node11781;
	wire [4-1:0] node11785;
	wire [4-1:0] node11786;
	wire [4-1:0] node11787;
	wire [4-1:0] node11788;
	wire [4-1:0] node11789;
	wire [4-1:0] node11794;
	wire [4-1:0] node11795;
	wire [4-1:0] node11799;
	wire [4-1:0] node11800;
	wire [4-1:0] node11801;
	wire [4-1:0] node11802;
	wire [4-1:0] node11806;
	wire [4-1:0] node11809;
	wire [4-1:0] node11811;
	wire [4-1:0] node11814;
	wire [4-1:0] node11815;
	wire [4-1:0] node11816;
	wire [4-1:0] node11817;
	wire [4-1:0] node11818;
	wire [4-1:0] node11820;
	wire [4-1:0] node11822;
	wire [4-1:0] node11824;
	wire [4-1:0] node11827;
	wire [4-1:0] node11828;
	wire [4-1:0] node11829;
	wire [4-1:0] node11831;
	wire [4-1:0] node11834;
	wire [4-1:0] node11836;
	wire [4-1:0] node11839;
	wire [4-1:0] node11840;
	wire [4-1:0] node11842;
	wire [4-1:0] node11845;
	wire [4-1:0] node11848;
	wire [4-1:0] node11849;
	wire [4-1:0] node11850;
	wire [4-1:0] node11851;
	wire [4-1:0] node11854;
	wire [4-1:0] node11858;
	wire [4-1:0] node11859;
	wire [4-1:0] node11860;
	wire [4-1:0] node11862;
	wire [4-1:0] node11865;
	wire [4-1:0] node11867;
	wire [4-1:0] node11870;
	wire [4-1:0] node11871;
	wire [4-1:0] node11873;
	wire [4-1:0] node11876;
	wire [4-1:0] node11879;
	wire [4-1:0] node11880;
	wire [4-1:0] node11881;
	wire [4-1:0] node11882;
	wire [4-1:0] node11883;
	wire [4-1:0] node11886;
	wire [4-1:0] node11888;
	wire [4-1:0] node11891;
	wire [4-1:0] node11892;
	wire [4-1:0] node11895;
	wire [4-1:0] node11898;
	wire [4-1:0] node11899;
	wire [4-1:0] node11900;
	wire [4-1:0] node11903;
	wire [4-1:0] node11906;
	wire [4-1:0] node11907;
	wire [4-1:0] node11909;
	wire [4-1:0] node11912;
	wire [4-1:0] node11913;
	wire [4-1:0] node11916;
	wire [4-1:0] node11919;
	wire [4-1:0] node11920;
	wire [4-1:0] node11921;
	wire [4-1:0] node11923;
	wire [4-1:0] node11924;
	wire [4-1:0] node11927;
	wire [4-1:0] node11930;
	wire [4-1:0] node11931;
	wire [4-1:0] node11934;
	wire [4-1:0] node11936;
	wire [4-1:0] node11939;
	wire [4-1:0] node11940;
	wire [4-1:0] node11941;
	wire [4-1:0] node11943;
	wire [4-1:0] node11946;
	wire [4-1:0] node11949;
	wire [4-1:0] node11950;
	wire [4-1:0] node11952;
	wire [4-1:0] node11955;
	wire [4-1:0] node11957;
	wire [4-1:0] node11960;
	wire [4-1:0] node11961;
	wire [4-1:0] node11962;
	wire [4-1:0] node11963;
	wire [4-1:0] node11964;
	wire [4-1:0] node11965;
	wire [4-1:0] node11968;
	wire [4-1:0] node11971;
	wire [4-1:0] node11973;
	wire [4-1:0] node11974;
	wire [4-1:0] node11977;
	wire [4-1:0] node11980;
	wire [4-1:0] node11981;
	wire [4-1:0] node11982;
	wire [4-1:0] node11984;
	wire [4-1:0] node11987;
	wire [4-1:0] node11989;
	wire [4-1:0] node11992;
	wire [4-1:0] node11994;
	wire [4-1:0] node11995;
	wire [4-1:0] node11998;
	wire [4-1:0] node12001;
	wire [4-1:0] node12002;
	wire [4-1:0] node12003;
	wire [4-1:0] node12004;
	wire [4-1:0] node12007;
	wire [4-1:0] node12010;
	wire [4-1:0] node12011;
	wire [4-1:0] node12015;
	wire [4-1:0] node12016;
	wire [4-1:0] node12017;
	wire [4-1:0] node12020;
	wire [4-1:0] node12023;
	wire [4-1:0] node12024;
	wire [4-1:0] node12027;
	wire [4-1:0] node12030;
	wire [4-1:0] node12031;
	wire [4-1:0] node12032;
	wire [4-1:0] node12033;
	wire [4-1:0] node12035;
	wire [4-1:0] node12038;
	wire [4-1:0] node12040;
	wire [4-1:0] node12043;
	wire [4-1:0] node12044;
	wire [4-1:0] node12046;
	wire [4-1:0] node12049;
	wire [4-1:0] node12050;
	wire [4-1:0] node12052;
	wire [4-1:0] node12056;
	wire [4-1:0] node12057;
	wire [4-1:0] node12058;
	wire [4-1:0] node12060;
	wire [4-1:0] node12062;
	wire [4-1:0] node12065;
	wire [4-1:0] node12066;
	wire [4-1:0] node12069;
	wire [4-1:0] node12072;
	wire [4-1:0] node12073;
	wire [4-1:0] node12074;
	wire [4-1:0] node12078;
	wire [4-1:0] node12079;
	wire [4-1:0] node12082;
	wire [4-1:0] node12084;
	wire [4-1:0] node12087;
	wire [4-1:0] node12088;
	wire [4-1:0] node12089;
	wire [4-1:0] node12090;
	wire [4-1:0] node12091;
	wire [4-1:0] node12092;
	wire [4-1:0] node12094;
	wire [4-1:0] node12097;
	wire [4-1:0] node12099;
	wire [4-1:0] node12102;
	wire [4-1:0] node12103;
	wire [4-1:0] node12105;
	wire [4-1:0] node12108;
	wire [4-1:0] node12110;
	wire [4-1:0] node12113;
	wire [4-1:0] node12114;
	wire [4-1:0] node12115;
	wire [4-1:0] node12116;
	wire [4-1:0] node12118;
	wire [4-1:0] node12121;
	wire [4-1:0] node12123;
	wire [4-1:0] node12126;
	wire [4-1:0] node12127;
	wire [4-1:0] node12129;
	wire [4-1:0] node12132;
	wire [4-1:0] node12134;
	wire [4-1:0] node12137;
	wire [4-1:0] node12138;
	wire [4-1:0] node12139;
	wire [4-1:0] node12140;
	wire [4-1:0] node12141;
	wire [4-1:0] node12144;
	wire [4-1:0] node12148;
	wire [4-1:0] node12150;
	wire [4-1:0] node12153;
	wire [4-1:0] node12154;
	wire [4-1:0] node12155;
	wire [4-1:0] node12158;
	wire [4-1:0] node12161;
	wire [4-1:0] node12162;
	wire [4-1:0] node12166;
	wire [4-1:0] node12167;
	wire [4-1:0] node12168;
	wire [4-1:0] node12169;
	wire [4-1:0] node12171;
	wire [4-1:0] node12174;
	wire [4-1:0] node12176;
	wire [4-1:0] node12179;
	wire [4-1:0] node12180;
	wire [4-1:0] node12182;
	wire [4-1:0] node12185;
	wire [4-1:0] node12187;
	wire [4-1:0] node12190;
	wire [4-1:0] node12191;
	wire [4-1:0] node12192;
	wire [4-1:0] node12193;
	wire [4-1:0] node12194;
	wire [4-1:0] node12195;
	wire [4-1:0] node12198;
	wire [4-1:0] node12201;
	wire [4-1:0] node12202;
	wire [4-1:0] node12206;
	wire [4-1:0] node12207;
	wire [4-1:0] node12208;
	wire [4-1:0] node12213;
	wire [4-1:0] node12214;
	wire [4-1:0] node12215;
	wire [4-1:0] node12218;
	wire [4-1:0] node12221;
	wire [4-1:0] node12222;
	wire [4-1:0] node12223;
	wire [4-1:0] node12228;
	wire [4-1:0] node12229;
	wire [4-1:0] node12230;
	wire [4-1:0] node12231;
	wire [4-1:0] node12234;
	wire [4-1:0] node12237;
	wire [4-1:0] node12238;
	wire [4-1:0] node12241;
	wire [4-1:0] node12244;
	wire [4-1:0] node12245;
	wire [4-1:0] node12246;
	wire [4-1:0] node12247;
	wire [4-1:0] node12250;
	wire [4-1:0] node12253;
	wire [4-1:0] node12254;
	wire [4-1:0] node12257;
	wire [4-1:0] node12260;
	wire [4-1:0] node12262;
	wire [4-1:0] node12265;
	wire [4-1:0] node12266;
	wire [4-1:0] node12267;
	wire [4-1:0] node12268;
	wire [4-1:0] node12269;
	wire [4-1:0] node12272;
	wire [4-1:0] node12275;
	wire [4-1:0] node12276;
	wire [4-1:0] node12277;
	wire [4-1:0] node12278;
	wire [4-1:0] node12281;
	wire [4-1:0] node12284;
	wire [4-1:0] node12285;
	wire [4-1:0] node12286;
	wire [4-1:0] node12289;
	wire [4-1:0] node12292;
	wire [4-1:0] node12293;
	wire [4-1:0] node12296;
	wire [4-1:0] node12299;
	wire [4-1:0] node12300;
	wire [4-1:0] node12303;
	wire [4-1:0] node12306;
	wire [4-1:0] node12307;
	wire [4-1:0] node12308;
	wire [4-1:0] node12309;
	wire [4-1:0] node12310;
	wire [4-1:0] node12314;
	wire [4-1:0] node12315;
	wire [4-1:0] node12316;
	wire [4-1:0] node12320;
	wire [4-1:0] node12321;
	wire [4-1:0] node12325;
	wire [4-1:0] node12326;
	wire [4-1:0] node12327;
	wire [4-1:0] node12328;
	wire [4-1:0] node12331;
	wire [4-1:0] node12334;
	wire [4-1:0] node12336;
	wire [4-1:0] node12339;
	wire [4-1:0] node12340;
	wire [4-1:0] node12341;
	wire [4-1:0] node12344;
	wire [4-1:0] node12347;
	wire [4-1:0] node12349;
	wire [4-1:0] node12352;
	wire [4-1:0] node12353;
	wire [4-1:0] node12354;
	wire [4-1:0] node12355;
	wire [4-1:0] node12356;
	wire [4-1:0] node12359;
	wire [4-1:0] node12362;
	wire [4-1:0] node12364;
	wire [4-1:0] node12367;
	wire [4-1:0] node12368;
	wire [4-1:0] node12372;
	wire [4-1:0] node12373;
	wire [4-1:0] node12376;
	wire [4-1:0] node12379;
	wire [4-1:0] node12380;
	wire [4-1:0] node12381;
	wire [4-1:0] node12382;
	wire [4-1:0] node12383;
	wire [4-1:0] node12387;
	wire [4-1:0] node12388;
	wire [4-1:0] node12392;
	wire [4-1:0] node12393;
	wire [4-1:0] node12394;
	wire [4-1:0] node12398;
	wire [4-1:0] node12399;
	wire [4-1:0] node12403;
	wire [4-1:0] node12404;
	wire [4-1:0] node12405;
	wire [4-1:0] node12406;
	wire [4-1:0] node12407;
	wire [4-1:0] node12410;
	wire [4-1:0] node12413;
	wire [4-1:0] node12414;
	wire [4-1:0] node12418;
	wire [4-1:0] node12419;
	wire [4-1:0] node12422;
	wire [4-1:0] node12425;
	wire [4-1:0] node12426;
	wire [4-1:0] node12427;
	wire [4-1:0] node12428;
	wire [4-1:0] node12431;
	wire [4-1:0] node12434;
	wire [4-1:0] node12435;
	wire [4-1:0] node12436;
	wire [4-1:0] node12440;
	wire [4-1:0] node12441;
	wire [4-1:0] node12445;
	wire [4-1:0] node12446;
	wire [4-1:0] node12449;
	wire [4-1:0] node12452;
	wire [4-1:0] node12453;
	wire [4-1:0] node12454;
	wire [4-1:0] node12455;
	wire [4-1:0] node12456;
	wire [4-1:0] node12457;
	wire [4-1:0] node12458;
	wire [4-1:0] node12459;
	wire [4-1:0] node12460;
	wire [4-1:0] node12461;
	wire [4-1:0] node12464;
	wire [4-1:0] node12467;
	wire [4-1:0] node12468;
	wire [4-1:0] node12470;
	wire [4-1:0] node12471;
	wire [4-1:0] node12474;
	wire [4-1:0] node12477;
	wire [4-1:0] node12478;
	wire [4-1:0] node12481;
	wire [4-1:0] node12484;
	wire [4-1:0] node12485;
	wire [4-1:0] node12486;
	wire [4-1:0] node12488;
	wire [4-1:0] node12489;
	wire [4-1:0] node12493;
	wire [4-1:0] node12495;
	wire [4-1:0] node12498;
	wire [4-1:0] node12499;
	wire [4-1:0] node12501;
	wire [4-1:0] node12504;
	wire [4-1:0] node12505;
	wire [4-1:0] node12508;
	wire [4-1:0] node12511;
	wire [4-1:0] node12512;
	wire [4-1:0] node12513;
	wire [4-1:0] node12514;
	wire [4-1:0] node12515;
	wire [4-1:0] node12518;
	wire [4-1:0] node12521;
	wire [4-1:0] node12522;
	wire [4-1:0] node12525;
	wire [4-1:0] node12528;
	wire [4-1:0] node12529;
	wire [4-1:0] node12530;
	wire [4-1:0] node12533;
	wire [4-1:0] node12536;
	wire [4-1:0] node12537;
	wire [4-1:0] node12538;
	wire [4-1:0] node12541;
	wire [4-1:0] node12545;
	wire [4-1:0] node12546;
	wire [4-1:0] node12547;
	wire [4-1:0] node12548;
	wire [4-1:0] node12551;
	wire [4-1:0] node12554;
	wire [4-1:0] node12555;
	wire [4-1:0] node12558;
	wire [4-1:0] node12561;
	wire [4-1:0] node12562;
	wire [4-1:0] node12564;
	wire [4-1:0] node12567;
	wire [4-1:0] node12568;
	wire [4-1:0] node12571;
	wire [4-1:0] node12574;
	wire [4-1:0] node12575;
	wire [4-1:0] node12576;
	wire [4-1:0] node12577;
	wire [4-1:0] node12578;
	wire [4-1:0] node12580;
	wire [4-1:0] node12583;
	wire [4-1:0] node12585;
	wire [4-1:0] node12588;
	wire [4-1:0] node12589;
	wire [4-1:0] node12590;
	wire [4-1:0] node12594;
	wire [4-1:0] node12596;
	wire [4-1:0] node12599;
	wire [4-1:0] node12600;
	wire [4-1:0] node12601;
	wire [4-1:0] node12602;
	wire [4-1:0] node12603;
	wire [4-1:0] node12606;
	wire [4-1:0] node12610;
	wire [4-1:0] node12611;
	wire [4-1:0] node12613;
	wire [4-1:0] node12616;
	wire [4-1:0] node12617;
	wire [4-1:0] node12620;
	wire [4-1:0] node12623;
	wire [4-1:0] node12624;
	wire [4-1:0] node12626;
	wire [4-1:0] node12627;
	wire [4-1:0] node12630;
	wire [4-1:0] node12634;
	wire [4-1:0] node12635;
	wire [4-1:0] node12636;
	wire [4-1:0] node12637;
	wire [4-1:0] node12640;
	wire [4-1:0] node12642;
	wire [4-1:0] node12645;
	wire [4-1:0] node12646;
	wire [4-1:0] node12648;
	wire [4-1:0] node12651;
	wire [4-1:0] node12653;
	wire [4-1:0] node12656;
	wire [4-1:0] node12657;
	wire [4-1:0] node12659;
	wire [4-1:0] node12661;
	wire [4-1:0] node12664;
	wire [4-1:0] node12665;
	wire [4-1:0] node12667;
	wire [4-1:0] node12670;
	wire [4-1:0] node12672;
	wire [4-1:0] node12675;
	wire [4-1:0] node12676;
	wire [4-1:0] node12677;
	wire [4-1:0] node12678;
	wire [4-1:0] node12679;
	wire [4-1:0] node12682;
	wire [4-1:0] node12685;
	wire [4-1:0] node12686;
	wire [4-1:0] node12687;
	wire [4-1:0] node12690;
	wire [4-1:0] node12693;
	wire [4-1:0] node12694;
	wire [4-1:0] node12695;
	wire [4-1:0] node12696;
	wire [4-1:0] node12700;
	wire [4-1:0] node12702;
	wire [4-1:0] node12705;
	wire [4-1:0] node12706;
	wire [4-1:0] node12708;
	wire [4-1:0] node12711;
	wire [4-1:0] node12712;
	wire [4-1:0] node12716;
	wire [4-1:0] node12717;
	wire [4-1:0] node12718;
	wire [4-1:0] node12719;
	wire [4-1:0] node12722;
	wire [4-1:0] node12725;
	wire [4-1:0] node12726;
	wire [4-1:0] node12729;
	wire [4-1:0] node12732;
	wire [4-1:0] node12733;
	wire [4-1:0] node12734;
	wire [4-1:0] node12737;
	wire [4-1:0] node12740;
	wire [4-1:0] node12741;
	wire [4-1:0] node12744;
	wire [4-1:0] node12747;
	wire [4-1:0] node12748;
	wire [4-1:0] node12749;
	wire [4-1:0] node12750;
	wire [4-1:0] node12751;
	wire [4-1:0] node12752;
	wire [4-1:0] node12755;
	wire [4-1:0] node12756;
	wire [4-1:0] node12760;
	wire [4-1:0] node12761;
	wire [4-1:0] node12764;
	wire [4-1:0] node12767;
	wire [4-1:0] node12768;
	wire [4-1:0] node12770;
	wire [4-1:0] node12771;
	wire [4-1:0] node12774;
	wire [4-1:0] node12777;
	wire [4-1:0] node12778;
	wire [4-1:0] node12781;
	wire [4-1:0] node12784;
	wire [4-1:0] node12785;
	wire [4-1:0] node12786;
	wire [4-1:0] node12789;
	wire [4-1:0] node12792;
	wire [4-1:0] node12793;
	wire [4-1:0] node12796;
	wire [4-1:0] node12799;
	wire [4-1:0] node12800;
	wire [4-1:0] node12801;
	wire [4-1:0] node12804;
	wire [4-1:0] node12807;
	wire [4-1:0] node12808;
	wire [4-1:0] node12809;
	wire [4-1:0] node12810;
	wire [4-1:0] node12811;
	wire [4-1:0] node12814;
	wire [4-1:0] node12818;
	wire [4-1:0] node12820;
	wire [4-1:0] node12823;
	wire [4-1:0] node12824;
	wire [4-1:0] node12825;
	wire [4-1:0] node12828;
	wire [4-1:0] node12831;
	wire [4-1:0] node12832;
	wire [4-1:0] node12834;
	wire [4-1:0] node12838;
	wire [4-1:0] node12839;
	wire [4-1:0] node12840;
	wire [4-1:0] node12841;
	wire [4-1:0] node12842;
	wire [4-1:0] node12843;
	wire [4-1:0] node12844;
	wire [4-1:0] node12845;
	wire [4-1:0] node12848;
	wire [4-1:0] node12851;
	wire [4-1:0] node12852;
	wire [4-1:0] node12855;
	wire [4-1:0] node12858;
	wire [4-1:0] node12859;
	wire [4-1:0] node12860;
	wire [4-1:0] node12861;
	wire [4-1:0] node12865;
	wire [4-1:0] node12866;
	wire [4-1:0] node12870;
	wire [4-1:0] node12871;
	wire [4-1:0] node12874;
	wire [4-1:0] node12877;
	wire [4-1:0] node12878;
	wire [4-1:0] node12879;
	wire [4-1:0] node12881;
	wire [4-1:0] node12884;
	wire [4-1:0] node12885;
	wire [4-1:0] node12888;
	wire [4-1:0] node12891;
	wire [4-1:0] node12892;
	wire [4-1:0] node12893;
	wire [4-1:0] node12896;
	wire [4-1:0] node12899;
	wire [4-1:0] node12900;
	wire [4-1:0] node12903;
	wire [4-1:0] node12906;
	wire [4-1:0] node12907;
	wire [4-1:0] node12908;
	wire [4-1:0] node12909;
	wire [4-1:0] node12910;
	wire [4-1:0] node12911;
	wire [4-1:0] node12914;
	wire [4-1:0] node12917;
	wire [4-1:0] node12920;
	wire [4-1:0] node12923;
	wire [4-1:0] node12924;
	wire [4-1:0] node12926;
	wire [4-1:0] node12927;
	wire [4-1:0] node12930;
	wire [4-1:0] node12933;
	wire [4-1:0] node12935;
	wire [4-1:0] node12937;
	wire [4-1:0] node12940;
	wire [4-1:0] node12941;
	wire [4-1:0] node12942;
	wire [4-1:0] node12944;
	wire [4-1:0] node12945;
	wire [4-1:0] node12948;
	wire [4-1:0] node12951;
	wire [4-1:0] node12952;
	wire [4-1:0] node12953;
	wire [4-1:0] node12956;
	wire [4-1:0] node12960;
	wire [4-1:0] node12961;
	wire [4-1:0] node12962;
	wire [4-1:0] node12964;
	wire [4-1:0] node12967;
	wire [4-1:0] node12968;
	wire [4-1:0] node12971;
	wire [4-1:0] node12974;
	wire [4-1:0] node12975;
	wire [4-1:0] node12976;
	wire [4-1:0] node12981;
	wire [4-1:0] node12982;
	wire [4-1:0] node12983;
	wire [4-1:0] node12984;
	wire [4-1:0] node12985;
	wire [4-1:0] node12988;
	wire [4-1:0] node12990;
	wire [4-1:0] node12993;
	wire [4-1:0] node12994;
	wire [4-1:0] node12996;
	wire [4-1:0] node12999;
	wire [4-1:0] node13001;
	wire [4-1:0] node13004;
	wire [4-1:0] node13005;
	wire [4-1:0] node13006;
	wire [4-1:0] node13007;
	wire [4-1:0] node13010;
	wire [4-1:0] node13013;
	wire [4-1:0] node13015;
	wire [4-1:0] node13018;
	wire [4-1:0] node13019;
	wire [4-1:0] node13020;
	wire [4-1:0] node13021;
	wire [4-1:0] node13024;
	wire [4-1:0] node13027;
	wire [4-1:0] node13029;
	wire [4-1:0] node13032;
	wire [4-1:0] node13033;
	wire [4-1:0] node13037;
	wire [4-1:0] node13038;
	wire [4-1:0] node13039;
	wire [4-1:0] node13041;
	wire [4-1:0] node13044;
	wire [4-1:0] node13045;
	wire [4-1:0] node13047;
	wire [4-1:0] node13050;
	wire [4-1:0] node13052;
	wire [4-1:0] node13055;
	wire [4-1:0] node13056;
	wire [4-1:0] node13057;
	wire [4-1:0] node13059;
	wire [4-1:0] node13062;
	wire [4-1:0] node13063;
	wire [4-1:0] node13064;
	wire [4-1:0] node13067;
	wire [4-1:0] node13070;
	wire [4-1:0] node13072;
	wire [4-1:0] node13075;
	wire [4-1:0] node13076;
	wire [4-1:0] node13077;
	wire [4-1:0] node13080;
	wire [4-1:0] node13083;
	wire [4-1:0] node13084;
	wire [4-1:0] node13085;
	wire [4-1:0] node13088;
	wire [4-1:0] node13092;
	wire [4-1:0] node13093;
	wire [4-1:0] node13094;
	wire [4-1:0] node13095;
	wire [4-1:0] node13096;
	wire [4-1:0] node13097;
	wire [4-1:0] node13098;
	wire [4-1:0] node13099;
	wire [4-1:0] node13102;
	wire [4-1:0] node13106;
	wire [4-1:0] node13108;
	wire [4-1:0] node13111;
	wire [4-1:0] node13112;
	wire [4-1:0] node13114;
	wire [4-1:0] node13115;
	wire [4-1:0] node13118;
	wire [4-1:0] node13121;
	wire [4-1:0] node13122;
	wire [4-1:0] node13125;
	wire [4-1:0] node13128;
	wire [4-1:0] node13129;
	wire [4-1:0] node13130;
	wire [4-1:0] node13131;
	wire [4-1:0] node13134;
	wire [4-1:0] node13135;
	wire [4-1:0] node13138;
	wire [4-1:0] node13141;
	wire [4-1:0] node13142;
	wire [4-1:0] node13145;
	wire [4-1:0] node13148;
	wire [4-1:0] node13149;
	wire [4-1:0] node13151;
	wire [4-1:0] node13152;
	wire [4-1:0] node13155;
	wire [4-1:0] node13158;
	wire [4-1:0] node13159;
	wire [4-1:0] node13161;
	wire [4-1:0] node13164;
	wire [4-1:0] node13165;
	wire [4-1:0] node13168;
	wire [4-1:0] node13171;
	wire [4-1:0] node13172;
	wire [4-1:0] node13173;
	wire [4-1:0] node13174;
	wire [4-1:0] node13175;
	wire [4-1:0] node13176;
	wire [4-1:0] node13179;
	wire [4-1:0] node13182;
	wire [4-1:0] node13183;
	wire [4-1:0] node13187;
	wire [4-1:0] node13188;
	wire [4-1:0] node13189;
	wire [4-1:0] node13192;
	wire [4-1:0] node13195;
	wire [4-1:0] node13197;
	wire [4-1:0] node13200;
	wire [4-1:0] node13201;
	wire [4-1:0] node13202;
	wire [4-1:0] node13205;
	wire [4-1:0] node13207;
	wire [4-1:0] node13210;
	wire [4-1:0] node13211;
	wire [4-1:0] node13212;
	wire [4-1:0] node13215;
	wire [4-1:0] node13218;
	wire [4-1:0] node13220;
	wire [4-1:0] node13223;
	wire [4-1:0] node13224;
	wire [4-1:0] node13225;
	wire [4-1:0] node13226;
	wire [4-1:0] node13229;
	wire [4-1:0] node13232;
	wire [4-1:0] node13233;
	wire [4-1:0] node13236;
	wire [4-1:0] node13239;
	wire [4-1:0] node13240;
	wire [4-1:0] node13241;
	wire [4-1:0] node13245;
	wire [4-1:0] node13246;
	wire [4-1:0] node13248;
	wire [4-1:0] node13251;
	wire [4-1:0] node13254;
	wire [4-1:0] node13255;
	wire [4-1:0] node13256;
	wire [4-1:0] node13257;
	wire [4-1:0] node13258;
	wire [4-1:0] node13259;
	wire [4-1:0] node13260;
	wire [4-1:0] node13265;
	wire [4-1:0] node13267;
	wire [4-1:0] node13268;
	wire [4-1:0] node13272;
	wire [4-1:0] node13273;
	wire [4-1:0] node13274;
	wire [4-1:0] node13277;
	wire [4-1:0] node13279;
	wire [4-1:0] node13282;
	wire [4-1:0] node13283;
	wire [4-1:0] node13286;
	wire [4-1:0] node13289;
	wire [4-1:0] node13290;
	wire [4-1:0] node13291;
	wire [4-1:0] node13292;
	wire [4-1:0] node13293;
	wire [4-1:0] node13296;
	wire [4-1:0] node13299;
	wire [4-1:0] node13300;
	wire [4-1:0] node13303;
	wire [4-1:0] node13306;
	wire [4-1:0] node13307;
	wire [4-1:0] node13311;
	wire [4-1:0] node13312;
	wire [4-1:0] node13313;
	wire [4-1:0] node13314;
	wire [4-1:0] node13317;
	wire [4-1:0] node13321;
	wire [4-1:0] node13322;
	wire [4-1:0] node13323;
	wire [4-1:0] node13326;
	wire [4-1:0] node13330;
	wire [4-1:0] node13331;
	wire [4-1:0] node13332;
	wire [4-1:0] node13333;
	wire [4-1:0] node13334;
	wire [4-1:0] node13335;
	wire [4-1:0] node13338;
	wire [4-1:0] node13342;
	wire [4-1:0] node13343;
	wire [4-1:0] node13345;
	wire [4-1:0] node13349;
	wire [4-1:0] node13350;
	wire [4-1:0] node13351;
	wire [4-1:0] node13354;
	wire [4-1:0] node13358;
	wire [4-1:0] node13359;
	wire [4-1:0] node13360;
	wire [4-1:0] node13361;
	wire [4-1:0] node13363;
	wire [4-1:0] node13366;
	wire [4-1:0] node13368;
	wire [4-1:0] node13371;
	wire [4-1:0] node13372;
	wire [4-1:0] node13374;
	wire [4-1:0] node13377;
	wire [4-1:0] node13379;
	wire [4-1:0] node13382;
	wire [4-1:0] node13383;
	wire [4-1:0] node13384;
	wire [4-1:0] node13387;
	wire [4-1:0] node13390;
	wire [4-1:0] node13391;
	wire [4-1:0] node13394;
	wire [4-1:0] node13397;
	wire [4-1:0] node13398;
	wire [4-1:0] node13399;
	wire [4-1:0] node13400;
	wire [4-1:0] node13401;
	wire [4-1:0] node13402;
	wire [4-1:0] node13403;
	wire [4-1:0] node13404;
	wire [4-1:0] node13405;
	wire [4-1:0] node13408;
	wire [4-1:0] node13411;
	wire [4-1:0] node13413;
	wire [4-1:0] node13416;
	wire [4-1:0] node13417;
	wire [4-1:0] node13419;
	wire [4-1:0] node13422;
	wire [4-1:0] node13423;
	wire [4-1:0] node13426;
	wire [4-1:0] node13429;
	wire [4-1:0] node13430;
	wire [4-1:0] node13431;
	wire [4-1:0] node13432;
	wire [4-1:0] node13433;
	wire [4-1:0] node13436;
	wire [4-1:0] node13439;
	wire [4-1:0] node13440;
	wire [4-1:0] node13444;
	wire [4-1:0] node13446;
	wire [4-1:0] node13448;
	wire [4-1:0] node13451;
	wire [4-1:0] node13452;
	wire [4-1:0] node13453;
	wire [4-1:0] node13456;
	wire [4-1:0] node13459;
	wire [4-1:0] node13460;
	wire [4-1:0] node13461;
	wire [4-1:0] node13464;
	wire [4-1:0] node13468;
	wire [4-1:0] node13469;
	wire [4-1:0] node13470;
	wire [4-1:0] node13471;
	wire [4-1:0] node13475;
	wire [4-1:0] node13476;
	wire [4-1:0] node13478;
	wire [4-1:0] node13482;
	wire [4-1:0] node13483;
	wire [4-1:0] node13484;
	wire [4-1:0] node13485;
	wire [4-1:0] node13488;
	wire [4-1:0] node13491;
	wire [4-1:0] node13492;
	wire [4-1:0] node13496;
	wire [4-1:0] node13497;
	wire [4-1:0] node13498;
	wire [4-1:0] node13499;
	wire [4-1:0] node13503;
	wire [4-1:0] node13505;
	wire [4-1:0] node13508;
	wire [4-1:0] node13509;
	wire [4-1:0] node13512;
	wire [4-1:0] node13515;
	wire [4-1:0] node13516;
	wire [4-1:0] node13517;
	wire [4-1:0] node13518;
	wire [4-1:0] node13519;
	wire [4-1:0] node13520;
	wire [4-1:0] node13521;
	wire [4-1:0] node13524;
	wire [4-1:0] node13527;
	wire [4-1:0] node13528;
	wire [4-1:0] node13531;
	wire [4-1:0] node13534;
	wire [4-1:0] node13536;
	wire [4-1:0] node13539;
	wire [4-1:0] node13540;
	wire [4-1:0] node13541;
	wire [4-1:0] node13542;
	wire [4-1:0] node13546;
	wire [4-1:0] node13547;
	wire [4-1:0] node13550;
	wire [4-1:0] node13553;
	wire [4-1:0] node13554;
	wire [4-1:0] node13557;
	wire [4-1:0] node13560;
	wire [4-1:0] node13561;
	wire [4-1:0] node13562;
	wire [4-1:0] node13563;
	wire [4-1:0] node13566;
	wire [4-1:0] node13569;
	wire [4-1:0] node13570;
	wire [4-1:0] node13573;
	wire [4-1:0] node13576;
	wire [4-1:0] node13577;
	wire [4-1:0] node13578;
	wire [4-1:0] node13579;
	wire [4-1:0] node13583;
	wire [4-1:0] node13584;
	wire [4-1:0] node13588;
	wire [4-1:0] node13589;
	wire [4-1:0] node13590;
	wire [4-1:0] node13594;
	wire [4-1:0] node13595;
	wire [4-1:0] node13598;
	wire [4-1:0] node13601;
	wire [4-1:0] node13602;
	wire [4-1:0] node13603;
	wire [4-1:0] node13604;
	wire [4-1:0] node13605;
	wire [4-1:0] node13608;
	wire [4-1:0] node13611;
	wire [4-1:0] node13612;
	wire [4-1:0] node13615;
	wire [4-1:0] node13618;
	wire [4-1:0] node13619;
	wire [4-1:0] node13620;
	wire [4-1:0] node13621;
	wire [4-1:0] node13625;
	wire [4-1:0] node13627;
	wire [4-1:0] node13630;
	wire [4-1:0] node13631;
	wire [4-1:0] node13632;
	wire [4-1:0] node13637;
	wire [4-1:0] node13638;
	wire [4-1:0] node13639;
	wire [4-1:0] node13640;
	wire [4-1:0] node13643;
	wire [4-1:0] node13646;
	wire [4-1:0] node13647;
	wire [4-1:0] node13650;
	wire [4-1:0] node13653;
	wire [4-1:0] node13654;
	wire [4-1:0] node13655;
	wire [4-1:0] node13658;
	wire [4-1:0] node13661;
	wire [4-1:0] node13662;
	wire [4-1:0] node13665;
	wire [4-1:0] node13668;
	wire [4-1:0] node13669;
	wire [4-1:0] node13670;
	wire [4-1:0] node13671;
	wire [4-1:0] node13672;
	wire [4-1:0] node13673;
	wire [4-1:0] node13674;
	wire [4-1:0] node13678;
	wire [4-1:0] node13679;
	wire [4-1:0] node13682;
	wire [4-1:0] node13685;
	wire [4-1:0] node13686;
	wire [4-1:0] node13687;
	wire [4-1:0] node13688;
	wire [4-1:0] node13691;
	wire [4-1:0] node13694;
	wire [4-1:0] node13695;
	wire [4-1:0] node13698;
	wire [4-1:0] node13701;
	wire [4-1:0] node13703;
	wire [4-1:0] node13704;
	wire [4-1:0] node13707;
	wire [4-1:0] node13710;
	wire [4-1:0] node13711;
	wire [4-1:0] node13712;
	wire [4-1:0] node13713;
	wire [4-1:0] node13717;
	wire [4-1:0] node13718;
	wire [4-1:0] node13721;
	wire [4-1:0] node13724;
	wire [4-1:0] node13725;
	wire [4-1:0] node13726;
	wire [4-1:0] node13727;
	wire [4-1:0] node13730;
	wire [4-1:0] node13733;
	wire [4-1:0] node13734;
	wire [4-1:0] node13737;
	wire [4-1:0] node13740;
	wire [4-1:0] node13741;
	wire [4-1:0] node13744;
	wire [4-1:0] node13747;
	wire [4-1:0] node13748;
	wire [4-1:0] node13749;
	wire [4-1:0] node13752;
	wire [4-1:0] node13755;
	wire [4-1:0] node13756;
	wire [4-1:0] node13757;
	wire [4-1:0] node13758;
	wire [4-1:0] node13762;
	wire [4-1:0] node13763;
	wire [4-1:0] node13765;
	wire [4-1:0] node13768;
	wire [4-1:0] node13769;
	wire [4-1:0] node13772;
	wire [4-1:0] node13775;
	wire [4-1:0] node13776;
	wire [4-1:0] node13779;
	wire [4-1:0] node13782;
	wire [4-1:0] node13783;
	wire [4-1:0] node13784;
	wire [4-1:0] node13785;
	wire [4-1:0] node13788;
	wire [4-1:0] node13791;
	wire [4-1:0] node13792;
	wire [4-1:0] node13793;
	wire [4-1:0] node13794;
	wire [4-1:0] node13797;
	wire [4-1:0] node13800;
	wire [4-1:0] node13802;
	wire [4-1:0] node13804;
	wire [4-1:0] node13807;
	wire [4-1:0] node13809;
	wire [4-1:0] node13810;
	wire [4-1:0] node13813;
	wire [4-1:0] node13816;
	wire [4-1:0] node13817;
	wire [4-1:0] node13818;
	wire [4-1:0] node13819;
	wire [4-1:0] node13820;
	wire [4-1:0] node13821;
	wire [4-1:0] node13825;
	wire [4-1:0] node13826;
	wire [4-1:0] node13829;
	wire [4-1:0] node13832;
	wire [4-1:0] node13833;
	wire [4-1:0] node13836;
	wire [4-1:0] node13839;
	wire [4-1:0] node13840;
	wire [4-1:0] node13841;
	wire [4-1:0] node13842;
	wire [4-1:0] node13845;
	wire [4-1:0] node13848;
	wire [4-1:0] node13849;
	wire [4-1:0] node13852;
	wire [4-1:0] node13855;
	wire [4-1:0] node13856;
	wire [4-1:0] node13859;
	wire [4-1:0] node13862;
	wire [4-1:0] node13863;
	wire [4-1:0] node13864;
	wire [4-1:0] node13865;
	wire [4-1:0] node13869;
	wire [4-1:0] node13870;
	wire [4-1:0] node13873;
	wire [4-1:0] node13876;
	wire [4-1:0] node13877;
	wire [4-1:0] node13878;
	wire [4-1:0] node13881;
	wire [4-1:0] node13884;
	wire [4-1:0] node13885;
	wire [4-1:0] node13886;
	wire [4-1:0] node13890;
	wire [4-1:0] node13891;
	wire [4-1:0] node13894;
	wire [4-1:0] node13897;
	wire [4-1:0] node13898;
	wire [4-1:0] node13899;
	wire [4-1:0] node13900;
	wire [4-1:0] node13901;
	wire [4-1:0] node13902;
	wire [4-1:0] node13903;
	wire [4-1:0] node13904;
	wire [4-1:0] node13907;
	wire [4-1:0] node13910;
	wire [4-1:0] node13911;
	wire [4-1:0] node13913;
	wire [4-1:0] node13916;
	wire [4-1:0] node13917;
	wire [4-1:0] node13920;
	wire [4-1:0] node13923;
	wire [4-1:0] node13924;
	wire [4-1:0] node13926;
	wire [4-1:0] node13929;
	wire [4-1:0] node13930;
	wire [4-1:0] node13931;
	wire [4-1:0] node13934;
	wire [4-1:0] node13937;
	wire [4-1:0] node13938;
	wire [4-1:0] node13941;
	wire [4-1:0] node13944;
	wire [4-1:0] node13945;
	wire [4-1:0] node13946;
	wire [4-1:0] node13947;
	wire [4-1:0] node13949;
	wire [4-1:0] node13952;
	wire [4-1:0] node13955;
	wire [4-1:0] node13956;
	wire [4-1:0] node13959;
	wire [4-1:0] node13962;
	wire [4-1:0] node13963;
	wire [4-1:0] node13964;
	wire [4-1:0] node13965;
	wire [4-1:0] node13969;
	wire [4-1:0] node13971;
	wire [4-1:0] node13974;
	wire [4-1:0] node13975;
	wire [4-1:0] node13976;
	wire [4-1:0] node13981;
	wire [4-1:0] node13982;
	wire [4-1:0] node13983;
	wire [4-1:0] node13984;
	wire [4-1:0] node13985;
	wire [4-1:0] node13986;
	wire [4-1:0] node13989;
	wire [4-1:0] node13992;
	wire [4-1:0] node13993;
	wire [4-1:0] node13996;
	wire [4-1:0] node13999;
	wire [4-1:0] node14000;
	wire [4-1:0] node14003;
	wire [4-1:0] node14006;
	wire [4-1:0] node14007;
	wire [4-1:0] node14008;
	wire [4-1:0] node14009;
	wire [4-1:0] node14012;
	wire [4-1:0] node14015;
	wire [4-1:0] node14016;
	wire [4-1:0] node14020;
	wire [4-1:0] node14021;
	wire [4-1:0] node14022;
	wire [4-1:0] node14025;
	wire [4-1:0] node14028;
	wire [4-1:0] node14029;
	wire [4-1:0] node14033;
	wire [4-1:0] node14034;
	wire [4-1:0] node14035;
	wire [4-1:0] node14036;
	wire [4-1:0] node14039;
	wire [4-1:0] node14042;
	wire [4-1:0] node14043;
	wire [4-1:0] node14044;
	wire [4-1:0] node14048;
	wire [4-1:0] node14050;
	wire [4-1:0] node14053;
	wire [4-1:0] node14054;
	wire [4-1:0] node14056;
	wire [4-1:0] node14059;
	wire [4-1:0] node14060;
	wire [4-1:0] node14062;
	wire [4-1:0] node14065;
	wire [4-1:0] node14066;
	wire [4-1:0] node14069;
	wire [4-1:0] node14072;
	wire [4-1:0] node14073;
	wire [4-1:0] node14074;
	wire [4-1:0] node14075;
	wire [4-1:0] node14076;
	wire [4-1:0] node14079;
	wire [4-1:0] node14082;
	wire [4-1:0] node14083;
	wire [4-1:0] node14086;
	wire [4-1:0] node14089;
	wire [4-1:0] node14090;
	wire [4-1:0] node14091;
	wire [4-1:0] node14092;
	wire [4-1:0] node14093;
	wire [4-1:0] node14096;
	wire [4-1:0] node14099;
	wire [4-1:0] node14101;
	wire [4-1:0] node14104;
	wire [4-1:0] node14105;
	wire [4-1:0] node14108;
	wire [4-1:0] node14111;
	wire [4-1:0] node14112;
	wire [4-1:0] node14115;
	wire [4-1:0] node14118;
	wire [4-1:0] node14119;
	wire [4-1:0] node14120;
	wire [4-1:0] node14121;
	wire [4-1:0] node14122;
	wire [4-1:0] node14124;
	wire [4-1:0] node14128;
	wire [4-1:0] node14129;
	wire [4-1:0] node14130;
	wire [4-1:0] node14134;
	wire [4-1:0] node14136;
	wire [4-1:0] node14139;
	wire [4-1:0] node14140;
	wire [4-1:0] node14142;
	wire [4-1:0] node14143;
	wire [4-1:0] node14146;
	wire [4-1:0] node14149;
	wire [4-1:0] node14150;
	wire [4-1:0] node14153;
	wire [4-1:0] node14154;
	wire [4-1:0] node14157;
	wire [4-1:0] node14160;
	wire [4-1:0] node14161;
	wire [4-1:0] node14162;
	wire [4-1:0] node14163;
	wire [4-1:0] node14164;
	wire [4-1:0] node14167;
	wire [4-1:0] node14170;
	wire [4-1:0] node14172;
	wire [4-1:0] node14175;
	wire [4-1:0] node14177;
	wire [4-1:0] node14178;
	wire [4-1:0] node14181;
	wire [4-1:0] node14184;
	wire [4-1:0] node14185;
	wire [4-1:0] node14186;
	wire [4-1:0] node14187;
	wire [4-1:0] node14190;
	wire [4-1:0] node14193;
	wire [4-1:0] node14194;
	wire [4-1:0] node14197;
	wire [4-1:0] node14200;
	wire [4-1:0] node14201;
	wire [4-1:0] node14202;
	wire [4-1:0] node14205;
	wire [4-1:0] node14208;
	wire [4-1:0] node14209;
	wire [4-1:0] node14212;
	wire [4-1:0] node14215;
	wire [4-1:0] node14216;
	wire [4-1:0] node14217;
	wire [4-1:0] node14218;
	wire [4-1:0] node14219;
	wire [4-1:0] node14220;
	wire [4-1:0] node14221;
	wire [4-1:0] node14224;
	wire [4-1:0] node14226;
	wire [4-1:0] node14229;
	wire [4-1:0] node14230;
	wire [4-1:0] node14231;
	wire [4-1:0] node14235;
	wire [4-1:0] node14238;
	wire [4-1:0] node14239;
	wire [4-1:0] node14240;
	wire [4-1:0] node14241;
	wire [4-1:0] node14244;
	wire [4-1:0] node14248;
	wire [4-1:0] node14249;
	wire [4-1:0] node14250;
	wire [4-1:0] node14253;
	wire [4-1:0] node14256;
	wire [4-1:0] node14257;
	wire [4-1:0] node14260;
	wire [4-1:0] node14263;
	wire [4-1:0] node14264;
	wire [4-1:0] node14265;
	wire [4-1:0] node14267;
	wire [4-1:0] node14269;
	wire [4-1:0] node14272;
	wire [4-1:0] node14274;
	wire [4-1:0] node14275;
	wire [4-1:0] node14278;
	wire [4-1:0] node14281;
	wire [4-1:0] node14282;
	wire [4-1:0] node14283;
	wire [4-1:0] node14284;
	wire [4-1:0] node14287;
	wire [4-1:0] node14290;
	wire [4-1:0] node14291;
	wire [4-1:0] node14294;
	wire [4-1:0] node14297;
	wire [4-1:0] node14298;
	wire [4-1:0] node14300;
	wire [4-1:0] node14303;
	wire [4-1:0] node14305;
	wire [4-1:0] node14308;
	wire [4-1:0] node14309;
	wire [4-1:0] node14310;
	wire [4-1:0] node14312;
	wire [4-1:0] node14313;
	wire [4-1:0] node14316;
	wire [4-1:0] node14319;
	wire [4-1:0] node14320;
	wire [4-1:0] node14321;
	wire [4-1:0] node14322;
	wire [4-1:0] node14325;
	wire [4-1:0] node14328;
	wire [4-1:0] node14330;
	wire [4-1:0] node14333;
	wire [4-1:0] node14334;
	wire [4-1:0] node14336;
	wire [4-1:0] node14339;
	wire [4-1:0] node14340;
	wire [4-1:0] node14343;
	wire [4-1:0] node14346;
	wire [4-1:0] node14347;
	wire [4-1:0] node14348;
	wire [4-1:0] node14349;
	wire [4-1:0] node14350;
	wire [4-1:0] node14353;
	wire [4-1:0] node14356;
	wire [4-1:0] node14357;
	wire [4-1:0] node14360;
	wire [4-1:0] node14363;
	wire [4-1:0] node14364;
	wire [4-1:0] node14366;
	wire [4-1:0] node14369;
	wire [4-1:0] node14370;
	wire [4-1:0] node14373;
	wire [4-1:0] node14376;
	wire [4-1:0] node14377;
	wire [4-1:0] node14379;
	wire [4-1:0] node14382;
	wire [4-1:0] node14384;
	wire [4-1:0] node14387;
	wire [4-1:0] node14388;
	wire [4-1:0] node14389;
	wire [4-1:0] node14390;
	wire [4-1:0] node14391;
	wire [4-1:0] node14392;
	wire [4-1:0] node14395;
	wire [4-1:0] node14399;
	wire [4-1:0] node14400;
	wire [4-1:0] node14401;
	wire [4-1:0] node14404;
	wire [4-1:0] node14407;
	wire [4-1:0] node14408;
	wire [4-1:0] node14411;
	wire [4-1:0] node14414;
	wire [4-1:0] node14415;
	wire [4-1:0] node14416;
	wire [4-1:0] node14418;
	wire [4-1:0] node14421;
	wire [4-1:0] node14423;
	wire [4-1:0] node14424;
	wire [4-1:0] node14427;
	wire [4-1:0] node14430;
	wire [4-1:0] node14431;
	wire [4-1:0] node14434;
	wire [4-1:0] node14437;
	wire [4-1:0] node14438;
	wire [4-1:0] node14439;
	wire [4-1:0] node14440;
	wire [4-1:0] node14441;
	wire [4-1:0] node14443;
	wire [4-1:0] node14446;
	wire [4-1:0] node14447;
	wire [4-1:0] node14451;
	wire [4-1:0] node14452;
	wire [4-1:0] node14456;
	wire [4-1:0] node14457;
	wire [4-1:0] node14460;
	wire [4-1:0] node14463;
	wire [4-1:0] node14464;
	wire [4-1:0] node14465;
	wire [4-1:0] node14466;
	wire [4-1:0] node14469;
	wire [4-1:0] node14472;
	wire [4-1:0] node14474;
	wire [4-1:0] node14475;
	wire [4-1:0] node14478;
	wire [4-1:0] node14481;
	wire [4-1:0] node14482;
	wire [4-1:0] node14483;
	wire [4-1:0] node14486;
	wire [4-1:0] node14489;
	wire [4-1:0] node14490;
	wire [4-1:0] node14493;
	wire [4-1:0] node14496;
	wire [4-1:0] node14497;
	wire [4-1:0] node14498;
	wire [4-1:0] node14499;
	wire [4-1:0] node14500;
	wire [4-1:0] node14501;
	wire [4-1:0] node14502;
	wire [4-1:0] node14503;
	wire [4-1:0] node14504;
	wire [4-1:0] node14505;
	wire [4-1:0] node14506;
	wire [4-1:0] node14511;
	wire [4-1:0] node14513;
	wire [4-1:0] node14514;
	wire [4-1:0] node14517;
	wire [4-1:0] node14520;
	wire [4-1:0] node14521;
	wire [4-1:0] node14522;
	wire [4-1:0] node14523;
	wire [4-1:0] node14526;
	wire [4-1:0] node14529;
	wire [4-1:0] node14531;
	wire [4-1:0] node14534;
	wire [4-1:0] node14536;
	wire [4-1:0] node14537;
	wire [4-1:0] node14540;
	wire [4-1:0] node14543;
	wire [4-1:0] node14544;
	wire [4-1:0] node14545;
	wire [4-1:0] node14547;
	wire [4-1:0] node14548;
	wire [4-1:0] node14552;
	wire [4-1:0] node14553;
	wire [4-1:0] node14554;
	wire [4-1:0] node14557;
	wire [4-1:0] node14560;
	wire [4-1:0] node14561;
	wire [4-1:0] node14565;
	wire [4-1:0] node14566;
	wire [4-1:0] node14567;
	wire [4-1:0] node14569;
	wire [4-1:0] node14572;
	wire [4-1:0] node14573;
	wire [4-1:0] node14576;
	wire [4-1:0] node14579;
	wire [4-1:0] node14582;
	wire [4-1:0] node14583;
	wire [4-1:0] node14584;
	wire [4-1:0] node14585;
	wire [4-1:0] node14586;
	wire [4-1:0] node14589;
	wire [4-1:0] node14592;
	wire [4-1:0] node14593;
	wire [4-1:0] node14594;
	wire [4-1:0] node14598;
	wire [4-1:0] node14599;
	wire [4-1:0] node14603;
	wire [4-1:0] node14604;
	wire [4-1:0] node14605;
	wire [4-1:0] node14607;
	wire [4-1:0] node14610;
	wire [4-1:0] node14612;
	wire [4-1:0] node14615;
	wire [4-1:0] node14616;
	wire [4-1:0] node14619;
	wire [4-1:0] node14622;
	wire [4-1:0] node14623;
	wire [4-1:0] node14624;
	wire [4-1:0] node14625;
	wire [4-1:0] node14626;
	wire [4-1:0] node14629;
	wire [4-1:0] node14632;
	wire [4-1:0] node14633;
	wire [4-1:0] node14637;
	wire [4-1:0] node14638;
	wire [4-1:0] node14639;
	wire [4-1:0] node14643;
	wire [4-1:0] node14644;
	wire [4-1:0] node14648;
	wire [4-1:0] node14649;
	wire [4-1:0] node14650;
	wire [4-1:0] node14651;
	wire [4-1:0] node14656;
	wire [4-1:0] node14657;
	wire [4-1:0] node14660;
	wire [4-1:0] node14663;
	wire [4-1:0] node14664;
	wire [4-1:0] node14665;
	wire [4-1:0] node14666;
	wire [4-1:0] node14667;
	wire [4-1:0] node14668;
	wire [4-1:0] node14671;
	wire [4-1:0] node14674;
	wire [4-1:0] node14676;
	wire [4-1:0] node14677;
	wire [4-1:0] node14681;
	wire [4-1:0] node14682;
	wire [4-1:0] node14684;
	wire [4-1:0] node14687;
	wire [4-1:0] node14689;
	wire [4-1:0] node14692;
	wire [4-1:0] node14693;
	wire [4-1:0] node14694;
	wire [4-1:0] node14695;
	wire [4-1:0] node14698;
	wire [4-1:0] node14701;
	wire [4-1:0] node14703;
	wire [4-1:0] node14705;
	wire [4-1:0] node14708;
	wire [4-1:0] node14709;
	wire [4-1:0] node14710;
	wire [4-1:0] node14713;
	wire [4-1:0] node14716;
	wire [4-1:0] node14718;
	wire [4-1:0] node14721;
	wire [4-1:0] node14722;
	wire [4-1:0] node14723;
	wire [4-1:0] node14725;
	wire [4-1:0] node14726;
	wire [4-1:0] node14729;
	wire [4-1:0] node14732;
	wire [4-1:0] node14733;
	wire [4-1:0] node14734;
	wire [4-1:0] node14735;
	wire [4-1:0] node14739;
	wire [4-1:0] node14740;
	wire [4-1:0] node14744;
	wire [4-1:0] node14745;
	wire [4-1:0] node14746;
	wire [4-1:0] node14751;
	wire [4-1:0] node14752;
	wire [4-1:0] node14753;
	wire [4-1:0] node14754;
	wire [4-1:0] node14755;
	wire [4-1:0] node14758;
	wire [4-1:0] node14762;
	wire [4-1:0] node14763;
	wire [4-1:0] node14764;
	wire [4-1:0] node14768;
	wire [4-1:0] node14770;
	wire [4-1:0] node14773;
	wire [4-1:0] node14774;
	wire [4-1:0] node14775;
	wire [4-1:0] node14778;
	wire [4-1:0] node14781;
	wire [4-1:0] node14782;
	wire [4-1:0] node14783;
	wire [4-1:0] node14786;
	wire [4-1:0] node14789;
	wire [4-1:0] node14790;
	wire [4-1:0] node14794;
	wire [4-1:0] node14795;
	wire [4-1:0] node14796;
	wire [4-1:0] node14797;
	wire [4-1:0] node14798;
	wire [4-1:0] node14799;
	wire [4-1:0] node14802;
	wire [4-1:0] node14805;
	wire [4-1:0] node14806;
	wire [4-1:0] node14807;
	wire [4-1:0] node14811;
	wire [4-1:0] node14812;
	wire [4-1:0] node14813;
	wire [4-1:0] node14816;
	wire [4-1:0] node14819;
	wire [4-1:0] node14820;
	wire [4-1:0] node14824;
	wire [4-1:0] node14825;
	wire [4-1:0] node14826;
	wire [4-1:0] node14827;
	wire [4-1:0] node14828;
	wire [4-1:0] node14831;
	wire [4-1:0] node14834;
	wire [4-1:0] node14836;
	wire [4-1:0] node14839;
	wire [4-1:0] node14840;
	wire [4-1:0] node14841;
	wire [4-1:0] node14844;
	wire [4-1:0] node14847;
	wire [4-1:0] node14848;
	wire [4-1:0] node14851;
	wire [4-1:0] node14854;
	wire [4-1:0] node14855;
	wire [4-1:0] node14859;
	wire [4-1:0] node14860;
	wire [4-1:0] node14861;
	wire [4-1:0] node14863;
	wire [4-1:0] node14866;
	wire [4-1:0] node14868;
	wire [4-1:0] node14871;
	wire [4-1:0] node14872;
	wire [4-1:0] node14874;
	wire [4-1:0] node14877;
	wire [4-1:0] node14879;
	wire [4-1:0] node14882;
	wire [4-1:0] node14883;
	wire [4-1:0] node14884;
	wire [4-1:0] node14885;
	wire [4-1:0] node14886;
	wire [4-1:0] node14888;
	wire [4-1:0] node14891;
	wire [4-1:0] node14893;
	wire [4-1:0] node14896;
	wire [4-1:0] node14897;
	wire [4-1:0] node14901;
	wire [4-1:0] node14902;
	wire [4-1:0] node14904;
	wire [4-1:0] node14907;
	wire [4-1:0] node14908;
	wire [4-1:0] node14910;
	wire [4-1:0] node14913;
	wire [4-1:0] node14915;
	wire [4-1:0] node14918;
	wire [4-1:0] node14919;
	wire [4-1:0] node14920;
	wire [4-1:0] node14921;
	wire [4-1:0] node14923;
	wire [4-1:0] node14926;
	wire [4-1:0] node14928;
	wire [4-1:0] node14931;
	wire [4-1:0] node14932;
	wire [4-1:0] node14934;
	wire [4-1:0] node14937;
	wire [4-1:0] node14939;
	wire [4-1:0] node14942;
	wire [4-1:0] node14943;
	wire [4-1:0] node14944;
	wire [4-1:0] node14947;
	wire [4-1:0] node14950;
	wire [4-1:0] node14951;
	wire [4-1:0] node14953;
	wire [4-1:0] node14956;
	wire [4-1:0] node14957;
	wire [4-1:0] node14960;
	wire [4-1:0] node14963;
	wire [4-1:0] node14964;
	wire [4-1:0] node14965;
	wire [4-1:0] node14966;
	wire [4-1:0] node14967;
	wire [4-1:0] node14968;
	wire [4-1:0] node14969;
	wire [4-1:0] node14970;
	wire [4-1:0] node14973;
	wire [4-1:0] node14976;
	wire [4-1:0] node14977;
	wire [4-1:0] node14980;
	wire [4-1:0] node14983;
	wire [4-1:0] node14984;
	wire [4-1:0] node14987;
	wire [4-1:0] node14990;
	wire [4-1:0] node14991;
	wire [4-1:0] node14992;
	wire [4-1:0] node14993;
	wire [4-1:0] node14997;
	wire [4-1:0] node14998;
	wire [4-1:0] node15002;
	wire [4-1:0] node15003;
	wire [4-1:0] node15004;
	wire [4-1:0] node15005;
	wire [4-1:0] node15008;
	wire [4-1:0] node15012;
	wire [4-1:0] node15013;
	wire [4-1:0] node15014;
	wire [4-1:0] node15017;
	wire [4-1:0] node15021;
	wire [4-1:0] node15022;
	wire [4-1:0] node15023;
	wire [4-1:0] node15024;
	wire [4-1:0] node15026;
	wire [4-1:0] node15027;
	wire [4-1:0] node15030;
	wire [4-1:0] node15033;
	wire [4-1:0] node15034;
	wire [4-1:0] node15037;
	wire [4-1:0] node15040;
	wire [4-1:0] node15041;
	wire [4-1:0] node15044;
	wire [4-1:0] node15047;
	wire [4-1:0] node15048;
	wire [4-1:0] node15051;
	wire [4-1:0] node15052;
	wire [4-1:0] node15053;
	wire [4-1:0] node15054;
	wire [4-1:0] node15058;
	wire [4-1:0] node15059;
	wire [4-1:0] node15064;
	wire [4-1:0] node15065;
	wire [4-1:0] node15066;
	wire [4-1:0] node15067;
	wire [4-1:0] node15068;
	wire [4-1:0] node15069;
	wire [4-1:0] node15070;
	wire [4-1:0] node15073;
	wire [4-1:0] node15076;
	wire [4-1:0] node15077;
	wire [4-1:0] node15080;
	wire [4-1:0] node15083;
	wire [4-1:0] node15084;
	wire [4-1:0] node15085;
	wire [4-1:0] node15088;
	wire [4-1:0] node15091;
	wire [4-1:0] node15092;
	wire [4-1:0] node15095;
	wire [4-1:0] node15098;
	wire [4-1:0] node15099;
	wire [4-1:0] node15102;
	wire [4-1:0] node15105;
	wire [4-1:0] node15106;
	wire [4-1:0] node15107;
	wire [4-1:0] node15108;
	wire [4-1:0] node15109;
	wire [4-1:0] node15113;
	wire [4-1:0] node15114;
	wire [4-1:0] node15117;
	wire [4-1:0] node15120;
	wire [4-1:0] node15122;
	wire [4-1:0] node15125;
	wire [4-1:0] node15126;
	wire [4-1:0] node15128;
	wire [4-1:0] node15129;
	wire [4-1:0] node15133;
	wire [4-1:0] node15134;
	wire [4-1:0] node15135;
	wire [4-1:0] node15139;
	wire [4-1:0] node15140;
	wire [4-1:0] node15144;
	wire [4-1:0] node15145;
	wire [4-1:0] node15146;
	wire [4-1:0] node15148;
	wire [4-1:0] node15149;
	wire [4-1:0] node15153;
	wire [4-1:0] node15155;
	wire [4-1:0] node15156;
	wire [4-1:0] node15160;
	wire [4-1:0] node15161;
	wire [4-1:0] node15162;
	wire [4-1:0] node15163;
	wire [4-1:0] node15165;
	wire [4-1:0] node15168;
	wire [4-1:0] node15170;
	wire [4-1:0] node15174;
	wire [4-1:0] node15175;
	wire [4-1:0] node15176;
	wire [4-1:0] node15179;
	wire [4-1:0] node15182;
	wire [4-1:0] node15184;
	wire [4-1:0] node15187;
	wire [4-1:0] node15188;
	wire [4-1:0] node15189;
	wire [4-1:0] node15190;
	wire [4-1:0] node15191;
	wire [4-1:0] node15192;
	wire [4-1:0] node15193;
	wire [4-1:0] node15197;
	wire [4-1:0] node15198;
	wire [4-1:0] node15202;
	wire [4-1:0] node15203;
	wire [4-1:0] node15204;
	wire [4-1:0] node15205;
	wire [4-1:0] node15209;
	wire [4-1:0] node15210;
	wire [4-1:0] node15214;
	wire [4-1:0] node15215;
	wire [4-1:0] node15216;
	wire [4-1:0] node15221;
	wire [4-1:0] node15222;
	wire [4-1:0] node15223;
	wire [4-1:0] node15224;
	wire [4-1:0] node15225;
	wire [4-1:0] node15229;
	wire [4-1:0] node15230;
	wire [4-1:0] node15233;
	wire [4-1:0] node15236;
	wire [4-1:0] node15237;
	wire [4-1:0] node15238;
	wire [4-1:0] node15241;
	wire [4-1:0] node15245;
	wire [4-1:0] node15246;
	wire [4-1:0] node15247;
	wire [4-1:0] node15250;
	wire [4-1:0] node15253;
	wire [4-1:0] node15254;
	wire [4-1:0] node15257;
	wire [4-1:0] node15260;
	wire [4-1:0] node15261;
	wire [4-1:0] node15262;
	wire [4-1:0] node15263;
	wire [4-1:0] node15264;
	wire [4-1:0] node15265;
	wire [4-1:0] node15269;
	wire [4-1:0] node15270;
	wire [4-1:0] node15273;
	wire [4-1:0] node15276;
	wire [4-1:0] node15277;
	wire [4-1:0] node15279;
	wire [4-1:0] node15282;
	wire [4-1:0] node15285;
	wire [4-1:0] node15286;
	wire [4-1:0] node15288;
	wire [4-1:0] node15291;
	wire [4-1:0] node15293;
	wire [4-1:0] node15294;
	wire [4-1:0] node15298;
	wire [4-1:0] node15299;
	wire [4-1:0] node15300;
	wire [4-1:0] node15301;
	wire [4-1:0] node15305;
	wire [4-1:0] node15306;
	wire [4-1:0] node15310;
	wire [4-1:0] node15312;
	wire [4-1:0] node15313;
	wire [4-1:0] node15317;
	wire [4-1:0] node15318;
	wire [4-1:0] node15319;
	wire [4-1:0] node15320;
	wire [4-1:0] node15321;
	wire [4-1:0] node15322;
	wire [4-1:0] node15324;
	wire [4-1:0] node15328;
	wire [4-1:0] node15329;
	wire [4-1:0] node15332;
	wire [4-1:0] node15335;
	wire [4-1:0] node15336;
	wire [4-1:0] node15337;
	wire [4-1:0] node15338;
	wire [4-1:0] node15342;
	wire [4-1:0] node15343;
	wire [4-1:0] node15347;
	wire [4-1:0] node15348;
	wire [4-1:0] node15352;
	wire [4-1:0] node15353;
	wire [4-1:0] node15354;
	wire [4-1:0] node15356;
	wire [4-1:0] node15357;
	wire [4-1:0] node15360;
	wire [4-1:0] node15363;
	wire [4-1:0] node15364;
	wire [4-1:0] node15365;
	wire [4-1:0] node15368;
	wire [4-1:0] node15372;
	wire [4-1:0] node15373;
	wire [4-1:0] node15376;
	wire [4-1:0] node15379;
	wire [4-1:0] node15380;
	wire [4-1:0] node15381;
	wire [4-1:0] node15382;
	wire [4-1:0] node15383;
	wire [4-1:0] node15384;
	wire [4-1:0] node15387;
	wire [4-1:0] node15390;
	wire [4-1:0] node15392;
	wire [4-1:0] node15395;
	wire [4-1:0] node15396;
	wire [4-1:0] node15399;
	wire [4-1:0] node15402;
	wire [4-1:0] node15403;
	wire [4-1:0] node15405;
	wire [4-1:0] node15406;
	wire [4-1:0] node15410;
	wire [4-1:0] node15411;
	wire [4-1:0] node15415;
	wire [4-1:0] node15416;
	wire [4-1:0] node15417;
	wire [4-1:0] node15418;
	wire [4-1:0] node15422;
	wire [4-1:0] node15423;
	wire [4-1:0] node15427;
	wire [4-1:0] node15428;
	wire [4-1:0] node15429;
	wire [4-1:0] node15433;
	wire [4-1:0] node15434;
	wire [4-1:0] node15438;
	wire [4-1:0] node15439;
	wire [4-1:0] node15440;
	wire [4-1:0] node15441;
	wire [4-1:0] node15442;
	wire [4-1:0] node15443;
	wire [4-1:0] node15444;
	wire [4-1:0] node15445;
	wire [4-1:0] node15446;
	wire [4-1:0] node15447;
	wire [4-1:0] node15450;
	wire [4-1:0] node15453;
	wire [4-1:0] node15456;
	wire [4-1:0] node15457;
	wire [4-1:0] node15459;
	wire [4-1:0] node15462;
	wire [4-1:0] node15463;
	wire [4-1:0] node15466;
	wire [4-1:0] node15469;
	wire [4-1:0] node15470;
	wire [4-1:0] node15471;
	wire [4-1:0] node15474;
	wire [4-1:0] node15476;
	wire [4-1:0] node15479;
	wire [4-1:0] node15480;
	wire [4-1:0] node15481;
	wire [4-1:0] node15484;
	wire [4-1:0] node15487;
	wire [4-1:0] node15488;
	wire [4-1:0] node15492;
	wire [4-1:0] node15493;
	wire [4-1:0] node15494;
	wire [4-1:0] node15495;
	wire [4-1:0] node15496;
	wire [4-1:0] node15499;
	wire [4-1:0] node15503;
	wire [4-1:0] node15504;
	wire [4-1:0] node15505;
	wire [4-1:0] node15508;
	wire [4-1:0] node15511;
	wire [4-1:0] node15512;
	wire [4-1:0] node15515;
	wire [4-1:0] node15518;
	wire [4-1:0] node15519;
	wire [4-1:0] node15520;
	wire [4-1:0] node15521;
	wire [4-1:0] node15524;
	wire [4-1:0] node15527;
	wire [4-1:0] node15528;
	wire [4-1:0] node15531;
	wire [4-1:0] node15534;
	wire [4-1:0] node15536;
	wire [4-1:0] node15538;
	wire [4-1:0] node15541;
	wire [4-1:0] node15542;
	wire [4-1:0] node15543;
	wire [4-1:0] node15544;
	wire [4-1:0] node15545;
	wire [4-1:0] node15546;
	wire [4-1:0] node15550;
	wire [4-1:0] node15551;
	wire [4-1:0] node15554;
	wire [4-1:0] node15557;
	wire [4-1:0] node15558;
	wire [4-1:0] node15560;
	wire [4-1:0] node15563;
	wire [4-1:0] node15564;
	wire [4-1:0] node15567;
	wire [4-1:0] node15570;
	wire [4-1:0] node15571;
	wire [4-1:0] node15572;
	wire [4-1:0] node15574;
	wire [4-1:0] node15578;
	wire [4-1:0] node15579;
	wire [4-1:0] node15580;
	wire [4-1:0] node15583;
	wire [4-1:0] node15586;
	wire [4-1:0] node15587;
	wire [4-1:0] node15590;
	wire [4-1:0] node15593;
	wire [4-1:0] node15594;
	wire [4-1:0] node15595;
	wire [4-1:0] node15596;
	wire [4-1:0] node15599;
	wire [4-1:0] node15600;
	wire [4-1:0] node15603;
	wire [4-1:0] node15606;
	wire [4-1:0] node15608;
	wire [4-1:0] node15610;
	wire [4-1:0] node15613;
	wire [4-1:0] node15614;
	wire [4-1:0] node15615;
	wire [4-1:0] node15616;
	wire [4-1:0] node15620;
	wire [4-1:0] node15621;
	wire [4-1:0] node15624;
	wire [4-1:0] node15627;
	wire [4-1:0] node15628;
	wire [4-1:0] node15629;
	wire [4-1:0] node15632;
	wire [4-1:0] node15636;
	wire [4-1:0] node15637;
	wire [4-1:0] node15638;
	wire [4-1:0] node15639;
	wire [4-1:0] node15640;
	wire [4-1:0] node15643;
	wire [4-1:0] node15644;
	wire [4-1:0] node15645;
	wire [4-1:0] node15648;
	wire [4-1:0] node15651;
	wire [4-1:0] node15652;
	wire [4-1:0] node15655;
	wire [4-1:0] node15658;
	wire [4-1:0] node15659;
	wire [4-1:0] node15660;
	wire [4-1:0] node15663;
	wire [4-1:0] node15666;
	wire [4-1:0] node15668;
	wire [4-1:0] node15669;
	wire [4-1:0] node15673;
	wire [4-1:0] node15674;
	wire [4-1:0] node15675;
	wire [4-1:0] node15677;
	wire [4-1:0] node15679;
	wire [4-1:0] node15682;
	wire [4-1:0] node15683;
	wire [4-1:0] node15686;
	wire [4-1:0] node15689;
	wire [4-1:0] node15690;
	wire [4-1:0] node15692;
	wire [4-1:0] node15695;
	wire [4-1:0] node15696;
	wire [4-1:0] node15699;
	wire [4-1:0] node15702;
	wire [4-1:0] node15703;
	wire [4-1:0] node15704;
	wire [4-1:0] node15705;
	wire [4-1:0] node15706;
	wire [4-1:0] node15707;
	wire [4-1:0] node15711;
	wire [4-1:0] node15712;
	wire [4-1:0] node15715;
	wire [4-1:0] node15718;
	wire [4-1:0] node15719;
	wire [4-1:0] node15720;
	wire [4-1:0] node15725;
	wire [4-1:0] node15726;
	wire [4-1:0] node15727;
	wire [4-1:0] node15728;
	wire [4-1:0] node15731;
	wire [4-1:0] node15734;
	wire [4-1:0] node15735;
	wire [4-1:0] node15739;
	wire [4-1:0] node15740;
	wire [4-1:0] node15741;
	wire [4-1:0] node15744;
	wire [4-1:0] node15748;
	wire [4-1:0] node15749;
	wire [4-1:0] node15750;
	wire [4-1:0] node15751;
	wire [4-1:0] node15755;
	wire [4-1:0] node15756;
	wire [4-1:0] node15759;
	wire [4-1:0] node15762;
	wire [4-1:0] node15763;
	wire [4-1:0] node15764;
	wire [4-1:0] node15767;
	wire [4-1:0] node15770;
	wire [4-1:0] node15771;
	wire [4-1:0] node15774;
	wire [4-1:0] node15777;
	wire [4-1:0] node15778;
	wire [4-1:0] node15779;
	wire [4-1:0] node15780;
	wire [4-1:0] node15781;
	wire [4-1:0] node15782;
	wire [4-1:0] node15783;
	wire [4-1:0] node15785;
	wire [4-1:0] node15788;
	wire [4-1:0] node15792;
	wire [4-1:0] node15793;
	wire [4-1:0] node15794;
	wire [4-1:0] node15797;
	wire [4-1:0] node15800;
	wire [4-1:0] node15801;
	wire [4-1:0] node15804;
	wire [4-1:0] node15807;
	wire [4-1:0] node15808;
	wire [4-1:0] node15809;
	wire [4-1:0] node15810;
	wire [4-1:0] node15813;
	wire [4-1:0] node15817;
	wire [4-1:0] node15818;
	wire [4-1:0] node15819;
	wire [4-1:0] node15822;
	wire [4-1:0] node15825;
	wire [4-1:0] node15826;
	wire [4-1:0] node15827;
	wire [4-1:0] node15830;
	wire [4-1:0] node15833;
	wire [4-1:0] node15834;
	wire [4-1:0] node15837;
	wire [4-1:0] node15840;
	wire [4-1:0] node15841;
	wire [4-1:0] node15842;
	wire [4-1:0] node15843;
	wire [4-1:0] node15845;
	wire [4-1:0] node15846;
	wire [4-1:0] node15849;
	wire [4-1:0] node15852;
	wire [4-1:0] node15853;
	wire [4-1:0] node15857;
	wire [4-1:0] node15858;
	wire [4-1:0] node15859;
	wire [4-1:0] node15862;
	wire [4-1:0] node15863;
	wire [4-1:0] node15867;
	wire [4-1:0] node15869;
	wire [4-1:0] node15872;
	wire [4-1:0] node15873;
	wire [4-1:0] node15874;
	wire [4-1:0] node15875;
	wire [4-1:0] node15880;
	wire [4-1:0] node15881;
	wire [4-1:0] node15882;
	wire [4-1:0] node15886;
	wire [4-1:0] node15887;
	wire [4-1:0] node15891;
	wire [4-1:0] node15892;
	wire [4-1:0] node15893;
	wire [4-1:0] node15894;
	wire [4-1:0] node15895;
	wire [4-1:0] node15896;
	wire [4-1:0] node15898;
	wire [4-1:0] node15901;
	wire [4-1:0] node15902;
	wire [4-1:0] node15906;
	wire [4-1:0] node15907;
	wire [4-1:0] node15908;
	wire [4-1:0] node15911;
	wire [4-1:0] node15915;
	wire [4-1:0] node15916;
	wire [4-1:0] node15918;
	wire [4-1:0] node15921;
	wire [4-1:0] node15922;
	wire [4-1:0] node15923;
	wire [4-1:0] node15926;
	wire [4-1:0] node15929;
	wire [4-1:0] node15930;
	wire [4-1:0] node15934;
	wire [4-1:0] node15935;
	wire [4-1:0] node15936;
	wire [4-1:0] node15937;
	wire [4-1:0] node15940;
	wire [4-1:0] node15943;
	wire [4-1:0] node15944;
	wire [4-1:0] node15948;
	wire [4-1:0] node15949;
	wire [4-1:0] node15950;
	wire [4-1:0] node15953;
	wire [4-1:0] node15956;
	wire [4-1:0] node15957;
	wire [4-1:0] node15958;
	wire [4-1:0] node15961;
	wire [4-1:0] node15964;
	wire [4-1:0] node15965;
	wire [4-1:0] node15968;
	wire [4-1:0] node15971;
	wire [4-1:0] node15972;
	wire [4-1:0] node15973;
	wire [4-1:0] node15974;
	wire [4-1:0] node15976;
	wire [4-1:0] node15977;
	wire [4-1:0] node15981;
	wire [4-1:0] node15982;
	wire [4-1:0] node15985;
	wire [4-1:0] node15988;
	wire [4-1:0] node15989;
	wire [4-1:0] node15990;
	wire [4-1:0] node15991;
	wire [4-1:0] node15994;
	wire [4-1:0] node15997;
	wire [4-1:0] node16000;
	wire [4-1:0] node16002;
	wire [4-1:0] node16005;
	wire [4-1:0] node16006;
	wire [4-1:0] node16007;
	wire [4-1:0] node16008;
	wire [4-1:0] node16009;
	wire [4-1:0] node16012;
	wire [4-1:0] node16015;
	wire [4-1:0] node16017;
	wire [4-1:0] node16020;
	wire [4-1:0] node16021;
	wire [4-1:0] node16022;
	wire [4-1:0] node16025;
	wire [4-1:0] node16028;
	wire [4-1:0] node16030;
	wire [4-1:0] node16033;
	wire [4-1:0] node16034;
	wire [4-1:0] node16035;
	wire [4-1:0] node16038;
	wire [4-1:0] node16039;
	wire [4-1:0] node16043;
	wire [4-1:0] node16044;
	wire [4-1:0] node16047;
	wire [4-1:0] node16050;
	wire [4-1:0] node16051;
	wire [4-1:0] node16052;
	wire [4-1:0] node16053;
	wire [4-1:0] node16054;
	wire [4-1:0] node16055;
	wire [4-1:0] node16056;
	wire [4-1:0] node16057;
	wire [4-1:0] node16058;
	wire [4-1:0] node16062;
	wire [4-1:0] node16063;
	wire [4-1:0] node16067;
	wire [4-1:0] node16068;
	wire [4-1:0] node16072;
	wire [4-1:0] node16074;
	wire [4-1:0] node16075;
	wire [4-1:0] node16076;
	wire [4-1:0] node16081;
	wire [4-1:0] node16082;
	wire [4-1:0] node16083;
	wire [4-1:0] node16084;
	wire [4-1:0] node16088;
	wire [4-1:0] node16089;
	wire [4-1:0] node16093;
	wire [4-1:0] node16094;
	wire [4-1:0] node16095;
	wire [4-1:0] node16099;
	wire [4-1:0] node16100;
	wire [4-1:0] node16104;
	wire [4-1:0] node16105;
	wire [4-1:0] node16106;
	wire [4-1:0] node16107;
	wire [4-1:0] node16108;
	wire [4-1:0] node16112;
	wire [4-1:0] node16113;
	wire [4-1:0] node16116;
	wire [4-1:0] node16119;
	wire [4-1:0] node16120;
	wire [4-1:0] node16121;
	wire [4-1:0] node16122;
	wire [4-1:0] node16127;
	wire [4-1:0] node16128;
	wire [4-1:0] node16132;
	wire [4-1:0] node16133;
	wire [4-1:0] node16134;
	wire [4-1:0] node16135;
	wire [4-1:0] node16139;
	wire [4-1:0] node16140;
	wire [4-1:0] node16144;
	wire [4-1:0] node16145;
	wire [4-1:0] node16146;
	wire [4-1:0] node16150;
	wire [4-1:0] node16151;
	wire [4-1:0] node16155;
	wire [4-1:0] node16156;
	wire [4-1:0] node16157;
	wire [4-1:0] node16158;
	wire [4-1:0] node16159;
	wire [4-1:0] node16160;
	wire [4-1:0] node16161;
	wire [4-1:0] node16164;
	wire [4-1:0] node16167;
	wire [4-1:0] node16168;
	wire [4-1:0] node16171;
	wire [4-1:0] node16174;
	wire [4-1:0] node16175;
	wire [4-1:0] node16179;
	wire [4-1:0] node16180;
	wire [4-1:0] node16181;
	wire [4-1:0] node16182;
	wire [4-1:0] node16187;
	wire [4-1:0] node16189;
	wire [4-1:0] node16190;
	wire [4-1:0] node16193;
	wire [4-1:0] node16196;
	wire [4-1:0] node16197;
	wire [4-1:0] node16198;
	wire [4-1:0] node16199;
	wire [4-1:0] node16203;
	wire [4-1:0] node16204;
	wire [4-1:0] node16207;
	wire [4-1:0] node16210;
	wire [4-1:0] node16211;
	wire [4-1:0] node16213;
	wire [4-1:0] node16216;
	wire [4-1:0] node16217;
	wire [4-1:0] node16220;
	wire [4-1:0] node16223;
	wire [4-1:0] node16224;
	wire [4-1:0] node16225;
	wire [4-1:0] node16226;
	wire [4-1:0] node16228;
	wire [4-1:0] node16231;
	wire [4-1:0] node16232;
	wire [4-1:0] node16235;
	wire [4-1:0] node16238;
	wire [4-1:0] node16240;
	wire [4-1:0] node16242;
	wire [4-1:0] node16243;
	wire [4-1:0] node16247;
	wire [4-1:0] node16248;
	wire [4-1:0] node16249;
	wire [4-1:0] node16250;
	wire [4-1:0] node16252;
	wire [4-1:0] node16255;
	wire [4-1:0] node16256;
	wire [4-1:0] node16259;
	wire [4-1:0] node16262;
	wire [4-1:0] node16263;
	wire [4-1:0] node16264;
	wire [4-1:0] node16267;
	wire [4-1:0] node16270;
	wire [4-1:0] node16272;
	wire [4-1:0] node16275;
	wire [4-1:0] node16277;
	wire [4-1:0] node16278;
	wire [4-1:0] node16280;
	wire [4-1:0] node16283;
	wire [4-1:0] node16285;
	wire [4-1:0] node16288;
	wire [4-1:0] node16289;
	wire [4-1:0] node16290;
	wire [4-1:0] node16291;
	wire [4-1:0] node16292;
	wire [4-1:0] node16293;
	wire [4-1:0] node16295;
	wire [4-1:0] node16298;
	wire [4-1:0] node16299;
	wire [4-1:0] node16300;
	wire [4-1:0] node16304;
	wire [4-1:0] node16305;
	wire [4-1:0] node16309;
	wire [4-1:0] node16310;
	wire [4-1:0] node16312;
	wire [4-1:0] node16313;
	wire [4-1:0] node16316;
	wire [4-1:0] node16319;
	wire [4-1:0] node16320;
	wire [4-1:0] node16322;
	wire [4-1:0] node16326;
	wire [4-1:0] node16327;
	wire [4-1:0] node16328;
	wire [4-1:0] node16330;
	wire [4-1:0] node16332;
	wire [4-1:0] node16335;
	wire [4-1:0] node16336;
	wire [4-1:0] node16337;
	wire [4-1:0] node16340;
	wire [4-1:0] node16343;
	wire [4-1:0] node16344;
	wire [4-1:0] node16347;
	wire [4-1:0] node16350;
	wire [4-1:0] node16351;
	wire [4-1:0] node16353;
	wire [4-1:0] node16355;
	wire [4-1:0] node16358;
	wire [4-1:0] node16359;
	wire [4-1:0] node16362;
	wire [4-1:0] node16365;
	wire [4-1:0] node16366;
	wire [4-1:0] node16367;
	wire [4-1:0] node16368;
	wire [4-1:0] node16369;
	wire [4-1:0] node16372;
	wire [4-1:0] node16375;
	wire [4-1:0] node16376;
	wire [4-1:0] node16377;
	wire [4-1:0] node16380;
	wire [4-1:0] node16384;
	wire [4-1:0] node16385;
	wire [4-1:0] node16386;
	wire [4-1:0] node16387;
	wire [4-1:0] node16391;
	wire [4-1:0] node16392;
	wire [4-1:0] node16396;
	wire [4-1:0] node16397;
	wire [4-1:0] node16398;
	wire [4-1:0] node16402;
	wire [4-1:0] node16405;
	wire [4-1:0] node16406;
	wire [4-1:0] node16407;
	wire [4-1:0] node16408;
	wire [4-1:0] node16409;
	wire [4-1:0] node16413;
	wire [4-1:0] node16414;
	wire [4-1:0] node16418;
	wire [4-1:0] node16419;
	wire [4-1:0] node16422;
	wire [4-1:0] node16423;
	wire [4-1:0] node16427;
	wire [4-1:0] node16428;
	wire [4-1:0] node16429;
	wire [4-1:0] node16431;
	wire [4-1:0] node16434;
	wire [4-1:0] node16437;
	wire [4-1:0] node16438;
	wire [4-1:0] node16439;
	wire [4-1:0] node16443;
	wire [4-1:0] node16446;
	wire [4-1:0] node16447;
	wire [4-1:0] node16448;
	wire [4-1:0] node16449;
	wire [4-1:0] node16450;
	wire [4-1:0] node16452;
	wire [4-1:0] node16453;
	wire [4-1:0] node16456;
	wire [4-1:0] node16459;
	wire [4-1:0] node16460;
	wire [4-1:0] node16463;
	wire [4-1:0] node16466;
	wire [4-1:0] node16467;
	wire [4-1:0] node16468;
	wire [4-1:0] node16469;
	wire [4-1:0] node16473;
	wire [4-1:0] node16476;
	wire [4-1:0] node16477;
	wire [4-1:0] node16481;
	wire [4-1:0] node16482;
	wire [4-1:0] node16483;
	wire [4-1:0] node16484;
	wire [4-1:0] node16485;
	wire [4-1:0] node16489;
	wire [4-1:0] node16490;
	wire [4-1:0] node16494;
	wire [4-1:0] node16495;
	wire [4-1:0] node16496;
	wire [4-1:0] node16500;
	wire [4-1:0] node16501;
	wire [4-1:0] node16505;
	wire [4-1:0] node16506;
	wire [4-1:0] node16507;
	wire [4-1:0] node16510;
	wire [4-1:0] node16513;
	wire [4-1:0] node16514;
	wire [4-1:0] node16518;
	wire [4-1:0] node16519;
	wire [4-1:0] node16520;
	wire [4-1:0] node16521;
	wire [4-1:0] node16522;
	wire [4-1:0] node16523;
	wire [4-1:0] node16527;
	wire [4-1:0] node16528;
	wire [4-1:0] node16532;
	wire [4-1:0] node16533;
	wire [4-1:0] node16534;
	wire [4-1:0] node16538;
	wire [4-1:0] node16539;
	wire [4-1:0] node16543;
	wire [4-1:0] node16544;
	wire [4-1:0] node16546;
	wire [4-1:0] node16549;
	wire [4-1:0] node16550;
	wire [4-1:0] node16551;
	wire [4-1:0] node16556;
	wire [4-1:0] node16557;
	wire [4-1:0] node16558;
	wire [4-1:0] node16559;
	wire [4-1:0] node16560;
	wire [4-1:0] node16564;
	wire [4-1:0] node16567;
	wire [4-1:0] node16568;
	wire [4-1:0] node16572;
	wire [4-1:0] node16573;
	wire [4-1:0] node16575;
	wire [4-1:0] node16578;
	wire [4-1:0] node16579;
	wire [4-1:0] node16582;
	wire [4-1:0] node16585;
	wire [4-1:0] node16586;
	wire [4-1:0] node16587;
	wire [4-1:0] node16588;
	wire [4-1:0] node16589;
	wire [4-1:0] node16590;
	wire [4-1:0] node16591;
	wire [4-1:0] node16592;
	wire [4-1:0] node16593;
	wire [4-1:0] node16594;
	wire [4-1:0] node16595;
	wire [4-1:0] node16596;
	wire [4-1:0] node16597;
	wire [4-1:0] node16600;
	wire [4-1:0] node16603;
	wire [4-1:0] node16604;
	wire [4-1:0] node16607;
	wire [4-1:0] node16610;
	wire [4-1:0] node16611;
	wire [4-1:0] node16614;
	wire [4-1:0] node16617;
	wire [4-1:0] node16618;
	wire [4-1:0] node16619;
	wire [4-1:0] node16622;
	wire [4-1:0] node16624;
	wire [4-1:0] node16627;
	wire [4-1:0] node16628;
	wire [4-1:0] node16629;
	wire [4-1:0] node16632;
	wire [4-1:0] node16635;
	wire [4-1:0] node16636;
	wire [4-1:0] node16639;
	wire [4-1:0] node16642;
	wire [4-1:0] node16643;
	wire [4-1:0] node16644;
	wire [4-1:0] node16645;
	wire [4-1:0] node16646;
	wire [4-1:0] node16649;
	wire [4-1:0] node16652;
	wire [4-1:0] node16654;
	wire [4-1:0] node16657;
	wire [4-1:0] node16658;
	wire [4-1:0] node16660;
	wire [4-1:0] node16663;
	wire [4-1:0] node16664;
	wire [4-1:0] node16667;
	wire [4-1:0] node16670;
	wire [4-1:0] node16671;
	wire [4-1:0] node16672;
	wire [4-1:0] node16674;
	wire [4-1:0] node16675;
	wire [4-1:0] node16679;
	wire [4-1:0] node16680;
	wire [4-1:0] node16681;
	wire [4-1:0] node16684;
	wire [4-1:0] node16688;
	wire [4-1:0] node16689;
	wire [4-1:0] node16690;
	wire [4-1:0] node16691;
	wire [4-1:0] node16694;
	wire [4-1:0] node16697;
	wire [4-1:0] node16698;
	wire [4-1:0] node16701;
	wire [4-1:0] node16704;
	wire [4-1:0] node16705;
	wire [4-1:0] node16708;
	wire [4-1:0] node16711;
	wire [4-1:0] node16712;
	wire [4-1:0] node16713;
	wire [4-1:0] node16714;
	wire [4-1:0] node16715;
	wire [4-1:0] node16717;
	wire [4-1:0] node16719;
	wire [4-1:0] node16722;
	wire [4-1:0] node16723;
	wire [4-1:0] node16725;
	wire [4-1:0] node16728;
	wire [4-1:0] node16730;
	wire [4-1:0] node16733;
	wire [4-1:0] node16734;
	wire [4-1:0] node16735;
	wire [4-1:0] node16738;
	wire [4-1:0] node16741;
	wire [4-1:0] node16742;
	wire [4-1:0] node16745;
	wire [4-1:0] node16748;
	wire [4-1:0] node16749;
	wire [4-1:0] node16750;
	wire [4-1:0] node16751;
	wire [4-1:0] node16752;
	wire [4-1:0] node16757;
	wire [4-1:0] node16759;
	wire [4-1:0] node16761;
	wire [4-1:0] node16764;
	wire [4-1:0] node16765;
	wire [4-1:0] node16766;
	wire [4-1:0] node16768;
	wire [4-1:0] node16771;
	wire [4-1:0] node16772;
	wire [4-1:0] node16775;
	wire [4-1:0] node16778;
	wire [4-1:0] node16779;
	wire [4-1:0] node16780;
	wire [4-1:0] node16783;
	wire [4-1:0] node16787;
	wire [4-1:0] node16788;
	wire [4-1:0] node16789;
	wire [4-1:0] node16790;
	wire [4-1:0] node16791;
	wire [4-1:0] node16792;
	wire [4-1:0] node16795;
	wire [4-1:0] node16798;
	wire [4-1:0] node16800;
	wire [4-1:0] node16803;
	wire [4-1:0] node16804;
	wire [4-1:0] node16805;
	wire [4-1:0] node16810;
	wire [4-1:0] node16811;
	wire [4-1:0] node16812;
	wire [4-1:0] node16815;
	wire [4-1:0] node16818;
	wire [4-1:0] node16819;
	wire [4-1:0] node16822;
	wire [4-1:0] node16825;
	wire [4-1:0] node16826;
	wire [4-1:0] node16827;
	wire [4-1:0] node16828;
	wire [4-1:0] node16829;
	wire [4-1:0] node16833;
	wire [4-1:0] node16835;
	wire [4-1:0] node16838;
	wire [4-1:0] node16839;
	wire [4-1:0] node16841;
	wire [4-1:0] node16845;
	wire [4-1:0] node16846;
	wire [4-1:0] node16848;
	wire [4-1:0] node16849;
	wire [4-1:0] node16852;
	wire [4-1:0] node16855;
	wire [4-1:0] node16856;
	wire [4-1:0] node16857;
	wire [4-1:0] node16860;
	wire [4-1:0] node16863;
	wire [4-1:0] node16864;
	wire [4-1:0] node16867;
	wire [4-1:0] node16870;
	wire [4-1:0] node16871;
	wire [4-1:0] node16872;
	wire [4-1:0] node16873;
	wire [4-1:0] node16874;
	wire [4-1:0] node16875;
	wire [4-1:0] node16876;
	wire [4-1:0] node16877;
	wire [4-1:0] node16882;
	wire [4-1:0] node16883;
	wire [4-1:0] node16887;
	wire [4-1:0] node16888;
	wire [4-1:0] node16889;
	wire [4-1:0] node16894;
	wire [4-1:0] node16895;
	wire [4-1:0] node16896;
	wire [4-1:0] node16897;
	wire [4-1:0] node16898;
	wire [4-1:0] node16902;
	wire [4-1:0] node16903;
	wire [4-1:0] node16907;
	wire [4-1:0] node16908;
	wire [4-1:0] node16912;
	wire [4-1:0] node16913;
	wire [4-1:0] node16915;
	wire [4-1:0] node16916;
	wire [4-1:0] node16920;
	wire [4-1:0] node16923;
	wire [4-1:0] node16924;
	wire [4-1:0] node16925;
	wire [4-1:0] node16926;
	wire [4-1:0] node16927;
	wire [4-1:0] node16930;
	wire [4-1:0] node16933;
	wire [4-1:0] node16934;
	wire [4-1:0] node16936;
	wire [4-1:0] node16939;
	wire [4-1:0] node16940;
	wire [4-1:0] node16944;
	wire [4-1:0] node16945;
	wire [4-1:0] node16948;
	wire [4-1:0] node16951;
	wire [4-1:0] node16952;
	wire [4-1:0] node16953;
	wire [4-1:0] node16955;
	wire [4-1:0] node16956;
	wire [4-1:0] node16960;
	wire [4-1:0] node16961;
	wire [4-1:0] node16962;
	wire [4-1:0] node16966;
	wire [4-1:0] node16969;
	wire [4-1:0] node16970;
	wire [4-1:0] node16971;
	wire [4-1:0] node16973;
	wire [4-1:0] node16976;
	wire [4-1:0] node16977;
	wire [4-1:0] node16981;
	wire [4-1:0] node16982;
	wire [4-1:0] node16986;
	wire [4-1:0] node16987;
	wire [4-1:0] node16988;
	wire [4-1:0] node16989;
	wire [4-1:0] node16990;
	wire [4-1:0] node16992;
	wire [4-1:0] node16995;
	wire [4-1:0] node16996;
	wire [4-1:0] node16997;
	wire [4-1:0] node17000;
	wire [4-1:0] node17003;
	wire [4-1:0] node17004;
	wire [4-1:0] node17007;
	wire [4-1:0] node17010;
	wire [4-1:0] node17011;
	wire [4-1:0] node17012;
	wire [4-1:0] node17015;
	wire [4-1:0] node17018;
	wire [4-1:0] node17019;
	wire [4-1:0] node17022;
	wire [4-1:0] node17025;
	wire [4-1:0] node17026;
	wire [4-1:0] node17027;
	wire [4-1:0] node17028;
	wire [4-1:0] node17030;
	wire [4-1:0] node17034;
	wire [4-1:0] node17036;
	wire [4-1:0] node17039;
	wire [4-1:0] node17040;
	wire [4-1:0] node17042;
	wire [4-1:0] node17044;
	wire [4-1:0] node17047;
	wire [4-1:0] node17049;
	wire [4-1:0] node17052;
	wire [4-1:0] node17053;
	wire [4-1:0] node17054;
	wire [4-1:0] node17055;
	wire [4-1:0] node17056;
	wire [4-1:0] node17060;
	wire [4-1:0] node17061;
	wire [4-1:0] node17062;
	wire [4-1:0] node17065;
	wire [4-1:0] node17068;
	wire [4-1:0] node17069;
	wire [4-1:0] node17072;
	wire [4-1:0] node17075;
	wire [4-1:0] node17076;
	wire [4-1:0] node17077;
	wire [4-1:0] node17080;
	wire [4-1:0] node17083;
	wire [4-1:0] node17084;
	wire [4-1:0] node17087;
	wire [4-1:0] node17090;
	wire [4-1:0] node17091;
	wire [4-1:0] node17092;
	wire [4-1:0] node17093;
	wire [4-1:0] node17094;
	wire [4-1:0] node17097;
	wire [4-1:0] node17100;
	wire [4-1:0] node17101;
	wire [4-1:0] node17104;
	wire [4-1:0] node17107;
	wire [4-1:0] node17108;
	wire [4-1:0] node17111;
	wire [4-1:0] node17114;
	wire [4-1:0] node17115;
	wire [4-1:0] node17116;
	wire [4-1:0] node17117;
	wire [4-1:0] node17120;
	wire [4-1:0] node17123;
	wire [4-1:0] node17124;
	wire [4-1:0] node17127;
	wire [4-1:0] node17130;
	wire [4-1:0] node17131;
	wire [4-1:0] node17134;
	wire [4-1:0] node17135;
	wire [4-1:0] node17139;
	wire [4-1:0] node17140;
	wire [4-1:0] node17141;
	wire [4-1:0] node17142;
	wire [4-1:0] node17143;
	wire [4-1:0] node17144;
	wire [4-1:0] node17145;
	wire [4-1:0] node17146;
	wire [4-1:0] node17147;
	wire [4-1:0] node17152;
	wire [4-1:0] node17153;
	wire [4-1:0] node17157;
	wire [4-1:0] node17159;
	wire [4-1:0] node17162;
	wire [4-1:0] node17163;
	wire [4-1:0] node17164;
	wire [4-1:0] node17166;
	wire [4-1:0] node17167;
	wire [4-1:0] node17171;
	wire [4-1:0] node17172;
	wire [4-1:0] node17175;
	wire [4-1:0] node17178;
	wire [4-1:0] node17179;
	wire [4-1:0] node17181;
	wire [4-1:0] node17182;
	wire [4-1:0] node17185;
	wire [4-1:0] node17188;
	wire [4-1:0] node17189;
	wire [4-1:0] node17192;
	wire [4-1:0] node17195;
	wire [4-1:0] node17196;
	wire [4-1:0] node17197;
	wire [4-1:0] node17198;
	wire [4-1:0] node17199;
	wire [4-1:0] node17203;
	wire [4-1:0] node17204;
	wire [4-1:0] node17208;
	wire [4-1:0] node17209;
	wire [4-1:0] node17211;
	wire [4-1:0] node17214;
	wire [4-1:0] node17215;
	wire [4-1:0] node17219;
	wire [4-1:0] node17220;
	wire [4-1:0] node17221;
	wire [4-1:0] node17222;
	wire [4-1:0] node17223;
	wire [4-1:0] node17226;
	wire [4-1:0] node17229;
	wire [4-1:0] node17230;
	wire [4-1:0] node17233;
	wire [4-1:0] node17236;
	wire [4-1:0] node17237;
	wire [4-1:0] node17240;
	wire [4-1:0] node17243;
	wire [4-1:0] node17244;
	wire [4-1:0] node17245;
	wire [4-1:0] node17249;
	wire [4-1:0] node17250;
	wire [4-1:0] node17251;
	wire [4-1:0] node17256;
	wire [4-1:0] node17257;
	wire [4-1:0] node17258;
	wire [4-1:0] node17259;
	wire [4-1:0] node17260;
	wire [4-1:0] node17261;
	wire [4-1:0] node17265;
	wire [4-1:0] node17266;
	wire [4-1:0] node17270;
	wire [4-1:0] node17271;
	wire [4-1:0] node17272;
	wire [4-1:0] node17276;
	wire [4-1:0] node17277;
	wire [4-1:0] node17281;
	wire [4-1:0] node17282;
	wire [4-1:0] node17283;
	wire [4-1:0] node17284;
	wire [4-1:0] node17285;
	wire [4-1:0] node17288;
	wire [4-1:0] node17292;
	wire [4-1:0] node17293;
	wire [4-1:0] node17297;
	wire [4-1:0] node17298;
	wire [4-1:0] node17299;
	wire [4-1:0] node17300;
	wire [4-1:0] node17304;
	wire [4-1:0] node17307;
	wire [4-1:0] node17309;
	wire [4-1:0] node17310;
	wire [4-1:0] node17314;
	wire [4-1:0] node17315;
	wire [4-1:0] node17316;
	wire [4-1:0] node17317;
	wire [4-1:0] node17318;
	wire [4-1:0] node17322;
	wire [4-1:0] node17323;
	wire [4-1:0] node17327;
	wire [4-1:0] node17328;
	wire [4-1:0] node17329;
	wire [4-1:0] node17333;
	wire [4-1:0] node17334;
	wire [4-1:0] node17338;
	wire [4-1:0] node17339;
	wire [4-1:0] node17340;
	wire [4-1:0] node17341;
	wire [4-1:0] node17342;
	wire [4-1:0] node17346;
	wire [4-1:0] node17347;
	wire [4-1:0] node17351;
	wire [4-1:0] node17354;
	wire [4-1:0] node17355;
	wire [4-1:0] node17357;
	wire [4-1:0] node17358;
	wire [4-1:0] node17361;
	wire [4-1:0] node17364;
	wire [4-1:0] node17365;
	wire [4-1:0] node17369;
	wire [4-1:0] node17370;
	wire [4-1:0] node17371;
	wire [4-1:0] node17372;
	wire [4-1:0] node17373;
	wire [4-1:0] node17374;
	wire [4-1:0] node17376;
	wire [4-1:0] node17377;
	wire [4-1:0] node17380;
	wire [4-1:0] node17384;
	wire [4-1:0] node17385;
	wire [4-1:0] node17387;
	wire [4-1:0] node17388;
	wire [4-1:0] node17392;
	wire [4-1:0] node17393;
	wire [4-1:0] node17395;
	wire [4-1:0] node17399;
	wire [4-1:0] node17400;
	wire [4-1:0] node17401;
	wire [4-1:0] node17402;
	wire [4-1:0] node17403;
	wire [4-1:0] node17406;
	wire [4-1:0] node17409;
	wire [4-1:0] node17411;
	wire [4-1:0] node17414;
	wire [4-1:0] node17415;
	wire [4-1:0] node17418;
	wire [4-1:0] node17421;
	wire [4-1:0] node17422;
	wire [4-1:0] node17423;
	wire [4-1:0] node17426;
	wire [4-1:0] node17429;
	wire [4-1:0] node17430;
	wire [4-1:0] node17432;
	wire [4-1:0] node17436;
	wire [4-1:0] node17437;
	wire [4-1:0] node17438;
	wire [4-1:0] node17439;
	wire [4-1:0] node17441;
	wire [4-1:0] node17444;
	wire [4-1:0] node17446;
	wire [4-1:0] node17447;
	wire [4-1:0] node17450;
	wire [4-1:0] node17453;
	wire [4-1:0] node17454;
	wire [4-1:0] node17457;
	wire [4-1:0] node17458;
	wire [4-1:0] node17459;
	wire [4-1:0] node17462;
	wire [4-1:0] node17465;
	wire [4-1:0] node17466;
	wire [4-1:0] node17470;
	wire [4-1:0] node17471;
	wire [4-1:0] node17472;
	wire [4-1:0] node17473;
	wire [4-1:0] node17476;
	wire [4-1:0] node17479;
	wire [4-1:0] node17480;
	wire [4-1:0] node17483;
	wire [4-1:0] node17486;
	wire [4-1:0] node17487;
	wire [4-1:0] node17488;
	wire [4-1:0] node17492;
	wire [4-1:0] node17494;
	wire [4-1:0] node17496;
	wire [4-1:0] node17499;
	wire [4-1:0] node17500;
	wire [4-1:0] node17501;
	wire [4-1:0] node17502;
	wire [4-1:0] node17503;
	wire [4-1:0] node17506;
	wire [4-1:0] node17509;
	wire [4-1:0] node17510;
	wire [4-1:0] node17511;
	wire [4-1:0] node17514;
	wire [4-1:0] node17517;
	wire [4-1:0] node17518;
	wire [4-1:0] node17521;
	wire [4-1:0] node17524;
	wire [4-1:0] node17525;
	wire [4-1:0] node17526;
	wire [4-1:0] node17529;
	wire [4-1:0] node17532;
	wire [4-1:0] node17533;
	wire [4-1:0] node17534;
	wire [4-1:0] node17535;
	wire [4-1:0] node17538;
	wire [4-1:0] node17542;
	wire [4-1:0] node17543;
	wire [4-1:0] node17546;
	wire [4-1:0] node17549;
	wire [4-1:0] node17550;
	wire [4-1:0] node17551;
	wire [4-1:0] node17552;
	wire [4-1:0] node17555;
	wire [4-1:0] node17558;
	wire [4-1:0] node17559;
	wire [4-1:0] node17560;
	wire [4-1:0] node17561;
	wire [4-1:0] node17565;
	wire [4-1:0] node17566;
	wire [4-1:0] node17569;
	wire [4-1:0] node17572;
	wire [4-1:0] node17574;
	wire [4-1:0] node17577;
	wire [4-1:0] node17578;
	wire [4-1:0] node17579;
	wire [4-1:0] node17582;
	wire [4-1:0] node17585;
	wire [4-1:0] node17586;
	wire [4-1:0] node17587;
	wire [4-1:0] node17588;
	wire [4-1:0] node17591;
	wire [4-1:0] node17595;
	wire [4-1:0] node17596;
	wire [4-1:0] node17597;
	wire [4-1:0] node17601;
	wire [4-1:0] node17604;
	wire [4-1:0] node17605;
	wire [4-1:0] node17606;
	wire [4-1:0] node17607;
	wire [4-1:0] node17608;
	wire [4-1:0] node17609;
	wire [4-1:0] node17610;
	wire [4-1:0] node17611;
	wire [4-1:0] node17612;
	wire [4-1:0] node17615;
	wire [4-1:0] node17618;
	wire [4-1:0] node17620;
	wire [4-1:0] node17621;
	wire [4-1:0] node17624;
	wire [4-1:0] node17627;
	wire [4-1:0] node17628;
	wire [4-1:0] node17629;
	wire [4-1:0] node17632;
	wire [4-1:0] node17635;
	wire [4-1:0] node17636;
	wire [4-1:0] node17638;
	wire [4-1:0] node17641;
	wire [4-1:0] node17644;
	wire [4-1:0] node17645;
	wire [4-1:0] node17646;
	wire [4-1:0] node17647;
	wire [4-1:0] node17651;
	wire [4-1:0] node17652;
	wire [4-1:0] node17653;
	wire [4-1:0] node17658;
	wire [4-1:0] node17659;
	wire [4-1:0] node17660;
	wire [4-1:0] node17663;
	wire [4-1:0] node17666;
	wire [4-1:0] node17667;
	wire [4-1:0] node17671;
	wire [4-1:0] node17672;
	wire [4-1:0] node17673;
	wire [4-1:0] node17674;
	wire [4-1:0] node17675;
	wire [4-1:0] node17679;
	wire [4-1:0] node17680;
	wire [4-1:0] node17681;
	wire [4-1:0] node17684;
	wire [4-1:0] node17688;
	wire [4-1:0] node17689;
	wire [4-1:0] node17690;
	wire [4-1:0] node17691;
	wire [4-1:0] node17694;
	wire [4-1:0] node17697;
	wire [4-1:0] node17698;
	wire [4-1:0] node17702;
	wire [4-1:0] node17703;
	wire [4-1:0] node17707;
	wire [4-1:0] node17708;
	wire [4-1:0] node17709;
	wire [4-1:0] node17710;
	wire [4-1:0] node17713;
	wire [4-1:0] node17716;
	wire [4-1:0] node17718;
	wire [4-1:0] node17721;
	wire [4-1:0] node17722;
	wire [4-1:0] node17723;
	wire [4-1:0] node17726;
	wire [4-1:0] node17729;
	wire [4-1:0] node17730;
	wire [4-1:0] node17733;
	wire [4-1:0] node17736;
	wire [4-1:0] node17737;
	wire [4-1:0] node17738;
	wire [4-1:0] node17739;
	wire [4-1:0] node17740;
	wire [4-1:0] node17742;
	wire [4-1:0] node17743;
	wire [4-1:0] node17746;
	wire [4-1:0] node17749;
	wire [4-1:0] node17750;
	wire [4-1:0] node17751;
	wire [4-1:0] node17755;
	wire [4-1:0] node17757;
	wire [4-1:0] node17760;
	wire [4-1:0] node17761;
	wire [4-1:0] node17762;
	wire [4-1:0] node17766;
	wire [4-1:0] node17767;
	wire [4-1:0] node17770;
	wire [4-1:0] node17771;
	wire [4-1:0] node17775;
	wire [4-1:0] node17776;
	wire [4-1:0] node17777;
	wire [4-1:0] node17778;
	wire [4-1:0] node17779;
	wire [4-1:0] node17783;
	wire [4-1:0] node17784;
	wire [4-1:0] node17787;
	wire [4-1:0] node17790;
	wire [4-1:0] node17791;
	wire [4-1:0] node17792;
	wire [4-1:0] node17795;
	wire [4-1:0] node17798;
	wire [4-1:0] node17799;
	wire [4-1:0] node17802;
	wire [4-1:0] node17805;
	wire [4-1:0] node17806;
	wire [4-1:0] node17808;
	wire [4-1:0] node17809;
	wire [4-1:0] node17812;
	wire [4-1:0] node17816;
	wire [4-1:0] node17817;
	wire [4-1:0] node17818;
	wire [4-1:0] node17819;
	wire [4-1:0] node17820;
	wire [4-1:0] node17822;
	wire [4-1:0] node17826;
	wire [4-1:0] node17827;
	wire [4-1:0] node17828;
	wire [4-1:0] node17832;
	wire [4-1:0] node17833;
	wire [4-1:0] node17836;
	wire [4-1:0] node17839;
	wire [4-1:0] node17840;
	wire [4-1:0] node17841;
	wire [4-1:0] node17845;
	wire [4-1:0] node17846;
	wire [4-1:0] node17849;
	wire [4-1:0] node17852;
	wire [4-1:0] node17853;
	wire [4-1:0] node17854;
	wire [4-1:0] node17855;
	wire [4-1:0] node17856;
	wire [4-1:0] node17859;
	wire [4-1:0] node17862;
	wire [4-1:0] node17865;
	wire [4-1:0] node17866;
	wire [4-1:0] node17869;
	wire [4-1:0] node17872;
	wire [4-1:0] node17873;
	wire [4-1:0] node17874;
	wire [4-1:0] node17877;
	wire [4-1:0] node17878;
	wire [4-1:0] node17882;
	wire [4-1:0] node17883;
	wire [4-1:0] node17884;
	wire [4-1:0] node17887;
	wire [4-1:0] node17890;
	wire [4-1:0] node17891;
	wire [4-1:0] node17894;
	wire [4-1:0] node17897;
	wire [4-1:0] node17898;
	wire [4-1:0] node17899;
	wire [4-1:0] node17900;
	wire [4-1:0] node17901;
	wire [4-1:0] node17902;
	wire [4-1:0] node17904;
	wire [4-1:0] node17905;
	wire [4-1:0] node17908;
	wire [4-1:0] node17911;
	wire [4-1:0] node17912;
	wire [4-1:0] node17913;
	wire [4-1:0] node17917;
	wire [4-1:0] node17918;
	wire [4-1:0] node17921;
	wire [4-1:0] node17924;
	wire [4-1:0] node17925;
	wire [4-1:0] node17929;
	wire [4-1:0] node17930;
	wire [4-1:0] node17931;
	wire [4-1:0] node17932;
	wire [4-1:0] node17933;
	wire [4-1:0] node17936;
	wire [4-1:0] node17939;
	wire [4-1:0] node17940;
	wire [4-1:0] node17943;
	wire [4-1:0] node17946;
	wire [4-1:0] node17947;
	wire [4-1:0] node17951;
	wire [4-1:0] node17952;
	wire [4-1:0] node17954;
	wire [4-1:0] node17957;
	wire [4-1:0] node17958;
	wire [4-1:0] node17959;
	wire [4-1:0] node17963;
	wire [4-1:0] node17964;
	wire [4-1:0] node17968;
	wire [4-1:0] node17969;
	wire [4-1:0] node17970;
	wire [4-1:0] node17971;
	wire [4-1:0] node17972;
	wire [4-1:0] node17976;
	wire [4-1:0] node17977;
	wire [4-1:0] node17980;
	wire [4-1:0] node17983;
	wire [4-1:0] node17984;
	wire [4-1:0] node17987;
	wire [4-1:0] node17990;
	wire [4-1:0] node17991;
	wire [4-1:0] node17992;
	wire [4-1:0] node17993;
	wire [4-1:0] node17995;
	wire [4-1:0] node17998;
	wire [4-1:0] node17999;
	wire [4-1:0] node18002;
	wire [4-1:0] node18005;
	wire [4-1:0] node18006;
	wire [4-1:0] node18007;
	wire [4-1:0] node18010;
	wire [4-1:0] node18014;
	wire [4-1:0] node18015;
	wire [4-1:0] node18016;
	wire [4-1:0] node18017;
	wire [4-1:0] node18020;
	wire [4-1:0] node18023;
	wire [4-1:0] node18024;
	wire [4-1:0] node18027;
	wire [4-1:0] node18030;
	wire [4-1:0] node18031;
	wire [4-1:0] node18033;
	wire [4-1:0] node18036;
	wire [4-1:0] node18037;
	wire [4-1:0] node18040;
	wire [4-1:0] node18043;
	wire [4-1:0] node18044;
	wire [4-1:0] node18045;
	wire [4-1:0] node18046;
	wire [4-1:0] node18047;
	wire [4-1:0] node18048;
	wire [4-1:0] node18051;
	wire [4-1:0] node18054;
	wire [4-1:0] node18055;
	wire [4-1:0] node18056;
	wire [4-1:0] node18059;
	wire [4-1:0] node18062;
	wire [4-1:0] node18063;
	wire [4-1:0] node18066;
	wire [4-1:0] node18069;
	wire [4-1:0] node18070;
	wire [4-1:0] node18073;
	wire [4-1:0] node18076;
	wire [4-1:0] node18077;
	wire [4-1:0] node18078;
	wire [4-1:0] node18080;
	wire [4-1:0] node18081;
	wire [4-1:0] node18086;
	wire [4-1:0] node18087;
	wire [4-1:0] node18088;
	wire [4-1:0] node18089;
	wire [4-1:0] node18092;
	wire [4-1:0] node18095;
	wire [4-1:0] node18096;
	wire [4-1:0] node18099;
	wire [4-1:0] node18102;
	wire [4-1:0] node18103;
	wire [4-1:0] node18106;
	wire [4-1:0] node18109;
	wire [4-1:0] node18110;
	wire [4-1:0] node18111;
	wire [4-1:0] node18112;
	wire [4-1:0] node18113;
	wire [4-1:0] node18116;
	wire [4-1:0] node18119;
	wire [4-1:0] node18120;
	wire [4-1:0] node18123;
	wire [4-1:0] node18126;
	wire [4-1:0] node18127;
	wire [4-1:0] node18128;
	wire [4-1:0] node18131;
	wire [4-1:0] node18134;
	wire [4-1:0] node18135;
	wire [4-1:0] node18137;
	wire [4-1:0] node18140;
	wire [4-1:0] node18141;
	wire [4-1:0] node18145;
	wire [4-1:0] node18146;
	wire [4-1:0] node18147;
	wire [4-1:0] node18148;
	wire [4-1:0] node18149;
	wire [4-1:0] node18152;
	wire [4-1:0] node18156;
	wire [4-1:0] node18158;
	wire [4-1:0] node18161;
	wire [4-1:0] node18162;
	wire [4-1:0] node18163;
	wire [4-1:0] node18167;
	wire [4-1:0] node18168;
	wire [4-1:0] node18172;
	wire [4-1:0] node18173;
	wire [4-1:0] node18174;
	wire [4-1:0] node18175;
	wire [4-1:0] node18176;
	wire [4-1:0] node18177;
	wire [4-1:0] node18178;
	wire [4-1:0] node18179;
	wire [4-1:0] node18183;
	wire [4-1:0] node18184;
	wire [4-1:0] node18188;
	wire [4-1:0] node18189;
	wire [4-1:0] node18190;
	wire [4-1:0] node18194;
	wire [4-1:0] node18195;
	wire [4-1:0] node18199;
	wire [4-1:0] node18200;
	wire [4-1:0] node18201;
	wire [4-1:0] node18202;
	wire [4-1:0] node18203;
	wire [4-1:0] node18206;
	wire [4-1:0] node18210;
	wire [4-1:0] node18211;
	wire [4-1:0] node18212;
	wire [4-1:0] node18217;
	wire [4-1:0] node18218;
	wire [4-1:0] node18219;
	wire [4-1:0] node18220;
	wire [4-1:0] node18225;
	wire [4-1:0] node18226;
	wire [4-1:0] node18227;
	wire [4-1:0] node18232;
	wire [4-1:0] node18233;
	wire [4-1:0] node18234;
	wire [4-1:0] node18235;
	wire [4-1:0] node18236;
	wire [4-1:0] node18240;
	wire [4-1:0] node18241;
	wire [4-1:0] node18245;
	wire [4-1:0] node18246;
	wire [4-1:0] node18247;
	wire [4-1:0] node18251;
	wire [4-1:0] node18252;
	wire [4-1:0] node18256;
	wire [4-1:0] node18257;
	wire [4-1:0] node18258;
	wire [4-1:0] node18259;
	wire [4-1:0] node18260;
	wire [4-1:0] node18264;
	wire [4-1:0] node18265;
	wire [4-1:0] node18269;
	wire [4-1:0] node18270;
	wire [4-1:0] node18274;
	wire [4-1:0] node18275;
	wire [4-1:0] node18277;
	wire [4-1:0] node18278;
	wire [4-1:0] node18281;
	wire [4-1:0] node18284;
	wire [4-1:0] node18285;
	wire [4-1:0] node18288;
	wire [4-1:0] node18291;
	wire [4-1:0] node18292;
	wire [4-1:0] node18293;
	wire [4-1:0] node18294;
	wire [4-1:0] node18295;
	wire [4-1:0] node18296;
	wire [4-1:0] node18300;
	wire [4-1:0] node18303;
	wire [4-1:0] node18305;
	wire [4-1:0] node18306;
	wire [4-1:0] node18310;
	wire [4-1:0] node18311;
	wire [4-1:0] node18312;
	wire [4-1:0] node18313;
	wire [4-1:0] node18314;
	wire [4-1:0] node18317;
	wire [4-1:0] node18321;
	wire [4-1:0] node18322;
	wire [4-1:0] node18325;
	wire [4-1:0] node18328;
	wire [4-1:0] node18329;
	wire [4-1:0] node18330;
	wire [4-1:0] node18332;
	wire [4-1:0] node18335;
	wire [4-1:0] node18337;
	wire [4-1:0] node18340;
	wire [4-1:0] node18341;
	wire [4-1:0] node18344;
	wire [4-1:0] node18347;
	wire [4-1:0] node18348;
	wire [4-1:0] node18349;
	wire [4-1:0] node18350;
	wire [4-1:0] node18351;
	wire [4-1:0] node18352;
	wire [4-1:0] node18355;
	wire [4-1:0] node18358;
	wire [4-1:0] node18360;
	wire [4-1:0] node18363;
	wire [4-1:0] node18364;
	wire [4-1:0] node18368;
	wire [4-1:0] node18369;
	wire [4-1:0] node18371;
	wire [4-1:0] node18373;
	wire [4-1:0] node18376;
	wire [4-1:0] node18377;
	wire [4-1:0] node18378;
	wire [4-1:0] node18382;
	wire [4-1:0] node18383;
	wire [4-1:0] node18386;
	wire [4-1:0] node18389;
	wire [4-1:0] node18390;
	wire [4-1:0] node18391;
	wire [4-1:0] node18393;
	wire [4-1:0] node18394;
	wire [4-1:0] node18397;
	wire [4-1:0] node18400;
	wire [4-1:0] node18401;
	wire [4-1:0] node18402;
	wire [4-1:0] node18407;
	wire [4-1:0] node18408;
	wire [4-1:0] node18409;
	wire [4-1:0] node18410;
	wire [4-1:0] node18413;
	wire [4-1:0] node18417;
	wire [4-1:0] node18418;
	wire [4-1:0] node18419;
	wire [4-1:0] node18423;
	wire [4-1:0] node18426;
	wire [4-1:0] node18427;
	wire [4-1:0] node18428;
	wire [4-1:0] node18429;
	wire [4-1:0] node18430;
	wire [4-1:0] node18431;
	wire [4-1:0] node18432;
	wire [4-1:0] node18436;
	wire [4-1:0] node18437;
	wire [4-1:0] node18440;
	wire [4-1:0] node18443;
	wire [4-1:0] node18445;
	wire [4-1:0] node18446;
	wire [4-1:0] node18448;
	wire [4-1:0] node18451;
	wire [4-1:0] node18453;
	wire [4-1:0] node18456;
	wire [4-1:0] node18457;
	wire [4-1:0] node18458;
	wire [4-1:0] node18460;
	wire [4-1:0] node18461;
	wire [4-1:0] node18464;
	wire [4-1:0] node18467;
	wire [4-1:0] node18468;
	wire [4-1:0] node18471;
	wire [4-1:0] node18474;
	wire [4-1:0] node18475;
	wire [4-1:0] node18477;
	wire [4-1:0] node18478;
	wire [4-1:0] node18481;
	wire [4-1:0] node18484;
	wire [4-1:0] node18487;
	wire [4-1:0] node18488;
	wire [4-1:0] node18489;
	wire [4-1:0] node18490;
	wire [4-1:0] node18491;
	wire [4-1:0] node18492;
	wire [4-1:0] node18495;
	wire [4-1:0] node18498;
	wire [4-1:0] node18499;
	wire [4-1:0] node18502;
	wire [4-1:0] node18505;
	wire [4-1:0] node18506;
	wire [4-1:0] node18510;
	wire [4-1:0] node18511;
	wire [4-1:0] node18512;
	wire [4-1:0] node18513;
	wire [4-1:0] node18516;
	wire [4-1:0] node18520;
	wire [4-1:0] node18521;
	wire [4-1:0] node18523;
	wire [4-1:0] node18526;
	wire [4-1:0] node18528;
	wire [4-1:0] node18531;
	wire [4-1:0] node18532;
	wire [4-1:0] node18533;
	wire [4-1:0] node18534;
	wire [4-1:0] node18537;
	wire [4-1:0] node18540;
	wire [4-1:0] node18541;
	wire [4-1:0] node18544;
	wire [4-1:0] node18547;
	wire [4-1:0] node18548;
	wire [4-1:0] node18550;
	wire [4-1:0] node18551;
	wire [4-1:0] node18554;
	wire [4-1:0] node18557;
	wire [4-1:0] node18558;
	wire [4-1:0] node18559;
	wire [4-1:0] node18562;
	wire [4-1:0] node18566;
	wire [4-1:0] node18567;
	wire [4-1:0] node18568;
	wire [4-1:0] node18569;
	wire [4-1:0] node18570;
	wire [4-1:0] node18573;
	wire [4-1:0] node18576;
	wire [4-1:0] node18577;
	wire [4-1:0] node18579;
	wire [4-1:0] node18582;
	wire [4-1:0] node18584;
	wire [4-1:0] node18587;
	wire [4-1:0] node18588;
	wire [4-1:0] node18589;
	wire [4-1:0] node18591;
	wire [4-1:0] node18592;
	wire [4-1:0] node18595;
	wire [4-1:0] node18598;
	wire [4-1:0] node18599;
	wire [4-1:0] node18603;
	wire [4-1:0] node18604;
	wire [4-1:0] node18605;
	wire [4-1:0] node18607;
	wire [4-1:0] node18611;
	wire [4-1:0] node18612;
	wire [4-1:0] node18615;
	wire [4-1:0] node18618;
	wire [4-1:0] node18619;
	wire [4-1:0] node18620;
	wire [4-1:0] node18621;
	wire [4-1:0] node18623;
	wire [4-1:0] node18624;
	wire [4-1:0] node18627;
	wire [4-1:0] node18630;
	wire [4-1:0] node18631;
	wire [4-1:0] node18634;
	wire [4-1:0] node18637;
	wire [4-1:0] node18638;
	wire [4-1:0] node18639;
	wire [4-1:0] node18642;
	wire [4-1:0] node18645;
	wire [4-1:0] node18646;
	wire [4-1:0] node18648;
	wire [4-1:0] node18652;
	wire [4-1:0] node18653;
	wire [4-1:0] node18654;
	wire [4-1:0] node18655;
	wire [4-1:0] node18659;
	wire [4-1:0] node18660;
	wire [4-1:0] node18663;
	wire [4-1:0] node18666;
	wire [4-1:0] node18667;
	wire [4-1:0] node18670;
	wire [4-1:0] node18671;
	wire [4-1:0] node18674;
	wire [4-1:0] node18677;
	wire [4-1:0] node18678;
	wire [4-1:0] node18679;
	wire [4-1:0] node18680;
	wire [4-1:0] node18681;
	wire [4-1:0] node18682;
	wire [4-1:0] node18683;
	wire [4-1:0] node18684;
	wire [4-1:0] node18685;
	wire [4-1:0] node18686;
	wire [4-1:0] node18690;
	wire [4-1:0] node18691;
	wire [4-1:0] node18695;
	wire [4-1:0] node18696;
	wire [4-1:0] node18699;
	wire [4-1:0] node18700;
	wire [4-1:0] node18704;
	wire [4-1:0] node18705;
	wire [4-1:0] node18706;
	wire [4-1:0] node18707;
	wire [4-1:0] node18710;
	wire [4-1:0] node18711;
	wire [4-1:0] node18715;
	wire [4-1:0] node18718;
	wire [4-1:0] node18720;
	wire [4-1:0] node18721;
	wire [4-1:0] node18722;
	wire [4-1:0] node18725;
	wire [4-1:0] node18728;
	wire [4-1:0] node18729;
	wire [4-1:0] node18732;
	wire [4-1:0] node18735;
	wire [4-1:0] node18736;
	wire [4-1:0] node18737;
	wire [4-1:0] node18738;
	wire [4-1:0] node18739;
	wire [4-1:0] node18742;
	wire [4-1:0] node18745;
	wire [4-1:0] node18747;
	wire [4-1:0] node18748;
	wire [4-1:0] node18751;
	wire [4-1:0] node18754;
	wire [4-1:0] node18755;
	wire [4-1:0] node18756;
	wire [4-1:0] node18759;
	wire [4-1:0] node18762;
	wire [4-1:0] node18764;
	wire [4-1:0] node18767;
	wire [4-1:0] node18768;
	wire [4-1:0] node18769;
	wire [4-1:0] node18771;
	wire [4-1:0] node18774;
	wire [4-1:0] node18777;
	wire [4-1:0] node18778;
	wire [4-1:0] node18779;
	wire [4-1:0] node18780;
	wire [4-1:0] node18783;
	wire [4-1:0] node18787;
	wire [4-1:0] node18788;
	wire [4-1:0] node18789;
	wire [4-1:0] node18792;
	wire [4-1:0] node18796;
	wire [4-1:0] node18797;
	wire [4-1:0] node18798;
	wire [4-1:0] node18799;
	wire [4-1:0] node18801;
	wire [4-1:0] node18802;
	wire [4-1:0] node18803;
	wire [4-1:0] node18806;
	wire [4-1:0] node18809;
	wire [4-1:0] node18810;
	wire [4-1:0] node18813;
	wire [4-1:0] node18816;
	wire [4-1:0] node18817;
	wire [4-1:0] node18818;
	wire [4-1:0] node18821;
	wire [4-1:0] node18824;
	wire [4-1:0] node18825;
	wire [4-1:0] node18828;
	wire [4-1:0] node18831;
	wire [4-1:0] node18832;
	wire [4-1:0] node18833;
	wire [4-1:0] node18834;
	wire [4-1:0] node18835;
	wire [4-1:0] node18839;
	wire [4-1:0] node18840;
	wire [4-1:0] node18844;
	wire [4-1:0] node18847;
	wire [4-1:0] node18848;
	wire [4-1:0] node18849;
	wire [4-1:0] node18850;
	wire [4-1:0] node18853;
	wire [4-1:0] node18857;
	wire [4-1:0] node18858;
	wire [4-1:0] node18859;
	wire [4-1:0] node18862;
	wire [4-1:0] node18866;
	wire [4-1:0] node18867;
	wire [4-1:0] node18868;
	wire [4-1:0] node18869;
	wire [4-1:0] node18870;
	wire [4-1:0] node18871;
	wire [4-1:0] node18874;
	wire [4-1:0] node18877;
	wire [4-1:0] node18879;
	wire [4-1:0] node18883;
	wire [4-1:0] node18884;
	wire [4-1:0] node18885;
	wire [4-1:0] node18886;
	wire [4-1:0] node18889;
	wire [4-1:0] node18893;
	wire [4-1:0] node18894;
	wire [4-1:0] node18897;
	wire [4-1:0] node18900;
	wire [4-1:0] node18901;
	wire [4-1:0] node18902;
	wire [4-1:0] node18903;
	wire [4-1:0] node18904;
	wire [4-1:0] node18909;
	wire [4-1:0] node18911;
	wire [4-1:0] node18914;
	wire [4-1:0] node18915;
	wire [4-1:0] node18916;
	wire [4-1:0] node18918;
	wire [4-1:0] node18921;
	wire [4-1:0] node18923;
	wire [4-1:0] node18926;
	wire [4-1:0] node18927;
	wire [4-1:0] node18930;
	wire [4-1:0] node18933;
	wire [4-1:0] node18934;
	wire [4-1:0] node18935;
	wire [4-1:0] node18936;
	wire [4-1:0] node18937;
	wire [4-1:0] node18938;
	wire [4-1:0] node18939;
	wire [4-1:0] node18943;
	wire [4-1:0] node18944;
	wire [4-1:0] node18948;
	wire [4-1:0] node18949;
	wire [4-1:0] node18950;
	wire [4-1:0] node18954;
	wire [4-1:0] node18955;
	wire [4-1:0] node18959;
	wire [4-1:0] node18960;
	wire [4-1:0] node18961;
	wire [4-1:0] node18962;
	wire [4-1:0] node18963;
	wire [4-1:0] node18966;
	wire [4-1:0] node18970;
	wire [4-1:0] node18971;
	wire [4-1:0] node18972;
	wire [4-1:0] node18976;
	wire [4-1:0] node18978;
	wire [4-1:0] node18981;
	wire [4-1:0] node18982;
	wire [4-1:0] node18983;
	wire [4-1:0] node18986;
	wire [4-1:0] node18987;
	wire [4-1:0] node18991;
	wire [4-1:0] node18994;
	wire [4-1:0] node18995;
	wire [4-1:0] node18996;
	wire [4-1:0] node18997;
	wire [4-1:0] node18998;
	wire [4-1:0] node18999;
	wire [4-1:0] node19003;
	wire [4-1:0] node19005;
	wire [4-1:0] node19008;
	wire [4-1:0] node19010;
	wire [4-1:0] node19012;
	wire [4-1:0] node19015;
	wire [4-1:0] node19016;
	wire [4-1:0] node19017;
	wire [4-1:0] node19020;
	wire [4-1:0] node19023;
	wire [4-1:0] node19024;
	wire [4-1:0] node19025;
	wire [4-1:0] node19028;
	wire [4-1:0] node19031;
	wire [4-1:0] node19032;
	wire [4-1:0] node19035;
	wire [4-1:0] node19038;
	wire [4-1:0] node19039;
	wire [4-1:0] node19040;
	wire [4-1:0] node19041;
	wire [4-1:0] node19042;
	wire [4-1:0] node19046;
	wire [4-1:0] node19048;
	wire [4-1:0] node19051;
	wire [4-1:0] node19052;
	wire [4-1:0] node19055;
	wire [4-1:0] node19058;
	wire [4-1:0] node19059;
	wire [4-1:0] node19062;
	wire [4-1:0] node19063;
	wire [4-1:0] node19064;
	wire [4-1:0] node19069;
	wire [4-1:0] node19070;
	wire [4-1:0] node19071;
	wire [4-1:0] node19072;
	wire [4-1:0] node19073;
	wire [4-1:0] node19074;
	wire [4-1:0] node19078;
	wire [4-1:0] node19079;
	wire [4-1:0] node19083;
	wire [4-1:0] node19084;
	wire [4-1:0] node19085;
	wire [4-1:0] node19089;
	wire [4-1:0] node19090;
	wire [4-1:0] node19094;
	wire [4-1:0] node19095;
	wire [4-1:0] node19096;
	wire [4-1:0] node19097;
	wire [4-1:0] node19101;
	wire [4-1:0] node19103;
	wire [4-1:0] node19106;
	wire [4-1:0] node19107;
	wire [4-1:0] node19108;
	wire [4-1:0] node19109;
	wire [4-1:0] node19113;
	wire [4-1:0] node19114;
	wire [4-1:0] node19117;
	wire [4-1:0] node19120;
	wire [4-1:0] node19122;
	wire [4-1:0] node19123;
	wire [4-1:0] node19126;
	wire [4-1:0] node19129;
	wire [4-1:0] node19130;
	wire [4-1:0] node19131;
	wire [4-1:0] node19132;
	wire [4-1:0] node19133;
	wire [4-1:0] node19134;
	wire [4-1:0] node19138;
	wire [4-1:0] node19139;
	wire [4-1:0] node19143;
	wire [4-1:0] node19144;
	wire [4-1:0] node19147;
	wire [4-1:0] node19150;
	wire [4-1:0] node19151;
	wire [4-1:0] node19154;
	wire [4-1:0] node19157;
	wire [4-1:0] node19158;
	wire [4-1:0] node19159;
	wire [4-1:0] node19161;
	wire [4-1:0] node19162;
	wire [4-1:0] node19166;
	wire [4-1:0] node19167;
	wire [4-1:0] node19171;
	wire [4-1:0] node19172;
	wire [4-1:0] node19173;
	wire [4-1:0] node19174;
	wire [4-1:0] node19177;
	wire [4-1:0] node19180;
	wire [4-1:0] node19181;
	wire [4-1:0] node19185;
	wire [4-1:0] node19186;
	wire [4-1:0] node19187;
	wire [4-1:0] node19190;
	wire [4-1:0] node19194;
	wire [4-1:0] node19195;
	wire [4-1:0] node19196;
	wire [4-1:0] node19197;
	wire [4-1:0] node19198;
	wire [4-1:0] node19199;
	wire [4-1:0] node19200;
	wire [4-1:0] node19201;
	wire [4-1:0] node19204;
	wire [4-1:0] node19207;
	wire [4-1:0] node19208;
	wire [4-1:0] node19211;
	wire [4-1:0] node19214;
	wire [4-1:0] node19215;
	wire [4-1:0] node19216;
	wire [4-1:0] node19217;
	wire [4-1:0] node19220;
	wire [4-1:0] node19223;
	wire [4-1:0] node19224;
	wire [4-1:0] node19227;
	wire [4-1:0] node19230;
	wire [4-1:0] node19232;
	wire [4-1:0] node19235;
	wire [4-1:0] node19236;
	wire [4-1:0] node19237;
	wire [4-1:0] node19238;
	wire [4-1:0] node19240;
	wire [4-1:0] node19243;
	wire [4-1:0] node19244;
	wire [4-1:0] node19247;
	wire [4-1:0] node19250;
	wire [4-1:0] node19252;
	wire [4-1:0] node19255;
	wire [4-1:0] node19256;
	wire [4-1:0] node19258;
	wire [4-1:0] node19259;
	wire [4-1:0] node19262;
	wire [4-1:0] node19265;
	wire [4-1:0] node19267;
	wire [4-1:0] node19268;
	wire [4-1:0] node19271;
	wire [4-1:0] node19274;
	wire [4-1:0] node19275;
	wire [4-1:0] node19276;
	wire [4-1:0] node19277;
	wire [4-1:0] node19278;
	wire [4-1:0] node19279;
	wire [4-1:0] node19282;
	wire [4-1:0] node19285;
	wire [4-1:0] node19287;
	wire [4-1:0] node19290;
	wire [4-1:0] node19291;
	wire [4-1:0] node19294;
	wire [4-1:0] node19297;
	wire [4-1:0] node19298;
	wire [4-1:0] node19299;
	wire [4-1:0] node19300;
	wire [4-1:0] node19303;
	wire [4-1:0] node19306;
	wire [4-1:0] node19308;
	wire [4-1:0] node19312;
	wire [4-1:0] node19313;
	wire [4-1:0] node19314;
	wire [4-1:0] node19317;
	wire [4-1:0] node19318;
	wire [4-1:0] node19321;
	wire [4-1:0] node19322;
	wire [4-1:0] node19326;
	wire [4-1:0] node19327;
	wire [4-1:0] node19329;
	wire [4-1:0] node19331;
	wire [4-1:0] node19334;
	wire [4-1:0] node19335;
	wire [4-1:0] node19337;
	wire [4-1:0] node19341;
	wire [4-1:0] node19342;
	wire [4-1:0] node19343;
	wire [4-1:0] node19344;
	wire [4-1:0] node19345;
	wire [4-1:0] node19346;
	wire [4-1:0] node19349;
	wire [4-1:0] node19352;
	wire [4-1:0] node19353;
	wire [4-1:0] node19356;
	wire [4-1:0] node19359;
	wire [4-1:0] node19360;
	wire [4-1:0] node19363;
	wire [4-1:0] node19366;
	wire [4-1:0] node19367;
	wire [4-1:0] node19368;
	wire [4-1:0] node19369;
	wire [4-1:0] node19373;
	wire [4-1:0] node19374;
	wire [4-1:0] node19378;
	wire [4-1:0] node19379;
	wire [4-1:0] node19380;
	wire [4-1:0] node19381;
	wire [4-1:0] node19385;
	wire [4-1:0] node19386;
	wire [4-1:0] node19390;
	wire [4-1:0] node19391;
	wire [4-1:0] node19394;
	wire [4-1:0] node19397;
	wire [4-1:0] node19398;
	wire [4-1:0] node19399;
	wire [4-1:0] node19400;
	wire [4-1:0] node19401;
	wire [4-1:0] node19405;
	wire [4-1:0] node19406;
	wire [4-1:0] node19410;
	wire [4-1:0] node19411;
	wire [4-1:0] node19412;
	wire [4-1:0] node19413;
	wire [4-1:0] node19416;
	wire [4-1:0] node19419;
	wire [4-1:0] node19420;
	wire [4-1:0] node19423;
	wire [4-1:0] node19426;
	wire [4-1:0] node19427;
	wire [4-1:0] node19430;
	wire [4-1:0] node19433;
	wire [4-1:0] node19434;
	wire [4-1:0] node19435;
	wire [4-1:0] node19436;
	wire [4-1:0] node19437;
	wire [4-1:0] node19441;
	wire [4-1:0] node19444;
	wire [4-1:0] node19445;
	wire [4-1:0] node19446;
	wire [4-1:0] node19450;
	wire [4-1:0] node19453;
	wire [4-1:0] node19454;
	wire [4-1:0] node19455;
	wire [4-1:0] node19459;
	wire [4-1:0] node19460;
	wire [4-1:0] node19461;
	wire [4-1:0] node19465;
	wire [4-1:0] node19466;
	wire [4-1:0] node19470;
	wire [4-1:0] node19471;
	wire [4-1:0] node19472;
	wire [4-1:0] node19473;
	wire [4-1:0] node19474;
	wire [4-1:0] node19475;
	wire [4-1:0] node19476;
	wire [4-1:0] node19478;
	wire [4-1:0] node19481;
	wire [4-1:0] node19484;
	wire [4-1:0] node19486;
	wire [4-1:0] node19488;
	wire [4-1:0] node19491;
	wire [4-1:0] node19492;
	wire [4-1:0] node19493;
	wire [4-1:0] node19496;
	wire [4-1:0] node19499;
	wire [4-1:0] node19501;
	wire [4-1:0] node19502;
	wire [4-1:0] node19505;
	wire [4-1:0] node19508;
	wire [4-1:0] node19509;
	wire [4-1:0] node19510;
	wire [4-1:0] node19513;
	wire [4-1:0] node19515;
	wire [4-1:0] node19518;
	wire [4-1:0] node19519;
	wire [4-1:0] node19521;
	wire [4-1:0] node19524;
	wire [4-1:0] node19526;
	wire [4-1:0] node19529;
	wire [4-1:0] node19530;
	wire [4-1:0] node19531;
	wire [4-1:0] node19532;
	wire [4-1:0] node19533;
	wire [4-1:0] node19536;
	wire [4-1:0] node19539;
	wire [4-1:0] node19540;
	wire [4-1:0] node19542;
	wire [4-1:0] node19545;
	wire [4-1:0] node19546;
	wire [4-1:0] node19549;
	wire [4-1:0] node19552;
	wire [4-1:0] node19553;
	wire [4-1:0] node19554;
	wire [4-1:0] node19556;
	wire [4-1:0] node19559;
	wire [4-1:0] node19562;
	wire [4-1:0] node19564;
	wire [4-1:0] node19566;
	wire [4-1:0] node19569;
	wire [4-1:0] node19570;
	wire [4-1:0] node19571;
	wire [4-1:0] node19573;
	wire [4-1:0] node19576;
	wire [4-1:0] node19578;
	wire [4-1:0] node19581;
	wire [4-1:0] node19583;
	wire [4-1:0] node19585;
	wire [4-1:0] node19588;
	wire [4-1:0] node19589;
	wire [4-1:0] node19590;
	wire [4-1:0] node19591;
	wire [4-1:0] node19592;
	wire [4-1:0] node19593;
	wire [4-1:0] node19596;
	wire [4-1:0] node19599;
	wire [4-1:0] node19600;
	wire [4-1:0] node19601;
	wire [4-1:0] node19604;
	wire [4-1:0] node19608;
	wire [4-1:0] node19609;
	wire [4-1:0] node19611;
	wire [4-1:0] node19613;
	wire [4-1:0] node19616;
	wire [4-1:0] node19617;
	wire [4-1:0] node19619;
	wire [4-1:0] node19622;
	wire [4-1:0] node19624;
	wire [4-1:0] node19627;
	wire [4-1:0] node19628;
	wire [4-1:0] node19629;
	wire [4-1:0] node19630;
	wire [4-1:0] node19633;
	wire [4-1:0] node19636;
	wire [4-1:0] node19637;
	wire [4-1:0] node19639;
	wire [4-1:0] node19642;
	wire [4-1:0] node19644;
	wire [4-1:0] node19647;
	wire [4-1:0] node19648;
	wire [4-1:0] node19649;
	wire [4-1:0] node19652;
	wire [4-1:0] node19655;
	wire [4-1:0] node19656;
	wire [4-1:0] node19659;
	wire [4-1:0] node19662;
	wire [4-1:0] node19663;
	wire [4-1:0] node19664;
	wire [4-1:0] node19665;
	wire [4-1:0] node19667;
	wire [4-1:0] node19668;
	wire [4-1:0] node19671;
	wire [4-1:0] node19674;
	wire [4-1:0] node19675;
	wire [4-1:0] node19678;
	wire [4-1:0] node19680;
	wire [4-1:0] node19683;
	wire [4-1:0] node19684;
	wire [4-1:0] node19685;
	wire [4-1:0] node19686;
	wire [4-1:0] node19689;
	wire [4-1:0] node19693;
	wire [4-1:0] node19694;
	wire [4-1:0] node19695;
	wire [4-1:0] node19698;
	wire [4-1:0] node19701;
	wire [4-1:0] node19702;
	wire [4-1:0] node19705;
	wire [4-1:0] node19708;
	wire [4-1:0] node19709;
	wire [4-1:0] node19710;
	wire [4-1:0] node19711;
	wire [4-1:0] node19712;
	wire [4-1:0] node19715;
	wire [4-1:0] node19718;
	wire [4-1:0] node19719;
	wire [4-1:0] node19723;
	wire [4-1:0] node19724;
	wire [4-1:0] node19726;
	wire [4-1:0] node19729;
	wire [4-1:0] node19730;
	wire [4-1:0] node19733;
	wire [4-1:0] node19736;
	wire [4-1:0] node19737;
	wire [4-1:0] node19738;
	wire [4-1:0] node19741;
	wire [4-1:0] node19744;
	wire [4-1:0] node19745;
	wire [4-1:0] node19748;
	wire [4-1:0] node19751;
	wire [4-1:0] node19752;
	wire [4-1:0] node19753;
	wire [4-1:0] node19754;
	wire [4-1:0] node19755;
	wire [4-1:0] node19756;
	wire [4-1:0] node19757;
	wire [4-1:0] node19758;
	wire [4-1:0] node19759;
	wire [4-1:0] node19760;
	wire [4-1:0] node19763;
	wire [4-1:0] node19767;
	wire [4-1:0] node19768;
	wire [4-1:0] node19769;
	wire [4-1:0] node19772;
	wire [4-1:0] node19775;
	wire [4-1:0] node19776;
	wire [4-1:0] node19779;
	wire [4-1:0] node19782;
	wire [4-1:0] node19783;
	wire [4-1:0] node19784;
	wire [4-1:0] node19787;
	wire [4-1:0] node19790;
	wire [4-1:0] node19791;
	wire [4-1:0] node19794;
	wire [4-1:0] node19797;
	wire [4-1:0] node19798;
	wire [4-1:0] node19799;
	wire [4-1:0] node19800;
	wire [4-1:0] node19804;
	wire [4-1:0] node19805;
	wire [4-1:0] node19808;
	wire [4-1:0] node19811;
	wire [4-1:0] node19812;
	wire [4-1:0] node19815;
	wire [4-1:0] node19818;
	wire [4-1:0] node19819;
	wire [4-1:0] node19820;
	wire [4-1:0] node19821;
	wire [4-1:0] node19822;
	wire [4-1:0] node19825;
	wire [4-1:0] node19828;
	wire [4-1:0] node19829;
	wire [4-1:0] node19832;
	wire [4-1:0] node19835;
	wire [4-1:0] node19836;
	wire [4-1:0] node19837;
	wire [4-1:0] node19840;
	wire [4-1:0] node19843;
	wire [4-1:0] node19844;
	wire [4-1:0] node19845;
	wire [4-1:0] node19848;
	wire [4-1:0] node19851;
	wire [4-1:0] node19853;
	wire [4-1:0] node19856;
	wire [4-1:0] node19857;
	wire [4-1:0] node19858;
	wire [4-1:0] node19860;
	wire [4-1:0] node19861;
	wire [4-1:0] node19864;
	wire [4-1:0] node19867;
	wire [4-1:0] node19868;
	wire [4-1:0] node19869;
	wire [4-1:0] node19873;
	wire [4-1:0] node19875;
	wire [4-1:0] node19878;
	wire [4-1:0] node19879;
	wire [4-1:0] node19880;
	wire [4-1:0] node19883;
	wire [4-1:0] node19886;
	wire [4-1:0] node19888;
	wire [4-1:0] node19891;
	wire [4-1:0] node19892;
	wire [4-1:0] node19893;
	wire [4-1:0] node19894;
	wire [4-1:0] node19895;
	wire [4-1:0] node19896;
	wire [4-1:0] node19897;
	wire [4-1:0] node19900;
	wire [4-1:0] node19904;
	wire [4-1:0] node19906;
	wire [4-1:0] node19907;
	wire [4-1:0] node19910;
	wire [4-1:0] node19913;
	wire [4-1:0] node19914;
	wire [4-1:0] node19916;
	wire [4-1:0] node19918;
	wire [4-1:0] node19921;
	wire [4-1:0] node19922;
	wire [4-1:0] node19923;
	wire [4-1:0] node19927;
	wire [4-1:0] node19930;
	wire [4-1:0] node19931;
	wire [4-1:0] node19932;
	wire [4-1:0] node19933;
	wire [4-1:0] node19934;
	wire [4-1:0] node19937;
	wire [4-1:0] node19940;
	wire [4-1:0] node19941;
	wire [4-1:0] node19945;
	wire [4-1:0] node19946;
	wire [4-1:0] node19947;
	wire [4-1:0] node19950;
	wire [4-1:0] node19954;
	wire [4-1:0] node19955;
	wire [4-1:0] node19956;
	wire [4-1:0] node19957;
	wire [4-1:0] node19960;
	wire [4-1:0] node19963;
	wire [4-1:0] node19964;
	wire [4-1:0] node19967;
	wire [4-1:0] node19970;
	wire [4-1:0] node19971;
	wire [4-1:0] node19973;
	wire [4-1:0] node19977;
	wire [4-1:0] node19978;
	wire [4-1:0] node19979;
	wire [4-1:0] node19980;
	wire [4-1:0] node19981;
	wire [4-1:0] node19982;
	wire [4-1:0] node19987;
	wire [4-1:0] node19988;
	wire [4-1:0] node19991;
	wire [4-1:0] node19994;
	wire [4-1:0] node19995;
	wire [4-1:0] node19996;
	wire [4-1:0] node19997;
	wire [4-1:0] node20000;
	wire [4-1:0] node20004;
	wire [4-1:0] node20005;
	wire [4-1:0] node20008;
	wire [4-1:0] node20011;
	wire [4-1:0] node20012;
	wire [4-1:0] node20013;
	wire [4-1:0] node20014;
	wire [4-1:0] node20017;
	wire [4-1:0] node20020;
	wire [4-1:0] node20021;
	wire [4-1:0] node20022;
	wire [4-1:0] node20025;
	wire [4-1:0] node20028;
	wire [4-1:0] node20030;
	wire [4-1:0] node20033;
	wire [4-1:0] node20034;
	wire [4-1:0] node20035;
	wire [4-1:0] node20038;
	wire [4-1:0] node20041;
	wire [4-1:0] node20043;
	wire [4-1:0] node20046;
	wire [4-1:0] node20047;
	wire [4-1:0] node20048;
	wire [4-1:0] node20049;
	wire [4-1:0] node20050;
	wire [4-1:0] node20051;
	wire [4-1:0] node20053;
	wire [4-1:0] node20056;
	wire [4-1:0] node20057;
	wire [4-1:0] node20058;
	wire [4-1:0] node20061;
	wire [4-1:0] node20064;
	wire [4-1:0] node20065;
	wire [4-1:0] node20068;
	wire [4-1:0] node20071;
	wire [4-1:0] node20072;
	wire [4-1:0] node20073;
	wire [4-1:0] node20077;
	wire [4-1:0] node20078;
	wire [4-1:0] node20081;
	wire [4-1:0] node20084;
	wire [4-1:0] node20085;
	wire [4-1:0] node20086;
	wire [4-1:0] node20087;
	wire [4-1:0] node20088;
	wire [4-1:0] node20093;
	wire [4-1:0] node20094;
	wire [4-1:0] node20098;
	wire [4-1:0] node20099;
	wire [4-1:0] node20101;
	wire [4-1:0] node20102;
	wire [4-1:0] node20105;
	wire [4-1:0] node20108;
	wire [4-1:0] node20109;
	wire [4-1:0] node20110;
	wire [4-1:0] node20113;
	wire [4-1:0] node20117;
	wire [4-1:0] node20118;
	wire [4-1:0] node20119;
	wire [4-1:0] node20120;
	wire [4-1:0] node20121;
	wire [4-1:0] node20125;
	wire [4-1:0] node20126;
	wire [4-1:0] node20130;
	wire [4-1:0] node20131;
	wire [4-1:0] node20132;
	wire [4-1:0] node20136;
	wire [4-1:0] node20137;
	wire [4-1:0] node20141;
	wire [4-1:0] node20142;
	wire [4-1:0] node20143;
	wire [4-1:0] node20144;
	wire [4-1:0] node20145;
	wire [4-1:0] node20149;
	wire [4-1:0] node20150;
	wire [4-1:0] node20153;
	wire [4-1:0] node20156;
	wire [4-1:0] node20157;
	wire [4-1:0] node20160;
	wire [4-1:0] node20163;
	wire [4-1:0] node20164;
	wire [4-1:0] node20165;
	wire [4-1:0] node20166;
	wire [4-1:0] node20169;
	wire [4-1:0] node20173;
	wire [4-1:0] node20174;
	wire [4-1:0] node20177;
	wire [4-1:0] node20180;
	wire [4-1:0] node20181;
	wire [4-1:0] node20182;
	wire [4-1:0] node20183;
	wire [4-1:0] node20184;
	wire [4-1:0] node20185;
	wire [4-1:0] node20188;
	wire [4-1:0] node20191;
	wire [4-1:0] node20192;
	wire [4-1:0] node20195;
	wire [4-1:0] node20198;
	wire [4-1:0] node20199;
	wire [4-1:0] node20201;
	wire [4-1:0] node20204;
	wire [4-1:0] node20205;
	wire [4-1:0] node20208;
	wire [4-1:0] node20211;
	wire [4-1:0] node20212;
	wire [4-1:0] node20213;
	wire [4-1:0] node20214;
	wire [4-1:0] node20215;
	wire [4-1:0] node20218;
	wire [4-1:0] node20222;
	wire [4-1:0] node20223;
	wire [4-1:0] node20226;
	wire [4-1:0] node20229;
	wire [4-1:0] node20230;
	wire [4-1:0] node20231;
	wire [4-1:0] node20232;
	wire [4-1:0] node20236;
	wire [4-1:0] node20237;
	wire [4-1:0] node20241;
	wire [4-1:0] node20243;
	wire [4-1:0] node20246;
	wire [4-1:0] node20247;
	wire [4-1:0] node20248;
	wire [4-1:0] node20249;
	wire [4-1:0] node20251;
	wire [4-1:0] node20254;
	wire [4-1:0] node20256;
	wire [4-1:0] node20257;
	wire [4-1:0] node20261;
	wire [4-1:0] node20262;
	wire [4-1:0] node20263;
	wire [4-1:0] node20264;
	wire [4-1:0] node20268;
	wire [4-1:0] node20269;
	wire [4-1:0] node20273;
	wire [4-1:0] node20274;
	wire [4-1:0] node20275;
	wire [4-1:0] node20279;
	wire [4-1:0] node20282;
	wire [4-1:0] node20283;
	wire [4-1:0] node20284;
	wire [4-1:0] node20286;
	wire [4-1:0] node20287;
	wire [4-1:0] node20291;
	wire [4-1:0] node20293;
	wire [4-1:0] node20294;
	wire [4-1:0] node20298;
	wire [4-1:0] node20299;
	wire [4-1:0] node20300;
	wire [4-1:0] node20301;
	wire [4-1:0] node20304;
	wire [4-1:0] node20307;
	wire [4-1:0] node20308;
	wire [4-1:0] node20311;
	wire [4-1:0] node20314;
	wire [4-1:0] node20315;
	wire [4-1:0] node20318;
	wire [4-1:0] node20321;
	wire [4-1:0] node20322;
	wire [4-1:0] node20323;
	wire [4-1:0] node20324;
	wire [4-1:0] node20325;
	wire [4-1:0] node20326;
	wire [4-1:0] node20327;
	wire [4-1:0] node20328;
	wire [4-1:0] node20332;
	wire [4-1:0] node20333;
	wire [4-1:0] node20337;
	wire [4-1:0] node20338;
	wire [4-1:0] node20339;
	wire [4-1:0] node20343;
	wire [4-1:0] node20344;
	wire [4-1:0] node20348;
	wire [4-1:0] node20349;
	wire [4-1:0] node20350;
	wire [4-1:0] node20351;
	wire [4-1:0] node20352;
	wire [4-1:0] node20355;
	wire [4-1:0] node20359;
	wire [4-1:0] node20360;
	wire [4-1:0] node20362;
	wire [4-1:0] node20365;
	wire [4-1:0] node20367;
	wire [4-1:0] node20370;
	wire [4-1:0] node20371;
	wire [4-1:0] node20372;
	wire [4-1:0] node20375;
	wire [4-1:0] node20376;
	wire [4-1:0] node20380;
	wire [4-1:0] node20382;
	wire [4-1:0] node20385;
	wire [4-1:0] node20386;
	wire [4-1:0] node20387;
	wire [4-1:0] node20389;
	wire [4-1:0] node20390;
	wire [4-1:0] node20394;
	wire [4-1:0] node20395;
	wire [4-1:0] node20396;
	wire [4-1:0] node20400;
	wire [4-1:0] node20401;
	wire [4-1:0] node20405;
	wire [4-1:0] node20406;
	wire [4-1:0] node20407;
	wire [4-1:0] node20408;
	wire [4-1:0] node20410;
	wire [4-1:0] node20413;
	wire [4-1:0] node20414;
	wire [4-1:0] node20418;
	wire [4-1:0] node20419;
	wire [4-1:0] node20422;
	wire [4-1:0] node20425;
	wire [4-1:0] node20426;
	wire [4-1:0] node20427;
	wire [4-1:0] node20428;
	wire [4-1:0] node20433;
	wire [4-1:0] node20435;
	wire [4-1:0] node20436;
	wire [4-1:0] node20440;
	wire [4-1:0] node20441;
	wire [4-1:0] node20442;
	wire [4-1:0] node20443;
	wire [4-1:0] node20444;
	wire [4-1:0] node20445;
	wire [4-1:0] node20449;
	wire [4-1:0] node20450;
	wire [4-1:0] node20454;
	wire [4-1:0] node20455;
	wire [4-1:0] node20456;
	wire [4-1:0] node20460;
	wire [4-1:0] node20461;
	wire [4-1:0] node20465;
	wire [4-1:0] node20466;
	wire [4-1:0] node20467;
	wire [4-1:0] node20469;
	wire [4-1:0] node20470;
	wire [4-1:0] node20474;
	wire [4-1:0] node20475;
	wire [4-1:0] node20476;
	wire [4-1:0] node20479;
	wire [4-1:0] node20483;
	wire [4-1:0] node20484;
	wire [4-1:0] node20485;
	wire [4-1:0] node20486;
	wire [4-1:0] node20491;
	wire [4-1:0] node20494;
	wire [4-1:0] node20495;
	wire [4-1:0] node20496;
	wire [4-1:0] node20497;
	wire [4-1:0] node20498;
	wire [4-1:0] node20501;
	wire [4-1:0] node20504;
	wire [4-1:0] node20505;
	wire [4-1:0] node20506;
	wire [4-1:0] node20509;
	wire [4-1:0] node20512;
	wire [4-1:0] node20513;
	wire [4-1:0] node20516;
	wire [4-1:0] node20519;
	wire [4-1:0] node20520;
	wire [4-1:0] node20523;
	wire [4-1:0] node20526;
	wire [4-1:0] node20527;
	wire [4-1:0] node20528;
	wire [4-1:0] node20529;
	wire [4-1:0] node20530;
	wire [4-1:0] node20533;
	wire [4-1:0] node20537;
	wire [4-1:0] node20538;
	wire [4-1:0] node20541;
	wire [4-1:0] node20544;
	wire [4-1:0] node20545;
	wire [4-1:0] node20546;
	wire [4-1:0] node20547;
	wire [4-1:0] node20550;
	wire [4-1:0] node20554;
	wire [4-1:0] node20556;
	wire [4-1:0] node20559;
	wire [4-1:0] node20560;
	wire [4-1:0] node20561;
	wire [4-1:0] node20562;
	wire [4-1:0] node20563;
	wire [4-1:0] node20564;
	wire [4-1:0] node20565;
	wire [4-1:0] node20568;
	wire [4-1:0] node20571;
	wire [4-1:0] node20572;
	wire [4-1:0] node20576;
	wire [4-1:0] node20577;
	wire [4-1:0] node20578;
	wire [4-1:0] node20579;
	wire [4-1:0] node20582;
	wire [4-1:0] node20585;
	wire [4-1:0] node20586;
	wire [4-1:0] node20590;
	wire [4-1:0] node20591;
	wire [4-1:0] node20594;
	wire [4-1:0] node20597;
	wire [4-1:0] node20598;
	wire [4-1:0] node20599;
	wire [4-1:0] node20601;
	wire [4-1:0] node20602;
	wire [4-1:0] node20605;
	wire [4-1:0] node20608;
	wire [4-1:0] node20609;
	wire [4-1:0] node20612;
	wire [4-1:0] node20615;
	wire [4-1:0] node20616;
	wire [4-1:0] node20617;
	wire [4-1:0] node20618;
	wire [4-1:0] node20622;
	wire [4-1:0] node20623;
	wire [4-1:0] node20627;
	wire [4-1:0] node20628;
	wire [4-1:0] node20632;
	wire [4-1:0] node20633;
	wire [4-1:0] node20634;
	wire [4-1:0] node20635;
	wire [4-1:0] node20636;
	wire [4-1:0] node20637;
	wire [4-1:0] node20640;
	wire [4-1:0] node20643;
	wire [4-1:0] node20644;
	wire [4-1:0] node20647;
	wire [4-1:0] node20650;
	wire [4-1:0] node20651;
	wire [4-1:0] node20652;
	wire [4-1:0] node20655;
	wire [4-1:0] node20658;
	wire [4-1:0] node20659;
	wire [4-1:0] node20662;
	wire [4-1:0] node20665;
	wire [4-1:0] node20666;
	wire [4-1:0] node20667;
	wire [4-1:0] node20668;
	wire [4-1:0] node20672;
	wire [4-1:0] node20675;
	wire [4-1:0] node20676;
	wire [4-1:0] node20678;
	wire [4-1:0] node20682;
	wire [4-1:0] node20683;
	wire [4-1:0] node20684;
	wire [4-1:0] node20685;
	wire [4-1:0] node20689;
	wire [4-1:0] node20691;
	wire [4-1:0] node20694;
	wire [4-1:0] node20695;
	wire [4-1:0] node20696;
	wire [4-1:0] node20697;
	wire [4-1:0] node20700;
	wire [4-1:0] node20703;
	wire [4-1:0] node20704;
	wire [4-1:0] node20707;
	wire [4-1:0] node20710;
	wire [4-1:0] node20711;
	wire [4-1:0] node20712;
	wire [4-1:0] node20716;
	wire [4-1:0] node20717;
	wire [4-1:0] node20720;
	wire [4-1:0] node20723;
	wire [4-1:0] node20724;
	wire [4-1:0] node20725;
	wire [4-1:0] node20726;
	wire [4-1:0] node20727;
	wire [4-1:0] node20728;
	wire [4-1:0] node20729;
	wire [4-1:0] node20733;
	wire [4-1:0] node20734;
	wire [4-1:0] node20738;
	wire [4-1:0] node20739;
	wire [4-1:0] node20742;
	wire [4-1:0] node20745;
	wire [4-1:0] node20746;
	wire [4-1:0] node20747;
	wire [4-1:0] node20750;
	wire [4-1:0] node20753;
	wire [4-1:0] node20754;
	wire [4-1:0] node20758;
	wire [4-1:0] node20759;
	wire [4-1:0] node20760;
	wire [4-1:0] node20761;
	wire [4-1:0] node20762;
	wire [4-1:0] node20765;
	wire [4-1:0] node20769;
	wire [4-1:0] node20770;
	wire [4-1:0] node20773;
	wire [4-1:0] node20774;
	wire [4-1:0] node20778;
	wire [4-1:0] node20779;
	wire [4-1:0] node20780;
	wire [4-1:0] node20784;
	wire [4-1:0] node20786;
	wire [4-1:0] node20789;
	wire [4-1:0] node20790;
	wire [4-1:0] node20791;
	wire [4-1:0] node20792;
	wire [4-1:0] node20793;
	wire [4-1:0] node20796;
	wire [4-1:0] node20799;
	wire [4-1:0] node20800;
	wire [4-1:0] node20803;
	wire [4-1:0] node20806;
	wire [4-1:0] node20807;
	wire [4-1:0] node20808;
	wire [4-1:0] node20811;
	wire [4-1:0] node20814;
	wire [4-1:0] node20815;
	wire [4-1:0] node20819;
	wire [4-1:0] node20820;
	wire [4-1:0] node20821;
	wire [4-1:0] node20822;
	wire [4-1:0] node20823;
	wire [4-1:0] node20827;
	wire [4-1:0] node20828;
	wire [4-1:0] node20832;
	wire [4-1:0] node20833;
	wire [4-1:0] node20834;
	wire [4-1:0] node20839;
	wire [4-1:0] node20840;
	wire [4-1:0] node20842;
	wire [4-1:0] node20843;
	wire [4-1:0] node20847;
	wire [4-1:0] node20848;
	wire [4-1:0] node20851;
	wire [4-1:0] node20854;
	wire [4-1:0] node20855;
	wire [4-1:0] node20856;
	wire [4-1:0] node20857;
	wire [4-1:0] node20858;
	wire [4-1:0] node20859;
	wire [4-1:0] node20860;
	wire [4-1:0] node20861;
	wire [4-1:0] node20862;
	wire [4-1:0] node20863;
	wire [4-1:0] node20865;
	wire [4-1:0] node20866;
	wire [4-1:0] node20869;
	wire [4-1:0] node20872;
	wire [4-1:0] node20874;
	wire [4-1:0] node20875;
	wire [4-1:0] node20879;
	wire [4-1:0] node20880;
	wire [4-1:0] node20881;
	wire [4-1:0] node20884;
	wire [4-1:0] node20887;
	wire [4-1:0] node20888;
	wire [4-1:0] node20892;
	wire [4-1:0] node20893;
	wire [4-1:0] node20895;
	wire [4-1:0] node20897;
	wire [4-1:0] node20898;
	wire [4-1:0] node20901;
	wire [4-1:0] node20904;
	wire [4-1:0] node20905;
	wire [4-1:0] node20907;
	wire [4-1:0] node20908;
	wire [4-1:0] node20911;
	wire [4-1:0] node20914;
	wire [4-1:0] node20917;
	wire [4-1:0] node20918;
	wire [4-1:0] node20919;
	wire [4-1:0] node20920;
	wire [4-1:0] node20921;
	wire [4-1:0] node20923;
	wire [4-1:0] node20926;
	wire [4-1:0] node20928;
	wire [4-1:0] node20931;
	wire [4-1:0] node20932;
	wire [4-1:0] node20934;
	wire [4-1:0] node20938;
	wire [4-1:0] node20939;
	wire [4-1:0] node20940;
	wire [4-1:0] node20943;
	wire [4-1:0] node20946;
	wire [4-1:0] node20947;
	wire [4-1:0] node20949;
	wire [4-1:0] node20953;
	wire [4-1:0] node20954;
	wire [4-1:0] node20955;
	wire [4-1:0] node20956;
	wire [4-1:0] node20960;
	wire [4-1:0] node20961;
	wire [4-1:0] node20963;
	wire [4-1:0] node20966;
	wire [4-1:0] node20968;
	wire [4-1:0] node20971;
	wire [4-1:0] node20972;
	wire [4-1:0] node20973;
	wire [4-1:0] node20974;
	wire [4-1:0] node20977;
	wire [4-1:0] node20980;
	wire [4-1:0] node20982;
	wire [4-1:0] node20985;
	wire [4-1:0] node20986;
	wire [4-1:0] node20987;
	wire [4-1:0] node20990;
	wire [4-1:0] node20994;
	wire [4-1:0] node20995;
	wire [4-1:0] node20996;
	wire [4-1:0] node20997;
	wire [4-1:0] node20998;
	wire [4-1:0] node20999;
	wire [4-1:0] node21003;
	wire [4-1:0] node21004;
	wire [4-1:0] node21007;
	wire [4-1:0] node21010;
	wire [4-1:0] node21011;
	wire [4-1:0] node21012;
	wire [4-1:0] node21015;
	wire [4-1:0] node21018;
	wire [4-1:0] node21019;
	wire [4-1:0] node21020;
	wire [4-1:0] node21024;
	wire [4-1:0] node21025;
	wire [4-1:0] node21029;
	wire [4-1:0] node21030;
	wire [4-1:0] node21031;
	wire [4-1:0] node21033;
	wire [4-1:0] node21036;
	wire [4-1:0] node21037;
	wire [4-1:0] node21039;
	wire [4-1:0] node21042;
	wire [4-1:0] node21045;
	wire [4-1:0] node21046;
	wire [4-1:0] node21047;
	wire [4-1:0] node21049;
	wire [4-1:0] node21052;
	wire [4-1:0] node21053;
	wire [4-1:0] node21056;
	wire [4-1:0] node21059;
	wire [4-1:0] node21060;
	wire [4-1:0] node21063;
	wire [4-1:0] node21066;
	wire [4-1:0] node21067;
	wire [4-1:0] node21068;
	wire [4-1:0] node21069;
	wire [4-1:0] node21071;
	wire [4-1:0] node21072;
	wire [4-1:0] node21075;
	wire [4-1:0] node21078;
	wire [4-1:0] node21079;
	wire [4-1:0] node21080;
	wire [4-1:0] node21083;
	wire [4-1:0] node21086;
	wire [4-1:0] node21087;
	wire [4-1:0] node21091;
	wire [4-1:0] node21092;
	wire [4-1:0] node21093;
	wire [4-1:0] node21096;
	wire [4-1:0] node21099;
	wire [4-1:0] node21100;
	wire [4-1:0] node21103;
	wire [4-1:0] node21104;
	wire [4-1:0] node21108;
	wire [4-1:0] node21109;
	wire [4-1:0] node21110;
	wire [4-1:0] node21111;
	wire [4-1:0] node21112;
	wire [4-1:0] node21116;
	wire [4-1:0] node21117;
	wire [4-1:0] node21121;
	wire [4-1:0] node21123;
	wire [4-1:0] node21124;
	wire [4-1:0] node21128;
	wire [4-1:0] node21129;
	wire [4-1:0] node21130;
	wire [4-1:0] node21132;
	wire [4-1:0] node21135;
	wire [4-1:0] node21137;
	wire [4-1:0] node21140;
	wire [4-1:0] node21141;
	wire [4-1:0] node21144;
	wire [4-1:0] node21147;
	wire [4-1:0] node21148;
	wire [4-1:0] node21149;
	wire [4-1:0] node21150;
	wire [4-1:0] node21151;
	wire [4-1:0] node21153;
	wire [4-1:0] node21154;
	wire [4-1:0] node21157;
	wire [4-1:0] node21159;
	wire [4-1:0] node21162;
	wire [4-1:0] node21163;
	wire [4-1:0] node21164;
	wire [4-1:0] node21166;
	wire [4-1:0] node21170;
	wire [4-1:0] node21171;
	wire [4-1:0] node21174;
	wire [4-1:0] node21176;
	wire [4-1:0] node21179;
	wire [4-1:0] node21180;
	wire [4-1:0] node21181;
	wire [4-1:0] node21182;
	wire [4-1:0] node21185;
	wire [4-1:0] node21188;
	wire [4-1:0] node21189;
	wire [4-1:0] node21191;
	wire [4-1:0] node21194;
	wire [4-1:0] node21196;
	wire [4-1:0] node21199;
	wire [4-1:0] node21200;
	wire [4-1:0] node21201;
	wire [4-1:0] node21203;
	wire [4-1:0] node21206;
	wire [4-1:0] node21208;
	wire [4-1:0] node21211;
	wire [4-1:0] node21212;
	wire [4-1:0] node21215;
	wire [4-1:0] node21217;
	wire [4-1:0] node21220;
	wire [4-1:0] node21221;
	wire [4-1:0] node21222;
	wire [4-1:0] node21223;
	wire [4-1:0] node21224;
	wire [4-1:0] node21227;
	wire [4-1:0] node21230;
	wire [4-1:0] node21231;
	wire [4-1:0] node21235;
	wire [4-1:0] node21237;
	wire [4-1:0] node21238;
	wire [4-1:0] node21239;
	wire [4-1:0] node21243;
	wire [4-1:0] node21245;
	wire [4-1:0] node21248;
	wire [4-1:0] node21249;
	wire [4-1:0] node21250;
	wire [4-1:0] node21252;
	wire [4-1:0] node21255;
	wire [4-1:0] node21257;
	wire [4-1:0] node21260;
	wire [4-1:0] node21261;
	wire [4-1:0] node21263;
	wire [4-1:0] node21265;
	wire [4-1:0] node21268;
	wire [4-1:0] node21271;
	wire [4-1:0] node21272;
	wire [4-1:0] node21273;
	wire [4-1:0] node21274;
	wire [4-1:0] node21275;
	wire [4-1:0] node21276;
	wire [4-1:0] node21278;
	wire [4-1:0] node21282;
	wire [4-1:0] node21283;
	wire [4-1:0] node21285;
	wire [4-1:0] node21288;
	wire [4-1:0] node21290;
	wire [4-1:0] node21293;
	wire [4-1:0] node21294;
	wire [4-1:0] node21295;
	wire [4-1:0] node21297;
	wire [4-1:0] node21301;
	wire [4-1:0] node21302;
	wire [4-1:0] node21306;
	wire [4-1:0] node21307;
	wire [4-1:0] node21308;
	wire [4-1:0] node21309;
	wire [4-1:0] node21311;
	wire [4-1:0] node21314;
	wire [4-1:0] node21316;
	wire [4-1:0] node21319;
	wire [4-1:0] node21320;
	wire [4-1:0] node21323;
	wire [4-1:0] node21325;
	wire [4-1:0] node21328;
	wire [4-1:0] node21329;
	wire [4-1:0] node21331;
	wire [4-1:0] node21333;
	wire [4-1:0] node21337;
	wire [4-1:0] node21338;
	wire [4-1:0] node21339;
	wire [4-1:0] node21340;
	wire [4-1:0] node21341;
	wire [4-1:0] node21343;
	wire [4-1:0] node21346;
	wire [4-1:0] node21348;
	wire [4-1:0] node21351;
	wire [4-1:0] node21352;
	wire [4-1:0] node21356;
	wire [4-1:0] node21357;
	wire [4-1:0] node21358;
	wire [4-1:0] node21362;
	wire [4-1:0] node21363;
	wire [4-1:0] node21367;
	wire [4-1:0] node21368;
	wire [4-1:0] node21369;
	wire [4-1:0] node21370;
	wire [4-1:0] node21373;
	wire [4-1:0] node21375;
	wire [4-1:0] node21378;
	wire [4-1:0] node21379;
	wire [4-1:0] node21383;
	wire [4-1:0] node21384;
	wire [4-1:0] node21385;
	wire [4-1:0] node21388;
	wire [4-1:0] node21391;
	wire [4-1:0] node21392;
	wire [4-1:0] node21393;
	wire [4-1:0] node21396;
	wire [4-1:0] node21399;
	wire [4-1:0] node21401;
	wire [4-1:0] node21404;
	wire [4-1:0] node21405;
	wire [4-1:0] node21406;
	wire [4-1:0] node21407;
	wire [4-1:0] node21408;
	wire [4-1:0] node21409;
	wire [4-1:0] node21410;
	wire [4-1:0] node21411;
	wire [4-1:0] node21414;
	wire [4-1:0] node21417;
	wire [4-1:0] node21418;
	wire [4-1:0] node21421;
	wire [4-1:0] node21424;
	wire [4-1:0] node21425;
	wire [4-1:0] node21426;
	wire [4-1:0] node21427;
	wire [4-1:0] node21430;
	wire [4-1:0] node21433;
	wire [4-1:0] node21435;
	wire [4-1:0] node21438;
	wire [4-1:0] node21440;
	wire [4-1:0] node21441;
	wire [4-1:0] node21444;
	wire [4-1:0] node21447;
	wire [4-1:0] node21448;
	wire [4-1:0] node21449;
	wire [4-1:0] node21450;
	wire [4-1:0] node21451;
	wire [4-1:0] node21454;
	wire [4-1:0] node21457;
	wire [4-1:0] node21458;
	wire [4-1:0] node21461;
	wire [4-1:0] node21464;
	wire [4-1:0] node21465;
	wire [4-1:0] node21468;
	wire [4-1:0] node21471;
	wire [4-1:0] node21472;
	wire [4-1:0] node21474;
	wire [4-1:0] node21475;
	wire [4-1:0] node21478;
	wire [4-1:0] node21481;
	wire [4-1:0] node21483;
	wire [4-1:0] node21485;
	wire [4-1:0] node21488;
	wire [4-1:0] node21489;
	wire [4-1:0] node21490;
	wire [4-1:0] node21491;
	wire [4-1:0] node21492;
	wire [4-1:0] node21495;
	wire [4-1:0] node21498;
	wire [4-1:0] node21500;
	wire [4-1:0] node21501;
	wire [4-1:0] node21504;
	wire [4-1:0] node21507;
	wire [4-1:0] node21508;
	wire [4-1:0] node21509;
	wire [4-1:0] node21512;
	wire [4-1:0] node21515;
	wire [4-1:0] node21516;
	wire [4-1:0] node21517;
	wire [4-1:0] node21521;
	wire [4-1:0] node21523;
	wire [4-1:0] node21526;
	wire [4-1:0] node21527;
	wire [4-1:0] node21528;
	wire [4-1:0] node21529;
	wire [4-1:0] node21532;
	wire [4-1:0] node21535;
	wire [4-1:0] node21536;
	wire [4-1:0] node21539;
	wire [4-1:0] node21542;
	wire [4-1:0] node21543;
	wire [4-1:0] node21545;
	wire [4-1:0] node21548;
	wire [4-1:0] node21549;
	wire [4-1:0] node21552;
	wire [4-1:0] node21555;
	wire [4-1:0] node21556;
	wire [4-1:0] node21557;
	wire [4-1:0] node21558;
	wire [4-1:0] node21559;
	wire [4-1:0] node21562;
	wire [4-1:0] node21564;
	wire [4-1:0] node21567;
	wire [4-1:0] node21568;
	wire [4-1:0] node21569;
	wire [4-1:0] node21572;
	wire [4-1:0] node21575;
	wire [4-1:0] node21576;
	wire [4-1:0] node21579;
	wire [4-1:0] node21582;
	wire [4-1:0] node21583;
	wire [4-1:0] node21584;
	wire [4-1:0] node21587;
	wire [4-1:0] node21589;
	wire [4-1:0] node21592;
	wire [4-1:0] node21593;
	wire [4-1:0] node21594;
	wire [4-1:0] node21597;
	wire [4-1:0] node21600;
	wire [4-1:0] node21601;
	wire [4-1:0] node21604;
	wire [4-1:0] node21607;
	wire [4-1:0] node21608;
	wire [4-1:0] node21609;
	wire [4-1:0] node21610;
	wire [4-1:0] node21613;
	wire [4-1:0] node21616;
	wire [4-1:0] node21617;
	wire [4-1:0] node21618;
	wire [4-1:0] node21621;
	wire [4-1:0] node21624;
	wire [4-1:0] node21625;
	wire [4-1:0] node21626;
	wire [4-1:0] node21629;
	wire [4-1:0] node21632;
	wire [4-1:0] node21634;
	wire [4-1:0] node21637;
	wire [4-1:0] node21638;
	wire [4-1:0] node21639;
	wire [4-1:0] node21642;
	wire [4-1:0] node21644;
	wire [4-1:0] node21647;
	wire [4-1:0] node21648;
	wire [4-1:0] node21649;
	wire [4-1:0] node21653;
	wire [4-1:0] node21654;
	wire [4-1:0] node21655;
	wire [4-1:0] node21658;
	wire [4-1:0] node21661;
	wire [4-1:0] node21663;
	wire [4-1:0] node21666;
	wire [4-1:0] node21667;
	wire [4-1:0] node21668;
	wire [4-1:0] node21669;
	wire [4-1:0] node21670;
	wire [4-1:0] node21671;
	wire [4-1:0] node21672;
	wire [4-1:0] node21677;
	wire [4-1:0] node21678;
	wire [4-1:0] node21680;
	wire [4-1:0] node21683;
	wire [4-1:0] node21685;
	wire [4-1:0] node21688;
	wire [4-1:0] node21689;
	wire [4-1:0] node21690;
	wire [4-1:0] node21692;
	wire [4-1:0] node21695;
	wire [4-1:0] node21697;
	wire [4-1:0] node21700;
	wire [4-1:0] node21701;
	wire [4-1:0] node21703;
	wire [4-1:0] node21706;
	wire [4-1:0] node21709;
	wire [4-1:0] node21710;
	wire [4-1:0] node21711;
	wire [4-1:0] node21713;
	wire [4-1:0] node21715;
	wire [4-1:0] node21718;
	wire [4-1:0] node21719;
	wire [4-1:0] node21721;
	wire [4-1:0] node21724;
	wire [4-1:0] node21726;
	wire [4-1:0] node21729;
	wire [4-1:0] node21730;
	wire [4-1:0] node21731;
	wire [4-1:0] node21732;
	wire [4-1:0] node21735;
	wire [4-1:0] node21738;
	wire [4-1:0] node21739;
	wire [4-1:0] node21742;
	wire [4-1:0] node21745;
	wire [4-1:0] node21747;
	wire [4-1:0] node21748;
	wire [4-1:0] node21752;
	wire [4-1:0] node21753;
	wire [4-1:0] node21754;
	wire [4-1:0] node21755;
	wire [4-1:0] node21756;
	wire [4-1:0] node21757;
	wire [4-1:0] node21760;
	wire [4-1:0] node21763;
	wire [4-1:0] node21766;
	wire [4-1:0] node21767;
	wire [4-1:0] node21768;
	wire [4-1:0] node21771;
	wire [4-1:0] node21774;
	wire [4-1:0] node21775;
	wire [4-1:0] node21778;
	wire [4-1:0] node21781;
	wire [4-1:0] node21782;
	wire [4-1:0] node21783;
	wire [4-1:0] node21784;
	wire [4-1:0] node21785;
	wire [4-1:0] node21789;
	wire [4-1:0] node21791;
	wire [4-1:0] node21794;
	wire [4-1:0] node21795;
	wire [4-1:0] node21798;
	wire [4-1:0] node21801;
	wire [4-1:0] node21802;
	wire [4-1:0] node21804;
	wire [4-1:0] node21807;
	wire [4-1:0] node21808;
	wire [4-1:0] node21809;
	wire [4-1:0] node21812;
	wire [4-1:0] node21815;
	wire [4-1:0] node21816;
	wire [4-1:0] node21820;
	wire [4-1:0] node21821;
	wire [4-1:0] node21822;
	wire [4-1:0] node21823;
	wire [4-1:0] node21824;
	wire [4-1:0] node21828;
	wire [4-1:0] node21829;
	wire [4-1:0] node21832;
	wire [4-1:0] node21835;
	wire [4-1:0] node21836;
	wire [4-1:0] node21837;
	wire [4-1:0] node21841;
	wire [4-1:0] node21844;
	wire [4-1:0] node21845;
	wire [4-1:0] node21846;
	wire [4-1:0] node21847;
	wire [4-1:0] node21850;
	wire [4-1:0] node21853;
	wire [4-1:0] node21854;
	wire [4-1:0] node21857;
	wire [4-1:0] node21860;
	wire [4-1:0] node21861;
	wire [4-1:0] node21862;
	wire [4-1:0] node21866;
	wire [4-1:0] node21869;
	wire [4-1:0] node21870;
	wire [4-1:0] node21871;
	wire [4-1:0] node21872;
	wire [4-1:0] node21873;
	wire [4-1:0] node21874;
	wire [4-1:0] node21875;
	wire [4-1:0] node21876;
	wire [4-1:0] node21879;
	wire [4-1:0] node21882;
	wire [4-1:0] node21883;
	wire [4-1:0] node21886;
	wire [4-1:0] node21889;
	wire [4-1:0] node21890;
	wire [4-1:0] node21891;
	wire [4-1:0] node21894;
	wire [4-1:0] node21897;
	wire [4-1:0] node21898;
	wire [4-1:0] node21900;
	wire [4-1:0] node21901;
	wire [4-1:0] node21904;
	wire [4-1:0] node21908;
	wire [4-1:0] node21909;
	wire [4-1:0] node21910;
	wire [4-1:0] node21911;
	wire [4-1:0] node21912;
	wire [4-1:0] node21916;
	wire [4-1:0] node21917;
	wire [4-1:0] node21918;
	wire [4-1:0] node21921;
	wire [4-1:0] node21924;
	wire [4-1:0] node21925;
	wire [4-1:0] node21929;
	wire [4-1:0] node21930;
	wire [4-1:0] node21931;
	wire [4-1:0] node21933;
	wire [4-1:0] node21936;
	wire [4-1:0] node21938;
	wire [4-1:0] node21941;
	wire [4-1:0] node21942;
	wire [4-1:0] node21945;
	wire [4-1:0] node21948;
	wire [4-1:0] node21949;
	wire [4-1:0] node21950;
	wire [4-1:0] node21951;
	wire [4-1:0] node21952;
	wire [4-1:0] node21955;
	wire [4-1:0] node21958;
	wire [4-1:0] node21959;
	wire [4-1:0] node21962;
	wire [4-1:0] node21965;
	wire [4-1:0] node21966;
	wire [4-1:0] node21968;
	wire [4-1:0] node21971;
	wire [4-1:0] node21973;
	wire [4-1:0] node21976;
	wire [4-1:0] node21977;
	wire [4-1:0] node21980;
	wire [4-1:0] node21983;
	wire [4-1:0] node21984;
	wire [4-1:0] node21985;
	wire [4-1:0] node21986;
	wire [4-1:0] node21987;
	wire [4-1:0] node21988;
	wire [4-1:0] node21991;
	wire [4-1:0] node21993;
	wire [4-1:0] node21996;
	wire [4-1:0] node21997;
	wire [4-1:0] node22000;
	wire [4-1:0] node22002;
	wire [4-1:0] node22005;
	wire [4-1:0] node22006;
	wire [4-1:0] node22007;
	wire [4-1:0] node22010;
	wire [4-1:0] node22012;
	wire [4-1:0] node22015;
	wire [4-1:0] node22018;
	wire [4-1:0] node22019;
	wire [4-1:0] node22020;
	wire [4-1:0] node22021;
	wire [4-1:0] node22022;
	wire [4-1:0] node22025;
	wire [4-1:0] node22028;
	wire [4-1:0] node22029;
	wire [4-1:0] node22033;
	wire [4-1:0] node22034;
	wire [4-1:0] node22035;
	wire [4-1:0] node22038;
	wire [4-1:0] node22041;
	wire [4-1:0] node22043;
	wire [4-1:0] node22046;
	wire [4-1:0] node22047;
	wire [4-1:0] node22048;
	wire [4-1:0] node22049;
	wire [4-1:0] node22052;
	wire [4-1:0] node22055;
	wire [4-1:0] node22056;
	wire [4-1:0] node22059;
	wire [4-1:0] node22062;
	wire [4-1:0] node22064;
	wire [4-1:0] node22066;
	wire [4-1:0] node22069;
	wire [4-1:0] node22070;
	wire [4-1:0] node22071;
	wire [4-1:0] node22072;
	wire [4-1:0] node22073;
	wire [4-1:0] node22076;
	wire [4-1:0] node22078;
	wire [4-1:0] node22081;
	wire [4-1:0] node22082;
	wire [4-1:0] node22085;
	wire [4-1:0] node22088;
	wire [4-1:0] node22089;
	wire [4-1:0] node22090;
	wire [4-1:0] node22091;
	wire [4-1:0] node22094;
	wire [4-1:0] node22097;
	wire [4-1:0] node22098;
	wire [4-1:0] node22101;
	wire [4-1:0] node22104;
	wire [4-1:0] node22105;
	wire [4-1:0] node22108;
	wire [4-1:0] node22111;
	wire [4-1:0] node22112;
	wire [4-1:0] node22113;
	wire [4-1:0] node22114;
	wire [4-1:0] node22116;
	wire [4-1:0] node22119;
	wire [4-1:0] node22120;
	wire [4-1:0] node22123;
	wire [4-1:0] node22126;
	wire [4-1:0] node22127;
	wire [4-1:0] node22130;
	wire [4-1:0] node22133;
	wire [4-1:0] node22134;
	wire [4-1:0] node22135;
	wire [4-1:0] node22137;
	wire [4-1:0] node22140;
	wire [4-1:0] node22142;
	wire [4-1:0] node22145;
	wire [4-1:0] node22146;
	wire [4-1:0] node22149;
	wire [4-1:0] node22152;
	wire [4-1:0] node22153;
	wire [4-1:0] node22154;
	wire [4-1:0] node22155;
	wire [4-1:0] node22156;
	wire [4-1:0] node22157;
	wire [4-1:0] node22158;
	wire [4-1:0] node22161;
	wire [4-1:0] node22163;
	wire [4-1:0] node22166;
	wire [4-1:0] node22168;
	wire [4-1:0] node22170;
	wire [4-1:0] node22173;
	wire [4-1:0] node22174;
	wire [4-1:0] node22175;
	wire [4-1:0] node22178;
	wire [4-1:0] node22179;
	wire [4-1:0] node22183;
	wire [4-1:0] node22185;
	wire [4-1:0] node22186;
	wire [4-1:0] node22190;
	wire [4-1:0] node22191;
	wire [4-1:0] node22192;
	wire [4-1:0] node22193;
	wire [4-1:0] node22195;
	wire [4-1:0] node22198;
	wire [4-1:0] node22201;
	wire [4-1:0] node22202;
	wire [4-1:0] node22203;
	wire [4-1:0] node22207;
	wire [4-1:0] node22208;
	wire [4-1:0] node22211;
	wire [4-1:0] node22214;
	wire [4-1:0] node22215;
	wire [4-1:0] node22217;
	wire [4-1:0] node22219;
	wire [4-1:0] node22223;
	wire [4-1:0] node22224;
	wire [4-1:0] node22225;
	wire [4-1:0] node22226;
	wire [4-1:0] node22227;
	wire [4-1:0] node22230;
	wire [4-1:0] node22232;
	wire [4-1:0] node22235;
	wire [4-1:0] node22236;
	wire [4-1:0] node22238;
	wire [4-1:0] node22241;
	wire [4-1:0] node22242;
	wire [4-1:0] node22246;
	wire [4-1:0] node22247;
	wire [4-1:0] node22248;
	wire [4-1:0] node22249;
	wire [4-1:0] node22253;
	wire [4-1:0] node22254;
	wire [4-1:0] node22258;
	wire [4-1:0] node22261;
	wire [4-1:0] node22262;
	wire [4-1:0] node22263;
	wire [4-1:0] node22264;
	wire [4-1:0] node22266;
	wire [4-1:0] node22269;
	wire [4-1:0] node22270;
	wire [4-1:0] node22273;
	wire [4-1:0] node22276;
	wire [4-1:0] node22277;
	wire [4-1:0] node22279;
	wire [4-1:0] node22282;
	wire [4-1:0] node22284;
	wire [4-1:0] node22287;
	wire [4-1:0] node22288;
	wire [4-1:0] node22290;
	wire [4-1:0] node22293;
	wire [4-1:0] node22294;
	wire [4-1:0] node22295;
	wire [4-1:0] node22298;
	wire [4-1:0] node22301;
	wire [4-1:0] node22302;
	wire [4-1:0] node22305;
	wire [4-1:0] node22308;
	wire [4-1:0] node22309;
	wire [4-1:0] node22310;
	wire [4-1:0] node22311;
	wire [4-1:0] node22312;
	wire [4-1:0] node22313;
	wire [4-1:0] node22316;
	wire [4-1:0] node22319;
	wire [4-1:0] node22320;
	wire [4-1:0] node22321;
	wire [4-1:0] node22325;
	wire [4-1:0] node22326;
	wire [4-1:0] node22330;
	wire [4-1:0] node22331;
	wire [4-1:0] node22332;
	wire [4-1:0] node22333;
	wire [4-1:0] node22338;
	wire [4-1:0] node22339;
	wire [4-1:0] node22342;
	wire [4-1:0] node22345;
	wire [4-1:0] node22346;
	wire [4-1:0] node22347;
	wire [4-1:0] node22348;
	wire [4-1:0] node22351;
	wire [4-1:0] node22354;
	wire [4-1:0] node22355;
	wire [4-1:0] node22359;
	wire [4-1:0] node22360;
	wire [4-1:0] node22361;
	wire [4-1:0] node22362;
	wire [4-1:0] node22366;
	wire [4-1:0] node22369;
	wire [4-1:0] node22371;
	wire [4-1:0] node22372;
	wire [4-1:0] node22376;
	wire [4-1:0] node22377;
	wire [4-1:0] node22378;
	wire [4-1:0] node22379;
	wire [4-1:0] node22380;
	wire [4-1:0] node22383;
	wire [4-1:0] node22384;
	wire [4-1:0] node22387;
	wire [4-1:0] node22390;
	wire [4-1:0] node22391;
	wire [4-1:0] node22392;
	wire [4-1:0] node22396;
	wire [4-1:0] node22397;
	wire [4-1:0] node22400;
	wire [4-1:0] node22403;
	wire [4-1:0] node22404;
	wire [4-1:0] node22405;
	wire [4-1:0] node22407;
	wire [4-1:0] node22410;
	wire [4-1:0] node22411;
	wire [4-1:0] node22414;
	wire [4-1:0] node22417;
	wire [4-1:0] node22418;
	wire [4-1:0] node22419;
	wire [4-1:0] node22422;
	wire [4-1:0] node22426;
	wire [4-1:0] node22427;
	wire [4-1:0] node22428;
	wire [4-1:0] node22429;
	wire [4-1:0] node22430;
	wire [4-1:0] node22434;
	wire [4-1:0] node22436;
	wire [4-1:0] node22439;
	wire [4-1:0] node22441;
	wire [4-1:0] node22444;
	wire [4-1:0] node22445;
	wire [4-1:0] node22446;
	wire [4-1:0] node22448;
	wire [4-1:0] node22452;
	wire [4-1:0] node22453;
	wire [4-1:0] node22456;
	wire [4-1:0] node22459;
	wire [4-1:0] node22460;
	wire [4-1:0] node22461;
	wire [4-1:0] node22462;
	wire [4-1:0] node22463;
	wire [4-1:0] node22464;
	wire [4-1:0] node22465;
	wire [4-1:0] node22468;
	wire [4-1:0] node22470;
	wire [4-1:0] node22473;
	wire [4-1:0] node22474;
	wire [4-1:0] node22477;
	wire [4-1:0] node22479;
	wire [4-1:0] node22482;
	wire [4-1:0] node22483;
	wire [4-1:0] node22484;
	wire [4-1:0] node22485;
	wire [4-1:0] node22489;
	wire [4-1:0] node22490;
	wire [4-1:0] node22492;
	wire [4-1:0] node22495;
	wire [4-1:0] node22496;
	wire [4-1:0] node22499;
	wire [4-1:0] node22502;
	wire [4-1:0] node22503;
	wire [4-1:0] node22504;
	wire [4-1:0] node22505;
	wire [4-1:0] node22509;
	wire [4-1:0] node22510;
	wire [4-1:0] node22513;
	wire [4-1:0] node22516;
	wire [4-1:0] node22517;
	wire [4-1:0] node22519;
	wire [4-1:0] node22523;
	wire [4-1:0] node22524;
	wire [4-1:0] node22525;
	wire [4-1:0] node22527;
	wire [4-1:0] node22530;
	wire [4-1:0] node22532;
	wire [4-1:0] node22535;
	wire [4-1:0] node22536;
	wire [4-1:0] node22538;
	wire [4-1:0] node22541;
	wire [4-1:0] node22543;
	wire [4-1:0] node22546;
	wire [4-1:0] node22547;
	wire [4-1:0] node22548;
	wire [4-1:0] node22549;
	wire [4-1:0] node22551;
	wire [4-1:0] node22552;
	wire [4-1:0] node22555;
	wire [4-1:0] node22558;
	wire [4-1:0] node22559;
	wire [4-1:0] node22560;
	wire [4-1:0] node22561;
	wire [4-1:0] node22564;
	wire [4-1:0] node22567;
	wire [4-1:0] node22569;
	wire [4-1:0] node22572;
	wire [4-1:0] node22573;
	wire [4-1:0] node22575;
	wire [4-1:0] node22578;
	wire [4-1:0] node22579;
	wire [4-1:0] node22582;
	wire [4-1:0] node22585;
	wire [4-1:0] node22586;
	wire [4-1:0] node22587;
	wire [4-1:0] node22589;
	wire [4-1:0] node22590;
	wire [4-1:0] node22594;
	wire [4-1:0] node22595;
	wire [4-1:0] node22598;
	wire [4-1:0] node22601;
	wire [4-1:0] node22602;
	wire [4-1:0] node22604;
	wire [4-1:0] node22607;
	wire [4-1:0] node22608;
	wire [4-1:0] node22609;
	wire [4-1:0] node22613;
	wire [4-1:0] node22614;
	wire [4-1:0] node22618;
	wire [4-1:0] node22619;
	wire [4-1:0] node22620;
	wire [4-1:0] node22621;
	wire [4-1:0] node22625;
	wire [4-1:0] node22628;
	wire [4-1:0] node22629;
	wire [4-1:0] node22630;
	wire [4-1:0] node22634;
	wire [4-1:0] node22635;
	wire [4-1:0] node22639;
	wire [4-1:0] node22640;
	wire [4-1:0] node22641;
	wire [4-1:0] node22642;
	wire [4-1:0] node22643;
	wire [4-1:0] node22644;
	wire [4-1:0] node22646;
	wire [4-1:0] node22649;
	wire [4-1:0] node22651;
	wire [4-1:0] node22654;
	wire [4-1:0] node22655;
	wire [4-1:0] node22659;
	wire [4-1:0] node22660;
	wire [4-1:0] node22661;
	wire [4-1:0] node22662;
	wire [4-1:0] node22665;
	wire [4-1:0] node22669;
	wire [4-1:0] node22670;
	wire [4-1:0] node22671;
	wire [4-1:0] node22675;
	wire [4-1:0] node22676;
	wire [4-1:0] node22680;
	wire [4-1:0] node22681;
	wire [4-1:0] node22682;
	wire [4-1:0] node22683;
	wire [4-1:0] node22687;
	wire [4-1:0] node22688;
	wire [4-1:0] node22692;
	wire [4-1:0] node22693;
	wire [4-1:0] node22694;
	wire [4-1:0] node22698;
	wire [4-1:0] node22699;
	wire [4-1:0] node22703;
	wire [4-1:0] node22704;
	wire [4-1:0] node22705;
	wire [4-1:0] node22706;
	wire [4-1:0] node22707;
	wire [4-1:0] node22708;
	wire [4-1:0] node22709;
	wire [4-1:0] node22712;
	wire [4-1:0] node22715;
	wire [4-1:0] node22716;
	wire [4-1:0] node22719;
	wire [4-1:0] node22722;
	wire [4-1:0] node22724;
	wire [4-1:0] node22725;
	wire [4-1:0] node22728;
	wire [4-1:0] node22731;
	wire [4-1:0] node22732;
	wire [4-1:0] node22735;
	wire [4-1:0] node22738;
	wire [4-1:0] node22739;
	wire [4-1:0] node22740;
	wire [4-1:0] node22741;
	wire [4-1:0] node22745;
	wire [4-1:0] node22747;
	wire [4-1:0] node22750;
	wire [4-1:0] node22751;
	wire [4-1:0] node22752;
	wire [4-1:0] node22755;
	wire [4-1:0] node22758;
	wire [4-1:0] node22759;
	wire [4-1:0] node22762;
	wire [4-1:0] node22765;
	wire [4-1:0] node22766;
	wire [4-1:0] node22767;
	wire [4-1:0] node22768;
	wire [4-1:0] node22771;
	wire [4-1:0] node22774;
	wire [4-1:0] node22775;
	wire [4-1:0] node22778;
	wire [4-1:0] node22781;
	wire [4-1:0] node22782;
	wire [4-1:0] node22785;
	wire [4-1:0] node22788;
	wire [4-1:0] node22789;
	wire [4-1:0] node22790;
	wire [4-1:0] node22791;
	wire [4-1:0] node22792;
	wire [4-1:0] node22793;
	wire [4-1:0] node22794;
	wire [4-1:0] node22795;
	wire [4-1:0] node22796;
	wire [4-1:0] node22797;
	wire [4-1:0] node22801;
	wire [4-1:0] node22802;
	wire [4-1:0] node22803;
	wire [4-1:0] node22807;
	wire [4-1:0] node22808;
	wire [4-1:0] node22812;
	wire [4-1:0] node22814;
	wire [4-1:0] node22815;
	wire [4-1:0] node22818;
	wire [4-1:0] node22821;
	wire [4-1:0] node22822;
	wire [4-1:0] node22823;
	wire [4-1:0] node22825;
	wire [4-1:0] node22828;
	wire [4-1:0] node22830;
	wire [4-1:0] node22833;
	wire [4-1:0] node22834;
	wire [4-1:0] node22835;
	wire [4-1:0] node22838;
	wire [4-1:0] node22841;
	wire [4-1:0] node22842;
	wire [4-1:0] node22845;
	wire [4-1:0] node22847;
	wire [4-1:0] node22850;
	wire [4-1:0] node22851;
	wire [4-1:0] node22852;
	wire [4-1:0] node22853;
	wire [4-1:0] node22854;
	wire [4-1:0] node22855;
	wire [4-1:0] node22859;
	wire [4-1:0] node22860;
	wire [4-1:0] node22863;
	wire [4-1:0] node22866;
	wire [4-1:0] node22868;
	wire [4-1:0] node22870;
	wire [4-1:0] node22873;
	wire [4-1:0] node22874;
	wire [4-1:0] node22875;
	wire [4-1:0] node22878;
	wire [4-1:0] node22881;
	wire [4-1:0] node22882;
	wire [4-1:0] node22883;
	wire [4-1:0] node22888;
	wire [4-1:0] node22889;
	wire [4-1:0] node22890;
	wire [4-1:0] node22891;
	wire [4-1:0] node22894;
	wire [4-1:0] node22897;
	wire [4-1:0] node22898;
	wire [4-1:0] node22899;
	wire [4-1:0] node22902;
	wire [4-1:0] node22905;
	wire [4-1:0] node22906;
	wire [4-1:0] node22909;
	wire [4-1:0] node22912;
	wire [4-1:0] node22913;
	wire [4-1:0] node22914;
	wire [4-1:0] node22917;
	wire [4-1:0] node22920;
	wire [4-1:0] node22921;
	wire [4-1:0] node22922;
	wire [4-1:0] node22926;
	wire [4-1:0] node22929;
	wire [4-1:0] node22930;
	wire [4-1:0] node22931;
	wire [4-1:0] node22932;
	wire [4-1:0] node22933;
	wire [4-1:0] node22934;
	wire [4-1:0] node22935;
	wire [4-1:0] node22940;
	wire [4-1:0] node22941;
	wire [4-1:0] node22942;
	wire [4-1:0] node22946;
	wire [4-1:0] node22947;
	wire [4-1:0] node22950;
	wire [4-1:0] node22953;
	wire [4-1:0] node22954;
	wire [4-1:0] node22955;
	wire [4-1:0] node22957;
	wire [4-1:0] node22960;
	wire [4-1:0] node22961;
	wire [4-1:0] node22965;
	wire [4-1:0] node22966;
	wire [4-1:0] node22968;
	wire [4-1:0] node22971;
	wire [4-1:0] node22972;
	wire [4-1:0] node22976;
	wire [4-1:0] node22977;
	wire [4-1:0] node22978;
	wire [4-1:0] node22980;
	wire [4-1:0] node22981;
	wire [4-1:0] node22984;
	wire [4-1:0] node22987;
	wire [4-1:0] node22988;
	wire [4-1:0] node22991;
	wire [4-1:0] node22994;
	wire [4-1:0] node22995;
	wire [4-1:0] node22996;
	wire [4-1:0] node22997;
	wire [4-1:0] node23000;
	wire [4-1:0] node23003;
	wire [4-1:0] node23004;
	wire [4-1:0] node23008;
	wire [4-1:0] node23009;
	wire [4-1:0] node23012;
	wire [4-1:0] node23015;
	wire [4-1:0] node23016;
	wire [4-1:0] node23017;
	wire [4-1:0] node23018;
	wire [4-1:0] node23019;
	wire [4-1:0] node23020;
	wire [4-1:0] node23024;
	wire [4-1:0] node23025;
	wire [4-1:0] node23028;
	wire [4-1:0] node23031;
	wire [4-1:0] node23032;
	wire [4-1:0] node23035;
	wire [4-1:0] node23038;
	wire [4-1:0] node23039;
	wire [4-1:0] node23040;
	wire [4-1:0] node23041;
	wire [4-1:0] node23044;
	wire [4-1:0] node23047;
	wire [4-1:0] node23048;
	wire [4-1:0] node23051;
	wire [4-1:0] node23054;
	wire [4-1:0] node23055;
	wire [4-1:0] node23058;
	wire [4-1:0] node23061;
	wire [4-1:0] node23062;
	wire [4-1:0] node23063;
	wire [4-1:0] node23066;
	wire [4-1:0] node23069;
	wire [4-1:0] node23070;
	wire [4-1:0] node23071;
	wire [4-1:0] node23074;
	wire [4-1:0] node23077;
	wire [4-1:0] node23078;
	wire [4-1:0] node23081;
	wire [4-1:0] node23084;
	wire [4-1:0] node23085;
	wire [4-1:0] node23086;
	wire [4-1:0] node23087;
	wire [4-1:0] node23088;
	wire [4-1:0] node23089;
	wire [4-1:0] node23090;
	wire [4-1:0] node23093;
	wire [4-1:0] node23096;
	wire [4-1:0] node23097;
	wire [4-1:0] node23098;
	wire [4-1:0] node23101;
	wire [4-1:0] node23104;
	wire [4-1:0] node23105;
	wire [4-1:0] node23109;
	wire [4-1:0] node23110;
	wire [4-1:0] node23111;
	wire [4-1:0] node23112;
	wire [4-1:0] node23115;
	wire [4-1:0] node23118;
	wire [4-1:0] node23120;
	wire [4-1:0] node23123;
	wire [4-1:0] node23125;
	wire [4-1:0] node23128;
	wire [4-1:0] node23129;
	wire [4-1:0] node23130;
	wire [4-1:0] node23131;
	wire [4-1:0] node23132;
	wire [4-1:0] node23136;
	wire [4-1:0] node23138;
	wire [4-1:0] node23141;
	wire [4-1:0] node23142;
	wire [4-1:0] node23143;
	wire [4-1:0] node23146;
	wire [4-1:0] node23149;
	wire [4-1:0] node23151;
	wire [4-1:0] node23154;
	wire [4-1:0] node23155;
	wire [4-1:0] node23156;
	wire [4-1:0] node23157;
	wire [4-1:0] node23160;
	wire [4-1:0] node23163;
	wire [4-1:0] node23164;
	wire [4-1:0] node23167;
	wire [4-1:0] node23170;
	wire [4-1:0] node23171;
	wire [4-1:0] node23172;
	wire [4-1:0] node23176;
	wire [4-1:0] node23177;
	wire [4-1:0] node23180;
	wire [4-1:0] node23183;
	wire [4-1:0] node23184;
	wire [4-1:0] node23185;
	wire [4-1:0] node23186;
	wire [4-1:0] node23187;
	wire [4-1:0] node23188;
	wire [4-1:0] node23191;
	wire [4-1:0] node23194;
	wire [4-1:0] node23196;
	wire [4-1:0] node23199;
	wire [4-1:0] node23201;
	wire [4-1:0] node23202;
	wire [4-1:0] node23205;
	wire [4-1:0] node23208;
	wire [4-1:0] node23209;
	wire [4-1:0] node23210;
	wire [4-1:0] node23213;
	wire [4-1:0] node23214;
	wire [4-1:0] node23217;
	wire [4-1:0] node23220;
	wire [4-1:0] node23222;
	wire [4-1:0] node23223;
	wire [4-1:0] node23226;
	wire [4-1:0] node23229;
	wire [4-1:0] node23230;
	wire [4-1:0] node23231;
	wire [4-1:0] node23232;
	wire [4-1:0] node23233;
	wire [4-1:0] node23236;
	wire [4-1:0] node23239;
	wire [4-1:0] node23240;
	wire [4-1:0] node23243;
	wire [4-1:0] node23246;
	wire [4-1:0] node23247;
	wire [4-1:0] node23248;
	wire [4-1:0] node23252;
	wire [4-1:0] node23255;
	wire [4-1:0] node23256;
	wire [4-1:0] node23257;
	wire [4-1:0] node23261;
	wire [4-1:0] node23262;
	wire [4-1:0] node23263;
	wire [4-1:0] node23266;
	wire [4-1:0] node23269;
	wire [4-1:0] node23272;
	wire [4-1:0] node23273;
	wire [4-1:0] node23274;
	wire [4-1:0] node23275;
	wire [4-1:0] node23276;
	wire [4-1:0] node23277;
	wire [4-1:0] node23279;
	wire [4-1:0] node23282;
	wire [4-1:0] node23285;
	wire [4-1:0] node23286;
	wire [4-1:0] node23288;
	wire [4-1:0] node23291;
	wire [4-1:0] node23293;
	wire [4-1:0] node23296;
	wire [4-1:0] node23297;
	wire [4-1:0] node23299;
	wire [4-1:0] node23300;
	wire [4-1:0] node23303;
	wire [4-1:0] node23306;
	wire [4-1:0] node23307;
	wire [4-1:0] node23308;
	wire [4-1:0] node23311;
	wire [4-1:0] node23314;
	wire [4-1:0] node23315;
	wire [4-1:0] node23318;
	wire [4-1:0] node23321;
	wire [4-1:0] node23322;
	wire [4-1:0] node23323;
	wire [4-1:0] node23324;
	wire [4-1:0] node23328;
	wire [4-1:0] node23329;
	wire [4-1:0] node23332;
	wire [4-1:0] node23335;
	wire [4-1:0] node23336;
	wire [4-1:0] node23337;
	wire [4-1:0] node23340;
	wire [4-1:0] node23343;
	wire [4-1:0] node23345;
	wire [4-1:0] node23348;
	wire [4-1:0] node23349;
	wire [4-1:0] node23350;
	wire [4-1:0] node23351;
	wire [4-1:0] node23352;
	wire [4-1:0] node23353;
	wire [4-1:0] node23357;
	wire [4-1:0] node23360;
	wire [4-1:0] node23361;
	wire [4-1:0] node23362;
	wire [4-1:0] node23366;
	wire [4-1:0] node23367;
	wire [4-1:0] node23371;
	wire [4-1:0] node23372;
	wire [4-1:0] node23373;
	wire [4-1:0] node23374;
	wire [4-1:0] node23378;
	wire [4-1:0] node23379;
	wire [4-1:0] node23383;
	wire [4-1:0] node23385;
	wire [4-1:0] node23388;
	wire [4-1:0] node23389;
	wire [4-1:0] node23390;
	wire [4-1:0] node23391;
	wire [4-1:0] node23394;
	wire [4-1:0] node23398;
	wire [4-1:0] node23399;
	wire [4-1:0] node23400;
	wire [4-1:0] node23404;
	wire [4-1:0] node23405;
	wire [4-1:0] node23409;
	wire [4-1:0] node23410;
	wire [4-1:0] node23411;
	wire [4-1:0] node23412;
	wire [4-1:0] node23413;
	wire [4-1:0] node23414;
	wire [4-1:0] node23416;
	wire [4-1:0] node23417;
	wire [4-1:0] node23418;
	wire [4-1:0] node23422;
	wire [4-1:0] node23423;
	wire [4-1:0] node23427;
	wire [4-1:0] node23428;
	wire [4-1:0] node23431;
	wire [4-1:0] node23433;
	wire [4-1:0] node23436;
	wire [4-1:0] node23437;
	wire [4-1:0] node23438;
	wire [4-1:0] node23441;
	wire [4-1:0] node23444;
	wire [4-1:0] node23445;
	wire [4-1:0] node23446;
	wire [4-1:0] node23447;
	wire [4-1:0] node23450;
	wire [4-1:0] node23454;
	wire [4-1:0] node23455;
	wire [4-1:0] node23458;
	wire [4-1:0] node23461;
	wire [4-1:0] node23462;
	wire [4-1:0] node23463;
	wire [4-1:0] node23466;
	wire [4-1:0] node23469;
	wire [4-1:0] node23470;
	wire [4-1:0] node23471;
	wire [4-1:0] node23474;
	wire [4-1:0] node23477;
	wire [4-1:0] node23478;
	wire [4-1:0] node23481;
	wire [4-1:0] node23484;
	wire [4-1:0] node23485;
	wire [4-1:0] node23486;
	wire [4-1:0] node23487;
	wire [4-1:0] node23488;
	wire [4-1:0] node23490;
	wire [4-1:0] node23493;
	wire [4-1:0] node23495;
	wire [4-1:0] node23498;
	wire [4-1:0] node23499;
	wire [4-1:0] node23501;
	wire [4-1:0] node23504;
	wire [4-1:0] node23506;
	wire [4-1:0] node23509;
	wire [4-1:0] node23510;
	wire [4-1:0] node23511;
	wire [4-1:0] node23512;
	wire [4-1:0] node23515;
	wire [4-1:0] node23518;
	wire [4-1:0] node23519;
	wire [4-1:0] node23522;
	wire [4-1:0] node23525;
	wire [4-1:0] node23526;
	wire [4-1:0] node23529;
	wire [4-1:0] node23532;
	wire [4-1:0] node23533;
	wire [4-1:0] node23534;
	wire [4-1:0] node23535;
	wire [4-1:0] node23536;
	wire [4-1:0] node23539;
	wire [4-1:0] node23542;
	wire [4-1:0] node23543;
	wire [4-1:0] node23546;
	wire [4-1:0] node23549;
	wire [4-1:0] node23550;
	wire [4-1:0] node23553;
	wire [4-1:0] node23556;
	wire [4-1:0] node23557;
	wire [4-1:0] node23558;
	wire [4-1:0] node23559;
	wire [4-1:0] node23560;
	wire [4-1:0] node23563;
	wire [4-1:0] node23567;
	wire [4-1:0] node23568;
	wire [4-1:0] node23571;
	wire [4-1:0] node23574;
	wire [4-1:0] node23575;
	wire [4-1:0] node23576;
	wire [4-1:0] node23577;
	wire [4-1:0] node23580;
	wire [4-1:0] node23584;
	wire [4-1:0] node23585;
	wire [4-1:0] node23588;
	wire [4-1:0] node23591;
	wire [4-1:0] node23592;
	wire [4-1:0] node23593;
	wire [4-1:0] node23594;
	wire [4-1:0] node23595;
	wire [4-1:0] node23596;
	wire [4-1:0] node23598;
	wire [4-1:0] node23601;
	wire [4-1:0] node23602;
	wire [4-1:0] node23603;
	wire [4-1:0] node23607;
	wire [4-1:0] node23609;
	wire [4-1:0] node23612;
	wire [4-1:0] node23613;
	wire [4-1:0] node23614;
	wire [4-1:0] node23618;
	wire [4-1:0] node23621;
	wire [4-1:0] node23622;
	wire [4-1:0] node23623;
	wire [4-1:0] node23625;
	wire [4-1:0] node23627;
	wire [4-1:0] node23630;
	wire [4-1:0] node23631;
	wire [4-1:0] node23632;
	wire [4-1:0] node23635;
	wire [4-1:0] node23638;
	wire [4-1:0] node23639;
	wire [4-1:0] node23642;
	wire [4-1:0] node23645;
	wire [4-1:0] node23646;
	wire [4-1:0] node23647;
	wire [4-1:0] node23648;
	wire [4-1:0] node23653;
	wire [4-1:0] node23655;
	wire [4-1:0] node23658;
	wire [4-1:0] node23659;
	wire [4-1:0] node23660;
	wire [4-1:0] node23661;
	wire [4-1:0] node23662;
	wire [4-1:0] node23663;
	wire [4-1:0] node23667;
	wire [4-1:0] node23668;
	wire [4-1:0] node23672;
	wire [4-1:0] node23673;
	wire [4-1:0] node23676;
	wire [4-1:0] node23677;
	wire [4-1:0] node23681;
	wire [4-1:0] node23682;
	wire [4-1:0] node23683;
	wire [4-1:0] node23684;
	wire [4-1:0] node23687;
	wire [4-1:0] node23690;
	wire [4-1:0] node23691;
	wire [4-1:0] node23694;
	wire [4-1:0] node23697;
	wire [4-1:0] node23698;
	wire [4-1:0] node23701;
	wire [4-1:0] node23704;
	wire [4-1:0] node23705;
	wire [4-1:0] node23706;
	wire [4-1:0] node23707;
	wire [4-1:0] node23711;
	wire [4-1:0] node23712;
	wire [4-1:0] node23713;
	wire [4-1:0] node23716;
	wire [4-1:0] node23720;
	wire [4-1:0] node23721;
	wire [4-1:0] node23724;
	wire [4-1:0] node23727;
	wire [4-1:0] node23728;
	wire [4-1:0] node23729;
	wire [4-1:0] node23730;
	wire [4-1:0] node23731;
	wire [4-1:0] node23732;
	wire [4-1:0] node23733;
	wire [4-1:0] node23736;
	wire [4-1:0] node23739;
	wire [4-1:0] node23740;
	wire [4-1:0] node23743;
	wire [4-1:0] node23746;
	wire [4-1:0] node23747;
	wire [4-1:0] node23748;
	wire [4-1:0] node23751;
	wire [4-1:0] node23754;
	wire [4-1:0] node23755;
	wire [4-1:0] node23758;
	wire [4-1:0] node23761;
	wire [4-1:0] node23762;
	wire [4-1:0] node23765;
	wire [4-1:0] node23768;
	wire [4-1:0] node23769;
	wire [4-1:0] node23770;
	wire [4-1:0] node23771;
	wire [4-1:0] node23774;
	wire [4-1:0] node23777;
	wire [4-1:0] node23778;
	wire [4-1:0] node23781;
	wire [4-1:0] node23784;
	wire [4-1:0] node23785;
	wire [4-1:0] node23787;
	wire [4-1:0] node23790;
	wire [4-1:0] node23791;
	wire [4-1:0] node23794;
	wire [4-1:0] node23797;
	wire [4-1:0] node23798;
	wire [4-1:0] node23799;
	wire [4-1:0] node23800;
	wire [4-1:0] node23801;
	wire [4-1:0] node23803;
	wire [4-1:0] node23806;
	wire [4-1:0] node23807;
	wire [4-1:0] node23810;
	wire [4-1:0] node23813;
	wire [4-1:0] node23814;
	wire [4-1:0] node23817;
	wire [4-1:0] node23820;
	wire [4-1:0] node23822;
	wire [4-1:0] node23825;
	wire [4-1:0] node23826;
	wire [4-1:0] node23829;
	wire [4-1:0] node23832;
	wire [4-1:0] node23833;
	wire [4-1:0] node23834;
	wire [4-1:0] node23835;
	wire [4-1:0] node23836;
	wire [4-1:0] node23837;
	wire [4-1:0] node23838;
	wire [4-1:0] node23839;
	wire [4-1:0] node23840;
	wire [4-1:0] node23843;
	wire [4-1:0] node23846;
	wire [4-1:0] node23847;
	wire [4-1:0] node23848;
	wire [4-1:0] node23851;
	wire [4-1:0] node23854;
	wire [4-1:0] node23856;
	wire [4-1:0] node23859;
	wire [4-1:0] node23860;
	wire [4-1:0] node23861;
	wire [4-1:0] node23862;
	wire [4-1:0] node23866;
	wire [4-1:0] node23868;
	wire [4-1:0] node23871;
	wire [4-1:0] node23873;
	wire [4-1:0] node23874;
	wire [4-1:0] node23877;
	wire [4-1:0] node23880;
	wire [4-1:0] node23881;
	wire [4-1:0] node23882;
	wire [4-1:0] node23884;
	wire [4-1:0] node23887;
	wire [4-1:0] node23889;
	wire [4-1:0] node23892;
	wire [4-1:0] node23893;
	wire [4-1:0] node23895;
	wire [4-1:0] node23899;
	wire [4-1:0] node23900;
	wire [4-1:0] node23901;
	wire [4-1:0] node23902;
	wire [4-1:0] node23903;
	wire [4-1:0] node23905;
	wire [4-1:0] node23908;
	wire [4-1:0] node23910;
	wire [4-1:0] node23913;
	wire [4-1:0] node23915;
	wire [4-1:0] node23917;
	wire [4-1:0] node23920;
	wire [4-1:0] node23921;
	wire [4-1:0] node23922;
	wire [4-1:0] node23926;
	wire [4-1:0] node23927;
	wire [4-1:0] node23929;
	wire [4-1:0] node23932;
	wire [4-1:0] node23935;
	wire [4-1:0] node23936;
	wire [4-1:0] node23938;
	wire [4-1:0] node23939;
	wire [4-1:0] node23942;
	wire [4-1:0] node23945;
	wire [4-1:0] node23946;
	wire [4-1:0] node23949;
	wire [4-1:0] node23952;
	wire [4-1:0] node23953;
	wire [4-1:0] node23954;
	wire [4-1:0] node23955;
	wire [4-1:0] node23956;
	wire [4-1:0] node23957;
	wire [4-1:0] node23960;
	wire [4-1:0] node23963;
	wire [4-1:0] node23964;
	wire [4-1:0] node23965;
	wire [4-1:0] node23968;
	wire [4-1:0] node23972;
	wire [4-1:0] node23973;
	wire [4-1:0] node23974;
	wire [4-1:0] node23975;
	wire [4-1:0] node23979;
	wire [4-1:0] node23982;
	wire [4-1:0] node23983;
	wire [4-1:0] node23984;
	wire [4-1:0] node23988;
	wire [4-1:0] node23989;
	wire [4-1:0] node23993;
	wire [4-1:0] node23994;
	wire [4-1:0] node23995;
	wire [4-1:0] node23996;
	wire [4-1:0] node23999;
	wire [4-1:0] node24002;
	wire [4-1:0] node24003;
	wire [4-1:0] node24006;
	wire [4-1:0] node24009;
	wire [4-1:0] node24010;
	wire [4-1:0] node24011;
	wire [4-1:0] node24013;
	wire [4-1:0] node24016;
	wire [4-1:0] node24017;
	wire [4-1:0] node24021;
	wire [4-1:0] node24022;
	wire [4-1:0] node24025;
	wire [4-1:0] node24028;
	wire [4-1:0] node24029;
	wire [4-1:0] node24030;
	wire [4-1:0] node24031;
	wire [4-1:0] node24032;
	wire [4-1:0] node24034;
	wire [4-1:0] node24038;
	wire [4-1:0] node24039;
	wire [4-1:0] node24042;
	wire [4-1:0] node24045;
	wire [4-1:0] node24046;
	wire [4-1:0] node24047;
	wire [4-1:0] node24048;
	wire [4-1:0] node24051;
	wire [4-1:0] node24055;
	wire [4-1:0] node24057;
	wire [4-1:0] node24060;
	wire [4-1:0] node24061;
	wire [4-1:0] node24062;
	wire [4-1:0] node24064;
	wire [4-1:0] node24065;
	wire [4-1:0] node24068;
	wire [4-1:0] node24071;
	wire [4-1:0] node24072;
	wire [4-1:0] node24075;
	wire [4-1:0] node24078;
	wire [4-1:0] node24079;
	wire [4-1:0] node24082;
	wire [4-1:0] node24085;
	wire [4-1:0] node24086;
	wire [4-1:0] node24087;
	wire [4-1:0] node24088;
	wire [4-1:0] node24089;
	wire [4-1:0] node24090;
	wire [4-1:0] node24091;
	wire [4-1:0] node24093;
	wire [4-1:0] node24097;
	wire [4-1:0] node24099;
	wire [4-1:0] node24102;
	wire [4-1:0] node24103;
	wire [4-1:0] node24104;
	wire [4-1:0] node24105;
	wire [4-1:0] node24110;
	wire [4-1:0] node24111;
	wire [4-1:0] node24113;
	wire [4-1:0] node24116;
	wire [4-1:0] node24118;
	wire [4-1:0] node24121;
	wire [4-1:0] node24122;
	wire [4-1:0] node24123;
	wire [4-1:0] node24124;
	wire [4-1:0] node24126;
	wire [4-1:0] node24129;
	wire [4-1:0] node24130;
	wire [4-1:0] node24134;
	wire [4-1:0] node24135;
	wire [4-1:0] node24138;
	wire [4-1:0] node24141;
	wire [4-1:0] node24142;
	wire [4-1:0] node24143;
	wire [4-1:0] node24144;
	wire [4-1:0] node24149;
	wire [4-1:0] node24150;
	wire [4-1:0] node24151;
	wire [4-1:0] node24156;
	wire [4-1:0] node24157;
	wire [4-1:0] node24158;
	wire [4-1:0] node24159;
	wire [4-1:0] node24160;
	wire [4-1:0] node24163;
	wire [4-1:0] node24164;
	wire [4-1:0] node24167;
	wire [4-1:0] node24170;
	wire [4-1:0] node24171;
	wire [4-1:0] node24174;
	wire [4-1:0] node24176;
	wire [4-1:0] node24179;
	wire [4-1:0] node24180;
	wire [4-1:0] node24181;
	wire [4-1:0] node24182;
	wire [4-1:0] node24185;
	wire [4-1:0] node24188;
	wire [4-1:0] node24189;
	wire [4-1:0] node24192;
	wire [4-1:0] node24195;
	wire [4-1:0] node24196;
	wire [4-1:0] node24197;
	wire [4-1:0] node24200;
	wire [4-1:0] node24204;
	wire [4-1:0] node24205;
	wire [4-1:0] node24206;
	wire [4-1:0] node24208;
	wire [4-1:0] node24211;
	wire [4-1:0] node24214;
	wire [4-1:0] node24215;
	wire [4-1:0] node24216;
	wire [4-1:0] node24219;
	wire [4-1:0] node24222;
	wire [4-1:0] node24224;
	wire [4-1:0] node24225;
	wire [4-1:0] node24228;
	wire [4-1:0] node24231;
	wire [4-1:0] node24232;
	wire [4-1:0] node24233;
	wire [4-1:0] node24234;
	wire [4-1:0] node24235;
	wire [4-1:0] node24236;
	wire [4-1:0] node24237;
	wire [4-1:0] node24241;
	wire [4-1:0] node24244;
	wire [4-1:0] node24245;
	wire [4-1:0] node24248;
	wire [4-1:0] node24251;
	wire [4-1:0] node24252;
	wire [4-1:0] node24253;
	wire [4-1:0] node24254;
	wire [4-1:0] node24257;
	wire [4-1:0] node24261;
	wire [4-1:0] node24262;
	wire [4-1:0] node24265;
	wire [4-1:0] node24266;
	wire [4-1:0] node24270;
	wire [4-1:0] node24271;
	wire [4-1:0] node24272;
	wire [4-1:0] node24274;
	wire [4-1:0] node24275;
	wire [4-1:0] node24278;
	wire [4-1:0] node24281;
	wire [4-1:0] node24282;
	wire [4-1:0] node24283;
	wire [4-1:0] node24286;
	wire [4-1:0] node24290;
	wire [4-1:0] node24291;
	wire [4-1:0] node24292;
	wire [4-1:0] node24294;
	wire [4-1:0] node24297;
	wire [4-1:0] node24298;
	wire [4-1:0] node24301;
	wire [4-1:0] node24304;
	wire [4-1:0] node24305;
	wire [4-1:0] node24306;
	wire [4-1:0] node24311;
	wire [4-1:0] node24312;
	wire [4-1:0] node24313;
	wire [4-1:0] node24314;
	wire [4-1:0] node24316;
	wire [4-1:0] node24317;
	wire [4-1:0] node24321;
	wire [4-1:0] node24322;
	wire [4-1:0] node24323;
	wire [4-1:0] node24326;
	wire [4-1:0] node24329;
	wire [4-1:0] node24330;
	wire [4-1:0] node24334;
	wire [4-1:0] node24335;
	wire [4-1:0] node24337;
	wire [4-1:0] node24340;
	wire [4-1:0] node24341;
	wire [4-1:0] node24343;
	wire [4-1:0] node24346;
	wire [4-1:0] node24347;
	wire [4-1:0] node24350;
	wire [4-1:0] node24353;
	wire [4-1:0] node24354;
	wire [4-1:0] node24355;
	wire [4-1:0] node24356;
	wire [4-1:0] node24359;
	wire [4-1:0] node24362;
	wire [4-1:0] node24363;
	wire [4-1:0] node24364;
	wire [4-1:0] node24367;
	wire [4-1:0] node24370;
	wire [4-1:0] node24372;
	wire [4-1:0] node24375;
	wire [4-1:0] node24376;
	wire [4-1:0] node24379;
	wire [4-1:0] node24382;
	wire [4-1:0] node24383;
	wire [4-1:0] node24384;
	wire [4-1:0] node24385;
	wire [4-1:0] node24386;
	wire [4-1:0] node24387;
	wire [4-1:0] node24388;
	wire [4-1:0] node24389;
	wire [4-1:0] node24393;
	wire [4-1:0] node24394;
	wire [4-1:0] node24397;
	wire [4-1:0] node24400;
	wire [4-1:0] node24401;
	wire [4-1:0] node24402;
	wire [4-1:0] node24405;
	wire [4-1:0] node24408;
	wire [4-1:0] node24409;
	wire [4-1:0] node24410;
	wire [4-1:0] node24413;
	wire [4-1:0] node24416;
	wire [4-1:0] node24418;
	wire [4-1:0] node24421;
	wire [4-1:0] node24422;
	wire [4-1:0] node24423;
	wire [4-1:0] node24426;
	wire [4-1:0] node24428;
	wire [4-1:0] node24431;
	wire [4-1:0] node24432;
	wire [4-1:0] node24433;
	wire [4-1:0] node24434;
	wire [4-1:0] node24439;
	wire [4-1:0] node24440;
	wire [4-1:0] node24441;
	wire [4-1:0] node24445;
	wire [4-1:0] node24446;
	wire [4-1:0] node24450;
	wire [4-1:0] node24451;
	wire [4-1:0] node24452;
	wire [4-1:0] node24453;
	wire [4-1:0] node24454;
	wire [4-1:0] node24457;
	wire [4-1:0] node24460;
	wire [4-1:0] node24461;
	wire [4-1:0] node24464;
	wire [4-1:0] node24467;
	wire [4-1:0] node24468;
	wire [4-1:0] node24469;
	wire [4-1:0] node24472;
	wire [4-1:0] node24475;
	wire [4-1:0] node24476;
	wire [4-1:0] node24477;
	wire [4-1:0] node24480;
	wire [4-1:0] node24483;
	wire [4-1:0] node24484;
	wire [4-1:0] node24487;
	wire [4-1:0] node24490;
	wire [4-1:0] node24491;
	wire [4-1:0] node24492;
	wire [4-1:0] node24494;
	wire [4-1:0] node24495;
	wire [4-1:0] node24498;
	wire [4-1:0] node24501;
	wire [4-1:0] node24502;
	wire [4-1:0] node24503;
	wire [4-1:0] node24507;
	wire [4-1:0] node24509;
	wire [4-1:0] node24512;
	wire [4-1:0] node24513;
	wire [4-1:0] node24514;
	wire [4-1:0] node24518;
	wire [4-1:0] node24521;
	wire [4-1:0] node24522;
	wire [4-1:0] node24523;
	wire [4-1:0] node24524;
	wire [4-1:0] node24525;
	wire [4-1:0] node24528;
	wire [4-1:0] node24531;
	wire [4-1:0] node24532;
	wire [4-1:0] node24533;
	wire [4-1:0] node24535;
	wire [4-1:0] node24538;
	wire [4-1:0] node24539;
	wire [4-1:0] node24542;
	wire [4-1:0] node24545;
	wire [4-1:0] node24546;
	wire [4-1:0] node24549;
	wire [4-1:0] node24552;
	wire [4-1:0] node24553;
	wire [4-1:0] node24554;
	wire [4-1:0] node24555;
	wire [4-1:0] node24558;
	wire [4-1:0] node24562;
	wire [4-1:0] node24563;
	wire [4-1:0] node24564;
	wire [4-1:0] node24568;
	wire [4-1:0] node24569;
	wire [4-1:0] node24572;
	wire [4-1:0] node24575;
	wire [4-1:0] node24576;
	wire [4-1:0] node24577;
	wire [4-1:0] node24578;
	wire [4-1:0] node24579;
	wire [4-1:0] node24583;
	wire [4-1:0] node24584;
	wire [4-1:0] node24587;
	wire [4-1:0] node24590;
	wire [4-1:0] node24591;
	wire [4-1:0] node24592;
	wire [4-1:0] node24595;
	wire [4-1:0] node24598;
	wire [4-1:0] node24599;
	wire [4-1:0] node24602;
	wire [4-1:0] node24605;
	wire [4-1:0] node24606;
	wire [4-1:0] node24607;
	wire [4-1:0] node24609;
	wire [4-1:0] node24610;
	wire [4-1:0] node24613;
	wire [4-1:0] node24616;
	wire [4-1:0] node24617;
	wire [4-1:0] node24620;
	wire [4-1:0] node24623;
	wire [4-1:0] node24624;
	wire [4-1:0] node24625;
	wire [4-1:0] node24626;
	wire [4-1:0] node24629;
	wire [4-1:0] node24632;
	wire [4-1:0] node24633;
	wire [4-1:0] node24636;
	wire [4-1:0] node24639;
	wire [4-1:0] node24641;
	wire [4-1:0] node24644;
	wire [4-1:0] node24645;
	wire [4-1:0] node24646;
	wire [4-1:0] node24647;
	wire [4-1:0] node24648;
	wire [4-1:0] node24649;
	wire [4-1:0] node24651;
	wire [4-1:0] node24654;
	wire [4-1:0] node24656;
	wire [4-1:0] node24659;
	wire [4-1:0] node24661;
	wire [4-1:0] node24663;
	wire [4-1:0] node24666;
	wire [4-1:0] node24667;
	wire [4-1:0] node24668;
	wire [4-1:0] node24671;
	wire [4-1:0] node24673;
	wire [4-1:0] node24676;
	wire [4-1:0] node24677;
	wire [4-1:0] node24681;
	wire [4-1:0] node24682;
	wire [4-1:0] node24683;
	wire [4-1:0] node24684;
	wire [4-1:0] node24688;
	wire [4-1:0] node24689;
	wire [4-1:0] node24693;
	wire [4-1:0] node24694;
	wire [4-1:0] node24695;
	wire [4-1:0] node24699;
	wire [4-1:0] node24700;
	wire [4-1:0] node24704;
	wire [4-1:0] node24705;
	wire [4-1:0] node24706;
	wire [4-1:0] node24707;
	wire [4-1:0] node24708;
	wire [4-1:0] node24712;
	wire [4-1:0] node24713;
	wire [4-1:0] node24717;
	wire [4-1:0] node24718;
	wire [4-1:0] node24719;
	wire [4-1:0] node24723;
	wire [4-1:0] node24724;
	wire [4-1:0] node24728;
	wire [4-1:0] node24729;
	wire [4-1:0] node24730;
	wire [4-1:0] node24731;
	wire [4-1:0] node24732;
	wire [4-1:0] node24736;
	wire [4-1:0] node24737;
	wire [4-1:0] node24741;
	wire [4-1:0] node24742;
	wire [4-1:0] node24743;
	wire [4-1:0] node24748;
	wire [4-1:0] node24749;
	wire [4-1:0] node24750;
	wire [4-1:0] node24751;
	wire [4-1:0] node24752;
	wire [4-1:0] node24755;
	wire [4-1:0] node24759;
	wire [4-1:0] node24760;
	wire [4-1:0] node24763;
	wire [4-1:0] node24766;
	wire [4-1:0] node24767;
	wire [4-1:0] node24768;
	wire [4-1:0] node24769;
	wire [4-1:0] node24772;
	wire [4-1:0] node24775;
	wire [4-1:0] node24777;
	wire [4-1:0] node24780;
	wire [4-1:0] node24781;
	wire [4-1:0] node24785;
	wire [4-1:0] node24786;
	wire [4-1:0] node24787;
	wire [4-1:0] node24788;
	wire [4-1:0] node24789;
	wire [4-1:0] node24790;
	wire [4-1:0] node24791;
	wire [4-1:0] node24792;
	wire [4-1:0] node24793;
	wire [4-1:0] node24794;
	wire [4-1:0] node24795;
	wire [4-1:0] node24797;
	wire [4-1:0] node24800;
	wire [4-1:0] node24803;
	wire [4-1:0] node24804;
	wire [4-1:0] node24806;
	wire [4-1:0] node24809;
	wire [4-1:0] node24810;
	wire [4-1:0] node24814;
	wire [4-1:0] node24815;
	wire [4-1:0] node24816;
	wire [4-1:0] node24817;
	wire [4-1:0] node24821;
	wire [4-1:0] node24822;
	wire [4-1:0] node24825;
	wire [4-1:0] node24827;
	wire [4-1:0] node24830;
	wire [4-1:0] node24831;
	wire [4-1:0] node24832;
	wire [4-1:0] node24834;
	wire [4-1:0] node24837;
	wire [4-1:0] node24840;
	wire [4-1:0] node24842;
	wire [4-1:0] node24845;
	wire [4-1:0] node24846;
	wire [4-1:0] node24847;
	wire [4-1:0] node24848;
	wire [4-1:0] node24849;
	wire [4-1:0] node24853;
	wire [4-1:0] node24854;
	wire [4-1:0] node24855;
	wire [4-1:0] node24859;
	wire [4-1:0] node24861;
	wire [4-1:0] node24864;
	wire [4-1:0] node24865;
	wire [4-1:0] node24866;
	wire [4-1:0] node24868;
	wire [4-1:0] node24871;
	wire [4-1:0] node24873;
	wire [4-1:0] node24876;
	wire [4-1:0] node24877;
	wire [4-1:0] node24881;
	wire [4-1:0] node24882;
	wire [4-1:0] node24883;
	wire [4-1:0] node24885;
	wire [4-1:0] node24887;
	wire [4-1:0] node24890;
	wire [4-1:0] node24891;
	wire [4-1:0] node24894;
	wire [4-1:0] node24897;
	wire [4-1:0] node24898;
	wire [4-1:0] node24899;
	wire [4-1:0] node24902;
	wire [4-1:0] node24905;
	wire [4-1:0] node24906;
	wire [4-1:0] node24908;
	wire [4-1:0] node24911;
	wire [4-1:0] node24912;
	wire [4-1:0] node24915;
	wire [4-1:0] node24918;
	wire [4-1:0] node24919;
	wire [4-1:0] node24920;
	wire [4-1:0] node24921;
	wire [4-1:0] node24922;
	wire [4-1:0] node24923;
	wire [4-1:0] node24925;
	wire [4-1:0] node24929;
	wire [4-1:0] node24930;
	wire [4-1:0] node24934;
	wire [4-1:0] node24935;
	wire [4-1:0] node24937;
	wire [4-1:0] node24939;
	wire [4-1:0] node24942;
	wire [4-1:0] node24943;
	wire [4-1:0] node24947;
	wire [4-1:0] node24948;
	wire [4-1:0] node24949;
	wire [4-1:0] node24950;
	wire [4-1:0] node24952;
	wire [4-1:0] node24955;
	wire [4-1:0] node24957;
	wire [4-1:0] node24960;
	wire [4-1:0] node24962;
	wire [4-1:0] node24963;
	wire [4-1:0] node24966;
	wire [4-1:0] node24969;
	wire [4-1:0] node24970;
	wire [4-1:0] node24971;
	wire [4-1:0] node24973;
	wire [4-1:0] node24977;
	wire [4-1:0] node24978;
	wire [4-1:0] node24982;
	wire [4-1:0] node24983;
	wire [4-1:0] node24984;
	wire [4-1:0] node24985;
	wire [4-1:0] node24987;
	wire [4-1:0] node24988;
	wire [4-1:0] node24991;
	wire [4-1:0] node24994;
	wire [4-1:0] node24995;
	wire [4-1:0] node24996;
	wire [4-1:0] node24999;
	wire [4-1:0] node25002;
	wire [4-1:0] node25003;
	wire [4-1:0] node25006;
	wire [4-1:0] node25009;
	wire [4-1:0] node25010;
	wire [4-1:0] node25011;
	wire [4-1:0] node25013;
	wire [4-1:0] node25016;
	wire [4-1:0] node25018;
	wire [4-1:0] node25021;
	wire [4-1:0] node25022;
	wire [4-1:0] node25026;
	wire [4-1:0] node25027;
	wire [4-1:0] node25028;
	wire [4-1:0] node25029;
	wire [4-1:0] node25031;
	wire [4-1:0] node25035;
	wire [4-1:0] node25037;
	wire [4-1:0] node25039;
	wire [4-1:0] node25042;
	wire [4-1:0] node25043;
	wire [4-1:0] node25044;
	wire [4-1:0] node25046;
	wire [4-1:0] node25049;
	wire [4-1:0] node25052;
	wire [4-1:0] node25053;
	wire [4-1:0] node25056;
	wire [4-1:0] node25058;
	wire [4-1:0] node25061;
	wire [4-1:0] node25062;
	wire [4-1:0] node25063;
	wire [4-1:0] node25064;
	wire [4-1:0] node25065;
	wire [4-1:0] node25067;
	wire [4-1:0] node25070;
	wire [4-1:0] node25071;
	wire [4-1:0] node25072;
	wire [4-1:0] node25073;
	wire [4-1:0] node25076;
	wire [4-1:0] node25080;
	wire [4-1:0] node25081;
	wire [4-1:0] node25084;
	wire [4-1:0] node25087;
	wire [4-1:0] node25088;
	wire [4-1:0] node25089;
	wire [4-1:0] node25090;
	wire [4-1:0] node25093;
	wire [4-1:0] node25097;
	wire [4-1:0] node25098;
	wire [4-1:0] node25100;
	wire [4-1:0] node25103;
	wire [4-1:0] node25104;
	wire [4-1:0] node25107;
	wire [4-1:0] node25110;
	wire [4-1:0] node25111;
	wire [4-1:0] node25112;
	wire [4-1:0] node25113;
	wire [4-1:0] node25116;
	wire [4-1:0] node25118;
	wire [4-1:0] node25121;
	wire [4-1:0] node25122;
	wire [4-1:0] node25123;
	wire [4-1:0] node25127;
	wire [4-1:0] node25128;
	wire [4-1:0] node25129;
	wire [4-1:0] node25132;
	wire [4-1:0] node25135;
	wire [4-1:0] node25136;
	wire [4-1:0] node25139;
	wire [4-1:0] node25142;
	wire [4-1:0] node25143;
	wire [4-1:0] node25144;
	wire [4-1:0] node25147;
	wire [4-1:0] node25149;
	wire [4-1:0] node25152;
	wire [4-1:0] node25153;
	wire [4-1:0] node25154;
	wire [4-1:0] node25157;
	wire [4-1:0] node25160;
	wire [4-1:0] node25161;
	wire [4-1:0] node25164;
	wire [4-1:0] node25167;
	wire [4-1:0] node25168;
	wire [4-1:0] node25169;
	wire [4-1:0] node25170;
	wire [4-1:0] node25171;
	wire [4-1:0] node25172;
	wire [4-1:0] node25175;
	wire [4-1:0] node25178;
	wire [4-1:0] node25179;
	wire [4-1:0] node25180;
	wire [4-1:0] node25183;
	wire [4-1:0] node25186;
	wire [4-1:0] node25187;
	wire [4-1:0] node25190;
	wire [4-1:0] node25193;
	wire [4-1:0] node25194;
	wire [4-1:0] node25195;
	wire [4-1:0] node25196;
	wire [4-1:0] node25199;
	wire [4-1:0] node25202;
	wire [4-1:0] node25204;
	wire [4-1:0] node25207;
	wire [4-1:0] node25208;
	wire [4-1:0] node25211;
	wire [4-1:0] node25212;
	wire [4-1:0] node25215;
	wire [4-1:0] node25218;
	wire [4-1:0] node25219;
	wire [4-1:0] node25220;
	wire [4-1:0] node25221;
	wire [4-1:0] node25223;
	wire [4-1:0] node25226;
	wire [4-1:0] node25228;
	wire [4-1:0] node25231;
	wire [4-1:0] node25234;
	wire [4-1:0] node25235;
	wire [4-1:0] node25236;
	wire [4-1:0] node25237;
	wire [4-1:0] node25241;
	wire [4-1:0] node25244;
	wire [4-1:0] node25245;
	wire [4-1:0] node25246;
	wire [4-1:0] node25250;
	wire [4-1:0] node25251;
	wire [4-1:0] node25255;
	wire [4-1:0] node25256;
	wire [4-1:0] node25257;
	wire [4-1:0] node25258;
	wire [4-1:0] node25259;
	wire [4-1:0] node25260;
	wire [4-1:0] node25264;
	wire [4-1:0] node25265;
	wire [4-1:0] node25268;
	wire [4-1:0] node25271;
	wire [4-1:0] node25272;
	wire [4-1:0] node25273;
	wire [4-1:0] node25276;
	wire [4-1:0] node25279;
	wire [4-1:0] node25281;
	wire [4-1:0] node25284;
	wire [4-1:0] node25285;
	wire [4-1:0] node25286;
	wire [4-1:0] node25288;
	wire [4-1:0] node25292;
	wire [4-1:0] node25293;
	wire [4-1:0] node25294;
	wire [4-1:0] node25299;
	wire [4-1:0] node25300;
	wire [4-1:0] node25301;
	wire [4-1:0] node25302;
	wire [4-1:0] node25304;
	wire [4-1:0] node25308;
	wire [4-1:0] node25309;
	wire [4-1:0] node25312;
	wire [4-1:0] node25315;
	wire [4-1:0] node25316;
	wire [4-1:0] node25317;
	wire [4-1:0] node25318;
	wire [4-1:0] node25322;
	wire [4-1:0] node25323;
	wire [4-1:0] node25327;
	wire [4-1:0] node25328;
	wire [4-1:0] node25329;
	wire [4-1:0] node25332;
	wire [4-1:0] node25336;
	wire [4-1:0] node25337;
	wire [4-1:0] node25338;
	wire [4-1:0] node25339;
	wire [4-1:0] node25340;
	wire [4-1:0] node25341;
	wire [4-1:0] node25342;
	wire [4-1:0] node25345;
	wire [4-1:0] node25348;
	wire [4-1:0] node25349;
	wire [4-1:0] node25351;
	wire [4-1:0] node25352;
	wire [4-1:0] node25355;
	wire [4-1:0] node25358;
	wire [4-1:0] node25359;
	wire [4-1:0] node25360;
	wire [4-1:0] node25363;
	wire [4-1:0] node25366;
	wire [4-1:0] node25367;
	wire [4-1:0] node25370;
	wire [4-1:0] node25373;
	wire [4-1:0] node25374;
	wire [4-1:0] node25375;
	wire [4-1:0] node25377;
	wire [4-1:0] node25380;
	wire [4-1:0] node25382;
	wire [4-1:0] node25385;
	wire [4-1:0] node25386;
	wire [4-1:0] node25388;
	wire [4-1:0] node25391;
	wire [4-1:0] node25393;
	wire [4-1:0] node25396;
	wire [4-1:0] node25397;
	wire [4-1:0] node25398;
	wire [4-1:0] node25399;
	wire [4-1:0] node25401;
	wire [4-1:0] node25404;
	wire [4-1:0] node25406;
	wire [4-1:0] node25409;
	wire [4-1:0] node25410;
	wire [4-1:0] node25412;
	wire [4-1:0] node25415;
	wire [4-1:0] node25417;
	wire [4-1:0] node25420;
	wire [4-1:0] node25421;
	wire [4-1:0] node25422;
	wire [4-1:0] node25424;
	wire [4-1:0] node25427;
	wire [4-1:0] node25429;
	wire [4-1:0] node25432;
	wire [4-1:0] node25433;
	wire [4-1:0] node25435;
	wire [4-1:0] node25438;
	wire [4-1:0] node25440;
	wire [4-1:0] node25443;
	wire [4-1:0] node25444;
	wire [4-1:0] node25445;
	wire [4-1:0] node25446;
	wire [4-1:0] node25447;
	wire [4-1:0] node25448;
	wire [4-1:0] node25451;
	wire [4-1:0] node25454;
	wire [4-1:0] node25455;
	wire [4-1:0] node25458;
	wire [4-1:0] node25461;
	wire [4-1:0] node25462;
	wire [4-1:0] node25463;
	wire [4-1:0] node25466;
	wire [4-1:0] node25469;
	wire [4-1:0] node25470;
	wire [4-1:0] node25473;
	wire [4-1:0] node25476;
	wire [4-1:0] node25477;
	wire [4-1:0] node25478;
	wire [4-1:0] node25482;
	wire [4-1:0] node25483;
	wire [4-1:0] node25484;
	wire [4-1:0] node25487;
	wire [4-1:0] node25490;
	wire [4-1:0] node25491;
	wire [4-1:0] node25494;
	wire [4-1:0] node25497;
	wire [4-1:0] node25498;
	wire [4-1:0] node25499;
	wire [4-1:0] node25500;
	wire [4-1:0] node25502;
	wire [4-1:0] node25505;
	wire [4-1:0] node25507;
	wire [4-1:0] node25510;
	wire [4-1:0] node25511;
	wire [4-1:0] node25513;
	wire [4-1:0] node25516;
	wire [4-1:0] node25519;
	wire [4-1:0] node25520;
	wire [4-1:0] node25521;
	wire [4-1:0] node25522;
	wire [4-1:0] node25525;
	wire [4-1:0] node25528;
	wire [4-1:0] node25530;
	wire [4-1:0] node25531;
	wire [4-1:0] node25534;
	wire [4-1:0] node25537;
	wire [4-1:0] node25538;
	wire [4-1:0] node25539;
	wire [4-1:0] node25541;
	wire [4-1:0] node25544;
	wire [4-1:0] node25547;
	wire [4-1:0] node25548;
	wire [4-1:0] node25550;
	wire [4-1:0] node25553;
	wire [4-1:0] node25556;
	wire [4-1:0] node25557;
	wire [4-1:0] node25558;
	wire [4-1:0] node25559;
	wire [4-1:0] node25560;
	wire [4-1:0] node25561;
	wire [4-1:0] node25563;
	wire [4-1:0] node25566;
	wire [4-1:0] node25568;
	wire [4-1:0] node25571;
	wire [4-1:0] node25573;
	wire [4-1:0] node25574;
	wire [4-1:0] node25576;
	wire [4-1:0] node25579;
	wire [4-1:0] node25580;
	wire [4-1:0] node25584;
	wire [4-1:0] node25585;
	wire [4-1:0] node25586;
	wire [4-1:0] node25588;
	wire [4-1:0] node25591;
	wire [4-1:0] node25593;
	wire [4-1:0] node25596;
	wire [4-1:0] node25597;
	wire [4-1:0] node25599;
	wire [4-1:0] node25602;
	wire [4-1:0] node25604;
	wire [4-1:0] node25607;
	wire [4-1:0] node25608;
	wire [4-1:0] node25609;
	wire [4-1:0] node25610;
	wire [4-1:0] node25612;
	wire [4-1:0] node25615;
	wire [4-1:0] node25617;
	wire [4-1:0] node25620;
	wire [4-1:0] node25621;
	wire [4-1:0] node25624;
	wire [4-1:0] node25626;
	wire [4-1:0] node25629;
	wire [4-1:0] node25630;
	wire [4-1:0] node25631;
	wire [4-1:0] node25633;
	wire [4-1:0] node25636;
	wire [4-1:0] node25638;
	wire [4-1:0] node25641;
	wire [4-1:0] node25642;
	wire [4-1:0] node25644;
	wire [4-1:0] node25647;
	wire [4-1:0] node25649;
	wire [4-1:0] node25652;
	wire [4-1:0] node25653;
	wire [4-1:0] node25654;
	wire [4-1:0] node25655;
	wire [4-1:0] node25656;
	wire [4-1:0] node25658;
	wire [4-1:0] node25661;
	wire [4-1:0] node25663;
	wire [4-1:0] node25666;
	wire [4-1:0] node25667;
	wire [4-1:0] node25669;
	wire [4-1:0] node25673;
	wire [4-1:0] node25674;
	wire [4-1:0] node25675;
	wire [4-1:0] node25677;
	wire [4-1:0] node25680;
	wire [4-1:0] node25682;
	wire [4-1:0] node25685;
	wire [4-1:0] node25686;
	wire [4-1:0] node25688;
	wire [4-1:0] node25691;
	wire [4-1:0] node25693;
	wire [4-1:0] node25696;
	wire [4-1:0] node25697;
	wire [4-1:0] node25698;
	wire [4-1:0] node25699;
	wire [4-1:0] node25701;
	wire [4-1:0] node25704;
	wire [4-1:0] node25706;
	wire [4-1:0] node25709;
	wire [4-1:0] node25710;
	wire [4-1:0] node25712;
	wire [4-1:0] node25715;
	wire [4-1:0] node25717;
	wire [4-1:0] node25720;
	wire [4-1:0] node25721;
	wire [4-1:0] node25722;
	wire [4-1:0] node25723;
	wire [4-1:0] node25726;
	wire [4-1:0] node25729;
	wire [4-1:0] node25730;
	wire [4-1:0] node25732;
	wire [4-1:0] node25735;
	wire [4-1:0] node25737;
	wire [4-1:0] node25740;
	wire [4-1:0] node25741;
	wire [4-1:0] node25742;
	wire [4-1:0] node25745;
	wire [4-1:0] node25748;
	wire [4-1:0] node25749;
	wire [4-1:0] node25752;
	wire [4-1:0] node25755;
	wire [4-1:0] node25756;
	wire [4-1:0] node25757;
	wire [4-1:0] node25758;
	wire [4-1:0] node25759;
	wire [4-1:0] node25760;
	wire [4-1:0] node25761;
	wire [4-1:0] node25762;
	wire [4-1:0] node25763;
	wire [4-1:0] node25764;
	wire [4-1:0] node25768;
	wire [4-1:0] node25769;
	wire [4-1:0] node25772;
	wire [4-1:0] node25775;
	wire [4-1:0] node25777;
	wire [4-1:0] node25778;
	wire [4-1:0] node25781;
	wire [4-1:0] node25784;
	wire [4-1:0] node25785;
	wire [4-1:0] node25786;
	wire [4-1:0] node25789;
	wire [4-1:0] node25791;
	wire [4-1:0] node25794;
	wire [4-1:0] node25795;
	wire [4-1:0] node25799;
	wire [4-1:0] node25800;
	wire [4-1:0] node25801;
	wire [4-1:0] node25802;
	wire [4-1:0] node25804;
	wire [4-1:0] node25808;
	wire [4-1:0] node25809;
	wire [4-1:0] node25812;
	wire [4-1:0] node25814;
	wire [4-1:0] node25817;
	wire [4-1:0] node25818;
	wire [4-1:0] node25819;
	wire [4-1:0] node25821;
	wire [4-1:0] node25824;
	wire [4-1:0] node25826;
	wire [4-1:0] node25829;
	wire [4-1:0] node25831;
	wire [4-1:0] node25834;
	wire [4-1:0] node25835;
	wire [4-1:0] node25836;
	wire [4-1:0] node25837;
	wire [4-1:0] node25839;
	wire [4-1:0] node25842;
	wire [4-1:0] node25844;
	wire [4-1:0] node25847;
	wire [4-1:0] node25848;
	wire [4-1:0] node25850;
	wire [4-1:0] node25851;
	wire [4-1:0] node25855;
	wire [4-1:0] node25856;
	wire [4-1:0] node25858;
	wire [4-1:0] node25861;
	wire [4-1:0] node25863;
	wire [4-1:0] node25866;
	wire [4-1:0] node25867;
	wire [4-1:0] node25868;
	wire [4-1:0] node25869;
	wire [4-1:0] node25871;
	wire [4-1:0] node25874;
	wire [4-1:0] node25876;
	wire [4-1:0] node25879;
	wire [4-1:0] node25880;
	wire [4-1:0] node25883;
	wire [4-1:0] node25885;
	wire [4-1:0] node25888;
	wire [4-1:0] node25889;
	wire [4-1:0] node25890;
	wire [4-1:0] node25891;
	wire [4-1:0] node25894;
	wire [4-1:0] node25898;
	wire [4-1:0] node25899;
	wire [4-1:0] node25900;
	wire [4-1:0] node25903;
	wire [4-1:0] node25906;
	wire [4-1:0] node25908;
	wire [4-1:0] node25911;
	wire [4-1:0] node25912;
	wire [4-1:0] node25913;
	wire [4-1:0] node25914;
	wire [4-1:0] node25915;
	wire [4-1:0] node25918;
	wire [4-1:0] node25921;
	wire [4-1:0] node25922;
	wire [4-1:0] node25923;
	wire [4-1:0] node25925;
	wire [4-1:0] node25928;
	wire [4-1:0] node25929;
	wire [4-1:0] node25932;
	wire [4-1:0] node25935;
	wire [4-1:0] node25936;
	wire [4-1:0] node25937;
	wire [4-1:0] node25940;
	wire [4-1:0] node25944;
	wire [4-1:0] node25945;
	wire [4-1:0] node25946;
	wire [4-1:0] node25949;
	wire [4-1:0] node25952;
	wire [4-1:0] node25953;
	wire [4-1:0] node25955;
	wire [4-1:0] node25956;
	wire [4-1:0] node25960;
	wire [4-1:0] node25961;
	wire [4-1:0] node25964;
	wire [4-1:0] node25967;
	wire [4-1:0] node25968;
	wire [4-1:0] node25969;
	wire [4-1:0] node25970;
	wire [4-1:0] node25972;
	wire [4-1:0] node25974;
	wire [4-1:0] node25977;
	wire [4-1:0] node25978;
	wire [4-1:0] node25980;
	wire [4-1:0] node25983;
	wire [4-1:0] node25985;
	wire [4-1:0] node25988;
	wire [4-1:0] node25989;
	wire [4-1:0] node25990;
	wire [4-1:0] node25992;
	wire [4-1:0] node25995;
	wire [4-1:0] node25997;
	wire [4-1:0] node26000;
	wire [4-1:0] node26001;
	wire [4-1:0] node26005;
	wire [4-1:0] node26006;
	wire [4-1:0] node26007;
	wire [4-1:0] node26008;
	wire [4-1:0] node26010;
	wire [4-1:0] node26013;
	wire [4-1:0] node26015;
	wire [4-1:0] node26019;
	wire [4-1:0] node26020;
	wire [4-1:0] node26021;
	wire [4-1:0] node26024;
	wire [4-1:0] node26027;
	wire [4-1:0] node26029;
	wire [4-1:0] node26030;
	wire [4-1:0] node26033;
	wire [4-1:0] node26036;
	wire [4-1:0] node26037;
	wire [4-1:0] node26038;
	wire [4-1:0] node26039;
	wire [4-1:0] node26040;
	wire [4-1:0] node26041;
	wire [4-1:0] node26042;
	wire [4-1:0] node26045;
	wire [4-1:0] node26048;
	wire [4-1:0] node26049;
	wire [4-1:0] node26052;
	wire [4-1:0] node26055;
	wire [4-1:0] node26056;
	wire [4-1:0] node26057;
	wire [4-1:0] node26060;
	wire [4-1:0] node26063;
	wire [4-1:0] node26064;
	wire [4-1:0] node26067;
	wire [4-1:0] node26070;
	wire [4-1:0] node26071;
	wire [4-1:0] node26072;
	wire [4-1:0] node26073;
	wire [4-1:0] node26077;
	wire [4-1:0] node26078;
	wire [4-1:0] node26082;
	wire [4-1:0] node26083;
	wire [4-1:0] node26084;
	wire [4-1:0] node26085;
	wire [4-1:0] node26089;
	wire [4-1:0] node26090;
	wire [4-1:0] node26093;
	wire [4-1:0] node26096;
	wire [4-1:0] node26097;
	wire [4-1:0] node26100;
	wire [4-1:0] node26103;
	wire [4-1:0] node26104;
	wire [4-1:0] node26105;
	wire [4-1:0] node26106;
	wire [4-1:0] node26107;
	wire [4-1:0] node26110;
	wire [4-1:0] node26113;
	wire [4-1:0] node26114;
	wire [4-1:0] node26118;
	wire [4-1:0] node26119;
	wire [4-1:0] node26121;
	wire [4-1:0] node26122;
	wire [4-1:0] node26125;
	wire [4-1:0] node26128;
	wire [4-1:0] node26129;
	wire [4-1:0] node26131;
	wire [4-1:0] node26134;
	wire [4-1:0] node26135;
	wire [4-1:0] node26138;
	wire [4-1:0] node26141;
	wire [4-1:0] node26142;
	wire [4-1:0] node26143;
	wire [4-1:0] node26144;
	wire [4-1:0] node26145;
	wire [4-1:0] node26150;
	wire [4-1:0] node26151;
	wire [4-1:0] node26152;
	wire [4-1:0] node26155;
	wire [4-1:0] node26158;
	wire [4-1:0] node26160;
	wire [4-1:0] node26163;
	wire [4-1:0] node26164;
	wire [4-1:0] node26165;
	wire [4-1:0] node26168;
	wire [4-1:0] node26171;
	wire [4-1:0] node26172;
	wire [4-1:0] node26175;
	wire [4-1:0] node26178;
	wire [4-1:0] node26179;
	wire [4-1:0] node26180;
	wire [4-1:0] node26181;
	wire [4-1:0] node26182;
	wire [4-1:0] node26183;
	wire [4-1:0] node26185;
	wire [4-1:0] node26188;
	wire [4-1:0] node26189;
	wire [4-1:0] node26193;
	wire [4-1:0] node26195;
	wire [4-1:0] node26198;
	wire [4-1:0] node26199;
	wire [4-1:0] node26200;
	wire [4-1:0] node26204;
	wire [4-1:0] node26205;
	wire [4-1:0] node26208;
	wire [4-1:0] node26211;
	wire [4-1:0] node26212;
	wire [4-1:0] node26213;
	wire [4-1:0] node26215;
	wire [4-1:0] node26216;
	wire [4-1:0] node26219;
	wire [4-1:0] node26222;
	wire [4-1:0] node26224;
	wire [4-1:0] node26227;
	wire [4-1:0] node26228;
	wire [4-1:0] node26231;
	wire [4-1:0] node26234;
	wire [4-1:0] node26235;
	wire [4-1:0] node26236;
	wire [4-1:0] node26237;
	wire [4-1:0] node26238;
	wire [4-1:0] node26240;
	wire [4-1:0] node26244;
	wire [4-1:0] node26245;
	wire [4-1:0] node26248;
	wire [4-1:0] node26251;
	wire [4-1:0] node26252;
	wire [4-1:0] node26253;
	wire [4-1:0] node26256;
	wire [4-1:0] node26259;
	wire [4-1:0] node26260;
	wire [4-1:0] node26263;
	wire [4-1:0] node26266;
	wire [4-1:0] node26267;
	wire [4-1:0] node26268;
	wire [4-1:0] node26269;
	wire [4-1:0] node26273;
	wire [4-1:0] node26275;
	wire [4-1:0] node26276;
	wire [4-1:0] node26280;
	wire [4-1:0] node26281;
	wire [4-1:0] node26284;
	wire [4-1:0] node26287;
	wire [4-1:0] node26288;
	wire [4-1:0] node26289;
	wire [4-1:0] node26290;
	wire [4-1:0] node26291;
	wire [4-1:0] node26292;
	wire [4-1:0] node26293;
	wire [4-1:0] node26295;
	wire [4-1:0] node26299;
	wire [4-1:0] node26300;
	wire [4-1:0] node26302;
	wire [4-1:0] node26305;
	wire [4-1:0] node26307;
	wire [4-1:0] node26310;
	wire [4-1:0] node26311;
	wire [4-1:0] node26312;
	wire [4-1:0] node26313;
	wire [4-1:0] node26314;
	wire [4-1:0] node26317;
	wire [4-1:0] node26321;
	wire [4-1:0] node26323;
	wire [4-1:0] node26324;
	wire [4-1:0] node26328;
	wire [4-1:0] node26329;
	wire [4-1:0] node26330;
	wire [4-1:0] node26333;
	wire [4-1:0] node26335;
	wire [4-1:0] node26338;
	wire [4-1:0] node26339;
	wire [4-1:0] node26340;
	wire [4-1:0] node26343;
	wire [4-1:0] node26346;
	wire [4-1:0] node26347;
	wire [4-1:0] node26350;
	wire [4-1:0] node26353;
	wire [4-1:0] node26354;
	wire [4-1:0] node26355;
	wire [4-1:0] node26356;
	wire [4-1:0] node26359;
	wire [4-1:0] node26362;
	wire [4-1:0] node26363;
	wire [4-1:0] node26365;
	wire [4-1:0] node26369;
	wire [4-1:0] node26370;
	wire [4-1:0] node26371;
	wire [4-1:0] node26373;
	wire [4-1:0] node26376;
	wire [4-1:0] node26378;
	wire [4-1:0] node26380;
	wire [4-1:0] node26383;
	wire [4-1:0] node26384;
	wire [4-1:0] node26385;
	wire [4-1:0] node26388;
	wire [4-1:0] node26391;
	wire [4-1:0] node26393;
	wire [4-1:0] node26395;
	wire [4-1:0] node26398;
	wire [4-1:0] node26399;
	wire [4-1:0] node26400;
	wire [4-1:0] node26401;
	wire [4-1:0] node26403;
	wire [4-1:0] node26406;
	wire [4-1:0] node26408;
	wire [4-1:0] node26410;
	wire [4-1:0] node26411;
	wire [4-1:0] node26414;
	wire [4-1:0] node26417;
	wire [4-1:0] node26418;
	wire [4-1:0] node26419;
	wire [4-1:0] node26420;
	wire [4-1:0] node26422;
	wire [4-1:0] node26426;
	wire [4-1:0] node26427;
	wire [4-1:0] node26428;
	wire [4-1:0] node26431;
	wire [4-1:0] node26434;
	wire [4-1:0] node26435;
	wire [4-1:0] node26439;
	wire [4-1:0] node26440;
	wire [4-1:0] node26441;
	wire [4-1:0] node26444;
	wire [4-1:0] node26447;
	wire [4-1:0] node26448;
	wire [4-1:0] node26449;
	wire [4-1:0] node26452;
	wire [4-1:0] node26455;
	wire [4-1:0] node26456;
	wire [4-1:0] node26459;
	wire [4-1:0] node26462;
	wire [4-1:0] node26463;
	wire [4-1:0] node26464;
	wire [4-1:0] node26465;
	wire [4-1:0] node26469;
	wire [4-1:0] node26470;
	wire [4-1:0] node26474;
	wire [4-1:0] node26475;
	wire [4-1:0] node26476;
	wire [4-1:0] node26480;
	wire [4-1:0] node26481;
	wire [4-1:0] node26485;
	wire [4-1:0] node26486;
	wire [4-1:0] node26487;
	wire [4-1:0] node26488;
	wire [4-1:0] node26489;
	wire [4-1:0] node26490;
	wire [4-1:0] node26492;
	wire [4-1:0] node26495;
	wire [4-1:0] node26497;
	wire [4-1:0] node26500;
	wire [4-1:0] node26501;
	wire [4-1:0] node26503;
	wire [4-1:0] node26506;
	wire [4-1:0] node26508;
	wire [4-1:0] node26511;
	wire [4-1:0] node26512;
	wire [4-1:0] node26513;
	wire [4-1:0] node26514;
	wire [4-1:0] node26518;
	wire [4-1:0] node26519;
	wire [4-1:0] node26523;
	wire [4-1:0] node26524;
	wire [4-1:0] node26525;
	wire [4-1:0] node26528;
	wire [4-1:0] node26532;
	wire [4-1:0] node26533;
	wire [4-1:0] node26534;
	wire [4-1:0] node26536;
	wire [4-1:0] node26537;
	wire [4-1:0] node26538;
	wire [4-1:0] node26543;
	wire [4-1:0] node26544;
	wire [4-1:0] node26545;
	wire [4-1:0] node26548;
	wire [4-1:0] node26551;
	wire [4-1:0] node26552;
	wire [4-1:0] node26555;
	wire [4-1:0] node26558;
	wire [4-1:0] node26559;
	wire [4-1:0] node26562;
	wire [4-1:0] node26565;
	wire [4-1:0] node26566;
	wire [4-1:0] node26567;
	wire [4-1:0] node26568;
	wire [4-1:0] node26569;
	wire [4-1:0] node26570;
	wire [4-1:0] node26572;
	wire [4-1:0] node26575;
	wire [4-1:0] node26576;
	wire [4-1:0] node26579;
	wire [4-1:0] node26582;
	wire [4-1:0] node26583;
	wire [4-1:0] node26587;
	wire [4-1:0] node26588;
	wire [4-1:0] node26589;
	wire [4-1:0] node26590;
	wire [4-1:0] node26594;
	wire [4-1:0] node26595;
	wire [4-1:0] node26598;
	wire [4-1:0] node26601;
	wire [4-1:0] node26602;
	wire [4-1:0] node26605;
	wire [4-1:0] node26608;
	wire [4-1:0] node26609;
	wire [4-1:0] node26610;
	wire [4-1:0] node26611;
	wire [4-1:0] node26615;
	wire [4-1:0] node26616;
	wire [4-1:0] node26620;
	wire [4-1:0] node26621;
	wire [4-1:0] node26622;
	wire [4-1:0] node26626;
	wire [4-1:0] node26629;
	wire [4-1:0] node26630;
	wire [4-1:0] node26631;
	wire [4-1:0] node26632;
	wire [4-1:0] node26637;
	wire [4-1:0] node26638;
	wire [4-1:0] node26639;
	wire [4-1:0] node26643;
	wire [4-1:0] node26644;
	wire [4-1:0] node26648;
	wire [4-1:0] node26649;
	wire [4-1:0] node26650;
	wire [4-1:0] node26651;
	wire [4-1:0] node26652;
	wire [4-1:0] node26653;
	wire [4-1:0] node26654;
	wire [4-1:0] node26655;
	wire [4-1:0] node26656;
	wire [4-1:0] node26657;
	wire [4-1:0] node26658;
	wire [4-1:0] node26663;
	wire [4-1:0] node26664;
	wire [4-1:0] node26667;
	wire [4-1:0] node26670;
	wire [4-1:0] node26672;
	wire [4-1:0] node26673;
	wire [4-1:0] node26675;
	wire [4-1:0] node26678;
	wire [4-1:0] node26679;
	wire [4-1:0] node26683;
	wire [4-1:0] node26684;
	wire [4-1:0] node26685;
	wire [4-1:0] node26686;
	wire [4-1:0] node26689;
	wire [4-1:0] node26693;
	wire [4-1:0] node26694;
	wire [4-1:0] node26695;
	wire [4-1:0] node26698;
	wire [4-1:0] node26700;
	wire [4-1:0] node26703;
	wire [4-1:0] node26704;
	wire [4-1:0] node26706;
	wire [4-1:0] node26709;
	wire [4-1:0] node26712;
	wire [4-1:0] node26713;
	wire [4-1:0] node26714;
	wire [4-1:0] node26715;
	wire [4-1:0] node26716;
	wire [4-1:0] node26717;
	wire [4-1:0] node26721;
	wire [4-1:0] node26722;
	wire [4-1:0] node26725;
	wire [4-1:0] node26728;
	wire [4-1:0] node26729;
	wire [4-1:0] node26731;
	wire [4-1:0] node26735;
	wire [4-1:0] node26736;
	wire [4-1:0] node26738;
	wire [4-1:0] node26740;
	wire [4-1:0] node26743;
	wire [4-1:0] node26744;
	wire [4-1:0] node26746;
	wire [4-1:0] node26749;
	wire [4-1:0] node26752;
	wire [4-1:0] node26753;
	wire [4-1:0] node26754;
	wire [4-1:0] node26755;
	wire [4-1:0] node26758;
	wire [4-1:0] node26762;
	wire [4-1:0] node26763;
	wire [4-1:0] node26764;
	wire [4-1:0] node26766;
	wire [4-1:0] node26769;
	wire [4-1:0] node26770;
	wire [4-1:0] node26773;
	wire [4-1:0] node26776;
	wire [4-1:0] node26778;
	wire [4-1:0] node26779;
	wire [4-1:0] node26782;
	wire [4-1:0] node26785;
	wire [4-1:0] node26786;
	wire [4-1:0] node26787;
	wire [4-1:0] node26788;
	wire [4-1:0] node26789;
	wire [4-1:0] node26792;
	wire [4-1:0] node26794;
	wire [4-1:0] node26797;
	wire [4-1:0] node26798;
	wire [4-1:0] node26800;
	wire [4-1:0] node26803;
	wire [4-1:0] node26805;
	wire [4-1:0] node26808;
	wire [4-1:0] node26809;
	wire [4-1:0] node26810;
	wire [4-1:0] node26813;
	wire [4-1:0] node26814;
	wire [4-1:0] node26818;
	wire [4-1:0] node26819;
	wire [4-1:0] node26820;
	wire [4-1:0] node26823;
	wire [4-1:0] node26824;
	wire [4-1:0] node26828;
	wire [4-1:0] node26829;
	wire [4-1:0] node26830;
	wire [4-1:0] node26834;
	wire [4-1:0] node26835;
	wire [4-1:0] node26839;
	wire [4-1:0] node26840;
	wire [4-1:0] node26841;
	wire [4-1:0] node26842;
	wire [4-1:0] node26843;
	wire [4-1:0] node26846;
	wire [4-1:0] node26849;
	wire [4-1:0] node26850;
	wire [4-1:0] node26852;
	wire [4-1:0] node26855;
	wire [4-1:0] node26857;
	wire [4-1:0] node26860;
	wire [4-1:0] node26861;
	wire [4-1:0] node26862;
	wire [4-1:0] node26865;
	wire [4-1:0] node26868;
	wire [4-1:0] node26869;
	wire [4-1:0] node26872;
	wire [4-1:0] node26875;
	wire [4-1:0] node26876;
	wire [4-1:0] node26878;
	wire [4-1:0] node26879;
	wire [4-1:0] node26880;
	wire [4-1:0] node26885;
	wire [4-1:0] node26886;
	wire [4-1:0] node26887;
	wire [4-1:0] node26888;
	wire [4-1:0] node26891;
	wire [4-1:0] node26894;
	wire [4-1:0] node26895;
	wire [4-1:0] node26898;
	wire [4-1:0] node26901;
	wire [4-1:0] node26903;
	wire [4-1:0] node26904;
	wire [4-1:0] node26908;
	wire [4-1:0] node26909;
	wire [4-1:0] node26910;
	wire [4-1:0] node26911;
	wire [4-1:0] node26912;
	wire [4-1:0] node26913;
	wire [4-1:0] node26914;
	wire [4-1:0] node26917;
	wire [4-1:0] node26920;
	wire [4-1:0] node26921;
	wire [4-1:0] node26923;
	wire [4-1:0] node26926;
	wire [4-1:0] node26928;
	wire [4-1:0] node26931;
	wire [4-1:0] node26932;
	wire [4-1:0] node26933;
	wire [4-1:0] node26936;
	wire [4-1:0] node26939;
	wire [4-1:0] node26940;
	wire [4-1:0] node26941;
	wire [4-1:0] node26944;
	wire [4-1:0] node26947;
	wire [4-1:0] node26949;
	wire [4-1:0] node26952;
	wire [4-1:0] node26953;
	wire [4-1:0] node26954;
	wire [4-1:0] node26956;
	wire [4-1:0] node26959;
	wire [4-1:0] node26961;
	wire [4-1:0] node26964;
	wire [4-1:0] node26965;
	wire [4-1:0] node26967;
	wire [4-1:0] node26970;
	wire [4-1:0] node26972;
	wire [4-1:0] node26975;
	wire [4-1:0] node26976;
	wire [4-1:0] node26977;
	wire [4-1:0] node26978;
	wire [4-1:0] node26979;
	wire [4-1:0] node26982;
	wire [4-1:0] node26985;
	wire [4-1:0] node26987;
	wire [4-1:0] node26990;
	wire [4-1:0] node26991;
	wire [4-1:0] node26992;
	wire [4-1:0] node26995;
	wire [4-1:0] node26998;
	wire [4-1:0] node26999;
	wire [4-1:0] node27002;
	wire [4-1:0] node27005;
	wire [4-1:0] node27006;
	wire [4-1:0] node27007;
	wire [4-1:0] node27008;
	wire [4-1:0] node27012;
	wire [4-1:0] node27013;
	wire [4-1:0] node27017;
	wire [4-1:0] node27018;
	wire [4-1:0] node27019;
	wire [4-1:0] node27023;
	wire [4-1:0] node27026;
	wire [4-1:0] node27027;
	wire [4-1:0] node27028;
	wire [4-1:0] node27029;
	wire [4-1:0] node27030;
	wire [4-1:0] node27031;
	wire [4-1:0] node27034;
	wire [4-1:0] node27036;
	wire [4-1:0] node27039;
	wire [4-1:0] node27041;
	wire [4-1:0] node27042;
	wire [4-1:0] node27045;
	wire [4-1:0] node27048;
	wire [4-1:0] node27049;
	wire [4-1:0] node27051;
	wire [4-1:0] node27052;
	wire [4-1:0] node27055;
	wire [4-1:0] node27058;
	wire [4-1:0] node27059;
	wire [4-1:0] node27063;
	wire [4-1:0] node27064;
	wire [4-1:0] node27065;
	wire [4-1:0] node27066;
	wire [4-1:0] node27067;
	wire [4-1:0] node27070;
	wire [4-1:0] node27073;
	wire [4-1:0] node27075;
	wire [4-1:0] node27079;
	wire [4-1:0] node27080;
	wire [4-1:0] node27083;
	wire [4-1:0] node27086;
	wire [4-1:0] node27087;
	wire [4-1:0] node27088;
	wire [4-1:0] node27089;
	wire [4-1:0] node27090;
	wire [4-1:0] node27091;
	wire [4-1:0] node27095;
	wire [4-1:0] node27096;
	wire [4-1:0] node27100;
	wire [4-1:0] node27101;
	wire [4-1:0] node27104;
	wire [4-1:0] node27107;
	wire [4-1:0] node27108;
	wire [4-1:0] node27109;
	wire [4-1:0] node27110;
	wire [4-1:0] node27113;
	wire [4-1:0] node27116;
	wire [4-1:0] node27117;
	wire [4-1:0] node27120;
	wire [4-1:0] node27123;
	wire [4-1:0] node27124;
	wire [4-1:0] node27128;
	wire [4-1:0] node27129;
	wire [4-1:0] node27130;
	wire [4-1:0] node27131;
	wire [4-1:0] node27132;
	wire [4-1:0] node27135;
	wire [4-1:0] node27138;
	wire [4-1:0] node27140;
	wire [4-1:0] node27143;
	wire [4-1:0] node27144;
	wire [4-1:0] node27147;
	wire [4-1:0] node27150;
	wire [4-1:0] node27151;
	wire [4-1:0] node27154;
	wire [4-1:0] node27157;
	wire [4-1:0] node27158;
	wire [4-1:0] node27159;
	wire [4-1:0] node27160;
	wire [4-1:0] node27161;
	wire [4-1:0] node27162;
	wire [4-1:0] node27163;
	wire [4-1:0] node27164;
	wire [4-1:0] node27165;
	wire [4-1:0] node27168;
	wire [4-1:0] node27171;
	wire [4-1:0] node27172;
	wire [4-1:0] node27176;
	wire [4-1:0] node27177;
	wire [4-1:0] node27178;
	wire [4-1:0] node27183;
	wire [4-1:0] node27184;
	wire [4-1:0] node27186;
	wire [4-1:0] node27188;
	wire [4-1:0] node27191;
	wire [4-1:0] node27194;
	wire [4-1:0] node27195;
	wire [4-1:0] node27196;
	wire [4-1:0] node27197;
	wire [4-1:0] node27200;
	wire [4-1:0] node27203;
	wire [4-1:0] node27204;
	wire [4-1:0] node27207;
	wire [4-1:0] node27210;
	wire [4-1:0] node27211;
	wire [4-1:0] node27212;
	wire [4-1:0] node27213;
	wire [4-1:0] node27217;
	wire [4-1:0] node27220;
	wire [4-1:0] node27221;
	wire [4-1:0] node27225;
	wire [4-1:0] node27226;
	wire [4-1:0] node27227;
	wire [4-1:0] node27228;
	wire [4-1:0] node27229;
	wire [4-1:0] node27233;
	wire [4-1:0] node27234;
	wire [4-1:0] node27235;
	wire [4-1:0] node27239;
	wire [4-1:0] node27240;
	wire [4-1:0] node27243;
	wire [4-1:0] node27246;
	wire [4-1:0] node27247;
	wire [4-1:0] node27248;
	wire [4-1:0] node27251;
	wire [4-1:0] node27252;
	wire [4-1:0] node27256;
	wire [4-1:0] node27257;
	wire [4-1:0] node27260;
	wire [4-1:0] node27263;
	wire [4-1:0] node27264;
	wire [4-1:0] node27265;
	wire [4-1:0] node27266;
	wire [4-1:0] node27267;
	wire [4-1:0] node27271;
	wire [4-1:0] node27272;
	wire [4-1:0] node27276;
	wire [4-1:0] node27277;
	wire [4-1:0] node27281;
	wire [4-1:0] node27282;
	wire [4-1:0] node27285;
	wire [4-1:0] node27287;
	wire [4-1:0] node27290;
	wire [4-1:0] node27291;
	wire [4-1:0] node27292;
	wire [4-1:0] node27293;
	wire [4-1:0] node27294;
	wire [4-1:0] node27295;
	wire [4-1:0] node27298;
	wire [4-1:0] node27301;
	wire [4-1:0] node27302;
	wire [4-1:0] node27303;
	wire [4-1:0] node27306;
	wire [4-1:0] node27309;
	wire [4-1:0] node27311;
	wire [4-1:0] node27314;
	wire [4-1:0] node27315;
	wire [4-1:0] node27316;
	wire [4-1:0] node27318;
	wire [4-1:0] node27321;
	wire [4-1:0] node27322;
	wire [4-1:0] node27326;
	wire [4-1:0] node27327;
	wire [4-1:0] node27331;
	wire [4-1:0] node27332;
	wire [4-1:0] node27333;
	wire [4-1:0] node27335;
	wire [4-1:0] node27336;
	wire [4-1:0] node27339;
	wire [4-1:0] node27342;
	wire [4-1:0] node27343;
	wire [4-1:0] node27344;
	wire [4-1:0] node27347;
	wire [4-1:0] node27350;
	wire [4-1:0] node27351;
	wire [4-1:0] node27354;
	wire [4-1:0] node27357;
	wire [4-1:0] node27358;
	wire [4-1:0] node27359;
	wire [4-1:0] node27362;
	wire [4-1:0] node27365;
	wire [4-1:0] node27366;
	wire [4-1:0] node27370;
	wire [4-1:0] node27371;
	wire [4-1:0] node27372;
	wire [4-1:0] node27373;
	wire [4-1:0] node27376;
	wire [4-1:0] node27377;
	wire [4-1:0] node27380;
	wire [4-1:0] node27381;
	wire [4-1:0] node27385;
	wire [4-1:0] node27386;
	wire [4-1:0] node27387;
	wire [4-1:0] node27389;
	wire [4-1:0] node27392;
	wire [4-1:0] node27393;
	wire [4-1:0] node27396;
	wire [4-1:0] node27399;
	wire [4-1:0] node27400;
	wire [4-1:0] node27403;
	wire [4-1:0] node27406;
	wire [4-1:0] node27407;
	wire [4-1:0] node27408;
	wire [4-1:0] node27409;
	wire [4-1:0] node27413;
	wire [4-1:0] node27414;
	wire [4-1:0] node27418;
	wire [4-1:0] node27419;
	wire [4-1:0] node27422;
	wire [4-1:0] node27423;
	wire [4-1:0] node27427;
	wire [4-1:0] node27428;
	wire [4-1:0] node27429;
	wire [4-1:0] node27430;
	wire [4-1:0] node27431;
	wire [4-1:0] node27432;
	wire [4-1:0] node27434;
	wire [4-1:0] node27435;
	wire [4-1:0] node27438;
	wire [4-1:0] node27441;
	wire [4-1:0] node27442;
	wire [4-1:0] node27443;
	wire [4-1:0] node27446;
	wire [4-1:0] node27449;
	wire [4-1:0] node27450;
	wire [4-1:0] node27453;
	wire [4-1:0] node27456;
	wire [4-1:0] node27457;
	wire [4-1:0] node27458;
	wire [4-1:0] node27459;
	wire [4-1:0] node27462;
	wire [4-1:0] node27466;
	wire [4-1:0] node27467;
	wire [4-1:0] node27469;
	wire [4-1:0] node27472;
	wire [4-1:0] node27473;
	wire [4-1:0] node27476;
	wire [4-1:0] node27479;
	wire [4-1:0] node27480;
	wire [4-1:0] node27481;
	wire [4-1:0] node27482;
	wire [4-1:0] node27483;
	wire [4-1:0] node27486;
	wire [4-1:0] node27489;
	wire [4-1:0] node27490;
	wire [4-1:0] node27494;
	wire [4-1:0] node27495;
	wire [4-1:0] node27498;
	wire [4-1:0] node27500;
	wire [4-1:0] node27503;
	wire [4-1:0] node27504;
	wire [4-1:0] node27505;
	wire [4-1:0] node27509;
	wire [4-1:0] node27510;
	wire [4-1:0] node27512;
	wire [4-1:0] node27516;
	wire [4-1:0] node27517;
	wire [4-1:0] node27518;
	wire [4-1:0] node27519;
	wire [4-1:0] node27520;
	wire [4-1:0] node27523;
	wire [4-1:0] node27526;
	wire [4-1:0] node27527;
	wire [4-1:0] node27530;
	wire [4-1:0] node27533;
	wire [4-1:0] node27534;
	wire [4-1:0] node27536;
	wire [4-1:0] node27537;
	wire [4-1:0] node27541;
	wire [4-1:0] node27542;
	wire [4-1:0] node27545;
	wire [4-1:0] node27548;
	wire [4-1:0] node27549;
	wire [4-1:0] node27550;
	wire [4-1:0] node27551;
	wire [4-1:0] node27554;
	wire [4-1:0] node27557;
	wire [4-1:0] node27559;
	wire [4-1:0] node27562;
	wire [4-1:0] node27563;
	wire [4-1:0] node27564;
	wire [4-1:0] node27567;
	wire [4-1:0] node27570;
	wire [4-1:0] node27571;
	wire [4-1:0] node27573;
	wire [4-1:0] node27576;
	wire [4-1:0] node27578;
	wire [4-1:0] node27581;
	wire [4-1:0] node27582;
	wire [4-1:0] node27583;
	wire [4-1:0] node27584;
	wire [4-1:0] node27585;
	wire [4-1:0] node27586;
	wire [4-1:0] node27587;
	wire [4-1:0] node27590;
	wire [4-1:0] node27593;
	wire [4-1:0] node27594;
	wire [4-1:0] node27597;
	wire [4-1:0] node27600;
	wire [4-1:0] node27601;
	wire [4-1:0] node27603;
	wire [4-1:0] node27606;
	wire [4-1:0] node27607;
	wire [4-1:0] node27610;
	wire [4-1:0] node27613;
	wire [4-1:0] node27614;
	wire [4-1:0] node27615;
	wire [4-1:0] node27617;
	wire [4-1:0] node27620;
	wire [4-1:0] node27622;
	wire [4-1:0] node27625;
	wire [4-1:0] node27626;
	wire [4-1:0] node27627;
	wire [4-1:0] node27632;
	wire [4-1:0] node27633;
	wire [4-1:0] node27634;
	wire [4-1:0] node27635;
	wire [4-1:0] node27636;
	wire [4-1:0] node27639;
	wire [4-1:0] node27642;
	wire [4-1:0] node27643;
	wire [4-1:0] node27646;
	wire [4-1:0] node27649;
	wire [4-1:0] node27650;
	wire [4-1:0] node27653;
	wire [4-1:0] node27656;
	wire [4-1:0] node27657;
	wire [4-1:0] node27658;
	wire [4-1:0] node27660;
	wire [4-1:0] node27663;
	wire [4-1:0] node27666;
	wire [4-1:0] node27667;
	wire [4-1:0] node27668;
	wire [4-1:0] node27672;
	wire [4-1:0] node27675;
	wire [4-1:0] node27676;
	wire [4-1:0] node27677;
	wire [4-1:0] node27678;
	wire [4-1:0] node27679;
	wire [4-1:0] node27680;
	wire [4-1:0] node27683;
	wire [4-1:0] node27687;
	wire [4-1:0] node27688;
	wire [4-1:0] node27691;
	wire [4-1:0] node27694;
	wire [4-1:0] node27695;
	wire [4-1:0] node27696;
	wire [4-1:0] node27699;
	wire [4-1:0] node27702;
	wire [4-1:0] node27703;
	wire [4-1:0] node27704;
	wire [4-1:0] node27708;
	wire [4-1:0] node27710;
	wire [4-1:0] node27713;
	wire [4-1:0] node27714;
	wire [4-1:0] node27715;
	wire [4-1:0] node27716;
	wire [4-1:0] node27719;
	wire [4-1:0] node27722;
	wire [4-1:0] node27723;
	wire [4-1:0] node27725;
	wire [4-1:0] node27728;
	wire [4-1:0] node27729;
	wire [4-1:0] node27733;
	wire [4-1:0] node27734;
	wire [4-1:0] node27736;
	wire [4-1:0] node27739;
	wire [4-1:0] node27740;
	wire [4-1:0] node27742;
	wire [4-1:0] node27745;
	wire [4-1:0] node27747;
	wire [4-1:0] node27750;
	wire [4-1:0] node27751;
	wire [4-1:0] node27752;
	wire [4-1:0] node27753;
	wire [4-1:0] node27754;
	wire [4-1:0] node27755;
	wire [4-1:0] node27756;
	wire [4-1:0] node27757;
	wire [4-1:0] node27758;
	wire [4-1:0] node27761;
	wire [4-1:0] node27764;
	wire [4-1:0] node27765;
	wire [4-1:0] node27768;
	wire [4-1:0] node27771;
	wire [4-1:0] node27773;
	wire [4-1:0] node27774;
	wire [4-1:0] node27775;
	wire [4-1:0] node27778;
	wire [4-1:0] node27781;
	wire [4-1:0] node27782;
	wire [4-1:0] node27786;
	wire [4-1:0] node27787;
	wire [4-1:0] node27788;
	wire [4-1:0] node27791;
	wire [4-1:0] node27792;
	wire [4-1:0] node27793;
	wire [4-1:0] node27796;
	wire [4-1:0] node27800;
	wire [4-1:0] node27801;
	wire [4-1:0] node27802;
	wire [4-1:0] node27803;
	wire [4-1:0] node27807;
	wire [4-1:0] node27808;
	wire [4-1:0] node27811;
	wire [4-1:0] node27814;
	wire [4-1:0] node27816;
	wire [4-1:0] node27818;
	wire [4-1:0] node27821;
	wire [4-1:0] node27822;
	wire [4-1:0] node27823;
	wire [4-1:0] node27824;
	wire [4-1:0] node27825;
	wire [4-1:0] node27826;
	wire [4-1:0] node27829;
	wire [4-1:0] node27832;
	wire [4-1:0] node27833;
	wire [4-1:0] node27836;
	wire [4-1:0] node27839;
	wire [4-1:0] node27840;
	wire [4-1:0] node27841;
	wire [4-1:0] node27845;
	wire [4-1:0] node27846;
	wire [4-1:0] node27850;
	wire [4-1:0] node27851;
	wire [4-1:0] node27852;
	wire [4-1:0] node27855;
	wire [4-1:0] node27858;
	wire [4-1:0] node27859;
	wire [4-1:0] node27863;
	wire [4-1:0] node27864;
	wire [4-1:0] node27865;
	wire [4-1:0] node27866;
	wire [4-1:0] node27867;
	wire [4-1:0] node27870;
	wire [4-1:0] node27873;
	wire [4-1:0] node27874;
	wire [4-1:0] node27878;
	wire [4-1:0] node27881;
	wire [4-1:0] node27882;
	wire [4-1:0] node27883;
	wire [4-1:0] node27884;
	wire [4-1:0] node27887;
	wire [4-1:0] node27890;
	wire [4-1:0] node27892;
	wire [4-1:0] node27895;
	wire [4-1:0] node27897;
	wire [4-1:0] node27898;
	wire [4-1:0] node27901;
	wire [4-1:0] node27904;
	wire [4-1:0] node27905;
	wire [4-1:0] node27906;
	wire [4-1:0] node27907;
	wire [4-1:0] node27908;
	wire [4-1:0] node27909;
	wire [4-1:0] node27910;
	wire [4-1:0] node27915;
	wire [4-1:0] node27916;
	wire [4-1:0] node27917;
	wire [4-1:0] node27920;
	wire [4-1:0] node27923;
	wire [4-1:0] node27925;
	wire [4-1:0] node27928;
	wire [4-1:0] node27929;
	wire [4-1:0] node27930;
	wire [4-1:0] node27931;
	wire [4-1:0] node27934;
	wire [4-1:0] node27938;
	wire [4-1:0] node27939;
	wire [4-1:0] node27942;
	wire [4-1:0] node27945;
	wire [4-1:0] node27946;
	wire [4-1:0] node27947;
	wire [4-1:0] node27948;
	wire [4-1:0] node27949;
	wire [4-1:0] node27953;
	wire [4-1:0] node27956;
	wire [4-1:0] node27957;
	wire [4-1:0] node27960;
	wire [4-1:0] node27963;
	wire [4-1:0] node27964;
	wire [4-1:0] node27965;
	wire [4-1:0] node27966;
	wire [4-1:0] node27970;
	wire [4-1:0] node27973;
	wire [4-1:0] node27974;
	wire [4-1:0] node27976;
	wire [4-1:0] node27979;
	wire [4-1:0] node27980;
	wire [4-1:0] node27983;
	wire [4-1:0] node27986;
	wire [4-1:0] node27987;
	wire [4-1:0] node27988;
	wire [4-1:0] node27989;
	wire [4-1:0] node27990;
	wire [4-1:0] node27994;
	wire [4-1:0] node27997;
	wire [4-1:0] node27998;
	wire [4-1:0] node27999;
	wire [4-1:0] node28003;
	wire [4-1:0] node28006;
	wire [4-1:0] node28007;
	wire [4-1:0] node28008;
	wire [4-1:0] node28010;
	wire [4-1:0] node28013;
	wire [4-1:0] node28014;
	wire [4-1:0] node28015;
	wire [4-1:0] node28018;
	wire [4-1:0] node28021;
	wire [4-1:0] node28022;
	wire [4-1:0] node28025;
	wire [4-1:0] node28028;
	wire [4-1:0] node28029;
	wire [4-1:0] node28030;
	wire [4-1:0] node28034;
	wire [4-1:0] node28037;
	wire [4-1:0] node28038;
	wire [4-1:0] node28039;
	wire [4-1:0] node28040;
	wire [4-1:0] node28041;
	wire [4-1:0] node28042;
	wire [4-1:0] node28043;
	wire [4-1:0] node28046;
	wire [4-1:0] node28050;
	wire [4-1:0] node28051;
	wire [4-1:0] node28052;
	wire [4-1:0] node28054;
	wire [4-1:0] node28058;
	wire [4-1:0] node28059;
	wire [4-1:0] node28062;
	wire [4-1:0] node28065;
	wire [4-1:0] node28066;
	wire [4-1:0] node28067;
	wire [4-1:0] node28068;
	wire [4-1:0] node28069;
	wire [4-1:0] node28072;
	wire [4-1:0] node28076;
	wire [4-1:0] node28077;
	wire [4-1:0] node28078;
	wire [4-1:0] node28081;
	wire [4-1:0] node28085;
	wire [4-1:0] node28086;
	wire [4-1:0] node28087;
	wire [4-1:0] node28090;
	wire [4-1:0] node28093;
	wire [4-1:0] node28095;
	wire [4-1:0] node28098;
	wire [4-1:0] node28099;
	wire [4-1:0] node28100;
	wire [4-1:0] node28101;
	wire [4-1:0] node28102;
	wire [4-1:0] node28105;
	wire [4-1:0] node28108;
	wire [4-1:0] node28109;
	wire [4-1:0] node28110;
	wire [4-1:0] node28113;
	wire [4-1:0] node28116;
	wire [4-1:0] node28118;
	wire [4-1:0] node28121;
	wire [4-1:0] node28122;
	wire [4-1:0] node28123;
	wire [4-1:0] node28126;
	wire [4-1:0] node28129;
	wire [4-1:0] node28130;
	wire [4-1:0] node28133;
	wire [4-1:0] node28136;
	wire [4-1:0] node28137;
	wire [4-1:0] node28138;
	wire [4-1:0] node28139;
	wire [4-1:0] node28140;
	wire [4-1:0] node28143;
	wire [4-1:0] node28146;
	wire [4-1:0] node28147;
	wire [4-1:0] node28151;
	wire [4-1:0] node28152;
	wire [4-1:0] node28153;
	wire [4-1:0] node28156;
	wire [4-1:0] node28159;
	wire [4-1:0] node28160;
	wire [4-1:0] node28164;
	wire [4-1:0] node28165;
	wire [4-1:0] node28166;
	wire [4-1:0] node28169;
	wire [4-1:0] node28172;
	wire [4-1:0] node28173;
	wire [4-1:0] node28176;
	wire [4-1:0] node28179;
	wire [4-1:0] node28180;
	wire [4-1:0] node28181;
	wire [4-1:0] node28182;
	wire [4-1:0] node28183;
	wire [4-1:0] node28184;
	wire [4-1:0] node28185;
	wire [4-1:0] node28188;
	wire [4-1:0] node28191;
	wire [4-1:0] node28192;
	wire [4-1:0] node28195;
	wire [4-1:0] node28198;
	wire [4-1:0] node28199;
	wire [4-1:0] node28201;
	wire [4-1:0] node28204;
	wire [4-1:0] node28205;
	wire [4-1:0] node28208;
	wire [4-1:0] node28211;
	wire [4-1:0] node28212;
	wire [4-1:0] node28213;
	wire [4-1:0] node28214;
	wire [4-1:0] node28217;
	wire [4-1:0] node28220;
	wire [4-1:0] node28221;
	wire [4-1:0] node28224;
	wire [4-1:0] node28227;
	wire [4-1:0] node28228;
	wire [4-1:0] node28229;
	wire [4-1:0] node28232;
	wire [4-1:0] node28235;
	wire [4-1:0] node28236;
	wire [4-1:0] node28239;
	wire [4-1:0] node28242;
	wire [4-1:0] node28243;
	wire [4-1:0] node28244;
	wire [4-1:0] node28245;
	wire [4-1:0] node28248;
	wire [4-1:0] node28251;
	wire [4-1:0] node28252;
	wire [4-1:0] node28253;
	wire [4-1:0] node28257;
	wire [4-1:0] node28260;
	wire [4-1:0] node28261;
	wire [4-1:0] node28262;
	wire [4-1:0] node28263;
	wire [4-1:0] node28267;
	wire [4-1:0] node28268;
	wire [4-1:0] node28271;
	wire [4-1:0] node28274;
	wire [4-1:0] node28275;
	wire [4-1:0] node28276;
	wire [4-1:0] node28280;
	wire [4-1:0] node28283;
	wire [4-1:0] node28284;
	wire [4-1:0] node28285;
	wire [4-1:0] node28286;
	wire [4-1:0] node28287;
	wire [4-1:0] node28291;
	wire [4-1:0] node28292;
	wire [4-1:0] node28294;
	wire [4-1:0] node28297;
	wire [4-1:0] node28298;
	wire [4-1:0] node28301;
	wire [4-1:0] node28304;
	wire [4-1:0] node28305;
	wire [4-1:0] node28306;
	wire [4-1:0] node28307;
	wire [4-1:0] node28310;
	wire [4-1:0] node28313;
	wire [4-1:0] node28314;
	wire [4-1:0] node28317;
	wire [4-1:0] node28320;
	wire [4-1:0] node28321;
	wire [4-1:0] node28324;
	wire [4-1:0] node28327;
	wire [4-1:0] node28328;
	wire [4-1:0] node28329;
	wire [4-1:0] node28330;
	wire [4-1:0] node28332;
	wire [4-1:0] node28336;
	wire [4-1:0] node28337;
	wire [4-1:0] node28338;
	wire [4-1:0] node28342;
	wire [4-1:0] node28345;
	wire [4-1:0] node28346;
	wire [4-1:0] node28347;
	wire [4-1:0] node28348;
	wire [4-1:0] node28352;
	wire [4-1:0] node28353;
	wire [4-1:0] node28357;
	wire [4-1:0] node28358;
	wire [4-1:0] node28361;
	wire [4-1:0] node28364;
	wire [4-1:0] node28365;
	wire [4-1:0] node28366;
	wire [4-1:0] node28367;
	wire [4-1:0] node28368;
	wire [4-1:0] node28369;
	wire [4-1:0] node28370;
	wire [4-1:0] node28371;
	wire [4-1:0] node28374;
	wire [4-1:0] node28376;
	wire [4-1:0] node28379;
	wire [4-1:0] node28380;
	wire [4-1:0] node28381;
	wire [4-1:0] node28384;
	wire [4-1:0] node28387;
	wire [4-1:0] node28388;
	wire [4-1:0] node28391;
	wire [4-1:0] node28394;
	wire [4-1:0] node28395;
	wire [4-1:0] node28396;
	wire [4-1:0] node28397;
	wire [4-1:0] node28400;
	wire [4-1:0] node28403;
	wire [4-1:0] node28404;
	wire [4-1:0] node28407;
	wire [4-1:0] node28410;
	wire [4-1:0] node28411;
	wire [4-1:0] node28415;
	wire [4-1:0] node28416;
	wire [4-1:0] node28417;
	wire [4-1:0] node28418;
	wire [4-1:0] node28422;
	wire [4-1:0] node28423;
	wire [4-1:0] node28427;
	wire [4-1:0] node28428;
	wire [4-1:0] node28429;
	wire [4-1:0] node28433;
	wire [4-1:0] node28436;
	wire [4-1:0] node28437;
	wire [4-1:0] node28438;
	wire [4-1:0] node28439;
	wire [4-1:0] node28440;
	wire [4-1:0] node28444;
	wire [4-1:0] node28447;
	wire [4-1:0] node28448;
	wire [4-1:0] node28449;
	wire [4-1:0] node28453;
	wire [4-1:0] node28454;
	wire [4-1:0] node28458;
	wire [4-1:0] node28459;
	wire [4-1:0] node28460;
	wire [4-1:0] node28461;
	wire [4-1:0] node28464;
	wire [4-1:0] node28467;
	wire [4-1:0] node28468;
	wire [4-1:0] node28471;
	wire [4-1:0] node28474;
	wire [4-1:0] node28475;
	wire [4-1:0] node28479;
	wire [4-1:0] node28480;
	wire [4-1:0] node28481;
	wire [4-1:0] node28482;
	wire [4-1:0] node28483;
	wire [4-1:0] node28484;
	wire [4-1:0] node28485;
	wire [4-1:0] node28488;
	wire [4-1:0] node28491;
	wire [4-1:0] node28492;
	wire [4-1:0] node28496;
	wire [4-1:0] node28497;
	wire [4-1:0] node28500;
	wire [4-1:0] node28503;
	wire [4-1:0] node28504;
	wire [4-1:0] node28505;
	wire [4-1:0] node28507;
	wire [4-1:0] node28510;
	wire [4-1:0] node28511;
	wire [4-1:0] node28515;
	wire [4-1:0] node28517;
	wire [4-1:0] node28520;
	wire [4-1:0] node28521;
	wire [4-1:0] node28522;
	wire [4-1:0] node28523;
	wire [4-1:0] node28527;
	wire [4-1:0] node28529;
	wire [4-1:0] node28530;
	wire [4-1:0] node28534;
	wire [4-1:0] node28535;
	wire [4-1:0] node28536;
	wire [4-1:0] node28540;
	wire [4-1:0] node28541;
	wire [4-1:0] node28545;
	wire [4-1:0] node28546;
	wire [4-1:0] node28547;
	wire [4-1:0] node28548;
	wire [4-1:0] node28549;
	wire [4-1:0] node28553;
	wire [4-1:0] node28554;
	wire [4-1:0] node28558;
	wire [4-1:0] node28560;
	wire [4-1:0] node28563;
	wire [4-1:0] node28564;
	wire [4-1:0] node28565;
	wire [4-1:0] node28566;
	wire [4-1:0] node28570;
	wire [4-1:0] node28571;
	wire [4-1:0] node28575;
	wire [4-1:0] node28576;
	wire [4-1:0] node28577;
	wire [4-1:0] node28581;
	wire [4-1:0] node28582;
	wire [4-1:0] node28586;
	wire [4-1:0] node28587;
	wire [4-1:0] node28588;
	wire [4-1:0] node28589;
	wire [4-1:0] node28590;
	wire [4-1:0] node28591;
	wire [4-1:0] node28593;
	wire [4-1:0] node28594;
	wire [4-1:0] node28597;
	wire [4-1:0] node28600;
	wire [4-1:0] node28601;
	wire [4-1:0] node28602;
	wire [4-1:0] node28605;
	wire [4-1:0] node28608;
	wire [4-1:0] node28609;
	wire [4-1:0] node28612;
	wire [4-1:0] node28615;
	wire [4-1:0] node28616;
	wire [4-1:0] node28617;
	wire [4-1:0] node28618;
	wire [4-1:0] node28623;
	wire [4-1:0] node28624;
	wire [4-1:0] node28625;
	wire [4-1:0] node28629;
	wire [4-1:0] node28630;
	wire [4-1:0] node28634;
	wire [4-1:0] node28635;
	wire [4-1:0] node28636;
	wire [4-1:0] node28637;
	wire [4-1:0] node28641;
	wire [4-1:0] node28644;
	wire [4-1:0] node28645;
	wire [4-1:0] node28646;
	wire [4-1:0] node28650;
	wire [4-1:0] node28651;
	wire [4-1:0] node28655;
	wire [4-1:0] node28656;
	wire [4-1:0] node28657;
	wire [4-1:0] node28658;
	wire [4-1:0] node28659;
	wire [4-1:0] node28663;
	wire [4-1:0] node28664;
	wire [4-1:0] node28668;
	wire [4-1:0] node28669;
	wire [4-1:0] node28670;
	wire [4-1:0] node28674;
	wire [4-1:0] node28675;
	wire [4-1:0] node28679;
	wire [4-1:0] node28680;
	wire [4-1:0] node28681;
	wire [4-1:0] node28682;
	wire [4-1:0] node28686;
	wire [4-1:0] node28687;
	wire [4-1:0] node28691;
	wire [4-1:0] node28692;
	wire [4-1:0] node28693;
	wire [4-1:0] node28697;
	wire [4-1:0] node28698;
	wire [4-1:0] node28702;
	wire [4-1:0] node28703;
	wire [4-1:0] node28704;
	wire [4-1:0] node28705;
	wire [4-1:0] node28706;
	wire [4-1:0] node28707;
	wire [4-1:0] node28711;
	wire [4-1:0] node28712;
	wire [4-1:0] node28716;
	wire [4-1:0] node28717;
	wire [4-1:0] node28720;
	wire [4-1:0] node28721;
	wire [4-1:0] node28725;
	wire [4-1:0] node28726;
	wire [4-1:0] node28727;
	wire [4-1:0] node28728;
	wire [4-1:0] node28732;
	wire [4-1:0] node28733;
	wire [4-1:0] node28737;
	wire [4-1:0] node28738;
	wire [4-1:0] node28739;
	wire [4-1:0] node28743;
	wire [4-1:0] node28744;
	wire [4-1:0] node28748;
	wire [4-1:0] node28749;
	wire [4-1:0] node28750;
	wire [4-1:0] node28751;
	wire [4-1:0] node28752;
	wire [4-1:0] node28756;
	wire [4-1:0] node28757;
	wire [4-1:0] node28761;
	wire [4-1:0] node28762;
	wire [4-1:0] node28763;
	wire [4-1:0] node28767;
	wire [4-1:0] node28770;
	wire [4-1:0] node28771;
	wire [4-1:0] node28772;
	wire [4-1:0] node28773;
	wire [4-1:0] node28774;
	wire [4-1:0] node28777;
	wire [4-1:0] node28780;
	wire [4-1:0] node28782;
	wire [4-1:0] node28785;
	wire [4-1:0] node28786;
	wire [4-1:0] node28788;
	wire [4-1:0] node28791;
	wire [4-1:0] node28792;
	wire [4-1:0] node28795;
	wire [4-1:0] node28798;
	wire [4-1:0] node28799;
	wire [4-1:0] node28800;
	wire [4-1:0] node28803;
	wire [4-1:0] node28806;
	wire [4-1:0] node28808;
	wire [4-1:0] node28811;
	wire [4-1:0] node28812;
	wire [4-1:0] node28813;
	wire [4-1:0] node28814;
	wire [4-1:0] node28815;
	wire [4-1:0] node28816;
	wire [4-1:0] node28817;
	wire [4-1:0] node28818;
	wire [4-1:0] node28819;
	wire [4-1:0] node28820;
	wire [4-1:0] node28821;
	wire [4-1:0] node28822;
	wire [4-1:0] node28825;
	wire [4-1:0] node28828;
	wire [4-1:0] node28829;
	wire [4-1:0] node28832;
	wire [4-1:0] node28835;
	wire [4-1:0] node28836;
	wire [4-1:0] node28837;
	wire [4-1:0] node28841;
	wire [4-1:0] node28843;
	wire [4-1:0] node28846;
	wire [4-1:0] node28847;
	wire [4-1:0] node28849;
	wire [4-1:0] node28852;
	wire [4-1:0] node28853;
	wire [4-1:0] node28856;
	wire [4-1:0] node28857;
	wire [4-1:0] node28860;
	wire [4-1:0] node28863;
	wire [4-1:0] node28864;
	wire [4-1:0] node28865;
	wire [4-1:0] node28866;
	wire [4-1:0] node28867;
	wire [4-1:0] node28870;
	wire [4-1:0] node28873;
	wire [4-1:0] node28874;
	wire [4-1:0] node28877;
	wire [4-1:0] node28880;
	wire [4-1:0] node28881;
	wire [4-1:0] node28882;
	wire [4-1:0] node28885;
	wire [4-1:0] node28888;
	wire [4-1:0] node28889;
	wire [4-1:0] node28893;
	wire [4-1:0] node28894;
	wire [4-1:0] node28895;
	wire [4-1:0] node28896;
	wire [4-1:0] node28900;
	wire [4-1:0] node28901;
	wire [4-1:0] node28904;
	wire [4-1:0] node28907;
	wire [4-1:0] node28908;
	wire [4-1:0] node28909;
	wire [4-1:0] node28912;
	wire [4-1:0] node28916;
	wire [4-1:0] node28917;
	wire [4-1:0] node28918;
	wire [4-1:0] node28919;
	wire [4-1:0] node28921;
	wire [4-1:0] node28922;
	wire [4-1:0] node28925;
	wire [4-1:0] node28928;
	wire [4-1:0] node28929;
	wire [4-1:0] node28930;
	wire [4-1:0] node28933;
	wire [4-1:0] node28936;
	wire [4-1:0] node28939;
	wire [4-1:0] node28940;
	wire [4-1:0] node28941;
	wire [4-1:0] node28942;
	wire [4-1:0] node28946;
	wire [4-1:0] node28949;
	wire [4-1:0] node28950;
	wire [4-1:0] node28953;
	wire [4-1:0] node28954;
	wire [4-1:0] node28957;
	wire [4-1:0] node28960;
	wire [4-1:0] node28961;
	wire [4-1:0] node28962;
	wire [4-1:0] node28963;
	wire [4-1:0] node28964;
	wire [4-1:0] node28968;
	wire [4-1:0] node28970;
	wire [4-1:0] node28973;
	wire [4-1:0] node28975;
	wire [4-1:0] node28976;
	wire [4-1:0] node28980;
	wire [4-1:0] node28982;
	wire [4-1:0] node28983;
	wire [4-1:0] node28984;
	wire [4-1:0] node28987;
	wire [4-1:0] node28991;
	wire [4-1:0] node28992;
	wire [4-1:0] node28993;
	wire [4-1:0] node28994;
	wire [4-1:0] node28995;
	wire [4-1:0] node28996;
	wire [4-1:0] node28999;
	wire [4-1:0] node29002;
	wire [4-1:0] node29003;
	wire [4-1:0] node29005;
	wire [4-1:0] node29008;
	wire [4-1:0] node29010;
	wire [4-1:0] node29013;
	wire [4-1:0] node29014;
	wire [4-1:0] node29016;
	wire [4-1:0] node29018;
	wire [4-1:0] node29021;
	wire [4-1:0] node29023;
	wire [4-1:0] node29024;
	wire [4-1:0] node29028;
	wire [4-1:0] node29029;
	wire [4-1:0] node29031;
	wire [4-1:0] node29033;
	wire [4-1:0] node29036;
	wire [4-1:0] node29037;
	wire [4-1:0] node29038;
	wire [4-1:0] node29041;
	wire [4-1:0] node29042;
	wire [4-1:0] node29045;
	wire [4-1:0] node29048;
	wire [4-1:0] node29049;
	wire [4-1:0] node29051;
	wire [4-1:0] node29054;
	wire [4-1:0] node29057;
	wire [4-1:0] node29058;
	wire [4-1:0] node29059;
	wire [4-1:0] node29060;
	wire [4-1:0] node29061;
	wire [4-1:0] node29064;
	wire [4-1:0] node29067;
	wire [4-1:0] node29068;
	wire [4-1:0] node29069;
	wire [4-1:0] node29074;
	wire [4-1:0] node29075;
	wire [4-1:0] node29076;
	wire [4-1:0] node29077;
	wire [4-1:0] node29080;
	wire [4-1:0] node29083;
	wire [4-1:0] node29084;
	wire [4-1:0] node29087;
	wire [4-1:0] node29090;
	wire [4-1:0] node29091;
	wire [4-1:0] node29092;
	wire [4-1:0] node29095;
	wire [4-1:0] node29098;
	wire [4-1:0] node29099;
	wire [4-1:0] node29103;
	wire [4-1:0] node29104;
	wire [4-1:0] node29105;
	wire [4-1:0] node29106;
	wire [4-1:0] node29108;
	wire [4-1:0] node29111;
	wire [4-1:0] node29114;
	wire [4-1:0] node29115;
	wire [4-1:0] node29119;
	wire [4-1:0] node29120;
	wire [4-1:0] node29122;
	wire [4-1:0] node29123;
	wire [4-1:0] node29126;
	wire [4-1:0] node29129;
	wire [4-1:0] node29130;
	wire [4-1:0] node29132;
	wire [4-1:0] node29136;
	wire [4-1:0] node29137;
	wire [4-1:0] node29138;
	wire [4-1:0] node29139;
	wire [4-1:0] node29140;
	wire [4-1:0] node29141;
	wire [4-1:0] node29143;
	wire [4-1:0] node29146;
	wire [4-1:0] node29148;
	wire [4-1:0] node29151;
	wire [4-1:0] node29152;
	wire [4-1:0] node29154;
	wire [4-1:0] node29157;
	wire [4-1:0] node29159;
	wire [4-1:0] node29162;
	wire [4-1:0] node29163;
	wire [4-1:0] node29165;
	wire [4-1:0] node29166;
	wire [4-1:0] node29169;
	wire [4-1:0] node29172;
	wire [4-1:0] node29173;
	wire [4-1:0] node29175;
	wire [4-1:0] node29178;
	wire [4-1:0] node29180;
	wire [4-1:0] node29183;
	wire [4-1:0] node29184;
	wire [4-1:0] node29185;
	wire [4-1:0] node29186;
	wire [4-1:0] node29188;
	wire [4-1:0] node29191;
	wire [4-1:0] node29193;
	wire [4-1:0] node29196;
	wire [4-1:0] node29197;
	wire [4-1:0] node29199;
	wire [4-1:0] node29202;
	wire [4-1:0] node29205;
	wire [4-1:0] node29206;
	wire [4-1:0] node29207;
	wire [4-1:0] node29208;
	wire [4-1:0] node29212;
	wire [4-1:0] node29213;
	wire [4-1:0] node29217;
	wire [4-1:0] node29218;
	wire [4-1:0] node29219;
	wire [4-1:0] node29222;
	wire [4-1:0] node29223;
	wire [4-1:0] node29228;
	wire [4-1:0] node29229;
	wire [4-1:0] node29230;
	wire [4-1:0] node29231;
	wire [4-1:0] node29232;
	wire [4-1:0] node29234;
	wire [4-1:0] node29237;
	wire [4-1:0] node29239;
	wire [4-1:0] node29242;
	wire [4-1:0] node29243;
	wire [4-1:0] node29246;
	wire [4-1:0] node29248;
	wire [4-1:0] node29251;
	wire [4-1:0] node29252;
	wire [4-1:0] node29253;
	wire [4-1:0] node29256;
	wire [4-1:0] node29259;
	wire [4-1:0] node29260;
	wire [4-1:0] node29261;
	wire [4-1:0] node29263;
	wire [4-1:0] node29266;
	wire [4-1:0] node29267;
	wire [4-1:0] node29270;
	wire [4-1:0] node29274;
	wire [4-1:0] node29275;
	wire [4-1:0] node29276;
	wire [4-1:0] node29277;
	wire [4-1:0] node29278;
	wire [4-1:0] node29279;
	wire [4-1:0] node29284;
	wire [4-1:0] node29285;
	wire [4-1:0] node29289;
	wire [4-1:0] node29291;
	wire [4-1:0] node29294;
	wire [4-1:0] node29295;
	wire [4-1:0] node29296;
	wire [4-1:0] node29297;
	wire [4-1:0] node29300;
	wire [4-1:0] node29303;
	wire [4-1:0] node29305;
	wire [4-1:0] node29306;
	wire [4-1:0] node29309;
	wire [4-1:0] node29312;
	wire [4-1:0] node29313;
	wire [4-1:0] node29316;
	wire [4-1:0] node29319;
	wire [4-1:0] node29320;
	wire [4-1:0] node29321;
	wire [4-1:0] node29322;
	wire [4-1:0] node29323;
	wire [4-1:0] node29324;
	wire [4-1:0] node29325;
	wire [4-1:0] node29326;
	wire [4-1:0] node29328;
	wire [4-1:0] node29331;
	wire [4-1:0] node29333;
	wire [4-1:0] node29336;
	wire [4-1:0] node29337;
	wire [4-1:0] node29339;
	wire [4-1:0] node29342;
	wire [4-1:0] node29344;
	wire [4-1:0] node29347;
	wire [4-1:0] node29349;
	wire [4-1:0] node29350;
	wire [4-1:0] node29352;
	wire [4-1:0] node29355;
	wire [4-1:0] node29357;
	wire [4-1:0] node29360;
	wire [4-1:0] node29361;
	wire [4-1:0] node29362;
	wire [4-1:0] node29363;
	wire [4-1:0] node29367;
	wire [4-1:0] node29368;
	wire [4-1:0] node29370;
	wire [4-1:0] node29373;
	wire [4-1:0] node29374;
	wire [4-1:0] node29377;
	wire [4-1:0] node29380;
	wire [4-1:0] node29381;
	wire [4-1:0] node29383;
	wire [4-1:0] node29384;
	wire [4-1:0] node29387;
	wire [4-1:0] node29390;
	wire [4-1:0] node29391;
	wire [4-1:0] node29394;
	wire [4-1:0] node29397;
	wire [4-1:0] node29398;
	wire [4-1:0] node29399;
	wire [4-1:0] node29400;
	wire [4-1:0] node29401;
	wire [4-1:0] node29403;
	wire [4-1:0] node29407;
	wire [4-1:0] node29408;
	wire [4-1:0] node29409;
	wire [4-1:0] node29413;
	wire [4-1:0] node29416;
	wire [4-1:0] node29417;
	wire [4-1:0] node29418;
	wire [4-1:0] node29421;
	wire [4-1:0] node29422;
	wire [4-1:0] node29426;
	wire [4-1:0] node29427;
	wire [4-1:0] node29430;
	wire [4-1:0] node29431;
	wire [4-1:0] node29435;
	wire [4-1:0] node29436;
	wire [4-1:0] node29437;
	wire [4-1:0] node29438;
	wire [4-1:0] node29439;
	wire [4-1:0] node29443;
	wire [4-1:0] node29445;
	wire [4-1:0] node29448;
	wire [4-1:0] node29449;
	wire [4-1:0] node29450;
	wire [4-1:0] node29453;
	wire [4-1:0] node29456;
	wire [4-1:0] node29458;
	wire [4-1:0] node29461;
	wire [4-1:0] node29462;
	wire [4-1:0] node29463;
	wire [4-1:0] node29466;
	wire [4-1:0] node29467;
	wire [4-1:0] node29471;
	wire [4-1:0] node29472;
	wire [4-1:0] node29473;
	wire [4-1:0] node29477;
	wire [4-1:0] node29480;
	wire [4-1:0] node29481;
	wire [4-1:0] node29482;
	wire [4-1:0] node29483;
	wire [4-1:0] node29484;
	wire [4-1:0] node29485;
	wire [4-1:0] node29488;
	wire [4-1:0] node29491;
	wire [4-1:0] node29494;
	wire [4-1:0] node29495;
	wire [4-1:0] node29496;
	wire [4-1:0] node29497;
	wire [4-1:0] node29500;
	wire [4-1:0] node29503;
	wire [4-1:0] node29505;
	wire [4-1:0] node29508;
	wire [4-1:0] node29509;
	wire [4-1:0] node29510;
	wire [4-1:0] node29514;
	wire [4-1:0] node29516;
	wire [4-1:0] node29519;
	wire [4-1:0] node29520;
	wire [4-1:0] node29521;
	wire [4-1:0] node29522;
	wire [4-1:0] node29523;
	wire [4-1:0] node29526;
	wire [4-1:0] node29529;
	wire [4-1:0] node29530;
	wire [4-1:0] node29534;
	wire [4-1:0] node29535;
	wire [4-1:0] node29537;
	wire [4-1:0] node29540;
	wire [4-1:0] node29542;
	wire [4-1:0] node29545;
	wire [4-1:0] node29546;
	wire [4-1:0] node29547;
	wire [4-1:0] node29548;
	wire [4-1:0] node29551;
	wire [4-1:0] node29554;
	wire [4-1:0] node29556;
	wire [4-1:0] node29559;
	wire [4-1:0] node29560;
	wire [4-1:0] node29561;
	wire [4-1:0] node29565;
	wire [4-1:0] node29567;
	wire [4-1:0] node29570;
	wire [4-1:0] node29571;
	wire [4-1:0] node29572;
	wire [4-1:0] node29573;
	wire [4-1:0] node29574;
	wire [4-1:0] node29575;
	wire [4-1:0] node29579;
	wire [4-1:0] node29581;
	wire [4-1:0] node29584;
	wire [4-1:0] node29585;
	wire [4-1:0] node29586;
	wire [4-1:0] node29590;
	wire [4-1:0] node29591;
	wire [4-1:0] node29594;
	wire [4-1:0] node29597;
	wire [4-1:0] node29598;
	wire [4-1:0] node29599;
	wire [4-1:0] node29601;
	wire [4-1:0] node29604;
	wire [4-1:0] node29607;
	wire [4-1:0] node29608;
	wire [4-1:0] node29610;
	wire [4-1:0] node29613;
	wire [4-1:0] node29615;
	wire [4-1:0] node29618;
	wire [4-1:0] node29619;
	wire [4-1:0] node29620;
	wire [4-1:0] node29622;
	wire [4-1:0] node29624;
	wire [4-1:0] node29627;
	wire [4-1:0] node29628;
	wire [4-1:0] node29629;
	wire [4-1:0] node29632;
	wire [4-1:0] node29636;
	wire [4-1:0] node29637;
	wire [4-1:0] node29638;
	wire [4-1:0] node29639;
	wire [4-1:0] node29643;
	wire [4-1:0] node29645;
	wire [4-1:0] node29648;
	wire [4-1:0] node29649;
	wire [4-1:0] node29650;
	wire [4-1:0] node29653;
	wire [4-1:0] node29657;
	wire [4-1:0] node29658;
	wire [4-1:0] node29659;
	wire [4-1:0] node29660;
	wire [4-1:0] node29661;
	wire [4-1:0] node29662;
	wire [4-1:0] node29663;
	wire [4-1:0] node29666;
	wire [4-1:0] node29669;
	wire [4-1:0] node29671;
	wire [4-1:0] node29674;
	wire [4-1:0] node29675;
	wire [4-1:0] node29676;
	wire [4-1:0] node29679;
	wire [4-1:0] node29682;
	wire [4-1:0] node29683;
	wire [4-1:0] node29684;
	wire [4-1:0] node29687;
	wire [4-1:0] node29691;
	wire [4-1:0] node29692;
	wire [4-1:0] node29693;
	wire [4-1:0] node29694;
	wire [4-1:0] node29696;
	wire [4-1:0] node29699;
	wire [4-1:0] node29700;
	wire [4-1:0] node29703;
	wire [4-1:0] node29706;
	wire [4-1:0] node29707;
	wire [4-1:0] node29710;
	wire [4-1:0] node29711;
	wire [4-1:0] node29714;
	wire [4-1:0] node29717;
	wire [4-1:0] node29718;
	wire [4-1:0] node29719;
	wire [4-1:0] node29721;
	wire [4-1:0] node29724;
	wire [4-1:0] node29726;
	wire [4-1:0] node29729;
	wire [4-1:0] node29730;
	wire [4-1:0] node29731;
	wire [4-1:0] node29734;
	wire [4-1:0] node29737;
	wire [4-1:0] node29738;
	wire [4-1:0] node29741;
	wire [4-1:0] node29744;
	wire [4-1:0] node29745;
	wire [4-1:0] node29746;
	wire [4-1:0] node29747;
	wire [4-1:0] node29748;
	wire [4-1:0] node29750;
	wire [4-1:0] node29753;
	wire [4-1:0] node29754;
	wire [4-1:0] node29757;
	wire [4-1:0] node29760;
	wire [4-1:0] node29761;
	wire [4-1:0] node29762;
	wire [4-1:0] node29765;
	wire [4-1:0] node29768;
	wire [4-1:0] node29770;
	wire [4-1:0] node29773;
	wire [4-1:0] node29774;
	wire [4-1:0] node29775;
	wire [4-1:0] node29776;
	wire [4-1:0] node29780;
	wire [4-1:0] node29781;
	wire [4-1:0] node29784;
	wire [4-1:0] node29787;
	wire [4-1:0] node29788;
	wire [4-1:0] node29789;
	wire [4-1:0] node29792;
	wire [4-1:0] node29795;
	wire [4-1:0] node29796;
	wire [4-1:0] node29799;
	wire [4-1:0] node29802;
	wire [4-1:0] node29803;
	wire [4-1:0] node29804;
	wire [4-1:0] node29805;
	wire [4-1:0] node29808;
	wire [4-1:0] node29811;
	wire [4-1:0] node29812;
	wire [4-1:0] node29813;
	wire [4-1:0] node29816;
	wire [4-1:0] node29820;
	wire [4-1:0] node29821;
	wire [4-1:0] node29822;
	wire [4-1:0] node29823;
	wire [4-1:0] node29826;
	wire [4-1:0] node29829;
	wire [4-1:0] node29831;
	wire [4-1:0] node29834;
	wire [4-1:0] node29836;
	wire [4-1:0] node29837;
	wire [4-1:0] node29841;
	wire [4-1:0] node29842;
	wire [4-1:0] node29843;
	wire [4-1:0] node29844;
	wire [4-1:0] node29845;
	wire [4-1:0] node29846;
	wire [4-1:0] node29847;
	wire [4-1:0] node29850;
	wire [4-1:0] node29855;
	wire [4-1:0] node29856;
	wire [4-1:0] node29857;
	wire [4-1:0] node29858;
	wire [4-1:0] node29861;
	wire [4-1:0] node29864;
	wire [4-1:0] node29866;
	wire [4-1:0] node29869;
	wire [4-1:0] node29870;
	wire [4-1:0] node29871;
	wire [4-1:0] node29874;
	wire [4-1:0] node29877;
	wire [4-1:0] node29878;
	wire [4-1:0] node29881;
	wire [4-1:0] node29884;
	wire [4-1:0] node29885;
	wire [4-1:0] node29886;
	wire [4-1:0] node29887;
	wire [4-1:0] node29888;
	wire [4-1:0] node29892;
	wire [4-1:0] node29893;
	wire [4-1:0] node29896;
	wire [4-1:0] node29899;
	wire [4-1:0] node29900;
	wire [4-1:0] node29901;
	wire [4-1:0] node29904;
	wire [4-1:0] node29908;
	wire [4-1:0] node29909;
	wire [4-1:0] node29911;
	wire [4-1:0] node29914;
	wire [4-1:0] node29916;
	wire [4-1:0] node29919;
	wire [4-1:0] node29920;
	wire [4-1:0] node29921;
	wire [4-1:0] node29922;
	wire [4-1:0] node29923;
	wire [4-1:0] node29925;
	wire [4-1:0] node29928;
	wire [4-1:0] node29930;
	wire [4-1:0] node29933;
	wire [4-1:0] node29935;
	wire [4-1:0] node29936;
	wire [4-1:0] node29939;
	wire [4-1:0] node29942;
	wire [4-1:0] node29943;
	wire [4-1:0] node29944;
	wire [4-1:0] node29947;
	wire [4-1:0] node29950;
	wire [4-1:0] node29952;
	wire [4-1:0] node29955;
	wire [4-1:0] node29956;
	wire [4-1:0] node29957;
	wire [4-1:0] node29960;
	wire [4-1:0] node29963;
	wire [4-1:0] node29964;
	wire [4-1:0] node29965;
	wire [4-1:0] node29968;
	wire [4-1:0] node29971;
	wire [4-1:0] node29972;
	wire [4-1:0] node29975;
	wire [4-1:0] node29978;
	wire [4-1:0] node29979;
	wire [4-1:0] node29980;
	wire [4-1:0] node29981;
	wire [4-1:0] node29982;
	wire [4-1:0] node29983;
	wire [4-1:0] node29984;
	wire [4-1:0] node29985;
	wire [4-1:0] node29986;
	wire [4-1:0] node29988;
	wire [4-1:0] node29991;
	wire [4-1:0] node29993;
	wire [4-1:0] node29996;
	wire [4-1:0] node29997;
	wire [4-1:0] node30000;
	wire [4-1:0] node30002;
	wire [4-1:0] node30005;
	wire [4-1:0] node30006;
	wire [4-1:0] node30008;
	wire [4-1:0] node30011;
	wire [4-1:0] node30012;
	wire [4-1:0] node30013;
	wire [4-1:0] node30017;
	wire [4-1:0] node30018;
	wire [4-1:0] node30022;
	wire [4-1:0] node30023;
	wire [4-1:0] node30024;
	wire [4-1:0] node30025;
	wire [4-1:0] node30026;
	wire [4-1:0] node30029;
	wire [4-1:0] node30032;
	wire [4-1:0] node30034;
	wire [4-1:0] node30037;
	wire [4-1:0] node30038;
	wire [4-1:0] node30039;
	wire [4-1:0] node30043;
	wire [4-1:0] node30046;
	wire [4-1:0] node30047;
	wire [4-1:0] node30048;
	wire [4-1:0] node30049;
	wire [4-1:0] node30052;
	wire [4-1:0] node30055;
	wire [4-1:0] node30057;
	wire [4-1:0] node30060;
	wire [4-1:0] node30062;
	wire [4-1:0] node30065;
	wire [4-1:0] node30066;
	wire [4-1:0] node30067;
	wire [4-1:0] node30068;
	wire [4-1:0] node30069;
	wire [4-1:0] node30072;
	wire [4-1:0] node30075;
	wire [4-1:0] node30076;
	wire [4-1:0] node30077;
	wire [4-1:0] node30080;
	wire [4-1:0] node30083;
	wire [4-1:0] node30084;
	wire [4-1:0] node30087;
	wire [4-1:0] node30090;
	wire [4-1:0] node30091;
	wire [4-1:0] node30092;
	wire [4-1:0] node30095;
	wire [4-1:0] node30097;
	wire [4-1:0] node30100;
	wire [4-1:0] node30101;
	wire [4-1:0] node30103;
	wire [4-1:0] node30106;
	wire [4-1:0] node30107;
	wire [4-1:0] node30111;
	wire [4-1:0] node30112;
	wire [4-1:0] node30113;
	wire [4-1:0] node30114;
	wire [4-1:0] node30117;
	wire [4-1:0] node30118;
	wire [4-1:0] node30122;
	wire [4-1:0] node30123;
	wire [4-1:0] node30126;
	wire [4-1:0] node30129;
	wire [4-1:0] node30130;
	wire [4-1:0] node30131;
	wire [4-1:0] node30132;
	wire [4-1:0] node30135;
	wire [4-1:0] node30138;
	wire [4-1:0] node30141;
	wire [4-1:0] node30142;
	wire [4-1:0] node30145;
	wire [4-1:0] node30148;
	wire [4-1:0] node30149;
	wire [4-1:0] node30150;
	wire [4-1:0] node30151;
	wire [4-1:0] node30152;
	wire [4-1:0] node30154;
	wire [4-1:0] node30157;
	wire [4-1:0] node30158;
	wire [4-1:0] node30160;
	wire [4-1:0] node30163;
	wire [4-1:0] node30166;
	wire [4-1:0] node30167;
	wire [4-1:0] node30168;
	wire [4-1:0] node30171;
	wire [4-1:0] node30172;
	wire [4-1:0] node30176;
	wire [4-1:0] node30177;
	wire [4-1:0] node30181;
	wire [4-1:0] node30182;
	wire [4-1:0] node30183;
	wire [4-1:0] node30185;
	wire [4-1:0] node30186;
	wire [4-1:0] node30189;
	wire [4-1:0] node30192;
	wire [4-1:0] node30193;
	wire [4-1:0] node30194;
	wire [4-1:0] node30197;
	wire [4-1:0] node30200;
	wire [4-1:0] node30201;
	wire [4-1:0] node30205;
	wire [4-1:0] node30206;
	wire [4-1:0] node30207;
	wire [4-1:0] node30211;
	wire [4-1:0] node30212;
	wire [4-1:0] node30214;
	wire [4-1:0] node30217;
	wire [4-1:0] node30220;
	wire [4-1:0] node30221;
	wire [4-1:0] node30222;
	wire [4-1:0] node30223;
	wire [4-1:0] node30224;
	wire [4-1:0] node30227;
	wire [4-1:0] node30230;
	wire [4-1:0] node30231;
	wire [4-1:0] node30232;
	wire [4-1:0] node30236;
	wire [4-1:0] node30237;
	wire [4-1:0] node30240;
	wire [4-1:0] node30243;
	wire [4-1:0] node30244;
	wire [4-1:0] node30245;
	wire [4-1:0] node30246;
	wire [4-1:0] node30249;
	wire [4-1:0] node30252;
	wire [4-1:0] node30253;
	wire [4-1:0] node30257;
	wire [4-1:0] node30258;
	wire [4-1:0] node30259;
	wire [4-1:0] node30264;
	wire [4-1:0] node30265;
	wire [4-1:0] node30266;
	wire [4-1:0] node30268;
	wire [4-1:0] node30271;
	wire [4-1:0] node30272;
	wire [4-1:0] node30273;
	wire [4-1:0] node30277;
	wire [4-1:0] node30278;
	wire [4-1:0] node30281;
	wire [4-1:0] node30284;
	wire [4-1:0] node30285;
	wire [4-1:0] node30287;
	wire [4-1:0] node30289;
	wire [4-1:0] node30292;
	wire [4-1:0] node30293;
	wire [4-1:0] node30295;
	wire [4-1:0] node30298;
	wire [4-1:0] node30300;
	wire [4-1:0] node30303;
	wire [4-1:0] node30304;
	wire [4-1:0] node30305;
	wire [4-1:0] node30306;
	wire [4-1:0] node30307;
	wire [4-1:0] node30308;
	wire [4-1:0] node30309;
	wire [4-1:0] node30312;
	wire [4-1:0] node30315;
	wire [4-1:0] node30317;
	wire [4-1:0] node30320;
	wire [4-1:0] node30321;
	wire [4-1:0] node30323;
	wire [4-1:0] node30326;
	wire [4-1:0] node30329;
	wire [4-1:0] node30330;
	wire [4-1:0] node30333;
	wire [4-1:0] node30334;
	wire [4-1:0] node30336;
	wire [4-1:0] node30339;
	wire [4-1:0] node30340;
	wire [4-1:0] node30344;
	wire [4-1:0] node30345;
	wire [4-1:0] node30346;
	wire [4-1:0] node30347;
	wire [4-1:0] node30348;
	wire [4-1:0] node30349;
	wire [4-1:0] node30352;
	wire [4-1:0] node30355;
	wire [4-1:0] node30356;
	wire [4-1:0] node30359;
	wire [4-1:0] node30362;
	wire [4-1:0] node30363;
	wire [4-1:0] node30364;
	wire [4-1:0] node30367;
	wire [4-1:0] node30371;
	wire [4-1:0] node30372;
	wire [4-1:0] node30373;
	wire [4-1:0] node30376;
	wire [4-1:0] node30379;
	wire [4-1:0] node30380;
	wire [4-1:0] node30381;
	wire [4-1:0] node30384;
	wire [4-1:0] node30387;
	wire [4-1:0] node30388;
	wire [4-1:0] node30392;
	wire [4-1:0] node30393;
	wire [4-1:0] node30394;
	wire [4-1:0] node30397;
	wire [4-1:0] node30399;
	wire [4-1:0] node30402;
	wire [4-1:0] node30403;
	wire [4-1:0] node30404;
	wire [4-1:0] node30408;
	wire [4-1:0] node30409;
	wire [4-1:0] node30412;
	wire [4-1:0] node30415;
	wire [4-1:0] node30416;
	wire [4-1:0] node30417;
	wire [4-1:0] node30418;
	wire [4-1:0] node30419;
	wire [4-1:0] node30421;
	wire [4-1:0] node30424;
	wire [4-1:0] node30427;
	wire [4-1:0] node30428;
	wire [4-1:0] node30430;
	wire [4-1:0] node30433;
	wire [4-1:0] node30435;
	wire [4-1:0] node30438;
	wire [4-1:0] node30439;
	wire [4-1:0] node30440;
	wire [4-1:0] node30441;
	wire [4-1:0] node30444;
	wire [4-1:0] node30447;
	wire [4-1:0] node30448;
	wire [4-1:0] node30451;
	wire [4-1:0] node30454;
	wire [4-1:0] node30455;
	wire [4-1:0] node30458;
	wire [4-1:0] node30461;
	wire [4-1:0] node30462;
	wire [4-1:0] node30463;
	wire [4-1:0] node30464;
	wire [4-1:0] node30465;
	wire [4-1:0] node30468;
	wire [4-1:0] node30471;
	wire [4-1:0] node30472;
	wire [4-1:0] node30476;
	wire [4-1:0] node30477;
	wire [4-1:0] node30480;
	wire [4-1:0] node30483;
	wire [4-1:0] node30484;
	wire [4-1:0] node30485;
	wire [4-1:0] node30486;
	wire [4-1:0] node30487;
	wire [4-1:0] node30491;
	wire [4-1:0] node30494;
	wire [4-1:0] node30495;
	wire [4-1:0] node30496;
	wire [4-1:0] node30501;
	wire [4-1:0] node30502;
	wire [4-1:0] node30503;
	wire [4-1:0] node30507;
	wire [4-1:0] node30510;
	wire [4-1:0] node30511;
	wire [4-1:0] node30512;
	wire [4-1:0] node30513;
	wire [4-1:0] node30514;
	wire [4-1:0] node30515;
	wire [4-1:0] node30516;
	wire [4-1:0] node30517;
	wire [4-1:0] node30521;
	wire [4-1:0] node30522;
	wire [4-1:0] node30523;
	wire [4-1:0] node30526;
	wire [4-1:0] node30530;
	wire [4-1:0] node30531;
	wire [4-1:0] node30532;
	wire [4-1:0] node30534;
	wire [4-1:0] node30538;
	wire [4-1:0] node30540;
	wire [4-1:0] node30541;
	wire [4-1:0] node30545;
	wire [4-1:0] node30546;
	wire [4-1:0] node30547;
	wire [4-1:0] node30549;
	wire [4-1:0] node30550;
	wire [4-1:0] node30554;
	wire [4-1:0] node30555;
	wire [4-1:0] node30557;
	wire [4-1:0] node30560;
	wire [4-1:0] node30561;
	wire [4-1:0] node30565;
	wire [4-1:0] node30566;
	wire [4-1:0] node30567;
	wire [4-1:0] node30569;
	wire [4-1:0] node30572;
	wire [4-1:0] node30575;
	wire [4-1:0] node30576;
	wire [4-1:0] node30577;
	wire [4-1:0] node30581;
	wire [4-1:0] node30584;
	wire [4-1:0] node30585;
	wire [4-1:0] node30586;
	wire [4-1:0] node30587;
	wire [4-1:0] node30588;
	wire [4-1:0] node30592;
	wire [4-1:0] node30593;
	wire [4-1:0] node30595;
	wire [4-1:0] node30598;
	wire [4-1:0] node30599;
	wire [4-1:0] node30602;
	wire [4-1:0] node30605;
	wire [4-1:0] node30606;
	wire [4-1:0] node30607;
	wire [4-1:0] node30608;
	wire [4-1:0] node30611;
	wire [4-1:0] node30615;
	wire [4-1:0] node30617;
	wire [4-1:0] node30618;
	wire [4-1:0] node30621;
	wire [4-1:0] node30624;
	wire [4-1:0] node30625;
	wire [4-1:0] node30626;
	wire [4-1:0] node30627;
	wire [4-1:0] node30630;
	wire [4-1:0] node30631;
	wire [4-1:0] node30635;
	wire [4-1:0] node30636;
	wire [4-1:0] node30639;
	wire [4-1:0] node30642;
	wire [4-1:0] node30643;
	wire [4-1:0] node30644;
	wire [4-1:0] node30647;
	wire [4-1:0] node30648;
	wire [4-1:0] node30652;
	wire [4-1:0] node30653;
	wire [4-1:0] node30656;
	wire [4-1:0] node30659;
	wire [4-1:0] node30660;
	wire [4-1:0] node30661;
	wire [4-1:0] node30662;
	wire [4-1:0] node30663;
	wire [4-1:0] node30665;
	wire [4-1:0] node30666;
	wire [4-1:0] node30669;
	wire [4-1:0] node30672;
	wire [4-1:0] node30673;
	wire [4-1:0] node30676;
	wire [4-1:0] node30679;
	wire [4-1:0] node30680;
	wire [4-1:0] node30681;
	wire [4-1:0] node30684;
	wire [4-1:0] node30687;
	wire [4-1:0] node30690;
	wire [4-1:0] node30691;
	wire [4-1:0] node30692;
	wire [4-1:0] node30694;
	wire [4-1:0] node30696;
	wire [4-1:0] node30699;
	wire [4-1:0] node30700;
	wire [4-1:0] node30701;
	wire [4-1:0] node30704;
	wire [4-1:0] node30707;
	wire [4-1:0] node30710;
	wire [4-1:0] node30711;
	wire [4-1:0] node30712;
	wire [4-1:0] node30713;
	wire [4-1:0] node30717;
	wire [4-1:0] node30718;
	wire [4-1:0] node30721;
	wire [4-1:0] node30724;
	wire [4-1:0] node30726;
	wire [4-1:0] node30727;
	wire [4-1:0] node30730;
	wire [4-1:0] node30733;
	wire [4-1:0] node30734;
	wire [4-1:0] node30735;
	wire [4-1:0] node30736;
	wire [4-1:0] node30737;
	wire [4-1:0] node30738;
	wire [4-1:0] node30741;
	wire [4-1:0] node30744;
	wire [4-1:0] node30746;
	wire [4-1:0] node30749;
	wire [4-1:0] node30750;
	wire [4-1:0] node30751;
	wire [4-1:0] node30756;
	wire [4-1:0] node30757;
	wire [4-1:0] node30758;
	wire [4-1:0] node30759;
	wire [4-1:0] node30762;
	wire [4-1:0] node30766;
	wire [4-1:0] node30767;
	wire [4-1:0] node30770;
	wire [4-1:0] node30773;
	wire [4-1:0] node30774;
	wire [4-1:0] node30775;
	wire [4-1:0] node30778;
	wire [4-1:0] node30779;
	wire [4-1:0] node30780;
	wire [4-1:0] node30783;
	wire [4-1:0] node30786;
	wire [4-1:0] node30787;
	wire [4-1:0] node30790;
	wire [4-1:0] node30793;
	wire [4-1:0] node30794;
	wire [4-1:0] node30795;
	wire [4-1:0] node30796;
	wire [4-1:0] node30799;
	wire [4-1:0] node30803;
	wire [4-1:0] node30804;
	wire [4-1:0] node30807;
	wire [4-1:0] node30810;
	wire [4-1:0] node30811;
	wire [4-1:0] node30812;
	wire [4-1:0] node30813;
	wire [4-1:0] node30814;
	wire [4-1:0] node30815;
	wire [4-1:0] node30818;
	wire [4-1:0] node30820;
	wire [4-1:0] node30823;
	wire [4-1:0] node30824;
	wire [4-1:0] node30826;
	wire [4-1:0] node30829;
	wire [4-1:0] node30830;
	wire [4-1:0] node30833;
	wire [4-1:0] node30836;
	wire [4-1:0] node30837;
	wire [4-1:0] node30838;
	wire [4-1:0] node30839;
	wire [4-1:0] node30842;
	wire [4-1:0] node30845;
	wire [4-1:0] node30846;
	wire [4-1:0] node30850;
	wire [4-1:0] node30851;
	wire [4-1:0] node30853;
	wire [4-1:0] node30854;
	wire [4-1:0] node30857;
	wire [4-1:0] node30860;
	wire [4-1:0] node30861;
	wire [4-1:0] node30862;
	wire [4-1:0] node30866;
	wire [4-1:0] node30867;
	wire [4-1:0] node30870;
	wire [4-1:0] node30873;
	wire [4-1:0] node30874;
	wire [4-1:0] node30875;
	wire [4-1:0] node30876;
	wire [4-1:0] node30877;
	wire [4-1:0] node30880;
	wire [4-1:0] node30883;
	wire [4-1:0] node30884;
	wire [4-1:0] node30887;
	wire [4-1:0] node30890;
	wire [4-1:0] node30891;
	wire [4-1:0] node30892;
	wire [4-1:0] node30895;
	wire [4-1:0] node30898;
	wire [4-1:0] node30899;
	wire [4-1:0] node30902;
	wire [4-1:0] node30905;
	wire [4-1:0] node30906;
	wire [4-1:0] node30907;
	wire [4-1:0] node30909;
	wire [4-1:0] node30910;
	wire [4-1:0] node30913;
	wire [4-1:0] node30916;
	wire [4-1:0] node30918;
	wire [4-1:0] node30921;
	wire [4-1:0] node30922;
	wire [4-1:0] node30925;
	wire [4-1:0] node30928;
	wire [4-1:0] node30929;
	wire [4-1:0] node30930;
	wire [4-1:0] node30931;
	wire [4-1:0] node30932;
	wire [4-1:0] node30933;
	wire [4-1:0] node30936;
	wire [4-1:0] node30939;
	wire [4-1:0] node30940;
	wire [4-1:0] node30941;
	wire [4-1:0] node30945;
	wire [4-1:0] node30947;
	wire [4-1:0] node30950;
	wire [4-1:0] node30951;
	wire [4-1:0] node30952;
	wire [4-1:0] node30956;
	wire [4-1:0] node30957;
	wire [4-1:0] node30959;
	wire [4-1:0] node30962;
	wire [4-1:0] node30964;
	wire [4-1:0] node30967;
	wire [4-1:0] node30968;
	wire [4-1:0] node30969;
	wire [4-1:0] node30971;
	wire [4-1:0] node30974;
	wire [4-1:0] node30976;
	wire [4-1:0] node30979;
	wire [4-1:0] node30980;
	wire [4-1:0] node30981;
	wire [4-1:0] node30984;
	wire [4-1:0] node30987;
	wire [4-1:0] node30988;
	wire [4-1:0] node30991;
	wire [4-1:0] node30994;
	wire [4-1:0] node30995;
	wire [4-1:0] node30996;
	wire [4-1:0] node30997;
	wire [4-1:0] node30998;
	wire [4-1:0] node31001;
	wire [4-1:0] node31004;
	wire [4-1:0] node31006;
	wire [4-1:0] node31009;
	wire [4-1:0] node31010;
	wire [4-1:0] node31011;
	wire [4-1:0] node31015;
	wire [4-1:0] node31016;
	wire [4-1:0] node31017;
	wire [4-1:0] node31020;
	wire [4-1:0] node31023;
	wire [4-1:0] node31024;
	wire [4-1:0] node31027;
	wire [4-1:0] node31030;
	wire [4-1:0] node31031;
	wire [4-1:0] node31032;
	wire [4-1:0] node31033;
	wire [4-1:0] node31036;
	wire [4-1:0] node31039;
	wire [4-1:0] node31041;
	wire [4-1:0] node31044;
	wire [4-1:0] node31045;
	wire [4-1:0] node31046;
	wire [4-1:0] node31047;
	wire [4-1:0] node31050;
	wire [4-1:0] node31053;
	wire [4-1:0] node31055;
	wire [4-1:0] node31058;
	wire [4-1:0] node31060;
	wire [4-1:0] node31063;
	wire [4-1:0] node31064;
	wire [4-1:0] node31065;
	wire [4-1:0] node31066;
	wire [4-1:0] node31067;
	wire [4-1:0] node31068;
	wire [4-1:0] node31069;
	wire [4-1:0] node31070;
	wire [4-1:0] node31071;
	wire [4-1:0] node31072;
	wire [4-1:0] node31073;
	wire [4-1:0] node31076;
	wire [4-1:0] node31079;
	wire [4-1:0] node31080;
	wire [4-1:0] node31083;
	wire [4-1:0] node31086;
	wire [4-1:0] node31088;
	wire [4-1:0] node31091;
	wire [4-1:0] node31092;
	wire [4-1:0] node31093;
	wire [4-1:0] node31094;
	wire [4-1:0] node31098;
	wire [4-1:0] node31100;
	wire [4-1:0] node31103;
	wire [4-1:0] node31104;
	wire [4-1:0] node31105;
	wire [4-1:0] node31110;
	wire [4-1:0] node31111;
	wire [4-1:0] node31112;
	wire [4-1:0] node31114;
	wire [4-1:0] node31116;
	wire [4-1:0] node31119;
	wire [4-1:0] node31120;
	wire [4-1:0] node31121;
	wire [4-1:0] node31124;
	wire [4-1:0] node31127;
	wire [4-1:0] node31128;
	wire [4-1:0] node31132;
	wire [4-1:0] node31133;
	wire [4-1:0] node31134;
	wire [4-1:0] node31136;
	wire [4-1:0] node31139;
	wire [4-1:0] node31141;
	wire [4-1:0] node31144;
	wire [4-1:0] node31145;
	wire [4-1:0] node31146;
	wire [4-1:0] node31150;
	wire [4-1:0] node31151;
	wire [4-1:0] node31154;
	wire [4-1:0] node31157;
	wire [4-1:0] node31158;
	wire [4-1:0] node31159;
	wire [4-1:0] node31160;
	wire [4-1:0] node31161;
	wire [4-1:0] node31163;
	wire [4-1:0] node31167;
	wire [4-1:0] node31168;
	wire [4-1:0] node31169;
	wire [4-1:0] node31173;
	wire [4-1:0] node31176;
	wire [4-1:0] node31177;
	wire [4-1:0] node31178;
	wire [4-1:0] node31179;
	wire [4-1:0] node31182;
	wire [4-1:0] node31186;
	wire [4-1:0] node31188;
	wire [4-1:0] node31189;
	wire [4-1:0] node31192;
	wire [4-1:0] node31195;
	wire [4-1:0] node31196;
	wire [4-1:0] node31197;
	wire [4-1:0] node31200;
	wire [4-1:0] node31202;
	wire [4-1:0] node31203;
	wire [4-1:0] node31206;
	wire [4-1:0] node31209;
	wire [4-1:0] node31210;
	wire [4-1:0] node31211;
	wire [4-1:0] node31212;
	wire [4-1:0] node31216;
	wire [4-1:0] node31218;
	wire [4-1:0] node31221;
	wire [4-1:0] node31222;
	wire [4-1:0] node31223;
	wire [4-1:0] node31227;
	wire [4-1:0] node31229;
	wire [4-1:0] node31232;
	wire [4-1:0] node31233;
	wire [4-1:0] node31234;
	wire [4-1:0] node31235;
	wire [4-1:0] node31236;
	wire [4-1:0] node31237;
	wire [4-1:0] node31240;
	wire [4-1:0] node31243;
	wire [4-1:0] node31245;
	wire [4-1:0] node31248;
	wire [4-1:0] node31249;
	wire [4-1:0] node31250;
	wire [4-1:0] node31251;
	wire [4-1:0] node31254;
	wire [4-1:0] node31257;
	wire [4-1:0] node31258;
	wire [4-1:0] node31261;
	wire [4-1:0] node31264;
	wire [4-1:0] node31265;
	wire [4-1:0] node31268;
	wire [4-1:0] node31271;
	wire [4-1:0] node31272;
	wire [4-1:0] node31273;
	wire [4-1:0] node31274;
	wire [4-1:0] node31275;
	wire [4-1:0] node31278;
	wire [4-1:0] node31281;
	wire [4-1:0] node31282;
	wire [4-1:0] node31285;
	wire [4-1:0] node31288;
	wire [4-1:0] node31289;
	wire [4-1:0] node31290;
	wire [4-1:0] node31294;
	wire [4-1:0] node31295;
	wire [4-1:0] node31299;
	wire [4-1:0] node31300;
	wire [4-1:0] node31302;
	wire [4-1:0] node31303;
	wire [4-1:0] node31306;
	wire [4-1:0] node31309;
	wire [4-1:0] node31310;
	wire [4-1:0] node31311;
	wire [4-1:0] node31314;
	wire [4-1:0] node31318;
	wire [4-1:0] node31319;
	wire [4-1:0] node31320;
	wire [4-1:0] node31321;
	wire [4-1:0] node31322;
	wire [4-1:0] node31323;
	wire [4-1:0] node31326;
	wire [4-1:0] node31329;
	wire [4-1:0] node31330;
	wire [4-1:0] node31333;
	wire [4-1:0] node31336;
	wire [4-1:0] node31337;
	wire [4-1:0] node31338;
	wire [4-1:0] node31342;
	wire [4-1:0] node31345;
	wire [4-1:0] node31346;
	wire [4-1:0] node31347;
	wire [4-1:0] node31350;
	wire [4-1:0] node31353;
	wire [4-1:0] node31354;
	wire [4-1:0] node31356;
	wire [4-1:0] node31359;
	wire [4-1:0] node31360;
	wire [4-1:0] node31364;
	wire [4-1:0] node31365;
	wire [4-1:0] node31366;
	wire [4-1:0] node31367;
	wire [4-1:0] node31368;
	wire [4-1:0] node31373;
	wire [4-1:0] node31374;
	wire [4-1:0] node31375;
	wire [4-1:0] node31378;
	wire [4-1:0] node31381;
	wire [4-1:0] node31383;
	wire [4-1:0] node31386;
	wire [4-1:0] node31387;
	wire [4-1:0] node31388;
	wire [4-1:0] node31389;
	wire [4-1:0] node31392;
	wire [4-1:0] node31396;
	wire [4-1:0] node31397;
	wire [4-1:0] node31398;
	wire [4-1:0] node31401;
	wire [4-1:0] node31404;
	wire [4-1:0] node31405;
	wire [4-1:0] node31408;
	wire [4-1:0] node31411;
	wire [4-1:0] node31412;
	wire [4-1:0] node31413;
	wire [4-1:0] node31414;
	wire [4-1:0] node31415;
	wire [4-1:0] node31416;
	wire [4-1:0] node31417;
	wire [4-1:0] node31418;
	wire [4-1:0] node31421;
	wire [4-1:0] node31424;
	wire [4-1:0] node31425;
	wire [4-1:0] node31429;
	wire [4-1:0] node31430;
	wire [4-1:0] node31432;
	wire [4-1:0] node31436;
	wire [4-1:0] node31437;
	wire [4-1:0] node31438;
	wire [4-1:0] node31442;
	wire [4-1:0] node31443;
	wire [4-1:0] node31447;
	wire [4-1:0] node31448;
	wire [4-1:0] node31449;
	wire [4-1:0] node31450;
	wire [4-1:0] node31454;
	wire [4-1:0] node31455;
	wire [4-1:0] node31459;
	wire [4-1:0] node31460;
	wire [4-1:0] node31461;
	wire [4-1:0] node31465;
	wire [4-1:0] node31466;
	wire [4-1:0] node31470;
	wire [4-1:0] node31471;
	wire [4-1:0] node31472;
	wire [4-1:0] node31473;
	wire [4-1:0] node31474;
	wire [4-1:0] node31475;
	wire [4-1:0] node31480;
	wire [4-1:0] node31482;
	wire [4-1:0] node31485;
	wire [4-1:0] node31486;
	wire [4-1:0] node31488;
	wire [4-1:0] node31491;
	wire [4-1:0] node31493;
	wire [4-1:0] node31496;
	wire [4-1:0] node31497;
	wire [4-1:0] node31498;
	wire [4-1:0] node31499;
	wire [4-1:0] node31502;
	wire [4-1:0] node31505;
	wire [4-1:0] node31506;
	wire [4-1:0] node31509;
	wire [4-1:0] node31512;
	wire [4-1:0] node31513;
	wire [4-1:0] node31515;
	wire [4-1:0] node31516;
	wire [4-1:0] node31520;
	wire [4-1:0] node31521;
	wire [4-1:0] node31522;
	wire [4-1:0] node31527;
	wire [4-1:0] node31528;
	wire [4-1:0] node31529;
	wire [4-1:0] node31530;
	wire [4-1:0] node31531;
	wire [4-1:0] node31532;
	wire [4-1:0] node31533;
	wire [4-1:0] node31538;
	wire [4-1:0] node31539;
	wire [4-1:0] node31540;
	wire [4-1:0] node31544;
	wire [4-1:0] node31545;
	wire [4-1:0] node31549;
	wire [4-1:0] node31550;
	wire [4-1:0] node31551;
	wire [4-1:0] node31552;
	wire [4-1:0] node31555;
	wire [4-1:0] node31559;
	wire [4-1:0] node31560;
	wire [4-1:0] node31563;
	wire [4-1:0] node31566;
	wire [4-1:0] node31567;
	wire [4-1:0] node31568;
	wire [4-1:0] node31569;
	wire [4-1:0] node31571;
	wire [4-1:0] node31574;
	wire [4-1:0] node31576;
	wire [4-1:0] node31579;
	wire [4-1:0] node31580;
	wire [4-1:0] node31583;
	wire [4-1:0] node31586;
	wire [4-1:0] node31587;
	wire [4-1:0] node31588;
	wire [4-1:0] node31591;
	wire [4-1:0] node31594;
	wire [4-1:0] node31595;
	wire [4-1:0] node31596;
	wire [4-1:0] node31599;
	wire [4-1:0] node31603;
	wire [4-1:0] node31604;
	wire [4-1:0] node31605;
	wire [4-1:0] node31606;
	wire [4-1:0] node31607;
	wire [4-1:0] node31608;
	wire [4-1:0] node31611;
	wire [4-1:0] node31614;
	wire [4-1:0] node31615;
	wire [4-1:0] node31619;
	wire [4-1:0] node31620;
	wire [4-1:0] node31622;
	wire [4-1:0] node31625;
	wire [4-1:0] node31626;
	wire [4-1:0] node31629;
	wire [4-1:0] node31632;
	wire [4-1:0] node31633;
	wire [4-1:0] node31637;
	wire [4-1:0] node31638;
	wire [4-1:0] node31640;
	wire [4-1:0] node31642;
	wire [4-1:0] node31644;
	wire [4-1:0] node31647;
	wire [4-1:0] node31648;
	wire [4-1:0] node31649;
	wire [4-1:0] node31652;
	wire [4-1:0] node31655;
	wire [4-1:0] node31656;
	wire [4-1:0] node31659;
	wire [4-1:0] node31662;
	wire [4-1:0] node31663;
	wire [4-1:0] node31664;
	wire [4-1:0] node31665;
	wire [4-1:0] node31666;
	wire [4-1:0] node31667;
	wire [4-1:0] node31668;
	wire [4-1:0] node31671;
	wire [4-1:0] node31672;
	wire [4-1:0] node31673;
	wire [4-1:0] node31676;
	wire [4-1:0] node31680;
	wire [4-1:0] node31681;
	wire [4-1:0] node31682;
	wire [4-1:0] node31683;
	wire [4-1:0] node31686;
	wire [4-1:0] node31689;
	wire [4-1:0] node31691;
	wire [4-1:0] node31694;
	wire [4-1:0] node31695;
	wire [4-1:0] node31697;
	wire [4-1:0] node31700;
	wire [4-1:0] node31701;
	wire [4-1:0] node31705;
	wire [4-1:0] node31706;
	wire [4-1:0] node31707;
	wire [4-1:0] node31708;
	wire [4-1:0] node31709;
	wire [4-1:0] node31712;
	wire [4-1:0] node31715;
	wire [4-1:0] node31717;
	wire [4-1:0] node31720;
	wire [4-1:0] node31721;
	wire [4-1:0] node31722;
	wire [4-1:0] node31725;
	wire [4-1:0] node31728;
	wire [4-1:0] node31730;
	wire [4-1:0] node31733;
	wire [4-1:0] node31734;
	wire [4-1:0] node31735;
	wire [4-1:0] node31736;
	wire [4-1:0] node31739;
	wire [4-1:0] node31742;
	wire [4-1:0] node31743;
	wire [4-1:0] node31747;
	wire [4-1:0] node31748;
	wire [4-1:0] node31751;
	wire [4-1:0] node31753;
	wire [4-1:0] node31756;
	wire [4-1:0] node31757;
	wire [4-1:0] node31758;
	wire [4-1:0] node31759;
	wire [4-1:0] node31760;
	wire [4-1:0] node31761;
	wire [4-1:0] node31764;
	wire [4-1:0] node31767;
	wire [4-1:0] node31768;
	wire [4-1:0] node31772;
	wire [4-1:0] node31773;
	wire [4-1:0] node31775;
	wire [4-1:0] node31778;
	wire [4-1:0] node31779;
	wire [4-1:0] node31782;
	wire [4-1:0] node31785;
	wire [4-1:0] node31786;
	wire [4-1:0] node31788;
	wire [4-1:0] node31789;
	wire [4-1:0] node31793;
	wire [4-1:0] node31794;
	wire [4-1:0] node31797;
	wire [4-1:0] node31798;
	wire [4-1:0] node31802;
	wire [4-1:0] node31803;
	wire [4-1:0] node31804;
	wire [4-1:0] node31806;
	wire [4-1:0] node31807;
	wire [4-1:0] node31810;
	wire [4-1:0] node31813;
	wire [4-1:0] node31814;
	wire [4-1:0] node31815;
	wire [4-1:0] node31819;
	wire [4-1:0] node31820;
	wire [4-1:0] node31823;
	wire [4-1:0] node31826;
	wire [4-1:0] node31827;
	wire [4-1:0] node31828;
	wire [4-1:0] node31830;
	wire [4-1:0] node31833;
	wire [4-1:0] node31834;
	wire [4-1:0] node31838;
	wire [4-1:0] node31839;
	wire [4-1:0] node31840;
	wire [4-1:0] node31843;
	wire [4-1:0] node31846;
	wire [4-1:0] node31847;
	wire [4-1:0] node31850;
	wire [4-1:0] node31853;
	wire [4-1:0] node31854;
	wire [4-1:0] node31855;
	wire [4-1:0] node31856;
	wire [4-1:0] node31857;
	wire [4-1:0] node31858;
	wire [4-1:0] node31861;
	wire [4-1:0] node31864;
	wire [4-1:0] node31865;
	wire [4-1:0] node31868;
	wire [4-1:0] node31871;
	wire [4-1:0] node31872;
	wire [4-1:0] node31874;
	wire [4-1:0] node31875;
	wire [4-1:0] node31878;
	wire [4-1:0] node31881;
	wire [4-1:0] node31882;
	wire [4-1:0] node31886;
	wire [4-1:0] node31887;
	wire [4-1:0] node31888;
	wire [4-1:0] node31889;
	wire [4-1:0] node31890;
	wire [4-1:0] node31894;
	wire [4-1:0] node31895;
	wire [4-1:0] node31898;
	wire [4-1:0] node31901;
	wire [4-1:0] node31902;
	wire [4-1:0] node31906;
	wire [4-1:0] node31907;
	wire [4-1:0] node31908;
	wire [4-1:0] node31909;
	wire [4-1:0] node31913;
	wire [4-1:0] node31914;
	wire [4-1:0] node31917;
	wire [4-1:0] node31920;
	wire [4-1:0] node31922;
	wire [4-1:0] node31923;
	wire [4-1:0] node31926;
	wire [4-1:0] node31929;
	wire [4-1:0] node31930;
	wire [4-1:0] node31931;
	wire [4-1:0] node31932;
	wire [4-1:0] node31933;
	wire [4-1:0] node31936;
	wire [4-1:0] node31939;
	wire [4-1:0] node31940;
	wire [4-1:0] node31943;
	wire [4-1:0] node31946;
	wire [4-1:0] node31947;
	wire [4-1:0] node31948;
	wire [4-1:0] node31951;
	wire [4-1:0] node31954;
	wire [4-1:0] node31955;
	wire [4-1:0] node31958;
	wire [4-1:0] node31961;
	wire [4-1:0] node31962;
	wire [4-1:0] node31963;
	wire [4-1:0] node31965;
	wire [4-1:0] node31968;
	wire [4-1:0] node31969;
	wire [4-1:0] node31972;
	wire [4-1:0] node31975;
	wire [4-1:0] node31976;
	wire [4-1:0] node31977;
	wire [4-1:0] node31980;
	wire [4-1:0] node31983;
	wire [4-1:0] node31984;
	wire [4-1:0] node31985;
	wire [4-1:0] node31988;
	wire [4-1:0] node31992;
	wire [4-1:0] node31993;
	wire [4-1:0] node31994;
	wire [4-1:0] node31995;
	wire [4-1:0] node31996;
	wire [4-1:0] node31997;
	wire [4-1:0] node31998;
	wire [4-1:0] node32001;
	wire [4-1:0] node32002;
	wire [4-1:0] node32006;
	wire [4-1:0] node32008;
	wire [4-1:0] node32011;
	wire [4-1:0] node32012;
	wire [4-1:0] node32013;
	wire [4-1:0] node32014;
	wire [4-1:0] node32017;
	wire [4-1:0] node32022;
	wire [4-1:0] node32023;
	wire [4-1:0] node32024;
	wire [4-1:0] node32025;
	wire [4-1:0] node32026;
	wire [4-1:0] node32030;
	wire [4-1:0] node32031;
	wire [4-1:0] node32035;
	wire [4-1:0] node32036;
	wire [4-1:0] node32037;
	wire [4-1:0] node32041;
	wire [4-1:0] node32042;
	wire [4-1:0] node32046;
	wire [4-1:0] node32047;
	wire [4-1:0] node32048;
	wire [4-1:0] node32049;
	wire [4-1:0] node32052;
	wire [4-1:0] node32055;
	wire [4-1:0] node32056;
	wire [4-1:0] node32059;
	wire [4-1:0] node32062;
	wire [4-1:0] node32063;
	wire [4-1:0] node32064;
	wire [4-1:0] node32067;
	wire [4-1:0] node32071;
	wire [4-1:0] node32072;
	wire [4-1:0] node32073;
	wire [4-1:0] node32074;
	wire [4-1:0] node32076;
	wire [4-1:0] node32079;
	wire [4-1:0] node32080;
	wire [4-1:0] node32081;
	wire [4-1:0] node32085;
	wire [4-1:0] node32086;
	wire [4-1:0] node32090;
	wire [4-1:0] node32091;
	wire [4-1:0] node32093;
	wire [4-1:0] node32094;
	wire [4-1:0] node32097;
	wire [4-1:0] node32100;
	wire [4-1:0] node32102;
	wire [4-1:0] node32105;
	wire [4-1:0] node32106;
	wire [4-1:0] node32107;
	wire [4-1:0] node32108;
	wire [4-1:0] node32112;
	wire [4-1:0] node32113;
	wire [4-1:0] node32117;
	wire [4-1:0] node32118;
	wire [4-1:0] node32119;
	wire [4-1:0] node32123;
	wire [4-1:0] node32124;
	wire [4-1:0] node32128;
	wire [4-1:0] node32129;
	wire [4-1:0] node32130;
	wire [4-1:0] node32131;
	wire [4-1:0] node32132;
	wire [4-1:0] node32134;
	wire [4-1:0] node32137;
	wire [4-1:0] node32139;
	wire [4-1:0] node32142;
	wire [4-1:0] node32143;
	wire [4-1:0] node32144;
	wire [4-1:0] node32145;
	wire [4-1:0] node32149;
	wire [4-1:0] node32152;
	wire [4-1:0] node32153;
	wire [4-1:0] node32156;
	wire [4-1:0] node32157;
	wire [4-1:0] node32161;
	wire [4-1:0] node32162;
	wire [4-1:0] node32163;
	wire [4-1:0] node32164;
	wire [4-1:0] node32165;
	wire [4-1:0] node32168;
	wire [4-1:0] node32171;
	wire [4-1:0] node32172;
	wire [4-1:0] node32175;
	wire [4-1:0] node32178;
	wire [4-1:0] node32180;
	wire [4-1:0] node32183;
	wire [4-1:0] node32184;
	wire [4-1:0] node32185;
	wire [4-1:0] node32186;
	wire [4-1:0] node32189;
	wire [4-1:0] node32192;
	wire [4-1:0] node32194;
	wire [4-1:0] node32197;
	wire [4-1:0] node32198;
	wire [4-1:0] node32201;
	wire [4-1:0] node32204;
	wire [4-1:0] node32205;
	wire [4-1:0] node32206;
	wire [4-1:0] node32207;
	wire [4-1:0] node32209;
	wire [4-1:0] node32210;
	wire [4-1:0] node32213;
	wire [4-1:0] node32216;
	wire [4-1:0] node32217;
	wire [4-1:0] node32220;
	wire [4-1:0] node32223;
	wire [4-1:0] node32224;
	wire [4-1:0] node32227;
	wire [4-1:0] node32228;
	wire [4-1:0] node32229;
	wire [4-1:0] node32234;
	wire [4-1:0] node32235;
	wire [4-1:0] node32236;
	wire [4-1:0] node32237;
	wire [4-1:0] node32238;
	wire [4-1:0] node32241;
	wire [4-1:0] node32244;
	wire [4-1:0] node32245;
	wire [4-1:0] node32248;
	wire [4-1:0] node32251;
	wire [4-1:0] node32253;
	wire [4-1:0] node32256;
	wire [4-1:0] node32257;
	wire [4-1:0] node32260;
	wire [4-1:0] node32263;
	wire [4-1:0] node32264;
	wire [4-1:0] node32265;
	wire [4-1:0] node32266;
	wire [4-1:0] node32267;
	wire [4-1:0] node32268;
	wire [4-1:0] node32269;
	wire [4-1:0] node32270;
	wire [4-1:0] node32271;
	wire [4-1:0] node32272;
	wire [4-1:0] node32276;
	wire [4-1:0] node32279;
	wire [4-1:0] node32280;
	wire [4-1:0] node32281;
	wire [4-1:0] node32286;
	wire [4-1:0] node32287;
	wire [4-1:0] node32288;
	wire [4-1:0] node32289;
	wire [4-1:0] node32293;
	wire [4-1:0] node32296;
	wire [4-1:0] node32297;
	wire [4-1:0] node32298;
	wire [4-1:0] node32303;
	wire [4-1:0] node32304;
	wire [4-1:0] node32305;
	wire [4-1:0] node32307;
	wire [4-1:0] node32309;
	wire [4-1:0] node32312;
	wire [4-1:0] node32313;
	wire [4-1:0] node32316;
	wire [4-1:0] node32319;
	wire [4-1:0] node32320;
	wire [4-1:0] node32321;
	wire [4-1:0] node32322;
	wire [4-1:0] node32327;
	wire [4-1:0] node32328;
	wire [4-1:0] node32331;
	wire [4-1:0] node32334;
	wire [4-1:0] node32335;
	wire [4-1:0] node32336;
	wire [4-1:0] node32337;
	wire [4-1:0] node32338;
	wire [4-1:0] node32339;
	wire [4-1:0] node32342;
	wire [4-1:0] node32345;
	wire [4-1:0] node32346;
	wire [4-1:0] node32349;
	wire [4-1:0] node32352;
	wire [4-1:0] node32353;
	wire [4-1:0] node32356;
	wire [4-1:0] node32359;
	wire [4-1:0] node32360;
	wire [4-1:0] node32362;
	wire [4-1:0] node32365;
	wire [4-1:0] node32366;
	wire [4-1:0] node32370;
	wire [4-1:0] node32371;
	wire [4-1:0] node32372;
	wire [4-1:0] node32373;
	wire [4-1:0] node32377;
	wire [4-1:0] node32378;
	wire [4-1:0] node32381;
	wire [4-1:0] node32384;
	wire [4-1:0] node32385;
	wire [4-1:0] node32386;
	wire [4-1:0] node32387;
	wire [4-1:0] node32391;
	wire [4-1:0] node32392;
	wire [4-1:0] node32396;
	wire [4-1:0] node32397;
	wire [4-1:0] node32398;
	wire [4-1:0] node32403;
	wire [4-1:0] node32404;
	wire [4-1:0] node32405;
	wire [4-1:0] node32406;
	wire [4-1:0] node32407;
	wire [4-1:0] node32408;
	wire [4-1:0] node32410;
	wire [4-1:0] node32413;
	wire [4-1:0] node32414;
	wire [4-1:0] node32417;
	wire [4-1:0] node32420;
	wire [4-1:0] node32421;
	wire [4-1:0] node32424;
	wire [4-1:0] node32425;
	wire [4-1:0] node32429;
	wire [4-1:0] node32430;
	wire [4-1:0] node32431;
	wire [4-1:0] node32433;
	wire [4-1:0] node32437;
	wire [4-1:0] node32439;
	wire [4-1:0] node32440;
	wire [4-1:0] node32443;
	wire [4-1:0] node32446;
	wire [4-1:0] node32447;
	wire [4-1:0] node32448;
	wire [4-1:0] node32449;
	wire [4-1:0] node32451;
	wire [4-1:0] node32455;
	wire [4-1:0] node32457;
	wire [4-1:0] node32458;
	wire [4-1:0] node32461;
	wire [4-1:0] node32464;
	wire [4-1:0] node32465;
	wire [4-1:0] node32466;
	wire [4-1:0] node32467;
	wire [4-1:0] node32470;
	wire [4-1:0] node32473;
	wire [4-1:0] node32474;
	wire [4-1:0] node32477;
	wire [4-1:0] node32480;
	wire [4-1:0] node32481;
	wire [4-1:0] node32482;
	wire [4-1:0] node32485;
	wire [4-1:0] node32489;
	wire [4-1:0] node32490;
	wire [4-1:0] node32491;
	wire [4-1:0] node32492;
	wire [4-1:0] node32494;
	wire [4-1:0] node32496;
	wire [4-1:0] node32499;
	wire [4-1:0] node32500;
	wire [4-1:0] node32503;
	wire [4-1:0] node32506;
	wire [4-1:0] node32507;
	wire [4-1:0] node32508;
	wire [4-1:0] node32509;
	wire [4-1:0] node32514;
	wire [4-1:0] node32516;
	wire [4-1:0] node32519;
	wire [4-1:0] node32520;
	wire [4-1:0] node32521;
	wire [4-1:0] node32522;
	wire [4-1:0] node32523;
	wire [4-1:0] node32527;
	wire [4-1:0] node32528;
	wire [4-1:0] node32532;
	wire [4-1:0] node32533;
	wire [4-1:0] node32537;
	wire [4-1:0] node32538;
	wire [4-1:0] node32539;
	wire [4-1:0] node32540;
	wire [4-1:0] node32543;
	wire [4-1:0] node32546;
	wire [4-1:0] node32547;
	wire [4-1:0] node32551;
	wire [4-1:0] node32552;
	wire [4-1:0] node32555;
	wire [4-1:0] node32558;
	wire [4-1:0] node32559;
	wire [4-1:0] node32560;
	wire [4-1:0] node32561;
	wire [4-1:0] node32562;
	wire [4-1:0] node32563;
	wire [4-1:0] node32564;
	wire [4-1:0] node32567;
	wire [4-1:0] node32569;
	wire [4-1:0] node32572;
	wire [4-1:0] node32573;
	wire [4-1:0] node32574;
	wire [4-1:0] node32577;
	wire [4-1:0] node32581;
	wire [4-1:0] node32582;
	wire [4-1:0] node32583;
	wire [4-1:0] node32584;
	wire [4-1:0] node32587;
	wire [4-1:0] node32591;
	wire [4-1:0] node32592;
	wire [4-1:0] node32595;
	wire [4-1:0] node32598;
	wire [4-1:0] node32599;
	wire [4-1:0] node32600;
	wire [4-1:0] node32602;
	wire [4-1:0] node32603;
	wire [4-1:0] node32606;
	wire [4-1:0] node32609;
	wire [4-1:0] node32610;
	wire [4-1:0] node32613;
	wire [4-1:0] node32616;
	wire [4-1:0] node32617;
	wire [4-1:0] node32618;
	wire [4-1:0] node32619;
	wire [4-1:0] node32622;
	wire [4-1:0] node32626;
	wire [4-1:0] node32627;
	wire [4-1:0] node32630;
	wire [4-1:0] node32633;
	wire [4-1:0] node32634;
	wire [4-1:0] node32635;
	wire [4-1:0] node32636;
	wire [4-1:0] node32637;
	wire [4-1:0] node32638;
	wire [4-1:0] node32642;
	wire [4-1:0] node32643;
	wire [4-1:0] node32646;
	wire [4-1:0] node32649;
	wire [4-1:0] node32650;
	wire [4-1:0] node32654;
	wire [4-1:0] node32655;
	wire [4-1:0] node32656;
	wire [4-1:0] node32657;
	wire [4-1:0] node32660;
	wire [4-1:0] node32663;
	wire [4-1:0] node32665;
	wire [4-1:0] node32668;
	wire [4-1:0] node32669;
	wire [4-1:0] node32672;
	wire [4-1:0] node32675;
	wire [4-1:0] node32676;
	wire [4-1:0] node32677;
	wire [4-1:0] node32678;
	wire [4-1:0] node32679;
	wire [4-1:0] node32682;
	wire [4-1:0] node32685;
	wire [4-1:0] node32686;
	wire [4-1:0] node32689;
	wire [4-1:0] node32692;
	wire [4-1:0] node32693;
	wire [4-1:0] node32696;
	wire [4-1:0] node32699;
	wire [4-1:0] node32700;
	wire [4-1:0] node32701;
	wire [4-1:0] node32702;
	wire [4-1:0] node32706;
	wire [4-1:0] node32709;
	wire [4-1:0] node32711;
	wire [4-1:0] node32714;
	wire [4-1:0] node32715;
	wire [4-1:0] node32716;
	wire [4-1:0] node32717;
	wire [4-1:0] node32718;
	wire [4-1:0] node32719;
	wire [4-1:0] node32721;
	wire [4-1:0] node32725;
	wire [4-1:0] node32726;
	wire [4-1:0] node32727;
	wire [4-1:0] node32730;
	wire [4-1:0] node32733;
	wire [4-1:0] node32734;
	wire [4-1:0] node32737;
	wire [4-1:0] node32740;
	wire [4-1:0] node32741;
	wire [4-1:0] node32743;
	wire [4-1:0] node32744;
	wire [4-1:0] node32747;
	wire [4-1:0] node32750;
	wire [4-1:0] node32751;
	wire [4-1:0] node32753;
	wire [4-1:0] node32756;
	wire [4-1:0] node32757;
	wire [4-1:0] node32760;
	wire [4-1:0] node32763;
	wire [4-1:0] node32764;
	wire [4-1:0] node32765;
	wire [4-1:0] node32766;
	wire [4-1:0] node32769;
	wire [4-1:0] node32772;
	wire [4-1:0] node32775;
	wire [4-1:0] node32776;
	wire [4-1:0] node32777;
	wire [4-1:0] node32780;
	wire [4-1:0] node32783;
	wire [4-1:0] node32785;
	wire [4-1:0] node32786;
	wire [4-1:0] node32789;
	wire [4-1:0] node32792;
	wire [4-1:0] node32793;
	wire [4-1:0] node32794;
	wire [4-1:0] node32795;
	wire [4-1:0] node32797;
	wire [4-1:0] node32798;
	wire [4-1:0] node32801;
	wire [4-1:0] node32804;
	wire [4-1:0] node32805;
	wire [4-1:0] node32806;
	wire [4-1:0] node32810;
	wire [4-1:0] node32811;
	wire [4-1:0] node32815;
	wire [4-1:0] node32816;
	wire [4-1:0] node32817;
	wire [4-1:0] node32818;
	wire [4-1:0] node32822;
	wire [4-1:0] node32823;
	wire [4-1:0] node32826;
	wire [4-1:0] node32830;
	wire [4-1:0] node32831;
	wire [4-1:0] node32832;
	wire [4-1:0] node32833;
	wire [4-1:0] node32835;
	wire [4-1:0] node32839;
	wire [4-1:0] node32840;
	wire [4-1:0] node32841;
	wire [4-1:0] node32844;
	wire [4-1:0] node32847;
	wire [4-1:0] node32848;
	wire [4-1:0] node32852;
	wire [4-1:0] node32854;
	wire [4-1:0] node32855;
	wire [4-1:0] node32858;
	wire [4-1:0] node32861;
	wire [4-1:0] node32862;
	wire [4-1:0] node32863;
	wire [4-1:0] node32864;
	wire [4-1:0] node32865;
	wire [4-1:0] node32866;
	wire [4-1:0] node32867;
	wire [4-1:0] node32868;
	wire [4-1:0] node32869;
	wire [4-1:0] node32873;
	wire [4-1:0] node32874;
	wire [4-1:0] node32877;
	wire [4-1:0] node32880;
	wire [4-1:0] node32881;
	wire [4-1:0] node32884;
	wire [4-1:0] node32887;
	wire [4-1:0] node32888;
	wire [4-1:0] node32889;
	wire [4-1:0] node32890;
	wire [4-1:0] node32894;
	wire [4-1:0] node32896;
	wire [4-1:0] node32899;
	wire [4-1:0] node32900;
	wire [4-1:0] node32903;
	wire [4-1:0] node32906;
	wire [4-1:0] node32907;
	wire [4-1:0] node32908;
	wire [4-1:0] node32910;
	wire [4-1:0] node32911;
	wire [4-1:0] node32914;
	wire [4-1:0] node32917;
	wire [4-1:0] node32918;
	wire [4-1:0] node32921;
	wire [4-1:0] node32924;
	wire [4-1:0] node32925;
	wire [4-1:0] node32926;
	wire [4-1:0] node32927;
	wire [4-1:0] node32930;
	wire [4-1:0] node32934;
	wire [4-1:0] node32935;
	wire [4-1:0] node32938;
	wire [4-1:0] node32941;
	wire [4-1:0] node32942;
	wire [4-1:0] node32943;
	wire [4-1:0] node32944;
	wire [4-1:0] node32946;
	wire [4-1:0] node32947;
	wire [4-1:0] node32950;
	wire [4-1:0] node32953;
	wire [4-1:0] node32955;
	wire [4-1:0] node32958;
	wire [4-1:0] node32959;
	wire [4-1:0] node32961;
	wire [4-1:0] node32962;
	wire [4-1:0] node32966;
	wire [4-1:0] node32967;
	wire [4-1:0] node32968;
	wire [4-1:0] node32973;
	wire [4-1:0] node32974;
	wire [4-1:0] node32975;
	wire [4-1:0] node32976;
	wire [4-1:0] node32977;
	wire [4-1:0] node32981;
	wire [4-1:0] node32982;
	wire [4-1:0] node32985;
	wire [4-1:0] node32988;
	wire [4-1:0] node32990;
	wire [4-1:0] node32991;
	wire [4-1:0] node32994;
	wire [4-1:0] node32997;
	wire [4-1:0] node32998;
	wire [4-1:0] node32999;
	wire [4-1:0] node33000;
	wire [4-1:0] node33003;
	wire [4-1:0] node33006;
	wire [4-1:0] node33007;
	wire [4-1:0] node33011;
	wire [4-1:0] node33012;
	wire [4-1:0] node33013;
	wire [4-1:0] node33017;
	wire [4-1:0] node33019;
	wire [4-1:0] node33022;
	wire [4-1:0] node33023;
	wire [4-1:0] node33024;
	wire [4-1:0] node33025;
	wire [4-1:0] node33026;
	wire [4-1:0] node33028;
	wire [4-1:0] node33029;
	wire [4-1:0] node33034;
	wire [4-1:0] node33035;
	wire [4-1:0] node33036;
	wire [4-1:0] node33037;
	wire [4-1:0] node33040;
	wire [4-1:0] node33044;
	wire [4-1:0] node33045;
	wire [4-1:0] node33048;
	wire [4-1:0] node33051;
	wire [4-1:0] node33052;
	wire [4-1:0] node33053;
	wire [4-1:0] node33054;
	wire [4-1:0] node33058;
	wire [4-1:0] node33059;
	wire [4-1:0] node33063;
	wire [4-1:0] node33064;
	wire [4-1:0] node33065;
	wire [4-1:0] node33069;
	wire [4-1:0] node33072;
	wire [4-1:0] node33073;
	wire [4-1:0] node33074;
	wire [4-1:0] node33075;
	wire [4-1:0] node33076;
	wire [4-1:0] node33078;
	wire [4-1:0] node33081;
	wire [4-1:0] node33082;
	wire [4-1:0] node33085;
	wire [4-1:0] node33089;
	wire [4-1:0] node33090;
	wire [4-1:0] node33091;
	wire [4-1:0] node33094;
	wire [4-1:0] node33097;
	wire [4-1:0] node33098;
	wire [4-1:0] node33101;
	wire [4-1:0] node33104;
	wire [4-1:0] node33105;
	wire [4-1:0] node33106;
	wire [4-1:0] node33107;
	wire [4-1:0] node33111;
	wire [4-1:0] node33112;
	wire [4-1:0] node33114;
	wire [4-1:0] node33117;
	wire [4-1:0] node33118;
	wire [4-1:0] node33122;
	wire [4-1:0] node33123;
	wire [4-1:0] node33126;
	wire [4-1:0] node33129;
	wire [4-1:0] node33130;
	wire [4-1:0] node33131;
	wire [4-1:0] node33132;
	wire [4-1:0] node33133;
	wire [4-1:0] node33134;
	wire [4-1:0] node33135;
	wire [4-1:0] node33136;
	wire [4-1:0] node33140;
	wire [4-1:0] node33141;
	wire [4-1:0] node33144;
	wire [4-1:0] node33147;
	wire [4-1:0] node33148;
	wire [4-1:0] node33149;
	wire [4-1:0] node33152;
	wire [4-1:0] node33156;
	wire [4-1:0] node33157;
	wire [4-1:0] node33159;
	wire [4-1:0] node33162;
	wire [4-1:0] node33163;
	wire [4-1:0] node33166;
	wire [4-1:0] node33169;
	wire [4-1:0] node33170;
	wire [4-1:0] node33171;
	wire [4-1:0] node33172;
	wire [4-1:0] node33173;
	wire [4-1:0] node33177;
	wire [4-1:0] node33178;
	wire [4-1:0] node33182;
	wire [4-1:0] node33183;
	wire [4-1:0] node33184;
	wire [4-1:0] node33188;
	wire [4-1:0] node33189;
	wire [4-1:0] node33193;
	wire [4-1:0] node33194;
	wire [4-1:0] node33195;
	wire [4-1:0] node33196;
	wire [4-1:0] node33199;
	wire [4-1:0] node33202;
	wire [4-1:0] node33204;
	wire [4-1:0] node33207;
	wire [4-1:0] node33208;
	wire [4-1:0] node33212;
	wire [4-1:0] node33213;
	wire [4-1:0] node33214;
	wire [4-1:0] node33215;
	wire [4-1:0] node33216;
	wire [4-1:0] node33217;
	wire [4-1:0] node33221;
	wire [4-1:0] node33223;
	wire [4-1:0] node33226;
	wire [4-1:0] node33227;
	wire [4-1:0] node33228;
	wire [4-1:0] node33231;
	wire [4-1:0] node33234;
	wire [4-1:0] node33235;
	wire [4-1:0] node33238;
	wire [4-1:0] node33241;
	wire [4-1:0] node33242;
	wire [4-1:0] node33243;
	wire [4-1:0] node33244;
	wire [4-1:0] node33247;
	wire [4-1:0] node33250;
	wire [4-1:0] node33251;
	wire [4-1:0] node33254;
	wire [4-1:0] node33257;
	wire [4-1:0] node33258;
	wire [4-1:0] node33259;
	wire [4-1:0] node33262;
	wire [4-1:0] node33265;
	wire [4-1:0] node33266;
	wire [4-1:0] node33269;
	wire [4-1:0] node33272;
	wire [4-1:0] node33273;
	wire [4-1:0] node33274;
	wire [4-1:0] node33275;
	wire [4-1:0] node33277;
	wire [4-1:0] node33281;
	wire [4-1:0] node33282;
	wire [4-1:0] node33283;
	wire [4-1:0] node33287;
	wire [4-1:0] node33288;
	wire [4-1:0] node33291;
	wire [4-1:0] node33294;
	wire [4-1:0] node33295;
	wire [4-1:0] node33296;
	wire [4-1:0] node33298;
	wire [4-1:0] node33302;
	wire [4-1:0] node33303;
	wire [4-1:0] node33306;
	wire [4-1:0] node33307;
	wire [4-1:0] node33310;
	wire [4-1:0] node33313;
	wire [4-1:0] node33314;
	wire [4-1:0] node33315;
	wire [4-1:0] node33316;
	wire [4-1:0] node33317;
	wire [4-1:0] node33319;
	wire [4-1:0] node33320;
	wire [4-1:0] node33323;
	wire [4-1:0] node33326;
	wire [4-1:0] node33327;
	wire [4-1:0] node33330;
	wire [4-1:0] node33333;
	wire [4-1:0] node33334;
	wire [4-1:0] node33335;
	wire [4-1:0] node33336;
	wire [4-1:0] node33339;
	wire [4-1:0] node33342;
	wire [4-1:0] node33343;
	wire [4-1:0] node33346;
	wire [4-1:0] node33349;
	wire [4-1:0] node33350;
	wire [4-1:0] node33353;
	wire [4-1:0] node33355;
	wire [4-1:0] node33358;
	wire [4-1:0] node33359;
	wire [4-1:0] node33360;
	wire [4-1:0] node33362;
	wire [4-1:0] node33363;
	wire [4-1:0] node33366;
	wire [4-1:0] node33369;
	wire [4-1:0] node33370;
	wire [4-1:0] node33373;
	wire [4-1:0] node33376;
	wire [4-1:0] node33378;
	wire [4-1:0] node33379;
	wire [4-1:0] node33382;
	wire [4-1:0] node33385;
	wire [4-1:0] node33386;
	wire [4-1:0] node33387;
	wire [4-1:0] node33388;
	wire [4-1:0] node33389;
	wire [4-1:0] node33392;
	wire [4-1:0] node33395;
	wire [4-1:0] node33396;
	wire [4-1:0] node33399;
	wire [4-1:0] node33402;
	wire [4-1:0] node33403;
	wire [4-1:0] node33406;
	wire [4-1:0] node33409;
	wire [4-1:0] node33410;
	wire [4-1:0] node33411;
	wire [4-1:0] node33412;
	wire [4-1:0] node33413;
	wire [4-1:0] node33417;
	wire [4-1:0] node33419;
	wire [4-1:0] node33423;
	wire [4-1:0] node33424;
	wire [4-1:0] node33427;
	wire [4-1:0] node33430;
	wire [4-1:0] node33431;
	wire [4-1:0] node33432;
	wire [4-1:0] node33433;
	wire [4-1:0] node33434;
	wire [4-1:0] node33435;
	wire [4-1:0] node33436;
	wire [4-1:0] node33437;
	wire [4-1:0] node33438;
	wire [4-1:0] node33439;
	wire [4-1:0] node33440;
	wire [4-1:0] node33441;
	wire [4-1:0] node33442;
	wire [4-1:0] node33445;
	wire [4-1:0] node33447;
	wire [4-1:0] node33450;
	wire [4-1:0] node33451;
	wire [4-1:0] node33452;
	wire [4-1:0] node33456;
	wire [4-1:0] node33457;
	wire [4-1:0] node33459;
	wire [4-1:0] node33463;
	wire [4-1:0] node33464;
	wire [4-1:0] node33465;
	wire [4-1:0] node33466;
	wire [4-1:0] node33467;
	wire [4-1:0] node33470;
	wire [4-1:0] node33474;
	wire [4-1:0] node33475;
	wire [4-1:0] node33478;
	wire [4-1:0] node33481;
	wire [4-1:0] node33482;
	wire [4-1:0] node33483;
	wire [4-1:0] node33487;
	wire [4-1:0] node33488;
	wire [4-1:0] node33489;
	wire [4-1:0] node33492;
	wire [4-1:0] node33495;
	wire [4-1:0] node33497;
	wire [4-1:0] node33500;
	wire [4-1:0] node33501;
	wire [4-1:0] node33502;
	wire [4-1:0] node33503;
	wire [4-1:0] node33504;
	wire [4-1:0] node33507;
	wire [4-1:0] node33510;
	wire [4-1:0] node33512;
	wire [4-1:0] node33513;
	wire [4-1:0] node33516;
	wire [4-1:0] node33519;
	wire [4-1:0] node33520;
	wire [4-1:0] node33521;
	wire [4-1:0] node33524;
	wire [4-1:0] node33527;
	wire [4-1:0] node33528;
	wire [4-1:0] node33531;
	wire [4-1:0] node33534;
	wire [4-1:0] node33535;
	wire [4-1:0] node33536;
	wire [4-1:0] node33539;
	wire [4-1:0] node33541;
	wire [4-1:0] node33544;
	wire [4-1:0] node33545;
	wire [4-1:0] node33546;
	wire [4-1:0] node33547;
	wire [4-1:0] node33551;
	wire [4-1:0] node33554;
	wire [4-1:0] node33555;
	wire [4-1:0] node33556;
	wire [4-1:0] node33559;
	wire [4-1:0] node33562;
	wire [4-1:0] node33563;
	wire [4-1:0] node33567;
	wire [4-1:0] node33568;
	wire [4-1:0] node33569;
	wire [4-1:0] node33570;
	wire [4-1:0] node33571;
	wire [4-1:0] node33572;
	wire [4-1:0] node33575;
	wire [4-1:0] node33578;
	wire [4-1:0] node33579;
	wire [4-1:0] node33582;
	wire [4-1:0] node33585;
	wire [4-1:0] node33586;
	wire [4-1:0] node33589;
	wire [4-1:0] node33591;
	wire [4-1:0] node33594;
	wire [4-1:0] node33595;
	wire [4-1:0] node33596;
	wire [4-1:0] node33597;
	wire [4-1:0] node33600;
	wire [4-1:0] node33603;
	wire [4-1:0] node33604;
	wire [4-1:0] node33606;
	wire [4-1:0] node33609;
	wire [4-1:0] node33610;
	wire [4-1:0] node33614;
	wire [4-1:0] node33615;
	wire [4-1:0] node33618;
	wire [4-1:0] node33621;
	wire [4-1:0] node33622;
	wire [4-1:0] node33623;
	wire [4-1:0] node33624;
	wire [4-1:0] node33625;
	wire [4-1:0] node33626;
	wire [4-1:0] node33630;
	wire [4-1:0] node33631;
	wire [4-1:0] node33635;
	wire [4-1:0] node33636;
	wire [4-1:0] node33637;
	wire [4-1:0] node33640;
	wire [4-1:0] node33643;
	wire [4-1:0] node33644;
	wire [4-1:0] node33647;
	wire [4-1:0] node33650;
	wire [4-1:0] node33651;
	wire [4-1:0] node33654;
	wire [4-1:0] node33655;
	wire [4-1:0] node33656;
	wire [4-1:0] node33660;
	wire [4-1:0] node33662;
	wire [4-1:0] node33665;
	wire [4-1:0] node33666;
	wire [4-1:0] node33667;
	wire [4-1:0] node33668;
	wire [4-1:0] node33671;
	wire [4-1:0] node33672;
	wire [4-1:0] node33675;
	wire [4-1:0] node33678;
	wire [4-1:0] node33679;
	wire [4-1:0] node33681;
	wire [4-1:0] node33684;
	wire [4-1:0] node33687;
	wire [4-1:0] node33688;
	wire [4-1:0] node33690;
	wire [4-1:0] node33691;
	wire [4-1:0] node33695;
	wire [4-1:0] node33696;
	wire [4-1:0] node33698;
	wire [4-1:0] node33702;
	wire [4-1:0] node33703;
	wire [4-1:0] node33704;
	wire [4-1:0] node33705;
	wire [4-1:0] node33706;
	wire [4-1:0] node33709;
	wire [4-1:0] node33711;
	wire [4-1:0] node33714;
	wire [4-1:0] node33715;
	wire [4-1:0] node33716;
	wire [4-1:0] node33719;
	wire [4-1:0] node33722;
	wire [4-1:0] node33723;
	wire [4-1:0] node33724;
	wire [4-1:0] node33725;
	wire [4-1:0] node33728;
	wire [4-1:0] node33731;
	wire [4-1:0] node33732;
	wire [4-1:0] node33736;
	wire [4-1:0] node33737;
	wire [4-1:0] node33739;
	wire [4-1:0] node33742;
	wire [4-1:0] node33743;
	wire [4-1:0] node33746;
	wire [4-1:0] node33749;
	wire [4-1:0] node33750;
	wire [4-1:0] node33751;
	wire [4-1:0] node33754;
	wire [4-1:0] node33756;
	wire [4-1:0] node33759;
	wire [4-1:0] node33760;
	wire [4-1:0] node33761;
	wire [4-1:0] node33764;
	wire [4-1:0] node33767;
	wire [4-1:0] node33768;
	wire [4-1:0] node33769;
	wire [4-1:0] node33773;
	wire [4-1:0] node33774;
	wire [4-1:0] node33777;
	wire [4-1:0] node33780;
	wire [4-1:0] node33781;
	wire [4-1:0] node33782;
	wire [4-1:0] node33783;
	wire [4-1:0] node33784;
	wire [4-1:0] node33787;
	wire [4-1:0] node33790;
	wire [4-1:0] node33791;
	wire [4-1:0] node33794;
	wire [4-1:0] node33797;
	wire [4-1:0] node33798;
	wire [4-1:0] node33799;
	wire [4-1:0] node33802;
	wire [4-1:0] node33805;
	wire [4-1:0] node33806;
	wire [4-1:0] node33807;
	wire [4-1:0] node33812;
	wire [4-1:0] node33813;
	wire [4-1:0] node33814;
	wire [4-1:0] node33817;
	wire [4-1:0] node33819;
	wire [4-1:0] node33822;
	wire [4-1:0] node33823;
	wire [4-1:0] node33824;
	wire [4-1:0] node33827;
	wire [4-1:0] node33830;
	wire [4-1:0] node33831;
	wire [4-1:0] node33834;
	wire [4-1:0] node33837;
	wire [4-1:0] node33838;
	wire [4-1:0] node33839;
	wire [4-1:0] node33840;
	wire [4-1:0] node33841;
	wire [4-1:0] node33842;
	wire [4-1:0] node33843;
	wire [4-1:0] node33846;
	wire [4-1:0] node33849;
	wire [4-1:0] node33850;
	wire [4-1:0] node33851;
	wire [4-1:0] node33855;
	wire [4-1:0] node33856;
	wire [4-1:0] node33859;
	wire [4-1:0] node33862;
	wire [4-1:0] node33863;
	wire [4-1:0] node33864;
	wire [4-1:0] node33867;
	wire [4-1:0] node33869;
	wire [4-1:0] node33872;
	wire [4-1:0] node33873;
	wire [4-1:0] node33874;
	wire [4-1:0] node33878;
	wire [4-1:0] node33879;
	wire [4-1:0] node33882;
	wire [4-1:0] node33885;
	wire [4-1:0] node33886;
	wire [4-1:0] node33887;
	wire [4-1:0] node33888;
	wire [4-1:0] node33889;
	wire [4-1:0] node33892;
	wire [4-1:0] node33895;
	wire [4-1:0] node33896;
	wire [4-1:0] node33899;
	wire [4-1:0] node33902;
	wire [4-1:0] node33903;
	wire [4-1:0] node33904;
	wire [4-1:0] node33907;
	wire [4-1:0] node33910;
	wire [4-1:0] node33911;
	wire [4-1:0] node33913;
	wire [4-1:0] node33916;
	wire [4-1:0] node33917;
	wire [4-1:0] node33921;
	wire [4-1:0] node33922;
	wire [4-1:0] node33923;
	wire [4-1:0] node33926;
	wire [4-1:0] node33928;
	wire [4-1:0] node33931;
	wire [4-1:0] node33932;
	wire [4-1:0] node33933;
	wire [4-1:0] node33936;
	wire [4-1:0] node33939;
	wire [4-1:0] node33940;
	wire [4-1:0] node33943;
	wire [4-1:0] node33946;
	wire [4-1:0] node33947;
	wire [4-1:0] node33948;
	wire [4-1:0] node33949;
	wire [4-1:0] node33950;
	wire [4-1:0] node33953;
	wire [4-1:0] node33955;
	wire [4-1:0] node33958;
	wire [4-1:0] node33959;
	wire [4-1:0] node33962;
	wire [4-1:0] node33964;
	wire [4-1:0] node33967;
	wire [4-1:0] node33968;
	wire [4-1:0] node33969;
	wire [4-1:0] node33972;
	wire [4-1:0] node33973;
	wire [4-1:0] node33977;
	wire [4-1:0] node33978;
	wire [4-1:0] node33981;
	wire [4-1:0] node33983;
	wire [4-1:0] node33986;
	wire [4-1:0] node33987;
	wire [4-1:0] node33988;
	wire [4-1:0] node33989;
	wire [4-1:0] node33991;
	wire [4-1:0] node33992;
	wire [4-1:0] node33996;
	wire [4-1:0] node33997;
	wire [4-1:0] node34001;
	wire [4-1:0] node34002;
	wire [4-1:0] node34003;
	wire [4-1:0] node34006;
	wire [4-1:0] node34009;
	wire [4-1:0] node34010;
	wire [4-1:0] node34011;
	wire [4-1:0] node34014;
	wire [4-1:0] node34017;
	wire [4-1:0] node34018;
	wire [4-1:0] node34021;
	wire [4-1:0] node34024;
	wire [4-1:0] node34025;
	wire [4-1:0] node34026;
	wire [4-1:0] node34027;
	wire [4-1:0] node34031;
	wire [4-1:0] node34032;
	wire [4-1:0] node34033;
	wire [4-1:0] node34036;
	wire [4-1:0] node34039;
	wire [4-1:0] node34040;
	wire [4-1:0] node34044;
	wire [4-1:0] node34045;
	wire [4-1:0] node34046;
	wire [4-1:0] node34049;
	wire [4-1:0] node34052;
	wire [4-1:0] node34053;
	wire [4-1:0] node34056;
	wire [4-1:0] node34059;
	wire [4-1:0] node34060;
	wire [4-1:0] node34061;
	wire [4-1:0] node34062;
	wire [4-1:0] node34063;
	wire [4-1:0] node34066;
	wire [4-1:0] node34068;
	wire [4-1:0] node34071;
	wire [4-1:0] node34072;
	wire [4-1:0] node34073;
	wire [4-1:0] node34076;
	wire [4-1:0] node34079;
	wire [4-1:0] node34080;
	wire [4-1:0] node34083;
	wire [4-1:0] node34086;
	wire [4-1:0] node34087;
	wire [4-1:0] node34088;
	wire [4-1:0] node34091;
	wire [4-1:0] node34093;
	wire [4-1:0] node34096;
	wire [4-1:0] node34097;
	wire [4-1:0] node34098;
	wire [4-1:0] node34101;
	wire [4-1:0] node34104;
	wire [4-1:0] node34105;
	wire [4-1:0] node34106;
	wire [4-1:0] node34109;
	wire [4-1:0] node34112;
	wire [4-1:0] node34113;
	wire [4-1:0] node34117;
	wire [4-1:0] node34118;
	wire [4-1:0] node34119;
	wire [4-1:0] node34120;
	wire [4-1:0] node34123;
	wire [4-1:0] node34125;
	wire [4-1:0] node34128;
	wire [4-1:0] node34129;
	wire [4-1:0] node34130;
	wire [4-1:0] node34133;
	wire [4-1:0] node34136;
	wire [4-1:0] node34137;
	wire [4-1:0] node34138;
	wire [4-1:0] node34141;
	wire [4-1:0] node34144;
	wire [4-1:0] node34146;
	wire [4-1:0] node34147;
	wire [4-1:0] node34151;
	wire [4-1:0] node34152;
	wire [4-1:0] node34153;
	wire [4-1:0] node34156;
	wire [4-1:0] node34158;
	wire [4-1:0] node34161;
	wire [4-1:0] node34162;
	wire [4-1:0] node34163;
	wire [4-1:0] node34166;
	wire [4-1:0] node34169;
	wire [4-1:0] node34170;
	wire [4-1:0] node34173;
	wire [4-1:0] node34176;
	wire [4-1:0] node34177;
	wire [4-1:0] node34178;
	wire [4-1:0] node34179;
	wire [4-1:0] node34180;
	wire [4-1:0] node34181;
	wire [4-1:0] node34182;
	wire [4-1:0] node34183;
	wire [4-1:0] node34184;
	wire [4-1:0] node34188;
	wire [4-1:0] node34189;
	wire [4-1:0] node34192;
	wire [4-1:0] node34195;
	wire [4-1:0] node34196;
	wire [4-1:0] node34198;
	wire [4-1:0] node34201;
	wire [4-1:0] node34202;
	wire [4-1:0] node34203;
	wire [4-1:0] node34207;
	wire [4-1:0] node34208;
	wire [4-1:0] node34211;
	wire [4-1:0] node34214;
	wire [4-1:0] node34215;
	wire [4-1:0] node34216;
	wire [4-1:0] node34219;
	wire [4-1:0] node34221;
	wire [4-1:0] node34224;
	wire [4-1:0] node34225;
	wire [4-1:0] node34226;
	wire [4-1:0] node34229;
	wire [4-1:0] node34232;
	wire [4-1:0] node34234;
	wire [4-1:0] node34237;
	wire [4-1:0] node34238;
	wire [4-1:0] node34239;
	wire [4-1:0] node34240;
	wire [4-1:0] node34242;
	wire [4-1:0] node34246;
	wire [4-1:0] node34247;
	wire [4-1:0] node34249;
	wire [4-1:0] node34253;
	wire [4-1:0] node34254;
	wire [4-1:0] node34255;
	wire [4-1:0] node34258;
	wire [4-1:0] node34260;
	wire [4-1:0] node34263;
	wire [4-1:0] node34264;
	wire [4-1:0] node34265;
	wire [4-1:0] node34268;
	wire [4-1:0] node34272;
	wire [4-1:0] node34273;
	wire [4-1:0] node34274;
	wire [4-1:0] node34275;
	wire [4-1:0] node34276;
	wire [4-1:0] node34277;
	wire [4-1:0] node34280;
	wire [4-1:0] node34283;
	wire [4-1:0] node34284;
	wire [4-1:0] node34287;
	wire [4-1:0] node34290;
	wire [4-1:0] node34291;
	wire [4-1:0] node34292;
	wire [4-1:0] node34293;
	wire [4-1:0] node34296;
	wire [4-1:0] node34299;
	wire [4-1:0] node34300;
	wire [4-1:0] node34303;
	wire [4-1:0] node34306;
	wire [4-1:0] node34307;
	wire [4-1:0] node34311;
	wire [4-1:0] node34312;
	wire [4-1:0] node34313;
	wire [4-1:0] node34314;
	wire [4-1:0] node34317;
	wire [4-1:0] node34320;
	wire [4-1:0] node34321;
	wire [4-1:0] node34323;
	wire [4-1:0] node34327;
	wire [4-1:0] node34328;
	wire [4-1:0] node34330;
	wire [4-1:0] node34332;
	wire [4-1:0] node34335;
	wire [4-1:0] node34336;
	wire [4-1:0] node34337;
	wire [4-1:0] node34341;
	wire [4-1:0] node34342;
	wire [4-1:0] node34346;
	wire [4-1:0] node34347;
	wire [4-1:0] node34348;
	wire [4-1:0] node34349;
	wire [4-1:0] node34350;
	wire [4-1:0] node34351;
	wire [4-1:0] node34355;
	wire [4-1:0] node34357;
	wire [4-1:0] node34360;
	wire [4-1:0] node34361;
	wire [4-1:0] node34362;
	wire [4-1:0] node34366;
	wire [4-1:0] node34367;
	wire [4-1:0] node34371;
	wire [4-1:0] node34372;
	wire [4-1:0] node34373;
	wire [4-1:0] node34374;
	wire [4-1:0] node34377;
	wire [4-1:0] node34381;
	wire [4-1:0] node34382;
	wire [4-1:0] node34385;
	wire [4-1:0] node34388;
	wire [4-1:0] node34389;
	wire [4-1:0] node34390;
	wire [4-1:0] node34392;
	wire [4-1:0] node34393;
	wire [4-1:0] node34397;
	wire [4-1:0] node34399;
	wire [4-1:0] node34401;
	wire [4-1:0] node34404;
	wire [4-1:0] node34405;
	wire [4-1:0] node34406;
	wire [4-1:0] node34407;
	wire [4-1:0] node34412;
	wire [4-1:0] node34413;
	wire [4-1:0] node34416;
	wire [4-1:0] node34419;
	wire [4-1:0] node34420;
	wire [4-1:0] node34421;
	wire [4-1:0] node34422;
	wire [4-1:0] node34423;
	wire [4-1:0] node34424;
	wire [4-1:0] node34425;
	wire [4-1:0] node34428;
	wire [4-1:0] node34431;
	wire [4-1:0] node34433;
	wire [4-1:0] node34434;
	wire [4-1:0] node34437;
	wire [4-1:0] node34440;
	wire [4-1:0] node34441;
	wire [4-1:0] node34442;
	wire [4-1:0] node34445;
	wire [4-1:0] node34448;
	wire [4-1:0] node34450;
	wire [4-1:0] node34453;
	wire [4-1:0] node34454;
	wire [4-1:0] node34457;
	wire [4-1:0] node34460;
	wire [4-1:0] node34461;
	wire [4-1:0] node34462;
	wire [4-1:0] node34463;
	wire [4-1:0] node34464;
	wire [4-1:0] node34465;
	wire [4-1:0] node34468;
	wire [4-1:0] node34471;
	wire [4-1:0] node34472;
	wire [4-1:0] node34475;
	wire [4-1:0] node34478;
	wire [4-1:0] node34479;
	wire [4-1:0] node34480;
	wire [4-1:0] node34484;
	wire [4-1:0] node34486;
	wire [4-1:0] node34489;
	wire [4-1:0] node34490;
	wire [4-1:0] node34493;
	wire [4-1:0] node34496;
	wire [4-1:0] node34497;
	wire [4-1:0] node34498;
	wire [4-1:0] node34500;
	wire [4-1:0] node34503;
	wire [4-1:0] node34504;
	wire [4-1:0] node34507;
	wire [4-1:0] node34510;
	wire [4-1:0] node34511;
	wire [4-1:0] node34512;
	wire [4-1:0] node34513;
	wire [4-1:0] node34516;
	wire [4-1:0] node34519;
	wire [4-1:0] node34520;
	wire [4-1:0] node34523;
	wire [4-1:0] node34526;
	wire [4-1:0] node34527;
	wire [4-1:0] node34530;
	wire [4-1:0] node34533;
	wire [4-1:0] node34534;
	wire [4-1:0] node34535;
	wire [4-1:0] node34536;
	wire [4-1:0] node34537;
	wire [4-1:0] node34538;
	wire [4-1:0] node34539;
	wire [4-1:0] node34543;
	wire [4-1:0] node34544;
	wire [4-1:0] node34547;
	wire [4-1:0] node34550;
	wire [4-1:0] node34551;
	wire [4-1:0] node34552;
	wire [4-1:0] node34555;
	wire [4-1:0] node34558;
	wire [4-1:0] node34559;
	wire [4-1:0] node34562;
	wire [4-1:0] node34565;
	wire [4-1:0] node34566;
	wire [4-1:0] node34567;
	wire [4-1:0] node34568;
	wire [4-1:0] node34571;
	wire [4-1:0] node34574;
	wire [4-1:0] node34576;
	wire [4-1:0] node34579;
	wire [4-1:0] node34580;
	wire [4-1:0] node34581;
	wire [4-1:0] node34584;
	wire [4-1:0] node34588;
	wire [4-1:0] node34589;
	wire [4-1:0] node34590;
	wire [4-1:0] node34591;
	wire [4-1:0] node34592;
	wire [4-1:0] node34595;
	wire [4-1:0] node34598;
	wire [4-1:0] node34601;
	wire [4-1:0] node34602;
	wire [4-1:0] node34603;
	wire [4-1:0] node34608;
	wire [4-1:0] node34609;
	wire [4-1:0] node34610;
	wire [4-1:0] node34611;
	wire [4-1:0] node34614;
	wire [4-1:0] node34617;
	wire [4-1:0] node34619;
	wire [4-1:0] node34622;
	wire [4-1:0] node34623;
	wire [4-1:0] node34624;
	wire [4-1:0] node34627;
	wire [4-1:0] node34630;
	wire [4-1:0] node34631;
	wire [4-1:0] node34634;
	wire [4-1:0] node34637;
	wire [4-1:0] node34638;
	wire [4-1:0] node34639;
	wire [4-1:0] node34640;
	wire [4-1:0] node34641;
	wire [4-1:0] node34642;
	wire [4-1:0] node34645;
	wire [4-1:0] node34648;
	wire [4-1:0] node34649;
	wire [4-1:0] node34652;
	wire [4-1:0] node34655;
	wire [4-1:0] node34656;
	wire [4-1:0] node34659;
	wire [4-1:0] node34662;
	wire [4-1:0] node34663;
	wire [4-1:0] node34664;
	wire [4-1:0] node34665;
	wire [4-1:0] node34669;
	wire [4-1:0] node34671;
	wire [4-1:0] node34674;
	wire [4-1:0] node34675;
	wire [4-1:0] node34678;
	wire [4-1:0] node34681;
	wire [4-1:0] node34682;
	wire [4-1:0] node34683;
	wire [4-1:0] node34684;
	wire [4-1:0] node34685;
	wire [4-1:0] node34689;
	wire [4-1:0] node34690;
	wire [4-1:0] node34693;
	wire [4-1:0] node34696;
	wire [4-1:0] node34698;
	wire [4-1:0] node34701;
	wire [4-1:0] node34702;
	wire [4-1:0] node34705;
	wire [4-1:0] node34708;
	wire [4-1:0] node34709;
	wire [4-1:0] node34710;
	wire [4-1:0] node34711;
	wire [4-1:0] node34712;
	wire [4-1:0] node34713;
	wire [4-1:0] node34714;
	wire [4-1:0] node34717;
	wire [4-1:0] node34719;
	wire [4-1:0] node34722;
	wire [4-1:0] node34723;
	wire [4-1:0] node34725;
	wire [4-1:0] node34728;
	wire [4-1:0] node34730;
	wire [4-1:0] node34733;
	wire [4-1:0] node34734;
	wire [4-1:0] node34735;
	wire [4-1:0] node34737;
	wire [4-1:0] node34740;
	wire [4-1:0] node34741;
	wire [4-1:0] node34744;
	wire [4-1:0] node34747;
	wire [4-1:0] node34748;
	wire [4-1:0] node34749;
	wire [4-1:0] node34752;
	wire [4-1:0] node34755;
	wire [4-1:0] node34756;
	wire [4-1:0] node34759;
	wire [4-1:0] node34762;
	wire [4-1:0] node34763;
	wire [4-1:0] node34764;
	wire [4-1:0] node34765;
	wire [4-1:0] node34767;
	wire [4-1:0] node34770;
	wire [4-1:0] node34772;
	wire [4-1:0] node34775;
	wire [4-1:0] node34776;
	wire [4-1:0] node34778;
	wire [4-1:0] node34781;
	wire [4-1:0] node34783;
	wire [4-1:0] node34786;
	wire [4-1:0] node34787;
	wire [4-1:0] node34788;
	wire [4-1:0] node34789;
	wire [4-1:0] node34793;
	wire [4-1:0] node34794;
	wire [4-1:0] node34798;
	wire [4-1:0] node34799;
	wire [4-1:0] node34800;
	wire [4-1:0] node34804;
	wire [4-1:0] node34805;
	wire [4-1:0] node34809;
	wire [4-1:0] node34810;
	wire [4-1:0] node34811;
	wire [4-1:0] node34812;
	wire [4-1:0] node34813;
	wire [4-1:0] node34816;
	wire [4-1:0] node34818;
	wire [4-1:0] node34821;
	wire [4-1:0] node34822;
	wire [4-1:0] node34823;
	wire [4-1:0] node34826;
	wire [4-1:0] node34829;
	wire [4-1:0] node34830;
	wire [4-1:0] node34834;
	wire [4-1:0] node34835;
	wire [4-1:0] node34836;
	wire [4-1:0] node34837;
	wire [4-1:0] node34840;
	wire [4-1:0] node34843;
	wire [4-1:0] node34845;
	wire [4-1:0] node34848;
	wire [4-1:0] node34849;
	wire [4-1:0] node34850;
	wire [4-1:0] node34853;
	wire [4-1:0] node34856;
	wire [4-1:0] node34857;
	wire [4-1:0] node34859;
	wire [4-1:0] node34863;
	wire [4-1:0] node34864;
	wire [4-1:0] node34865;
	wire [4-1:0] node34866;
	wire [4-1:0] node34868;
	wire [4-1:0] node34870;
	wire [4-1:0] node34873;
	wire [4-1:0] node34874;
	wire [4-1:0] node34877;
	wire [4-1:0] node34880;
	wire [4-1:0] node34881;
	wire [4-1:0] node34882;
	wire [4-1:0] node34885;
	wire [4-1:0] node34888;
	wire [4-1:0] node34889;
	wire [4-1:0] node34892;
	wire [4-1:0] node34895;
	wire [4-1:0] node34896;
	wire [4-1:0] node34897;
	wire [4-1:0] node34900;
	wire [4-1:0] node34903;
	wire [4-1:0] node34904;
	wire [4-1:0] node34905;
	wire [4-1:0] node34908;
	wire [4-1:0] node34911;
	wire [4-1:0] node34912;
	wire [4-1:0] node34916;
	wire [4-1:0] node34917;
	wire [4-1:0] node34918;
	wire [4-1:0] node34919;
	wire [4-1:0] node34920;
	wire [4-1:0] node34923;
	wire [4-1:0] node34926;
	wire [4-1:0] node34927;
	wire [4-1:0] node34928;
	wire [4-1:0] node34929;
	wire [4-1:0] node34932;
	wire [4-1:0] node34935;
	wire [4-1:0] node34936;
	wire [4-1:0] node34939;
	wire [4-1:0] node34942;
	wire [4-1:0] node34943;
	wire [4-1:0] node34944;
	wire [4-1:0] node34947;
	wire [4-1:0] node34950;
	wire [4-1:0] node34951;
	wire [4-1:0] node34955;
	wire [4-1:0] node34956;
	wire [4-1:0] node34957;
	wire [4-1:0] node34960;
	wire [4-1:0] node34963;
	wire [4-1:0] node34964;
	wire [4-1:0] node34965;
	wire [4-1:0] node34968;
	wire [4-1:0] node34971;
	wire [4-1:0] node34973;
	wire [4-1:0] node34974;
	wire [4-1:0] node34978;
	wire [4-1:0] node34979;
	wire [4-1:0] node34980;
	wire [4-1:0] node34981;
	wire [4-1:0] node34982;
	wire [4-1:0] node34984;
	wire [4-1:0] node34987;
	wire [4-1:0] node34988;
	wire [4-1:0] node34989;
	wire [4-1:0] node34992;
	wire [4-1:0] node34996;
	wire [4-1:0] node34997;
	wire [4-1:0] node34998;
	wire [4-1:0] node35001;
	wire [4-1:0] node35004;
	wire [4-1:0] node35007;
	wire [4-1:0] node35008;
	wire [4-1:0] node35009;
	wire [4-1:0] node35010;
	wire [4-1:0] node35014;
	wire [4-1:0] node35015;
	wire [4-1:0] node35017;
	wire [4-1:0] node35020;
	wire [4-1:0] node35021;
	wire [4-1:0] node35024;
	wire [4-1:0] node35027;
	wire [4-1:0] node35028;
	wire [4-1:0] node35029;
	wire [4-1:0] node35033;
	wire [4-1:0] node35035;
	wire [4-1:0] node35038;
	wire [4-1:0] node35039;
	wire [4-1:0] node35040;
	wire [4-1:0] node35041;
	wire [4-1:0] node35044;
	wire [4-1:0] node35047;
	wire [4-1:0] node35048;
	wire [4-1:0] node35051;
	wire [4-1:0] node35054;
	wire [4-1:0] node35055;
	wire [4-1:0] node35056;
	wire [4-1:0] node35059;
	wire [4-1:0] node35062;
	wire [4-1:0] node35063;
	wire [4-1:0] node35064;
	wire [4-1:0] node35065;
	wire [4-1:0] node35068;
	wire [4-1:0] node35071;
	wire [4-1:0] node35073;
	wire [4-1:0] node35076;
	wire [4-1:0] node35078;
	wire [4-1:0] node35081;
	wire [4-1:0] node35082;
	wire [4-1:0] node35083;
	wire [4-1:0] node35084;
	wire [4-1:0] node35085;
	wire [4-1:0] node35086;
	wire [4-1:0] node35087;
	wire [4-1:0] node35088;
	wire [4-1:0] node35089;
	wire [4-1:0] node35091;
	wire [4-1:0] node35092;
	wire [4-1:0] node35095;
	wire [4-1:0] node35098;
	wire [4-1:0] node35099;
	wire [4-1:0] node35100;
	wire [4-1:0] node35103;
	wire [4-1:0] node35106;
	wire [4-1:0] node35107;
	wire [4-1:0] node35110;
	wire [4-1:0] node35113;
	wire [4-1:0] node35114;
	wire [4-1:0] node35117;
	wire [4-1:0] node35120;
	wire [4-1:0] node35121;
	wire [4-1:0] node35122;
	wire [4-1:0] node35123;
	wire [4-1:0] node35127;
	wire [4-1:0] node35128;
	wire [4-1:0] node35132;
	wire [4-1:0] node35133;
	wire [4-1:0] node35134;
	wire [4-1:0] node35138;
	wire [4-1:0] node35139;
	wire [4-1:0] node35143;
	wire [4-1:0] node35144;
	wire [4-1:0] node35145;
	wire [4-1:0] node35146;
	wire [4-1:0] node35150;
	wire [4-1:0] node35151;
	wire [4-1:0] node35152;
	wire [4-1:0] node35156;
	wire [4-1:0] node35157;
	wire [4-1:0] node35161;
	wire [4-1:0] node35162;
	wire [4-1:0] node35163;
	wire [4-1:0] node35165;
	wire [4-1:0] node35168;
	wire [4-1:0] node35169;
	wire [4-1:0] node35170;
	wire [4-1:0] node35174;
	wire [4-1:0] node35175;
	wire [4-1:0] node35179;
	wire [4-1:0] node35180;
	wire [4-1:0] node35181;
	wire [4-1:0] node35182;
	wire [4-1:0] node35185;
	wire [4-1:0] node35188;
	wire [4-1:0] node35190;
	wire [4-1:0] node35193;
	wire [4-1:0] node35194;
	wire [4-1:0] node35197;
	wire [4-1:0] node35200;
	wire [4-1:0] node35201;
	wire [4-1:0] node35202;
	wire [4-1:0] node35203;
	wire [4-1:0] node35204;
	wire [4-1:0] node35205;
	wire [4-1:0] node35206;
	wire [4-1:0] node35209;
	wire [4-1:0] node35212;
	wire [4-1:0] node35213;
	wire [4-1:0] node35217;
	wire [4-1:0] node35220;
	wire [4-1:0] node35221;
	wire [4-1:0] node35223;
	wire [4-1:0] node35226;
	wire [4-1:0] node35227;
	wire [4-1:0] node35228;
	wire [4-1:0] node35232;
	wire [4-1:0] node35233;
	wire [4-1:0] node35237;
	wire [4-1:0] node35238;
	wire [4-1:0] node35239;
	wire [4-1:0] node35240;
	wire [4-1:0] node35241;
	wire [4-1:0] node35244;
	wire [4-1:0] node35247;
	wire [4-1:0] node35249;
	wire [4-1:0] node35252;
	wire [4-1:0] node35253;
	wire [4-1:0] node35256;
	wire [4-1:0] node35259;
	wire [4-1:0] node35260;
	wire [4-1:0] node35261;
	wire [4-1:0] node35262;
	wire [4-1:0] node35266;
	wire [4-1:0] node35267;
	wire [4-1:0] node35271;
	wire [4-1:0] node35272;
	wire [4-1:0] node35273;
	wire [4-1:0] node35277;
	wire [4-1:0] node35279;
	wire [4-1:0] node35282;
	wire [4-1:0] node35283;
	wire [4-1:0] node35284;
	wire [4-1:0] node35285;
	wire [4-1:0] node35287;
	wire [4-1:0] node35290;
	wire [4-1:0] node35291;
	wire [4-1:0] node35292;
	wire [4-1:0] node35296;
	wire [4-1:0] node35299;
	wire [4-1:0] node35300;
	wire [4-1:0] node35302;
	wire [4-1:0] node35303;
	wire [4-1:0] node35307;
	wire [4-1:0] node35308;
	wire [4-1:0] node35309;
	wire [4-1:0] node35312;
	wire [4-1:0] node35315;
	wire [4-1:0] node35316;
	wire [4-1:0] node35320;
	wire [4-1:0] node35321;
	wire [4-1:0] node35322;
	wire [4-1:0] node35323;
	wire [4-1:0] node35324;
	wire [4-1:0] node35327;
	wire [4-1:0] node35331;
	wire [4-1:0] node35332;
	wire [4-1:0] node35335;
	wire [4-1:0] node35338;
	wire [4-1:0] node35339;
	wire [4-1:0] node35341;
	wire [4-1:0] node35344;
	wire [4-1:0] node35346;
	wire [4-1:0] node35349;
	wire [4-1:0] node35350;
	wire [4-1:0] node35351;
	wire [4-1:0] node35352;
	wire [4-1:0] node35353;
	wire [4-1:0] node35354;
	wire [4-1:0] node35355;
	wire [4-1:0] node35358;
	wire [4-1:0] node35359;
	wire [4-1:0] node35363;
	wire [4-1:0] node35364;
	wire [4-1:0] node35365;
	wire [4-1:0] node35368;
	wire [4-1:0] node35371;
	wire [4-1:0] node35372;
	wire [4-1:0] node35375;
	wire [4-1:0] node35378;
	wire [4-1:0] node35379;
	wire [4-1:0] node35380;
	wire [4-1:0] node35381;
	wire [4-1:0] node35386;
	wire [4-1:0] node35387;
	wire [4-1:0] node35390;
	wire [4-1:0] node35393;
	wire [4-1:0] node35394;
	wire [4-1:0] node35395;
	wire [4-1:0] node35396;
	wire [4-1:0] node35399;
	wire [4-1:0] node35400;
	wire [4-1:0] node35404;
	wire [4-1:0] node35405;
	wire [4-1:0] node35406;
	wire [4-1:0] node35409;
	wire [4-1:0] node35413;
	wire [4-1:0] node35414;
	wire [4-1:0] node35415;
	wire [4-1:0] node35417;
	wire [4-1:0] node35420;
	wire [4-1:0] node35423;
	wire [4-1:0] node35424;
	wire [4-1:0] node35425;
	wire [4-1:0] node35429;
	wire [4-1:0] node35430;
	wire [4-1:0] node35433;
	wire [4-1:0] node35436;
	wire [4-1:0] node35437;
	wire [4-1:0] node35438;
	wire [4-1:0] node35439;
	wire [4-1:0] node35441;
	wire [4-1:0] node35442;
	wire [4-1:0] node35445;
	wire [4-1:0] node35448;
	wire [4-1:0] node35449;
	wire [4-1:0] node35452;
	wire [4-1:0] node35455;
	wire [4-1:0] node35456;
	wire [4-1:0] node35457;
	wire [4-1:0] node35458;
	wire [4-1:0] node35462;
	wire [4-1:0] node35463;
	wire [4-1:0] node35466;
	wire [4-1:0] node35469;
	wire [4-1:0] node35471;
	wire [4-1:0] node35474;
	wire [4-1:0] node35475;
	wire [4-1:0] node35476;
	wire [4-1:0] node35478;
	wire [4-1:0] node35479;
	wire [4-1:0] node35482;
	wire [4-1:0] node35485;
	wire [4-1:0] node35487;
	wire [4-1:0] node35490;
	wire [4-1:0] node35491;
	wire [4-1:0] node35492;
	wire [4-1:0] node35493;
	wire [4-1:0] node35496;
	wire [4-1:0] node35500;
	wire [4-1:0] node35502;
	wire [4-1:0] node35505;
	wire [4-1:0] node35506;
	wire [4-1:0] node35507;
	wire [4-1:0] node35508;
	wire [4-1:0] node35510;
	wire [4-1:0] node35512;
	wire [4-1:0] node35513;
	wire [4-1:0] node35517;
	wire [4-1:0] node35518;
	wire [4-1:0] node35520;
	wire [4-1:0] node35523;
	wire [4-1:0] node35524;
	wire [4-1:0] node35527;
	wire [4-1:0] node35530;
	wire [4-1:0] node35531;
	wire [4-1:0] node35532;
	wire [4-1:0] node35533;
	wire [4-1:0] node35537;
	wire [4-1:0] node35538;
	wire [4-1:0] node35540;
	wire [4-1:0] node35543;
	wire [4-1:0] node35545;
	wire [4-1:0] node35548;
	wire [4-1:0] node35549;
	wire [4-1:0] node35550;
	wire [4-1:0] node35551;
	wire [4-1:0] node35555;
	wire [4-1:0] node35556;
	wire [4-1:0] node35560;
	wire [4-1:0] node35562;
	wire [4-1:0] node35563;
	wire [4-1:0] node35567;
	wire [4-1:0] node35568;
	wire [4-1:0] node35569;
	wire [4-1:0] node35570;
	wire [4-1:0] node35571;
	wire [4-1:0] node35575;
	wire [4-1:0] node35577;
	wire [4-1:0] node35578;
	wire [4-1:0] node35582;
	wire [4-1:0] node35583;
	wire [4-1:0] node35584;
	wire [4-1:0] node35585;
	wire [4-1:0] node35588;
	wire [4-1:0] node35592;
	wire [4-1:0] node35593;
	wire [4-1:0] node35596;
	wire [4-1:0] node35599;
	wire [4-1:0] node35600;
	wire [4-1:0] node35601;
	wire [4-1:0] node35603;
	wire [4-1:0] node35606;
	wire [4-1:0] node35607;
	wire [4-1:0] node35610;
	wire [4-1:0] node35613;
	wire [4-1:0] node35614;
	wire [4-1:0] node35615;
	wire [4-1:0] node35616;
	wire [4-1:0] node35619;
	wire [4-1:0] node35622;
	wire [4-1:0] node35623;
	wire [4-1:0] node35627;
	wire [4-1:0] node35628;
	wire [4-1:0] node35632;
	wire [4-1:0] node35633;
	wire [4-1:0] node35634;
	wire [4-1:0] node35635;
	wire [4-1:0] node35636;
	wire [4-1:0] node35637;
	wire [4-1:0] node35638;
	wire [4-1:0] node35639;
	wire [4-1:0] node35643;
	wire [4-1:0] node35644;
	wire [4-1:0] node35648;
	wire [4-1:0] node35649;
	wire [4-1:0] node35650;
	wire [4-1:0] node35654;
	wire [4-1:0] node35655;
	wire [4-1:0] node35659;
	wire [4-1:0] node35660;
	wire [4-1:0] node35661;
	wire [4-1:0] node35662;
	wire [4-1:0] node35666;
	wire [4-1:0] node35669;
	wire [4-1:0] node35670;
	wire [4-1:0] node35671;
	wire [4-1:0] node35675;
	wire [4-1:0] node35676;
	wire [4-1:0] node35680;
	wire [4-1:0] node35681;
	wire [4-1:0] node35682;
	wire [4-1:0] node35683;
	wire [4-1:0] node35684;
	wire [4-1:0] node35687;
	wire [4-1:0] node35690;
	wire [4-1:0] node35691;
	wire [4-1:0] node35692;
	wire [4-1:0] node35695;
	wire [4-1:0] node35698;
	wire [4-1:0] node35699;
	wire [4-1:0] node35702;
	wire [4-1:0] node35705;
	wire [4-1:0] node35706;
	wire [4-1:0] node35708;
	wire [4-1:0] node35711;
	wire [4-1:0] node35712;
	wire [4-1:0] node35715;
	wire [4-1:0] node35718;
	wire [4-1:0] node35719;
	wire [4-1:0] node35720;
	wire [4-1:0] node35721;
	wire [4-1:0] node35723;
	wire [4-1:0] node35727;
	wire [4-1:0] node35728;
	wire [4-1:0] node35729;
	wire [4-1:0] node35733;
	wire [4-1:0] node35735;
	wire [4-1:0] node35738;
	wire [4-1:0] node35739;
	wire [4-1:0] node35740;
	wire [4-1:0] node35741;
	wire [4-1:0] node35744;
	wire [4-1:0] node35747;
	wire [4-1:0] node35748;
	wire [4-1:0] node35751;
	wire [4-1:0] node35754;
	wire [4-1:0] node35755;
	wire [4-1:0] node35756;
	wire [4-1:0] node35760;
	wire [4-1:0] node35763;
	wire [4-1:0] node35764;
	wire [4-1:0] node35765;
	wire [4-1:0] node35766;
	wire [4-1:0] node35767;
	wire [4-1:0] node35768;
	wire [4-1:0] node35769;
	wire [4-1:0] node35774;
	wire [4-1:0] node35775;
	wire [4-1:0] node35776;
	wire [4-1:0] node35779;
	wire [4-1:0] node35782;
	wire [4-1:0] node35784;
	wire [4-1:0] node35787;
	wire [4-1:0] node35788;
	wire [4-1:0] node35789;
	wire [4-1:0] node35790;
	wire [4-1:0] node35794;
	wire [4-1:0] node35795;
	wire [4-1:0] node35799;
	wire [4-1:0] node35800;
	wire [4-1:0] node35801;
	wire [4-1:0] node35805;
	wire [4-1:0] node35806;
	wire [4-1:0] node35810;
	wire [4-1:0] node35811;
	wire [4-1:0] node35812;
	wire [4-1:0] node35814;
	wire [4-1:0] node35815;
	wire [4-1:0] node35818;
	wire [4-1:0] node35821;
	wire [4-1:0] node35822;
	wire [4-1:0] node35825;
	wire [4-1:0] node35828;
	wire [4-1:0] node35829;
	wire [4-1:0] node35830;
	wire [4-1:0] node35831;
	wire [4-1:0] node35836;
	wire [4-1:0] node35837;
	wire [4-1:0] node35838;
	wire [4-1:0] node35843;
	wire [4-1:0] node35844;
	wire [4-1:0] node35845;
	wire [4-1:0] node35846;
	wire [4-1:0] node35847;
	wire [4-1:0] node35848;
	wire [4-1:0] node35851;
	wire [4-1:0] node35855;
	wire [4-1:0] node35856;
	wire [4-1:0] node35859;
	wire [4-1:0] node35862;
	wire [4-1:0] node35863;
	wire [4-1:0] node35864;
	wire [4-1:0] node35865;
	wire [4-1:0] node35869;
	wire [4-1:0] node35870;
	wire [4-1:0] node35874;
	wire [4-1:0] node35876;
	wire [4-1:0] node35879;
	wire [4-1:0] node35880;
	wire [4-1:0] node35881;
	wire [4-1:0] node35882;
	wire [4-1:0] node35883;
	wire [4-1:0] node35886;
	wire [4-1:0] node35889;
	wire [4-1:0] node35890;
	wire [4-1:0] node35893;
	wire [4-1:0] node35896;
	wire [4-1:0] node35897;
	wire [4-1:0] node35898;
	wire [4-1:0] node35901;
	wire [4-1:0] node35905;
	wire [4-1:0] node35906;
	wire [4-1:0] node35908;
	wire [4-1:0] node35911;
	wire [4-1:0] node35912;
	wire [4-1:0] node35915;
	wire [4-1:0] node35918;
	wire [4-1:0] node35919;
	wire [4-1:0] node35920;
	wire [4-1:0] node35921;
	wire [4-1:0] node35922;
	wire [4-1:0] node35923;
	wire [4-1:0] node35924;
	wire [4-1:0] node35928;
	wire [4-1:0] node35929;
	wire [4-1:0] node35933;
	wire [4-1:0] node35934;
	wire [4-1:0] node35935;
	wire [4-1:0] node35939;
	wire [4-1:0] node35940;
	wire [4-1:0] node35944;
	wire [4-1:0] node35945;
	wire [4-1:0] node35946;
	wire [4-1:0] node35947;
	wire [4-1:0] node35951;
	wire [4-1:0] node35954;
	wire [4-1:0] node35956;
	wire [4-1:0] node35959;
	wire [4-1:0] node35960;
	wire [4-1:0] node35961;
	wire [4-1:0] node35962;
	wire [4-1:0] node35963;
	wire [4-1:0] node35966;
	wire [4-1:0] node35969;
	wire [4-1:0] node35970;
	wire [4-1:0] node35973;
	wire [4-1:0] node35976;
	wire [4-1:0] node35977;
	wire [4-1:0] node35980;
	wire [4-1:0] node35983;
	wire [4-1:0] node35984;
	wire [4-1:0] node35985;
	wire [4-1:0] node35986;
	wire [4-1:0] node35990;
	wire [4-1:0] node35991;
	wire [4-1:0] node35992;
	wire [4-1:0] node35997;
	wire [4-1:0] node35998;
	wire [4-1:0] node35999;
	wire [4-1:0] node36000;
	wire [4-1:0] node36003;
	wire [4-1:0] node36006;
	wire [4-1:0] node36007;
	wire [4-1:0] node36010;
	wire [4-1:0] node36013;
	wire [4-1:0] node36014;
	wire [4-1:0] node36017;
	wire [4-1:0] node36020;
	wire [4-1:0] node36021;
	wire [4-1:0] node36022;
	wire [4-1:0] node36023;
	wire [4-1:0] node36024;
	wire [4-1:0] node36027;
	wire [4-1:0] node36028;
	wire [4-1:0] node36029;
	wire [4-1:0] node36033;
	wire [4-1:0] node36034;
	wire [4-1:0] node36038;
	wire [4-1:0] node36039;
	wire [4-1:0] node36040;
	wire [4-1:0] node36041;
	wire [4-1:0] node36046;
	wire [4-1:0] node36047;
	wire [4-1:0] node36048;
	wire [4-1:0] node36051;
	wire [4-1:0] node36055;
	wire [4-1:0] node36056;
	wire [4-1:0] node36057;
	wire [4-1:0] node36058;
	wire [4-1:0] node36059;
	wire [4-1:0] node36062;
	wire [4-1:0] node36066;
	wire [4-1:0] node36068;
	wire [4-1:0] node36069;
	wire [4-1:0] node36072;
	wire [4-1:0] node36075;
	wire [4-1:0] node36076;
	wire [4-1:0] node36077;
	wire [4-1:0] node36078;
	wire [4-1:0] node36082;
	wire [4-1:0] node36083;
	wire [4-1:0] node36086;
	wire [4-1:0] node36089;
	wire [4-1:0] node36090;
	wire [4-1:0] node36091;
	wire [4-1:0] node36095;
	wire [4-1:0] node36096;
	wire [4-1:0] node36099;
	wire [4-1:0] node36102;
	wire [4-1:0] node36103;
	wire [4-1:0] node36104;
	wire [4-1:0] node36105;
	wire [4-1:0] node36106;
	wire [4-1:0] node36107;
	wire [4-1:0] node36110;
	wire [4-1:0] node36113;
	wire [4-1:0] node36115;
	wire [4-1:0] node36118;
	wire [4-1:0] node36119;
	wire [4-1:0] node36120;
	wire [4-1:0] node36123;
	wire [4-1:0] node36126;
	wire [4-1:0] node36127;
	wire [4-1:0] node36130;
	wire [4-1:0] node36133;
	wire [4-1:0] node36134;
	wire [4-1:0] node36135;
	wire [4-1:0] node36136;
	wire [4-1:0] node36139;
	wire [4-1:0] node36142;
	wire [4-1:0] node36143;
	wire [4-1:0] node36146;
	wire [4-1:0] node36149;
	wire [4-1:0] node36151;
	wire [4-1:0] node36152;
	wire [4-1:0] node36155;
	wire [4-1:0] node36158;
	wire [4-1:0] node36159;
	wire [4-1:0] node36160;
	wire [4-1:0] node36161;
	wire [4-1:0] node36164;
	wire [4-1:0] node36167;
	wire [4-1:0] node36168;
	wire [4-1:0] node36171;
	wire [4-1:0] node36174;
	wire [4-1:0] node36175;
	wire [4-1:0] node36176;
	wire [4-1:0] node36177;
	wire [4-1:0] node36180;
	wire [4-1:0] node36183;
	wire [4-1:0] node36184;
	wire [4-1:0] node36187;
	wire [4-1:0] node36190;
	wire [4-1:0] node36191;
	wire [4-1:0] node36192;
	wire [4-1:0] node36197;
	wire [4-1:0] node36198;
	wire [4-1:0] node36199;
	wire [4-1:0] node36200;
	wire [4-1:0] node36201;
	wire [4-1:0] node36202;
	wire [4-1:0] node36203;
	wire [4-1:0] node36204;
	wire [4-1:0] node36206;
	wire [4-1:0] node36207;
	wire [4-1:0] node36210;
	wire [4-1:0] node36213;
	wire [4-1:0] node36214;
	wire [4-1:0] node36216;
	wire [4-1:0] node36219;
	wire [4-1:0] node36220;
	wire [4-1:0] node36223;
	wire [4-1:0] node36226;
	wire [4-1:0] node36227;
	wire [4-1:0] node36228;
	wire [4-1:0] node36231;
	wire [4-1:0] node36232;
	wire [4-1:0] node36236;
	wire [4-1:0] node36237;
	wire [4-1:0] node36239;
	wire [4-1:0] node36242;
	wire [4-1:0] node36244;
	wire [4-1:0] node36247;
	wire [4-1:0] node36248;
	wire [4-1:0] node36249;
	wire [4-1:0] node36250;
	wire [4-1:0] node36252;
	wire [4-1:0] node36255;
	wire [4-1:0] node36256;
	wire [4-1:0] node36260;
	wire [4-1:0] node36261;
	wire [4-1:0] node36264;
	wire [4-1:0] node36267;
	wire [4-1:0] node36268;
	wire [4-1:0] node36269;
	wire [4-1:0] node36272;
	wire [4-1:0] node36275;
	wire [4-1:0] node36276;
	wire [4-1:0] node36280;
	wire [4-1:0] node36281;
	wire [4-1:0] node36282;
	wire [4-1:0] node36283;
	wire [4-1:0] node36285;
	wire [4-1:0] node36286;
	wire [4-1:0] node36290;
	wire [4-1:0] node36291;
	wire [4-1:0] node36292;
	wire [4-1:0] node36296;
	wire [4-1:0] node36299;
	wire [4-1:0] node36300;
	wire [4-1:0] node36301;
	wire [4-1:0] node36303;
	wire [4-1:0] node36306;
	wire [4-1:0] node36307;
	wire [4-1:0] node36311;
	wire [4-1:0] node36312;
	wire [4-1:0] node36315;
	wire [4-1:0] node36318;
	wire [4-1:0] node36319;
	wire [4-1:0] node36320;
	wire [4-1:0] node36323;
	wire [4-1:0] node36324;
	wire [4-1:0] node36325;
	wire [4-1:0] node36329;
	wire [4-1:0] node36330;
	wire [4-1:0] node36334;
	wire [4-1:0] node36335;
	wire [4-1:0] node36337;
	wire [4-1:0] node36340;
	wire [4-1:0] node36342;
	wire [4-1:0] node36345;
	wire [4-1:0] node36346;
	wire [4-1:0] node36347;
	wire [4-1:0] node36348;
	wire [4-1:0] node36349;
	wire [4-1:0] node36351;
	wire [4-1:0] node36354;
	wire [4-1:0] node36355;
	wire [4-1:0] node36358;
	wire [4-1:0] node36361;
	wire [4-1:0] node36362;
	wire [4-1:0] node36363;
	wire [4-1:0] node36368;
	wire [4-1:0] node36369;
	wire [4-1:0] node36370;
	wire [4-1:0] node36371;
	wire [4-1:0] node36372;
	wire [4-1:0] node36375;
	wire [4-1:0] node36378;
	wire [4-1:0] node36379;
	wire [4-1:0] node36382;
	wire [4-1:0] node36385;
	wire [4-1:0] node36386;
	wire [4-1:0] node36388;
	wire [4-1:0] node36391;
	wire [4-1:0] node36392;
	wire [4-1:0] node36395;
	wire [4-1:0] node36398;
	wire [4-1:0] node36399;
	wire [4-1:0] node36400;
	wire [4-1:0] node36403;
	wire [4-1:0] node36406;
	wire [4-1:0] node36407;
	wire [4-1:0] node36409;
	wire [4-1:0] node36413;
	wire [4-1:0] node36414;
	wire [4-1:0] node36415;
	wire [4-1:0] node36416;
	wire [4-1:0] node36417;
	wire [4-1:0] node36421;
	wire [4-1:0] node36422;
	wire [4-1:0] node36426;
	wire [4-1:0] node36427;
	wire [4-1:0] node36428;
	wire [4-1:0] node36432;
	wire [4-1:0] node36433;
	wire [4-1:0] node36437;
	wire [4-1:0] node36438;
	wire [4-1:0] node36439;
	wire [4-1:0] node36440;
	wire [4-1:0] node36444;
	wire [4-1:0] node36445;
	wire [4-1:0] node36448;
	wire [4-1:0] node36451;
	wire [4-1:0] node36452;
	wire [4-1:0] node36455;
	wire [4-1:0] node36458;
	wire [4-1:0] node36459;
	wire [4-1:0] node36460;
	wire [4-1:0] node36461;
	wire [4-1:0] node36462;
	wire [4-1:0] node36463;
	wire [4-1:0] node36465;
	wire [4-1:0] node36468;
	wire [4-1:0] node36469;
	wire [4-1:0] node36470;
	wire [4-1:0] node36473;
	wire [4-1:0] node36477;
	wire [4-1:0] node36478;
	wire [4-1:0] node36479;
	wire [4-1:0] node36480;
	wire [4-1:0] node36483;
	wire [4-1:0] node36486;
	wire [4-1:0] node36487;
	wire [4-1:0] node36490;
	wire [4-1:0] node36493;
	wire [4-1:0] node36494;
	wire [4-1:0] node36497;
	wire [4-1:0] node36500;
	wire [4-1:0] node36501;
	wire [4-1:0] node36502;
	wire [4-1:0] node36503;
	wire [4-1:0] node36505;
	wire [4-1:0] node36508;
	wire [4-1:0] node36509;
	wire [4-1:0] node36513;
	wire [4-1:0] node36514;
	wire [4-1:0] node36518;
	wire [4-1:0] node36519;
	wire [4-1:0] node36520;
	wire [4-1:0] node36521;
	wire [4-1:0] node36525;
	wire [4-1:0] node36526;
	wire [4-1:0] node36529;
	wire [4-1:0] node36532;
	wire [4-1:0] node36533;
	wire [4-1:0] node36537;
	wire [4-1:0] node36538;
	wire [4-1:0] node36539;
	wire [4-1:0] node36540;
	wire [4-1:0] node36541;
	wire [4-1:0] node36544;
	wire [4-1:0] node36547;
	wire [4-1:0] node36549;
	wire [4-1:0] node36550;
	wire [4-1:0] node36554;
	wire [4-1:0] node36555;
	wire [4-1:0] node36556;
	wire [4-1:0] node36557;
	wire [4-1:0] node36561;
	wire [4-1:0] node36564;
	wire [4-1:0] node36565;
	wire [4-1:0] node36566;
	wire [4-1:0] node36571;
	wire [4-1:0] node36572;
	wire [4-1:0] node36573;
	wire [4-1:0] node36575;
	wire [4-1:0] node36578;
	wire [4-1:0] node36579;
	wire [4-1:0] node36580;
	wire [4-1:0] node36584;
	wire [4-1:0] node36585;
	wire [4-1:0] node36589;
	wire [4-1:0] node36590;
	wire [4-1:0] node36591;
	wire [4-1:0] node36595;
	wire [4-1:0] node36596;
	wire [4-1:0] node36599;
	wire [4-1:0] node36602;
	wire [4-1:0] node36603;
	wire [4-1:0] node36604;
	wire [4-1:0] node36605;
	wire [4-1:0] node36606;
	wire [4-1:0] node36608;
	wire [4-1:0] node36609;
	wire [4-1:0] node36612;
	wire [4-1:0] node36615;
	wire [4-1:0] node36616;
	wire [4-1:0] node36620;
	wire [4-1:0] node36621;
	wire [4-1:0] node36622;
	wire [4-1:0] node36623;
	wire [4-1:0] node36626;
	wire [4-1:0] node36629;
	wire [4-1:0] node36630;
	wire [4-1:0] node36633;
	wire [4-1:0] node36636;
	wire [4-1:0] node36637;
	wire [4-1:0] node36638;
	wire [4-1:0] node36641;
	wire [4-1:0] node36645;
	wire [4-1:0] node36646;
	wire [4-1:0] node36648;
	wire [4-1:0] node36649;
	wire [4-1:0] node36650;
	wire [4-1:0] node36654;
	wire [4-1:0] node36655;
	wire [4-1:0] node36659;
	wire [4-1:0] node36660;
	wire [4-1:0] node36661;
	wire [4-1:0] node36665;
	wire [4-1:0] node36667;
	wire [4-1:0] node36670;
	wire [4-1:0] node36671;
	wire [4-1:0] node36672;
	wire [4-1:0] node36673;
	wire [4-1:0] node36676;
	wire [4-1:0] node36677;
	wire [4-1:0] node36678;
	wire [4-1:0] node36682;
	wire [4-1:0] node36683;
	wire [4-1:0] node36687;
	wire [4-1:0] node36688;
	wire [4-1:0] node36689;
	wire [4-1:0] node36691;
	wire [4-1:0] node36695;
	wire [4-1:0] node36696;
	wire [4-1:0] node36697;
	wire [4-1:0] node36701;
	wire [4-1:0] node36702;
	wire [4-1:0] node36706;
	wire [4-1:0] node36707;
	wire [4-1:0] node36708;
	wire [4-1:0] node36709;
	wire [4-1:0] node36713;
	wire [4-1:0] node36714;
	wire [4-1:0] node36718;
	wire [4-1:0] node36719;
	wire [4-1:0] node36720;
	wire [4-1:0] node36724;
	wire [4-1:0] node36725;
	wire [4-1:0] node36729;
	wire [4-1:0] node36730;
	wire [4-1:0] node36731;
	wire [4-1:0] node36732;
	wire [4-1:0] node36733;
	wire [4-1:0] node36734;
	wire [4-1:0] node36735;
	wire [4-1:0] node36736;
	wire [4-1:0] node36737;
	wire [4-1:0] node36742;
	wire [4-1:0] node36743;
	wire [4-1:0] node36746;
	wire [4-1:0] node36749;
	wire [4-1:0] node36750;
	wire [4-1:0] node36751;
	wire [4-1:0] node36752;
	wire [4-1:0] node36756;
	wire [4-1:0] node36757;
	wire [4-1:0] node36762;
	wire [4-1:0] node36763;
	wire [4-1:0] node36764;
	wire [4-1:0] node36765;
	wire [4-1:0] node36766;
	wire [4-1:0] node36769;
	wire [4-1:0] node36773;
	wire [4-1:0] node36774;
	wire [4-1:0] node36776;
	wire [4-1:0] node36780;
	wire [4-1:0] node36781;
	wire [4-1:0] node36782;
	wire [4-1:0] node36784;
	wire [4-1:0] node36787;
	wire [4-1:0] node36789;
	wire [4-1:0] node36792;
	wire [4-1:0] node36793;
	wire [4-1:0] node36794;
	wire [4-1:0] node36798;
	wire [4-1:0] node36801;
	wire [4-1:0] node36802;
	wire [4-1:0] node36803;
	wire [4-1:0] node36804;
	wire [4-1:0] node36805;
	wire [4-1:0] node36808;
	wire [4-1:0] node36809;
	wire [4-1:0] node36813;
	wire [4-1:0] node36814;
	wire [4-1:0] node36817;
	wire [4-1:0] node36818;
	wire [4-1:0] node36822;
	wire [4-1:0] node36823;
	wire [4-1:0] node36825;
	wire [4-1:0] node36826;
	wire [4-1:0] node36830;
	wire [4-1:0] node36831;
	wire [4-1:0] node36832;
	wire [4-1:0] node36836;
	wire [4-1:0] node36839;
	wire [4-1:0] node36840;
	wire [4-1:0] node36841;
	wire [4-1:0] node36842;
	wire [4-1:0] node36843;
	wire [4-1:0] node36846;
	wire [4-1:0] node36849;
	wire [4-1:0] node36850;
	wire [4-1:0] node36854;
	wire [4-1:0] node36855;
	wire [4-1:0] node36856;
	wire [4-1:0] node36859;
	wire [4-1:0] node36862;
	wire [4-1:0] node36863;
	wire [4-1:0] node36866;
	wire [4-1:0] node36869;
	wire [4-1:0] node36870;
	wire [4-1:0] node36871;
	wire [4-1:0] node36872;
	wire [4-1:0] node36875;
	wire [4-1:0] node36878;
	wire [4-1:0] node36880;
	wire [4-1:0] node36883;
	wire [4-1:0] node36884;
	wire [4-1:0] node36887;
	wire [4-1:0] node36890;
	wire [4-1:0] node36891;
	wire [4-1:0] node36892;
	wire [4-1:0] node36893;
	wire [4-1:0] node36894;
	wire [4-1:0] node36895;
	wire [4-1:0] node36896;
	wire [4-1:0] node36900;
	wire [4-1:0] node36901;
	wire [4-1:0] node36904;
	wire [4-1:0] node36907;
	wire [4-1:0] node36908;
	wire [4-1:0] node36911;
	wire [4-1:0] node36914;
	wire [4-1:0] node36915;
	wire [4-1:0] node36916;
	wire [4-1:0] node36917;
	wire [4-1:0] node36920;
	wire [4-1:0] node36923;
	wire [4-1:0] node36924;
	wire [4-1:0] node36928;
	wire [4-1:0] node36929;
	wire [4-1:0] node36930;
	wire [4-1:0] node36934;
	wire [4-1:0] node36935;
	wire [4-1:0] node36938;
	wire [4-1:0] node36941;
	wire [4-1:0] node36942;
	wire [4-1:0] node36943;
	wire [4-1:0] node36944;
	wire [4-1:0] node36945;
	wire [4-1:0] node36948;
	wire [4-1:0] node36952;
	wire [4-1:0] node36953;
	wire [4-1:0] node36954;
	wire [4-1:0] node36958;
	wire [4-1:0] node36959;
	wire [4-1:0] node36963;
	wire [4-1:0] node36964;
	wire [4-1:0] node36965;
	wire [4-1:0] node36966;
	wire [4-1:0] node36969;
	wire [4-1:0] node36972;
	wire [4-1:0] node36974;
	wire [4-1:0] node36977;
	wire [4-1:0] node36978;
	wire [4-1:0] node36980;
	wire [4-1:0] node36983;
	wire [4-1:0] node36984;
	wire [4-1:0] node36988;
	wire [4-1:0] node36989;
	wire [4-1:0] node36990;
	wire [4-1:0] node36991;
	wire [4-1:0] node36992;
	wire [4-1:0] node36993;
	wire [4-1:0] node36996;
	wire [4-1:0] node36999;
	wire [4-1:0] node37001;
	wire [4-1:0] node37004;
	wire [4-1:0] node37005;
	wire [4-1:0] node37007;
	wire [4-1:0] node37010;
	wire [4-1:0] node37012;
	wire [4-1:0] node37015;
	wire [4-1:0] node37016;
	wire [4-1:0] node37017;
	wire [4-1:0] node37018;
	wire [4-1:0] node37021;
	wire [4-1:0] node37024;
	wire [4-1:0] node37027;
	wire [4-1:0] node37029;
	wire [4-1:0] node37031;
	wire [4-1:0] node37034;
	wire [4-1:0] node37035;
	wire [4-1:0] node37036;
	wire [4-1:0] node37037;
	wire [4-1:0] node37038;
	wire [4-1:0] node37041;
	wire [4-1:0] node37044;
	wire [4-1:0] node37045;
	wire [4-1:0] node37048;
	wire [4-1:0] node37051;
	wire [4-1:0] node37052;
	wire [4-1:0] node37053;
	wire [4-1:0] node37056;
	wire [4-1:0] node37059;
	wire [4-1:0] node37062;
	wire [4-1:0] node37063;
	wire [4-1:0] node37064;
	wire [4-1:0] node37065;
	wire [4-1:0] node37068;
	wire [4-1:0] node37071;
	wire [4-1:0] node37072;
	wire [4-1:0] node37075;
	wire [4-1:0] node37078;
	wire [4-1:0] node37079;
	wire [4-1:0] node37081;
	wire [4-1:0] node37084;
	wire [4-1:0] node37085;
	wire [4-1:0] node37089;
	wire [4-1:0] node37090;
	wire [4-1:0] node37091;
	wire [4-1:0] node37092;
	wire [4-1:0] node37093;
	wire [4-1:0] node37094;
	wire [4-1:0] node37095;
	wire [4-1:0] node37096;
	wire [4-1:0] node37099;
	wire [4-1:0] node37103;
	wire [4-1:0] node37104;
	wire [4-1:0] node37107;
	wire [4-1:0] node37110;
	wire [4-1:0] node37111;
	wire [4-1:0] node37112;
	wire [4-1:0] node37113;
	wire [4-1:0] node37116;
	wire [4-1:0] node37120;
	wire [4-1:0] node37121;
	wire [4-1:0] node37124;
	wire [4-1:0] node37127;
	wire [4-1:0] node37128;
	wire [4-1:0] node37129;
	wire [4-1:0] node37130;
	wire [4-1:0] node37132;
	wire [4-1:0] node37135;
	wire [4-1:0] node37137;
	wire [4-1:0] node37140;
	wire [4-1:0] node37141;
	wire [4-1:0] node37142;
	wire [4-1:0] node37145;
	wire [4-1:0] node37148;
	wire [4-1:0] node37149;
	wire [4-1:0] node37152;
	wire [4-1:0] node37155;
	wire [4-1:0] node37156;
	wire [4-1:0] node37157;
	wire [4-1:0] node37158;
	wire [4-1:0] node37161;
	wire [4-1:0] node37164;
	wire [4-1:0] node37166;
	wire [4-1:0] node37169;
	wire [4-1:0] node37170;
	wire [4-1:0] node37171;
	wire [4-1:0] node37176;
	wire [4-1:0] node37177;
	wire [4-1:0] node37178;
	wire [4-1:0] node37179;
	wire [4-1:0] node37182;
	wire [4-1:0] node37183;
	wire [4-1:0] node37184;
	wire [4-1:0] node37188;
	wire [4-1:0] node37189;
	wire [4-1:0] node37193;
	wire [4-1:0] node37195;
	wire [4-1:0] node37196;
	wire [4-1:0] node37198;
	wire [4-1:0] node37202;
	wire [4-1:0] node37203;
	wire [4-1:0] node37204;
	wire [4-1:0] node37205;
	wire [4-1:0] node37206;
	wire [4-1:0] node37211;
	wire [4-1:0] node37212;
	wire [4-1:0] node37215;
	wire [4-1:0] node37216;
	wire [4-1:0] node37220;
	wire [4-1:0] node37221;
	wire [4-1:0] node37222;
	wire [4-1:0] node37223;
	wire [4-1:0] node37228;
	wire [4-1:0] node37230;
	wire [4-1:0] node37233;
	wire [4-1:0] node37234;
	wire [4-1:0] node37235;
	wire [4-1:0] node37236;
	wire [4-1:0] node37237;
	wire [4-1:0] node37239;
	wire [4-1:0] node37240;
	wire [4-1:0] node37244;
	wire [4-1:0] node37246;
	wire [4-1:0] node37247;
	wire [4-1:0] node37251;
	wire [4-1:0] node37252;
	wire [4-1:0] node37254;
	wire [4-1:0] node37256;
	wire [4-1:0] node37259;
	wire [4-1:0] node37260;
	wire [4-1:0] node37263;
	wire [4-1:0] node37266;
	wire [4-1:0] node37267;
	wire [4-1:0] node37268;
	wire [4-1:0] node37269;
	wire [4-1:0] node37270;
	wire [4-1:0] node37274;
	wire [4-1:0] node37275;
	wire [4-1:0] node37279;
	wire [4-1:0] node37280;
	wire [4-1:0] node37281;
	wire [4-1:0] node37286;
	wire [4-1:0] node37287;
	wire [4-1:0] node37288;
	wire [4-1:0] node37292;
	wire [4-1:0] node37293;
	wire [4-1:0] node37294;
	wire [4-1:0] node37298;
	wire [4-1:0] node37301;
	wire [4-1:0] node37302;
	wire [4-1:0] node37303;
	wire [4-1:0] node37304;
	wire [4-1:0] node37305;
	wire [4-1:0] node37306;
	wire [4-1:0] node37309;
	wire [4-1:0] node37313;
	wire [4-1:0] node37314;
	wire [4-1:0] node37316;
	wire [4-1:0] node37319;
	wire [4-1:0] node37320;
	wire [4-1:0] node37323;
	wire [4-1:0] node37326;
	wire [4-1:0] node37327;
	wire [4-1:0] node37330;
	wire [4-1:0] node37333;
	wire [4-1:0] node37334;
	wire [4-1:0] node37335;
	wire [4-1:0] node37336;
	wire [4-1:0] node37337;
	wire [4-1:0] node37340;
	wire [4-1:0] node37343;
	wire [4-1:0] node37344;
	wire [4-1:0] node37347;
	wire [4-1:0] node37350;
	wire [4-1:0] node37351;
	wire [4-1:0] node37353;
	wire [4-1:0] node37356;
	wire [4-1:0] node37358;
	wire [4-1:0] node37361;
	wire [4-1:0] node37362;
	wire [4-1:0] node37363;
	wire [4-1:0] node37364;
	wire [4-1:0] node37367;
	wire [4-1:0] node37371;
	wire [4-1:0] node37372;
	wire [4-1:0] node37374;
	wire [4-1:0] node37377;
	wire [4-1:0] node37379;
	wire [4-1:0] node37382;
	wire [4-1:0] node37383;
	wire [4-1:0] node37384;
	wire [4-1:0] node37385;
	wire [4-1:0] node37386;
	wire [4-1:0] node37387;
	wire [4-1:0] node37388;
	wire [4-1:0] node37389;
	wire [4-1:0] node37390;
	wire [4-1:0] node37391;
	wire [4-1:0] node37394;
	wire [4-1:0] node37397;
	wire [4-1:0] node37398;
	wire [4-1:0] node37401;
	wire [4-1:0] node37404;
	wire [4-1:0] node37405;
	wire [4-1:0] node37406;
	wire [4-1:0] node37409;
	wire [4-1:0] node37412;
	wire [4-1:0] node37413;
	wire [4-1:0] node37414;
	wire [4-1:0] node37418;
	wire [4-1:0] node37419;
	wire [4-1:0] node37422;
	wire [4-1:0] node37425;
	wire [4-1:0] node37426;
	wire [4-1:0] node37427;
	wire [4-1:0] node37428;
	wire [4-1:0] node37429;
	wire [4-1:0] node37430;
	wire [4-1:0] node37434;
	wire [4-1:0] node37435;
	wire [4-1:0] node37438;
	wire [4-1:0] node37441;
	wire [4-1:0] node37442;
	wire [4-1:0] node37443;
	wire [4-1:0] node37446;
	wire [4-1:0] node37450;
	wire [4-1:0] node37451;
	wire [4-1:0] node37452;
	wire [4-1:0] node37453;
	wire [4-1:0] node37457;
	wire [4-1:0] node37458;
	wire [4-1:0] node37462;
	wire [4-1:0] node37463;
	wire [4-1:0] node37464;
	wire [4-1:0] node37467;
	wire [4-1:0] node37470;
	wire [4-1:0] node37471;
	wire [4-1:0] node37474;
	wire [4-1:0] node37477;
	wire [4-1:0] node37478;
	wire [4-1:0] node37479;
	wire [4-1:0] node37480;
	wire [4-1:0] node37481;
	wire [4-1:0] node37484;
	wire [4-1:0] node37487;
	wire [4-1:0] node37488;
	wire [4-1:0] node37491;
	wire [4-1:0] node37494;
	wire [4-1:0] node37495;
	wire [4-1:0] node37496;
	wire [4-1:0] node37499;
	wire [4-1:0] node37502;
	wire [4-1:0] node37503;
	wire [4-1:0] node37506;
	wire [4-1:0] node37509;
	wire [4-1:0] node37510;
	wire [4-1:0] node37511;
	wire [4-1:0] node37512;
	wire [4-1:0] node37515;
	wire [4-1:0] node37519;
	wire [4-1:0] node37520;
	wire [4-1:0] node37522;
	wire [4-1:0] node37525;
	wire [4-1:0] node37526;
	wire [4-1:0] node37529;
	wire [4-1:0] node37532;
	wire [4-1:0] node37533;
	wire [4-1:0] node37534;
	wire [4-1:0] node37535;
	wire [4-1:0] node37536;
	wire [4-1:0] node37537;
	wire [4-1:0] node37539;
	wire [4-1:0] node37542;
	wire [4-1:0] node37544;
	wire [4-1:0] node37547;
	wire [4-1:0] node37548;
	wire [4-1:0] node37550;
	wire [4-1:0] node37554;
	wire [4-1:0] node37555;
	wire [4-1:0] node37556;
	wire [4-1:0] node37557;
	wire [4-1:0] node37560;
	wire [4-1:0] node37564;
	wire [4-1:0] node37565;
	wire [4-1:0] node37566;
	wire [4-1:0] node37571;
	wire [4-1:0] node37572;
	wire [4-1:0] node37573;
	wire [4-1:0] node37576;
	wire [4-1:0] node37577;
	wire [4-1:0] node37580;
	wire [4-1:0] node37582;
	wire [4-1:0] node37585;
	wire [4-1:0] node37586;
	wire [4-1:0] node37587;
	wire [4-1:0] node37590;
	wire [4-1:0] node37593;
	wire [4-1:0] node37594;
	wire [4-1:0] node37596;
	wire [4-1:0] node37599;
	wire [4-1:0] node37600;
	wire [4-1:0] node37603;
	wire [4-1:0] node37606;
	wire [4-1:0] node37607;
	wire [4-1:0] node37608;
	wire [4-1:0] node37609;
	wire [4-1:0] node37610;
	wire [4-1:0] node37612;
	wire [4-1:0] node37616;
	wire [4-1:0] node37617;
	wire [4-1:0] node37619;
	wire [4-1:0] node37622;
	wire [4-1:0] node37624;
	wire [4-1:0] node37627;
	wire [4-1:0] node37628;
	wire [4-1:0] node37630;
	wire [4-1:0] node37631;
	wire [4-1:0] node37634;
	wire [4-1:0] node37637;
	wire [4-1:0] node37638;
	wire [4-1:0] node37639;
	wire [4-1:0] node37642;
	wire [4-1:0] node37646;
	wire [4-1:0] node37647;
	wire [4-1:0] node37648;
	wire [4-1:0] node37649;
	wire [4-1:0] node37652;
	wire [4-1:0] node37654;
	wire [4-1:0] node37657;
	wire [4-1:0] node37658;
	wire [4-1:0] node37660;
	wire [4-1:0] node37663;
	wire [4-1:0] node37665;
	wire [4-1:0] node37668;
	wire [4-1:0] node37669;
	wire [4-1:0] node37670;
	wire [4-1:0] node37674;
	wire [4-1:0] node37675;
	wire [4-1:0] node37676;
	wire [4-1:0] node37679;
	wire [4-1:0] node37682;
	wire [4-1:0] node37683;
	wire [4-1:0] node37687;
	wire [4-1:0] node37688;
	wire [4-1:0] node37689;
	wire [4-1:0] node37690;
	wire [4-1:0] node37691;
	wire [4-1:0] node37692;
	wire [4-1:0] node37693;
	wire [4-1:0] node37697;
	wire [4-1:0] node37698;
	wire [4-1:0] node37699;
	wire [4-1:0] node37702;
	wire [4-1:0] node37705;
	wire [4-1:0] node37706;
	wire [4-1:0] node37709;
	wire [4-1:0] node37712;
	wire [4-1:0] node37713;
	wire [4-1:0] node37715;
	wire [4-1:0] node37716;
	wire [4-1:0] node37719;
	wire [4-1:0] node37722;
	wire [4-1:0] node37723;
	wire [4-1:0] node37725;
	wire [4-1:0] node37728;
	wire [4-1:0] node37730;
	wire [4-1:0] node37733;
	wire [4-1:0] node37734;
	wire [4-1:0] node37735;
	wire [4-1:0] node37737;
	wire [4-1:0] node37739;
	wire [4-1:0] node37742;
	wire [4-1:0] node37744;
	wire [4-1:0] node37747;
	wire [4-1:0] node37749;
	wire [4-1:0] node37752;
	wire [4-1:0] node37753;
	wire [4-1:0] node37754;
	wire [4-1:0] node37755;
	wire [4-1:0] node37756;
	wire [4-1:0] node37759;
	wire [4-1:0] node37762;
	wire [4-1:0] node37763;
	wire [4-1:0] node37766;
	wire [4-1:0] node37769;
	wire [4-1:0] node37770;
	wire [4-1:0] node37771;
	wire [4-1:0] node37775;
	wire [4-1:0] node37777;
	wire [4-1:0] node37780;
	wire [4-1:0] node37781;
	wire [4-1:0] node37782;
	wire [4-1:0] node37783;
	wire [4-1:0] node37786;
	wire [4-1:0] node37787;
	wire [4-1:0] node37792;
	wire [4-1:0] node37793;
	wire [4-1:0] node37794;
	wire [4-1:0] node37797;
	wire [4-1:0] node37800;
	wire [4-1:0] node37802;
	wire [4-1:0] node37804;
	wire [4-1:0] node37807;
	wire [4-1:0] node37808;
	wire [4-1:0] node37809;
	wire [4-1:0] node37810;
	wire [4-1:0] node37811;
	wire [4-1:0] node37812;
	wire [4-1:0] node37815;
	wire [4-1:0] node37818;
	wire [4-1:0] node37819;
	wire [4-1:0] node37822;
	wire [4-1:0] node37825;
	wire [4-1:0] node37826;
	wire [4-1:0] node37827;
	wire [4-1:0] node37828;
	wire [4-1:0] node37831;
	wire [4-1:0] node37835;
	wire [4-1:0] node37837;
	wire [4-1:0] node37838;
	wire [4-1:0] node37842;
	wire [4-1:0] node37843;
	wire [4-1:0] node37844;
	wire [4-1:0] node37846;
	wire [4-1:0] node37849;
	wire [4-1:0] node37850;
	wire [4-1:0] node37853;
	wire [4-1:0] node37856;
	wire [4-1:0] node37857;
	wire [4-1:0] node37858;
	wire [4-1:0] node37859;
	wire [4-1:0] node37864;
	wire [4-1:0] node37865;
	wire [4-1:0] node37868;
	wire [4-1:0] node37871;
	wire [4-1:0] node37872;
	wire [4-1:0] node37873;
	wire [4-1:0] node37874;
	wire [4-1:0] node37875;
	wire [4-1:0] node37876;
	wire [4-1:0] node37880;
	wire [4-1:0] node37881;
	wire [4-1:0] node37884;
	wire [4-1:0] node37887;
	wire [4-1:0] node37888;
	wire [4-1:0] node37889;
	wire [4-1:0] node37892;
	wire [4-1:0] node37895;
	wire [4-1:0] node37896;
	wire [4-1:0] node37900;
	wire [4-1:0] node37901;
	wire [4-1:0] node37903;
	wire [4-1:0] node37904;
	wire [4-1:0] node37907;
	wire [4-1:0] node37910;
	wire [4-1:0] node37911;
	wire [4-1:0] node37914;
	wire [4-1:0] node37917;
	wire [4-1:0] node37918;
	wire [4-1:0] node37919;
	wire [4-1:0] node37922;
	wire [4-1:0] node37925;
	wire [4-1:0] node37926;
	wire [4-1:0] node37928;
	wire [4-1:0] node37929;
	wire [4-1:0] node37932;
	wire [4-1:0] node37935;
	wire [4-1:0] node37936;
	wire [4-1:0] node37937;
	wire [4-1:0] node37940;
	wire [4-1:0] node37943;
	wire [4-1:0] node37944;
	wire [4-1:0] node37948;
	wire [4-1:0] node37949;
	wire [4-1:0] node37950;
	wire [4-1:0] node37951;
	wire [4-1:0] node37952;
	wire [4-1:0] node37953;
	wire [4-1:0] node37956;
	wire [4-1:0] node37959;
	wire [4-1:0] node37960;
	wire [4-1:0] node37961;
	wire [4-1:0] node37964;
	wire [4-1:0] node37967;
	wire [4-1:0] node37968;
	wire [4-1:0] node37969;
	wire [4-1:0] node37971;
	wire [4-1:0] node37975;
	wire [4-1:0] node37976;
	wire [4-1:0] node37979;
	wire [4-1:0] node37982;
	wire [4-1:0] node37983;
	wire [4-1:0] node37984;
	wire [4-1:0] node37985;
	wire [4-1:0] node37988;
	wire [4-1:0] node37991;
	wire [4-1:0] node37992;
	wire [4-1:0] node37993;
	wire [4-1:0] node37996;
	wire [4-1:0] node37999;
	wire [4-1:0] node38000;
	wire [4-1:0] node38003;
	wire [4-1:0] node38006;
	wire [4-1:0] node38007;
	wire [4-1:0] node38008;
	wire [4-1:0] node38010;
	wire [4-1:0] node38013;
	wire [4-1:0] node38014;
	wire [4-1:0] node38016;
	wire [4-1:0] node38019;
	wire [4-1:0] node38022;
	wire [4-1:0] node38023;
	wire [4-1:0] node38024;
	wire [4-1:0] node38027;
	wire [4-1:0] node38030;
	wire [4-1:0] node38031;
	wire [4-1:0] node38034;
	wire [4-1:0] node38037;
	wire [4-1:0] node38038;
	wire [4-1:0] node38039;
	wire [4-1:0] node38040;
	wire [4-1:0] node38041;
	wire [4-1:0] node38042;
	wire [4-1:0] node38046;
	wire [4-1:0] node38047;
	wire [4-1:0] node38050;
	wire [4-1:0] node38053;
	wire [4-1:0] node38054;
	wire [4-1:0] node38055;
	wire [4-1:0] node38058;
	wire [4-1:0] node38061;
	wire [4-1:0] node38062;
	wire [4-1:0] node38065;
	wire [4-1:0] node38068;
	wire [4-1:0] node38069;
	wire [4-1:0] node38070;
	wire [4-1:0] node38072;
	wire [4-1:0] node38075;
	wire [4-1:0] node38078;
	wire [4-1:0] node38079;
	wire [4-1:0] node38080;
	wire [4-1:0] node38083;
	wire [4-1:0] node38086;
	wire [4-1:0] node38087;
	wire [4-1:0] node38090;
	wire [4-1:0] node38093;
	wire [4-1:0] node38094;
	wire [4-1:0] node38095;
	wire [4-1:0] node38096;
	wire [4-1:0] node38097;
	wire [4-1:0] node38098;
	wire [4-1:0] node38102;
	wire [4-1:0] node38103;
	wire [4-1:0] node38107;
	wire [4-1:0] node38108;
	wire [4-1:0] node38111;
	wire [4-1:0] node38114;
	wire [4-1:0] node38115;
	wire [4-1:0] node38116;
	wire [4-1:0] node38117;
	wire [4-1:0] node38120;
	wire [4-1:0] node38123;
	wire [4-1:0] node38124;
	wire [4-1:0] node38127;
	wire [4-1:0] node38130;
	wire [4-1:0] node38131;
	wire [4-1:0] node38133;
	wire [4-1:0] node38136;
	wire [4-1:0] node38137;
	wire [4-1:0] node38140;
	wire [4-1:0] node38143;
	wire [4-1:0] node38144;
	wire [4-1:0] node38145;
	wire [4-1:0] node38146;
	wire [4-1:0] node38149;
	wire [4-1:0] node38152;
	wire [4-1:0] node38153;
	wire [4-1:0] node38156;
	wire [4-1:0] node38159;
	wire [4-1:0] node38160;
	wire [4-1:0] node38162;
	wire [4-1:0] node38163;
	wire [4-1:0] node38166;
	wire [4-1:0] node38169;
	wire [4-1:0] node38171;
	wire [4-1:0] node38173;
	wire [4-1:0] node38176;
	wire [4-1:0] node38177;
	wire [4-1:0] node38178;
	wire [4-1:0] node38179;
	wire [4-1:0] node38180;
	wire [4-1:0] node38181;
	wire [4-1:0] node38183;
	wire [4-1:0] node38186;
	wire [4-1:0] node38188;
	wire [4-1:0] node38191;
	wire [4-1:0] node38192;
	wire [4-1:0] node38194;
	wire [4-1:0] node38198;
	wire [4-1:0] node38199;
	wire [4-1:0] node38200;
	wire [4-1:0] node38202;
	wire [4-1:0] node38206;
	wire [4-1:0] node38207;
	wire [4-1:0] node38209;
	wire [4-1:0] node38212;
	wire [4-1:0] node38214;
	wire [4-1:0] node38217;
	wire [4-1:0] node38218;
	wire [4-1:0] node38219;
	wire [4-1:0] node38220;
	wire [4-1:0] node38222;
	wire [4-1:0] node38226;
	wire [4-1:0] node38227;
	wire [4-1:0] node38229;
	wire [4-1:0] node38232;
	wire [4-1:0] node38234;
	wire [4-1:0] node38237;
	wire [4-1:0] node38238;
	wire [4-1:0] node38240;
	wire [4-1:0] node38241;
	wire [4-1:0] node38244;
	wire [4-1:0] node38247;
	wire [4-1:0] node38248;
	wire [4-1:0] node38250;
	wire [4-1:0] node38253;
	wire [4-1:0] node38254;
	wire [4-1:0] node38257;
	wire [4-1:0] node38260;
	wire [4-1:0] node38261;
	wire [4-1:0] node38262;
	wire [4-1:0] node38263;
	wire [4-1:0] node38264;
	wire [4-1:0] node38265;
	wire [4-1:0] node38268;
	wire [4-1:0] node38271;
	wire [4-1:0] node38272;
	wire [4-1:0] node38275;
	wire [4-1:0] node38278;
	wire [4-1:0] node38279;
	wire [4-1:0] node38280;
	wire [4-1:0] node38283;
	wire [4-1:0] node38287;
	wire [4-1:0] node38288;
	wire [4-1:0] node38289;
	wire [4-1:0] node38290;
	wire [4-1:0] node38292;
	wire [4-1:0] node38295;
	wire [4-1:0] node38297;
	wire [4-1:0] node38300;
	wire [4-1:0] node38302;
	wire [4-1:0] node38303;
	wire [4-1:0] node38306;
	wire [4-1:0] node38309;
	wire [4-1:0] node38310;
	wire [4-1:0] node38311;
	wire [4-1:0] node38313;
	wire [4-1:0] node38316;
	wire [4-1:0] node38318;
	wire [4-1:0] node38321;
	wire [4-1:0] node38322;
	wire [4-1:0] node38325;
	wire [4-1:0] node38327;
	wire [4-1:0] node38330;
	wire [4-1:0] node38331;
	wire [4-1:0] node38332;
	wire [4-1:0] node38333;
	wire [4-1:0] node38334;
	wire [4-1:0] node38336;
	wire [4-1:0] node38339;
	wire [4-1:0] node38343;
	wire [4-1:0] node38344;
	wire [4-1:0] node38345;
	wire [4-1:0] node38348;
	wire [4-1:0] node38351;
	wire [4-1:0] node38352;
	wire [4-1:0] node38353;
	wire [4-1:0] node38356;
	wire [4-1:0] node38360;
	wire [4-1:0] node38361;
	wire [4-1:0] node38362;
	wire [4-1:0] node38364;
	wire [4-1:0] node38368;
	wire [4-1:0] node38369;
	wire [4-1:0] node38372;
	wire [4-1:0] node38374;
	wire [4-1:0] node38377;
	wire [4-1:0] node38378;
	wire [4-1:0] node38379;
	wire [4-1:0] node38380;
	wire [4-1:0] node38381;
	wire [4-1:0] node38382;
	wire [4-1:0] node38383;
	wire [4-1:0] node38384;
	wire [4-1:0] node38385;
	wire [4-1:0] node38388;
	wire [4-1:0] node38392;
	wire [4-1:0] node38393;
	wire [4-1:0] node38394;
	wire [4-1:0] node38397;
	wire [4-1:0] node38400;
	wire [4-1:0] node38401;
	wire [4-1:0] node38404;
	wire [4-1:0] node38407;
	wire [4-1:0] node38408;
	wire [4-1:0] node38409;
	wire [4-1:0] node38412;
	wire [4-1:0] node38414;
	wire [4-1:0] node38417;
	wire [4-1:0] node38418;
	wire [4-1:0] node38420;
	wire [4-1:0] node38423;
	wire [4-1:0] node38425;
	wire [4-1:0] node38428;
	wire [4-1:0] node38429;
	wire [4-1:0] node38430;
	wire [4-1:0] node38431;
	wire [4-1:0] node38432;
	wire [4-1:0] node38435;
	wire [4-1:0] node38438;
	wire [4-1:0] node38439;
	wire [4-1:0] node38442;
	wire [4-1:0] node38445;
	wire [4-1:0] node38446;
	wire [4-1:0] node38447;
	wire [4-1:0] node38448;
	wire [4-1:0] node38451;
	wire [4-1:0] node38454;
	wire [4-1:0] node38455;
	wire [4-1:0] node38458;
	wire [4-1:0] node38461;
	wire [4-1:0] node38463;
	wire [4-1:0] node38466;
	wire [4-1:0] node38467;
	wire [4-1:0] node38468;
	wire [4-1:0] node38469;
	wire [4-1:0] node38474;
	wire [4-1:0] node38475;
	wire [4-1:0] node38476;
	wire [4-1:0] node38480;
	wire [4-1:0] node38481;
	wire [4-1:0] node38485;
	wire [4-1:0] node38486;
	wire [4-1:0] node38487;
	wire [4-1:0] node38488;
	wire [4-1:0] node38489;
	wire [4-1:0] node38490;
	wire [4-1:0] node38493;
	wire [4-1:0] node38495;
	wire [4-1:0] node38498;
	wire [4-1:0] node38499;
	wire [4-1:0] node38502;
	wire [4-1:0] node38504;
	wire [4-1:0] node38507;
	wire [4-1:0] node38508;
	wire [4-1:0] node38509;
	wire [4-1:0] node38512;
	wire [4-1:0] node38515;
	wire [4-1:0] node38516;
	wire [4-1:0] node38519;
	wire [4-1:0] node38521;
	wire [4-1:0] node38524;
	wire [4-1:0] node38525;
	wire [4-1:0] node38526;
	wire [4-1:0] node38527;
	wire [4-1:0] node38530;
	wire [4-1:0] node38531;
	wire [4-1:0] node38534;
	wire [4-1:0] node38537;
	wire [4-1:0] node38538;
	wire [4-1:0] node38541;
	wire [4-1:0] node38544;
	wire [4-1:0] node38545;
	wire [4-1:0] node38546;
	wire [4-1:0] node38547;
	wire [4-1:0] node38550;
	wire [4-1:0] node38553;
	wire [4-1:0] node38556;
	wire [4-1:0] node38557;
	wire [4-1:0] node38558;
	wire [4-1:0] node38563;
	wire [4-1:0] node38564;
	wire [4-1:0] node38565;
	wire [4-1:0] node38566;
	wire [4-1:0] node38568;
	wire [4-1:0] node38571;
	wire [4-1:0] node38572;
	wire [4-1:0] node38573;
	wire [4-1:0] node38576;
	wire [4-1:0] node38579;
	wire [4-1:0] node38580;
	wire [4-1:0] node38583;
	wire [4-1:0] node38586;
	wire [4-1:0] node38587;
	wire [4-1:0] node38588;
	wire [4-1:0] node38592;
	wire [4-1:0] node38593;
	wire [4-1:0] node38596;
	wire [4-1:0] node38599;
	wire [4-1:0] node38600;
	wire [4-1:0] node38601;
	wire [4-1:0] node38602;
	wire [4-1:0] node38603;
	wire [4-1:0] node38606;
	wire [4-1:0] node38609;
	wire [4-1:0] node38610;
	wire [4-1:0] node38614;
	wire [4-1:0] node38615;
	wire [4-1:0] node38616;
	wire [4-1:0] node38619;
	wire [4-1:0] node38622;
	wire [4-1:0] node38623;
	wire [4-1:0] node38626;
	wire [4-1:0] node38629;
	wire [4-1:0] node38630;
	wire [4-1:0] node38631;
	wire [4-1:0] node38632;
	wire [4-1:0] node38636;
	wire [4-1:0] node38639;
	wire [4-1:0] node38641;
	wire [4-1:0] node38644;
	wire [4-1:0] node38645;
	wire [4-1:0] node38646;
	wire [4-1:0] node38647;
	wire [4-1:0] node38648;
	wire [4-1:0] node38649;
	wire [4-1:0] node38650;
	wire [4-1:0] node38652;
	wire [4-1:0] node38655;
	wire [4-1:0] node38657;
	wire [4-1:0] node38660;
	wire [4-1:0] node38661;
	wire [4-1:0] node38662;
	wire [4-1:0] node38665;
	wire [4-1:0] node38669;
	wire [4-1:0] node38670;
	wire [4-1:0] node38671;
	wire [4-1:0] node38672;
	wire [4-1:0] node38676;
	wire [4-1:0] node38677;
	wire [4-1:0] node38680;
	wire [4-1:0] node38683;
	wire [4-1:0] node38684;
	wire [4-1:0] node38685;
	wire [4-1:0] node38688;
	wire [4-1:0] node38691;
	wire [4-1:0] node38693;
	wire [4-1:0] node38696;
	wire [4-1:0] node38697;
	wire [4-1:0] node38698;
	wire [4-1:0] node38700;
	wire [4-1:0] node38703;
	wire [4-1:0] node38704;
	wire [4-1:0] node38706;
	wire [4-1:0] node38709;
	wire [4-1:0] node38711;
	wire [4-1:0] node38714;
	wire [4-1:0] node38715;
	wire [4-1:0] node38716;
	wire [4-1:0] node38719;
	wire [4-1:0] node38722;
	wire [4-1:0] node38724;
	wire [4-1:0] node38727;
	wire [4-1:0] node38728;
	wire [4-1:0] node38729;
	wire [4-1:0] node38730;
	wire [4-1:0] node38731;
	wire [4-1:0] node38732;
	wire [4-1:0] node38735;
	wire [4-1:0] node38739;
	wire [4-1:0] node38740;
	wire [4-1:0] node38741;
	wire [4-1:0] node38744;
	wire [4-1:0] node38747;
	wire [4-1:0] node38750;
	wire [4-1:0] node38751;
	wire [4-1:0] node38752;
	wire [4-1:0] node38753;
	wire [4-1:0] node38756;
	wire [4-1:0] node38759;
	wire [4-1:0] node38761;
	wire [4-1:0] node38764;
	wire [4-1:0] node38765;
	wire [4-1:0] node38767;
	wire [4-1:0] node38771;
	wire [4-1:0] node38772;
	wire [4-1:0] node38774;
	wire [4-1:0] node38775;
	wire [4-1:0] node38776;
	wire [4-1:0] node38779;
	wire [4-1:0] node38782;
	wire [4-1:0] node38784;
	wire [4-1:0] node38787;
	wire [4-1:0] node38788;
	wire [4-1:0] node38789;
	wire [4-1:0] node38790;
	wire [4-1:0] node38793;
	wire [4-1:0] node38797;
	wire [4-1:0] node38799;
	wire [4-1:0] node38802;
	wire [4-1:0] node38803;
	wire [4-1:0] node38804;
	wire [4-1:0] node38805;
	wire [4-1:0] node38806;
	wire [4-1:0] node38809;
	wire [4-1:0] node38811;
	wire [4-1:0] node38814;
	wire [4-1:0] node38815;
	wire [4-1:0] node38817;
	wire [4-1:0] node38820;
	wire [4-1:0] node38823;
	wire [4-1:0] node38824;
	wire [4-1:0] node38825;
	wire [4-1:0] node38826;
	wire [4-1:0] node38829;
	wire [4-1:0] node38832;
	wire [4-1:0] node38833;
	wire [4-1:0] node38837;
	wire [4-1:0] node38838;
	wire [4-1:0] node38839;
	wire [4-1:0] node38842;
	wire [4-1:0] node38845;
	wire [4-1:0] node38846;
	wire [4-1:0] node38849;
	wire [4-1:0] node38852;
	wire [4-1:0] node38853;
	wire [4-1:0] node38854;
	wire [4-1:0] node38855;
	wire [4-1:0] node38856;
	wire [4-1:0] node38859;
	wire [4-1:0] node38862;
	wire [4-1:0] node38863;
	wire [4-1:0] node38866;
	wire [4-1:0] node38869;
	wire [4-1:0] node38870;
	wire [4-1:0] node38871;
	wire [4-1:0] node38874;
	wire [4-1:0] node38877;
	wire [4-1:0] node38878;
	wire [4-1:0] node38879;
	wire [4-1:0] node38882;
	wire [4-1:0] node38886;
	wire [4-1:0] node38887;
	wire [4-1:0] node38888;
	wire [4-1:0] node38889;
	wire [4-1:0] node38891;
	wire [4-1:0] node38894;
	wire [4-1:0] node38895;
	wire [4-1:0] node38898;
	wire [4-1:0] node38901;
	wire [4-1:0] node38902;
	wire [4-1:0] node38905;
	wire [4-1:0] node38908;
	wire [4-1:0] node38909;
	wire [4-1:0] node38912;
	wire [4-1:0] node38915;
	wire [4-1:0] node38916;
	wire [4-1:0] node38917;
	wire [4-1:0] node38918;
	wire [4-1:0] node38919;
	wire [4-1:0] node38920;
	wire [4-1:0] node38921;
	wire [4-1:0] node38922;
	wire [4-1:0] node38926;
	wire [4-1:0] node38928;
	wire [4-1:0] node38931;
	wire [4-1:0] node38932;
	wire [4-1:0] node38933;
	wire [4-1:0] node38936;
	wire [4-1:0] node38939;
	wire [4-1:0] node38940;
	wire [4-1:0] node38943;
	wire [4-1:0] node38946;
	wire [4-1:0] node38947;
	wire [4-1:0] node38948;
	wire [4-1:0] node38949;
	wire [4-1:0] node38952;
	wire [4-1:0] node38955;
	wire [4-1:0] node38956;
	wire [4-1:0] node38959;
	wire [4-1:0] node38962;
	wire [4-1:0] node38963;
	wire [4-1:0] node38964;
	wire [4-1:0] node38968;
	wire [4-1:0] node38970;
	wire [4-1:0] node38972;
	wire [4-1:0] node38975;
	wire [4-1:0] node38976;
	wire [4-1:0] node38977;
	wire [4-1:0] node38978;
	wire [4-1:0] node38979;
	wire [4-1:0] node38980;
	wire [4-1:0] node38984;
	wire [4-1:0] node38985;
	wire [4-1:0] node38988;
	wire [4-1:0] node38991;
	wire [4-1:0] node38992;
	wire [4-1:0] node38994;
	wire [4-1:0] node38997;
	wire [4-1:0] node38998;
	wire [4-1:0] node39001;
	wire [4-1:0] node39004;
	wire [4-1:0] node39005;
	wire [4-1:0] node39006;
	wire [4-1:0] node39008;
	wire [4-1:0] node39011;
	wire [4-1:0] node39014;
	wire [4-1:0] node39015;
	wire [4-1:0] node39017;
	wire [4-1:0] node39020;
	wire [4-1:0] node39021;
	wire [4-1:0] node39025;
	wire [4-1:0] node39026;
	wire [4-1:0] node39027;
	wire [4-1:0] node39028;
	wire [4-1:0] node39031;
	wire [4-1:0] node39034;
	wire [4-1:0] node39035;
	wire [4-1:0] node39038;
	wire [4-1:0] node39041;
	wire [4-1:0] node39042;
	wire [4-1:0] node39044;
	wire [4-1:0] node39047;
	wire [4-1:0] node39048;
	wire [4-1:0] node39050;
	wire [4-1:0] node39054;
	wire [4-1:0] node39055;
	wire [4-1:0] node39056;
	wire [4-1:0] node39057;
	wire [4-1:0] node39058;
	wire [4-1:0] node39059;
	wire [4-1:0] node39062;
	wire [4-1:0] node39065;
	wire [4-1:0] node39067;
	wire [4-1:0] node39070;
	wire [4-1:0] node39071;
	wire [4-1:0] node39072;
	wire [4-1:0] node39075;
	wire [4-1:0] node39078;
	wire [4-1:0] node39079;
	wire [4-1:0] node39082;
	wire [4-1:0] node39085;
	wire [4-1:0] node39086;
	wire [4-1:0] node39087;
	wire [4-1:0] node39088;
	wire [4-1:0] node39091;
	wire [4-1:0] node39094;
	wire [4-1:0] node39096;
	wire [4-1:0] node39097;
	wire [4-1:0] node39100;
	wire [4-1:0] node39103;
	wire [4-1:0] node39104;
	wire [4-1:0] node39105;
	wire [4-1:0] node39107;
	wire [4-1:0] node39110;
	wire [4-1:0] node39111;
	wire [4-1:0] node39114;
	wire [4-1:0] node39118;
	wire [4-1:0] node39119;
	wire [4-1:0] node39120;
	wire [4-1:0] node39121;
	wire [4-1:0] node39122;
	wire [4-1:0] node39125;
	wire [4-1:0] node39128;
	wire [4-1:0] node39129;
	wire [4-1:0] node39131;
	wire [4-1:0] node39134;
	wire [4-1:0] node39135;
	wire [4-1:0] node39139;
	wire [4-1:0] node39140;
	wire [4-1:0] node39141;
	wire [4-1:0] node39144;
	wire [4-1:0] node39147;
	wire [4-1:0] node39148;
	wire [4-1:0] node39149;
	wire [4-1:0] node39152;
	wire [4-1:0] node39155;
	wire [4-1:0] node39156;
	wire [4-1:0] node39159;
	wire [4-1:0] node39162;
	wire [4-1:0] node39163;
	wire [4-1:0] node39164;
	wire [4-1:0] node39165;
	wire [4-1:0] node39168;
	wire [4-1:0] node39171;
	wire [4-1:0] node39172;
	wire [4-1:0] node39175;
	wire [4-1:0] node39178;
	wire [4-1:0] node39179;
	wire [4-1:0] node39181;
	wire [4-1:0] node39184;
	wire [4-1:0] node39185;
	wire [4-1:0] node39188;
	wire [4-1:0] node39191;
	wire [4-1:0] node39192;
	wire [4-1:0] node39193;
	wire [4-1:0] node39194;
	wire [4-1:0] node39195;
	wire [4-1:0] node39198;
	wire [4-1:0] node39201;
	wire [4-1:0] node39202;
	wire [4-1:0] node39203;
	wire [4-1:0] node39204;
	wire [4-1:0] node39205;
	wire [4-1:0] node39208;
	wire [4-1:0] node39212;
	wire [4-1:0] node39213;
	wire [4-1:0] node39216;
	wire [4-1:0] node39219;
	wire [4-1:0] node39220;
	wire [4-1:0] node39222;
	wire [4-1:0] node39224;
	wire [4-1:0] node39227;
	wire [4-1:0] node39228;
	wire [4-1:0] node39229;
	wire [4-1:0] node39232;
	wire [4-1:0] node39235;
	wire [4-1:0] node39237;
	wire [4-1:0] node39240;
	wire [4-1:0] node39241;
	wire [4-1:0] node39242;
	wire [4-1:0] node39243;
	wire [4-1:0] node39245;
	wire [4-1:0] node39248;
	wire [4-1:0] node39249;
	wire [4-1:0] node39250;
	wire [4-1:0] node39254;
	wire [4-1:0] node39255;
	wire [4-1:0] node39259;
	wire [4-1:0] node39260;
	wire [4-1:0] node39261;
	wire [4-1:0] node39262;
	wire [4-1:0] node39265;
	wire [4-1:0] node39268;
	wire [4-1:0] node39269;
	wire [4-1:0] node39273;
	wire [4-1:0] node39275;
	wire [4-1:0] node39276;
	wire [4-1:0] node39279;
	wire [4-1:0] node39282;
	wire [4-1:0] node39283;
	wire [4-1:0] node39285;
	wire [4-1:0] node39286;
	wire [4-1:0] node39287;
	wire [4-1:0] node39290;
	wire [4-1:0] node39294;
	wire [4-1:0] node39295;
	wire [4-1:0] node39296;
	wire [4-1:0] node39300;
	wire [4-1:0] node39301;
	wire [4-1:0] node39304;
	wire [4-1:0] node39307;
	wire [4-1:0] node39308;
	wire [4-1:0] node39309;
	wire [4-1:0] node39310;
	wire [4-1:0] node39311;
	wire [4-1:0] node39312;
	wire [4-1:0] node39316;
	wire [4-1:0] node39317;
	wire [4-1:0] node39321;
	wire [4-1:0] node39322;
	wire [4-1:0] node39323;
	wire [4-1:0] node39324;
	wire [4-1:0] node39327;
	wire [4-1:0] node39330;
	wire [4-1:0] node39331;
	wire [4-1:0] node39336;
	wire [4-1:0] node39337;
	wire [4-1:0] node39338;
	wire [4-1:0] node39339;
	wire [4-1:0] node39342;
	wire [4-1:0] node39345;
	wire [4-1:0] node39347;
	wire [4-1:0] node39350;
	wire [4-1:0] node39351;
	wire [4-1:0] node39354;
	wire [4-1:0] node39357;
	wire [4-1:0] node39358;
	wire [4-1:0] node39359;
	wire [4-1:0] node39361;
	wire [4-1:0] node39362;
	wire [4-1:0] node39363;
	wire [4-1:0] node39366;
	wire [4-1:0] node39369;
	wire [4-1:0] node39371;
	wire [4-1:0] node39374;
	wire [4-1:0] node39375;
	wire [4-1:0] node39376;
	wire [4-1:0] node39379;
	wire [4-1:0] node39382;
	wire [4-1:0] node39383;
	wire [4-1:0] node39385;
	wire [4-1:0] node39388;
	wire [4-1:0] node39389;
	wire [4-1:0] node39392;
	wire [4-1:0] node39395;
	wire [4-1:0] node39396;
	wire [4-1:0] node39397;
	wire [4-1:0] node39398;
	wire [4-1:0] node39402;
	wire [4-1:0] node39403;
	wire [4-1:0] node39407;
	wire [4-1:0] node39408;
	wire [4-1:0] node39411;
	wire [4-1:0] node39412;
	wire [4-1:0] node39416;
	wire [4-1:0] node39417;
	wire [4-1:0] node39418;
	wire [4-1:0] node39419;
	wire [4-1:0] node39420;
	wire [4-1:0] node39421;
	wire [4-1:0] node39422;
	wire [4-1:0] node39423;
	wire [4-1:0] node39424;
	wire [4-1:0] node39425;
	wire [4-1:0] node39428;
	wire [4-1:0] node39431;
	wire [4-1:0] node39434;
	wire [4-1:0] node39435;
	wire [4-1:0] node39436;
	wire [4-1:0] node39439;
	wire [4-1:0] node39442;
	wire [4-1:0] node39443;
	wire [4-1:0] node39446;
	wire [4-1:0] node39449;
	wire [4-1:0] node39450;
	wire [4-1:0] node39451;
	wire [4-1:0] node39452;
	wire [4-1:0] node39455;
	wire [4-1:0] node39458;
	wire [4-1:0] node39459;
	wire [4-1:0] node39460;
	wire [4-1:0] node39463;
	wire [4-1:0] node39466;
	wire [4-1:0] node39467;
	wire [4-1:0] node39470;
	wire [4-1:0] node39473;
	wire [4-1:0] node39474;
	wire [4-1:0] node39475;
	wire [4-1:0] node39476;
	wire [4-1:0] node39479;
	wire [4-1:0] node39482;
	wire [4-1:0] node39483;
	wire [4-1:0] node39486;
	wire [4-1:0] node39489;
	wire [4-1:0] node39490;
	wire [4-1:0] node39493;
	wire [4-1:0] node39496;
	wire [4-1:0] node39497;
	wire [4-1:0] node39498;
	wire [4-1:0] node39499;
	wire [4-1:0] node39500;
	wire [4-1:0] node39501;
	wire [4-1:0] node39504;
	wire [4-1:0] node39507;
	wire [4-1:0] node39508;
	wire [4-1:0] node39512;
	wire [4-1:0] node39513;
	wire [4-1:0] node39516;
	wire [4-1:0] node39518;
	wire [4-1:0] node39521;
	wire [4-1:0] node39522;
	wire [4-1:0] node39523;
	wire [4-1:0] node39524;
	wire [4-1:0] node39529;
	wire [4-1:0] node39530;
	wire [4-1:0] node39531;
	wire [4-1:0] node39535;
	wire [4-1:0] node39536;
	wire [4-1:0] node39540;
	wire [4-1:0] node39541;
	wire [4-1:0] node39542;
	wire [4-1:0] node39543;
	wire [4-1:0] node39544;
	wire [4-1:0] node39547;
	wire [4-1:0] node39550;
	wire [4-1:0] node39551;
	wire [4-1:0] node39555;
	wire [4-1:0] node39556;
	wire [4-1:0] node39558;
	wire [4-1:0] node39562;
	wire [4-1:0] node39563;
	wire [4-1:0] node39564;
	wire [4-1:0] node39565;
	wire [4-1:0] node39568;
	wire [4-1:0] node39571;
	wire [4-1:0] node39572;
	wire [4-1:0] node39575;
	wire [4-1:0] node39578;
	wire [4-1:0] node39579;
	wire [4-1:0] node39582;
	wire [4-1:0] node39585;
	wire [4-1:0] node39586;
	wire [4-1:0] node39587;
	wire [4-1:0] node39588;
	wire [4-1:0] node39589;
	wire [4-1:0] node39591;
	wire [4-1:0] node39594;
	wire [4-1:0] node39595;
	wire [4-1:0] node39596;
	wire [4-1:0] node39599;
	wire [4-1:0] node39602;
	wire [4-1:0] node39603;
	wire [4-1:0] node39606;
	wire [4-1:0] node39609;
	wire [4-1:0] node39610;
	wire [4-1:0] node39611;
	wire [4-1:0] node39614;
	wire [4-1:0] node39617;
	wire [4-1:0] node39618;
	wire [4-1:0] node39619;
	wire [4-1:0] node39622;
	wire [4-1:0] node39625;
	wire [4-1:0] node39626;
	wire [4-1:0] node39630;
	wire [4-1:0] node39631;
	wire [4-1:0] node39632;
	wire [4-1:0] node39633;
	wire [4-1:0] node39636;
	wire [4-1:0] node39637;
	wire [4-1:0] node39641;
	wire [4-1:0] node39642;
	wire [4-1:0] node39645;
	wire [4-1:0] node39648;
	wire [4-1:0] node39649;
	wire [4-1:0] node39650;
	wire [4-1:0] node39651;
	wire [4-1:0] node39655;
	wire [4-1:0] node39656;
	wire [4-1:0] node39659;
	wire [4-1:0] node39662;
	wire [4-1:0] node39663;
	wire [4-1:0] node39664;
	wire [4-1:0] node39668;
	wire [4-1:0] node39671;
	wire [4-1:0] node39672;
	wire [4-1:0] node39673;
	wire [4-1:0] node39674;
	wire [4-1:0] node39675;
	wire [4-1:0] node39678;
	wire [4-1:0] node39680;
	wire [4-1:0] node39684;
	wire [4-1:0] node39685;
	wire [4-1:0] node39686;
	wire [4-1:0] node39687;
	wire [4-1:0] node39690;
	wire [4-1:0] node39694;
	wire [4-1:0] node39695;
	wire [4-1:0] node39697;
	wire [4-1:0] node39700;
	wire [4-1:0] node39701;
	wire [4-1:0] node39704;
	wire [4-1:0] node39707;
	wire [4-1:0] node39708;
	wire [4-1:0] node39709;
	wire [4-1:0] node39710;
	wire [4-1:0] node39711;
	wire [4-1:0] node39714;
	wire [4-1:0] node39717;
	wire [4-1:0] node39718;
	wire [4-1:0] node39721;
	wire [4-1:0] node39724;
	wire [4-1:0] node39725;
	wire [4-1:0] node39726;
	wire [4-1:0] node39730;
	wire [4-1:0] node39732;
	wire [4-1:0] node39735;
	wire [4-1:0] node39736;
	wire [4-1:0] node39737;
	wire [4-1:0] node39738;
	wire [4-1:0] node39742;
	wire [4-1:0] node39743;
	wire [4-1:0] node39746;
	wire [4-1:0] node39749;
	wire [4-1:0] node39751;
	wire [4-1:0] node39754;
	wire [4-1:0] node39755;
	wire [4-1:0] node39756;
	wire [4-1:0] node39757;
	wire [4-1:0] node39758;
	wire [4-1:0] node39759;
	wire [4-1:0] node39760;
	wire [4-1:0] node39761;
	wire [4-1:0] node39764;
	wire [4-1:0] node39767;
	wire [4-1:0] node39768;
	wire [4-1:0] node39773;
	wire [4-1:0] node39774;
	wire [4-1:0] node39775;
	wire [4-1:0] node39776;
	wire [4-1:0] node39780;
	wire [4-1:0] node39781;
	wire [4-1:0] node39785;
	wire [4-1:0] node39786;
	wire [4-1:0] node39789;
	wire [4-1:0] node39792;
	wire [4-1:0] node39793;
	wire [4-1:0] node39794;
	wire [4-1:0] node39795;
	wire [4-1:0] node39798;
	wire [4-1:0] node39801;
	wire [4-1:0] node39802;
	wire [4-1:0] node39806;
	wire [4-1:0] node39807;
	wire [4-1:0] node39808;
	wire [4-1:0] node39812;
	wire [4-1:0] node39813;
	wire [4-1:0] node39817;
	wire [4-1:0] node39818;
	wire [4-1:0] node39819;
	wire [4-1:0] node39820;
	wire [4-1:0] node39821;
	wire [4-1:0] node39823;
	wire [4-1:0] node39826;
	wire [4-1:0] node39827;
	wire [4-1:0] node39831;
	wire [4-1:0] node39832;
	wire [4-1:0] node39834;
	wire [4-1:0] node39837;
	wire [4-1:0] node39840;
	wire [4-1:0] node39841;
	wire [4-1:0] node39843;
	wire [4-1:0] node39846;
	wire [4-1:0] node39847;
	wire [4-1:0] node39848;
	wire [4-1:0] node39853;
	wire [4-1:0] node39854;
	wire [4-1:0] node39855;
	wire [4-1:0] node39856;
	wire [4-1:0] node39859;
	wire [4-1:0] node39862;
	wire [4-1:0] node39865;
	wire [4-1:0] node39866;
	wire [4-1:0] node39867;
	wire [4-1:0] node39871;
	wire [4-1:0] node39872;
	wire [4-1:0] node39876;
	wire [4-1:0] node39877;
	wire [4-1:0] node39878;
	wire [4-1:0] node39879;
	wire [4-1:0] node39880;
	wire [4-1:0] node39881;
	wire [4-1:0] node39885;
	wire [4-1:0] node39886;
	wire [4-1:0] node39889;
	wire [4-1:0] node39892;
	wire [4-1:0] node39893;
	wire [4-1:0] node39894;
	wire [4-1:0] node39897;
	wire [4-1:0] node39900;
	wire [4-1:0] node39901;
	wire [4-1:0] node39904;
	wire [4-1:0] node39907;
	wire [4-1:0] node39908;
	wire [4-1:0] node39909;
	wire [4-1:0] node39910;
	wire [4-1:0] node39913;
	wire [4-1:0] node39914;
	wire [4-1:0] node39918;
	wire [4-1:0] node39919;
	wire [4-1:0] node39920;
	wire [4-1:0] node39924;
	wire [4-1:0] node39925;
	wire [4-1:0] node39929;
	wire [4-1:0] node39930;
	wire [4-1:0] node39931;
	wire [4-1:0] node39932;
	wire [4-1:0] node39935;
	wire [4-1:0] node39939;
	wire [4-1:0] node39940;
	wire [4-1:0] node39941;
	wire [4-1:0] node39944;
	wire [4-1:0] node39947;
	wire [4-1:0] node39948;
	wire [4-1:0] node39951;
	wire [4-1:0] node39954;
	wire [4-1:0] node39955;
	wire [4-1:0] node39956;
	wire [4-1:0] node39957;
	wire [4-1:0] node39958;
	wire [4-1:0] node39959;
	wire [4-1:0] node39964;
	wire [4-1:0] node39965;
	wire [4-1:0] node39966;
	wire [4-1:0] node39971;
	wire [4-1:0] node39972;
	wire [4-1:0] node39973;
	wire [4-1:0] node39974;
	wire [4-1:0] node39978;
	wire [4-1:0] node39979;
	wire [4-1:0] node39983;
	wire [4-1:0] node39984;
	wire [4-1:0] node39986;
	wire [4-1:0] node39989;
	wire [4-1:0] node39991;
	wire [4-1:0] node39994;
	wire [4-1:0] node39995;
	wire [4-1:0] node39996;
	wire [4-1:0] node39998;
	wire [4-1:0] node40001;
	wire [4-1:0] node40002;
	wire [4-1:0] node40005;
	wire [4-1:0] node40008;
	wire [4-1:0] node40009;
	wire [4-1:0] node40010;
	wire [4-1:0] node40011;
	wire [4-1:0] node40014;
	wire [4-1:0] node40018;
	wire [4-1:0] node40019;
	wire [4-1:0] node40023;
	wire [4-1:0] node40024;
	wire [4-1:0] node40025;
	wire [4-1:0] node40026;
	wire [4-1:0] node40027;
	wire [4-1:0] node40028;
	wire [4-1:0] node40029;
	wire [4-1:0] node40031;
	wire [4-1:0] node40032;
	wire [4-1:0] node40035;
	wire [4-1:0] node40038;
	wire [4-1:0] node40040;
	wire [4-1:0] node40043;
	wire [4-1:0] node40044;
	wire [4-1:0] node40045;
	wire [4-1:0] node40048;
	wire [4-1:0] node40051;
	wire [4-1:0] node40052;
	wire [4-1:0] node40055;
	wire [4-1:0] node40058;
	wire [4-1:0] node40059;
	wire [4-1:0] node40060;
	wire [4-1:0] node40062;
	wire [4-1:0] node40065;
	wire [4-1:0] node40066;
	wire [4-1:0] node40067;
	wire [4-1:0] node40070;
	wire [4-1:0] node40074;
	wire [4-1:0] node40075;
	wire [4-1:0] node40077;
	wire [4-1:0] node40080;
	wire [4-1:0] node40081;
	wire [4-1:0] node40084;
	wire [4-1:0] node40087;
	wire [4-1:0] node40088;
	wire [4-1:0] node40089;
	wire [4-1:0] node40090;
	wire [4-1:0] node40091;
	wire [4-1:0] node40092;
	wire [4-1:0] node40095;
	wire [4-1:0] node40098;
	wire [4-1:0] node40099;
	wire [4-1:0] node40103;
	wire [4-1:0] node40104;
	wire [4-1:0] node40106;
	wire [4-1:0] node40109;
	wire [4-1:0] node40110;
	wire [4-1:0] node40114;
	wire [4-1:0] node40115;
	wire [4-1:0] node40116;
	wire [4-1:0] node40119;
	wire [4-1:0] node40122;
	wire [4-1:0] node40123;
	wire [4-1:0] node40125;
	wire [4-1:0] node40128;
	wire [4-1:0] node40130;
	wire [4-1:0] node40133;
	wire [4-1:0] node40134;
	wire [4-1:0] node40135;
	wire [4-1:0] node40136;
	wire [4-1:0] node40139;
	wire [4-1:0] node40142;
	wire [4-1:0] node40143;
	wire [4-1:0] node40147;
	wire [4-1:0] node40148;
	wire [4-1:0] node40150;
	wire [4-1:0] node40151;
	wire [4-1:0] node40155;
	wire [4-1:0] node40157;
	wire [4-1:0] node40160;
	wire [4-1:0] node40161;
	wire [4-1:0] node40162;
	wire [4-1:0] node40163;
	wire [4-1:0] node40164;
	wire [4-1:0] node40165;
	wire [4-1:0] node40168;
	wire [4-1:0] node40171;
	wire [4-1:0] node40172;
	wire [4-1:0] node40175;
	wire [4-1:0] node40178;
	wire [4-1:0] node40179;
	wire [4-1:0] node40180;
	wire [4-1:0] node40184;
	wire [4-1:0] node40186;
	wire [4-1:0] node40187;
	wire [4-1:0] node40190;
	wire [4-1:0] node40193;
	wire [4-1:0] node40194;
	wire [4-1:0] node40195;
	wire [4-1:0] node40196;
	wire [4-1:0] node40197;
	wire [4-1:0] node40200;
	wire [4-1:0] node40203;
	wire [4-1:0] node40205;
	wire [4-1:0] node40208;
	wire [4-1:0] node40209;
	wire [4-1:0] node40212;
	wire [4-1:0] node40215;
	wire [4-1:0] node40216;
	wire [4-1:0] node40219;
	wire [4-1:0] node40222;
	wire [4-1:0] node40223;
	wire [4-1:0] node40224;
	wire [4-1:0] node40225;
	wire [4-1:0] node40226;
	wire [4-1:0] node40228;
	wire [4-1:0] node40231;
	wire [4-1:0] node40233;
	wire [4-1:0] node40236;
	wire [4-1:0] node40237;
	wire [4-1:0] node40238;
	wire [4-1:0] node40243;
	wire [4-1:0] node40244;
	wire [4-1:0] node40245;
	wire [4-1:0] node40246;
	wire [4-1:0] node40250;
	wire [4-1:0] node40251;
	wire [4-1:0] node40255;
	wire [4-1:0] node40256;
	wire [4-1:0] node40257;
	wire [4-1:0] node40260;
	wire [4-1:0] node40263;
	wire [4-1:0] node40264;
	wire [4-1:0] node40268;
	wire [4-1:0] node40269;
	wire [4-1:0] node40270;
	wire [4-1:0] node40272;
	wire [4-1:0] node40273;
	wire [4-1:0] node40277;
	wire [4-1:0] node40280;
	wire [4-1:0] node40281;
	wire [4-1:0] node40282;
	wire [4-1:0] node40285;
	wire [4-1:0] node40288;
	wire [4-1:0] node40289;
	wire [4-1:0] node40290;
	wire [4-1:0] node40293;
	wire [4-1:0] node40296;
	wire [4-1:0] node40297;
	wire [4-1:0] node40301;
	wire [4-1:0] node40302;
	wire [4-1:0] node40303;
	wire [4-1:0] node40304;
	wire [4-1:0] node40305;
	wire [4-1:0] node40306;
	wire [4-1:0] node40309;
	wire [4-1:0] node40310;
	wire [4-1:0] node40311;
	wire [4-1:0] node40314;
	wire [4-1:0] node40317;
	wire [4-1:0] node40318;
	wire [4-1:0] node40322;
	wire [4-1:0] node40323;
	wire [4-1:0] node40325;
	wire [4-1:0] node40328;
	wire [4-1:0] node40329;
	wire [4-1:0] node40330;
	wire [4-1:0] node40333;
	wire [4-1:0] node40336;
	wire [4-1:0] node40338;
	wire [4-1:0] node40341;
	wire [4-1:0] node40342;
	wire [4-1:0] node40343;
	wire [4-1:0] node40344;
	wire [4-1:0] node40345;
	wire [4-1:0] node40348;
	wire [4-1:0] node40351;
	wire [4-1:0] node40352;
	wire [4-1:0] node40355;
	wire [4-1:0] node40358;
	wire [4-1:0] node40359;
	wire [4-1:0] node40360;
	wire [4-1:0] node40364;
	wire [4-1:0] node40365;
	wire [4-1:0] node40368;
	wire [4-1:0] node40371;
	wire [4-1:0] node40372;
	wire [4-1:0] node40373;
	wire [4-1:0] node40375;
	wire [4-1:0] node40378;
	wire [4-1:0] node40379;
	wire [4-1:0] node40382;
	wire [4-1:0] node40385;
	wire [4-1:0] node40386;
	wire [4-1:0] node40387;
	wire [4-1:0] node40390;
	wire [4-1:0] node40393;
	wire [4-1:0] node40396;
	wire [4-1:0] node40397;
	wire [4-1:0] node40398;
	wire [4-1:0] node40399;
	wire [4-1:0] node40400;
	wire [4-1:0] node40403;
	wire [4-1:0] node40405;
	wire [4-1:0] node40408;
	wire [4-1:0] node40409;
	wire [4-1:0] node40411;
	wire [4-1:0] node40415;
	wire [4-1:0] node40416;
	wire [4-1:0] node40417;
	wire [4-1:0] node40418;
	wire [4-1:0] node40421;
	wire [4-1:0] node40425;
	wire [4-1:0] node40426;
	wire [4-1:0] node40427;
	wire [4-1:0] node40430;
	wire [4-1:0] node40433;
	wire [4-1:0] node40434;
	wire [4-1:0] node40437;
	wire [4-1:0] node40440;
	wire [4-1:0] node40441;
	wire [4-1:0] node40442;
	wire [4-1:0] node40443;
	wire [4-1:0] node40444;
	wire [4-1:0] node40448;
	wire [4-1:0] node40449;
	wire [4-1:0] node40453;
	wire [4-1:0] node40454;
	wire [4-1:0] node40457;
	wire [4-1:0] node40458;
	wire [4-1:0] node40462;
	wire [4-1:0] node40463;
	wire [4-1:0] node40464;
	wire [4-1:0] node40465;
	wire [4-1:0] node40468;
	wire [4-1:0] node40472;
	wire [4-1:0] node40474;
	wire [4-1:0] node40477;
	wire [4-1:0] node40478;
	wire [4-1:0] node40479;
	wire [4-1:0] node40480;
	wire [4-1:0] node40481;
	wire [4-1:0] node40482;
	wire [4-1:0] node40485;
	wire [4-1:0] node40488;
	wire [4-1:0] node40489;
	wire [4-1:0] node40492;
	wire [4-1:0] node40495;
	wire [4-1:0] node40496;
	wire [4-1:0] node40497;
	wire [4-1:0] node40500;
	wire [4-1:0] node40503;
	wire [4-1:0] node40504;
	wire [4-1:0] node40507;
	wire [4-1:0] node40510;
	wire [4-1:0] node40511;
	wire [4-1:0] node40512;
	wire [4-1:0] node40513;
	wire [4-1:0] node40517;
	wire [4-1:0] node40518;
	wire [4-1:0] node40521;
	wire [4-1:0] node40524;
	wire [4-1:0] node40525;
	wire [4-1:0] node40526;
	wire [4-1:0] node40530;
	wire [4-1:0] node40533;
	wire [4-1:0] node40534;
	wire [4-1:0] node40535;
	wire [4-1:0] node40536;
	wire [4-1:0] node40538;
	wire [4-1:0] node40539;
	wire [4-1:0] node40542;
	wire [4-1:0] node40545;
	wire [4-1:0] node40546;
	wire [4-1:0] node40549;
	wire [4-1:0] node40552;
	wire [4-1:0] node40553;
	wire [4-1:0] node40554;
	wire [4-1:0] node40558;
	wire [4-1:0] node40561;
	wire [4-1:0] node40562;
	wire [4-1:0] node40563;
	wire [4-1:0] node40565;
	wire [4-1:0] node40568;
	wire [4-1:0] node40569;
	wire [4-1:0] node40572;
	wire [4-1:0] node40575;
	wire [4-1:0] node40576;
	wire [4-1:0] node40577;
	wire [4-1:0] node40581;
	wire [4-1:0] node40584;
	wire [4-1:0] node40585;
	wire [4-1:0] node40586;
	wire [4-1:0] node40587;
	wire [4-1:0] node40588;
	wire [4-1:0] node40589;
	wire [4-1:0] node40590;
	wire [4-1:0] node40591;
	wire [4-1:0] node40593;
	wire [4-1:0] node40594;
	wire [4-1:0] node40597;
	wire [4-1:0] node40600;
	wire [4-1:0] node40601;
	wire [4-1:0] node40602;
	wire [4-1:0] node40605;
	wire [4-1:0] node40608;
	wire [4-1:0] node40610;
	wire [4-1:0] node40613;
	wire [4-1:0] node40614;
	wire [4-1:0] node40615;
	wire [4-1:0] node40618;
	wire [4-1:0] node40621;
	wire [4-1:0] node40622;
	wire [4-1:0] node40623;
	wire [4-1:0] node40627;
	wire [4-1:0] node40628;
	wire [4-1:0] node40631;
	wire [4-1:0] node40634;
	wire [4-1:0] node40635;
	wire [4-1:0] node40636;
	wire [4-1:0] node40637;
	wire [4-1:0] node40638;
	wire [4-1:0] node40641;
	wire [4-1:0] node40644;
	wire [4-1:0] node40645;
	wire [4-1:0] node40649;
	wire [4-1:0] node40651;
	wire [4-1:0] node40653;
	wire [4-1:0] node40656;
	wire [4-1:0] node40657;
	wire [4-1:0] node40658;
	wire [4-1:0] node40661;
	wire [4-1:0] node40664;
	wire [4-1:0] node40665;
	wire [4-1:0] node40668;
	wire [4-1:0] node40670;
	wire [4-1:0] node40673;
	wire [4-1:0] node40674;
	wire [4-1:0] node40675;
	wire [4-1:0] node40676;
	wire [4-1:0] node40677;
	wire [4-1:0] node40680;
	wire [4-1:0] node40683;
	wire [4-1:0] node40685;
	wire [4-1:0] node40688;
	wire [4-1:0] node40689;
	wire [4-1:0] node40690;
	wire [4-1:0] node40694;
	wire [4-1:0] node40695;
	wire [4-1:0] node40696;
	wire [4-1:0] node40699;
	wire [4-1:0] node40702;
	wire [4-1:0] node40703;
	wire [4-1:0] node40706;
	wire [4-1:0] node40709;
	wire [4-1:0] node40710;
	wire [4-1:0] node40711;
	wire [4-1:0] node40712;
	wire [4-1:0] node40714;
	wire [4-1:0] node40717;
	wire [4-1:0] node40718;
	wire [4-1:0] node40722;
	wire [4-1:0] node40723;
	wire [4-1:0] node40726;
	wire [4-1:0] node40729;
	wire [4-1:0] node40730;
	wire [4-1:0] node40731;
	wire [4-1:0] node40732;
	wire [4-1:0] node40735;
	wire [4-1:0] node40738;
	wire [4-1:0] node40739;
	wire [4-1:0] node40742;
	wire [4-1:0] node40745;
	wire [4-1:0] node40746;
	wire [4-1:0] node40748;
	wire [4-1:0] node40751;
	wire [4-1:0] node40752;
	wire [4-1:0] node40755;
	wire [4-1:0] node40758;
	wire [4-1:0] node40759;
	wire [4-1:0] node40760;
	wire [4-1:0] node40761;
	wire [4-1:0] node40762;
	wire [4-1:0] node40763;
	wire [4-1:0] node40764;
	wire [4-1:0] node40768;
	wire [4-1:0] node40770;
	wire [4-1:0] node40773;
	wire [4-1:0] node40774;
	wire [4-1:0] node40777;
	wire [4-1:0] node40780;
	wire [4-1:0] node40781;
	wire [4-1:0] node40783;
	wire [4-1:0] node40786;
	wire [4-1:0] node40787;
	wire [4-1:0] node40790;
	wire [4-1:0] node40793;
	wire [4-1:0] node40794;
	wire [4-1:0] node40795;
	wire [4-1:0] node40796;
	wire [4-1:0] node40797;
	wire [4-1:0] node40800;
	wire [4-1:0] node40804;
	wire [4-1:0] node40805;
	wire [4-1:0] node40807;
	wire [4-1:0] node40810;
	wire [4-1:0] node40811;
	wire [4-1:0] node40814;
	wire [4-1:0] node40817;
	wire [4-1:0] node40818;
	wire [4-1:0] node40819;
	wire [4-1:0] node40822;
	wire [4-1:0] node40824;
	wire [4-1:0] node40827;
	wire [4-1:0] node40828;
	wire [4-1:0] node40831;
	wire [4-1:0] node40834;
	wire [4-1:0] node40835;
	wire [4-1:0] node40836;
	wire [4-1:0] node40837;
	wire [4-1:0] node40838;
	wire [4-1:0] node40842;
	wire [4-1:0] node40845;
	wire [4-1:0] node40846;
	wire [4-1:0] node40847;
	wire [4-1:0] node40851;
	wire [4-1:0] node40854;
	wire [4-1:0] node40855;
	wire [4-1:0] node40856;
	wire [4-1:0] node40857;
	wire [4-1:0] node40861;
	wire [4-1:0] node40864;
	wire [4-1:0] node40865;
	wire [4-1:0] node40866;
	wire [4-1:0] node40870;
	wire [4-1:0] node40873;
	wire [4-1:0] node40874;
	wire [4-1:0] node40875;
	wire [4-1:0] node40876;
	wire [4-1:0] node40877;
	wire [4-1:0] node40878;
	wire [4-1:0] node40879;
	wire [4-1:0] node40883;
	wire [4-1:0] node40884;
	wire [4-1:0] node40887;
	wire [4-1:0] node40890;
	wire [4-1:0] node40891;
	wire [4-1:0] node40894;
	wire [4-1:0] node40897;
	wire [4-1:0] node40898;
	wire [4-1:0] node40899;
	wire [4-1:0] node40900;
	wire [4-1:0] node40903;
	wire [4-1:0] node40906;
	wire [4-1:0] node40908;
	wire [4-1:0] node40909;
	wire [4-1:0] node40913;
	wire [4-1:0] node40914;
	wire [4-1:0] node40916;
	wire [4-1:0] node40917;
	wire [4-1:0] node40920;
	wire [4-1:0] node40923;
	wire [4-1:0] node40924;
	wire [4-1:0] node40925;
	wire [4-1:0] node40928;
	wire [4-1:0] node40932;
	wire [4-1:0] node40933;
	wire [4-1:0] node40934;
	wire [4-1:0] node40935;
	wire [4-1:0] node40936;
	wire [4-1:0] node40937;
	wire [4-1:0] node40940;
	wire [4-1:0] node40944;
	wire [4-1:0] node40945;
	wire [4-1:0] node40947;
	wire [4-1:0] node40950;
	wire [4-1:0] node40952;
	wire [4-1:0] node40955;
	wire [4-1:0] node40956;
	wire [4-1:0] node40957;
	wire [4-1:0] node40959;
	wire [4-1:0] node40962;
	wire [4-1:0] node40963;
	wire [4-1:0] node40966;
	wire [4-1:0] node40969;
	wire [4-1:0] node40970;
	wire [4-1:0] node40971;
	wire [4-1:0] node40974;
	wire [4-1:0] node40978;
	wire [4-1:0] node40979;
	wire [4-1:0] node40980;
	wire [4-1:0] node40981;
	wire [4-1:0] node40983;
	wire [4-1:0] node40986;
	wire [4-1:0] node40987;
	wire [4-1:0] node40991;
	wire [4-1:0] node40992;
	wire [4-1:0] node40994;
	wire [4-1:0] node40998;
	wire [4-1:0] node40999;
	wire [4-1:0] node41000;
	wire [4-1:0] node41003;
	wire [4-1:0] node41007;
	wire [4-1:0] node41008;
	wire [4-1:0] node41009;
	wire [4-1:0] node41010;
	wire [4-1:0] node41011;
	wire [4-1:0] node41012;
	wire [4-1:0] node41013;
	wire [4-1:0] node41017;
	wire [4-1:0] node41019;
	wire [4-1:0] node41022;
	wire [4-1:0] node41023;
	wire [4-1:0] node41026;
	wire [4-1:0] node41029;
	wire [4-1:0] node41030;
	wire [4-1:0] node41031;
	wire [4-1:0] node41032;
	wire [4-1:0] node41037;
	wire [4-1:0] node41038;
	wire [4-1:0] node41041;
	wire [4-1:0] node41044;
	wire [4-1:0] node41045;
	wire [4-1:0] node41046;
	wire [4-1:0] node41047;
	wire [4-1:0] node41048;
	wire [4-1:0] node41051;
	wire [4-1:0] node41054;
	wire [4-1:0] node41055;
	wire [4-1:0] node41059;
	wire [4-1:0] node41060;
	wire [4-1:0] node41063;
	wire [4-1:0] node41066;
	wire [4-1:0] node41067;
	wire [4-1:0] node41068;
	wire [4-1:0] node41069;
	wire [4-1:0] node41072;
	wire [4-1:0] node41075;
	wire [4-1:0] node41076;
	wire [4-1:0] node41079;
	wire [4-1:0] node41082;
	wire [4-1:0] node41083;
	wire [4-1:0] node41086;
	wire [4-1:0] node41089;
	wire [4-1:0] node41090;
	wire [4-1:0] node41091;
	wire [4-1:0] node41092;
	wire [4-1:0] node41094;
	wire [4-1:0] node41097;
	wire [4-1:0] node41098;
	wire [4-1:0] node41099;
	wire [4-1:0] node41102;
	wire [4-1:0] node41105;
	wire [4-1:0] node41107;
	wire [4-1:0] node41110;
	wire [4-1:0] node41111;
	wire [4-1:0] node41112;
	wire [4-1:0] node41114;
	wire [4-1:0] node41117;
	wire [4-1:0] node41119;
	wire [4-1:0] node41123;
	wire [4-1:0] node41124;
	wire [4-1:0] node41125;
	wire [4-1:0] node41126;
	wire [4-1:0] node41130;
	wire [4-1:0] node41131;
	wire [4-1:0] node41134;
	wire [4-1:0] node41137;
	wire [4-1:0] node41138;
	wire [4-1:0] node41141;
	wire [4-1:0] node41142;
	wire [4-1:0] node41145;
	wire [4-1:0] node41146;
	wire [4-1:0] node41150;
	wire [4-1:0] node41151;
	wire [4-1:0] node41152;
	wire [4-1:0] node41153;
	wire [4-1:0] node41154;
	wire [4-1:0] node41155;
	wire [4-1:0] node41156;
	wire [4-1:0] node41157;
	wire [4-1:0] node41159;
	wire [4-1:0] node41163;
	wire [4-1:0] node41164;
	wire [4-1:0] node41167;
	wire [4-1:0] node41169;
	wire [4-1:0] node41172;
	wire [4-1:0] node41173;
	wire [4-1:0] node41174;
	wire [4-1:0] node41177;
	wire [4-1:0] node41180;
	wire [4-1:0] node41181;
	wire [4-1:0] node41183;
	wire [4-1:0] node41187;
	wire [4-1:0] node41188;
	wire [4-1:0] node41190;
	wire [4-1:0] node41191;
	wire [4-1:0] node41194;
	wire [4-1:0] node41197;
	wire [4-1:0] node41198;
	wire [4-1:0] node41200;
	wire [4-1:0] node41203;
	wire [4-1:0] node41206;
	wire [4-1:0] node41207;
	wire [4-1:0] node41208;
	wire [4-1:0] node41211;
	wire [4-1:0] node41214;
	wire [4-1:0] node41215;
	wire [4-1:0] node41216;
	wire [4-1:0] node41219;
	wire [4-1:0] node41222;
	wire [4-1:0] node41223;
	wire [4-1:0] node41226;
	wire [4-1:0] node41229;
	wire [4-1:0] node41230;
	wire [4-1:0] node41231;
	wire [4-1:0] node41232;
	wire [4-1:0] node41233;
	wire [4-1:0] node41236;
	wire [4-1:0] node41238;
	wire [4-1:0] node41241;
	wire [4-1:0] node41242;
	wire [4-1:0] node41244;
	wire [4-1:0] node41247;
	wire [4-1:0] node41249;
	wire [4-1:0] node41252;
	wire [4-1:0] node41253;
	wire [4-1:0] node41254;
	wire [4-1:0] node41256;
	wire [4-1:0] node41258;
	wire [4-1:0] node41261;
	wire [4-1:0] node41262;
	wire [4-1:0] node41263;
	wire [4-1:0] node41268;
	wire [4-1:0] node41269;
	wire [4-1:0] node41270;
	wire [4-1:0] node41273;
	wire [4-1:0] node41276;
	wire [4-1:0] node41278;
	wire [4-1:0] node41281;
	wire [4-1:0] node41282;
	wire [4-1:0] node41283;
	wire [4-1:0] node41284;
	wire [4-1:0] node41285;
	wire [4-1:0] node41288;
	wire [4-1:0] node41291;
	wire [4-1:0] node41292;
	wire [4-1:0] node41293;
	wire [4-1:0] node41296;
	wire [4-1:0] node41299;
	wire [4-1:0] node41301;
	wire [4-1:0] node41304;
	wire [4-1:0] node41305;
	wire [4-1:0] node41306;
	wire [4-1:0] node41310;
	wire [4-1:0] node41312;
	wire [4-1:0] node41313;
	wire [4-1:0] node41316;
	wire [4-1:0] node41319;
	wire [4-1:0] node41320;
	wire [4-1:0] node41321;
	wire [4-1:0] node41322;
	wire [4-1:0] node41325;
	wire [4-1:0] node41328;
	wire [4-1:0] node41329;
	wire [4-1:0] node41332;
	wire [4-1:0] node41335;
	wire [4-1:0] node41336;
	wire [4-1:0] node41337;
	wire [4-1:0] node41340;
	wire [4-1:0] node41343;
	wire [4-1:0] node41344;
	wire [4-1:0] node41346;
	wire [4-1:0] node41349;
	wire [4-1:0] node41351;
	wire [4-1:0] node41354;
	wire [4-1:0] node41355;
	wire [4-1:0] node41356;
	wire [4-1:0] node41357;
	wire [4-1:0] node41358;
	wire [4-1:0] node41359;
	wire [4-1:0] node41361;
	wire [4-1:0] node41364;
	wire [4-1:0] node41366;
	wire [4-1:0] node41369;
	wire [4-1:0] node41370;
	wire [4-1:0] node41372;
	wire [4-1:0] node41375;
	wire [4-1:0] node41377;
	wire [4-1:0] node41380;
	wire [4-1:0] node41381;
	wire [4-1:0] node41382;
	wire [4-1:0] node41385;
	wire [4-1:0] node41386;
	wire [4-1:0] node41390;
	wire [4-1:0] node41391;
	wire [4-1:0] node41392;
	wire [4-1:0] node41397;
	wire [4-1:0] node41398;
	wire [4-1:0] node41399;
	wire [4-1:0] node41400;
	wire [4-1:0] node41401;
	wire [4-1:0] node41402;
	wire [4-1:0] node41405;
	wire [4-1:0] node41408;
	wire [4-1:0] node41409;
	wire [4-1:0] node41413;
	wire [4-1:0] node41415;
	wire [4-1:0] node41416;
	wire [4-1:0] node41419;
	wire [4-1:0] node41422;
	wire [4-1:0] node41423;
	wire [4-1:0] node41424;
	wire [4-1:0] node41425;
	wire [4-1:0] node41428;
	wire [4-1:0] node41432;
	wire [4-1:0] node41433;
	wire [4-1:0] node41434;
	wire [4-1:0] node41437;
	wire [4-1:0] node41441;
	wire [4-1:0] node41442;
	wire [4-1:0] node41443;
	wire [4-1:0] node41446;
	wire [4-1:0] node41449;
	wire [4-1:0] node41450;
	wire [4-1:0] node41453;
	wire [4-1:0] node41456;
	wire [4-1:0] node41457;
	wire [4-1:0] node41458;
	wire [4-1:0] node41459;
	wire [4-1:0] node41460;
	wire [4-1:0] node41461;
	wire [4-1:0] node41464;
	wire [4-1:0] node41468;
	wire [4-1:0] node41469;
	wire [4-1:0] node41470;
	wire [4-1:0] node41471;
	wire [4-1:0] node41474;
	wire [4-1:0] node41478;
	wire [4-1:0] node41479;
	wire [4-1:0] node41480;
	wire [4-1:0] node41483;
	wire [4-1:0] node41486;
	wire [4-1:0] node41487;
	wire [4-1:0] node41490;
	wire [4-1:0] node41493;
	wire [4-1:0] node41494;
	wire [4-1:0] node41495;
	wire [4-1:0] node41496;
	wire [4-1:0] node41500;
	wire [4-1:0] node41501;
	wire [4-1:0] node41505;
	wire [4-1:0] node41506;
	wire [4-1:0] node41507;
	wire [4-1:0] node41511;
	wire [4-1:0] node41512;
	wire [4-1:0] node41516;
	wire [4-1:0] node41517;
	wire [4-1:0] node41518;
	wire [4-1:0] node41519;
	wire [4-1:0] node41523;
	wire [4-1:0] node41524;
	wire [4-1:0] node41528;
	wire [4-1:0] node41529;
	wire [4-1:0] node41530;
	wire [4-1:0] node41534;
	wire [4-1:0] node41535;
	wire [4-1:0] node41539;
	wire [4-1:0] node41540;
	wire [4-1:0] node41541;
	wire [4-1:0] node41542;
	wire [4-1:0] node41543;
	wire [4-1:0] node41544;
	wire [4-1:0] node41545;
	wire [4-1:0] node41546;
	wire [4-1:0] node41547;
	wire [4-1:0] node41548;
	wire [4-1:0] node41549;
	wire [4-1:0] node41550;
	wire [4-1:0] node41553;
	wire [4-1:0] node41556;
	wire [4-1:0] node41558;
	wire [4-1:0] node41559;
	wire [4-1:0] node41562;
	wire [4-1:0] node41565;
	wire [4-1:0] node41566;
	wire [4-1:0] node41569;
	wire [4-1:0] node41570;
	wire [4-1:0] node41574;
	wire [4-1:0] node41575;
	wire [4-1:0] node41576;
	wire [4-1:0] node41579;
	wire [4-1:0] node41580;
	wire [4-1:0] node41583;
	wire [4-1:0] node41585;
	wire [4-1:0] node41588;
	wire [4-1:0] node41589;
	wire [4-1:0] node41590;
	wire [4-1:0] node41592;
	wire [4-1:0] node41596;
	wire [4-1:0] node41599;
	wire [4-1:0] node41600;
	wire [4-1:0] node41601;
	wire [4-1:0] node41602;
	wire [4-1:0] node41604;
	wire [4-1:0] node41607;
	wire [4-1:0] node41608;
	wire [4-1:0] node41610;
	wire [4-1:0] node41614;
	wire [4-1:0] node41615;
	wire [4-1:0] node41616;
	wire [4-1:0] node41618;
	wire [4-1:0] node41621;
	wire [4-1:0] node41624;
	wire [4-1:0] node41626;
	wire [4-1:0] node41628;
	wire [4-1:0] node41631;
	wire [4-1:0] node41632;
	wire [4-1:0] node41633;
	wire [4-1:0] node41634;
	wire [4-1:0] node41636;
	wire [4-1:0] node41639;
	wire [4-1:0] node41641;
	wire [4-1:0] node41644;
	wire [4-1:0] node41645;
	wire [4-1:0] node41649;
	wire [4-1:0] node41650;
	wire [4-1:0] node41651;
	wire [4-1:0] node41655;
	wire [4-1:0] node41657;
	wire [4-1:0] node41659;
	wire [4-1:0] node41662;
	wire [4-1:0] node41663;
	wire [4-1:0] node41664;
	wire [4-1:0] node41665;
	wire [4-1:0] node41666;
	wire [4-1:0] node41667;
	wire [4-1:0] node41668;
	wire [4-1:0] node41673;
	wire [4-1:0] node41674;
	wire [4-1:0] node41675;
	wire [4-1:0] node41679;
	wire [4-1:0] node41680;
	wire [4-1:0] node41683;
	wire [4-1:0] node41686;
	wire [4-1:0] node41687;
	wire [4-1:0] node41688;
	wire [4-1:0] node41691;
	wire [4-1:0] node41695;
	wire [4-1:0] node41696;
	wire [4-1:0] node41697;
	wire [4-1:0] node41698;
	wire [4-1:0] node41701;
	wire [4-1:0] node41704;
	wire [4-1:0] node41705;
	wire [4-1:0] node41706;
	wire [4-1:0] node41709;
	wire [4-1:0] node41712;
	wire [4-1:0] node41713;
	wire [4-1:0] node41716;
	wire [4-1:0] node41719;
	wire [4-1:0] node41720;
	wire [4-1:0] node41722;
	wire [4-1:0] node41725;
	wire [4-1:0] node41727;
	wire [4-1:0] node41730;
	wire [4-1:0] node41731;
	wire [4-1:0] node41732;
	wire [4-1:0] node41733;
	wire [4-1:0] node41734;
	wire [4-1:0] node41735;
	wire [4-1:0] node41739;
	wire [4-1:0] node41742;
	wire [4-1:0] node41743;
	wire [4-1:0] node41744;
	wire [4-1:0] node41747;
	wire [4-1:0] node41750;
	wire [4-1:0] node41751;
	wire [4-1:0] node41755;
	wire [4-1:0] node41756;
	wire [4-1:0] node41757;
	wire [4-1:0] node41758;
	wire [4-1:0] node41761;
	wire [4-1:0] node41765;
	wire [4-1:0] node41767;
	wire [4-1:0] node41768;
	wire [4-1:0] node41772;
	wire [4-1:0] node41773;
	wire [4-1:0] node41774;
	wire [4-1:0] node41775;
	wire [4-1:0] node41776;
	wire [4-1:0] node41779;
	wire [4-1:0] node41782;
	wire [4-1:0] node41784;
	wire [4-1:0] node41787;
	wire [4-1:0] node41789;
	wire [4-1:0] node41792;
	wire [4-1:0] node41793;
	wire [4-1:0] node41794;
	wire [4-1:0] node41797;
	wire [4-1:0] node41800;
	wire [4-1:0] node41802;
	wire [4-1:0] node41805;
	wire [4-1:0] node41806;
	wire [4-1:0] node41807;
	wire [4-1:0] node41808;
	wire [4-1:0] node41809;
	wire [4-1:0] node41810;
	wire [4-1:0] node41811;
	wire [4-1:0] node41814;
	wire [4-1:0] node41815;
	wire [4-1:0] node41818;
	wire [4-1:0] node41821;
	wire [4-1:0] node41822;
	wire [4-1:0] node41823;
	wire [4-1:0] node41827;
	wire [4-1:0] node41829;
	wire [4-1:0] node41832;
	wire [4-1:0] node41833;
	wire [4-1:0] node41834;
	wire [4-1:0] node41835;
	wire [4-1:0] node41838;
	wire [4-1:0] node41841;
	wire [4-1:0] node41842;
	wire [4-1:0] node41846;
	wire [4-1:0] node41847;
	wire [4-1:0] node41848;
	wire [4-1:0] node41852;
	wire [4-1:0] node41854;
	wire [4-1:0] node41857;
	wire [4-1:0] node41858;
	wire [4-1:0] node41859;
	wire [4-1:0] node41860;
	wire [4-1:0] node41861;
	wire [4-1:0] node41864;
	wire [4-1:0] node41867;
	wire [4-1:0] node41868;
	wire [4-1:0] node41872;
	wire [4-1:0] node41874;
	wire [4-1:0] node41875;
	wire [4-1:0] node41878;
	wire [4-1:0] node41881;
	wire [4-1:0] node41882;
	wire [4-1:0] node41883;
	wire [4-1:0] node41884;
	wire [4-1:0] node41887;
	wire [4-1:0] node41890;
	wire [4-1:0] node41893;
	wire [4-1:0] node41894;
	wire [4-1:0] node41895;
	wire [4-1:0] node41898;
	wire [4-1:0] node41901;
	wire [4-1:0] node41902;
	wire [4-1:0] node41905;
	wire [4-1:0] node41908;
	wire [4-1:0] node41909;
	wire [4-1:0] node41910;
	wire [4-1:0] node41911;
	wire [4-1:0] node41912;
	wire [4-1:0] node41913;
	wire [4-1:0] node41916;
	wire [4-1:0] node41920;
	wire [4-1:0] node41922;
	wire [4-1:0] node41923;
	wire [4-1:0] node41926;
	wire [4-1:0] node41929;
	wire [4-1:0] node41930;
	wire [4-1:0] node41931;
	wire [4-1:0] node41932;
	wire [4-1:0] node41935;
	wire [4-1:0] node41938;
	wire [4-1:0] node41941;
	wire [4-1:0] node41942;
	wire [4-1:0] node41943;
	wire [4-1:0] node41946;
	wire [4-1:0] node41949;
	wire [4-1:0] node41950;
	wire [4-1:0] node41953;
	wire [4-1:0] node41956;
	wire [4-1:0] node41957;
	wire [4-1:0] node41958;
	wire [4-1:0] node41959;
	wire [4-1:0] node41963;
	wire [4-1:0] node41965;
	wire [4-1:0] node41966;
	wire [4-1:0] node41969;
	wire [4-1:0] node41972;
	wire [4-1:0] node41973;
	wire [4-1:0] node41974;
	wire [4-1:0] node41975;
	wire [4-1:0] node41978;
	wire [4-1:0] node41981;
	wire [4-1:0] node41982;
	wire [4-1:0] node41985;
	wire [4-1:0] node41988;
	wire [4-1:0] node41989;
	wire [4-1:0] node41992;
	wire [4-1:0] node41995;
	wire [4-1:0] node41996;
	wire [4-1:0] node41997;
	wire [4-1:0] node41998;
	wire [4-1:0] node41999;
	wire [4-1:0] node42001;
	wire [4-1:0] node42004;
	wire [4-1:0] node42005;
	wire [4-1:0] node42008;
	wire [4-1:0] node42011;
	wire [4-1:0] node42012;
	wire [4-1:0] node42013;
	wire [4-1:0] node42016;
	wire [4-1:0] node42019;
	wire [4-1:0] node42022;
	wire [4-1:0] node42023;
	wire [4-1:0] node42024;
	wire [4-1:0] node42025;
	wire [4-1:0] node42029;
	wire [4-1:0] node42031;
	wire [4-1:0] node42034;
	wire [4-1:0] node42035;
	wire [4-1:0] node42036;
	wire [4-1:0] node42040;
	wire [4-1:0] node42042;
	wire [4-1:0] node42043;
	wire [4-1:0] node42046;
	wire [4-1:0] node42049;
	wire [4-1:0] node42050;
	wire [4-1:0] node42051;
	wire [4-1:0] node42052;
	wire [4-1:0] node42053;
	wire [4-1:0] node42054;
	wire [4-1:0] node42057;
	wire [4-1:0] node42060;
	wire [4-1:0] node42061;
	wire [4-1:0] node42064;
	wire [4-1:0] node42067;
	wire [4-1:0] node42068;
	wire [4-1:0] node42070;
	wire [4-1:0] node42073;
	wire [4-1:0] node42074;
	wire [4-1:0] node42078;
	wire [4-1:0] node42079;
	wire [4-1:0] node42080;
	wire [4-1:0] node42081;
	wire [4-1:0] node42085;
	wire [4-1:0] node42086;
	wire [4-1:0] node42089;
	wire [4-1:0] node42092;
	wire [4-1:0] node42093;
	wire [4-1:0] node42094;
	wire [4-1:0] node42097;
	wire [4-1:0] node42100;
	wire [4-1:0] node42101;
	wire [4-1:0] node42104;
	wire [4-1:0] node42107;
	wire [4-1:0] node42108;
	wire [4-1:0] node42109;
	wire [4-1:0] node42110;
	wire [4-1:0] node42112;
	wire [4-1:0] node42115;
	wire [4-1:0] node42116;
	wire [4-1:0] node42119;
	wire [4-1:0] node42122;
	wire [4-1:0] node42123;
	wire [4-1:0] node42124;
	wire [4-1:0] node42127;
	wire [4-1:0] node42130;
	wire [4-1:0] node42131;
	wire [4-1:0] node42135;
	wire [4-1:0] node42136;
	wire [4-1:0] node42138;
	wire [4-1:0] node42139;
	wire [4-1:0] node42143;
	wire [4-1:0] node42144;
	wire [4-1:0] node42145;
	wire [4-1:0] node42149;
	wire [4-1:0] node42150;
	wire [4-1:0] node42153;
	wire [4-1:0] node42156;
	wire [4-1:0] node42157;
	wire [4-1:0] node42158;
	wire [4-1:0] node42159;
	wire [4-1:0] node42160;
	wire [4-1:0] node42161;
	wire [4-1:0] node42163;
	wire [4-1:0] node42166;
	wire [4-1:0] node42168;
	wire [4-1:0] node42171;
	wire [4-1:0] node42172;
	wire [4-1:0] node42174;
	wire [4-1:0] node42177;
	wire [4-1:0] node42179;
	wire [4-1:0] node42182;
	wire [4-1:0] node42183;
	wire [4-1:0] node42184;
	wire [4-1:0] node42185;
	wire [4-1:0] node42187;
	wire [4-1:0] node42190;
	wire [4-1:0] node42192;
	wire [4-1:0] node42195;
	wire [4-1:0] node42196;
	wire [4-1:0] node42198;
	wire [4-1:0] node42201;
	wire [4-1:0] node42203;
	wire [4-1:0] node42206;
	wire [4-1:0] node42207;
	wire [4-1:0] node42208;
	wire [4-1:0] node42209;
	wire [4-1:0] node42212;
	wire [4-1:0] node42215;
	wire [4-1:0] node42217;
	wire [4-1:0] node42220;
	wire [4-1:0] node42221;
	wire [4-1:0] node42222;
	wire [4-1:0] node42223;
	wire [4-1:0] node42226;
	wire [4-1:0] node42229;
	wire [4-1:0] node42230;
	wire [4-1:0] node42233;
	wire [4-1:0] node42236;
	wire [4-1:0] node42237;
	wire [4-1:0] node42238;
	wire [4-1:0] node42241;
	wire [4-1:0] node42244;
	wire [4-1:0] node42245;
	wire [4-1:0] node42249;
	wire [4-1:0] node42250;
	wire [4-1:0] node42251;
	wire [4-1:0] node42252;
	wire [4-1:0] node42253;
	wire [4-1:0] node42255;
	wire [4-1:0] node42258;
	wire [4-1:0] node42260;
	wire [4-1:0] node42263;
	wire [4-1:0] node42266;
	wire [4-1:0] node42267;
	wire [4-1:0] node42268;
	wire [4-1:0] node42269;
	wire [4-1:0] node42272;
	wire [4-1:0] node42275;
	wire [4-1:0] node42276;
	wire [4-1:0] node42277;
	wire [4-1:0] node42280;
	wire [4-1:0] node42283;
	wire [4-1:0] node42284;
	wire [4-1:0] node42287;
	wire [4-1:0] node42290;
	wire [4-1:0] node42291;
	wire [4-1:0] node42292;
	wire [4-1:0] node42295;
	wire [4-1:0] node42298;
	wire [4-1:0] node42299;
	wire [4-1:0] node42302;
	wire [4-1:0] node42305;
	wire [4-1:0] node42306;
	wire [4-1:0] node42307;
	wire [4-1:0] node42308;
	wire [4-1:0] node42310;
	wire [4-1:0] node42313;
	wire [4-1:0] node42315;
	wire [4-1:0] node42318;
	wire [4-1:0] node42319;
	wire [4-1:0] node42321;
	wire [4-1:0] node42324;
	wire [4-1:0] node42327;
	wire [4-1:0] node42328;
	wire [4-1:0] node42329;
	wire [4-1:0] node42330;
	wire [4-1:0] node42334;
	wire [4-1:0] node42335;
	wire [4-1:0] node42339;
	wire [4-1:0] node42340;
	wire [4-1:0] node42341;
	wire [4-1:0] node42342;
	wire [4-1:0] node42345;
	wire [4-1:0] node42348;
	wire [4-1:0] node42349;
	wire [4-1:0] node42353;
	wire [4-1:0] node42356;
	wire [4-1:0] node42357;
	wire [4-1:0] node42358;
	wire [4-1:0] node42359;
	wire [4-1:0] node42360;
	wire [4-1:0] node42363;
	wire [4-1:0] node42366;
	wire [4-1:0] node42367;
	wire [4-1:0] node42368;
	wire [4-1:0] node42369;
	wire [4-1:0] node42373;
	wire [4-1:0] node42374;
	wire [4-1:0] node42377;
	wire [4-1:0] node42380;
	wire [4-1:0] node42381;
	wire [4-1:0] node42384;
	wire [4-1:0] node42387;
	wire [4-1:0] node42388;
	wire [4-1:0] node42389;
	wire [4-1:0] node42390;
	wire [4-1:0] node42391;
	wire [4-1:0] node42394;
	wire [4-1:0] node42397;
	wire [4-1:0] node42399;
	wire [4-1:0] node42400;
	wire [4-1:0] node42403;
	wire [4-1:0] node42406;
	wire [4-1:0] node42407;
	wire [4-1:0] node42408;
	wire [4-1:0] node42411;
	wire [4-1:0] node42414;
	wire [4-1:0] node42415;
	wire [4-1:0] node42416;
	wire [4-1:0] node42419;
	wire [4-1:0] node42422;
	wire [4-1:0] node42423;
	wire [4-1:0] node42426;
	wire [4-1:0] node42429;
	wire [4-1:0] node42430;
	wire [4-1:0] node42431;
	wire [4-1:0] node42433;
	wire [4-1:0] node42434;
	wire [4-1:0] node42437;
	wire [4-1:0] node42440;
	wire [4-1:0] node42441;
	wire [4-1:0] node42444;
	wire [4-1:0] node42447;
	wire [4-1:0] node42448;
	wire [4-1:0] node42451;
	wire [4-1:0] node42454;
	wire [4-1:0] node42455;
	wire [4-1:0] node42456;
	wire [4-1:0] node42457;
	wire [4-1:0] node42458;
	wire [4-1:0] node42459;
	wire [4-1:0] node42460;
	wire [4-1:0] node42463;
	wire [4-1:0] node42467;
	wire [4-1:0] node42468;
	wire [4-1:0] node42471;
	wire [4-1:0] node42474;
	wire [4-1:0] node42476;
	wire [4-1:0] node42477;
	wire [4-1:0] node42479;
	wire [4-1:0] node42482;
	wire [4-1:0] node42483;
	wire [4-1:0] node42487;
	wire [4-1:0] node42488;
	wire [4-1:0] node42489;
	wire [4-1:0] node42490;
	wire [4-1:0] node42494;
	wire [4-1:0] node42495;
	wire [4-1:0] node42499;
	wire [4-1:0] node42500;
	wire [4-1:0] node42501;
	wire [4-1:0] node42505;
	wire [4-1:0] node42506;
	wire [4-1:0] node42510;
	wire [4-1:0] node42511;
	wire [4-1:0] node42512;
	wire [4-1:0] node42513;
	wire [4-1:0] node42514;
	wire [4-1:0] node42518;
	wire [4-1:0] node42520;
	wire [4-1:0] node42523;
	wire [4-1:0] node42524;
	wire [4-1:0] node42525;
	wire [4-1:0] node42529;
	wire [4-1:0] node42530;
	wire [4-1:0] node42534;
	wire [4-1:0] node42535;
	wire [4-1:0] node42536;
	wire [4-1:0] node42537;
	wire [4-1:0] node42541;
	wire [4-1:0] node42542;
	wire [4-1:0] node42546;
	wire [4-1:0] node42547;
	wire [4-1:0] node42550;
	wire [4-1:0] node42551;
	wire [4-1:0] node42555;
	wire [4-1:0] node42556;
	wire [4-1:0] node42557;
	wire [4-1:0] node42558;
	wire [4-1:0] node42559;
	wire [4-1:0] node42560;
	wire [4-1:0] node42561;
	wire [4-1:0] node42563;
	wire [4-1:0] node42564;
	wire [4-1:0] node42567;
	wire [4-1:0] node42570;
	wire [4-1:0] node42571;
	wire [4-1:0] node42572;
	wire [4-1:0] node42575;
	wire [4-1:0] node42578;
	wire [4-1:0] node42579;
	wire [4-1:0] node42580;
	wire [4-1:0] node42584;
	wire [4-1:0] node42587;
	wire [4-1:0] node42588;
	wire [4-1:0] node42589;
	wire [4-1:0] node42591;
	wire [4-1:0] node42594;
	wire [4-1:0] node42595;
	wire [4-1:0] node42597;
	wire [4-1:0] node42601;
	wire [4-1:0] node42602;
	wire [4-1:0] node42603;
	wire [4-1:0] node42606;
	wire [4-1:0] node42609;
	wire [4-1:0] node42610;
	wire [4-1:0] node42611;
	wire [4-1:0] node42614;
	wire [4-1:0] node42617;
	wire [4-1:0] node42618;
	wire [4-1:0] node42621;
	wire [4-1:0] node42624;
	wire [4-1:0] node42625;
	wire [4-1:0] node42626;
	wire [4-1:0] node42627;
	wire [4-1:0] node42629;
	wire [4-1:0] node42632;
	wire [4-1:0] node42634;
	wire [4-1:0] node42637;
	wire [4-1:0] node42638;
	wire [4-1:0] node42640;
	wire [4-1:0] node42643;
	wire [4-1:0] node42645;
	wire [4-1:0] node42648;
	wire [4-1:0] node42649;
	wire [4-1:0] node42650;
	wire [4-1:0] node42651;
	wire [4-1:0] node42652;
	wire [4-1:0] node42655;
	wire [4-1:0] node42658;
	wire [4-1:0] node42659;
	wire [4-1:0] node42662;
	wire [4-1:0] node42665;
	wire [4-1:0] node42666;
	wire [4-1:0] node42669;
	wire [4-1:0] node42672;
	wire [4-1:0] node42673;
	wire [4-1:0] node42674;
	wire [4-1:0] node42677;
	wire [4-1:0] node42680;
	wire [4-1:0] node42681;
	wire [4-1:0] node42684;
	wire [4-1:0] node42687;
	wire [4-1:0] node42688;
	wire [4-1:0] node42689;
	wire [4-1:0] node42690;
	wire [4-1:0] node42691;
	wire [4-1:0] node42692;
	wire [4-1:0] node42693;
	wire [4-1:0] node42696;
	wire [4-1:0] node42699;
	wire [4-1:0] node42700;
	wire [4-1:0] node42704;
	wire [4-1:0] node42705;
	wire [4-1:0] node42706;
	wire [4-1:0] node42709;
	wire [4-1:0] node42712;
	wire [4-1:0] node42713;
	wire [4-1:0] node42717;
	wire [4-1:0] node42718;
	wire [4-1:0] node42719;
	wire [4-1:0] node42720;
	wire [4-1:0] node42723;
	wire [4-1:0] node42726;
	wire [4-1:0] node42727;
	wire [4-1:0] node42730;
	wire [4-1:0] node42733;
	wire [4-1:0] node42735;
	wire [4-1:0] node42737;
	wire [4-1:0] node42740;
	wire [4-1:0] node42741;
	wire [4-1:0] node42742;
	wire [4-1:0] node42743;
	wire [4-1:0] node42745;
	wire [4-1:0] node42748;
	wire [4-1:0] node42749;
	wire [4-1:0] node42752;
	wire [4-1:0] node42755;
	wire [4-1:0] node42756;
	wire [4-1:0] node42758;
	wire [4-1:0] node42761;
	wire [4-1:0] node42762;
	wire [4-1:0] node42766;
	wire [4-1:0] node42767;
	wire [4-1:0] node42768;
	wire [4-1:0] node42769;
	wire [4-1:0] node42772;
	wire [4-1:0] node42775;
	wire [4-1:0] node42776;
	wire [4-1:0] node42779;
	wire [4-1:0] node42782;
	wire [4-1:0] node42784;
	wire [4-1:0] node42786;
	wire [4-1:0] node42789;
	wire [4-1:0] node42790;
	wire [4-1:0] node42791;
	wire [4-1:0] node42792;
	wire [4-1:0] node42793;
	wire [4-1:0] node42794;
	wire [4-1:0] node42797;
	wire [4-1:0] node42800;
	wire [4-1:0] node42801;
	wire [4-1:0] node42804;
	wire [4-1:0] node42807;
	wire [4-1:0] node42808;
	wire [4-1:0] node42809;
	wire [4-1:0] node42813;
	wire [4-1:0] node42816;
	wire [4-1:0] node42817;
	wire [4-1:0] node42818;
	wire [4-1:0] node42819;
	wire [4-1:0] node42823;
	wire [4-1:0] node42824;
	wire [4-1:0] node42828;
	wire [4-1:0] node42829;
	wire [4-1:0] node42831;
	wire [4-1:0] node42834;
	wire [4-1:0] node42835;
	wire [4-1:0] node42839;
	wire [4-1:0] node42840;
	wire [4-1:0] node42841;
	wire [4-1:0] node42842;
	wire [4-1:0] node42843;
	wire [4-1:0] node42846;
	wire [4-1:0] node42849;
	wire [4-1:0] node42850;
	wire [4-1:0] node42853;
	wire [4-1:0] node42856;
	wire [4-1:0] node42857;
	wire [4-1:0] node42858;
	wire [4-1:0] node42861;
	wire [4-1:0] node42864;
	wire [4-1:0] node42866;
	wire [4-1:0] node42869;
	wire [4-1:0] node42870;
	wire [4-1:0] node42872;
	wire [4-1:0] node42873;
	wire [4-1:0] node42876;
	wire [4-1:0] node42879;
	wire [4-1:0] node42880;
	wire [4-1:0] node42881;
	wire [4-1:0] node42885;
	wire [4-1:0] node42886;
	wire [4-1:0] node42889;
	wire [4-1:0] node42892;
	wire [4-1:0] node42893;
	wire [4-1:0] node42894;
	wire [4-1:0] node42895;
	wire [4-1:0] node42896;
	wire [4-1:0] node42897;
	wire [4-1:0] node42898;
	wire [4-1:0] node42900;
	wire [4-1:0] node42903;
	wire [4-1:0] node42905;
	wire [4-1:0] node42909;
	wire [4-1:0] node42910;
	wire [4-1:0] node42911;
	wire [4-1:0] node42913;
	wire [4-1:0] node42917;
	wire [4-1:0] node42918;
	wire [4-1:0] node42919;
	wire [4-1:0] node42924;
	wire [4-1:0] node42925;
	wire [4-1:0] node42926;
	wire [4-1:0] node42927;
	wire [4-1:0] node42930;
	wire [4-1:0] node42932;
	wire [4-1:0] node42935;
	wire [4-1:0] node42937;
	wire [4-1:0] node42940;
	wire [4-1:0] node42941;
	wire [4-1:0] node42942;
	wire [4-1:0] node42945;
	wire [4-1:0] node42948;
	wire [4-1:0] node42949;
	wire [4-1:0] node42950;
	wire [4-1:0] node42953;
	wire [4-1:0] node42957;
	wire [4-1:0] node42958;
	wire [4-1:0] node42959;
	wire [4-1:0] node42960;
	wire [4-1:0] node42961;
	wire [4-1:0] node42965;
	wire [4-1:0] node42966;
	wire [4-1:0] node42968;
	wire [4-1:0] node42971;
	wire [4-1:0] node42974;
	wire [4-1:0] node42975;
	wire [4-1:0] node42978;
	wire [4-1:0] node42979;
	wire [4-1:0] node42980;
	wire [4-1:0] node42984;
	wire [4-1:0] node42987;
	wire [4-1:0] node42988;
	wire [4-1:0] node42989;
	wire [4-1:0] node42990;
	wire [4-1:0] node42991;
	wire [4-1:0] node42994;
	wire [4-1:0] node42998;
	wire [4-1:0] node42999;
	wire [4-1:0] node43000;
	wire [4-1:0] node43004;
	wire [4-1:0] node43005;
	wire [4-1:0] node43009;
	wire [4-1:0] node43010;
	wire [4-1:0] node43011;
	wire [4-1:0] node43012;
	wire [4-1:0] node43015;
	wire [4-1:0] node43018;
	wire [4-1:0] node43019;
	wire [4-1:0] node43023;
	wire [4-1:0] node43025;
	wire [4-1:0] node43027;
	wire [4-1:0] node43030;
	wire [4-1:0] node43031;
	wire [4-1:0] node43032;
	wire [4-1:0] node43033;
	wire [4-1:0] node43034;
	wire [4-1:0] node43035;
	wire [4-1:0] node43038;
	wire [4-1:0] node43041;
	wire [4-1:0] node43044;
	wire [4-1:0] node43045;
	wire [4-1:0] node43046;
	wire [4-1:0] node43047;
	wire [4-1:0] node43051;
	wire [4-1:0] node43054;
	wire [4-1:0] node43055;
	wire [4-1:0] node43056;
	wire [4-1:0] node43060;
	wire [4-1:0] node43061;
	wire [4-1:0] node43065;
	wire [4-1:0] node43066;
	wire [4-1:0] node43067;
	wire [4-1:0] node43068;
	wire [4-1:0] node43071;
	wire [4-1:0] node43074;
	wire [4-1:0] node43075;
	wire [4-1:0] node43078;
	wire [4-1:0] node43081;
	wire [4-1:0] node43082;
	wire [4-1:0] node43083;
	wire [4-1:0] node43086;
	wire [4-1:0] node43089;
	wire [4-1:0] node43090;
	wire [4-1:0] node43093;
	wire [4-1:0] node43096;
	wire [4-1:0] node43097;
	wire [4-1:0] node43098;
	wire [4-1:0] node43099;
	wire [4-1:0] node43101;
	wire [4-1:0] node43104;
	wire [4-1:0] node43105;
	wire [4-1:0] node43108;
	wire [4-1:0] node43111;
	wire [4-1:0] node43112;
	wire [4-1:0] node43113;
	wire [4-1:0] node43116;
	wire [4-1:0] node43119;
	wire [4-1:0] node43120;
	wire [4-1:0] node43123;
	wire [4-1:0] node43126;
	wire [4-1:0] node43127;
	wire [4-1:0] node43128;
	wire [4-1:0] node43129;
	wire [4-1:0] node43133;
	wire [4-1:0] node43136;
	wire [4-1:0] node43137;
	wire [4-1:0] node43138;
	wire [4-1:0] node43142;
	wire [4-1:0] node43145;
	wire [4-1:0] node43146;
	wire [4-1:0] node43147;
	wire [4-1:0] node43148;
	wire [4-1:0] node43149;
	wire [4-1:0] node43150;
	wire [4-1:0] node43151;
	wire [4-1:0] node43153;
	wire [4-1:0] node43156;
	wire [4-1:0] node43158;
	wire [4-1:0] node43161;
	wire [4-1:0] node43162;
	wire [4-1:0] node43164;
	wire [4-1:0] node43167;
	wire [4-1:0] node43169;
	wire [4-1:0] node43172;
	wire [4-1:0] node43173;
	wire [4-1:0] node43174;
	wire [4-1:0] node43175;
	wire [4-1:0] node43178;
	wire [4-1:0] node43181;
	wire [4-1:0] node43183;
	wire [4-1:0] node43186;
	wire [4-1:0] node43188;
	wire [4-1:0] node43190;
	wire [4-1:0] node43191;
	wire [4-1:0] node43194;
	wire [4-1:0] node43197;
	wire [4-1:0] node43198;
	wire [4-1:0] node43199;
	wire [4-1:0] node43200;
	wire [4-1:0] node43203;
	wire [4-1:0] node43206;
	wire [4-1:0] node43207;
	wire [4-1:0] node43209;
	wire [4-1:0] node43212;
	wire [4-1:0] node43213;
	wire [4-1:0] node43214;
	wire [4-1:0] node43217;
	wire [4-1:0] node43220;
	wire [4-1:0] node43222;
	wire [4-1:0] node43225;
	wire [4-1:0] node43226;
	wire [4-1:0] node43227;
	wire [4-1:0] node43228;
	wire [4-1:0] node43232;
	wire [4-1:0] node43233;
	wire [4-1:0] node43234;
	wire [4-1:0] node43237;
	wire [4-1:0] node43241;
	wire [4-1:0] node43242;
	wire [4-1:0] node43243;
	wire [4-1:0] node43244;
	wire [4-1:0] node43247;
	wire [4-1:0] node43252;
	wire [4-1:0] node43253;
	wire [4-1:0] node43254;
	wire [4-1:0] node43255;
	wire [4-1:0] node43256;
	wire [4-1:0] node43258;
	wire [4-1:0] node43262;
	wire [4-1:0] node43263;
	wire [4-1:0] node43265;
	wire [4-1:0] node43268;
	wire [4-1:0] node43270;
	wire [4-1:0] node43273;
	wire [4-1:0] node43274;
	wire [4-1:0] node43275;
	wire [4-1:0] node43276;
	wire [4-1:0] node43280;
	wire [4-1:0] node43281;
	wire [4-1:0] node43285;
	wire [4-1:0] node43286;
	wire [4-1:0] node43287;
	wire [4-1:0] node43291;
	wire [4-1:0] node43292;
	wire [4-1:0] node43296;
	wire [4-1:0] node43297;
	wire [4-1:0] node43298;
	wire [4-1:0] node43299;
	wire [4-1:0] node43300;
	wire [4-1:0] node43301;
	wire [4-1:0] node43305;
	wire [4-1:0] node43306;
	wire [4-1:0] node43310;
	wire [4-1:0] node43311;
	wire [4-1:0] node43312;
	wire [4-1:0] node43316;
	wire [4-1:0] node43317;
	wire [4-1:0] node43321;
	wire [4-1:0] node43322;
	wire [4-1:0] node43324;
	wire [4-1:0] node43325;
	wire [4-1:0] node43329;
	wire [4-1:0] node43330;
	wire [4-1:0] node43331;
	wire [4-1:0] node43336;
	wire [4-1:0] node43337;
	wire [4-1:0] node43338;
	wire [4-1:0] node43339;
	wire [4-1:0] node43340;
	wire [4-1:0] node43344;
	wire [4-1:0] node43345;
	wire [4-1:0] node43348;
	wire [4-1:0] node43351;
	wire [4-1:0] node43352;
	wire [4-1:0] node43355;
	wire [4-1:0] node43358;
	wire [4-1:0] node43359;
	wire [4-1:0] node43362;
	wire [4-1:0] node43365;
	wire [4-1:0] node43366;
	wire [4-1:0] node43367;
	wire [4-1:0] node43368;
	wire [4-1:0] node43369;
	wire [4-1:0] node43370;
	wire [4-1:0] node43371;
	wire [4-1:0] node43373;
	wire [4-1:0] node43376;
	wire [4-1:0] node43378;
	wire [4-1:0] node43381;
	wire [4-1:0] node43382;
	wire [4-1:0] node43384;
	wire [4-1:0] node43387;
	wire [4-1:0] node43389;
	wire [4-1:0] node43392;
	wire [4-1:0] node43393;
	wire [4-1:0] node43394;
	wire [4-1:0] node43398;
	wire [4-1:0] node43399;
	wire [4-1:0] node43400;
	wire [4-1:0] node43404;
	wire [4-1:0] node43405;
	wire [4-1:0] node43409;
	wire [4-1:0] node43410;
	wire [4-1:0] node43411;
	wire [4-1:0] node43412;
	wire [4-1:0] node43414;
	wire [4-1:0] node43417;
	wire [4-1:0] node43419;
	wire [4-1:0] node43422;
	wire [4-1:0] node43423;
	wire [4-1:0] node43425;
	wire [4-1:0] node43429;
	wire [4-1:0] node43430;
	wire [4-1:0] node43433;
	wire [4-1:0] node43436;
	wire [4-1:0] node43437;
	wire [4-1:0] node43438;
	wire [4-1:0] node43439;
	wire [4-1:0] node43440;
	wire [4-1:0] node43443;
	wire [4-1:0] node43446;
	wire [4-1:0] node43448;
	wire [4-1:0] node43449;
	wire [4-1:0] node43453;
	wire [4-1:0] node43454;
	wire [4-1:0] node43455;
	wire [4-1:0] node43458;
	wire [4-1:0] node43461;
	wire [4-1:0] node43462;
	wire [4-1:0] node43463;
	wire [4-1:0] node43466;
	wire [4-1:0] node43469;
	wire [4-1:0] node43470;
	wire [4-1:0] node43473;
	wire [4-1:0] node43476;
	wire [4-1:0] node43477;
	wire [4-1:0] node43478;
	wire [4-1:0] node43481;
	wire [4-1:0] node43484;
	wire [4-1:0] node43485;
	wire [4-1:0] node43488;
	wire [4-1:0] node43491;
	wire [4-1:0] node43492;
	wire [4-1:0] node43493;
	wire [4-1:0] node43494;
	wire [4-1:0] node43495;
	wire [4-1:0] node43496;
	wire [4-1:0] node43500;
	wire [4-1:0] node43503;
	wire [4-1:0] node43504;
	wire [4-1:0] node43505;
	wire [4-1:0] node43509;
	wire [4-1:0] node43510;
	wire [4-1:0] node43514;
	wire [4-1:0] node43515;
	wire [4-1:0] node43516;
	wire [4-1:0] node43517;
	wire [4-1:0] node43518;
	wire [4-1:0] node43521;
	wire [4-1:0] node43524;
	wire [4-1:0] node43525;
	wire [4-1:0] node43528;
	wire [4-1:0] node43531;
	wire [4-1:0] node43532;
	wire [4-1:0] node43535;
	wire [4-1:0] node43538;
	wire [4-1:0] node43539;
	wire [4-1:0] node43541;
	wire [4-1:0] node43542;
	wire [4-1:0] node43546;
	wire [4-1:0] node43547;
	wire [4-1:0] node43550;
	wire [4-1:0] node43553;
	wire [4-1:0] node43554;
	wire [4-1:0] node43555;
	wire [4-1:0] node43556;
	wire [4-1:0] node43557;
	wire [4-1:0] node43558;
	wire [4-1:0] node43561;
	wire [4-1:0] node43565;
	wire [4-1:0] node43566;
	wire [4-1:0] node43567;
	wire [4-1:0] node43570;
	wire [4-1:0] node43574;
	wire [4-1:0] node43575;
	wire [4-1:0] node43576;
	wire [4-1:0] node43578;
	wire [4-1:0] node43581;
	wire [4-1:0] node43583;
	wire [4-1:0] node43586;
	wire [4-1:0] node43588;
	wire [4-1:0] node43589;
	wire [4-1:0] node43592;
	wire [4-1:0] node43595;
	wire [4-1:0] node43596;
	wire [4-1:0] node43599;
	wire [4-1:0] node43602;
	wire [4-1:0] node43603;
	wire [4-1:0] node43604;
	wire [4-1:0] node43605;
	wire [4-1:0] node43606;
	wire [4-1:0] node43607;
	wire [4-1:0] node43608;
	wire [4-1:0] node43609;
	wire [4-1:0] node43610;
	wire [4-1:0] node43611;
	wire [4-1:0] node43612;
	wire [4-1:0] node43615;
	wire [4-1:0] node43618;
	wire [4-1:0] node43619;
	wire [4-1:0] node43623;
	wire [4-1:0] node43624;
	wire [4-1:0] node43625;
	wire [4-1:0] node43628;
	wire [4-1:0] node43631;
	wire [4-1:0] node43633;
	wire [4-1:0] node43636;
	wire [4-1:0] node43637;
	wire [4-1:0] node43639;
	wire [4-1:0] node43640;
	wire [4-1:0] node43643;
	wire [4-1:0] node43646;
	wire [4-1:0] node43647;
	wire [4-1:0] node43649;
	wire [4-1:0] node43652;
	wire [4-1:0] node43653;
	wire [4-1:0] node43656;
	wire [4-1:0] node43659;
	wire [4-1:0] node43660;
	wire [4-1:0] node43661;
	wire [4-1:0] node43663;
	wire [4-1:0] node43665;
	wire [4-1:0] node43668;
	wire [4-1:0] node43670;
	wire [4-1:0] node43672;
	wire [4-1:0] node43675;
	wire [4-1:0] node43676;
	wire [4-1:0] node43677;
	wire [4-1:0] node43681;
	wire [4-1:0] node43684;
	wire [4-1:0] node43685;
	wire [4-1:0] node43686;
	wire [4-1:0] node43687;
	wire [4-1:0] node43688;
	wire [4-1:0] node43689;
	wire [4-1:0] node43692;
	wire [4-1:0] node43695;
	wire [4-1:0] node43696;
	wire [4-1:0] node43699;
	wire [4-1:0] node43702;
	wire [4-1:0] node43703;
	wire [4-1:0] node43704;
	wire [4-1:0] node43708;
	wire [4-1:0] node43710;
	wire [4-1:0] node43713;
	wire [4-1:0] node43714;
	wire [4-1:0] node43715;
	wire [4-1:0] node43716;
	wire [4-1:0] node43720;
	wire [4-1:0] node43721;
	wire [4-1:0] node43725;
	wire [4-1:0] node43726;
	wire [4-1:0] node43727;
	wire [4-1:0] node43730;
	wire [4-1:0] node43733;
	wire [4-1:0] node43735;
	wire [4-1:0] node43738;
	wire [4-1:0] node43739;
	wire [4-1:0] node43740;
	wire [4-1:0] node43741;
	wire [4-1:0] node43742;
	wire [4-1:0] node43746;
	wire [4-1:0] node43748;
	wire [4-1:0] node43752;
	wire [4-1:0] node43753;
	wire [4-1:0] node43754;
	wire [4-1:0] node43757;
	wire [4-1:0] node43759;
	wire [4-1:0] node43762;
	wire [4-1:0] node43763;
	wire [4-1:0] node43764;
	wire [4-1:0] node43767;
	wire [4-1:0] node43770;
	wire [4-1:0] node43771;
	wire [4-1:0] node43774;
	wire [4-1:0] node43777;
	wire [4-1:0] node43778;
	wire [4-1:0] node43779;
	wire [4-1:0] node43780;
	wire [4-1:0] node43781;
	wire [4-1:0] node43782;
	wire [4-1:0] node43784;
	wire [4-1:0] node43787;
	wire [4-1:0] node43789;
	wire [4-1:0] node43792;
	wire [4-1:0] node43793;
	wire [4-1:0] node43795;
	wire [4-1:0] node43799;
	wire [4-1:0] node43800;
	wire [4-1:0] node43801;
	wire [4-1:0] node43803;
	wire [4-1:0] node43806;
	wire [4-1:0] node43808;
	wire [4-1:0] node43811;
	wire [4-1:0] node43812;
	wire [4-1:0] node43816;
	wire [4-1:0] node43817;
	wire [4-1:0] node43818;
	wire [4-1:0] node43819;
	wire [4-1:0] node43821;
	wire [4-1:0] node43825;
	wire [4-1:0] node43826;
	wire [4-1:0] node43829;
	wire [4-1:0] node43831;
	wire [4-1:0] node43834;
	wire [4-1:0] node43835;
	wire [4-1:0] node43837;
	wire [4-1:0] node43840;
	wire [4-1:0] node43841;
	wire [4-1:0] node43845;
	wire [4-1:0] node43846;
	wire [4-1:0] node43847;
	wire [4-1:0] node43848;
	wire [4-1:0] node43849;
	wire [4-1:0] node43852;
	wire [4-1:0] node43855;
	wire [4-1:0] node43857;
	wire [4-1:0] node43858;
	wire [4-1:0] node43862;
	wire [4-1:0] node43863;
	wire [4-1:0] node43866;
	wire [4-1:0] node43867;
	wire [4-1:0] node43870;
	wire [4-1:0] node43873;
	wire [4-1:0] node43874;
	wire [4-1:0] node43875;
	wire [4-1:0] node43877;
	wire [4-1:0] node43878;
	wire [4-1:0] node43882;
	wire [4-1:0] node43883;
	wire [4-1:0] node43886;
	wire [4-1:0] node43888;
	wire [4-1:0] node43891;
	wire [4-1:0] node43892;
	wire [4-1:0] node43893;
	wire [4-1:0] node43896;
	wire [4-1:0] node43899;
	wire [4-1:0] node43900;
	wire [4-1:0] node43901;
	wire [4-1:0] node43905;
	wire [4-1:0] node43907;
	wire [4-1:0] node43910;
	wire [4-1:0] node43911;
	wire [4-1:0] node43912;
	wire [4-1:0] node43913;
	wire [4-1:0] node43914;
	wire [4-1:0] node43915;
	wire [4-1:0] node43917;
	wire [4-1:0] node43920;
	wire [4-1:0] node43921;
	wire [4-1:0] node43922;
	wire [4-1:0] node43927;
	wire [4-1:0] node43928;
	wire [4-1:0] node43930;
	wire [4-1:0] node43933;
	wire [4-1:0] node43934;
	wire [4-1:0] node43936;
	wire [4-1:0] node43939;
	wire [4-1:0] node43942;
	wire [4-1:0] node43943;
	wire [4-1:0] node43945;
	wire [4-1:0] node43946;
	wire [4-1:0] node43948;
	wire [4-1:0] node43951;
	wire [4-1:0] node43953;
	wire [4-1:0] node43956;
	wire [4-1:0] node43957;
	wire [4-1:0] node43958;
	wire [4-1:0] node43960;
	wire [4-1:0] node43964;
	wire [4-1:0] node43965;
	wire [4-1:0] node43967;
	wire [4-1:0] node43970;
	wire [4-1:0] node43973;
	wire [4-1:0] node43974;
	wire [4-1:0] node43975;
	wire [4-1:0] node43976;
	wire [4-1:0] node43978;
	wire [4-1:0] node43980;
	wire [4-1:0] node43984;
	wire [4-1:0] node43985;
	wire [4-1:0] node43987;
	wire [4-1:0] node43988;
	wire [4-1:0] node43991;
	wire [4-1:0] node43994;
	wire [4-1:0] node43995;
	wire [4-1:0] node43998;
	wire [4-1:0] node44001;
	wire [4-1:0] node44002;
	wire [4-1:0] node44003;
	wire [4-1:0] node44004;
	wire [4-1:0] node44007;
	wire [4-1:0] node44010;
	wire [4-1:0] node44011;
	wire [4-1:0] node44012;
	wire [4-1:0] node44016;
	wire [4-1:0] node44017;
	wire [4-1:0] node44020;
	wire [4-1:0] node44023;
	wire [4-1:0] node44024;
	wire [4-1:0] node44027;
	wire [4-1:0] node44030;
	wire [4-1:0] node44031;
	wire [4-1:0] node44032;
	wire [4-1:0] node44033;
	wire [4-1:0] node44034;
	wire [4-1:0] node44035;
	wire [4-1:0] node44037;
	wire [4-1:0] node44040;
	wire [4-1:0] node44041;
	wire [4-1:0] node44044;
	wire [4-1:0] node44047;
	wire [4-1:0] node44048;
	wire [4-1:0] node44049;
	wire [4-1:0] node44052;
	wire [4-1:0] node44056;
	wire [4-1:0] node44057;
	wire [4-1:0] node44060;
	wire [4-1:0] node44061;
	wire [4-1:0] node44064;
	wire [4-1:0] node44067;
	wire [4-1:0] node44068;
	wire [4-1:0] node44069;
	wire [4-1:0] node44070;
	wire [4-1:0] node44072;
	wire [4-1:0] node44075;
	wire [4-1:0] node44078;
	wire [4-1:0] node44079;
	wire [4-1:0] node44082;
	wire [4-1:0] node44085;
	wire [4-1:0] node44086;
	wire [4-1:0] node44089;
	wire [4-1:0] node44092;
	wire [4-1:0] node44093;
	wire [4-1:0] node44094;
	wire [4-1:0] node44095;
	wire [4-1:0] node44097;
	wire [4-1:0] node44100;
	wire [4-1:0] node44101;
	wire [4-1:0] node44104;
	wire [4-1:0] node44107;
	wire [4-1:0] node44108;
	wire [4-1:0] node44109;
	wire [4-1:0] node44110;
	wire [4-1:0] node44114;
	wire [4-1:0] node44115;
	wire [4-1:0] node44119;
	wire [4-1:0] node44120;
	wire [4-1:0] node44121;
	wire [4-1:0] node44125;
	wire [4-1:0] node44128;
	wire [4-1:0] node44129;
	wire [4-1:0] node44130;
	wire [4-1:0] node44131;
	wire [4-1:0] node44134;
	wire [4-1:0] node44135;
	wire [4-1:0] node44139;
	wire [4-1:0] node44140;
	wire [4-1:0] node44141;
	wire [4-1:0] node44145;
	wire [4-1:0] node44146;
	wire [4-1:0] node44150;
	wire [4-1:0] node44151;
	wire [4-1:0] node44153;
	wire [4-1:0] node44154;
	wire [4-1:0] node44158;
	wire [4-1:0] node44160;
	wire [4-1:0] node44163;
	wire [4-1:0] node44164;
	wire [4-1:0] node44165;
	wire [4-1:0] node44166;
	wire [4-1:0] node44167;
	wire [4-1:0] node44168;
	wire [4-1:0] node44169;
	wire [4-1:0] node44171;
	wire [4-1:0] node44174;
	wire [4-1:0] node44176;
	wire [4-1:0] node44179;
	wire [4-1:0] node44180;
	wire [4-1:0] node44182;
	wire [4-1:0] node44186;
	wire [4-1:0] node44187;
	wire [4-1:0] node44189;
	wire [4-1:0] node44192;
	wire [4-1:0] node44194;
	wire [4-1:0] node44197;
	wire [4-1:0] node44198;
	wire [4-1:0] node44199;
	wire [4-1:0] node44200;
	wire [4-1:0] node44202;
	wire [4-1:0] node44205;
	wire [4-1:0] node44207;
	wire [4-1:0] node44210;
	wire [4-1:0] node44211;
	wire [4-1:0] node44212;
	wire [4-1:0] node44216;
	wire [4-1:0] node44217;
	wire [4-1:0] node44221;
	wire [4-1:0] node44222;
	wire [4-1:0] node44223;
	wire [4-1:0] node44227;
	wire [4-1:0] node44228;
	wire [4-1:0] node44232;
	wire [4-1:0] node44233;
	wire [4-1:0] node44234;
	wire [4-1:0] node44235;
	wire [4-1:0] node44237;
	wire [4-1:0] node44239;
	wire [4-1:0] node44242;
	wire [4-1:0] node44243;
	wire [4-1:0] node44244;
	wire [4-1:0] node44248;
	wire [4-1:0] node44249;
	wire [4-1:0] node44250;
	wire [4-1:0] node44254;
	wire [4-1:0] node44255;
	wire [4-1:0] node44259;
	wire [4-1:0] node44260;
	wire [4-1:0] node44261;
	wire [4-1:0] node44265;
	wire [4-1:0] node44266;
	wire [4-1:0] node44270;
	wire [4-1:0] node44271;
	wire [4-1:0] node44272;
	wire [4-1:0] node44273;
	wire [4-1:0] node44276;
	wire [4-1:0] node44277;
	wire [4-1:0] node44281;
	wire [4-1:0] node44282;
	wire [4-1:0] node44283;
	wire [4-1:0] node44286;
	wire [4-1:0] node44289;
	wire [4-1:0] node44290;
	wire [4-1:0] node44294;
	wire [4-1:0] node44295;
	wire [4-1:0] node44296;
	wire [4-1:0] node44300;
	wire [4-1:0] node44301;
	wire [4-1:0] node44305;
	wire [4-1:0] node44306;
	wire [4-1:0] node44307;
	wire [4-1:0] node44308;
	wire [4-1:0] node44309;
	wire [4-1:0] node44310;
	wire [4-1:0] node44311;
	wire [4-1:0] node44314;
	wire [4-1:0] node44317;
	wire [4-1:0] node44318;
	wire [4-1:0] node44321;
	wire [4-1:0] node44324;
	wire [4-1:0] node44325;
	wire [4-1:0] node44328;
	wire [4-1:0] node44331;
	wire [4-1:0] node44332;
	wire [4-1:0] node44333;
	wire [4-1:0] node44334;
	wire [4-1:0] node44338;
	wire [4-1:0] node44339;
	wire [4-1:0] node44343;
	wire [4-1:0] node44344;
	wire [4-1:0] node44345;
	wire [4-1:0] node44349;
	wire [4-1:0] node44350;
	wire [4-1:0] node44354;
	wire [4-1:0] node44355;
	wire [4-1:0] node44356;
	wire [4-1:0] node44357;
	wire [4-1:0] node44358;
	wire [4-1:0] node44362;
	wire [4-1:0] node44363;
	wire [4-1:0] node44367;
	wire [4-1:0] node44369;
	wire [4-1:0] node44370;
	wire [4-1:0] node44374;
	wire [4-1:0] node44375;
	wire [4-1:0] node44376;
	wire [4-1:0] node44377;
	wire [4-1:0] node44379;
	wire [4-1:0] node44382;
	wire [4-1:0] node44383;
	wire [4-1:0] node44386;
	wire [4-1:0] node44389;
	wire [4-1:0] node44390;
	wire [4-1:0] node44394;
	wire [4-1:0] node44395;
	wire [4-1:0] node44397;
	wire [4-1:0] node44398;
	wire [4-1:0] node44402;
	wire [4-1:0] node44403;
	wire [4-1:0] node44407;
	wire [4-1:0] node44408;
	wire [4-1:0] node44409;
	wire [4-1:0] node44410;
	wire [4-1:0] node44411;
	wire [4-1:0] node44413;
	wire [4-1:0] node44414;
	wire [4-1:0] node44418;
	wire [4-1:0] node44420;
	wire [4-1:0] node44423;
	wire [4-1:0] node44424;
	wire [4-1:0] node44425;
	wire [4-1:0] node44428;
	wire [4-1:0] node44429;
	wire [4-1:0] node44433;
	wire [4-1:0] node44434;
	wire [4-1:0] node44435;
	wire [4-1:0] node44438;
	wire [4-1:0] node44442;
	wire [4-1:0] node44443;
	wire [4-1:0] node44444;
	wire [4-1:0] node44445;
	wire [4-1:0] node44449;
	wire [4-1:0] node44452;
	wire [4-1:0] node44453;
	wire [4-1:0] node44454;
	wire [4-1:0] node44459;
	wire [4-1:0] node44460;
	wire [4-1:0] node44461;
	wire [4-1:0] node44462;
	wire [4-1:0] node44463;
	wire [4-1:0] node44467;
	wire [4-1:0] node44470;
	wire [4-1:0] node44471;
	wire [4-1:0] node44472;
	wire [4-1:0] node44476;
	wire [4-1:0] node44477;
	wire [4-1:0] node44481;
	wire [4-1:0] node44482;
	wire [4-1:0] node44483;
	wire [4-1:0] node44486;
	wire [4-1:0] node44487;
	wire [4-1:0] node44488;
	wire [4-1:0] node44492;
	wire [4-1:0] node44493;
	wire [4-1:0] node44497;
	wire [4-1:0] node44498;
	wire [4-1:0] node44499;
	wire [4-1:0] node44500;
	wire [4-1:0] node44503;
	wire [4-1:0] node44506;
	wire [4-1:0] node44508;
	wire [4-1:0] node44512;
	wire [4-1:0] node44513;
	wire [4-1:0] node44514;
	wire [4-1:0] node44515;
	wire [4-1:0] node44516;
	wire [4-1:0] node44517;
	wire [4-1:0] node44518;
	wire [4-1:0] node44519;
	wire [4-1:0] node44520;
	wire [4-1:0] node44521;
	wire [4-1:0] node44524;
	wire [4-1:0] node44527;
	wire [4-1:0] node44528;
	wire [4-1:0] node44532;
	wire [4-1:0] node44533;
	wire [4-1:0] node44536;
	wire [4-1:0] node44539;
	wire [4-1:0] node44540;
	wire [4-1:0] node44541;
	wire [4-1:0] node44542;
	wire [4-1:0] node44546;
	wire [4-1:0] node44549;
	wire [4-1:0] node44550;
	wire [4-1:0] node44551;
	wire [4-1:0] node44554;
	wire [4-1:0] node44557;
	wire [4-1:0] node44558;
	wire [4-1:0] node44561;
	wire [4-1:0] node44564;
	wire [4-1:0] node44565;
	wire [4-1:0] node44566;
	wire [4-1:0] node44567;
	wire [4-1:0] node44572;
	wire [4-1:0] node44573;
	wire [4-1:0] node44574;
	wire [4-1:0] node44575;
	wire [4-1:0] node44579;
	wire [4-1:0] node44582;
	wire [4-1:0] node44583;
	wire [4-1:0] node44584;
	wire [4-1:0] node44589;
	wire [4-1:0] node44590;
	wire [4-1:0] node44591;
	wire [4-1:0] node44592;
	wire [4-1:0] node44595;
	wire [4-1:0] node44596;
	wire [4-1:0] node44600;
	wire [4-1:0] node44601;
	wire [4-1:0] node44603;
	wire [4-1:0] node44606;
	wire [4-1:0] node44607;
	wire [4-1:0] node44610;
	wire [4-1:0] node44613;
	wire [4-1:0] node44614;
	wire [4-1:0] node44615;
	wire [4-1:0] node44617;
	wire [4-1:0] node44620;
	wire [4-1:0] node44621;
	wire [4-1:0] node44625;
	wire [4-1:0] node44626;
	wire [4-1:0] node44630;
	wire [4-1:0] node44631;
	wire [4-1:0] node44632;
	wire [4-1:0] node44633;
	wire [4-1:0] node44634;
	wire [4-1:0] node44635;
	wire [4-1:0] node44636;
	wire [4-1:0] node44640;
	wire [4-1:0] node44643;
	wire [4-1:0] node44644;
	wire [4-1:0] node44645;
	wire [4-1:0] node44648;
	wire [4-1:0] node44652;
	wire [4-1:0] node44653;
	wire [4-1:0] node44654;
	wire [4-1:0] node44655;
	wire [4-1:0] node44660;
	wire [4-1:0] node44662;
	wire [4-1:0] node44663;
	wire [4-1:0] node44667;
	wire [4-1:0] node44668;
	wire [4-1:0] node44669;
	wire [4-1:0] node44671;
	wire [4-1:0] node44672;
	wire [4-1:0] node44676;
	wire [4-1:0] node44677;
	wire [4-1:0] node44678;
	wire [4-1:0] node44682;
	wire [4-1:0] node44683;
	wire [4-1:0] node44687;
	wire [4-1:0] node44688;
	wire [4-1:0] node44689;
	wire [4-1:0] node44690;
	wire [4-1:0] node44694;
	wire [4-1:0] node44697;
	wire [4-1:0] node44698;
	wire [4-1:0] node44699;
	wire [4-1:0] node44702;
	wire [4-1:0] node44706;
	wire [4-1:0] node44707;
	wire [4-1:0] node44708;
	wire [4-1:0] node44709;
	wire [4-1:0] node44711;
	wire [4-1:0] node44712;
	wire [4-1:0] node44715;
	wire [4-1:0] node44718;
	wire [4-1:0] node44719;
	wire [4-1:0] node44720;
	wire [4-1:0] node44723;
	wire [4-1:0] node44726;
	wire [4-1:0] node44727;
	wire [4-1:0] node44731;
	wire [4-1:0] node44732;
	wire [4-1:0] node44733;
	wire [4-1:0] node44734;
	wire [4-1:0] node44738;
	wire [4-1:0] node44741;
	wire [4-1:0] node44743;
	wire [4-1:0] node44746;
	wire [4-1:0] node44747;
	wire [4-1:0] node44748;
	wire [4-1:0] node44749;
	wire [4-1:0] node44750;
	wire [4-1:0] node44754;
	wire [4-1:0] node44755;
	wire [4-1:0] node44758;
	wire [4-1:0] node44761;
	wire [4-1:0] node44762;
	wire [4-1:0] node44765;
	wire [4-1:0] node44768;
	wire [4-1:0] node44769;
	wire [4-1:0] node44772;
	wire [4-1:0] node44773;
	wire [4-1:0] node44774;
	wire [4-1:0] node44778;
	wire [4-1:0] node44779;
	wire [4-1:0] node44783;
	wire [4-1:0] node44784;
	wire [4-1:0] node44785;
	wire [4-1:0] node44786;
	wire [4-1:0] node44787;
	wire [4-1:0] node44788;
	wire [4-1:0] node44790;
	wire [4-1:0] node44791;
	wire [4-1:0] node44794;
	wire [4-1:0] node44797;
	wire [4-1:0] node44798;
	wire [4-1:0] node44800;
	wire [4-1:0] node44803;
	wire [4-1:0] node44805;
	wire [4-1:0] node44808;
	wire [4-1:0] node44809;
	wire [4-1:0] node44811;
	wire [4-1:0] node44812;
	wire [4-1:0] node44815;
	wire [4-1:0] node44818;
	wire [4-1:0] node44820;
	wire [4-1:0] node44823;
	wire [4-1:0] node44824;
	wire [4-1:0] node44826;
	wire [4-1:0] node44828;
	wire [4-1:0] node44830;
	wire [4-1:0] node44833;
	wire [4-1:0] node44834;
	wire [4-1:0] node44835;
	wire [4-1:0] node44838;
	wire [4-1:0] node44841;
	wire [4-1:0] node44842;
	wire [4-1:0] node44844;
	wire [4-1:0] node44848;
	wire [4-1:0] node44849;
	wire [4-1:0] node44850;
	wire [4-1:0] node44851;
	wire [4-1:0] node44853;
	wire [4-1:0] node44855;
	wire [4-1:0] node44858;
	wire [4-1:0] node44859;
	wire [4-1:0] node44860;
	wire [4-1:0] node44863;
	wire [4-1:0] node44866;
	wire [4-1:0] node44867;
	wire [4-1:0] node44871;
	wire [4-1:0] node44872;
	wire [4-1:0] node44873;
	wire [4-1:0] node44874;
	wire [4-1:0] node44879;
	wire [4-1:0] node44880;
	wire [4-1:0] node44881;
	wire [4-1:0] node44884;
	wire [4-1:0] node44888;
	wire [4-1:0] node44889;
	wire [4-1:0] node44890;
	wire [4-1:0] node44891;
	wire [4-1:0] node44892;
	wire [4-1:0] node44895;
	wire [4-1:0] node44898;
	wire [4-1:0] node44899;
	wire [4-1:0] node44902;
	wire [4-1:0] node44905;
	wire [4-1:0] node44906;
	wire [4-1:0] node44909;
	wire [4-1:0] node44912;
	wire [4-1:0] node44913;
	wire [4-1:0] node44914;
	wire [4-1:0] node44917;
	wire [4-1:0] node44920;
	wire [4-1:0] node44921;
	wire [4-1:0] node44925;
	wire [4-1:0] node44926;
	wire [4-1:0] node44927;
	wire [4-1:0] node44928;
	wire [4-1:0] node44929;
	wire [4-1:0] node44930;
	wire [4-1:0] node44931;
	wire [4-1:0] node44934;
	wire [4-1:0] node44938;
	wire [4-1:0] node44939;
	wire [4-1:0] node44940;
	wire [4-1:0] node44944;
	wire [4-1:0] node44945;
	wire [4-1:0] node44949;
	wire [4-1:0] node44950;
	wire [4-1:0] node44951;
	wire [4-1:0] node44954;
	wire [4-1:0] node44955;
	wire [4-1:0] node44959;
	wire [4-1:0] node44961;
	wire [4-1:0] node44964;
	wire [4-1:0] node44965;
	wire [4-1:0] node44966;
	wire [4-1:0] node44967;
	wire [4-1:0] node44968;
	wire [4-1:0] node44972;
	wire [4-1:0] node44973;
	wire [4-1:0] node44977;
	wire [4-1:0] node44978;
	wire [4-1:0] node44981;
	wire [4-1:0] node44982;
	wire [4-1:0] node44986;
	wire [4-1:0] node44987;
	wire [4-1:0] node44988;
	wire [4-1:0] node44989;
	wire [4-1:0] node44993;
	wire [4-1:0] node44994;
	wire [4-1:0] node44999;
	wire [4-1:0] node45000;
	wire [4-1:0] node45001;
	wire [4-1:0] node45002;
	wire [4-1:0] node45004;
	wire [4-1:0] node45007;
	wire [4-1:0] node45009;
	wire [4-1:0] node45012;
	wire [4-1:0] node45013;
	wire [4-1:0] node45014;
	wire [4-1:0] node45015;
	wire [4-1:0] node45019;
	wire [4-1:0] node45020;
	wire [4-1:0] node45024;
	wire [4-1:0] node45025;
	wire [4-1:0] node45029;
	wire [4-1:0] node45030;
	wire [4-1:0] node45031;
	wire [4-1:0] node45032;
	wire [4-1:0] node45033;
	wire [4-1:0] node45038;
	wire [4-1:0] node45039;
	wire [4-1:0] node45043;
	wire [4-1:0] node45044;
	wire [4-1:0] node45047;
	wire [4-1:0] node45050;
	wire [4-1:0] node45051;
	wire [4-1:0] node45052;
	wire [4-1:0] node45053;
	wire [4-1:0] node45054;
	wire [4-1:0] node45055;
	wire [4-1:0] node45056;
	wire [4-1:0] node45057;
	wire [4-1:0] node45060;
	wire [4-1:0] node45063;
	wire [4-1:0] node45064;
	wire [4-1:0] node45067;
	wire [4-1:0] node45070;
	wire [4-1:0] node45072;
	wire [4-1:0] node45073;
	wire [4-1:0] node45076;
	wire [4-1:0] node45079;
	wire [4-1:0] node45080;
	wire [4-1:0] node45081;
	wire [4-1:0] node45082;
	wire [4-1:0] node45086;
	wire [4-1:0] node45087;
	wire [4-1:0] node45091;
	wire [4-1:0] node45093;
	wire [4-1:0] node45094;
	wire [4-1:0] node45098;
	wire [4-1:0] node45099;
	wire [4-1:0] node45100;
	wire [4-1:0] node45101;
	wire [4-1:0] node45102;
	wire [4-1:0] node45106;
	wire [4-1:0] node45107;
	wire [4-1:0] node45111;
	wire [4-1:0] node45112;
	wire [4-1:0] node45113;
	wire [4-1:0] node45117;
	wire [4-1:0] node45118;
	wire [4-1:0] node45122;
	wire [4-1:0] node45123;
	wire [4-1:0] node45124;
	wire [4-1:0] node45125;
	wire [4-1:0] node45126;
	wire [4-1:0] node45131;
	wire [4-1:0] node45133;
	wire [4-1:0] node45136;
	wire [4-1:0] node45137;
	wire [4-1:0] node45138;
	wire [4-1:0] node45139;
	wire [4-1:0] node45142;
	wire [4-1:0] node45145;
	wire [4-1:0] node45146;
	wire [4-1:0] node45149;
	wire [4-1:0] node45152;
	wire [4-1:0] node45154;
	wire [4-1:0] node45157;
	wire [4-1:0] node45158;
	wire [4-1:0] node45159;
	wire [4-1:0] node45160;
	wire [4-1:0] node45161;
	wire [4-1:0] node45163;
	wire [4-1:0] node45166;
	wire [4-1:0] node45167;
	wire [4-1:0] node45170;
	wire [4-1:0] node45173;
	wire [4-1:0] node45174;
	wire [4-1:0] node45177;
	wire [4-1:0] node45180;
	wire [4-1:0] node45181;
	wire [4-1:0] node45182;
	wire [4-1:0] node45183;
	wire [4-1:0] node45187;
	wire [4-1:0] node45188;
	wire [4-1:0] node45192;
	wire [4-1:0] node45193;
	wire [4-1:0] node45194;
	wire [4-1:0] node45198;
	wire [4-1:0] node45199;
	wire [4-1:0] node45203;
	wire [4-1:0] node45204;
	wire [4-1:0] node45205;
	wire [4-1:0] node45206;
	wire [4-1:0] node45207;
	wire [4-1:0] node45211;
	wire [4-1:0] node45212;
	wire [4-1:0] node45216;
	wire [4-1:0] node45217;
	wire [4-1:0] node45218;
	wire [4-1:0] node45222;
	wire [4-1:0] node45223;
	wire [4-1:0] node45227;
	wire [4-1:0] node45228;
	wire [4-1:0] node45229;
	wire [4-1:0] node45230;
	wire [4-1:0] node45234;
	wire [4-1:0] node45235;
	wire [4-1:0] node45239;
	wire [4-1:0] node45240;
	wire [4-1:0] node45241;
	wire [4-1:0] node45245;
	wire [4-1:0] node45246;
	wire [4-1:0] node45250;
	wire [4-1:0] node45251;
	wire [4-1:0] node45252;
	wire [4-1:0] node45253;
	wire [4-1:0] node45254;
	wire [4-1:0] node45255;
	wire [4-1:0] node45256;
	wire [4-1:0] node45257;
	wire [4-1:0] node45260;
	wire [4-1:0] node45263;
	wire [4-1:0] node45264;
	wire [4-1:0] node45267;
	wire [4-1:0] node45270;
	wire [4-1:0] node45271;
	wire [4-1:0] node45272;
	wire [4-1:0] node45276;
	wire [4-1:0] node45279;
	wire [4-1:0] node45280;
	wire [4-1:0] node45282;
	wire [4-1:0] node45283;
	wire [4-1:0] node45287;
	wire [4-1:0] node45288;
	wire [4-1:0] node45289;
	wire [4-1:0] node45293;
	wire [4-1:0] node45296;
	wire [4-1:0] node45297;
	wire [4-1:0] node45298;
	wire [4-1:0] node45299;
	wire [4-1:0] node45303;
	wire [4-1:0] node45304;
	wire [4-1:0] node45305;
	wire [4-1:0] node45309;
	wire [4-1:0] node45310;
	wire [4-1:0] node45314;
	wire [4-1:0] node45315;
	wire [4-1:0] node45316;
	wire [4-1:0] node45317;
	wire [4-1:0] node45320;
	wire [4-1:0] node45324;
	wire [4-1:0] node45325;
	wire [4-1:0] node45328;
	wire [4-1:0] node45331;
	wire [4-1:0] node45332;
	wire [4-1:0] node45333;
	wire [4-1:0] node45334;
	wire [4-1:0] node45335;
	wire [4-1:0] node45336;
	wire [4-1:0] node45341;
	wire [4-1:0] node45342;
	wire [4-1:0] node45346;
	wire [4-1:0] node45347;
	wire [4-1:0] node45348;
	wire [4-1:0] node45351;
	wire [4-1:0] node45352;
	wire [4-1:0] node45356;
	wire [4-1:0] node45357;
	wire [4-1:0] node45358;
	wire [4-1:0] node45361;
	wire [4-1:0] node45365;
	wire [4-1:0] node45366;
	wire [4-1:0] node45367;
	wire [4-1:0] node45368;
	wire [4-1:0] node45369;
	wire [4-1:0] node45374;
	wire [4-1:0] node45375;
	wire [4-1:0] node45376;
	wire [4-1:0] node45381;
	wire [4-1:0] node45382;
	wire [4-1:0] node45383;
	wire [4-1:0] node45387;
	wire [4-1:0] node45388;
	wire [4-1:0] node45392;
	wire [4-1:0] node45393;
	wire [4-1:0] node45394;
	wire [4-1:0] node45395;
	wire [4-1:0] node45396;
	wire [4-1:0] node45397;
	wire [4-1:0] node45398;
	wire [4-1:0] node45401;
	wire [4-1:0] node45404;
	wire [4-1:0] node45405;
	wire [4-1:0] node45408;
	wire [4-1:0] node45411;
	wire [4-1:0] node45412;
	wire [4-1:0] node45415;
	wire [4-1:0] node45418;
	wire [4-1:0] node45419;
	wire [4-1:0] node45420;
	wire [4-1:0] node45421;
	wire [4-1:0] node45425;
	wire [4-1:0] node45428;
	wire [4-1:0] node45430;
	wire [4-1:0] node45433;
	wire [4-1:0] node45434;
	wire [4-1:0] node45435;
	wire [4-1:0] node45437;
	wire [4-1:0] node45438;
	wire [4-1:0] node45442;
	wire [4-1:0] node45443;
	wire [4-1:0] node45444;
	wire [4-1:0] node45448;
	wire [4-1:0] node45449;
	wire [4-1:0] node45453;
	wire [4-1:0] node45454;
	wire [4-1:0] node45456;
	wire [4-1:0] node45457;
	wire [4-1:0] node45461;
	wire [4-1:0] node45463;
	wire [4-1:0] node45466;
	wire [4-1:0] node45467;
	wire [4-1:0] node45468;
	wire [4-1:0] node45469;
	wire [4-1:0] node45470;
	wire [4-1:0] node45471;
	wire [4-1:0] node45475;
	wire [4-1:0] node45478;
	wire [4-1:0] node45479;
	wire [4-1:0] node45482;
	wire [4-1:0] node45483;
	wire [4-1:0] node45487;
	wire [4-1:0] node45488;
	wire [4-1:0] node45490;
	wire [4-1:0] node45493;
	wire [4-1:0] node45495;
	wire [4-1:0] node45496;
	wire [4-1:0] node45500;
	wire [4-1:0] node45501;
	wire [4-1:0] node45502;
	wire [4-1:0] node45504;
	wire [4-1:0] node45507;
	wire [4-1:0] node45508;
	wire [4-1:0] node45509;
	wire [4-1:0] node45514;
	wire [4-1:0] node45515;
	wire [4-1:0] node45516;
	wire [4-1:0] node45517;
	wire [4-1:0] node45520;
	wire [4-1:0] node45523;
	wire [4-1:0] node45524;
	wire [4-1:0] node45527;
	wire [4-1:0] node45530;
	wire [4-1:0] node45532;
	wire [4-1:0] node45533;
	wire [4-1:0] node45536;
	wire [4-1:0] node45539;
	wire [4-1:0] node45540;
	wire [4-1:0] node45541;
	wire [4-1:0] node45542;
	wire [4-1:0] node45543;
	wire [4-1:0] node45544;
	wire [4-1:0] node45545;
	wire [4-1:0] node45546;
	wire [4-1:0] node45547;
	wire [4-1:0] node45548;
	wire [4-1:0] node45550;
	wire [4-1:0] node45551;
	wire [4-1:0] node45554;
	wire [4-1:0] node45557;
	wire [4-1:0] node45558;
	wire [4-1:0] node45559;
	wire [4-1:0] node45563;
	wire [4-1:0] node45564;
	wire [4-1:0] node45567;
	wire [4-1:0] node45570;
	wire [4-1:0] node45571;
	wire [4-1:0] node45572;
	wire [4-1:0] node45573;
	wire [4-1:0] node45577;
	wire [4-1:0] node45579;
	wire [4-1:0] node45582;
	wire [4-1:0] node45583;
	wire [4-1:0] node45584;
	wire [4-1:0] node45588;
	wire [4-1:0] node45589;
	wire [4-1:0] node45593;
	wire [4-1:0] node45594;
	wire [4-1:0] node45595;
	wire [4-1:0] node45596;
	wire [4-1:0] node45599;
	wire [4-1:0] node45602;
	wire [4-1:0] node45603;
	wire [4-1:0] node45606;
	wire [4-1:0] node45609;
	wire [4-1:0] node45610;
	wire [4-1:0] node45611;
	wire [4-1:0] node45614;
	wire [4-1:0] node45617;
	wire [4-1:0] node45618;
	wire [4-1:0] node45621;
	wire [4-1:0] node45624;
	wire [4-1:0] node45625;
	wire [4-1:0] node45626;
	wire [4-1:0] node45627;
	wire [4-1:0] node45628;
	wire [4-1:0] node45629;
	wire [4-1:0] node45633;
	wire [4-1:0] node45634;
	wire [4-1:0] node45638;
	wire [4-1:0] node45639;
	wire [4-1:0] node45640;
	wire [4-1:0] node45643;
	wire [4-1:0] node45646;
	wire [4-1:0] node45649;
	wire [4-1:0] node45650;
	wire [4-1:0] node45651;
	wire [4-1:0] node45653;
	wire [4-1:0] node45656;
	wire [4-1:0] node45657;
	wire [4-1:0] node45660;
	wire [4-1:0] node45663;
	wire [4-1:0] node45664;
	wire [4-1:0] node45665;
	wire [4-1:0] node45668;
	wire [4-1:0] node45671;
	wire [4-1:0] node45672;
	wire [4-1:0] node45676;
	wire [4-1:0] node45677;
	wire [4-1:0] node45678;
	wire [4-1:0] node45679;
	wire [4-1:0] node45682;
	wire [4-1:0] node45685;
	wire [4-1:0] node45687;
	wire [4-1:0] node45688;
	wire [4-1:0] node45692;
	wire [4-1:0] node45693;
	wire [4-1:0] node45694;
	wire [4-1:0] node45697;
	wire [4-1:0] node45699;
	wire [4-1:0] node45702;
	wire [4-1:0] node45703;
	wire [4-1:0] node45706;
	wire [4-1:0] node45709;
	wire [4-1:0] node45710;
	wire [4-1:0] node45711;
	wire [4-1:0] node45712;
	wire [4-1:0] node45713;
	wire [4-1:0] node45715;
	wire [4-1:0] node45716;
	wire [4-1:0] node45720;
	wire [4-1:0] node45721;
	wire [4-1:0] node45724;
	wire [4-1:0] node45727;
	wire [4-1:0] node45728;
	wire [4-1:0] node45729;
	wire [4-1:0] node45730;
	wire [4-1:0] node45734;
	wire [4-1:0] node45735;
	wire [4-1:0] node45738;
	wire [4-1:0] node45741;
	wire [4-1:0] node45742;
	wire [4-1:0] node45745;
	wire [4-1:0] node45748;
	wire [4-1:0] node45749;
	wire [4-1:0] node45750;
	wire [4-1:0] node45751;
	wire [4-1:0] node45752;
	wire [4-1:0] node45755;
	wire [4-1:0] node45758;
	wire [4-1:0] node45759;
	wire [4-1:0] node45762;
	wire [4-1:0] node45765;
	wire [4-1:0] node45766;
	wire [4-1:0] node45769;
	wire [4-1:0] node45772;
	wire [4-1:0] node45773;
	wire [4-1:0] node45774;
	wire [4-1:0] node45775;
	wire [4-1:0] node45778;
	wire [4-1:0] node45781;
	wire [4-1:0] node45783;
	wire [4-1:0] node45786;
	wire [4-1:0] node45788;
	wire [4-1:0] node45791;
	wire [4-1:0] node45792;
	wire [4-1:0] node45793;
	wire [4-1:0] node45794;
	wire [4-1:0] node45795;
	wire [4-1:0] node45798;
	wire [4-1:0] node45801;
	wire [4-1:0] node45802;
	wire [4-1:0] node45806;
	wire [4-1:0] node45807;
	wire [4-1:0] node45808;
	wire [4-1:0] node45810;
	wire [4-1:0] node45813;
	wire [4-1:0] node45814;
	wire [4-1:0] node45817;
	wire [4-1:0] node45820;
	wire [4-1:0] node45822;
	wire [4-1:0] node45825;
	wire [4-1:0] node45826;
	wire [4-1:0] node45827;
	wire [4-1:0] node45828;
	wire [4-1:0] node45829;
	wire [4-1:0] node45832;
	wire [4-1:0] node45835;
	wire [4-1:0] node45836;
	wire [4-1:0] node45840;
	wire [4-1:0] node45841;
	wire [4-1:0] node45844;
	wire [4-1:0] node45847;
	wire [4-1:0] node45848;
	wire [4-1:0] node45849;
	wire [4-1:0] node45850;
	wire [4-1:0] node45855;
	wire [4-1:0] node45858;
	wire [4-1:0] node45859;
	wire [4-1:0] node45860;
	wire [4-1:0] node45861;
	wire [4-1:0] node45862;
	wire [4-1:0] node45863;
	wire [4-1:0] node45864;
	wire [4-1:0] node45866;
	wire [4-1:0] node45869;
	wire [4-1:0] node45870;
	wire [4-1:0] node45873;
	wire [4-1:0] node45876;
	wire [4-1:0] node45877;
	wire [4-1:0] node45880;
	wire [4-1:0] node45883;
	wire [4-1:0] node45884;
	wire [4-1:0] node45886;
	wire [4-1:0] node45889;
	wire [4-1:0] node45890;
	wire [4-1:0] node45891;
	wire [4-1:0] node45895;
	wire [4-1:0] node45898;
	wire [4-1:0] node45899;
	wire [4-1:0] node45900;
	wire [4-1:0] node45901;
	wire [4-1:0] node45904;
	wire [4-1:0] node45907;
	wire [4-1:0] node45908;
	wire [4-1:0] node45911;
	wire [4-1:0] node45914;
	wire [4-1:0] node45915;
	wire [4-1:0] node45916;
	wire [4-1:0] node45917;
	wire [4-1:0] node45920;
	wire [4-1:0] node45924;
	wire [4-1:0] node45925;
	wire [4-1:0] node45928;
	wire [4-1:0] node45931;
	wire [4-1:0] node45932;
	wire [4-1:0] node45933;
	wire [4-1:0] node45934;
	wire [4-1:0] node45936;
	wire [4-1:0] node45937;
	wire [4-1:0] node45941;
	wire [4-1:0] node45944;
	wire [4-1:0] node45945;
	wire [4-1:0] node45946;
	wire [4-1:0] node45947;
	wire [4-1:0] node45951;
	wire [4-1:0] node45953;
	wire [4-1:0] node45956;
	wire [4-1:0] node45957;
	wire [4-1:0] node45960;
	wire [4-1:0] node45963;
	wire [4-1:0] node45964;
	wire [4-1:0] node45965;
	wire [4-1:0] node45966;
	wire [4-1:0] node45970;
	wire [4-1:0] node45971;
	wire [4-1:0] node45974;
	wire [4-1:0] node45977;
	wire [4-1:0] node45978;
	wire [4-1:0] node45979;
	wire [4-1:0] node45980;
	wire [4-1:0] node45983;
	wire [4-1:0] node45986;
	wire [4-1:0] node45988;
	wire [4-1:0] node45991;
	wire [4-1:0] node45992;
	wire [4-1:0] node45993;
	wire [4-1:0] node45996;
	wire [4-1:0] node45999;
	wire [4-1:0] node46000;
	wire [4-1:0] node46003;
	wire [4-1:0] node46006;
	wire [4-1:0] node46007;
	wire [4-1:0] node46008;
	wire [4-1:0] node46009;
	wire [4-1:0] node46010;
	wire [4-1:0] node46012;
	wire [4-1:0] node46013;
	wire [4-1:0] node46018;
	wire [4-1:0] node46019;
	wire [4-1:0] node46020;
	wire [4-1:0] node46021;
	wire [4-1:0] node46025;
	wire [4-1:0] node46026;
	wire [4-1:0] node46030;
	wire [4-1:0] node46031;
	wire [4-1:0] node46032;
	wire [4-1:0] node46036;
	wire [4-1:0] node46037;
	wire [4-1:0] node46041;
	wire [4-1:0] node46042;
	wire [4-1:0] node46044;
	wire [4-1:0] node46045;
	wire [4-1:0] node46046;
	wire [4-1:0] node46050;
	wire [4-1:0] node46053;
	wire [4-1:0] node46054;
	wire [4-1:0] node46055;
	wire [4-1:0] node46056;
	wire [4-1:0] node46061;
	wire [4-1:0] node46062;
	wire [4-1:0] node46063;
	wire [4-1:0] node46068;
	wire [4-1:0] node46069;
	wire [4-1:0] node46070;
	wire [4-1:0] node46071;
	wire [4-1:0] node46072;
	wire [4-1:0] node46073;
	wire [4-1:0] node46078;
	wire [4-1:0] node46079;
	wire [4-1:0] node46083;
	wire [4-1:0] node46084;
	wire [4-1:0] node46085;
	wire [4-1:0] node46086;
	wire [4-1:0] node46091;
	wire [4-1:0] node46092;
	wire [4-1:0] node46095;
	wire [4-1:0] node46096;
	wire [4-1:0] node46100;
	wire [4-1:0] node46101;
	wire [4-1:0] node46102;
	wire [4-1:0] node46103;
	wire [4-1:0] node46104;
	wire [4-1:0] node46108;
	wire [4-1:0] node46111;
	wire [4-1:0] node46112;
	wire [4-1:0] node46113;
	wire [4-1:0] node46117;
	wire [4-1:0] node46118;
	wire [4-1:0] node46122;
	wire [4-1:0] node46123;
	wire [4-1:0] node46124;
	wire [4-1:0] node46125;
	wire [4-1:0] node46129;
	wire [4-1:0] node46132;
	wire [4-1:0] node46134;
	wire [4-1:0] node46135;
	wire [4-1:0] node46139;
	wire [4-1:0] node46140;
	wire [4-1:0] node46141;
	wire [4-1:0] node46142;
	wire [4-1:0] node46143;
	wire [4-1:0] node46144;
	wire [4-1:0] node46146;
	wire [4-1:0] node46147;
	wire [4-1:0] node46151;
	wire [4-1:0] node46152;
	wire [4-1:0] node46154;
	wire [4-1:0] node46156;
	wire [4-1:0] node46159;
	wire [4-1:0] node46161;
	wire [4-1:0] node46162;
	wire [4-1:0] node46165;
	wire [4-1:0] node46168;
	wire [4-1:0] node46169;
	wire [4-1:0] node46170;
	wire [4-1:0] node46171;
	wire [4-1:0] node46173;
	wire [4-1:0] node46176;
	wire [4-1:0] node46177;
	wire [4-1:0] node46180;
	wire [4-1:0] node46183;
	wire [4-1:0] node46184;
	wire [4-1:0] node46188;
	wire [4-1:0] node46189;
	wire [4-1:0] node46190;
	wire [4-1:0] node46193;
	wire [4-1:0] node46196;
	wire [4-1:0] node46198;
	wire [4-1:0] node46200;
	wire [4-1:0] node46203;
	wire [4-1:0] node46204;
	wire [4-1:0] node46205;
	wire [4-1:0] node46206;
	wire [4-1:0] node46207;
	wire [4-1:0] node46208;
	wire [4-1:0] node46211;
	wire [4-1:0] node46215;
	wire [4-1:0] node46216;
	wire [4-1:0] node46218;
	wire [4-1:0] node46221;
	wire [4-1:0] node46223;
	wire [4-1:0] node46226;
	wire [4-1:0] node46227;
	wire [4-1:0] node46228;
	wire [4-1:0] node46232;
	wire [4-1:0] node46233;
	wire [4-1:0] node46236;
	wire [4-1:0] node46239;
	wire [4-1:0] node46240;
	wire [4-1:0] node46241;
	wire [4-1:0] node46242;
	wire [4-1:0] node46243;
	wire [4-1:0] node46247;
	wire [4-1:0] node46248;
	wire [4-1:0] node46252;
	wire [4-1:0] node46254;
	wire [4-1:0] node46255;
	wire [4-1:0] node46258;
	wire [4-1:0] node46261;
	wire [4-1:0] node46262;
	wire [4-1:0] node46263;
	wire [4-1:0] node46266;
	wire [4-1:0] node46269;
	wire [4-1:0] node46270;
	wire [4-1:0] node46273;
	wire [4-1:0] node46276;
	wire [4-1:0] node46277;
	wire [4-1:0] node46278;
	wire [4-1:0] node46279;
	wire [4-1:0] node46280;
	wire [4-1:0] node46281;
	wire [4-1:0] node46282;
	wire [4-1:0] node46285;
	wire [4-1:0] node46289;
	wire [4-1:0] node46290;
	wire [4-1:0] node46291;
	wire [4-1:0] node46294;
	wire [4-1:0] node46298;
	wire [4-1:0] node46299;
	wire [4-1:0] node46300;
	wire [4-1:0] node46301;
	wire [4-1:0] node46305;
	wire [4-1:0] node46306;
	wire [4-1:0] node46309;
	wire [4-1:0] node46312;
	wire [4-1:0] node46313;
	wire [4-1:0] node46314;
	wire [4-1:0] node46317;
	wire [4-1:0] node46320;
	wire [4-1:0] node46321;
	wire [4-1:0] node46325;
	wire [4-1:0] node46326;
	wire [4-1:0] node46327;
	wire [4-1:0] node46329;
	wire [4-1:0] node46330;
	wire [4-1:0] node46334;
	wire [4-1:0] node46335;
	wire [4-1:0] node46338;
	wire [4-1:0] node46341;
	wire [4-1:0] node46343;
	wire [4-1:0] node46344;
	wire [4-1:0] node46345;
	wire [4-1:0] node46350;
	wire [4-1:0] node46351;
	wire [4-1:0] node46352;
	wire [4-1:0] node46353;
	wire [4-1:0] node46355;
	wire [4-1:0] node46356;
	wire [4-1:0] node46359;
	wire [4-1:0] node46362;
	wire [4-1:0] node46363;
	wire [4-1:0] node46364;
	wire [4-1:0] node46367;
	wire [4-1:0] node46370;
	wire [4-1:0] node46372;
	wire [4-1:0] node46375;
	wire [4-1:0] node46376;
	wire [4-1:0] node46379;
	wire [4-1:0] node46380;
	wire [4-1:0] node46381;
	wire [4-1:0] node46385;
	wire [4-1:0] node46388;
	wire [4-1:0] node46389;
	wire [4-1:0] node46390;
	wire [4-1:0] node46391;
	wire [4-1:0] node46392;
	wire [4-1:0] node46396;
	wire [4-1:0] node46397;
	wire [4-1:0] node46401;
	wire [4-1:0] node46402;
	wire [4-1:0] node46404;
	wire [4-1:0] node46407;
	wire [4-1:0] node46408;
	wire [4-1:0] node46411;
	wire [4-1:0] node46414;
	wire [4-1:0] node46415;
	wire [4-1:0] node46416;
	wire [4-1:0] node46417;
	wire [4-1:0] node46420;
	wire [4-1:0] node46424;
	wire [4-1:0] node46425;
	wire [4-1:0] node46426;
	wire [4-1:0] node46431;
	wire [4-1:0] node46432;
	wire [4-1:0] node46433;
	wire [4-1:0] node46434;
	wire [4-1:0] node46435;
	wire [4-1:0] node46436;
	wire [4-1:0] node46437;
	wire [4-1:0] node46438;
	wire [4-1:0] node46441;
	wire [4-1:0] node46445;
	wire [4-1:0] node46446;
	wire [4-1:0] node46448;
	wire [4-1:0] node46451;
	wire [4-1:0] node46452;
	wire [4-1:0] node46456;
	wire [4-1:0] node46457;
	wire [4-1:0] node46458;
	wire [4-1:0] node46459;
	wire [4-1:0] node46462;
	wire [4-1:0] node46465;
	wire [4-1:0] node46466;
	wire [4-1:0] node46469;
	wire [4-1:0] node46472;
	wire [4-1:0] node46473;
	wire [4-1:0] node46475;
	wire [4-1:0] node46478;
	wire [4-1:0] node46479;
	wire [4-1:0] node46482;
	wire [4-1:0] node46485;
	wire [4-1:0] node46486;
	wire [4-1:0] node46487;
	wire [4-1:0] node46488;
	wire [4-1:0] node46490;
	wire [4-1:0] node46493;
	wire [4-1:0] node46494;
	wire [4-1:0] node46498;
	wire [4-1:0] node46499;
	wire [4-1:0] node46500;
	wire [4-1:0] node46503;
	wire [4-1:0] node46506;
	wire [4-1:0] node46509;
	wire [4-1:0] node46510;
	wire [4-1:0] node46511;
	wire [4-1:0] node46512;
	wire [4-1:0] node46516;
	wire [4-1:0] node46517;
	wire [4-1:0] node46521;
	wire [4-1:0] node46522;
	wire [4-1:0] node46523;
	wire [4-1:0] node46526;
	wire [4-1:0] node46529;
	wire [4-1:0] node46530;
	wire [4-1:0] node46533;
	wire [4-1:0] node46536;
	wire [4-1:0] node46537;
	wire [4-1:0] node46538;
	wire [4-1:0] node46540;
	wire [4-1:0] node46541;
	wire [4-1:0] node46542;
	wire [4-1:0] node46546;
	wire [4-1:0] node46549;
	wire [4-1:0] node46550;
	wire [4-1:0] node46551;
	wire [4-1:0] node46555;
	wire [4-1:0] node46556;
	wire [4-1:0] node46557;
	wire [4-1:0] node46560;
	wire [4-1:0] node46564;
	wire [4-1:0] node46565;
	wire [4-1:0] node46566;
	wire [4-1:0] node46568;
	wire [4-1:0] node46571;
	wire [4-1:0] node46572;
	wire [4-1:0] node46575;
	wire [4-1:0] node46578;
	wire [4-1:0] node46579;
	wire [4-1:0] node46580;
	wire [4-1:0] node46581;
	wire [4-1:0] node46584;
	wire [4-1:0] node46587;
	wire [4-1:0] node46588;
	wire [4-1:0] node46591;
	wire [4-1:0] node46594;
	wire [4-1:0] node46595;
	wire [4-1:0] node46598;
	wire [4-1:0] node46601;
	wire [4-1:0] node46602;
	wire [4-1:0] node46603;
	wire [4-1:0] node46604;
	wire [4-1:0] node46605;
	wire [4-1:0] node46606;
	wire [4-1:0] node46607;
	wire [4-1:0] node46610;
	wire [4-1:0] node46613;
	wire [4-1:0] node46615;
	wire [4-1:0] node46618;
	wire [4-1:0] node46619;
	wire [4-1:0] node46622;
	wire [4-1:0] node46625;
	wire [4-1:0] node46626;
	wire [4-1:0] node46627;
	wire [4-1:0] node46628;
	wire [4-1:0] node46632;
	wire [4-1:0] node46633;
	wire [4-1:0] node46637;
	wire [4-1:0] node46638;
	wire [4-1:0] node46639;
	wire [4-1:0] node46643;
	wire [4-1:0] node46644;
	wire [4-1:0] node46648;
	wire [4-1:0] node46649;
	wire [4-1:0] node46650;
	wire [4-1:0] node46651;
	wire [4-1:0] node46652;
	wire [4-1:0] node46655;
	wire [4-1:0] node46658;
	wire [4-1:0] node46659;
	wire [4-1:0] node46663;
	wire [4-1:0] node46664;
	wire [4-1:0] node46667;
	wire [4-1:0] node46670;
	wire [4-1:0] node46671;
	wire [4-1:0] node46673;
	wire [4-1:0] node46674;
	wire [4-1:0] node46678;
	wire [4-1:0] node46679;
	wire [4-1:0] node46682;
	wire [4-1:0] node46685;
	wire [4-1:0] node46686;
	wire [4-1:0] node46688;
	wire [4-1:0] node46689;
	wire [4-1:0] node46691;
	wire [4-1:0] node46694;
	wire [4-1:0] node46695;
	wire [4-1:0] node46698;
	wire [4-1:0] node46701;
	wire [4-1:0] node46702;
	wire [4-1:0] node46703;
	wire [4-1:0] node46704;
	wire [4-1:0] node46705;
	wire [4-1:0] node46708;
	wire [4-1:0] node46712;
	wire [4-1:0] node46713;
	wire [4-1:0] node46717;
	wire [4-1:0] node46718;
	wire [4-1:0] node46720;
	wire [4-1:0] node46723;
	wire [4-1:0] node46724;
	wire [4-1:0] node46725;
	wire [4-1:0] node46729;
	wire [4-1:0] node46732;
	wire [4-1:0] node46733;
	wire [4-1:0] node46734;
	wire [4-1:0] node46735;
	wire [4-1:0] node46736;
	wire [4-1:0] node46737;
	wire [4-1:0] node46738;
	wire [4-1:0] node46739;
	wire [4-1:0] node46740;
	wire [4-1:0] node46743;
	wire [4-1:0] node46744;
	wire [4-1:0] node46747;
	wire [4-1:0] node46750;
	wire [4-1:0] node46751;
	wire [4-1:0] node46752;
	wire [4-1:0] node46757;
	wire [4-1:0] node46758;
	wire [4-1:0] node46759;
	wire [4-1:0] node46760;
	wire [4-1:0] node46763;
	wire [4-1:0] node46766;
	wire [4-1:0] node46767;
	wire [4-1:0] node46771;
	wire [4-1:0] node46772;
	wire [4-1:0] node46774;
	wire [4-1:0] node46777;
	wire [4-1:0] node46778;
	wire [4-1:0] node46781;
	wire [4-1:0] node46784;
	wire [4-1:0] node46785;
	wire [4-1:0] node46786;
	wire [4-1:0] node46788;
	wire [4-1:0] node46789;
	wire [4-1:0] node46792;
	wire [4-1:0] node46795;
	wire [4-1:0] node46796;
	wire [4-1:0] node46797;
	wire [4-1:0] node46800;
	wire [4-1:0] node46803;
	wire [4-1:0] node46804;
	wire [4-1:0] node46807;
	wire [4-1:0] node46810;
	wire [4-1:0] node46811;
	wire [4-1:0] node46812;
	wire [4-1:0] node46813;
	wire [4-1:0] node46816;
	wire [4-1:0] node46819;
	wire [4-1:0] node46821;
	wire [4-1:0] node46824;
	wire [4-1:0] node46825;
	wire [4-1:0] node46826;
	wire [4-1:0] node46830;
	wire [4-1:0] node46831;
	wire [4-1:0] node46834;
	wire [4-1:0] node46837;
	wire [4-1:0] node46838;
	wire [4-1:0] node46839;
	wire [4-1:0] node46840;
	wire [4-1:0] node46841;
	wire [4-1:0] node46842;
	wire [4-1:0] node46845;
	wire [4-1:0] node46848;
	wire [4-1:0] node46851;
	wire [4-1:0] node46852;
	wire [4-1:0] node46854;
	wire [4-1:0] node46857;
	wire [4-1:0] node46860;
	wire [4-1:0] node46861;
	wire [4-1:0] node46864;
	wire [4-1:0] node46865;
	wire [4-1:0] node46866;
	wire [4-1:0] node46869;
	wire [4-1:0] node46873;
	wire [4-1:0] node46874;
	wire [4-1:0] node46875;
	wire [4-1:0] node46878;
	wire [4-1:0] node46879;
	wire [4-1:0] node46882;
	wire [4-1:0] node46885;
	wire [4-1:0] node46886;
	wire [4-1:0] node46887;
	wire [4-1:0] node46890;
	wire [4-1:0] node46893;
	wire [4-1:0] node46894;
	wire [4-1:0] node46897;
	wire [4-1:0] node46900;
	wire [4-1:0] node46901;
	wire [4-1:0] node46902;
	wire [4-1:0] node46903;
	wire [4-1:0] node46904;
	wire [4-1:0] node46905;
	wire [4-1:0] node46906;
	wire [4-1:0] node46909;
	wire [4-1:0] node46913;
	wire [4-1:0] node46914;
	wire [4-1:0] node46915;
	wire [4-1:0] node46919;
	wire [4-1:0] node46920;
	wire [4-1:0] node46923;
	wire [4-1:0] node46926;
	wire [4-1:0] node46927;
	wire [4-1:0] node46930;
	wire [4-1:0] node46931;
	wire [4-1:0] node46932;
	wire [4-1:0] node46935;
	wire [4-1:0] node46938;
	wire [4-1:0] node46940;
	wire [4-1:0] node46943;
	wire [4-1:0] node46944;
	wire [4-1:0] node46945;
	wire [4-1:0] node46946;
	wire [4-1:0] node46947;
	wire [4-1:0] node46950;
	wire [4-1:0] node46953;
	wire [4-1:0] node46956;
	wire [4-1:0] node46957;
	wire [4-1:0] node46960;
	wire [4-1:0] node46962;
	wire [4-1:0] node46965;
	wire [4-1:0] node46966;
	wire [4-1:0] node46967;
	wire [4-1:0] node46968;
	wire [4-1:0] node46971;
	wire [4-1:0] node46974;
	wire [4-1:0] node46976;
	wire [4-1:0] node46979;
	wire [4-1:0] node46980;
	wire [4-1:0] node46983;
	wire [4-1:0] node46984;
	wire [4-1:0] node46988;
	wire [4-1:0] node46989;
	wire [4-1:0] node46990;
	wire [4-1:0] node46991;
	wire [4-1:0] node46992;
	wire [4-1:0] node46994;
	wire [4-1:0] node46997;
	wire [4-1:0] node46999;
	wire [4-1:0] node47002;
	wire [4-1:0] node47003;
	wire [4-1:0] node47004;
	wire [4-1:0] node47009;
	wire [4-1:0] node47010;
	wire [4-1:0] node47011;
	wire [4-1:0] node47014;
	wire [4-1:0] node47015;
	wire [4-1:0] node47018;
	wire [4-1:0] node47021;
	wire [4-1:0] node47022;
	wire [4-1:0] node47023;
	wire [4-1:0] node47027;
	wire [4-1:0] node47030;
	wire [4-1:0] node47031;
	wire [4-1:0] node47032;
	wire [4-1:0] node47034;
	wire [4-1:0] node47035;
	wire [4-1:0] node47038;
	wire [4-1:0] node47041;
	wire [4-1:0] node47042;
	wire [4-1:0] node47043;
	wire [4-1:0] node47046;
	wire [4-1:0] node47050;
	wire [4-1:0] node47051;
	wire [4-1:0] node47053;
	wire [4-1:0] node47054;
	wire [4-1:0] node47058;
	wire [4-1:0] node47059;
	wire [4-1:0] node47061;
	wire [4-1:0] node47064;
	wire [4-1:0] node47065;
	wire [4-1:0] node47068;
	wire [4-1:0] node47071;
	wire [4-1:0] node47072;
	wire [4-1:0] node47073;
	wire [4-1:0] node47074;
	wire [4-1:0] node47075;
	wire [4-1:0] node47076;
	wire [4-1:0] node47077;
	wire [4-1:0] node47078;
	wire [4-1:0] node47081;
	wire [4-1:0] node47085;
	wire [4-1:0] node47086;
	wire [4-1:0] node47087;
	wire [4-1:0] node47090;
	wire [4-1:0] node47093;
	wire [4-1:0] node47094;
	wire [4-1:0] node47097;
	wire [4-1:0] node47100;
	wire [4-1:0] node47101;
	wire [4-1:0] node47102;
	wire [4-1:0] node47104;
	wire [4-1:0] node47108;
	wire [4-1:0] node47109;
	wire [4-1:0] node47111;
	wire [4-1:0] node47114;
	wire [4-1:0] node47115;
	wire [4-1:0] node47118;
	wire [4-1:0] node47121;
	wire [4-1:0] node47122;
	wire [4-1:0] node47123;
	wire [4-1:0] node47125;
	wire [4-1:0] node47126;
	wire [4-1:0] node47129;
	wire [4-1:0] node47132;
	wire [4-1:0] node47133;
	wire [4-1:0] node47134;
	wire [4-1:0] node47137;
	wire [4-1:0] node47140;
	wire [4-1:0] node47142;
	wire [4-1:0] node47145;
	wire [4-1:0] node47146;
	wire [4-1:0] node47148;
	wire [4-1:0] node47149;
	wire [4-1:0] node47152;
	wire [4-1:0] node47155;
	wire [4-1:0] node47156;
	wire [4-1:0] node47157;
	wire [4-1:0] node47162;
	wire [4-1:0] node47163;
	wire [4-1:0] node47164;
	wire [4-1:0] node47165;
	wire [4-1:0] node47167;
	wire [4-1:0] node47168;
	wire [4-1:0] node47172;
	wire [4-1:0] node47173;
	wire [4-1:0] node47174;
	wire [4-1:0] node47177;
	wire [4-1:0] node47180;
	wire [4-1:0] node47181;
	wire [4-1:0] node47184;
	wire [4-1:0] node47187;
	wire [4-1:0] node47188;
	wire [4-1:0] node47190;
	wire [4-1:0] node47191;
	wire [4-1:0] node47194;
	wire [4-1:0] node47197;
	wire [4-1:0] node47198;
	wire [4-1:0] node47201;
	wire [4-1:0] node47204;
	wire [4-1:0] node47205;
	wire [4-1:0] node47206;
	wire [4-1:0] node47207;
	wire [4-1:0] node47208;
	wire [4-1:0] node47212;
	wire [4-1:0] node47215;
	wire [4-1:0] node47216;
	wire [4-1:0] node47217;
	wire [4-1:0] node47220;
	wire [4-1:0] node47224;
	wire [4-1:0] node47225;
	wire [4-1:0] node47228;
	wire [4-1:0] node47230;
	wire [4-1:0] node47233;
	wire [4-1:0] node47234;
	wire [4-1:0] node47235;
	wire [4-1:0] node47236;
	wire [4-1:0] node47237;
	wire [4-1:0] node47239;
	wire [4-1:0] node47240;
	wire [4-1:0] node47243;
	wire [4-1:0] node47246;
	wire [4-1:0] node47247;
	wire [4-1:0] node47250;
	wire [4-1:0] node47253;
	wire [4-1:0] node47254;
	wire [4-1:0] node47256;
	wire [4-1:0] node47257;
	wire [4-1:0] node47260;
	wire [4-1:0] node47263;
	wire [4-1:0] node47264;
	wire [4-1:0] node47267;
	wire [4-1:0] node47270;
	wire [4-1:0] node47271;
	wire [4-1:0] node47272;
	wire [4-1:0] node47273;
	wire [4-1:0] node47275;
	wire [4-1:0] node47278;
	wire [4-1:0] node47279;
	wire [4-1:0] node47282;
	wire [4-1:0] node47285;
	wire [4-1:0] node47286;
	wire [4-1:0] node47287;
	wire [4-1:0] node47290;
	wire [4-1:0] node47294;
	wire [4-1:0] node47295;
	wire [4-1:0] node47296;
	wire [4-1:0] node47297;
	wire [4-1:0] node47300;
	wire [4-1:0] node47304;
	wire [4-1:0] node47305;
	wire [4-1:0] node47307;
	wire [4-1:0] node47310;
	wire [4-1:0] node47312;
	wire [4-1:0] node47315;
	wire [4-1:0] node47316;
	wire [4-1:0] node47317;
	wire [4-1:0] node47318;
	wire [4-1:0] node47319;
	wire [4-1:0] node47321;
	wire [4-1:0] node47324;
	wire [4-1:0] node47325;
	wire [4-1:0] node47329;
	wire [4-1:0] node47330;
	wire [4-1:0] node47331;
	wire [4-1:0] node47334;
	wire [4-1:0] node47337;
	wire [4-1:0] node47338;
	wire [4-1:0] node47341;
	wire [4-1:0] node47344;
	wire [4-1:0] node47345;
	wire [4-1:0] node47346;
	wire [4-1:0] node47347;
	wire [4-1:0] node47351;
	wire [4-1:0] node47352;
	wire [4-1:0] node47355;
	wire [4-1:0] node47358;
	wire [4-1:0] node47359;
	wire [4-1:0] node47360;
	wire [4-1:0] node47364;
	wire [4-1:0] node47367;
	wire [4-1:0] node47368;
	wire [4-1:0] node47369;
	wire [4-1:0] node47370;
	wire [4-1:0] node47372;
	wire [4-1:0] node47375;
	wire [4-1:0] node47376;
	wire [4-1:0] node47379;
	wire [4-1:0] node47382;
	wire [4-1:0] node47383;
	wire [4-1:0] node47386;
	wire [4-1:0] node47389;
	wire [4-1:0] node47390;
	wire [4-1:0] node47391;
	wire [4-1:0] node47394;
	wire [4-1:0] node47397;
	wire [4-1:0] node47398;
	wire [4-1:0] node47401;
	wire [4-1:0] node47404;
	wire [4-1:0] node47405;
	wire [4-1:0] node47406;
	wire [4-1:0] node47407;
	wire [4-1:0] node47408;
	wire [4-1:0] node47409;
	wire [4-1:0] node47410;
	wire [4-1:0] node47412;
	wire [4-1:0] node47415;
	wire [4-1:0] node47417;
	wire [4-1:0] node47418;
	wire [4-1:0] node47421;
	wire [4-1:0] node47424;
	wire [4-1:0] node47425;
	wire [4-1:0] node47426;
	wire [4-1:0] node47427;
	wire [4-1:0] node47430;
	wire [4-1:0] node47433;
	wire [4-1:0] node47434;
	wire [4-1:0] node47437;
	wire [4-1:0] node47440;
	wire [4-1:0] node47442;
	wire [4-1:0] node47443;
	wire [4-1:0] node47447;
	wire [4-1:0] node47448;
	wire [4-1:0] node47449;
	wire [4-1:0] node47450;
	wire [4-1:0] node47453;
	wire [4-1:0] node47455;
	wire [4-1:0] node47458;
	wire [4-1:0] node47459;
	wire [4-1:0] node47460;
	wire [4-1:0] node47463;
	wire [4-1:0] node47466;
	wire [4-1:0] node47467;
	wire [4-1:0] node47470;
	wire [4-1:0] node47473;
	wire [4-1:0] node47474;
	wire [4-1:0] node47475;
	wire [4-1:0] node47476;
	wire [4-1:0] node47480;
	wire [4-1:0] node47483;
	wire [4-1:0] node47485;
	wire [4-1:0] node47486;
	wire [4-1:0] node47490;
	wire [4-1:0] node47491;
	wire [4-1:0] node47492;
	wire [4-1:0] node47493;
	wire [4-1:0] node47494;
	wire [4-1:0] node47497;
	wire [4-1:0] node47500;
	wire [4-1:0] node47501;
	wire [4-1:0] node47503;
	wire [4-1:0] node47506;
	wire [4-1:0] node47507;
	wire [4-1:0] node47510;
	wire [4-1:0] node47513;
	wire [4-1:0] node47514;
	wire [4-1:0] node47515;
	wire [4-1:0] node47519;
	wire [4-1:0] node47520;
	wire [4-1:0] node47523;
	wire [4-1:0] node47524;
	wire [4-1:0] node47527;
	wire [4-1:0] node47530;
	wire [4-1:0] node47531;
	wire [4-1:0] node47532;
	wire [4-1:0] node47534;
	wire [4-1:0] node47535;
	wire [4-1:0] node47538;
	wire [4-1:0] node47541;
	wire [4-1:0] node47542;
	wire [4-1:0] node47545;
	wire [4-1:0] node47548;
	wire [4-1:0] node47549;
	wire [4-1:0] node47550;
	wire [4-1:0] node47554;
	wire [4-1:0] node47555;
	wire [4-1:0] node47559;
	wire [4-1:0] node47560;
	wire [4-1:0] node47561;
	wire [4-1:0] node47562;
	wire [4-1:0] node47563;
	wire [4-1:0] node47564;
	wire [4-1:0] node47567;
	wire [4-1:0] node47570;
	wire [4-1:0] node47571;
	wire [4-1:0] node47574;
	wire [4-1:0] node47577;
	wire [4-1:0] node47578;
	wire [4-1:0] node47579;
	wire [4-1:0] node47580;
	wire [4-1:0] node47584;
	wire [4-1:0] node47585;
	wire [4-1:0] node47588;
	wire [4-1:0] node47591;
	wire [4-1:0] node47593;
	wire [4-1:0] node47594;
	wire [4-1:0] node47597;
	wire [4-1:0] node47600;
	wire [4-1:0] node47601;
	wire [4-1:0] node47602;
	wire [4-1:0] node47603;
	wire [4-1:0] node47606;
	wire [4-1:0] node47609;
	wire [4-1:0] node47610;
	wire [4-1:0] node47612;
	wire [4-1:0] node47615;
	wire [4-1:0] node47617;
	wire [4-1:0] node47620;
	wire [4-1:0] node47621;
	wire [4-1:0] node47622;
	wire [4-1:0] node47623;
	wire [4-1:0] node47626;
	wire [4-1:0] node47629;
	wire [4-1:0] node47631;
	wire [4-1:0] node47634;
	wire [4-1:0] node47635;
	wire [4-1:0] node47639;
	wire [4-1:0] node47640;
	wire [4-1:0] node47641;
	wire [4-1:0] node47642;
	wire [4-1:0] node47643;
	wire [4-1:0] node47646;
	wire [4-1:0] node47649;
	wire [4-1:0] node47651;
	wire [4-1:0] node47653;
	wire [4-1:0] node47656;
	wire [4-1:0] node47657;
	wire [4-1:0] node47659;
	wire [4-1:0] node47660;
	wire [4-1:0] node47663;
	wire [4-1:0] node47666;
	wire [4-1:0] node47667;
	wire [4-1:0] node47670;
	wire [4-1:0] node47673;
	wire [4-1:0] node47674;
	wire [4-1:0] node47675;
	wire [4-1:0] node47676;
	wire [4-1:0] node47679;
	wire [4-1:0] node47683;
	wire [4-1:0] node47684;
	wire [4-1:0] node47685;
	wire [4-1:0] node47687;
	wire [4-1:0] node47691;
	wire [4-1:0] node47693;
	wire [4-1:0] node47694;
	wire [4-1:0] node47697;
	wire [4-1:0] node47700;
	wire [4-1:0] node47701;
	wire [4-1:0] node47702;
	wire [4-1:0] node47703;
	wire [4-1:0] node47704;
	wire [4-1:0] node47705;
	wire [4-1:0] node47706;
	wire [4-1:0] node47707;
	wire [4-1:0] node47710;
	wire [4-1:0] node47713;
	wire [4-1:0] node47714;
	wire [4-1:0] node47718;
	wire [4-1:0] node47719;
	wire [4-1:0] node47720;
	wire [4-1:0] node47724;
	wire [4-1:0] node47726;
	wire [4-1:0] node47729;
	wire [4-1:0] node47730;
	wire [4-1:0] node47731;
	wire [4-1:0] node47732;
	wire [4-1:0] node47735;
	wire [4-1:0] node47738;
	wire [4-1:0] node47739;
	wire [4-1:0] node47742;
	wire [4-1:0] node47745;
	wire [4-1:0] node47746;
	wire [4-1:0] node47748;
	wire [4-1:0] node47751;
	wire [4-1:0] node47752;
	wire [4-1:0] node47755;
	wire [4-1:0] node47758;
	wire [4-1:0] node47759;
	wire [4-1:0] node47760;
	wire [4-1:0] node47761;
	wire [4-1:0] node47762;
	wire [4-1:0] node47766;
	wire [4-1:0] node47769;
	wire [4-1:0] node47770;
	wire [4-1:0] node47771;
	wire [4-1:0] node47776;
	wire [4-1:0] node47777;
	wire [4-1:0] node47778;
	wire [4-1:0] node47779;
	wire [4-1:0] node47783;
	wire [4-1:0] node47784;
	wire [4-1:0] node47787;
	wire [4-1:0] node47790;
	wire [4-1:0] node47791;
	wire [4-1:0] node47792;
	wire [4-1:0] node47795;
	wire [4-1:0] node47798;
	wire [4-1:0] node47799;
	wire [4-1:0] node47803;
	wire [4-1:0] node47804;
	wire [4-1:0] node47805;
	wire [4-1:0] node47806;
	wire [4-1:0] node47809;
	wire [4-1:0] node47810;
	wire [4-1:0] node47811;
	wire [4-1:0] node47814;
	wire [4-1:0] node47817;
	wire [4-1:0] node47819;
	wire [4-1:0] node47822;
	wire [4-1:0] node47823;
	wire [4-1:0] node47824;
	wire [4-1:0] node47828;
	wire [4-1:0] node47829;
	wire [4-1:0] node47831;
	wire [4-1:0] node47834;
	wire [4-1:0] node47835;
	wire [4-1:0] node47838;
	wire [4-1:0] node47841;
	wire [4-1:0] node47842;
	wire [4-1:0] node47843;
	wire [4-1:0] node47845;
	wire [4-1:0] node47847;
	wire [4-1:0] node47850;
	wire [4-1:0] node47851;
	wire [4-1:0] node47852;
	wire [4-1:0] node47856;
	wire [4-1:0] node47859;
	wire [4-1:0] node47860;
	wire [4-1:0] node47861;
	wire [4-1:0] node47862;
	wire [4-1:0] node47866;
	wire [4-1:0] node47867;
	wire [4-1:0] node47870;
	wire [4-1:0] node47873;
	wire [4-1:0] node47874;
	wire [4-1:0] node47875;
	wire [4-1:0] node47878;
	wire [4-1:0] node47881;
	wire [4-1:0] node47883;
	wire [4-1:0] node47886;
	wire [4-1:0] node47887;
	wire [4-1:0] node47888;
	wire [4-1:0] node47889;
	wire [4-1:0] node47890;
	wire [4-1:0] node47891;
	wire [4-1:0] node47892;
	wire [4-1:0] node47897;
	wire [4-1:0] node47898;
	wire [4-1:0] node47901;
	wire [4-1:0] node47904;
	wire [4-1:0] node47905;
	wire [4-1:0] node47906;
	wire [4-1:0] node47909;
	wire [4-1:0] node47912;
	wire [4-1:0] node47914;
	wire [4-1:0] node47915;
	wire [4-1:0] node47918;
	wire [4-1:0] node47921;
	wire [4-1:0] node47922;
	wire [4-1:0] node47923;
	wire [4-1:0] node47924;
	wire [4-1:0] node47928;
	wire [4-1:0] node47929;
	wire [4-1:0] node47932;
	wire [4-1:0] node47935;
	wire [4-1:0] node47936;
	wire [4-1:0] node47937;
	wire [4-1:0] node47939;
	wire [4-1:0] node47942;
	wire [4-1:0] node47943;
	wire [4-1:0] node47946;
	wire [4-1:0] node47949;
	wire [4-1:0] node47951;
	wire [4-1:0] node47952;
	wire [4-1:0] node47955;
	wire [4-1:0] node47958;
	wire [4-1:0] node47959;
	wire [4-1:0] node47960;
	wire [4-1:0] node47961;
	wire [4-1:0] node47962;
	wire [4-1:0] node47965;
	wire [4-1:0] node47968;
	wire [4-1:0] node47969;
	wire [4-1:0] node47972;
	wire [4-1:0] node47975;
	wire [4-1:0] node47976;
	wire [4-1:0] node47977;
	wire [4-1:0] node47980;
	wire [4-1:0] node47983;
	wire [4-1:0] node47984;
	wire [4-1:0] node47987;
	wire [4-1:0] node47990;
	wire [4-1:0] node47991;
	wire [4-1:0] node47992;
	wire [4-1:0] node47993;
	wire [4-1:0] node47996;
	wire [4-1:0] node47999;
	wire [4-1:0] node48000;
	wire [4-1:0] node48003;
	wire [4-1:0] node48006;
	wire [4-1:0] node48007;
	wire [4-1:0] node48008;
	wire [4-1:0] node48009;
	wire [4-1:0] node48012;
	wire [4-1:0] node48016;
	wire [4-1:0] node48017;
	wire [4-1:0] node48018;
	wire [4-1:0] node48022;
	wire [4-1:0] node48023;
	wire [4-1:0] node48026;
	wire [4-1:0] node48029;
	wire [4-1:0] node48030;
	wire [4-1:0] node48031;
	wire [4-1:0] node48032;
	wire [4-1:0] node48033;
	wire [4-1:0] node48034;
	wire [4-1:0] node48035;
	wire [4-1:0] node48036;
	wire [4-1:0] node48037;
	wire [4-1:0] node48038;
	wire [4-1:0] node48039;
	wire [4-1:0] node48042;
	wire [4-1:0] node48045;
	wire [4-1:0] node48047;
	wire [4-1:0] node48050;
	wire [4-1:0] node48051;
	wire [4-1:0] node48052;
	wire [4-1:0] node48055;
	wire [4-1:0] node48059;
	wire [4-1:0] node48060;
	wire [4-1:0] node48061;
	wire [4-1:0] node48064;
	wire [4-1:0] node48067;
	wire [4-1:0] node48068;
	wire [4-1:0] node48069;
	wire [4-1:0] node48072;
	wire [4-1:0] node48075;
	wire [4-1:0] node48076;
	wire [4-1:0] node48079;
	wire [4-1:0] node48082;
	wire [4-1:0] node48083;
	wire [4-1:0] node48084;
	wire [4-1:0] node48085;
	wire [4-1:0] node48088;
	wire [4-1:0] node48091;
	wire [4-1:0] node48092;
	wire [4-1:0] node48095;
	wire [4-1:0] node48098;
	wire [4-1:0] node48099;
	wire [4-1:0] node48100;
	wire [4-1:0] node48103;
	wire [4-1:0] node48106;
	wire [4-1:0] node48107;
	wire [4-1:0] node48110;
	wire [4-1:0] node48113;
	wire [4-1:0] node48114;
	wire [4-1:0] node48115;
	wire [4-1:0] node48116;
	wire [4-1:0] node48118;
	wire [4-1:0] node48119;
	wire [4-1:0] node48122;
	wire [4-1:0] node48125;
	wire [4-1:0] node48126;
	wire [4-1:0] node48127;
	wire [4-1:0] node48130;
	wire [4-1:0] node48133;
	wire [4-1:0] node48134;
	wire [4-1:0] node48137;
	wire [4-1:0] node48140;
	wire [4-1:0] node48141;
	wire [4-1:0] node48142;
	wire [4-1:0] node48145;
	wire [4-1:0] node48148;
	wire [4-1:0] node48149;
	wire [4-1:0] node48153;
	wire [4-1:0] node48154;
	wire [4-1:0] node48156;
	wire [4-1:0] node48157;
	wire [4-1:0] node48158;
	wire [4-1:0] node48161;
	wire [4-1:0] node48164;
	wire [4-1:0] node48165;
	wire [4-1:0] node48168;
	wire [4-1:0] node48171;
	wire [4-1:0] node48172;
	wire [4-1:0] node48173;
	wire [4-1:0] node48174;
	wire [4-1:0] node48178;
	wire [4-1:0] node48180;
	wire [4-1:0] node48183;
	wire [4-1:0] node48184;
	wire [4-1:0] node48187;
	wire [4-1:0] node48190;
	wire [4-1:0] node48191;
	wire [4-1:0] node48192;
	wire [4-1:0] node48193;
	wire [4-1:0] node48194;
	wire [4-1:0] node48195;
	wire [4-1:0] node48196;
	wire [4-1:0] node48200;
	wire [4-1:0] node48201;
	wire [4-1:0] node48204;
	wire [4-1:0] node48207;
	wire [4-1:0] node48208;
	wire [4-1:0] node48209;
	wire [4-1:0] node48212;
	wire [4-1:0] node48215;
	wire [4-1:0] node48216;
	wire [4-1:0] node48219;
	wire [4-1:0] node48222;
	wire [4-1:0] node48223;
	wire [4-1:0] node48224;
	wire [4-1:0] node48227;
	wire [4-1:0] node48228;
	wire [4-1:0] node48232;
	wire [4-1:0] node48235;
	wire [4-1:0] node48236;
	wire [4-1:0] node48237;
	wire [4-1:0] node48238;
	wire [4-1:0] node48240;
	wire [4-1:0] node48243;
	wire [4-1:0] node48244;
	wire [4-1:0] node48248;
	wire [4-1:0] node48249;
	wire [4-1:0] node48250;
	wire [4-1:0] node48254;
	wire [4-1:0] node48255;
	wire [4-1:0] node48258;
	wire [4-1:0] node48261;
	wire [4-1:0] node48262;
	wire [4-1:0] node48265;
	wire [4-1:0] node48266;
	wire [4-1:0] node48268;
	wire [4-1:0] node48271;
	wire [4-1:0] node48272;
	wire [4-1:0] node48275;
	wire [4-1:0] node48278;
	wire [4-1:0] node48279;
	wire [4-1:0] node48280;
	wire [4-1:0] node48281;
	wire [4-1:0] node48282;
	wire [4-1:0] node48285;
	wire [4-1:0] node48288;
	wire [4-1:0] node48289;
	wire [4-1:0] node48291;
	wire [4-1:0] node48294;
	wire [4-1:0] node48295;
	wire [4-1:0] node48298;
	wire [4-1:0] node48301;
	wire [4-1:0] node48302;
	wire [4-1:0] node48303;
	wire [4-1:0] node48304;
	wire [4-1:0] node48307;
	wire [4-1:0] node48310;
	wire [4-1:0] node48311;
	wire [4-1:0] node48314;
	wire [4-1:0] node48317;
	wire [4-1:0] node48318;
	wire [4-1:0] node48322;
	wire [4-1:0] node48323;
	wire [4-1:0] node48324;
	wire [4-1:0] node48325;
	wire [4-1:0] node48328;
	wire [4-1:0] node48331;
	wire [4-1:0] node48332;
	wire [4-1:0] node48335;
	wire [4-1:0] node48338;
	wire [4-1:0] node48339;
	wire [4-1:0] node48340;
	wire [4-1:0] node48343;
	wire [4-1:0] node48346;
	wire [4-1:0] node48347;
	wire [4-1:0] node48350;
	wire [4-1:0] node48353;
	wire [4-1:0] node48354;
	wire [4-1:0] node48355;
	wire [4-1:0] node48356;
	wire [4-1:0] node48357;
	wire [4-1:0] node48358;
	wire [4-1:0] node48360;
	wire [4-1:0] node48361;
	wire [4-1:0] node48364;
	wire [4-1:0] node48367;
	wire [4-1:0] node48368;
	wire [4-1:0] node48369;
	wire [4-1:0] node48372;
	wire [4-1:0] node48376;
	wire [4-1:0] node48377;
	wire [4-1:0] node48378;
	wire [4-1:0] node48379;
	wire [4-1:0] node48383;
	wire [4-1:0] node48384;
	wire [4-1:0] node48387;
	wire [4-1:0] node48390;
	wire [4-1:0] node48391;
	wire [4-1:0] node48394;
	wire [4-1:0] node48395;
	wire [4-1:0] node48398;
	wire [4-1:0] node48401;
	wire [4-1:0] node48402;
	wire [4-1:0] node48403;
	wire [4-1:0] node48404;
	wire [4-1:0] node48407;
	wire [4-1:0] node48410;
	wire [4-1:0] node48411;
	wire [4-1:0] node48414;
	wire [4-1:0] node48417;
	wire [4-1:0] node48418;
	wire [4-1:0] node48419;
	wire [4-1:0] node48422;
	wire [4-1:0] node48425;
	wire [4-1:0] node48426;
	wire [4-1:0] node48430;
	wire [4-1:0] node48431;
	wire [4-1:0] node48432;
	wire [4-1:0] node48433;
	wire [4-1:0] node48434;
	wire [4-1:0] node48437;
	wire [4-1:0] node48440;
	wire [4-1:0] node48441;
	wire [4-1:0] node48442;
	wire [4-1:0] node48446;
	wire [4-1:0] node48447;
	wire [4-1:0] node48450;
	wire [4-1:0] node48453;
	wire [4-1:0] node48454;
	wire [4-1:0] node48455;
	wire [4-1:0] node48456;
	wire [4-1:0] node48460;
	wire [4-1:0] node48461;
	wire [4-1:0] node48465;
	wire [4-1:0] node48467;
	wire [4-1:0] node48470;
	wire [4-1:0] node48471;
	wire [4-1:0] node48472;
	wire [4-1:0] node48474;
	wire [4-1:0] node48475;
	wire [4-1:0] node48478;
	wire [4-1:0] node48481;
	wire [4-1:0] node48482;
	wire [4-1:0] node48484;
	wire [4-1:0] node48487;
	wire [4-1:0] node48488;
	wire [4-1:0] node48492;
	wire [4-1:0] node48493;
	wire [4-1:0] node48494;
	wire [4-1:0] node48497;
	wire [4-1:0] node48498;
	wire [4-1:0] node48501;
	wire [4-1:0] node48504;
	wire [4-1:0] node48505;
	wire [4-1:0] node48506;
	wire [4-1:0] node48510;
	wire [4-1:0] node48511;
	wire [4-1:0] node48514;
	wire [4-1:0] node48517;
	wire [4-1:0] node48518;
	wire [4-1:0] node48519;
	wire [4-1:0] node48520;
	wire [4-1:0] node48521;
	wire [4-1:0] node48523;
	wire [4-1:0] node48526;
	wire [4-1:0] node48527;
	wire [4-1:0] node48530;
	wire [4-1:0] node48533;
	wire [4-1:0] node48534;
	wire [4-1:0] node48535;
	wire [4-1:0] node48538;
	wire [4-1:0] node48541;
	wire [4-1:0] node48542;
	wire [4-1:0] node48543;
	wire [4-1:0] node48546;
	wire [4-1:0] node48549;
	wire [4-1:0] node48550;
	wire [4-1:0] node48553;
	wire [4-1:0] node48556;
	wire [4-1:0] node48557;
	wire [4-1:0] node48558;
	wire [4-1:0] node48559;
	wire [4-1:0] node48562;
	wire [4-1:0] node48565;
	wire [4-1:0] node48566;
	wire [4-1:0] node48569;
	wire [4-1:0] node48572;
	wire [4-1:0] node48573;
	wire [4-1:0] node48574;
	wire [4-1:0] node48575;
	wire [4-1:0] node48578;
	wire [4-1:0] node48581;
	wire [4-1:0] node48582;
	wire [4-1:0] node48586;
	wire [4-1:0] node48587;
	wire [4-1:0] node48590;
	wire [4-1:0] node48593;
	wire [4-1:0] node48594;
	wire [4-1:0] node48595;
	wire [4-1:0] node48596;
	wire [4-1:0] node48597;
	wire [4-1:0] node48599;
	wire [4-1:0] node48602;
	wire [4-1:0] node48603;
	wire [4-1:0] node48606;
	wire [4-1:0] node48609;
	wire [4-1:0] node48610;
	wire [4-1:0] node48611;
	wire [4-1:0] node48616;
	wire [4-1:0] node48617;
	wire [4-1:0] node48619;
	wire [4-1:0] node48620;
	wire [4-1:0] node48623;
	wire [4-1:0] node48626;
	wire [4-1:0] node48627;
	wire [4-1:0] node48631;
	wire [4-1:0] node48632;
	wire [4-1:0] node48633;
	wire [4-1:0] node48635;
	wire [4-1:0] node48636;
	wire [4-1:0] node48639;
	wire [4-1:0] node48642;
	wire [4-1:0] node48644;
	wire [4-1:0] node48647;
	wire [4-1:0] node48648;
	wire [4-1:0] node48651;
	wire [4-1:0] node48652;
	wire [4-1:0] node48655;
	wire [4-1:0] node48658;
	wire [4-1:0] node48659;
	wire [4-1:0] node48660;
	wire [4-1:0] node48661;
	wire [4-1:0] node48662;
	wire [4-1:0] node48663;
	wire [4-1:0] node48664;
	wire [4-1:0] node48667;
	wire [4-1:0] node48670;
	wire [4-1:0] node48671;
	wire [4-1:0] node48672;
	wire [4-1:0] node48676;
	wire [4-1:0] node48677;
	wire [4-1:0] node48680;
	wire [4-1:0] node48683;
	wire [4-1:0] node48684;
	wire [4-1:0] node48685;
	wire [4-1:0] node48686;
	wire [4-1:0] node48689;
	wire [4-1:0] node48692;
	wire [4-1:0] node48693;
	wire [4-1:0] node48696;
	wire [4-1:0] node48699;
	wire [4-1:0] node48700;
	wire [4-1:0] node48703;
	wire [4-1:0] node48706;
	wire [4-1:0] node48707;
	wire [4-1:0] node48708;
	wire [4-1:0] node48709;
	wire [4-1:0] node48711;
	wire [4-1:0] node48713;
	wire [4-1:0] node48716;
	wire [4-1:0] node48717;
	wire [4-1:0] node48719;
	wire [4-1:0] node48722;
	wire [4-1:0] node48723;
	wire [4-1:0] node48726;
	wire [4-1:0] node48729;
	wire [4-1:0] node48730;
	wire [4-1:0] node48733;
	wire [4-1:0] node48736;
	wire [4-1:0] node48737;
	wire [4-1:0] node48738;
	wire [4-1:0] node48739;
	wire [4-1:0] node48742;
	wire [4-1:0] node48745;
	wire [4-1:0] node48746;
	wire [4-1:0] node48749;
	wire [4-1:0] node48752;
	wire [4-1:0] node48753;
	wire [4-1:0] node48754;
	wire [4-1:0] node48758;
	wire [4-1:0] node48759;
	wire [4-1:0] node48762;
	wire [4-1:0] node48765;
	wire [4-1:0] node48766;
	wire [4-1:0] node48767;
	wire [4-1:0] node48768;
	wire [4-1:0] node48769;
	wire [4-1:0] node48770;
	wire [4-1:0] node48773;
	wire [4-1:0] node48776;
	wire [4-1:0] node48777;
	wire [4-1:0] node48780;
	wire [4-1:0] node48783;
	wire [4-1:0] node48784;
	wire [4-1:0] node48787;
	wire [4-1:0] node48790;
	wire [4-1:0] node48791;
	wire [4-1:0] node48792;
	wire [4-1:0] node48795;
	wire [4-1:0] node48798;
	wire [4-1:0] node48799;
	wire [4-1:0] node48801;
	wire [4-1:0] node48804;
	wire [4-1:0] node48805;
	wire [4-1:0] node48808;
	wire [4-1:0] node48811;
	wire [4-1:0] node48812;
	wire [4-1:0] node48813;
	wire [4-1:0] node48814;
	wire [4-1:0] node48817;
	wire [4-1:0] node48820;
	wire [4-1:0] node48821;
	wire [4-1:0] node48822;
	wire [4-1:0] node48825;
	wire [4-1:0] node48828;
	wire [4-1:0] node48829;
	wire [4-1:0] node48832;
	wire [4-1:0] node48835;
	wire [4-1:0] node48836;
	wire [4-1:0] node48837;
	wire [4-1:0] node48838;
	wire [4-1:0] node48841;
	wire [4-1:0] node48844;
	wire [4-1:0] node48845;
	wire [4-1:0] node48848;
	wire [4-1:0] node48851;
	wire [4-1:0] node48852;
	wire [4-1:0] node48853;
	wire [4-1:0] node48856;
	wire [4-1:0] node48859;
	wire [4-1:0] node48860;
	wire [4-1:0] node48861;
	wire [4-1:0] node48866;
	wire [4-1:0] node48867;
	wire [4-1:0] node48868;
	wire [4-1:0] node48869;
	wire [4-1:0] node48870;
	wire [4-1:0] node48872;
	wire [4-1:0] node48873;
	wire [4-1:0] node48876;
	wire [4-1:0] node48879;
	wire [4-1:0] node48880;
	wire [4-1:0] node48883;
	wire [4-1:0] node48886;
	wire [4-1:0] node48887;
	wire [4-1:0] node48888;
	wire [4-1:0] node48889;
	wire [4-1:0] node48891;
	wire [4-1:0] node48895;
	wire [4-1:0] node48896;
	wire [4-1:0] node48899;
	wire [4-1:0] node48902;
	wire [4-1:0] node48903;
	wire [4-1:0] node48906;
	wire [4-1:0] node48909;
	wire [4-1:0] node48910;
	wire [4-1:0] node48911;
	wire [4-1:0] node48912;
	wire [4-1:0] node48915;
	wire [4-1:0] node48918;
	wire [4-1:0] node48919;
	wire [4-1:0] node48920;
	wire [4-1:0] node48923;
	wire [4-1:0] node48926;
	wire [4-1:0] node48927;
	wire [4-1:0] node48931;
	wire [4-1:0] node48932;
	wire [4-1:0] node48933;
	wire [4-1:0] node48934;
	wire [4-1:0] node48935;
	wire [4-1:0] node48938;
	wire [4-1:0] node48942;
	wire [4-1:0] node48944;
	wire [4-1:0] node48945;
	wire [4-1:0] node48948;
	wire [4-1:0] node48951;
	wire [4-1:0] node48952;
	wire [4-1:0] node48953;
	wire [4-1:0] node48957;
	wire [4-1:0] node48958;
	wire [4-1:0] node48959;
	wire [4-1:0] node48962;
	wire [4-1:0] node48965;
	wire [4-1:0] node48967;
	wire [4-1:0] node48970;
	wire [4-1:0] node48971;
	wire [4-1:0] node48972;
	wire [4-1:0] node48973;
	wire [4-1:0] node48974;
	wire [4-1:0] node48975;
	wire [4-1:0] node48978;
	wire [4-1:0] node48981;
	wire [4-1:0] node48982;
	wire [4-1:0] node48986;
	wire [4-1:0] node48987;
	wire [4-1:0] node48990;
	wire [4-1:0] node48993;
	wire [4-1:0] node48994;
	wire [4-1:0] node48995;
	wire [4-1:0] node48998;
	wire [4-1:0] node49001;
	wire [4-1:0] node49002;
	wire [4-1:0] node49003;
	wire [4-1:0] node49007;
	wire [4-1:0] node49008;
	wire [4-1:0] node49012;
	wire [4-1:0] node49013;
	wire [4-1:0] node49014;
	wire [4-1:0] node49015;
	wire [4-1:0] node49018;
	wire [4-1:0] node49021;
	wire [4-1:0] node49022;
	wire [4-1:0] node49024;
	wire [4-1:0] node49027;
	wire [4-1:0] node49028;
	wire [4-1:0] node49031;
	wire [4-1:0] node49034;
	wire [4-1:0] node49035;
	wire [4-1:0] node49036;
	wire [4-1:0] node49039;
	wire [4-1:0] node49042;
	wire [4-1:0] node49043;
	wire [4-1:0] node49044;
	wire [4-1:0] node49047;
	wire [4-1:0] node49050;
	wire [4-1:0] node49052;
	wire [4-1:0] node49053;
	wire [4-1:0] node49056;
	wire [4-1:0] node49059;
	wire [4-1:0] node49060;
	wire [4-1:0] node49061;
	wire [4-1:0] node49062;
	wire [4-1:0] node49063;
	wire [4-1:0] node49064;
	wire [4-1:0] node49065;
	wire [4-1:0] node49066;
	wire [4-1:0] node49067;
	wire [4-1:0] node49071;
	wire [4-1:0] node49072;
	wire [4-1:0] node49075;
	wire [4-1:0] node49078;
	wire [4-1:0] node49079;
	wire [4-1:0] node49080;
	wire [4-1:0] node49083;
	wire [4-1:0] node49086;
	wire [4-1:0] node49088;
	wire [4-1:0] node49091;
	wire [4-1:0] node49092;
	wire [4-1:0] node49093;
	wire [4-1:0] node49094;
	wire [4-1:0] node49095;
	wire [4-1:0] node49099;
	wire [4-1:0] node49102;
	wire [4-1:0] node49103;
	wire [4-1:0] node49104;
	wire [4-1:0] node49108;
	wire [4-1:0] node49111;
	wire [4-1:0] node49112;
	wire [4-1:0] node49113;
	wire [4-1:0] node49114;
	wire [4-1:0] node49118;
	wire [4-1:0] node49121;
	wire [4-1:0] node49122;
	wire [4-1:0] node49125;
	wire [4-1:0] node49126;
	wire [4-1:0] node49130;
	wire [4-1:0] node49131;
	wire [4-1:0] node49132;
	wire [4-1:0] node49133;
	wire [4-1:0] node49134;
	wire [4-1:0] node49136;
	wire [4-1:0] node49139;
	wire [4-1:0] node49140;
	wire [4-1:0] node49143;
	wire [4-1:0] node49147;
	wire [4-1:0] node49148;
	wire [4-1:0] node49151;
	wire [4-1:0] node49154;
	wire [4-1:0] node49155;
	wire [4-1:0] node49156;
	wire [4-1:0] node49159;
	wire [4-1:0] node49162;
	wire [4-1:0] node49163;
	wire [4-1:0] node49164;
	wire [4-1:0] node49167;
	wire [4-1:0] node49170;
	wire [4-1:0] node49171;
	wire [4-1:0] node49174;
	wire [4-1:0] node49177;
	wire [4-1:0] node49178;
	wire [4-1:0] node49179;
	wire [4-1:0] node49180;
	wire [4-1:0] node49181;
	wire [4-1:0] node49182;
	wire [4-1:0] node49185;
	wire [4-1:0] node49188;
	wire [4-1:0] node49189;
	wire [4-1:0] node49192;
	wire [4-1:0] node49195;
	wire [4-1:0] node49196;
	wire [4-1:0] node49198;
	wire [4-1:0] node49201;
	wire [4-1:0] node49202;
	wire [4-1:0] node49205;
	wire [4-1:0] node49208;
	wire [4-1:0] node49209;
	wire [4-1:0] node49210;
	wire [4-1:0] node49212;
	wire [4-1:0] node49215;
	wire [4-1:0] node49216;
	wire [4-1:0] node49219;
	wire [4-1:0] node49222;
	wire [4-1:0] node49223;
	wire [4-1:0] node49224;
	wire [4-1:0] node49227;
	wire [4-1:0] node49230;
	wire [4-1:0] node49231;
	wire [4-1:0] node49234;
	wire [4-1:0] node49237;
	wire [4-1:0] node49238;
	wire [4-1:0] node49239;
	wire [4-1:0] node49240;
	wire [4-1:0] node49241;
	wire [4-1:0] node49242;
	wire [4-1:0] node49246;
	wire [4-1:0] node49247;
	wire [4-1:0] node49251;
	wire [4-1:0] node49252;
	wire [4-1:0] node49255;
	wire [4-1:0] node49258;
	wire [4-1:0] node49259;
	wire [4-1:0] node49260;
	wire [4-1:0] node49261;
	wire [4-1:0] node49265;
	wire [4-1:0] node49266;
	wire [4-1:0] node49270;
	wire [4-1:0] node49271;
	wire [4-1:0] node49274;
	wire [4-1:0] node49277;
	wire [4-1:0] node49278;
	wire [4-1:0] node49279;
	wire [4-1:0] node49282;
	wire [4-1:0] node49285;
	wire [4-1:0] node49286;
	wire [4-1:0] node49289;
	wire [4-1:0] node49292;
	wire [4-1:0] node49293;
	wire [4-1:0] node49294;
	wire [4-1:0] node49295;
	wire [4-1:0] node49296;
	wire [4-1:0] node49297;
	wire [4-1:0] node49298;
	wire [4-1:0] node49302;
	wire [4-1:0] node49305;
	wire [4-1:0] node49306;
	wire [4-1:0] node49307;
	wire [4-1:0] node49311;
	wire [4-1:0] node49314;
	wire [4-1:0] node49315;
	wire [4-1:0] node49316;
	wire [4-1:0] node49317;
	wire [4-1:0] node49320;
	wire [4-1:0] node49323;
	wire [4-1:0] node49324;
	wire [4-1:0] node49327;
	wire [4-1:0] node49330;
	wire [4-1:0] node49331;
	wire [4-1:0] node49332;
	wire [4-1:0] node49334;
	wire [4-1:0] node49337;
	wire [4-1:0] node49338;
	wire [4-1:0] node49342;
	wire [4-1:0] node49343;
	wire [4-1:0] node49344;
	wire [4-1:0] node49348;
	wire [4-1:0] node49351;
	wire [4-1:0] node49352;
	wire [4-1:0] node49353;
	wire [4-1:0] node49354;
	wire [4-1:0] node49356;
	wire [4-1:0] node49359;
	wire [4-1:0] node49360;
	wire [4-1:0] node49363;
	wire [4-1:0] node49366;
	wire [4-1:0] node49367;
	wire [4-1:0] node49368;
	wire [4-1:0] node49371;
	wire [4-1:0] node49374;
	wire [4-1:0] node49375;
	wire [4-1:0] node49378;
	wire [4-1:0] node49381;
	wire [4-1:0] node49382;
	wire [4-1:0] node49383;
	wire [4-1:0] node49384;
	wire [4-1:0] node49388;
	wire [4-1:0] node49391;
	wire [4-1:0] node49392;
	wire [4-1:0] node49393;
	wire [4-1:0] node49394;
	wire [4-1:0] node49399;
	wire [4-1:0] node49400;
	wire [4-1:0] node49404;
	wire [4-1:0] node49405;
	wire [4-1:0] node49406;
	wire [4-1:0] node49407;
	wire [4-1:0] node49408;
	wire [4-1:0] node49409;
	wire [4-1:0] node49410;
	wire [4-1:0] node49414;
	wire [4-1:0] node49418;
	wire [4-1:0] node49419;
	wire [4-1:0] node49420;
	wire [4-1:0] node49424;
	wire [4-1:0] node49427;
	wire [4-1:0] node49428;
	wire [4-1:0] node49429;
	wire [4-1:0] node49430;
	wire [4-1:0] node49431;
	wire [4-1:0] node49434;
	wire [4-1:0] node49438;
	wire [4-1:0] node49439;
	wire [4-1:0] node49442;
	wire [4-1:0] node49445;
	wire [4-1:0] node49446;
	wire [4-1:0] node49447;
	wire [4-1:0] node49451;
	wire [4-1:0] node49454;
	wire [4-1:0] node49455;
	wire [4-1:0] node49456;
	wire [4-1:0] node49457;
	wire [4-1:0] node49458;
	wire [4-1:0] node49461;
	wire [4-1:0] node49464;
	wire [4-1:0] node49465;
	wire [4-1:0] node49468;
	wire [4-1:0] node49471;
	wire [4-1:0] node49472;
	wire [4-1:0] node49473;
	wire [4-1:0] node49476;
	wire [4-1:0] node49479;
	wire [4-1:0] node49480;
	wire [4-1:0] node49483;
	wire [4-1:0] node49486;
	wire [4-1:0] node49487;
	wire [4-1:0] node49488;
	wire [4-1:0] node49489;
	wire [4-1:0] node49492;
	wire [4-1:0] node49495;
	wire [4-1:0] node49497;
	wire [4-1:0] node49500;
	wire [4-1:0] node49501;
	wire [4-1:0] node49502;
	wire [4-1:0] node49506;
	wire [4-1:0] node49507;
	wire [4-1:0] node49511;
	wire [4-1:0] node49512;
	wire [4-1:0] node49513;
	wire [4-1:0] node49514;
	wire [4-1:0] node49515;
	wire [4-1:0] node49516;
	wire [4-1:0] node49517;
	wire [4-1:0] node49518;
	wire [4-1:0] node49522;
	wire [4-1:0] node49523;
	wire [4-1:0] node49526;
	wire [4-1:0] node49527;
	wire [4-1:0] node49531;
	wire [4-1:0] node49532;
	wire [4-1:0] node49535;
	wire [4-1:0] node49538;
	wire [4-1:0] node49539;
	wire [4-1:0] node49540;
	wire [4-1:0] node49541;
	wire [4-1:0] node49545;
	wire [4-1:0] node49548;
	wire [4-1:0] node49549;
	wire [4-1:0] node49550;
	wire [4-1:0] node49554;
	wire [4-1:0] node49557;
	wire [4-1:0] node49558;
	wire [4-1:0] node49559;
	wire [4-1:0] node49560;
	wire [4-1:0] node49561;
	wire [4-1:0] node49564;
	wire [4-1:0] node49567;
	wire [4-1:0] node49568;
	wire [4-1:0] node49571;
	wire [4-1:0] node49574;
	wire [4-1:0] node49575;
	wire [4-1:0] node49576;
	wire [4-1:0] node49579;
	wire [4-1:0] node49583;
	wire [4-1:0] node49584;
	wire [4-1:0] node49585;
	wire [4-1:0] node49588;
	wire [4-1:0] node49591;
	wire [4-1:0] node49592;
	wire [4-1:0] node49594;
	wire [4-1:0] node49597;
	wire [4-1:0] node49598;
	wire [4-1:0] node49601;
	wire [4-1:0] node49604;
	wire [4-1:0] node49605;
	wire [4-1:0] node49606;
	wire [4-1:0] node49607;
	wire [4-1:0] node49608;
	wire [4-1:0] node49612;
	wire [4-1:0] node49615;
	wire [4-1:0] node49616;
	wire [4-1:0] node49617;
	wire [4-1:0] node49621;
	wire [4-1:0] node49624;
	wire [4-1:0] node49625;
	wire [4-1:0] node49626;
	wire [4-1:0] node49627;
	wire [4-1:0] node49631;
	wire [4-1:0] node49634;
	wire [4-1:0] node49635;
	wire [4-1:0] node49636;
	wire [4-1:0] node49640;
	wire [4-1:0] node49643;
	wire [4-1:0] node49644;
	wire [4-1:0] node49645;
	wire [4-1:0] node49646;
	wire [4-1:0] node49647;
	wire [4-1:0] node49649;
	wire [4-1:0] node49650;
	wire [4-1:0] node49653;
	wire [4-1:0] node49656;
	wire [4-1:0] node49657;
	wire [4-1:0] node49658;
	wire [4-1:0] node49659;
	wire [4-1:0] node49662;
	wire [4-1:0] node49665;
	wire [4-1:0] node49666;
	wire [4-1:0] node49669;
	wire [4-1:0] node49672;
	wire [4-1:0] node49673;
	wire [4-1:0] node49676;
	wire [4-1:0] node49679;
	wire [4-1:0] node49680;
	wire [4-1:0] node49681;
	wire [4-1:0] node49684;
	wire [4-1:0] node49687;
	wire [4-1:0] node49688;
	wire [4-1:0] node49689;
	wire [4-1:0] node49692;
	wire [4-1:0] node49695;
	wire [4-1:0] node49696;
	wire [4-1:0] node49699;
	wire [4-1:0] node49702;
	wire [4-1:0] node49703;
	wire [4-1:0] node49704;
	wire [4-1:0] node49705;
	wire [4-1:0] node49706;
	wire [4-1:0] node49708;
	wire [4-1:0] node49711;
	wire [4-1:0] node49712;
	wire [4-1:0] node49716;
	wire [4-1:0] node49717;
	wire [4-1:0] node49721;
	wire [4-1:0] node49722;
	wire [4-1:0] node49723;
	wire [4-1:0] node49724;
	wire [4-1:0] node49727;
	wire [4-1:0] node49731;
	wire [4-1:0] node49732;
	wire [4-1:0] node49733;
	wire [4-1:0] node49737;
	wire [4-1:0] node49738;
	wire [4-1:0] node49741;
	wire [4-1:0] node49744;
	wire [4-1:0] node49745;
	wire [4-1:0] node49746;
	wire [4-1:0] node49748;
	wire [4-1:0] node49749;
	wire [4-1:0] node49752;
	wire [4-1:0] node49755;
	wire [4-1:0] node49756;
	wire [4-1:0] node49760;
	wire [4-1:0] node49761;
	wire [4-1:0] node49762;
	wire [4-1:0] node49764;
	wire [4-1:0] node49767;
	wire [4-1:0] node49769;
	wire [4-1:0] node49772;
	wire [4-1:0] node49773;
	wire [4-1:0] node49777;
	wire [4-1:0] node49778;
	wire [4-1:0] node49779;
	wire [4-1:0] node49780;
	wire [4-1:0] node49781;
	wire [4-1:0] node49782;
	wire [4-1:0] node49784;
	wire [4-1:0] node49787;
	wire [4-1:0] node49788;
	wire [4-1:0] node49792;
	wire [4-1:0] node49793;
	wire [4-1:0] node49794;
	wire [4-1:0] node49797;
	wire [4-1:0] node49800;
	wire [4-1:0] node49801;
	wire [4-1:0] node49804;
	wire [4-1:0] node49807;
	wire [4-1:0] node49808;
	wire [4-1:0] node49809;
	wire [4-1:0] node49812;
	wire [4-1:0] node49815;
	wire [4-1:0] node49816;
	wire [4-1:0] node49819;
	wire [4-1:0] node49822;
	wire [4-1:0] node49823;
	wire [4-1:0] node49826;
	wire [4-1:0] node49829;
	wire [4-1:0] node49830;
	wire [4-1:0] node49831;
	wire [4-1:0] node49832;
	wire [4-1:0] node49835;
	wire [4-1:0] node49838;
	wire [4-1:0] node49839;
	wire [4-1:0] node49842;
	wire [4-1:0] node49845;
	wire [4-1:0] node49846;
	wire [4-1:0] node49849;
	wire [4-1:0] node49852;
	wire [4-1:0] node49853;
	wire [4-1:0] node49854;
	wire [4-1:0] node49855;
	wire [4-1:0] node49856;
	wire [4-1:0] node49857;
	wire [4-1:0] node49858;
	wire [4-1:0] node49859;
	wire [4-1:0] node49860;
	wire [4-1:0] node49861;
	wire [4-1:0] node49862;
	wire [4-1:0] node49863;
	wire [4-1:0] node49864;
	wire [4-1:0] node49865;
	wire [4-1:0] node49868;
	wire [4-1:0] node49871;
	wire [4-1:0] node49872;
	wire [4-1:0] node49875;
	wire [4-1:0] node49878;
	wire [4-1:0] node49879;
	wire [4-1:0] node49881;
	wire [4-1:0] node49884;
	wire [4-1:0] node49886;
	wire [4-1:0] node49889;
	wire [4-1:0] node49890;
	wire [4-1:0] node49891;
	wire [4-1:0] node49892;
	wire [4-1:0] node49895;
	wire [4-1:0] node49898;
	wire [4-1:0] node49899;
	wire [4-1:0] node49902;
	wire [4-1:0] node49905;
	wire [4-1:0] node49906;
	wire [4-1:0] node49907;
	wire [4-1:0] node49911;
	wire [4-1:0] node49914;
	wire [4-1:0] node49915;
	wire [4-1:0] node49916;
	wire [4-1:0] node49917;
	wire [4-1:0] node49920;
	wire [4-1:0] node49923;
	wire [4-1:0] node49924;
	wire [4-1:0] node49926;
	wire [4-1:0] node49929;
	wire [4-1:0] node49930;
	wire [4-1:0] node49933;
	wire [4-1:0] node49936;
	wire [4-1:0] node49937;
	wire [4-1:0] node49938;
	wire [4-1:0] node49939;
	wire [4-1:0] node49943;
	wire [4-1:0] node49944;
	wire [4-1:0] node49947;
	wire [4-1:0] node49950;
	wire [4-1:0] node49951;
	wire [4-1:0] node49952;
	wire [4-1:0] node49956;
	wire [4-1:0] node49957;
	wire [4-1:0] node49960;
	wire [4-1:0] node49963;
	wire [4-1:0] node49964;
	wire [4-1:0] node49965;
	wire [4-1:0] node49966;
	wire [4-1:0] node49967;
	wire [4-1:0] node49968;
	wire [4-1:0] node49972;
	wire [4-1:0] node49973;
	wire [4-1:0] node49976;
	wire [4-1:0] node49979;
	wire [4-1:0] node49980;
	wire [4-1:0] node49981;
	wire [4-1:0] node49985;
	wire [4-1:0] node49987;
	wire [4-1:0] node49990;
	wire [4-1:0] node49991;
	wire [4-1:0] node49992;
	wire [4-1:0] node49993;
	wire [4-1:0] node49997;
	wire [4-1:0] node49998;
	wire [4-1:0] node50001;
	wire [4-1:0] node50004;
	wire [4-1:0] node50005;
	wire [4-1:0] node50007;
	wire [4-1:0] node50010;
	wire [4-1:0] node50011;
	wire [4-1:0] node50014;
	wire [4-1:0] node50017;
	wire [4-1:0] node50018;
	wire [4-1:0] node50019;
	wire [4-1:0] node50021;
	wire [4-1:0] node50023;
	wire [4-1:0] node50026;
	wire [4-1:0] node50027;
	wire [4-1:0] node50030;
	wire [4-1:0] node50033;
	wire [4-1:0] node50034;
	wire [4-1:0] node50035;
	wire [4-1:0] node50037;
	wire [4-1:0] node50040;
	wire [4-1:0] node50042;
	wire [4-1:0] node50045;
	wire [4-1:0] node50046;
	wire [4-1:0] node50047;
	wire [4-1:0] node50052;
	wire [4-1:0] node50053;
	wire [4-1:0] node50054;
	wire [4-1:0] node50055;
	wire [4-1:0] node50056;
	wire [4-1:0] node50057;
	wire [4-1:0] node50059;
	wire [4-1:0] node50062;
	wire [4-1:0] node50064;
	wire [4-1:0] node50067;
	wire [4-1:0] node50068;
	wire [4-1:0] node50069;
	wire [4-1:0] node50074;
	wire [4-1:0] node50075;
	wire [4-1:0] node50077;
	wire [4-1:0] node50078;
	wire [4-1:0] node50081;
	wire [4-1:0] node50084;
	wire [4-1:0] node50085;
	wire [4-1:0] node50088;
	wire [4-1:0] node50091;
	wire [4-1:0] node50092;
	wire [4-1:0] node50093;
	wire [4-1:0] node50095;
	wire [4-1:0] node50097;
	wire [4-1:0] node50100;
	wire [4-1:0] node50101;
	wire [4-1:0] node50102;
	wire [4-1:0] node50105;
	wire [4-1:0] node50109;
	wire [4-1:0] node50110;
	wire [4-1:0] node50112;
	wire [4-1:0] node50113;
	wire [4-1:0] node50116;
	wire [4-1:0] node50119;
	wire [4-1:0] node50121;
	wire [4-1:0] node50124;
	wire [4-1:0] node50125;
	wire [4-1:0] node50126;
	wire [4-1:0] node50127;
	wire [4-1:0] node50128;
	wire [4-1:0] node50131;
	wire [4-1:0] node50135;
	wire [4-1:0] node50136;
	wire [4-1:0] node50137;
	wire [4-1:0] node50140;
	wire [4-1:0] node50143;
	wire [4-1:0] node50144;
	wire [4-1:0] node50147;
	wire [4-1:0] node50150;
	wire [4-1:0] node50151;
	wire [4-1:0] node50152;
	wire [4-1:0] node50153;
	wire [4-1:0] node50156;
	wire [4-1:0] node50159;
	wire [4-1:0] node50160;
	wire [4-1:0] node50163;
	wire [4-1:0] node50166;
	wire [4-1:0] node50167;
	wire [4-1:0] node50169;
	wire [4-1:0] node50172;
	wire [4-1:0] node50174;
	wire [4-1:0] node50175;
	wire [4-1:0] node50178;
	wire [4-1:0] node50181;
	wire [4-1:0] node50182;
	wire [4-1:0] node50183;
	wire [4-1:0] node50184;
	wire [4-1:0] node50185;
	wire [4-1:0] node50186;
	wire [4-1:0] node50187;
	wire [4-1:0] node50190;
	wire [4-1:0] node50192;
	wire [4-1:0] node50195;
	wire [4-1:0] node50196;
	wire [4-1:0] node50199;
	wire [4-1:0] node50202;
	wire [4-1:0] node50204;
	wire [4-1:0] node50205;
	wire [4-1:0] node50206;
	wire [4-1:0] node50210;
	wire [4-1:0] node50213;
	wire [4-1:0] node50214;
	wire [4-1:0] node50215;
	wire [4-1:0] node50216;
	wire [4-1:0] node50217;
	wire [4-1:0] node50221;
	wire [4-1:0] node50224;
	wire [4-1:0] node50225;
	wire [4-1:0] node50226;
	wire [4-1:0] node50229;
	wire [4-1:0] node50232;
	wire [4-1:0] node50233;
	wire [4-1:0] node50237;
	wire [4-1:0] node50238;
	wire [4-1:0] node50239;
	wire [4-1:0] node50240;
	wire [4-1:0] node50243;
	wire [4-1:0] node50246;
	wire [4-1:0] node50247;
	wire [4-1:0] node50250;
	wire [4-1:0] node50253;
	wire [4-1:0] node50254;
	wire [4-1:0] node50255;
	wire [4-1:0] node50259;
	wire [4-1:0] node50260;
	wire [4-1:0] node50263;
	wire [4-1:0] node50266;
	wire [4-1:0] node50267;
	wire [4-1:0] node50268;
	wire [4-1:0] node50269;
	wire [4-1:0] node50271;
	wire [4-1:0] node50274;
	wire [4-1:0] node50275;
	wire [4-1:0] node50278;
	wire [4-1:0] node50281;
	wire [4-1:0] node50282;
	wire [4-1:0] node50283;
	wire [4-1:0] node50285;
	wire [4-1:0] node50288;
	wire [4-1:0] node50290;
	wire [4-1:0] node50293;
	wire [4-1:0] node50294;
	wire [4-1:0] node50295;
	wire [4-1:0] node50298;
	wire [4-1:0] node50301;
	wire [4-1:0] node50303;
	wire [4-1:0] node50306;
	wire [4-1:0] node50307;
	wire [4-1:0] node50308;
	wire [4-1:0] node50310;
	wire [4-1:0] node50312;
	wire [4-1:0] node50315;
	wire [4-1:0] node50316;
	wire [4-1:0] node50318;
	wire [4-1:0] node50321;
	wire [4-1:0] node50324;
	wire [4-1:0] node50325;
	wire [4-1:0] node50326;
	wire [4-1:0] node50327;
	wire [4-1:0] node50330;
	wire [4-1:0] node50333;
	wire [4-1:0] node50335;
	wire [4-1:0] node50338;
	wire [4-1:0] node50339;
	wire [4-1:0] node50340;
	wire [4-1:0] node50343;
	wire [4-1:0] node50346;
	wire [4-1:0] node50347;
	wire [4-1:0] node50350;
	wire [4-1:0] node50353;
	wire [4-1:0] node50354;
	wire [4-1:0] node50355;
	wire [4-1:0] node50356;
	wire [4-1:0] node50357;
	wire [4-1:0] node50358;
	wire [4-1:0] node50359;
	wire [4-1:0] node50362;
	wire [4-1:0] node50366;
	wire [4-1:0] node50367;
	wire [4-1:0] node50368;
	wire [4-1:0] node50371;
	wire [4-1:0] node50375;
	wire [4-1:0] node50376;
	wire [4-1:0] node50377;
	wire [4-1:0] node50378;
	wire [4-1:0] node50383;
	wire [4-1:0] node50384;
	wire [4-1:0] node50385;
	wire [4-1:0] node50388;
	wire [4-1:0] node50391;
	wire [4-1:0] node50392;
	wire [4-1:0] node50395;
	wire [4-1:0] node50398;
	wire [4-1:0] node50399;
	wire [4-1:0] node50400;
	wire [4-1:0] node50401;
	wire [4-1:0] node50402;
	wire [4-1:0] node50405;
	wire [4-1:0] node50408;
	wire [4-1:0] node50409;
	wire [4-1:0] node50412;
	wire [4-1:0] node50415;
	wire [4-1:0] node50416;
	wire [4-1:0] node50417;
	wire [4-1:0] node50420;
	wire [4-1:0] node50423;
	wire [4-1:0] node50425;
	wire [4-1:0] node50428;
	wire [4-1:0] node50429;
	wire [4-1:0] node50430;
	wire [4-1:0] node50431;
	wire [4-1:0] node50434;
	wire [4-1:0] node50437;
	wire [4-1:0] node50438;
	wire [4-1:0] node50442;
	wire [4-1:0] node50443;
	wire [4-1:0] node50444;
	wire [4-1:0] node50449;
	wire [4-1:0] node50450;
	wire [4-1:0] node50451;
	wire [4-1:0] node50452;
	wire [4-1:0] node50453;
	wire [4-1:0] node50456;
	wire [4-1:0] node50459;
	wire [4-1:0] node50460;
	wire [4-1:0] node50463;
	wire [4-1:0] node50465;
	wire [4-1:0] node50468;
	wire [4-1:0] node50469;
	wire [4-1:0] node50470;
	wire [4-1:0] node50474;
	wire [4-1:0] node50475;
	wire [4-1:0] node50476;
	wire [4-1:0] node50479;
	wire [4-1:0] node50482;
	wire [4-1:0] node50483;
	wire [4-1:0] node50486;
	wire [4-1:0] node50489;
	wire [4-1:0] node50490;
	wire [4-1:0] node50491;
	wire [4-1:0] node50492;
	wire [4-1:0] node50493;
	wire [4-1:0] node50496;
	wire [4-1:0] node50500;
	wire [4-1:0] node50501;
	wire [4-1:0] node50503;
	wire [4-1:0] node50506;
	wire [4-1:0] node50507;
	wire [4-1:0] node50510;
	wire [4-1:0] node50513;
	wire [4-1:0] node50514;
	wire [4-1:0] node50515;
	wire [4-1:0] node50518;
	wire [4-1:0] node50520;
	wire [4-1:0] node50523;
	wire [4-1:0] node50525;
	wire [4-1:0] node50527;
	wire [4-1:0] node50530;
	wire [4-1:0] node50531;
	wire [4-1:0] node50532;
	wire [4-1:0] node50533;
	wire [4-1:0] node50534;
	wire [4-1:0] node50535;
	wire [4-1:0] node50536;
	wire [4-1:0] node50537;
	wire [4-1:0] node50538;
	wire [4-1:0] node50542;
	wire [4-1:0] node50543;
	wire [4-1:0] node50546;
	wire [4-1:0] node50549;
	wire [4-1:0] node50551;
	wire [4-1:0] node50552;
	wire [4-1:0] node50556;
	wire [4-1:0] node50557;
	wire [4-1:0] node50558;
	wire [4-1:0] node50559;
	wire [4-1:0] node50562;
	wire [4-1:0] node50565;
	wire [4-1:0] node50567;
	wire [4-1:0] node50570;
	wire [4-1:0] node50571;
	wire [4-1:0] node50572;
	wire [4-1:0] node50575;
	wire [4-1:0] node50578;
	wire [4-1:0] node50579;
	wire [4-1:0] node50583;
	wire [4-1:0] node50584;
	wire [4-1:0] node50585;
	wire [4-1:0] node50587;
	wire [4-1:0] node50588;
	wire [4-1:0] node50591;
	wire [4-1:0] node50594;
	wire [4-1:0] node50595;
	wire [4-1:0] node50596;
	wire [4-1:0] node50599;
	wire [4-1:0] node50602;
	wire [4-1:0] node50604;
	wire [4-1:0] node50607;
	wire [4-1:0] node50608;
	wire [4-1:0] node50610;
	wire [4-1:0] node50611;
	wire [4-1:0] node50614;
	wire [4-1:0] node50617;
	wire [4-1:0] node50618;
	wire [4-1:0] node50619;
	wire [4-1:0] node50622;
	wire [4-1:0] node50625;
	wire [4-1:0] node50626;
	wire [4-1:0] node50629;
	wire [4-1:0] node50632;
	wire [4-1:0] node50633;
	wire [4-1:0] node50634;
	wire [4-1:0] node50635;
	wire [4-1:0] node50636;
	wire [4-1:0] node50637;
	wire [4-1:0] node50641;
	wire [4-1:0] node50642;
	wire [4-1:0] node50646;
	wire [4-1:0] node50647;
	wire [4-1:0] node50650;
	wire [4-1:0] node50652;
	wire [4-1:0] node50655;
	wire [4-1:0] node50656;
	wire [4-1:0] node50658;
	wire [4-1:0] node50661;
	wire [4-1:0] node50662;
	wire [4-1:0] node50665;
	wire [4-1:0] node50668;
	wire [4-1:0] node50669;
	wire [4-1:0] node50670;
	wire [4-1:0] node50671;
	wire [4-1:0] node50672;
	wire [4-1:0] node50675;
	wire [4-1:0] node50678;
	wire [4-1:0] node50679;
	wire [4-1:0] node50682;
	wire [4-1:0] node50685;
	wire [4-1:0] node50687;
	wire [4-1:0] node50688;
	wire [4-1:0] node50691;
	wire [4-1:0] node50694;
	wire [4-1:0] node50695;
	wire [4-1:0] node50696;
	wire [4-1:0] node50697;
	wire [4-1:0] node50701;
	wire [4-1:0] node50702;
	wire [4-1:0] node50706;
	wire [4-1:0] node50709;
	wire [4-1:0] node50710;
	wire [4-1:0] node50711;
	wire [4-1:0] node50712;
	wire [4-1:0] node50713;
	wire [4-1:0] node50714;
	wire [4-1:0] node50717;
	wire [4-1:0] node50720;
	wire [4-1:0] node50721;
	wire [4-1:0] node50724;
	wire [4-1:0] node50727;
	wire [4-1:0] node50728;
	wire [4-1:0] node50731;
	wire [4-1:0] node50733;
	wire [4-1:0] node50736;
	wire [4-1:0] node50737;
	wire [4-1:0] node50738;
	wire [4-1:0] node50741;
	wire [4-1:0] node50743;
	wire [4-1:0] node50746;
	wire [4-1:0] node50747;
	wire [4-1:0] node50748;
	wire [4-1:0] node50751;
	wire [4-1:0] node50754;
	wire [4-1:0] node50755;
	wire [4-1:0] node50758;
	wire [4-1:0] node50761;
	wire [4-1:0] node50762;
	wire [4-1:0] node50763;
	wire [4-1:0] node50764;
	wire [4-1:0] node50765;
	wire [4-1:0] node50768;
	wire [4-1:0] node50771;
	wire [4-1:0] node50772;
	wire [4-1:0] node50775;
	wire [4-1:0] node50778;
	wire [4-1:0] node50779;
	wire [4-1:0] node50780;
	wire [4-1:0] node50782;
	wire [4-1:0] node50786;
	wire [4-1:0] node50787;
	wire [4-1:0] node50790;
	wire [4-1:0] node50793;
	wire [4-1:0] node50794;
	wire [4-1:0] node50795;
	wire [4-1:0] node50796;
	wire [4-1:0] node50799;
	wire [4-1:0] node50802;
	wire [4-1:0] node50803;
	wire [4-1:0] node50806;
	wire [4-1:0] node50809;
	wire [4-1:0] node50810;
	wire [4-1:0] node50812;
	wire [4-1:0] node50813;
	wire [4-1:0] node50816;
	wire [4-1:0] node50819;
	wire [4-1:0] node50820;
	wire [4-1:0] node50823;
	wire [4-1:0] node50826;
	wire [4-1:0] node50827;
	wire [4-1:0] node50828;
	wire [4-1:0] node50829;
	wire [4-1:0] node50830;
	wire [4-1:0] node50831;
	wire [4-1:0] node50832;
	wire [4-1:0] node50833;
	wire [4-1:0] node50836;
	wire [4-1:0] node50839;
	wire [4-1:0] node50840;
	wire [4-1:0] node50844;
	wire [4-1:0] node50845;
	wire [4-1:0] node50846;
	wire [4-1:0] node50849;
	wire [4-1:0] node50853;
	wire [4-1:0] node50854;
	wire [4-1:0] node50855;
	wire [4-1:0] node50856;
	wire [4-1:0] node50859;
	wire [4-1:0] node50862;
	wire [4-1:0] node50864;
	wire [4-1:0] node50867;
	wire [4-1:0] node50869;
	wire [4-1:0] node50870;
	wire [4-1:0] node50874;
	wire [4-1:0] node50875;
	wire [4-1:0] node50876;
	wire [4-1:0] node50878;
	wire [4-1:0] node50880;
	wire [4-1:0] node50883;
	wire [4-1:0] node50884;
	wire [4-1:0] node50885;
	wire [4-1:0] node50889;
	wire [4-1:0] node50890;
	wire [4-1:0] node50894;
	wire [4-1:0] node50895;
	wire [4-1:0] node50896;
	wire [4-1:0] node50897;
	wire [4-1:0] node50900;
	wire [4-1:0] node50903;
	wire [4-1:0] node50904;
	wire [4-1:0] node50907;
	wire [4-1:0] node50910;
	wire [4-1:0] node50911;
	wire [4-1:0] node50912;
	wire [4-1:0] node50916;
	wire [4-1:0] node50918;
	wire [4-1:0] node50921;
	wire [4-1:0] node50922;
	wire [4-1:0] node50923;
	wire [4-1:0] node50924;
	wire [4-1:0] node50925;
	wire [4-1:0] node50926;
	wire [4-1:0] node50929;
	wire [4-1:0] node50932;
	wire [4-1:0] node50933;
	wire [4-1:0] node50937;
	wire [4-1:0] node50938;
	wire [4-1:0] node50939;
	wire [4-1:0] node50942;
	wire [4-1:0] node50945;
	wire [4-1:0] node50946;
	wire [4-1:0] node50949;
	wire [4-1:0] node50952;
	wire [4-1:0] node50953;
	wire [4-1:0] node50954;
	wire [4-1:0] node50955;
	wire [4-1:0] node50958;
	wire [4-1:0] node50961;
	wire [4-1:0] node50964;
	wire [4-1:0] node50965;
	wire [4-1:0] node50967;
	wire [4-1:0] node50971;
	wire [4-1:0] node50972;
	wire [4-1:0] node50973;
	wire [4-1:0] node50974;
	wire [4-1:0] node50975;
	wire [4-1:0] node50978;
	wire [4-1:0] node50981;
	wire [4-1:0] node50984;
	wire [4-1:0] node50985;
	wire [4-1:0] node50988;
	wire [4-1:0] node50990;
	wire [4-1:0] node50993;
	wire [4-1:0] node50994;
	wire [4-1:0] node50995;
	wire [4-1:0] node50996;
	wire [4-1:0] node50999;
	wire [4-1:0] node51002;
	wire [4-1:0] node51003;
	wire [4-1:0] node51006;
	wire [4-1:0] node51009;
	wire [4-1:0] node51010;
	wire [4-1:0] node51013;
	wire [4-1:0] node51016;
	wire [4-1:0] node51017;
	wire [4-1:0] node51018;
	wire [4-1:0] node51019;
	wire [4-1:0] node51020;
	wire [4-1:0] node51021;
	wire [4-1:0] node51022;
	wire [4-1:0] node51025;
	wire [4-1:0] node51029;
	wire [4-1:0] node51030;
	wire [4-1:0] node51033;
	wire [4-1:0] node51036;
	wire [4-1:0] node51037;
	wire [4-1:0] node51038;
	wire [4-1:0] node51041;
	wire [4-1:0] node51043;
	wire [4-1:0] node51046;
	wire [4-1:0] node51047;
	wire [4-1:0] node51050;
	wire [4-1:0] node51053;
	wire [4-1:0] node51054;
	wire [4-1:0] node51055;
	wire [4-1:0] node51058;
	wire [4-1:0] node51060;
	wire [4-1:0] node51063;
	wire [4-1:0] node51064;
	wire [4-1:0] node51066;
	wire [4-1:0] node51067;
	wire [4-1:0] node51070;
	wire [4-1:0] node51073;
	wire [4-1:0] node51074;
	wire [4-1:0] node51077;
	wire [4-1:0] node51080;
	wire [4-1:0] node51081;
	wire [4-1:0] node51082;
	wire [4-1:0] node51083;
	wire [4-1:0] node51085;
	wire [4-1:0] node51086;
	wire [4-1:0] node51090;
	wire [4-1:0] node51091;
	wire [4-1:0] node51092;
	wire [4-1:0] node51095;
	wire [4-1:0] node51099;
	wire [4-1:0] node51100;
	wire [4-1:0] node51101;
	wire [4-1:0] node51104;
	wire [4-1:0] node51107;
	wire [4-1:0] node51108;
	wire [4-1:0] node51111;
	wire [4-1:0] node51114;
	wire [4-1:0] node51115;
	wire [4-1:0] node51116;
	wire [4-1:0] node51117;
	wire [4-1:0] node51120;
	wire [4-1:0] node51121;
	wire [4-1:0] node51124;
	wire [4-1:0] node51127;
	wire [4-1:0] node51129;
	wire [4-1:0] node51130;
	wire [4-1:0] node51133;
	wire [4-1:0] node51136;
	wire [4-1:0] node51137;
	wire [4-1:0] node51140;
	wire [4-1:0] node51141;
	wire [4-1:0] node51142;
	wire [4-1:0] node51145;
	wire [4-1:0] node51149;
	wire [4-1:0] node51150;
	wire [4-1:0] node51151;
	wire [4-1:0] node51152;
	wire [4-1:0] node51153;
	wire [4-1:0] node51154;
	wire [4-1:0] node51155;
	wire [4-1:0] node51156;
	wire [4-1:0] node51157;
	wire [4-1:0] node51158;
	wire [4-1:0] node51162;
	wire [4-1:0] node51163;
	wire [4-1:0] node51166;
	wire [4-1:0] node51169;
	wire [4-1:0] node51170;
	wire [4-1:0] node51172;
	wire [4-1:0] node51175;
	wire [4-1:0] node51176;
	wire [4-1:0] node51180;
	wire [4-1:0] node51181;
	wire [4-1:0] node51183;
	wire [4-1:0] node51185;
	wire [4-1:0] node51188;
	wire [4-1:0] node51189;
	wire [4-1:0] node51191;
	wire [4-1:0] node51195;
	wire [4-1:0] node51196;
	wire [4-1:0] node51197;
	wire [4-1:0] node51198;
	wire [4-1:0] node51201;
	wire [4-1:0] node51204;
	wire [4-1:0] node51205;
	wire [4-1:0] node51208;
	wire [4-1:0] node51211;
	wire [4-1:0] node51212;
	wire [4-1:0] node51214;
	wire [4-1:0] node51217;
	wire [4-1:0] node51218;
	wire [4-1:0] node51222;
	wire [4-1:0] node51223;
	wire [4-1:0] node51224;
	wire [4-1:0] node51225;
	wire [4-1:0] node51226;
	wire [4-1:0] node51229;
	wire [4-1:0] node51232;
	wire [4-1:0] node51233;
	wire [4-1:0] node51236;
	wire [4-1:0] node51238;
	wire [4-1:0] node51241;
	wire [4-1:0] node51242;
	wire [4-1:0] node51243;
	wire [4-1:0] node51246;
	wire [4-1:0] node51249;
	wire [4-1:0] node51250;
	wire [4-1:0] node51253;
	wire [4-1:0] node51256;
	wire [4-1:0] node51257;
	wire [4-1:0] node51258;
	wire [4-1:0] node51259;
	wire [4-1:0] node51262;
	wire [4-1:0] node51265;
	wire [4-1:0] node51266;
	wire [4-1:0] node51269;
	wire [4-1:0] node51272;
	wire [4-1:0] node51273;
	wire [4-1:0] node51274;
	wire [4-1:0] node51277;
	wire [4-1:0] node51280;
	wire [4-1:0] node51281;
	wire [4-1:0] node51283;
	wire [4-1:0] node51286;
	wire [4-1:0] node51288;
	wire [4-1:0] node51291;
	wire [4-1:0] node51292;
	wire [4-1:0] node51293;
	wire [4-1:0] node51294;
	wire [4-1:0] node51295;
	wire [4-1:0] node51298;
	wire [4-1:0] node51301;
	wire [4-1:0] node51302;
	wire [4-1:0] node51303;
	wire [4-1:0] node51306;
	wire [4-1:0] node51309;
	wire [4-1:0] node51311;
	wire [4-1:0] node51312;
	wire [4-1:0] node51315;
	wire [4-1:0] node51318;
	wire [4-1:0] node51319;
	wire [4-1:0] node51320;
	wire [4-1:0] node51323;
	wire [4-1:0] node51326;
	wire [4-1:0] node51327;
	wire [4-1:0] node51330;
	wire [4-1:0] node51333;
	wire [4-1:0] node51334;
	wire [4-1:0] node51335;
	wire [4-1:0] node51336;
	wire [4-1:0] node51339;
	wire [4-1:0] node51342;
	wire [4-1:0] node51343;
	wire [4-1:0] node51346;
	wire [4-1:0] node51349;
	wire [4-1:0] node51350;
	wire [4-1:0] node51351;
	wire [4-1:0] node51354;
	wire [4-1:0] node51357;
	wire [4-1:0] node51358;
	wire [4-1:0] node51361;
	wire [4-1:0] node51364;
	wire [4-1:0] node51365;
	wire [4-1:0] node51366;
	wire [4-1:0] node51367;
	wire [4-1:0] node51368;
	wire [4-1:0] node51370;
	wire [4-1:0] node51371;
	wire [4-1:0] node51372;
	wire [4-1:0] node51376;
	wire [4-1:0] node51378;
	wire [4-1:0] node51381;
	wire [4-1:0] node51382;
	wire [4-1:0] node51383;
	wire [4-1:0] node51386;
	wire [4-1:0] node51389;
	wire [4-1:0] node51390;
	wire [4-1:0] node51392;
	wire [4-1:0] node51396;
	wire [4-1:0] node51397;
	wire [4-1:0] node51398;
	wire [4-1:0] node51399;
	wire [4-1:0] node51402;
	wire [4-1:0] node51405;
	wire [4-1:0] node51407;
	wire [4-1:0] node51410;
	wire [4-1:0] node51411;
	wire [4-1:0] node51413;
	wire [4-1:0] node51414;
	wire [4-1:0] node51417;
	wire [4-1:0] node51420;
	wire [4-1:0] node51421;
	wire [4-1:0] node51424;
	wire [4-1:0] node51427;
	wire [4-1:0] node51428;
	wire [4-1:0] node51429;
	wire [4-1:0] node51430;
	wire [4-1:0] node51433;
	wire [4-1:0] node51436;
	wire [4-1:0] node51437;
	wire [4-1:0] node51439;
	wire [4-1:0] node51440;
	wire [4-1:0] node51443;
	wire [4-1:0] node51447;
	wire [4-1:0] node51448;
	wire [4-1:0] node51450;
	wire [4-1:0] node51451;
	wire [4-1:0] node51453;
	wire [4-1:0] node51456;
	wire [4-1:0] node51459;
	wire [4-1:0] node51460;
	wire [4-1:0] node51462;
	wire [4-1:0] node51465;
	wire [4-1:0] node51466;
	wire [4-1:0] node51470;
	wire [4-1:0] node51471;
	wire [4-1:0] node51472;
	wire [4-1:0] node51473;
	wire [4-1:0] node51474;
	wire [4-1:0] node51477;
	wire [4-1:0] node51478;
	wire [4-1:0] node51481;
	wire [4-1:0] node51484;
	wire [4-1:0] node51486;
	wire [4-1:0] node51487;
	wire [4-1:0] node51490;
	wire [4-1:0] node51493;
	wire [4-1:0] node51494;
	wire [4-1:0] node51495;
	wire [4-1:0] node51496;
	wire [4-1:0] node51498;
	wire [4-1:0] node51501;
	wire [4-1:0] node51502;
	wire [4-1:0] node51505;
	wire [4-1:0] node51508;
	wire [4-1:0] node51509;
	wire [4-1:0] node51512;
	wire [4-1:0] node51515;
	wire [4-1:0] node51516;
	wire [4-1:0] node51517;
	wire [4-1:0] node51521;
	wire [4-1:0] node51522;
	wire [4-1:0] node51525;
	wire [4-1:0] node51528;
	wire [4-1:0] node51529;
	wire [4-1:0] node51530;
	wire [4-1:0] node51532;
	wire [4-1:0] node51533;
	wire [4-1:0] node51536;
	wire [4-1:0] node51539;
	wire [4-1:0] node51540;
	wire [4-1:0] node51541;
	wire [4-1:0] node51544;
	wire [4-1:0] node51547;
	wire [4-1:0] node51549;
	wire [4-1:0] node51552;
	wire [4-1:0] node51553;
	wire [4-1:0] node51554;
	wire [4-1:0] node51556;
	wire [4-1:0] node51559;
	wire [4-1:0] node51560;
	wire [4-1:0] node51562;
	wire [4-1:0] node51565;
	wire [4-1:0] node51567;
	wire [4-1:0] node51570;
	wire [4-1:0] node51571;
	wire [4-1:0] node51573;
	wire [4-1:0] node51576;
	wire [4-1:0] node51577;
	wire [4-1:0] node51580;
	wire [4-1:0] node51583;
	wire [4-1:0] node51584;
	wire [4-1:0] node51585;
	wire [4-1:0] node51586;
	wire [4-1:0] node51587;
	wire [4-1:0] node51588;
	wire [4-1:0] node51589;
	wire [4-1:0] node51590;
	wire [4-1:0] node51591;
	wire [4-1:0] node51594;
	wire [4-1:0] node51597;
	wire [4-1:0] node51598;
	wire [4-1:0] node51601;
	wire [4-1:0] node51605;
	wire [4-1:0] node51606;
	wire [4-1:0] node51607;
	wire [4-1:0] node51610;
	wire [4-1:0] node51613;
	wire [4-1:0] node51614;
	wire [4-1:0] node51617;
	wire [4-1:0] node51620;
	wire [4-1:0] node51621;
	wire [4-1:0] node51622;
	wire [4-1:0] node51624;
	wire [4-1:0] node51627;
	wire [4-1:0] node51630;
	wire [4-1:0] node51631;
	wire [4-1:0] node51632;
	wire [4-1:0] node51634;
	wire [4-1:0] node51637;
	wire [4-1:0] node51640;
	wire [4-1:0] node51641;
	wire [4-1:0] node51644;
	wire [4-1:0] node51647;
	wire [4-1:0] node51648;
	wire [4-1:0] node51649;
	wire [4-1:0] node51650;
	wire [4-1:0] node51652;
	wire [4-1:0] node51655;
	wire [4-1:0] node51656;
	wire [4-1:0] node51657;
	wire [4-1:0] node51660;
	wire [4-1:0] node51663;
	wire [4-1:0] node51665;
	wire [4-1:0] node51668;
	wire [4-1:0] node51669;
	wire [4-1:0] node51670;
	wire [4-1:0] node51671;
	wire [4-1:0] node51675;
	wire [4-1:0] node51676;
	wire [4-1:0] node51680;
	wire [4-1:0] node51681;
	wire [4-1:0] node51682;
	wire [4-1:0] node51686;
	wire [4-1:0] node51687;
	wire [4-1:0] node51690;
	wire [4-1:0] node51693;
	wire [4-1:0] node51694;
	wire [4-1:0] node51695;
	wire [4-1:0] node51696;
	wire [4-1:0] node51699;
	wire [4-1:0] node51702;
	wire [4-1:0] node51703;
	wire [4-1:0] node51704;
	wire [4-1:0] node51707;
	wire [4-1:0] node51711;
	wire [4-1:0] node51712;
	wire [4-1:0] node51713;
	wire [4-1:0] node51714;
	wire [4-1:0] node51718;
	wire [4-1:0] node51719;
	wire [4-1:0] node51723;
	wire [4-1:0] node51724;
	wire [4-1:0] node51727;
	wire [4-1:0] node51730;
	wire [4-1:0] node51731;
	wire [4-1:0] node51732;
	wire [4-1:0] node51733;
	wire [4-1:0] node51734;
	wire [4-1:0] node51735;
	wire [4-1:0] node51738;
	wire [4-1:0] node51741;
	wire [4-1:0] node51743;
	wire [4-1:0] node51746;
	wire [4-1:0] node51747;
	wire [4-1:0] node51750;
	wire [4-1:0] node51753;
	wire [4-1:0] node51754;
	wire [4-1:0] node51755;
	wire [4-1:0] node51758;
	wire [4-1:0] node51761;
	wire [4-1:0] node51762;
	wire [4-1:0] node51765;
	wire [4-1:0] node51768;
	wire [4-1:0] node51769;
	wire [4-1:0] node51770;
	wire [4-1:0] node51771;
	wire [4-1:0] node51772;
	wire [4-1:0] node51775;
	wire [4-1:0] node51776;
	wire [4-1:0] node51780;
	wire [4-1:0] node51781;
	wire [4-1:0] node51784;
	wire [4-1:0] node51786;
	wire [4-1:0] node51789;
	wire [4-1:0] node51790;
	wire [4-1:0] node51791;
	wire [4-1:0] node51792;
	wire [4-1:0] node51796;
	wire [4-1:0] node51797;
	wire [4-1:0] node51800;
	wire [4-1:0] node51803;
	wire [4-1:0] node51804;
	wire [4-1:0] node51805;
	wire [4-1:0] node51809;
	wire [4-1:0] node51811;
	wire [4-1:0] node51814;
	wire [4-1:0] node51815;
	wire [4-1:0] node51816;
	wire [4-1:0] node51817;
	wire [4-1:0] node51818;
	wire [4-1:0] node51821;
	wire [4-1:0] node51824;
	wire [4-1:0] node51825;
	wire [4-1:0] node51828;
	wire [4-1:0] node51831;
	wire [4-1:0] node51832;
	wire [4-1:0] node51834;
	wire [4-1:0] node51837;
	wire [4-1:0] node51839;
	wire [4-1:0] node51842;
	wire [4-1:0] node51843;
	wire [4-1:0] node51844;
	wire [4-1:0] node51845;
	wire [4-1:0] node51850;
	wire [4-1:0] node51851;
	wire [4-1:0] node51852;
	wire [4-1:0] node51856;
	wire [4-1:0] node51859;
	wire [4-1:0] node51860;
	wire [4-1:0] node51861;
	wire [4-1:0] node51862;
	wire [4-1:0] node51863;
	wire [4-1:0] node51864;
	wire [4-1:0] node51865;
	wire [4-1:0] node51866;
	wire [4-1:0] node51869;
	wire [4-1:0] node51873;
	wire [4-1:0] node51874;
	wire [4-1:0] node51875;
	wire [4-1:0] node51880;
	wire [4-1:0] node51881;
	wire [4-1:0] node51882;
	wire [4-1:0] node51886;
	wire [4-1:0] node51888;
	wire [4-1:0] node51891;
	wire [4-1:0] node51892;
	wire [4-1:0] node51893;
	wire [4-1:0] node51894;
	wire [4-1:0] node51897;
	wire [4-1:0] node51900;
	wire [4-1:0] node51902;
	wire [4-1:0] node51905;
	wire [4-1:0] node51906;
	wire [4-1:0] node51908;
	wire [4-1:0] node51911;
	wire [4-1:0] node51912;
	wire [4-1:0] node51915;
	wire [4-1:0] node51918;
	wire [4-1:0] node51919;
	wire [4-1:0] node51920;
	wire [4-1:0] node51921;
	wire [4-1:0] node51924;
	wire [4-1:0] node51927;
	wire [4-1:0] node51928;
	wire [4-1:0] node51929;
	wire [4-1:0] node51932;
	wire [4-1:0] node51935;
	wire [4-1:0] node51937;
	wire [4-1:0] node51940;
	wire [4-1:0] node51941;
	wire [4-1:0] node51942;
	wire [4-1:0] node51943;
	wire [4-1:0] node51944;
	wire [4-1:0] node51947;
	wire [4-1:0] node51951;
	wire [4-1:0] node51952;
	wire [4-1:0] node51953;
	wire [4-1:0] node51958;
	wire [4-1:0] node51959;
	wire [4-1:0] node51961;
	wire [4-1:0] node51962;
	wire [4-1:0] node51966;
	wire [4-1:0] node51967;
	wire [4-1:0] node51968;
	wire [4-1:0] node51973;
	wire [4-1:0] node51974;
	wire [4-1:0] node51975;
	wire [4-1:0] node51976;
	wire [4-1:0] node51977;
	wire [4-1:0] node51980;
	wire [4-1:0] node51983;
	wire [4-1:0] node51984;
	wire [4-1:0] node51987;
	wire [4-1:0] node51990;
	wire [4-1:0] node51991;
	wire [4-1:0] node51992;
	wire [4-1:0] node51993;
	wire [4-1:0] node51996;
	wire [4-1:0] node51999;
	wire [4-1:0] node52001;
	wire [4-1:0] node52004;
	wire [4-1:0] node52005;
	wire [4-1:0] node52008;
	wire [4-1:0] node52011;
	wire [4-1:0] node52012;
	wire [4-1:0] node52013;
	wire [4-1:0] node52014;
	wire [4-1:0] node52015;
	wire [4-1:0] node52016;
	wire [4-1:0] node52020;
	wire [4-1:0] node52021;
	wire [4-1:0] node52024;
	wire [4-1:0] node52027;
	wire [4-1:0] node52028;
	wire [4-1:0] node52029;
	wire [4-1:0] node52032;
	wire [4-1:0] node52035;
	wire [4-1:0] node52036;
	wire [4-1:0] node52039;
	wire [4-1:0] node52042;
	wire [4-1:0] node52043;
	wire [4-1:0] node52046;
	wire [4-1:0] node52049;
	wire [4-1:0] node52050;
	wire [4-1:0] node52051;
	wire [4-1:0] node52052;
	wire [4-1:0] node52055;
	wire [4-1:0] node52058;
	wire [4-1:0] node52060;
	wire [4-1:0] node52063;
	wire [4-1:0] node52064;
	wire [4-1:0] node52067;
	wire [4-1:0] node52070;
	wire [4-1:0] node52071;
	wire [4-1:0] node52072;
	wire [4-1:0] node52073;
	wire [4-1:0] node52074;
	wire [4-1:0] node52075;
	wire [4-1:0] node52076;
	wire [4-1:0] node52077;
	wire [4-1:0] node52078;
	wire [4-1:0] node52079;
	wire [4-1:0] node52080;
	wire [4-1:0] node52084;
	wire [4-1:0] node52087;
	wire [4-1:0] node52089;
	wire [4-1:0] node52090;
	wire [4-1:0] node52093;
	wire [4-1:0] node52096;
	wire [4-1:0] node52097;
	wire [4-1:0] node52098;
	wire [4-1:0] node52099;
	wire [4-1:0] node52103;
	wire [4-1:0] node52105;
	wire [4-1:0] node52108;
	wire [4-1:0] node52109;
	wire [4-1:0] node52110;
	wire [4-1:0] node52114;
	wire [4-1:0] node52115;
	wire [4-1:0] node52118;
	wire [4-1:0] node52121;
	wire [4-1:0] node52122;
	wire [4-1:0] node52123;
	wire [4-1:0] node52124;
	wire [4-1:0] node52127;
	wire [4-1:0] node52129;
	wire [4-1:0] node52132;
	wire [4-1:0] node52133;
	wire [4-1:0] node52134;
	wire [4-1:0] node52137;
	wire [4-1:0] node52140;
	wire [4-1:0] node52142;
	wire [4-1:0] node52145;
	wire [4-1:0] node52146;
	wire [4-1:0] node52147;
	wire [4-1:0] node52148;
	wire [4-1:0] node52151;
	wire [4-1:0] node52154;
	wire [4-1:0] node52155;
	wire [4-1:0] node52158;
	wire [4-1:0] node52161;
	wire [4-1:0] node52162;
	wire [4-1:0] node52163;
	wire [4-1:0] node52166;
	wire [4-1:0] node52170;
	wire [4-1:0] node52171;
	wire [4-1:0] node52172;
	wire [4-1:0] node52173;
	wire [4-1:0] node52174;
	wire [4-1:0] node52175;
	wire [4-1:0] node52178;
	wire [4-1:0] node52182;
	wire [4-1:0] node52183;
	wire [4-1:0] node52184;
	wire [4-1:0] node52188;
	wire [4-1:0] node52189;
	wire [4-1:0] node52192;
	wire [4-1:0] node52195;
	wire [4-1:0] node52196;
	wire [4-1:0] node52197;
	wire [4-1:0] node52201;
	wire [4-1:0] node52202;
	wire [4-1:0] node52205;
	wire [4-1:0] node52208;
	wire [4-1:0] node52209;
	wire [4-1:0] node52210;
	wire [4-1:0] node52211;
	wire [4-1:0] node52212;
	wire [4-1:0] node52216;
	wire [4-1:0] node52219;
	wire [4-1:0] node52220;
	wire [4-1:0] node52223;
	wire [4-1:0] node52225;
	wire [4-1:0] node52228;
	wire [4-1:0] node52229;
	wire [4-1:0] node52230;
	wire [4-1:0] node52231;
	wire [4-1:0] node52235;
	wire [4-1:0] node52238;
	wire [4-1:0] node52239;
	wire [4-1:0] node52242;
	wire [4-1:0] node52245;
	wire [4-1:0] node52246;
	wire [4-1:0] node52247;
	wire [4-1:0] node52248;
	wire [4-1:0] node52249;
	wire [4-1:0] node52250;
	wire [4-1:0] node52253;
	wire [4-1:0] node52256;
	wire [4-1:0] node52257;
	wire [4-1:0] node52258;
	wire [4-1:0] node52263;
	wire [4-1:0] node52264;
	wire [4-1:0] node52266;
	wire [4-1:0] node52268;
	wire [4-1:0] node52271;
	wire [4-1:0] node52272;
	wire [4-1:0] node52275;
	wire [4-1:0] node52278;
	wire [4-1:0] node52279;
	wire [4-1:0] node52280;
	wire [4-1:0] node52281;
	wire [4-1:0] node52282;
	wire [4-1:0] node52285;
	wire [4-1:0] node52288;
	wire [4-1:0] node52289;
	wire [4-1:0] node52292;
	wire [4-1:0] node52295;
	wire [4-1:0] node52297;
	wire [4-1:0] node52300;
	wire [4-1:0] node52301;
	wire [4-1:0] node52303;
	wire [4-1:0] node52304;
	wire [4-1:0] node52307;
	wire [4-1:0] node52310;
	wire [4-1:0] node52311;
	wire [4-1:0] node52315;
	wire [4-1:0] node52316;
	wire [4-1:0] node52317;
	wire [4-1:0] node52318;
	wire [4-1:0] node52320;
	wire [4-1:0] node52323;
	wire [4-1:0] node52324;
	wire [4-1:0] node52326;
	wire [4-1:0] node52329;
	wire [4-1:0] node52332;
	wire [4-1:0] node52333;
	wire [4-1:0] node52334;
	wire [4-1:0] node52338;
	wire [4-1:0] node52339;
	wire [4-1:0] node52342;
	wire [4-1:0] node52343;
	wire [4-1:0] node52347;
	wire [4-1:0] node52348;
	wire [4-1:0] node52349;
	wire [4-1:0] node52350;
	wire [4-1:0] node52351;
	wire [4-1:0] node52354;
	wire [4-1:0] node52357;
	wire [4-1:0] node52358;
	wire [4-1:0] node52362;
	wire [4-1:0] node52364;
	wire [4-1:0] node52367;
	wire [4-1:0] node52368;
	wire [4-1:0] node52370;
	wire [4-1:0] node52371;
	wire [4-1:0] node52375;
	wire [4-1:0] node52377;
	wire [4-1:0] node52380;
	wire [4-1:0] node52381;
	wire [4-1:0] node52382;
	wire [4-1:0] node52383;
	wire [4-1:0] node52384;
	wire [4-1:0] node52385;
	wire [4-1:0] node52387;
	wire [4-1:0] node52388;
	wire [4-1:0] node52391;
	wire [4-1:0] node52394;
	wire [4-1:0] node52396;
	wire [4-1:0] node52397;
	wire [4-1:0] node52401;
	wire [4-1:0] node52402;
	wire [4-1:0] node52403;
	wire [4-1:0] node52404;
	wire [4-1:0] node52407;
	wire [4-1:0] node52411;
	wire [4-1:0] node52413;
	wire [4-1:0] node52414;
	wire [4-1:0] node52417;
	wire [4-1:0] node52420;
	wire [4-1:0] node52421;
	wire [4-1:0] node52422;
	wire [4-1:0] node52423;
	wire [4-1:0] node52426;
	wire [4-1:0] node52428;
	wire [4-1:0] node52431;
	wire [4-1:0] node52433;
	wire [4-1:0] node52434;
	wire [4-1:0] node52438;
	wire [4-1:0] node52439;
	wire [4-1:0] node52442;
	wire [4-1:0] node52443;
	wire [4-1:0] node52446;
	wire [4-1:0] node52448;
	wire [4-1:0] node52451;
	wire [4-1:0] node52452;
	wire [4-1:0] node52453;
	wire [4-1:0] node52454;
	wire [4-1:0] node52456;
	wire [4-1:0] node52459;
	wire [4-1:0] node52460;
	wire [4-1:0] node52463;
	wire [4-1:0] node52466;
	wire [4-1:0] node52467;
	wire [4-1:0] node52468;
	wire [4-1:0] node52471;
	wire [4-1:0] node52474;
	wire [4-1:0] node52475;
	wire [4-1:0] node52479;
	wire [4-1:0] node52480;
	wire [4-1:0] node52481;
	wire [4-1:0] node52482;
	wire [4-1:0] node52483;
	wire [4-1:0] node52486;
	wire [4-1:0] node52489;
	wire [4-1:0] node52490;
	wire [4-1:0] node52494;
	wire [4-1:0] node52495;
	wire [4-1:0] node52499;
	wire [4-1:0] node52500;
	wire [4-1:0] node52501;
	wire [4-1:0] node52504;
	wire [4-1:0] node52507;
	wire [4-1:0] node52508;
	wire [4-1:0] node52509;
	wire [4-1:0] node52512;
	wire [4-1:0] node52516;
	wire [4-1:0] node52517;
	wire [4-1:0] node52518;
	wire [4-1:0] node52519;
	wire [4-1:0] node52520;
	wire [4-1:0] node52523;
	wire [4-1:0] node52526;
	wire [4-1:0] node52527;
	wire [4-1:0] node52530;
	wire [4-1:0] node52533;
	wire [4-1:0] node52534;
	wire [4-1:0] node52535;
	wire [4-1:0] node52536;
	wire [4-1:0] node52539;
	wire [4-1:0] node52542;
	wire [4-1:0] node52543;
	wire [4-1:0] node52546;
	wire [4-1:0] node52549;
	wire [4-1:0] node52550;
	wire [4-1:0] node52551;
	wire [4-1:0] node52555;
	wire [4-1:0] node52558;
	wire [4-1:0] node52559;
	wire [4-1:0] node52560;
	wire [4-1:0] node52561;
	wire [4-1:0] node52564;
	wire [4-1:0] node52567;
	wire [4-1:0] node52569;
	wire [4-1:0] node52572;
	wire [4-1:0] node52573;
	wire [4-1:0] node52574;
	wire [4-1:0] node52578;
	wire [4-1:0] node52581;
	wire [4-1:0] node52582;
	wire [4-1:0] node52583;
	wire [4-1:0] node52584;
	wire [4-1:0] node52585;
	wire [4-1:0] node52586;
	wire [4-1:0] node52587;
	wire [4-1:0] node52588;
	wire [4-1:0] node52589;
	wire [4-1:0] node52593;
	wire [4-1:0] node52594;
	wire [4-1:0] node52597;
	wire [4-1:0] node52600;
	wire [4-1:0] node52601;
	wire [4-1:0] node52603;
	wire [4-1:0] node52606;
	wire [4-1:0] node52608;
	wire [4-1:0] node52611;
	wire [4-1:0] node52612;
	wire [4-1:0] node52613;
	wire [4-1:0] node52616;
	wire [4-1:0] node52619;
	wire [4-1:0] node52620;
	wire [4-1:0] node52623;
	wire [4-1:0] node52626;
	wire [4-1:0] node52627;
	wire [4-1:0] node52628;
	wire [4-1:0] node52629;
	wire [4-1:0] node52631;
	wire [4-1:0] node52634;
	wire [4-1:0] node52635;
	wire [4-1:0] node52638;
	wire [4-1:0] node52641;
	wire [4-1:0] node52642;
	wire [4-1:0] node52645;
	wire [4-1:0] node52648;
	wire [4-1:0] node52649;
	wire [4-1:0] node52652;
	wire [4-1:0] node52655;
	wire [4-1:0] node52656;
	wire [4-1:0] node52657;
	wire [4-1:0] node52658;
	wire [4-1:0] node52659;
	wire [4-1:0] node52661;
	wire [4-1:0] node52665;
	wire [4-1:0] node52666;
	wire [4-1:0] node52669;
	wire [4-1:0] node52672;
	wire [4-1:0] node52673;
	wire [4-1:0] node52676;
	wire [4-1:0] node52679;
	wire [4-1:0] node52680;
	wire [4-1:0] node52681;
	wire [4-1:0] node52682;
	wire [4-1:0] node52685;
	wire [4-1:0] node52688;
	wire [4-1:0] node52689;
	wire [4-1:0] node52692;
	wire [4-1:0] node52695;
	wire [4-1:0] node52696;
	wire [4-1:0] node52699;
	wire [4-1:0] node52702;
	wire [4-1:0] node52703;
	wire [4-1:0] node52704;
	wire [4-1:0] node52705;
	wire [4-1:0] node52706;
	wire [4-1:0] node52707;
	wire [4-1:0] node52708;
	wire [4-1:0] node52711;
	wire [4-1:0] node52714;
	wire [4-1:0] node52715;
	wire [4-1:0] node52718;
	wire [4-1:0] node52721;
	wire [4-1:0] node52722;
	wire [4-1:0] node52723;
	wire [4-1:0] node52726;
	wire [4-1:0] node52729;
	wire [4-1:0] node52730;
	wire [4-1:0] node52734;
	wire [4-1:0] node52735;
	wire [4-1:0] node52736;
	wire [4-1:0] node52738;
	wire [4-1:0] node52741;
	wire [4-1:0] node52742;
	wire [4-1:0] node52745;
	wire [4-1:0] node52748;
	wire [4-1:0] node52749;
	wire [4-1:0] node52750;
	wire [4-1:0] node52753;
	wire [4-1:0] node52756;
	wire [4-1:0] node52757;
	wire [4-1:0] node52761;
	wire [4-1:0] node52762;
	wire [4-1:0] node52763;
	wire [4-1:0] node52764;
	wire [4-1:0] node52765;
	wire [4-1:0] node52768;
	wire [4-1:0] node52772;
	wire [4-1:0] node52774;
	wire [4-1:0] node52776;
	wire [4-1:0] node52779;
	wire [4-1:0] node52780;
	wire [4-1:0] node52783;
	wire [4-1:0] node52786;
	wire [4-1:0] node52787;
	wire [4-1:0] node52788;
	wire [4-1:0] node52789;
	wire [4-1:0] node52790;
	wire [4-1:0] node52791;
	wire [4-1:0] node52794;
	wire [4-1:0] node52798;
	wire [4-1:0] node52799;
	wire [4-1:0] node52800;
	wire [4-1:0] node52804;
	wire [4-1:0] node52806;
	wire [4-1:0] node52809;
	wire [4-1:0] node52810;
	wire [4-1:0] node52811;
	wire [4-1:0] node52812;
	wire [4-1:0] node52815;
	wire [4-1:0] node52818;
	wire [4-1:0] node52819;
	wire [4-1:0] node52822;
	wire [4-1:0] node52825;
	wire [4-1:0] node52826;
	wire [4-1:0] node52828;
	wire [4-1:0] node52831;
	wire [4-1:0] node52832;
	wire [4-1:0] node52836;
	wire [4-1:0] node52837;
	wire [4-1:0] node52838;
	wire [4-1:0] node52839;
	wire [4-1:0] node52840;
	wire [4-1:0] node52843;
	wire [4-1:0] node52846;
	wire [4-1:0] node52847;
	wire [4-1:0] node52851;
	wire [4-1:0] node52852;
	wire [4-1:0] node52856;
	wire [4-1:0] node52857;
	wire [4-1:0] node52860;
	wire [4-1:0] node52863;
	wire [4-1:0] node52864;
	wire [4-1:0] node52865;
	wire [4-1:0] node52866;
	wire [4-1:0] node52867;
	wire [4-1:0] node52868;
	wire [4-1:0] node52869;
	wire [4-1:0] node52873;
	wire [4-1:0] node52874;
	wire [4-1:0] node52878;
	wire [4-1:0] node52879;
	wire [4-1:0] node52880;
	wire [4-1:0] node52884;
	wire [4-1:0] node52885;
	wire [4-1:0] node52889;
	wire [4-1:0] node52890;
	wire [4-1:0] node52891;
	wire [4-1:0] node52893;
	wire [4-1:0] node52895;
	wire [4-1:0] node52898;
	wire [4-1:0] node52900;
	wire [4-1:0] node52903;
	wire [4-1:0] node52904;
	wire [4-1:0] node52907;
	wire [4-1:0] node52910;
	wire [4-1:0] node52911;
	wire [4-1:0] node52912;
	wire [4-1:0] node52913;
	wire [4-1:0] node52914;
	wire [4-1:0] node52918;
	wire [4-1:0] node52919;
	wire [4-1:0] node52923;
	wire [4-1:0] node52924;
	wire [4-1:0] node52925;
	wire [4-1:0] node52926;
	wire [4-1:0] node52931;
	wire [4-1:0] node52932;
	wire [4-1:0] node52936;
	wire [4-1:0] node52937;
	wire [4-1:0] node52938;
	wire [4-1:0] node52939;
	wire [4-1:0] node52940;
	wire [4-1:0] node52943;
	wire [4-1:0] node52946;
	wire [4-1:0] node52947;
	wire [4-1:0] node52950;
	wire [4-1:0] node52953;
	wire [4-1:0] node52954;
	wire [4-1:0] node52957;
	wire [4-1:0] node52960;
	wire [4-1:0] node52961;
	wire [4-1:0] node52964;
	wire [4-1:0] node52967;
	wire [4-1:0] node52968;
	wire [4-1:0] node52969;
	wire [4-1:0] node52970;
	wire [4-1:0] node52971;
	wire [4-1:0] node52972;
	wire [4-1:0] node52976;
	wire [4-1:0] node52977;
	wire [4-1:0] node52981;
	wire [4-1:0] node52982;
	wire [4-1:0] node52983;
	wire [4-1:0] node52987;
	wire [4-1:0] node52988;
	wire [4-1:0] node52992;
	wire [4-1:0] node52993;
	wire [4-1:0] node52994;
	wire [4-1:0] node52996;
	wire [4-1:0] node52999;
	wire [4-1:0] node53001;
	wire [4-1:0] node53002;
	wire [4-1:0] node53006;
	wire [4-1:0] node53007;
	wire [4-1:0] node53009;
	wire [4-1:0] node53011;
	wire [4-1:0] node53014;
	wire [4-1:0] node53015;
	wire [4-1:0] node53018;
	wire [4-1:0] node53021;
	wire [4-1:0] node53022;
	wire [4-1:0] node53023;
	wire [4-1:0] node53024;
	wire [4-1:0] node53025;
	wire [4-1:0] node53029;
	wire [4-1:0] node53030;
	wire [4-1:0] node53034;
	wire [4-1:0] node53035;
	wire [4-1:0] node53036;
	wire [4-1:0] node53040;
	wire [4-1:0] node53041;
	wire [4-1:0] node53045;
	wire [4-1:0] node53046;
	wire [4-1:0] node53047;
	wire [4-1:0] node53048;
	wire [4-1:0] node53052;
	wire [4-1:0] node53053;
	wire [4-1:0] node53057;
	wire [4-1:0] node53058;
	wire [4-1:0] node53059;
	wire [4-1:0] node53063;
	wire [4-1:0] node53064;
	wire [4-1:0] node53068;
	wire [4-1:0] node53069;
	wire [4-1:0] node53070;
	wire [4-1:0] node53071;
	wire [4-1:0] node53072;
	wire [4-1:0] node53073;
	wire [4-1:0] node53074;
	wire [4-1:0] node53075;
	wire [4-1:0] node53076;
	wire [4-1:0] node53077;
	wire [4-1:0] node53080;
	wire [4-1:0] node53083;
	wire [4-1:0] node53085;
	wire [4-1:0] node53088;
	wire [4-1:0] node53089;
	wire [4-1:0] node53090;
	wire [4-1:0] node53094;
	wire [4-1:0] node53096;
	wire [4-1:0] node53099;
	wire [4-1:0] node53100;
	wire [4-1:0] node53102;
	wire [4-1:0] node53103;
	wire [4-1:0] node53106;
	wire [4-1:0] node53109;
	wire [4-1:0] node53110;
	wire [4-1:0] node53111;
	wire [4-1:0] node53115;
	wire [4-1:0] node53116;
	wire [4-1:0] node53120;
	wire [4-1:0] node53121;
	wire [4-1:0] node53123;
	wire [4-1:0] node53124;
	wire [4-1:0] node53125;
	wire [4-1:0] node53128;
	wire [4-1:0] node53131;
	wire [4-1:0] node53133;
	wire [4-1:0] node53136;
	wire [4-1:0] node53137;
	wire [4-1:0] node53138;
	wire [4-1:0] node53139;
	wire [4-1:0] node53142;
	wire [4-1:0] node53146;
	wire [4-1:0] node53147;
	wire [4-1:0] node53151;
	wire [4-1:0] node53152;
	wire [4-1:0] node53153;
	wire [4-1:0] node53154;
	wire [4-1:0] node53156;
	wire [4-1:0] node53159;
	wire [4-1:0] node53160;
	wire [4-1:0] node53164;
	wire [4-1:0] node53165;
	wire [4-1:0] node53167;
	wire [4-1:0] node53170;
	wire [4-1:0] node53171;
	wire [4-1:0] node53172;
	wire [4-1:0] node53175;
	wire [4-1:0] node53178;
	wire [4-1:0] node53179;
	wire [4-1:0] node53182;
	wire [4-1:0] node53185;
	wire [4-1:0] node53186;
	wire [4-1:0] node53187;
	wire [4-1:0] node53188;
	wire [4-1:0] node53191;
	wire [4-1:0] node53194;
	wire [4-1:0] node53196;
	wire [4-1:0] node53198;
	wire [4-1:0] node53201;
	wire [4-1:0] node53202;
	wire [4-1:0] node53203;
	wire [4-1:0] node53207;
	wire [4-1:0] node53208;
	wire [4-1:0] node53210;
	wire [4-1:0] node53213;
	wire [4-1:0] node53215;
	wire [4-1:0] node53218;
	wire [4-1:0] node53219;
	wire [4-1:0] node53220;
	wire [4-1:0] node53221;
	wire [4-1:0] node53222;
	wire [4-1:0] node53223;
	wire [4-1:0] node53224;
	wire [4-1:0] node53228;
	wire [4-1:0] node53229;
	wire [4-1:0] node53232;
	wire [4-1:0] node53235;
	wire [4-1:0] node53236;
	wire [4-1:0] node53240;
	wire [4-1:0] node53241;
	wire [4-1:0] node53242;
	wire [4-1:0] node53245;
	wire [4-1:0] node53249;
	wire [4-1:0] node53250;
	wire [4-1:0] node53251;
	wire [4-1:0] node53252;
	wire [4-1:0] node53254;
	wire [4-1:0] node53259;
	wire [4-1:0] node53260;
	wire [4-1:0] node53263;
	wire [4-1:0] node53266;
	wire [4-1:0] node53267;
	wire [4-1:0] node53268;
	wire [4-1:0] node53270;
	wire [4-1:0] node53272;
	wire [4-1:0] node53275;
	wire [4-1:0] node53276;
	wire [4-1:0] node53277;
	wire [4-1:0] node53280;
	wire [4-1:0] node53283;
	wire [4-1:0] node53285;
	wire [4-1:0] node53286;
	wire [4-1:0] node53289;
	wire [4-1:0] node53292;
	wire [4-1:0] node53293;
	wire [4-1:0] node53294;
	wire [4-1:0] node53295;
	wire [4-1:0] node53298;
	wire [4-1:0] node53301;
	wire [4-1:0] node53302;
	wire [4-1:0] node53306;
	wire [4-1:0] node53307;
	wire [4-1:0] node53309;
	wire [4-1:0] node53312;
	wire [4-1:0] node53313;
	wire [4-1:0] node53317;
	wire [4-1:0] node53318;
	wire [4-1:0] node53319;
	wire [4-1:0] node53320;
	wire [4-1:0] node53321;
	wire [4-1:0] node53322;
	wire [4-1:0] node53323;
	wire [4-1:0] node53327;
	wire [4-1:0] node53328;
	wire [4-1:0] node53332;
	wire [4-1:0] node53333;
	wire [4-1:0] node53334;
	wire [4-1:0] node53339;
	wire [4-1:0] node53340;
	wire [4-1:0] node53341;
	wire [4-1:0] node53345;
	wire [4-1:0] node53346;
	wire [4-1:0] node53350;
	wire [4-1:0] node53351;
	wire [4-1:0] node53352;
	wire [4-1:0] node53354;
	wire [4-1:0] node53355;
	wire [4-1:0] node53359;
	wire [4-1:0] node53360;
	wire [4-1:0] node53361;
	wire [4-1:0] node53365;
	wire [4-1:0] node53366;
	wire [4-1:0] node53370;
	wire [4-1:0] node53371;
	wire [4-1:0] node53372;
	wire [4-1:0] node53374;
	wire [4-1:0] node53377;
	wire [4-1:0] node53378;
	wire [4-1:0] node53381;
	wire [4-1:0] node53384;
	wire [4-1:0] node53386;
	wire [4-1:0] node53387;
	wire [4-1:0] node53388;
	wire [4-1:0] node53392;
	wire [4-1:0] node53393;
	wire [4-1:0] node53397;
	wire [4-1:0] node53398;
	wire [4-1:0] node53399;
	wire [4-1:0] node53400;
	wire [4-1:0] node53401;
	wire [4-1:0] node53402;
	wire [4-1:0] node53406;
	wire [4-1:0] node53409;
	wire [4-1:0] node53410;
	wire [4-1:0] node53411;
	wire [4-1:0] node53415;
	wire [4-1:0] node53416;
	wire [4-1:0] node53420;
	wire [4-1:0] node53421;
	wire [4-1:0] node53422;
	wire [4-1:0] node53424;
	wire [4-1:0] node53426;
	wire [4-1:0] node53429;
	wire [4-1:0] node53431;
	wire [4-1:0] node53434;
	wire [4-1:0] node53435;
	wire [4-1:0] node53436;
	wire [4-1:0] node53437;
	wire [4-1:0] node53441;
	wire [4-1:0] node53442;
	wire [4-1:0] node53445;
	wire [4-1:0] node53448;
	wire [4-1:0] node53449;
	wire [4-1:0] node53452;
	wire [4-1:0] node53455;
	wire [4-1:0] node53456;
	wire [4-1:0] node53457;
	wire [4-1:0] node53458;
	wire [4-1:0] node53459;
	wire [4-1:0] node53463;
	wire [4-1:0] node53464;
	wire [4-1:0] node53468;
	wire [4-1:0] node53469;
	wire [4-1:0] node53470;
	wire [4-1:0] node53471;
	wire [4-1:0] node53476;
	wire [4-1:0] node53477;
	wire [4-1:0] node53481;
	wire [4-1:0] node53482;
	wire [4-1:0] node53483;
	wire [4-1:0] node53484;
	wire [4-1:0] node53488;
	wire [4-1:0] node53489;
	wire [4-1:0] node53493;
	wire [4-1:0] node53494;
	wire [4-1:0] node53495;
	wire [4-1:0] node53499;
	wire [4-1:0] node53500;
	wire [4-1:0] node53504;
	wire [4-1:0] node53505;
	wire [4-1:0] node53506;
	wire [4-1:0] node53507;
	wire [4-1:0] node53508;
	wire [4-1:0] node53509;
	wire [4-1:0] node53510;
	wire [4-1:0] node53511;
	wire [4-1:0] node53512;
	wire [4-1:0] node53516;
	wire [4-1:0] node53517;
	wire [4-1:0] node53521;
	wire [4-1:0] node53523;
	wire [4-1:0] node53526;
	wire [4-1:0] node53527;
	wire [4-1:0] node53528;
	wire [4-1:0] node53530;
	wire [4-1:0] node53533;
	wire [4-1:0] node53534;
	wire [4-1:0] node53537;
	wire [4-1:0] node53540;
	wire [4-1:0] node53541;
	wire [4-1:0] node53542;
	wire [4-1:0] node53545;
	wire [4-1:0] node53548;
	wire [4-1:0] node53549;
	wire [4-1:0] node53552;
	wire [4-1:0] node53555;
	wire [4-1:0] node53556;
	wire [4-1:0] node53557;
	wire [4-1:0] node53558;
	wire [4-1:0] node53559;
	wire [4-1:0] node53563;
	wire [4-1:0] node53566;
	wire [4-1:0] node53567;
	wire [4-1:0] node53570;
	wire [4-1:0] node53573;
	wire [4-1:0] node53574;
	wire [4-1:0] node53575;
	wire [4-1:0] node53576;
	wire [4-1:0] node53579;
	wire [4-1:0] node53582;
	wire [4-1:0] node53583;
	wire [4-1:0] node53586;
	wire [4-1:0] node53589;
	wire [4-1:0] node53590;
	wire [4-1:0] node53591;
	wire [4-1:0] node53594;
	wire [4-1:0] node53598;
	wire [4-1:0] node53599;
	wire [4-1:0] node53600;
	wire [4-1:0] node53601;
	wire [4-1:0] node53602;
	wire [4-1:0] node53603;
	wire [4-1:0] node53606;
	wire [4-1:0] node53609;
	wire [4-1:0] node53611;
	wire [4-1:0] node53614;
	wire [4-1:0] node53615;
	wire [4-1:0] node53617;
	wire [4-1:0] node53620;
	wire [4-1:0] node53621;
	wire [4-1:0] node53625;
	wire [4-1:0] node53626;
	wire [4-1:0] node53627;
	wire [4-1:0] node53628;
	wire [4-1:0] node53631;
	wire [4-1:0] node53634;
	wire [4-1:0] node53636;
	wire [4-1:0] node53639;
	wire [4-1:0] node53641;
	wire [4-1:0] node53642;
	wire [4-1:0] node53645;
	wire [4-1:0] node53648;
	wire [4-1:0] node53649;
	wire [4-1:0] node53650;
	wire [4-1:0] node53651;
	wire [4-1:0] node53654;
	wire [4-1:0] node53657;
	wire [4-1:0] node53658;
	wire [4-1:0] node53660;
	wire [4-1:0] node53664;
	wire [4-1:0] node53665;
	wire [4-1:0] node53666;
	wire [4-1:0] node53667;
	wire [4-1:0] node53671;
	wire [4-1:0] node53674;
	wire [4-1:0] node53675;
	wire [4-1:0] node53678;
	wire [4-1:0] node53681;
	wire [4-1:0] node53682;
	wire [4-1:0] node53683;
	wire [4-1:0] node53684;
	wire [4-1:0] node53685;
	wire [4-1:0] node53686;
	wire [4-1:0] node53689;
	wire [4-1:0] node53692;
	wire [4-1:0] node53693;
	wire [4-1:0] node53694;
	wire [4-1:0] node53698;
	wire [4-1:0] node53699;
	wire [4-1:0] node53703;
	wire [4-1:0] node53704;
	wire [4-1:0] node53706;
	wire [4-1:0] node53709;
	wire [4-1:0] node53710;
	wire [4-1:0] node53713;
	wire [4-1:0] node53716;
	wire [4-1:0] node53717;
	wire [4-1:0] node53718;
	wire [4-1:0] node53719;
	wire [4-1:0] node53720;
	wire [4-1:0] node53725;
	wire [4-1:0] node53727;
	wire [4-1:0] node53730;
	wire [4-1:0] node53731;
	wire [4-1:0] node53732;
	wire [4-1:0] node53733;
	wire [4-1:0] node53736;
	wire [4-1:0] node53739;
	wire [4-1:0] node53741;
	wire [4-1:0] node53744;
	wire [4-1:0] node53745;
	wire [4-1:0] node53749;
	wire [4-1:0] node53750;
	wire [4-1:0] node53751;
	wire [4-1:0] node53752;
	wire [4-1:0] node53754;
	wire [4-1:0] node53755;
	wire [4-1:0] node53759;
	wire [4-1:0] node53760;
	wire [4-1:0] node53761;
	wire [4-1:0] node53765;
	wire [4-1:0] node53766;
	wire [4-1:0] node53770;
	wire [4-1:0] node53771;
	wire [4-1:0] node53772;
	wire [4-1:0] node53776;
	wire [4-1:0] node53777;
	wire [4-1:0] node53778;
	wire [4-1:0] node53782;
	wire [4-1:0] node53785;
	wire [4-1:0] node53786;
	wire [4-1:0] node53787;
	wire [4-1:0] node53789;
	wire [4-1:0] node53790;
	wire [4-1:0] node53795;
	wire [4-1:0] node53796;
	wire [4-1:0] node53797;
	wire [4-1:0] node53798;
	wire [4-1:0] node53802;
	wire [4-1:0] node53803;
	wire [4-1:0] node53807;
	wire [4-1:0] node53808;
	wire [4-1:0] node53809;
	wire [4-1:0] node53814;
	wire [4-1:0] node53815;
	wire [4-1:0] node53816;
	wire [4-1:0] node53817;
	wire [4-1:0] node53818;
	wire [4-1:0] node53819;
	wire [4-1:0] node53820;
	wire [4-1:0] node53821;
	wire [4-1:0] node53824;
	wire [4-1:0] node53827;
	wire [4-1:0] node53828;
	wire [4-1:0] node53831;
	wire [4-1:0] node53834;
	wire [4-1:0] node53835;
	wire [4-1:0] node53839;
	wire [4-1:0] node53840;
	wire [4-1:0] node53841;
	wire [4-1:0] node53842;
	wire [4-1:0] node53845;
	wire [4-1:0] node53849;
	wire [4-1:0] node53850;
	wire [4-1:0] node53851;
	wire [4-1:0] node53855;
	wire [4-1:0] node53856;
	wire [4-1:0] node53859;
	wire [4-1:0] node53862;
	wire [4-1:0] node53863;
	wire [4-1:0] node53864;
	wire [4-1:0] node53865;
	wire [4-1:0] node53868;
	wire [4-1:0] node53871;
	wire [4-1:0] node53872;
	wire [4-1:0] node53873;
	wire [4-1:0] node53877;
	wire [4-1:0] node53880;
	wire [4-1:0] node53881;
	wire [4-1:0] node53882;
	wire [4-1:0] node53884;
	wire [4-1:0] node53888;
	wire [4-1:0] node53889;
	wire [4-1:0] node53891;
	wire [4-1:0] node53894;
	wire [4-1:0] node53895;
	wire [4-1:0] node53898;
	wire [4-1:0] node53901;
	wire [4-1:0] node53902;
	wire [4-1:0] node53903;
	wire [4-1:0] node53904;
	wire [4-1:0] node53905;
	wire [4-1:0] node53906;
	wire [4-1:0] node53909;
	wire [4-1:0] node53913;
	wire [4-1:0] node53914;
	wire [4-1:0] node53915;
	wire [4-1:0] node53920;
	wire [4-1:0] node53921;
	wire [4-1:0] node53922;
	wire [4-1:0] node53923;
	wire [4-1:0] node53928;
	wire [4-1:0] node53929;
	wire [4-1:0] node53930;
	wire [4-1:0] node53933;
	wire [4-1:0] node53936;
	wire [4-1:0] node53937;
	wire [4-1:0] node53940;
	wire [4-1:0] node53943;
	wire [4-1:0] node53944;
	wire [4-1:0] node53945;
	wire [4-1:0] node53946;
	wire [4-1:0] node53948;
	wire [4-1:0] node53952;
	wire [4-1:0] node53953;
	wire [4-1:0] node53955;
	wire [4-1:0] node53958;
	wire [4-1:0] node53960;
	wire [4-1:0] node53963;
	wire [4-1:0] node53964;
	wire [4-1:0] node53966;
	wire [4-1:0] node53969;
	wire [4-1:0] node53971;
	wire [4-1:0] node53974;
	wire [4-1:0] node53975;
	wire [4-1:0] node53976;
	wire [4-1:0] node53977;
	wire [4-1:0] node53978;
	wire [4-1:0] node53979;
	wire [4-1:0] node53981;
	wire [4-1:0] node53984;
	wire [4-1:0] node53987;
	wire [4-1:0] node53988;
	wire [4-1:0] node53989;
	wire [4-1:0] node53993;
	wire [4-1:0] node53996;
	wire [4-1:0] node53997;
	wire [4-1:0] node53998;
	wire [4-1:0] node54001;
	wire [4-1:0] node54004;
	wire [4-1:0] node54005;
	wire [4-1:0] node54006;
	wire [4-1:0] node54010;
	wire [4-1:0] node54013;
	wire [4-1:0] node54014;
	wire [4-1:0] node54015;
	wire [4-1:0] node54016;
	wire [4-1:0] node54019;
	wire [4-1:0] node54022;
	wire [4-1:0] node54024;
	wire [4-1:0] node54027;
	wire [4-1:0] node54028;
	wire [4-1:0] node54029;
	wire [4-1:0] node54032;
	wire [4-1:0] node54035;
	wire [4-1:0] node54036;
	wire [4-1:0] node54037;
	wire [4-1:0] node54041;
	wire [4-1:0] node54044;
	wire [4-1:0] node54045;
	wire [4-1:0] node54046;
	wire [4-1:0] node54047;
	wire [4-1:0] node54048;
	wire [4-1:0] node54049;
	wire [4-1:0] node54053;
	wire [4-1:0] node54056;
	wire [4-1:0] node54057;
	wire [4-1:0] node54061;
	wire [4-1:0] node54062;
	wire [4-1:0] node54063;
	wire [4-1:0] node54066;
	wire [4-1:0] node54069;
	wire [4-1:0] node54070;
	wire [4-1:0] node54072;
	wire [4-1:0] node54075;
	wire [4-1:0] node54078;
	wire [4-1:0] node54079;
	wire [4-1:0] node54080;
	wire [4-1:0] node54081;
	wire [4-1:0] node54082;
	wire [4-1:0] node54086;
	wire [4-1:0] node54089;
	wire [4-1:0] node54090;
	wire [4-1:0] node54091;
	wire [4-1:0] node54094;
	wire [4-1:0] node54098;
	wire [4-1:0] node54099;
	wire [4-1:0] node54100;
	wire [4-1:0] node54103;
	wire [4-1:0] node54106;
	wire [4-1:0] node54107;
	wire [4-1:0] node54110;
	wire [4-1:0] node54113;
	wire [4-1:0] node54114;
	wire [4-1:0] node54115;
	wire [4-1:0] node54116;
	wire [4-1:0] node54117;
	wire [4-1:0] node54118;
	wire [4-1:0] node54119;
	wire [4-1:0] node54120;
	wire [4-1:0] node54121;
	wire [4-1:0] node54122;
	wire [4-1:0] node54123;
	wire [4-1:0] node54124;
	wire [4-1:0] node54128;
	wire [4-1:0] node54129;
	wire [4-1:0] node54132;
	wire [4-1:0] node54135;
	wire [4-1:0] node54136;
	wire [4-1:0] node54137;
	wire [4-1:0] node54140;
	wire [4-1:0] node54144;
	wire [4-1:0] node54145;
	wire [4-1:0] node54146;
	wire [4-1:0] node54147;
	wire [4-1:0] node54150;
	wire [4-1:0] node54154;
	wire [4-1:0] node54155;
	wire [4-1:0] node54156;
	wire [4-1:0] node54159;
	wire [4-1:0] node54162;
	wire [4-1:0] node54163;
	wire [4-1:0] node54166;
	wire [4-1:0] node54169;
	wire [4-1:0] node54170;
	wire [4-1:0] node54171;
	wire [4-1:0] node54172;
	wire [4-1:0] node54175;
	wire [4-1:0] node54178;
	wire [4-1:0] node54179;
	wire [4-1:0] node54180;
	wire [4-1:0] node54184;
	wire [4-1:0] node54185;
	wire [4-1:0] node54188;
	wire [4-1:0] node54191;
	wire [4-1:0] node54192;
	wire [4-1:0] node54193;
	wire [4-1:0] node54194;
	wire [4-1:0] node54197;
	wire [4-1:0] node54200;
	wire [4-1:0] node54203;
	wire [4-1:0] node54204;
	wire [4-1:0] node54207;
	wire [4-1:0] node54209;
	wire [4-1:0] node54212;
	wire [4-1:0] node54213;
	wire [4-1:0] node54214;
	wire [4-1:0] node54215;
	wire [4-1:0] node54217;
	wire [4-1:0] node54220;
	wire [4-1:0] node54222;
	wire [4-1:0] node54225;
	wire [4-1:0] node54226;
	wire [4-1:0] node54227;
	wire [4-1:0] node54230;
	wire [4-1:0] node54233;
	wire [4-1:0] node54234;
	wire [4-1:0] node54237;
	wire [4-1:0] node54240;
	wire [4-1:0] node54241;
	wire [4-1:0] node54242;
	wire [4-1:0] node54243;
	wire [4-1:0] node54246;
	wire [4-1:0] node54249;
	wire [4-1:0] node54250;
	wire [4-1:0] node54253;
	wire [4-1:0] node54256;
	wire [4-1:0] node54257;
	wire [4-1:0] node54258;
	wire [4-1:0] node54261;
	wire [4-1:0] node54264;
	wire [4-1:0] node54265;
	wire [4-1:0] node54269;
	wire [4-1:0] node54270;
	wire [4-1:0] node54271;
	wire [4-1:0] node54272;
	wire [4-1:0] node54273;
	wire [4-1:0] node54274;
	wire [4-1:0] node54277;
	wire [4-1:0] node54278;
	wire [4-1:0] node54282;
	wire [4-1:0] node54285;
	wire [4-1:0] node54286;
	wire [4-1:0] node54287;
	wire [4-1:0] node54289;
	wire [4-1:0] node54292;
	wire [4-1:0] node54294;
	wire [4-1:0] node54297;
	wire [4-1:0] node54300;
	wire [4-1:0] node54301;
	wire [4-1:0] node54302;
	wire [4-1:0] node54303;
	wire [4-1:0] node54305;
	wire [4-1:0] node54309;
	wire [4-1:0] node54311;
	wire [4-1:0] node54314;
	wire [4-1:0] node54315;
	wire [4-1:0] node54316;
	wire [4-1:0] node54317;
	wire [4-1:0] node54321;
	wire [4-1:0] node54322;
	wire [4-1:0] node54326;
	wire [4-1:0] node54327;
	wire [4-1:0] node54328;
	wire [4-1:0] node54332;
	wire [4-1:0] node54335;
	wire [4-1:0] node54336;
	wire [4-1:0] node54337;
	wire [4-1:0] node54338;
	wire [4-1:0] node54340;
	wire [4-1:0] node54343;
	wire [4-1:0] node54344;
	wire [4-1:0] node54347;
	wire [4-1:0] node54348;
	wire [4-1:0] node54352;
	wire [4-1:0] node54353;
	wire [4-1:0] node54354;
	wire [4-1:0] node54356;
	wire [4-1:0] node54359;
	wire [4-1:0] node54361;
	wire [4-1:0] node54364;
	wire [4-1:0] node54365;
	wire [4-1:0] node54367;
	wire [4-1:0] node54370;
	wire [4-1:0] node54372;
	wire [4-1:0] node54375;
	wire [4-1:0] node54376;
	wire [4-1:0] node54377;
	wire [4-1:0] node54378;
	wire [4-1:0] node54379;
	wire [4-1:0] node54383;
	wire [4-1:0] node54386;
	wire [4-1:0] node54387;
	wire [4-1:0] node54388;
	wire [4-1:0] node54392;
	wire [4-1:0] node54393;
	wire [4-1:0] node54397;
	wire [4-1:0] node54398;
	wire [4-1:0] node54401;
	wire [4-1:0] node54403;
	wire [4-1:0] node54404;
	wire [4-1:0] node54407;
	wire [4-1:0] node54410;
	wire [4-1:0] node54411;
	wire [4-1:0] node54412;
	wire [4-1:0] node54413;
	wire [4-1:0] node54414;
	wire [4-1:0] node54415;
	wire [4-1:0] node54416;
	wire [4-1:0] node54418;
	wire [4-1:0] node54421;
	wire [4-1:0] node54423;
	wire [4-1:0] node54426;
	wire [4-1:0] node54427;
	wire [4-1:0] node54429;
	wire [4-1:0] node54432;
	wire [4-1:0] node54434;
	wire [4-1:0] node54437;
	wire [4-1:0] node54438;
	wire [4-1:0] node54439;
	wire [4-1:0] node54443;
	wire [4-1:0] node54445;
	wire [4-1:0] node54447;
	wire [4-1:0] node54450;
	wire [4-1:0] node54451;
	wire [4-1:0] node54452;
	wire [4-1:0] node54455;
	wire [4-1:0] node54456;
	wire [4-1:0] node54459;
	wire [4-1:0] node54462;
	wire [4-1:0] node54463;
	wire [4-1:0] node54465;
	wire [4-1:0] node54468;
	wire [4-1:0] node54470;
	wire [4-1:0] node54473;
	wire [4-1:0] node54474;
	wire [4-1:0] node54475;
	wire [4-1:0] node54476;
	wire [4-1:0] node54478;
	wire [4-1:0] node54481;
	wire [4-1:0] node54482;
	wire [4-1:0] node54485;
	wire [4-1:0] node54487;
	wire [4-1:0] node54490;
	wire [4-1:0] node54491;
	wire [4-1:0] node54492;
	wire [4-1:0] node54493;
	wire [4-1:0] node54497;
	wire [4-1:0] node54500;
	wire [4-1:0] node54502;
	wire [4-1:0] node54505;
	wire [4-1:0] node54506;
	wire [4-1:0] node54507;
	wire [4-1:0] node54508;
	wire [4-1:0] node54512;
	wire [4-1:0] node54513;
	wire [4-1:0] node54517;
	wire [4-1:0] node54518;
	wire [4-1:0] node54519;
	wire [4-1:0] node54523;
	wire [4-1:0] node54524;
	wire [4-1:0] node54528;
	wire [4-1:0] node54529;
	wire [4-1:0] node54530;
	wire [4-1:0] node54531;
	wire [4-1:0] node54532;
	wire [4-1:0] node54534;
	wire [4-1:0] node54537;
	wire [4-1:0] node54538;
	wire [4-1:0] node54539;
	wire [4-1:0] node54542;
	wire [4-1:0] node54545;
	wire [4-1:0] node54546;
	wire [4-1:0] node54549;
	wire [4-1:0] node54552;
	wire [4-1:0] node54553;
	wire [4-1:0] node54556;
	wire [4-1:0] node54557;
	wire [4-1:0] node54560;
	wire [4-1:0] node54563;
	wire [4-1:0] node54564;
	wire [4-1:0] node54565;
	wire [4-1:0] node54568;
	wire [4-1:0] node54569;
	wire [4-1:0] node54573;
	wire [4-1:0] node54574;
	wire [4-1:0] node54575;
	wire [4-1:0] node54580;
	wire [4-1:0] node54581;
	wire [4-1:0] node54582;
	wire [4-1:0] node54583;
	wire [4-1:0] node54585;
	wire [4-1:0] node54588;
	wire [4-1:0] node54589;
	wire [4-1:0] node54590;
	wire [4-1:0] node54594;
	wire [4-1:0] node54595;
	wire [4-1:0] node54599;
	wire [4-1:0] node54600;
	wire [4-1:0] node54601;
	wire [4-1:0] node54603;
	wire [4-1:0] node54607;
	wire [4-1:0] node54608;
	wire [4-1:0] node54612;
	wire [4-1:0] node54613;
	wire [4-1:0] node54614;
	wire [4-1:0] node54615;
	wire [4-1:0] node54616;
	wire [4-1:0] node54619;
	wire [4-1:0] node54622;
	wire [4-1:0] node54623;
	wire [4-1:0] node54627;
	wire [4-1:0] node54628;
	wire [4-1:0] node54631;
	wire [4-1:0] node54634;
	wire [4-1:0] node54635;
	wire [4-1:0] node54638;
	wire [4-1:0] node54641;
	wire [4-1:0] node54642;
	wire [4-1:0] node54643;
	wire [4-1:0] node54644;
	wire [4-1:0] node54645;
	wire [4-1:0] node54646;
	wire [4-1:0] node54647;
	wire [4-1:0] node54648;
	wire [4-1:0] node54651;
	wire [4-1:0] node54652;
	wire [4-1:0] node54655;
	wire [4-1:0] node54658;
	wire [4-1:0] node54659;
	wire [4-1:0] node54660;
	wire [4-1:0] node54663;
	wire [4-1:0] node54666;
	wire [4-1:0] node54667;
	wire [4-1:0] node54670;
	wire [4-1:0] node54673;
	wire [4-1:0] node54674;
	wire [4-1:0] node54676;
	wire [4-1:0] node54677;
	wire [4-1:0] node54681;
	wire [4-1:0] node54682;
	wire [4-1:0] node54683;
	wire [4-1:0] node54687;
	wire [4-1:0] node54688;
	wire [4-1:0] node54692;
	wire [4-1:0] node54693;
	wire [4-1:0] node54694;
	wire [4-1:0] node54695;
	wire [4-1:0] node54698;
	wire [4-1:0] node54701;
	wire [4-1:0] node54702;
	wire [4-1:0] node54705;
	wire [4-1:0] node54708;
	wire [4-1:0] node54709;
	wire [4-1:0] node54710;
	wire [4-1:0] node54713;
	wire [4-1:0] node54716;
	wire [4-1:0] node54717;
	wire [4-1:0] node54718;
	wire [4-1:0] node54722;
	wire [4-1:0] node54723;
	wire [4-1:0] node54726;
	wire [4-1:0] node54729;
	wire [4-1:0] node54730;
	wire [4-1:0] node54731;
	wire [4-1:0] node54732;
	wire [4-1:0] node54735;
	wire [4-1:0] node54738;
	wire [4-1:0] node54739;
	wire [4-1:0] node54740;
	wire [4-1:0] node54743;
	wire [4-1:0] node54746;
	wire [4-1:0] node54748;
	wire [4-1:0] node54749;
	wire [4-1:0] node54753;
	wire [4-1:0] node54754;
	wire [4-1:0] node54755;
	wire [4-1:0] node54756;
	wire [4-1:0] node54757;
	wire [4-1:0] node54760;
	wire [4-1:0] node54763;
	wire [4-1:0] node54765;
	wire [4-1:0] node54768;
	wire [4-1:0] node54770;
	wire [4-1:0] node54773;
	wire [4-1:0] node54774;
	wire [4-1:0] node54775;
	wire [4-1:0] node54778;
	wire [4-1:0] node54779;
	wire [4-1:0] node54783;
	wire [4-1:0] node54784;
	wire [4-1:0] node54787;
	wire [4-1:0] node54790;
	wire [4-1:0] node54791;
	wire [4-1:0] node54792;
	wire [4-1:0] node54793;
	wire [4-1:0] node54794;
	wire [4-1:0] node54795;
	wire [4-1:0] node54796;
	wire [4-1:0] node54800;
	wire [4-1:0] node54803;
	wire [4-1:0] node54804;
	wire [4-1:0] node54808;
	wire [4-1:0] node54809;
	wire [4-1:0] node54810;
	wire [4-1:0] node54811;
	wire [4-1:0] node54814;
	wire [4-1:0] node54817;
	wire [4-1:0] node54818;
	wire [4-1:0] node54821;
	wire [4-1:0] node54824;
	wire [4-1:0] node54825;
	wire [4-1:0] node54826;
	wire [4-1:0] node54829;
	wire [4-1:0] node54832;
	wire [4-1:0] node54833;
	wire [4-1:0] node54837;
	wire [4-1:0] node54838;
	wire [4-1:0] node54839;
	wire [4-1:0] node54840;
	wire [4-1:0] node54841;
	wire [4-1:0] node54844;
	wire [4-1:0] node54847;
	wire [4-1:0] node54849;
	wire [4-1:0] node54852;
	wire [4-1:0] node54854;
	wire [4-1:0] node54857;
	wire [4-1:0] node54858;
	wire [4-1:0] node54859;
	wire [4-1:0] node54862;
	wire [4-1:0] node54865;
	wire [4-1:0] node54867;
	wire [4-1:0] node54869;
	wire [4-1:0] node54872;
	wire [4-1:0] node54873;
	wire [4-1:0] node54874;
	wire [4-1:0] node54875;
	wire [4-1:0] node54877;
	wire [4-1:0] node54878;
	wire [4-1:0] node54881;
	wire [4-1:0] node54884;
	wire [4-1:0] node54885;
	wire [4-1:0] node54888;
	wire [4-1:0] node54890;
	wire [4-1:0] node54893;
	wire [4-1:0] node54894;
	wire [4-1:0] node54895;
	wire [4-1:0] node54896;
	wire [4-1:0] node54899;
	wire [4-1:0] node54902;
	wire [4-1:0] node54903;
	wire [4-1:0] node54906;
	wire [4-1:0] node54909;
	wire [4-1:0] node54910;
	wire [4-1:0] node54913;
	wire [4-1:0] node54916;
	wire [4-1:0] node54917;
	wire [4-1:0] node54918;
	wire [4-1:0] node54919;
	wire [4-1:0] node54921;
	wire [4-1:0] node54924;
	wire [4-1:0] node54926;
	wire [4-1:0] node54929;
	wire [4-1:0] node54930;
	wire [4-1:0] node54933;
	wire [4-1:0] node54935;
	wire [4-1:0] node54938;
	wire [4-1:0] node54939;
	wire [4-1:0] node54941;
	wire [4-1:0] node54944;
	wire [4-1:0] node54945;
	wire [4-1:0] node54946;
	wire [4-1:0] node54950;
	wire [4-1:0] node54953;
	wire [4-1:0] node54954;
	wire [4-1:0] node54955;
	wire [4-1:0] node54956;
	wire [4-1:0] node54957;
	wire [4-1:0] node54958;
	wire [4-1:0] node54960;
	wire [4-1:0] node54963;
	wire [4-1:0] node54964;
	wire [4-1:0] node54965;
	wire [4-1:0] node54968;
	wire [4-1:0] node54971;
	wire [4-1:0] node54973;
	wire [4-1:0] node54976;
	wire [4-1:0] node54977;
	wire [4-1:0] node54978;
	wire [4-1:0] node54981;
	wire [4-1:0] node54983;
	wire [4-1:0] node54986;
	wire [4-1:0] node54987;
	wire [4-1:0] node54989;
	wire [4-1:0] node54992;
	wire [4-1:0] node54994;
	wire [4-1:0] node54997;
	wire [4-1:0] node54998;
	wire [4-1:0] node54999;
	wire [4-1:0] node55000;
	wire [4-1:0] node55003;
	wire [4-1:0] node55006;
	wire [4-1:0] node55007;
	wire [4-1:0] node55010;
	wire [4-1:0] node55012;
	wire [4-1:0] node55015;
	wire [4-1:0] node55016;
	wire [4-1:0] node55017;
	wire [4-1:0] node55019;
	wire [4-1:0] node55022;
	wire [4-1:0] node55023;
	wire [4-1:0] node55026;
	wire [4-1:0] node55030;
	wire [4-1:0] node55031;
	wire [4-1:0] node55032;
	wire [4-1:0] node55033;
	wire [4-1:0] node55034;
	wire [4-1:0] node55037;
	wire [4-1:0] node55038;
	wire [4-1:0] node55042;
	wire [4-1:0] node55043;
	wire [4-1:0] node55045;
	wire [4-1:0] node55048;
	wire [4-1:0] node55049;
	wire [4-1:0] node55052;
	wire [4-1:0] node55055;
	wire [4-1:0] node55056;
	wire [4-1:0] node55059;
	wire [4-1:0] node55060;
	wire [4-1:0] node55063;
	wire [4-1:0] node55066;
	wire [4-1:0] node55067;
	wire [4-1:0] node55068;
	wire [4-1:0] node55069;
	wire [4-1:0] node55071;
	wire [4-1:0] node55074;
	wire [4-1:0] node55077;
	wire [4-1:0] node55078;
	wire [4-1:0] node55081;
	wire [4-1:0] node55082;
	wire [4-1:0] node55085;
	wire [4-1:0] node55088;
	wire [4-1:0] node55089;
	wire [4-1:0] node55091;
	wire [4-1:0] node55094;
	wire [4-1:0] node55095;
	wire [4-1:0] node55096;
	wire [4-1:0] node55100;
	wire [4-1:0] node55101;
	wire [4-1:0] node55104;
	wire [4-1:0] node55107;
	wire [4-1:0] node55108;
	wire [4-1:0] node55109;
	wire [4-1:0] node55110;
	wire [4-1:0] node55111;
	wire [4-1:0] node55112;
	wire [4-1:0] node55116;
	wire [4-1:0] node55117;
	wire [4-1:0] node55120;
	wire [4-1:0] node55123;
	wire [4-1:0] node55124;
	wire [4-1:0] node55125;
	wire [4-1:0] node55129;
	wire [4-1:0] node55132;
	wire [4-1:0] node55133;
	wire [4-1:0] node55134;
	wire [4-1:0] node55135;
	wire [4-1:0] node55138;
	wire [4-1:0] node55141;
	wire [4-1:0] node55142;
	wire [4-1:0] node55145;
	wire [4-1:0] node55148;
	wire [4-1:0] node55149;
	wire [4-1:0] node55150;
	wire [4-1:0] node55154;
	wire [4-1:0] node55157;
	wire [4-1:0] node55158;
	wire [4-1:0] node55159;
	wire [4-1:0] node55160;
	wire [4-1:0] node55161;
	wire [4-1:0] node55164;
	wire [4-1:0] node55167;
	wire [4-1:0] node55169;
	wire [4-1:0] node55172;
	wire [4-1:0] node55173;
	wire [4-1:0] node55174;
	wire [4-1:0] node55178;
	wire [4-1:0] node55181;
	wire [4-1:0] node55182;
	wire [4-1:0] node55183;
	wire [4-1:0] node55185;
	wire [4-1:0] node55186;
	wire [4-1:0] node55190;
	wire [4-1:0] node55192;
	wire [4-1:0] node55195;
	wire [4-1:0] node55196;
	wire [4-1:0] node55197;
	wire [4-1:0] node55200;
	wire [4-1:0] node55203;
	wire [4-1:0] node55204;
	wire [4-1:0] node55207;
	wire [4-1:0] node55210;
	wire [4-1:0] node55211;
	wire [4-1:0] node55212;
	wire [4-1:0] node55213;
	wire [4-1:0] node55214;
	wire [4-1:0] node55215;
	wire [4-1:0] node55216;
	wire [4-1:0] node55217;
	wire [4-1:0] node55218;
	wire [4-1:0] node55219;
	wire [4-1:0] node55222;
	wire [4-1:0] node55225;
	wire [4-1:0] node55226;
	wire [4-1:0] node55229;
	wire [4-1:0] node55232;
	wire [4-1:0] node55233;
	wire [4-1:0] node55237;
	wire [4-1:0] node55238;
	wire [4-1:0] node55239;
	wire [4-1:0] node55240;
	wire [4-1:0] node55243;
	wire [4-1:0] node55247;
	wire [4-1:0] node55248;
	wire [4-1:0] node55249;
	wire [4-1:0] node55252;
	wire [4-1:0] node55256;
	wire [4-1:0] node55257;
	wire [4-1:0] node55258;
	wire [4-1:0] node55260;
	wire [4-1:0] node55261;
	wire [4-1:0] node55264;
	wire [4-1:0] node55267;
	wire [4-1:0] node55268;
	wire [4-1:0] node55271;
	wire [4-1:0] node55274;
	wire [4-1:0] node55275;
	wire [4-1:0] node55277;
	wire [4-1:0] node55280;
	wire [4-1:0] node55281;
	wire [4-1:0] node55284;
	wire [4-1:0] node55287;
	wire [4-1:0] node55288;
	wire [4-1:0] node55289;
	wire [4-1:0] node55290;
	wire [4-1:0] node55291;
	wire [4-1:0] node55294;
	wire [4-1:0] node55295;
	wire [4-1:0] node55299;
	wire [4-1:0] node55300;
	wire [4-1:0] node55301;
	wire [4-1:0] node55304;
	wire [4-1:0] node55307;
	wire [4-1:0] node55308;
	wire [4-1:0] node55311;
	wire [4-1:0] node55314;
	wire [4-1:0] node55315;
	wire [4-1:0] node55317;
	wire [4-1:0] node55318;
	wire [4-1:0] node55321;
	wire [4-1:0] node55324;
	wire [4-1:0] node55325;
	wire [4-1:0] node55328;
	wire [4-1:0] node55331;
	wire [4-1:0] node55332;
	wire [4-1:0] node55333;
	wire [4-1:0] node55334;
	wire [4-1:0] node55338;
	wire [4-1:0] node55339;
	wire [4-1:0] node55343;
	wire [4-1:0] node55344;
	wire [4-1:0] node55345;
	wire [4-1:0] node55349;
	wire [4-1:0] node55350;
	wire [4-1:0] node55354;
	wire [4-1:0] node55355;
	wire [4-1:0] node55356;
	wire [4-1:0] node55357;
	wire [4-1:0] node55358;
	wire [4-1:0] node55359;
	wire [4-1:0] node55362;
	wire [4-1:0] node55365;
	wire [4-1:0] node55366;
	wire [4-1:0] node55368;
	wire [4-1:0] node55371;
	wire [4-1:0] node55373;
	wire [4-1:0] node55376;
	wire [4-1:0] node55377;
	wire [4-1:0] node55379;
	wire [4-1:0] node55380;
	wire [4-1:0] node55383;
	wire [4-1:0] node55386;
	wire [4-1:0] node55387;
	wire [4-1:0] node55391;
	wire [4-1:0] node55392;
	wire [4-1:0] node55393;
	wire [4-1:0] node55394;
	wire [4-1:0] node55398;
	wire [4-1:0] node55399;
	wire [4-1:0] node55403;
	wire [4-1:0] node55404;
	wire [4-1:0] node55405;
	wire [4-1:0] node55409;
	wire [4-1:0] node55410;
	wire [4-1:0] node55414;
	wire [4-1:0] node55415;
	wire [4-1:0] node55416;
	wire [4-1:0] node55417;
	wire [4-1:0] node55419;
	wire [4-1:0] node55422;
	wire [4-1:0] node55423;
	wire [4-1:0] node55425;
	wire [4-1:0] node55428;
	wire [4-1:0] node55431;
	wire [4-1:0] node55432;
	wire [4-1:0] node55434;
	wire [4-1:0] node55435;
	wire [4-1:0] node55438;
	wire [4-1:0] node55441;
	wire [4-1:0] node55442;
	wire [4-1:0] node55445;
	wire [4-1:0] node55448;
	wire [4-1:0] node55449;
	wire [4-1:0] node55450;
	wire [4-1:0] node55451;
	wire [4-1:0] node55455;
	wire [4-1:0] node55456;
	wire [4-1:0] node55460;
	wire [4-1:0] node55461;
	wire [4-1:0] node55462;
	wire [4-1:0] node55466;
	wire [4-1:0] node55467;
	wire [4-1:0] node55471;
	wire [4-1:0] node55472;
	wire [4-1:0] node55473;
	wire [4-1:0] node55474;
	wire [4-1:0] node55475;
	wire [4-1:0] node55476;
	wire [4-1:0] node55477;
	wire [4-1:0] node55478;
	wire [4-1:0] node55481;
	wire [4-1:0] node55484;
	wire [4-1:0] node55485;
	wire [4-1:0] node55488;
	wire [4-1:0] node55491;
	wire [4-1:0] node55492;
	wire [4-1:0] node55496;
	wire [4-1:0] node55497;
	wire [4-1:0] node55498;
	wire [4-1:0] node55499;
	wire [4-1:0] node55503;
	wire [4-1:0] node55506;
	wire [4-1:0] node55507;
	wire [4-1:0] node55511;
	wire [4-1:0] node55512;
	wire [4-1:0] node55513;
	wire [4-1:0] node55514;
	wire [4-1:0] node55515;
	wire [4-1:0] node55519;
	wire [4-1:0] node55522;
	wire [4-1:0] node55523;
	wire [4-1:0] node55525;
	wire [4-1:0] node55528;
	wire [4-1:0] node55531;
	wire [4-1:0] node55532;
	wire [4-1:0] node55533;
	wire [4-1:0] node55534;
	wire [4-1:0] node55538;
	wire [4-1:0] node55539;
	wire [4-1:0] node55542;
	wire [4-1:0] node55545;
	wire [4-1:0] node55546;
	wire [4-1:0] node55547;
	wire [4-1:0] node55550;
	wire [4-1:0] node55553;
	wire [4-1:0] node55555;
	wire [4-1:0] node55558;
	wire [4-1:0] node55559;
	wire [4-1:0] node55560;
	wire [4-1:0] node55561;
	wire [4-1:0] node55564;
	wire [4-1:0] node55566;
	wire [4-1:0] node55567;
	wire [4-1:0] node55571;
	wire [4-1:0] node55572;
	wire [4-1:0] node55573;
	wire [4-1:0] node55574;
	wire [4-1:0] node55578;
	wire [4-1:0] node55581;
	wire [4-1:0] node55582;
	wire [4-1:0] node55583;
	wire [4-1:0] node55587;
	wire [4-1:0] node55588;
	wire [4-1:0] node55592;
	wire [4-1:0] node55593;
	wire [4-1:0] node55594;
	wire [4-1:0] node55596;
	wire [4-1:0] node55597;
	wire [4-1:0] node55601;
	wire [4-1:0] node55602;
	wire [4-1:0] node55603;
	wire [4-1:0] node55607;
	wire [4-1:0] node55608;
	wire [4-1:0] node55612;
	wire [4-1:0] node55613;
	wire [4-1:0] node55614;
	wire [4-1:0] node55615;
	wire [4-1:0] node55619;
	wire [4-1:0] node55620;
	wire [4-1:0] node55624;
	wire [4-1:0] node55625;
	wire [4-1:0] node55626;
	wire [4-1:0] node55630;
	wire [4-1:0] node55631;
	wire [4-1:0] node55635;
	wire [4-1:0] node55636;
	wire [4-1:0] node55637;
	wire [4-1:0] node55638;
	wire [4-1:0] node55639;
	wire [4-1:0] node55641;
	wire [4-1:0] node55644;
	wire [4-1:0] node55645;
	wire [4-1:0] node55646;
	wire [4-1:0] node55649;
	wire [4-1:0] node55653;
	wire [4-1:0] node55654;
	wire [4-1:0] node55655;
	wire [4-1:0] node55657;
	wire [4-1:0] node55660;
	wire [4-1:0] node55661;
	wire [4-1:0] node55664;
	wire [4-1:0] node55667;
	wire [4-1:0] node55668;
	wire [4-1:0] node55671;
	wire [4-1:0] node55672;
	wire [4-1:0] node55675;
	wire [4-1:0] node55678;
	wire [4-1:0] node55679;
	wire [4-1:0] node55680;
	wire [4-1:0] node55681;
	wire [4-1:0] node55682;
	wire [4-1:0] node55686;
	wire [4-1:0] node55687;
	wire [4-1:0] node55691;
	wire [4-1:0] node55692;
	wire [4-1:0] node55694;
	wire [4-1:0] node55697;
	wire [4-1:0] node55698;
	wire [4-1:0] node55701;
	wire [4-1:0] node55704;
	wire [4-1:0] node55705;
	wire [4-1:0] node55706;
	wire [4-1:0] node55708;
	wire [4-1:0] node55711;
	wire [4-1:0] node55713;
	wire [4-1:0] node55716;
	wire [4-1:0] node55717;
	wire [4-1:0] node55718;
	wire [4-1:0] node55722;
	wire [4-1:0] node55723;
	wire [4-1:0] node55726;
	wire [4-1:0] node55729;
	wire [4-1:0] node55730;
	wire [4-1:0] node55731;
	wire [4-1:0] node55732;
	wire [4-1:0] node55733;
	wire [4-1:0] node55736;
	wire [4-1:0] node55739;
	wire [4-1:0] node55740;
	wire [4-1:0] node55744;
	wire [4-1:0] node55745;
	wire [4-1:0] node55746;
	wire [4-1:0] node55748;
	wire [4-1:0] node55752;
	wire [4-1:0] node55755;
	wire [4-1:0] node55756;
	wire [4-1:0] node55757;
	wire [4-1:0] node55758;
	wire [4-1:0] node55759;
	wire [4-1:0] node55762;
	wire [4-1:0] node55765;
	wire [4-1:0] node55767;
	wire [4-1:0] node55770;
	wire [4-1:0] node55771;
	wire [4-1:0] node55772;
	wire [4-1:0] node55775;
	wire [4-1:0] node55778;
	wire [4-1:0] node55781;
	wire [4-1:0] node55782;
	wire [4-1:0] node55783;
	wire [4-1:0] node55784;
	wire [4-1:0] node55788;
	wire [4-1:0] node55791;
	wire [4-1:0] node55794;
	wire [4-1:0] node55795;
	wire [4-1:0] node55796;
	wire [4-1:0] node55797;
	wire [4-1:0] node55798;
	wire [4-1:0] node55799;
	wire [4-1:0] node55800;
	wire [4-1:0] node55803;
	wire [4-1:0] node55805;
	wire [4-1:0] node55808;
	wire [4-1:0] node55809;
	wire [4-1:0] node55812;
	wire [4-1:0] node55814;
	wire [4-1:0] node55817;
	wire [4-1:0] node55818;
	wire [4-1:0] node55819;
	wire [4-1:0] node55821;
	wire [4-1:0] node55824;
	wire [4-1:0] node55825;
	wire [4-1:0] node55828;
	wire [4-1:0] node55831;
	wire [4-1:0] node55832;
	wire [4-1:0] node55833;
	wire [4-1:0] node55835;
	wire [4-1:0] node55838;
	wire [4-1:0] node55839;
	wire [4-1:0] node55842;
	wire [4-1:0] node55845;
	wire [4-1:0] node55848;
	wire [4-1:0] node55849;
	wire [4-1:0] node55850;
	wire [4-1:0] node55851;
	wire [4-1:0] node55852;
	wire [4-1:0] node55856;
	wire [4-1:0] node55857;
	wire [4-1:0] node55858;
	wire [4-1:0] node55861;
	wire [4-1:0] node55864;
	wire [4-1:0] node55866;
	wire [4-1:0] node55869;
	wire [4-1:0] node55870;
	wire [4-1:0] node55871;
	wire [4-1:0] node55874;
	wire [4-1:0] node55877;
	wire [4-1:0] node55878;
	wire [4-1:0] node55882;
	wire [4-1:0] node55883;
	wire [4-1:0] node55884;
	wire [4-1:0] node55885;
	wire [4-1:0] node55887;
	wire [4-1:0] node55890;
	wire [4-1:0] node55891;
	wire [4-1:0] node55894;
	wire [4-1:0] node55897;
	wire [4-1:0] node55899;
	wire [4-1:0] node55902;
	wire [4-1:0] node55903;
	wire [4-1:0] node55904;
	wire [4-1:0] node55907;
	wire [4-1:0] node55910;
	wire [4-1:0] node55912;
	wire [4-1:0] node55913;
	wire [4-1:0] node55916;
	wire [4-1:0] node55919;
	wire [4-1:0] node55920;
	wire [4-1:0] node55921;
	wire [4-1:0] node55922;
	wire [4-1:0] node55923;
	wire [4-1:0] node55925;
	wire [4-1:0] node55928;
	wire [4-1:0] node55929;
	wire [4-1:0] node55930;
	wire [4-1:0] node55933;
	wire [4-1:0] node55936;
	wire [4-1:0] node55937;
	wire [4-1:0] node55940;
	wire [4-1:0] node55943;
	wire [4-1:0] node55944;
	wire [4-1:0] node55945;
	wire [4-1:0] node55948;
	wire [4-1:0] node55951;
	wire [4-1:0] node55952;
	wire [4-1:0] node55955;
	wire [4-1:0] node55958;
	wire [4-1:0] node55959;
	wire [4-1:0] node55960;
	wire [4-1:0] node55961;
	wire [4-1:0] node55962;
	wire [4-1:0] node55965;
	wire [4-1:0] node55969;
	wire [4-1:0] node55971;
	wire [4-1:0] node55972;
	wire [4-1:0] node55976;
	wire [4-1:0] node55977;
	wire [4-1:0] node55980;
	wire [4-1:0] node55983;
	wire [4-1:0] node55984;
	wire [4-1:0] node55985;
	wire [4-1:0] node55986;
	wire [4-1:0] node55988;
	wire [4-1:0] node55989;
	wire [4-1:0] node55992;
	wire [4-1:0] node55996;
	wire [4-1:0] node55997;
	wire [4-1:0] node55998;
	wire [4-1:0] node55999;
	wire [4-1:0] node56004;
	wire [4-1:0] node56005;
	wire [4-1:0] node56008;
	wire [4-1:0] node56011;
	wire [4-1:0] node56012;
	wire [4-1:0] node56013;
	wire [4-1:0] node56014;
	wire [4-1:0] node56016;
	wire [4-1:0] node56019;
	wire [4-1:0] node56021;
	wire [4-1:0] node56024;
	wire [4-1:0] node56025;
	wire [4-1:0] node56026;
	wire [4-1:0] node56029;
	wire [4-1:0] node56033;
	wire [4-1:0] node56034;
	wire [4-1:0] node56035;
	wire [4-1:0] node56036;
	wire [4-1:0] node56040;
	wire [4-1:0] node56041;
	wire [4-1:0] node56045;
	wire [4-1:0] node56046;
	wire [4-1:0] node56049;
	wire [4-1:0] node56052;
	wire [4-1:0] node56053;
	wire [4-1:0] node56054;
	wire [4-1:0] node56055;
	wire [4-1:0] node56056;
	wire [4-1:0] node56057;
	wire [4-1:0] node56060;
	wire [4-1:0] node56063;
	wire [4-1:0] node56064;
	wire [4-1:0] node56067;
	wire [4-1:0] node56070;
	wire [4-1:0] node56071;
	wire [4-1:0] node56072;
	wire [4-1:0] node56076;
	wire [4-1:0] node56079;
	wire [4-1:0] node56080;
	wire [4-1:0] node56081;
	wire [4-1:0] node56082;
	wire [4-1:0] node56085;
	wire [4-1:0] node56088;
	wire [4-1:0] node56089;
	wire [4-1:0] node56092;
	wire [4-1:0] node56095;
	wire [4-1:0] node56096;
	wire [4-1:0] node56097;
	wire [4-1:0] node56101;
	wire [4-1:0] node56104;
	wire [4-1:0] node56105;
	wire [4-1:0] node56106;
	wire [4-1:0] node56107;
	wire [4-1:0] node56108;
	wire [4-1:0] node56109;
	wire [4-1:0] node56110;
	wire [4-1:0] node56113;
	wire [4-1:0] node56116;
	wire [4-1:0] node56117;
	wire [4-1:0] node56121;
	wire [4-1:0] node56122;
	wire [4-1:0] node56124;
	wire [4-1:0] node56128;
	wire [4-1:0] node56129;
	wire [4-1:0] node56132;
	wire [4-1:0] node56135;
	wire [4-1:0] node56136;
	wire [4-1:0] node56137;
	wire [4-1:0] node56141;
	wire [4-1:0] node56144;
	wire [4-1:0] node56145;
	wire [4-1:0] node56146;
	wire [4-1:0] node56147;
	wire [4-1:0] node56148;
	wire [4-1:0] node56151;
	wire [4-1:0] node56154;
	wire [4-1:0] node56155;
	wire [4-1:0] node56158;
	wire [4-1:0] node56161;
	wire [4-1:0] node56162;
	wire [4-1:0] node56165;
	wire [4-1:0] node56168;
	wire [4-1:0] node56169;
	wire [4-1:0] node56170;
	wire [4-1:0] node56173;
	wire [4-1:0] node56176;
	wire [4-1:0] node56177;
	wire [4-1:0] node56180;
	wire [4-1:0] node56183;
	wire [4-1:0] node56184;
	wire [4-1:0] node56185;
	wire [4-1:0] node56186;
	wire [4-1:0] node56187;
	wire [4-1:0] node56188;
	wire [4-1:0] node56189;
	wire [4-1:0] node56190;
	wire [4-1:0] node56191;
	wire [4-1:0] node56192;
	wire [4-1:0] node56195;
	wire [4-1:0] node56198;
	wire [4-1:0] node56200;
	wire [4-1:0] node56201;
	wire [4-1:0] node56204;
	wire [4-1:0] node56207;
	wire [4-1:0] node56208;
	wire [4-1:0] node56209;
	wire [4-1:0] node56212;
	wire [4-1:0] node56215;
	wire [4-1:0] node56216;
	wire [4-1:0] node56217;
	wire [4-1:0] node56220;
	wire [4-1:0] node56223;
	wire [4-1:0] node56224;
	wire [4-1:0] node56228;
	wire [4-1:0] node56229;
	wire [4-1:0] node56230;
	wire [4-1:0] node56232;
	wire [4-1:0] node56235;
	wire [4-1:0] node56237;
	wire [4-1:0] node56240;
	wire [4-1:0] node56241;
	wire [4-1:0] node56243;
	wire [4-1:0] node56246;
	wire [4-1:0] node56248;
	wire [4-1:0] node56251;
	wire [4-1:0] node56252;
	wire [4-1:0] node56253;
	wire [4-1:0] node56254;
	wire [4-1:0] node56255;
	wire [4-1:0] node56256;
	wire [4-1:0] node56260;
	wire [4-1:0] node56262;
	wire [4-1:0] node56266;
	wire [4-1:0] node56267;
	wire [4-1:0] node56269;
	wire [4-1:0] node56270;
	wire [4-1:0] node56274;
	wire [4-1:0] node56275;
	wire [4-1:0] node56278;
	wire [4-1:0] node56281;
	wire [4-1:0] node56282;
	wire [4-1:0] node56283;
	wire [4-1:0] node56284;
	wire [4-1:0] node56285;
	wire [4-1:0] node56288;
	wire [4-1:0] node56292;
	wire [4-1:0] node56293;
	wire [4-1:0] node56296;
	wire [4-1:0] node56299;
	wire [4-1:0] node56300;
	wire [4-1:0] node56303;
	wire [4-1:0] node56306;
	wire [4-1:0] node56307;
	wire [4-1:0] node56308;
	wire [4-1:0] node56309;
	wire [4-1:0] node56310;
	wire [4-1:0] node56311;
	wire [4-1:0] node56314;
	wire [4-1:0] node56316;
	wire [4-1:0] node56319;
	wire [4-1:0] node56320;
	wire [4-1:0] node56322;
	wire [4-1:0] node56326;
	wire [4-1:0] node56327;
	wire [4-1:0] node56328;
	wire [4-1:0] node56330;
	wire [4-1:0] node56333;
	wire [4-1:0] node56336;
	wire [4-1:0] node56337;
	wire [4-1:0] node56338;
	wire [4-1:0] node56341;
	wire [4-1:0] node56345;
	wire [4-1:0] node56346;
	wire [4-1:0] node56347;
	wire [4-1:0] node56348;
	wire [4-1:0] node56352;
	wire [4-1:0] node56353;
	wire [4-1:0] node56357;
	wire [4-1:0] node56358;
	wire [4-1:0] node56359;
	wire [4-1:0] node56360;
	wire [4-1:0] node56363;
	wire [4-1:0] node56368;
	wire [4-1:0] node56369;
	wire [4-1:0] node56370;
	wire [4-1:0] node56371;
	wire [4-1:0] node56372;
	wire [4-1:0] node56373;
	wire [4-1:0] node56376;
	wire [4-1:0] node56380;
	wire [4-1:0] node56381;
	wire [4-1:0] node56383;
	wire [4-1:0] node56386;
	wire [4-1:0] node56387;
	wire [4-1:0] node56390;
	wire [4-1:0] node56393;
	wire [4-1:0] node56394;
	wire [4-1:0] node56395;
	wire [4-1:0] node56396;
	wire [4-1:0] node56400;
	wire [4-1:0] node56403;
	wire [4-1:0] node56405;
	wire [4-1:0] node56406;
	wire [4-1:0] node56410;
	wire [4-1:0] node56411;
	wire [4-1:0] node56412;
	wire [4-1:0] node56413;
	wire [4-1:0] node56417;
	wire [4-1:0] node56418;
	wire [4-1:0] node56422;
	wire [4-1:0] node56423;
	wire [4-1:0] node56424;
	wire [4-1:0] node56428;
	wire [4-1:0] node56429;
	wire [4-1:0] node56433;
	wire [4-1:0] node56434;
	wire [4-1:0] node56435;
	wire [4-1:0] node56436;
	wire [4-1:0] node56437;
	wire [4-1:0] node56438;
	wire [4-1:0] node56439;
	wire [4-1:0] node56442;
	wire [4-1:0] node56445;
	wire [4-1:0] node56446;
	wire [4-1:0] node56448;
	wire [4-1:0] node56451;
	wire [4-1:0] node56452;
	wire [4-1:0] node56455;
	wire [4-1:0] node56458;
	wire [4-1:0] node56459;
	wire [4-1:0] node56460;
	wire [4-1:0] node56463;
	wire [4-1:0] node56466;
	wire [4-1:0] node56467;
	wire [4-1:0] node56468;
	wire [4-1:0] node56473;
	wire [4-1:0] node56474;
	wire [4-1:0] node56475;
	wire [4-1:0] node56476;
	wire [4-1:0] node56479;
	wire [4-1:0] node56482;
	wire [4-1:0] node56484;
	wire [4-1:0] node56486;
	wire [4-1:0] node56489;
	wire [4-1:0] node56490;
	wire [4-1:0] node56492;
	wire [4-1:0] node56495;
	wire [4-1:0] node56496;
	wire [4-1:0] node56499;
	wire [4-1:0] node56502;
	wire [4-1:0] node56503;
	wire [4-1:0] node56504;
	wire [4-1:0] node56505;
	wire [4-1:0] node56506;
	wire [4-1:0] node56509;
	wire [4-1:0] node56512;
	wire [4-1:0] node56513;
	wire [4-1:0] node56514;
	wire [4-1:0] node56517;
	wire [4-1:0] node56521;
	wire [4-1:0] node56522;
	wire [4-1:0] node56523;
	wire [4-1:0] node56524;
	wire [4-1:0] node56527;
	wire [4-1:0] node56530;
	wire [4-1:0] node56532;
	wire [4-1:0] node56535;
	wire [4-1:0] node56537;
	wire [4-1:0] node56540;
	wire [4-1:0] node56541;
	wire [4-1:0] node56542;
	wire [4-1:0] node56544;
	wire [4-1:0] node56545;
	wire [4-1:0] node56548;
	wire [4-1:0] node56551;
	wire [4-1:0] node56552;
	wire [4-1:0] node56554;
	wire [4-1:0] node56558;
	wire [4-1:0] node56559;
	wire [4-1:0] node56560;
	wire [4-1:0] node56561;
	wire [4-1:0] node56564;
	wire [4-1:0] node56569;
	wire [4-1:0] node56570;
	wire [4-1:0] node56571;
	wire [4-1:0] node56572;
	wire [4-1:0] node56573;
	wire [4-1:0] node56574;
	wire [4-1:0] node56575;
	wire [4-1:0] node56579;
	wire [4-1:0] node56582;
	wire [4-1:0] node56583;
	wire [4-1:0] node56585;
	wire [4-1:0] node56588;
	wire [4-1:0] node56589;
	wire [4-1:0] node56592;
	wire [4-1:0] node56595;
	wire [4-1:0] node56596;
	wire [4-1:0] node56597;
	wire [4-1:0] node56598;
	wire [4-1:0] node56601;
	wire [4-1:0] node56604;
	wire [4-1:0] node56607;
	wire [4-1:0] node56608;
	wire [4-1:0] node56609;
	wire [4-1:0] node56612;
	wire [4-1:0] node56615;
	wire [4-1:0] node56616;
	wire [4-1:0] node56619;
	wire [4-1:0] node56622;
	wire [4-1:0] node56623;
	wire [4-1:0] node56624;
	wire [4-1:0] node56626;
	wire [4-1:0] node56629;
	wire [4-1:0] node56630;
	wire [4-1:0] node56633;
	wire [4-1:0] node56636;
	wire [4-1:0] node56637;
	wire [4-1:0] node56638;
	wire [4-1:0] node56641;
	wire [4-1:0] node56644;
	wire [4-1:0] node56645;
	wire [4-1:0] node56648;
	wire [4-1:0] node56651;
	wire [4-1:0] node56652;
	wire [4-1:0] node56653;
	wire [4-1:0] node56654;
	wire [4-1:0] node56655;
	wire [4-1:0] node56658;
	wire [4-1:0] node56659;
	wire [4-1:0] node56663;
	wire [4-1:0] node56664;
	wire [4-1:0] node56667;
	wire [4-1:0] node56670;
	wire [4-1:0] node56671;
	wire [4-1:0] node56672;
	wire [4-1:0] node56673;
	wire [4-1:0] node56677;
	wire [4-1:0] node56680;
	wire [4-1:0] node56682;
	wire [4-1:0] node56685;
	wire [4-1:0] node56686;
	wire [4-1:0] node56687;
	wire [4-1:0] node56688;
	wire [4-1:0] node56689;
	wire [4-1:0] node56692;
	wire [4-1:0] node56695;
	wire [4-1:0] node56697;
	wire [4-1:0] node56700;
	wire [4-1:0] node56701;
	wire [4-1:0] node56705;
	wire [4-1:0] node56706;
	wire [4-1:0] node56707;
	wire [4-1:0] node56709;
	wire [4-1:0] node56713;
	wire [4-1:0] node56714;
	wire [4-1:0] node56715;
	wire [4-1:0] node56719;
	wire [4-1:0] node56720;
	wire [4-1:0] node56723;
	wire [4-1:0] node56726;
	wire [4-1:0] node56727;
	wire [4-1:0] node56728;
	wire [4-1:0] node56729;
	wire [4-1:0] node56730;
	wire [4-1:0] node56731;
	wire [4-1:0] node56732;
	wire [4-1:0] node56733;
	wire [4-1:0] node56736;
	wire [4-1:0] node56739;
	wire [4-1:0] node56740;
	wire [4-1:0] node56743;
	wire [4-1:0] node56746;
	wire [4-1:0] node56747;
	wire [4-1:0] node56748;
	wire [4-1:0] node56751;
	wire [4-1:0] node56754;
	wire [4-1:0] node56755;
	wire [4-1:0] node56756;
	wire [4-1:0] node56760;
	wire [4-1:0] node56761;
	wire [4-1:0] node56764;
	wire [4-1:0] node56767;
	wire [4-1:0] node56768;
	wire [4-1:0] node56769;
	wire [4-1:0] node56770;
	wire [4-1:0] node56774;
	wire [4-1:0] node56776;
	wire [4-1:0] node56779;
	wire [4-1:0] node56780;
	wire [4-1:0] node56781;
	wire [4-1:0] node56785;
	wire [4-1:0] node56786;
	wire [4-1:0] node56790;
	wire [4-1:0] node56791;
	wire [4-1:0] node56792;
	wire [4-1:0] node56793;
	wire [4-1:0] node56794;
	wire [4-1:0] node56798;
	wire [4-1:0] node56799;
	wire [4-1:0] node56803;
	wire [4-1:0] node56804;
	wire [4-1:0] node56806;
	wire [4-1:0] node56809;
	wire [4-1:0] node56810;
	wire [4-1:0] node56814;
	wire [4-1:0] node56815;
	wire [4-1:0] node56816;
	wire [4-1:0] node56817;
	wire [4-1:0] node56821;
	wire [4-1:0] node56822;
	wire [4-1:0] node56826;
	wire [4-1:0] node56827;
	wire [4-1:0] node56828;
	wire [4-1:0] node56832;
	wire [4-1:0] node56833;
	wire [4-1:0] node56837;
	wire [4-1:0] node56838;
	wire [4-1:0] node56839;
	wire [4-1:0] node56840;
	wire [4-1:0] node56842;
	wire [4-1:0] node56843;
	wire [4-1:0] node56847;
	wire [4-1:0] node56848;
	wire [4-1:0] node56850;
	wire [4-1:0] node56851;
	wire [4-1:0] node56855;
	wire [4-1:0] node56858;
	wire [4-1:0] node56859;
	wire [4-1:0] node56860;
	wire [4-1:0] node56861;
	wire [4-1:0] node56865;
	wire [4-1:0] node56868;
	wire [4-1:0] node56869;
	wire [4-1:0] node56870;
	wire [4-1:0] node56874;
	wire [4-1:0] node56877;
	wire [4-1:0] node56878;
	wire [4-1:0] node56879;
	wire [4-1:0] node56880;
	wire [4-1:0] node56881;
	wire [4-1:0] node56885;
	wire [4-1:0] node56886;
	wire [4-1:0] node56890;
	wire [4-1:0] node56892;
	wire [4-1:0] node56893;
	wire [4-1:0] node56897;
	wire [4-1:0] node56898;
	wire [4-1:0] node56899;
	wire [4-1:0] node56900;
	wire [4-1:0] node56903;
	wire [4-1:0] node56906;
	wire [4-1:0] node56907;
	wire [4-1:0] node56908;
	wire [4-1:0] node56911;
	wire [4-1:0] node56914;
	wire [4-1:0] node56915;
	wire [4-1:0] node56918;
	wire [4-1:0] node56921;
	wire [4-1:0] node56922;
	wire [4-1:0] node56925;
	wire [4-1:0] node56928;
	wire [4-1:0] node56929;
	wire [4-1:0] node56930;
	wire [4-1:0] node56931;
	wire [4-1:0] node56932;
	wire [4-1:0] node56933;
	wire [4-1:0] node56934;
	wire [4-1:0] node56938;
	wire [4-1:0] node56939;
	wire [4-1:0] node56943;
	wire [4-1:0] node56944;
	wire [4-1:0] node56945;
	wire [4-1:0] node56950;
	wire [4-1:0] node56951;
	wire [4-1:0] node56952;
	wire [4-1:0] node56953;
	wire [4-1:0] node56957;
	wire [4-1:0] node56958;
	wire [4-1:0] node56962;
	wire [4-1:0] node56963;
	wire [4-1:0] node56964;
	wire [4-1:0] node56968;
	wire [4-1:0] node56969;
	wire [4-1:0] node56973;
	wire [4-1:0] node56974;
	wire [4-1:0] node56975;
	wire [4-1:0] node56976;
	wire [4-1:0] node56979;
	wire [4-1:0] node56980;
	wire [4-1:0] node56984;
	wire [4-1:0] node56986;
	wire [4-1:0] node56989;
	wire [4-1:0] node56990;
	wire [4-1:0] node56992;
	wire [4-1:0] node56995;
	wire [4-1:0] node56996;
	wire [4-1:0] node56997;
	wire [4-1:0] node57001;
	wire [4-1:0] node57004;
	wire [4-1:0] node57005;
	wire [4-1:0] node57006;
	wire [4-1:0] node57007;
	wire [4-1:0] node57008;
	wire [4-1:0] node57009;
	wire [4-1:0] node57013;
	wire [4-1:0] node57014;
	wire [4-1:0] node57018;
	wire [4-1:0] node57020;
	wire [4-1:0] node57021;
	wire [4-1:0] node57025;
	wire [4-1:0] node57026;
	wire [4-1:0] node57027;
	wire [4-1:0] node57028;
	wire [4-1:0] node57032;
	wire [4-1:0] node57033;
	wire [4-1:0] node57037;
	wire [4-1:0] node57038;
	wire [4-1:0] node57039;
	wire [4-1:0] node57043;
	wire [4-1:0] node57044;
	wire [4-1:0] node57048;
	wire [4-1:0] node57049;
	wire [4-1:0] node57050;
	wire [4-1:0] node57052;
	wire [4-1:0] node57053;
	wire [4-1:0] node57057;
	wire [4-1:0] node57058;
	wire [4-1:0] node57059;
	wire [4-1:0] node57063;
	wire [4-1:0] node57064;
	wire [4-1:0] node57068;
	wire [4-1:0] node57069;
	wire [4-1:0] node57070;
	wire [4-1:0] node57073;
	wire [4-1:0] node57074;
	wire [4-1:0] node57078;
	wire [4-1:0] node57079;
	wire [4-1:0] node57080;
	wire [4-1:0] node57085;
	wire [4-1:0] node57086;
	wire [4-1:0] node57087;
	wire [4-1:0] node57088;
	wire [4-1:0] node57089;
	wire [4-1:0] node57090;
	wire [4-1:0] node57091;
	wire [4-1:0] node57092;
	wire [4-1:0] node57093;
	wire [4-1:0] node57094;
	wire [4-1:0] node57097;
	wire [4-1:0] node57100;
	wire [4-1:0] node57101;
	wire [4-1:0] node57105;
	wire [4-1:0] node57108;
	wire [4-1:0] node57109;
	wire [4-1:0] node57110;
	wire [4-1:0] node57113;
	wire [4-1:0] node57114;
	wire [4-1:0] node57117;
	wire [4-1:0] node57120;
	wire [4-1:0] node57121;
	wire [4-1:0] node57124;
	wire [4-1:0] node57125;
	wire [4-1:0] node57128;
	wire [4-1:0] node57131;
	wire [4-1:0] node57132;
	wire [4-1:0] node57133;
	wire [4-1:0] node57134;
	wire [4-1:0] node57135;
	wire [4-1:0] node57138;
	wire [4-1:0] node57141;
	wire [4-1:0] node57142;
	wire [4-1:0] node57145;
	wire [4-1:0] node57148;
	wire [4-1:0] node57149;
	wire [4-1:0] node57151;
	wire [4-1:0] node57154;
	wire [4-1:0] node57155;
	wire [4-1:0] node57158;
	wire [4-1:0] node57161;
	wire [4-1:0] node57162;
	wire [4-1:0] node57164;
	wire [4-1:0] node57166;
	wire [4-1:0] node57169;
	wire [4-1:0] node57170;
	wire [4-1:0] node57172;
	wire [4-1:0] node57175;
	wire [4-1:0] node57178;
	wire [4-1:0] node57179;
	wire [4-1:0] node57180;
	wire [4-1:0] node57181;
	wire [4-1:0] node57182;
	wire [4-1:0] node57183;
	wire [4-1:0] node57186;
	wire [4-1:0] node57189;
	wire [4-1:0] node57191;
	wire [4-1:0] node57194;
	wire [4-1:0] node57196;
	wire [4-1:0] node57197;
	wire [4-1:0] node57200;
	wire [4-1:0] node57203;
	wire [4-1:0] node57204;
	wire [4-1:0] node57205;
	wire [4-1:0] node57206;
	wire [4-1:0] node57209;
	wire [4-1:0] node57212;
	wire [4-1:0] node57213;
	wire [4-1:0] node57217;
	wire [4-1:0] node57218;
	wire [4-1:0] node57219;
	wire [4-1:0] node57222;
	wire [4-1:0] node57225;
	wire [4-1:0] node57226;
	wire [4-1:0] node57229;
	wire [4-1:0] node57232;
	wire [4-1:0] node57233;
	wire [4-1:0] node57234;
	wire [4-1:0] node57236;
	wire [4-1:0] node57237;
	wire [4-1:0] node57241;
	wire [4-1:0] node57242;
	wire [4-1:0] node57243;
	wire [4-1:0] node57246;
	wire [4-1:0] node57250;
	wire [4-1:0] node57251;
	wire [4-1:0] node57252;
	wire [4-1:0] node57254;
	wire [4-1:0] node57257;
	wire [4-1:0] node57258;
	wire [4-1:0] node57262;
	wire [4-1:0] node57263;
	wire [4-1:0] node57264;
	wire [4-1:0] node57267;
	wire [4-1:0] node57270;
	wire [4-1:0] node57271;
	wire [4-1:0] node57275;
	wire [4-1:0] node57276;
	wire [4-1:0] node57277;
	wire [4-1:0] node57278;
	wire [4-1:0] node57280;
	wire [4-1:0] node57281;
	wire [4-1:0] node57282;
	wire [4-1:0] node57285;
	wire [4-1:0] node57288;
	wire [4-1:0] node57289;
	wire [4-1:0] node57292;
	wire [4-1:0] node57295;
	wire [4-1:0] node57296;
	wire [4-1:0] node57298;
	wire [4-1:0] node57301;
	wire [4-1:0] node57303;
	wire [4-1:0] node57306;
	wire [4-1:0] node57307;
	wire [4-1:0] node57308;
	wire [4-1:0] node57310;
	wire [4-1:0] node57311;
	wire [4-1:0] node57314;
	wire [4-1:0] node57317;
	wire [4-1:0] node57319;
	wire [4-1:0] node57320;
	wire [4-1:0] node57324;
	wire [4-1:0] node57325;
	wire [4-1:0] node57326;
	wire [4-1:0] node57329;
	wire [4-1:0] node57332;
	wire [4-1:0] node57333;
	wire [4-1:0] node57336;
	wire [4-1:0] node57339;
	wire [4-1:0] node57340;
	wire [4-1:0] node57341;
	wire [4-1:0] node57342;
	wire [4-1:0] node57343;
	wire [4-1:0] node57347;
	wire [4-1:0] node57348;
	wire [4-1:0] node57352;
	wire [4-1:0] node57353;
	wire [4-1:0] node57354;
	wire [4-1:0] node57358;
	wire [4-1:0] node57359;
	wire [4-1:0] node57363;
	wire [4-1:0] node57364;
	wire [4-1:0] node57365;
	wire [4-1:0] node57366;
	wire [4-1:0] node57370;
	wire [4-1:0] node57371;
	wire [4-1:0] node57375;
	wire [4-1:0] node57376;
	wire [4-1:0] node57377;
	wire [4-1:0] node57382;
	wire [4-1:0] node57383;
	wire [4-1:0] node57384;
	wire [4-1:0] node57385;
	wire [4-1:0] node57386;
	wire [4-1:0] node57387;
	wire [4-1:0] node57388;
	wire [4-1:0] node57389;
	wire [4-1:0] node57394;
	wire [4-1:0] node57395;
	wire [4-1:0] node57396;
	wire [4-1:0] node57399;
	wire [4-1:0] node57403;
	wire [4-1:0] node57404;
	wire [4-1:0] node57407;
	wire [4-1:0] node57410;
	wire [4-1:0] node57411;
	wire [4-1:0] node57412;
	wire [4-1:0] node57414;
	wire [4-1:0] node57415;
	wire [4-1:0] node57419;
	wire [4-1:0] node57421;
	wire [4-1:0] node57424;
	wire [4-1:0] node57425;
	wire [4-1:0] node57426;
	wire [4-1:0] node57429;
	wire [4-1:0] node57432;
	wire [4-1:0] node57434;
	wire [4-1:0] node57437;
	wire [4-1:0] node57438;
	wire [4-1:0] node57439;
	wire [4-1:0] node57440;
	wire [4-1:0] node57441;
	wire [4-1:0] node57442;
	wire [4-1:0] node57445;
	wire [4-1:0] node57448;
	wire [4-1:0] node57449;
	wire [4-1:0] node57452;
	wire [4-1:0] node57455;
	wire [4-1:0] node57457;
	wire [4-1:0] node57458;
	wire [4-1:0] node57461;
	wire [4-1:0] node57464;
	wire [4-1:0] node57465;
	wire [4-1:0] node57467;
	wire [4-1:0] node57470;
	wire [4-1:0] node57471;
	wire [4-1:0] node57472;
	wire [4-1:0] node57475;
	wire [4-1:0] node57478;
	wire [4-1:0] node57479;
	wire [4-1:0] node57482;
	wire [4-1:0] node57485;
	wire [4-1:0] node57486;
	wire [4-1:0] node57487;
	wire [4-1:0] node57489;
	wire [4-1:0] node57490;
	wire [4-1:0] node57494;
	wire [4-1:0] node57495;
	wire [4-1:0] node57496;
	wire [4-1:0] node57499;
	wire [4-1:0] node57502;
	wire [4-1:0] node57503;
	wire [4-1:0] node57507;
	wire [4-1:0] node57508;
	wire [4-1:0] node57509;
	wire [4-1:0] node57510;
	wire [4-1:0] node57513;
	wire [4-1:0] node57516;
	wire [4-1:0] node57517;
	wire [4-1:0] node57520;
	wire [4-1:0] node57523;
	wire [4-1:0] node57524;
	wire [4-1:0] node57525;
	wire [4-1:0] node57528;
	wire [4-1:0] node57532;
	wire [4-1:0] node57533;
	wire [4-1:0] node57534;
	wire [4-1:0] node57535;
	wire [4-1:0] node57536;
	wire [4-1:0] node57537;
	wire [4-1:0] node57539;
	wire [4-1:0] node57543;
	wire [4-1:0] node57544;
	wire [4-1:0] node57545;
	wire [4-1:0] node57548;
	wire [4-1:0] node57551;
	wire [4-1:0] node57552;
	wire [4-1:0] node57556;
	wire [4-1:0] node57557;
	wire [4-1:0] node57559;
	wire [4-1:0] node57560;
	wire [4-1:0] node57563;
	wire [4-1:0] node57566;
	wire [4-1:0] node57567;
	wire [4-1:0] node57570;
	wire [4-1:0] node57573;
	wire [4-1:0] node57574;
	wire [4-1:0] node57575;
	wire [4-1:0] node57576;
	wire [4-1:0] node57577;
	wire [4-1:0] node57580;
	wire [4-1:0] node57583;
	wire [4-1:0] node57584;
	wire [4-1:0] node57587;
	wire [4-1:0] node57590;
	wire [4-1:0] node57591;
	wire [4-1:0] node57592;
	wire [4-1:0] node57596;
	wire [4-1:0] node57599;
	wire [4-1:0] node57600;
	wire [4-1:0] node57601;
	wire [4-1:0] node57604;
	wire [4-1:0] node57607;
	wire [4-1:0] node57609;
	wire [4-1:0] node57612;
	wire [4-1:0] node57613;
	wire [4-1:0] node57614;
	wire [4-1:0] node57615;
	wire [4-1:0] node57619;
	wire [4-1:0] node57620;
	wire [4-1:0] node57622;
	wire [4-1:0] node57623;
	wire [4-1:0] node57626;
	wire [4-1:0] node57629;
	wire [4-1:0] node57630;
	wire [4-1:0] node57633;
	wire [4-1:0] node57636;
	wire [4-1:0] node57637;
	wire [4-1:0] node57638;
	wire [4-1:0] node57639;
	wire [4-1:0] node57642;
	wire [4-1:0] node57645;
	wire [4-1:0] node57646;
	wire [4-1:0] node57649;
	wire [4-1:0] node57652;
	wire [4-1:0] node57653;
	wire [4-1:0] node57654;
	wire [4-1:0] node57657;
	wire [4-1:0] node57660;
	wire [4-1:0] node57661;
	wire [4-1:0] node57664;
	wire [4-1:0] node57667;
	wire [4-1:0] node57668;
	wire [4-1:0] node57669;
	wire [4-1:0] node57670;
	wire [4-1:0] node57671;
	wire [4-1:0] node57672;
	wire [4-1:0] node57673;
	wire [4-1:0] node57674;
	wire [4-1:0] node57677;
	wire [4-1:0] node57680;
	wire [4-1:0] node57681;
	wire [4-1:0] node57682;
	wire [4-1:0] node57685;
	wire [4-1:0] node57689;
	wire [4-1:0] node57691;
	wire [4-1:0] node57692;
	wire [4-1:0] node57694;
	wire [4-1:0] node57698;
	wire [4-1:0] node57699;
	wire [4-1:0] node57700;
	wire [4-1:0] node57701;
	wire [4-1:0] node57706;
	wire [4-1:0] node57707;
	wire [4-1:0] node57708;
	wire [4-1:0] node57712;
	wire [4-1:0] node57715;
	wire [4-1:0] node57716;
	wire [4-1:0] node57717;
	wire [4-1:0] node57718;
	wire [4-1:0] node57719;
	wire [4-1:0] node57720;
	wire [4-1:0] node57723;
	wire [4-1:0] node57726;
	wire [4-1:0] node57727;
	wire [4-1:0] node57730;
	wire [4-1:0] node57733;
	wire [4-1:0] node57734;
	wire [4-1:0] node57736;
	wire [4-1:0] node57739;
	wire [4-1:0] node57740;
	wire [4-1:0] node57743;
	wire [4-1:0] node57746;
	wire [4-1:0] node57747;
	wire [4-1:0] node57750;
	wire [4-1:0] node57753;
	wire [4-1:0] node57754;
	wire [4-1:0] node57755;
	wire [4-1:0] node57756;
	wire [4-1:0] node57760;
	wire [4-1:0] node57761;
	wire [4-1:0] node57765;
	wire [4-1:0] node57766;
	wire [4-1:0] node57767;
	wire [4-1:0] node57771;
	wire [4-1:0] node57772;
	wire [4-1:0] node57776;
	wire [4-1:0] node57777;
	wire [4-1:0] node57778;
	wire [4-1:0] node57779;
	wire [4-1:0] node57780;
	wire [4-1:0] node57781;
	wire [4-1:0] node57784;
	wire [4-1:0] node57787;
	wire [4-1:0] node57788;
	wire [4-1:0] node57791;
	wire [4-1:0] node57792;
	wire [4-1:0] node57796;
	wire [4-1:0] node57797;
	wire [4-1:0] node57798;
	wire [4-1:0] node57799;
	wire [4-1:0] node57803;
	wire [4-1:0] node57804;
	wire [4-1:0] node57808;
	wire [4-1:0] node57810;
	wire [4-1:0] node57813;
	wire [4-1:0] node57814;
	wire [4-1:0] node57815;
	wire [4-1:0] node57816;
	wire [4-1:0] node57820;
	wire [4-1:0] node57821;
	wire [4-1:0] node57825;
	wire [4-1:0] node57826;
	wire [4-1:0] node57827;
	wire [4-1:0] node57832;
	wire [4-1:0] node57833;
	wire [4-1:0] node57834;
	wire [4-1:0] node57836;
	wire [4-1:0] node57837;
	wire [4-1:0] node57841;
	wire [4-1:0] node57842;
	wire [4-1:0] node57843;
	wire [4-1:0] node57847;
	wire [4-1:0] node57848;
	wire [4-1:0] node57852;
	wire [4-1:0] node57853;
	wire [4-1:0] node57854;
	wire [4-1:0] node57855;
	wire [4-1:0] node57859;
	wire [4-1:0] node57860;
	wire [4-1:0] node57864;
	wire [4-1:0] node57865;
	wire [4-1:0] node57866;
	wire [4-1:0] node57870;
	wire [4-1:0] node57871;
	wire [4-1:0] node57875;
	wire [4-1:0] node57876;
	wire [4-1:0] node57877;
	wire [4-1:0] node57878;
	wire [4-1:0] node57879;
	wire [4-1:0] node57880;
	wire [4-1:0] node57881;
	wire [4-1:0] node57884;
	wire [4-1:0] node57887;
	wire [4-1:0] node57888;
	wire [4-1:0] node57891;
	wire [4-1:0] node57894;
	wire [4-1:0] node57895;
	wire [4-1:0] node57896;
	wire [4-1:0] node57899;
	wire [4-1:0] node57902;
	wire [4-1:0] node57903;
	wire [4-1:0] node57907;
	wire [4-1:0] node57908;
	wire [4-1:0] node57909;
	wire [4-1:0] node57910;
	wire [4-1:0] node57913;
	wire [4-1:0] node57916;
	wire [4-1:0] node57917;
	wire [4-1:0] node57920;
	wire [4-1:0] node57923;
	wire [4-1:0] node57924;
	wire [4-1:0] node57925;
	wire [4-1:0] node57928;
	wire [4-1:0] node57931;
	wire [4-1:0] node57932;
	wire [4-1:0] node57933;
	wire [4-1:0] node57936;
	wire [4-1:0] node57939;
	wire [4-1:0] node57941;
	wire [4-1:0] node57944;
	wire [4-1:0] node57945;
	wire [4-1:0] node57946;
	wire [4-1:0] node57947;
	wire [4-1:0] node57948;
	wire [4-1:0] node57951;
	wire [4-1:0] node57954;
	wire [4-1:0] node57956;
	wire [4-1:0] node57957;
	wire [4-1:0] node57960;
	wire [4-1:0] node57963;
	wire [4-1:0] node57964;
	wire [4-1:0] node57965;
	wire [4-1:0] node57966;
	wire [4-1:0] node57969;
	wire [4-1:0] node57972;
	wire [4-1:0] node57973;
	wire [4-1:0] node57976;
	wire [4-1:0] node57979;
	wire [4-1:0] node57980;
	wire [4-1:0] node57984;
	wire [4-1:0] node57985;
	wire [4-1:0] node57986;
	wire [4-1:0] node57989;
	wire [4-1:0] node57992;
	wire [4-1:0] node57993;
	wire [4-1:0] node57994;
	wire [4-1:0] node57997;
	wire [4-1:0] node58000;
	wire [4-1:0] node58001;
	wire [4-1:0] node58003;
	wire [4-1:0] node58006;
	wire [4-1:0] node58009;
	wire [4-1:0] node58010;
	wire [4-1:0] node58011;
	wire [4-1:0] node58012;
	wire [4-1:0] node58013;
	wire [4-1:0] node58017;
	wire [4-1:0] node58020;
	wire [4-1:0] node58021;
	wire [4-1:0] node58022;
	wire [4-1:0] node58026;
	wire [4-1:0] node58029;
	wire [4-1:0] node58030;
	wire [4-1:0] node58031;
	wire [4-1:0] node58032;
	wire [4-1:0] node58036;
	wire [4-1:0] node58039;
	wire [4-1:0] node58040;
	wire [4-1:0] node58041;
	wire [4-1:0] node58045;
	wire [4-1:0] node58046;
	wire [4-1:0] node58049;
	wire [4-1:0] node58052;
	wire [4-1:0] node58053;
	wire [4-1:0] node58054;
	wire [4-1:0] node58055;
	wire [4-1:0] node58056;
	wire [4-1:0] node58057;
	wire [4-1:0] node58058;
	wire [4-1:0] node58059;
	wire [4-1:0] node58060;
	wire [4-1:0] node58061;
	wire [4-1:0] node58062;
	wire [4-1:0] node58063;
	wire [4-1:0] node58066;
	wire [4-1:0] node58069;
	wire [4-1:0] node58070;
	wire [4-1:0] node58073;
	wire [4-1:0] node58075;
	wire [4-1:0] node58078;
	wire [4-1:0] node58079;
	wire [4-1:0] node58080;
	wire [4-1:0] node58082;
	wire [4-1:0] node58085;
	wire [4-1:0] node58088;
	wire [4-1:0] node58089;
	wire [4-1:0] node58092;
	wire [4-1:0] node58093;
	wire [4-1:0] node58097;
	wire [4-1:0] node58098;
	wire [4-1:0] node58099;
	wire [4-1:0] node58100;
	wire [4-1:0] node58102;
	wire [4-1:0] node58105;
	wire [4-1:0] node58106;
	wire [4-1:0] node58109;
	wire [4-1:0] node58112;
	wire [4-1:0] node58113;
	wire [4-1:0] node58116;
	wire [4-1:0] node58117;
	wire [4-1:0] node58120;
	wire [4-1:0] node58123;
	wire [4-1:0] node58124;
	wire [4-1:0] node58126;
	wire [4-1:0] node58127;
	wire [4-1:0] node58131;
	wire [4-1:0] node58132;
	wire [4-1:0] node58134;
	wire [4-1:0] node58138;
	wire [4-1:0] node58139;
	wire [4-1:0] node58140;
	wire [4-1:0] node58141;
	wire [4-1:0] node58143;
	wire [4-1:0] node58146;
	wire [4-1:0] node58147;
	wire [4-1:0] node58148;
	wire [4-1:0] node58152;
	wire [4-1:0] node58153;
	wire [4-1:0] node58156;
	wire [4-1:0] node58159;
	wire [4-1:0] node58160;
	wire [4-1:0] node58162;
	wire [4-1:0] node58164;
	wire [4-1:0] node58167;
	wire [4-1:0] node58169;
	wire [4-1:0] node58170;
	wire [4-1:0] node58173;
	wire [4-1:0] node58176;
	wire [4-1:0] node58177;
	wire [4-1:0] node58178;
	wire [4-1:0] node58179;
	wire [4-1:0] node58182;
	wire [4-1:0] node58185;
	wire [4-1:0] node58188;
	wire [4-1:0] node58190;
	wire [4-1:0] node58191;
	wire [4-1:0] node58192;
	wire [4-1:0] node58195;
	wire [4-1:0] node58199;
	wire [4-1:0] node58200;
	wire [4-1:0] node58201;
	wire [4-1:0] node58202;
	wire [4-1:0] node58203;
	wire [4-1:0] node58204;
	wire [4-1:0] node58205;
	wire [4-1:0] node58208;
	wire [4-1:0] node58211;
	wire [4-1:0] node58212;
	wire [4-1:0] node58215;
	wire [4-1:0] node58218;
	wire [4-1:0] node58219;
	wire [4-1:0] node58220;
	wire [4-1:0] node58223;
	wire [4-1:0] node58227;
	wire [4-1:0] node58228;
	wire [4-1:0] node58229;
	wire [4-1:0] node58230;
	wire [4-1:0] node58234;
	wire [4-1:0] node58237;
	wire [4-1:0] node58238;
	wire [4-1:0] node58239;
	wire [4-1:0] node58244;
	wire [4-1:0] node58245;
	wire [4-1:0] node58246;
	wire [4-1:0] node58247;
	wire [4-1:0] node58248;
	wire [4-1:0] node58251;
	wire [4-1:0] node58254;
	wire [4-1:0] node58256;
	wire [4-1:0] node58259;
	wire [4-1:0] node58260;
	wire [4-1:0] node58262;
	wire [4-1:0] node58265;
	wire [4-1:0] node58266;
	wire [4-1:0] node58270;
	wire [4-1:0] node58271;
	wire [4-1:0] node58272;
	wire [4-1:0] node58275;
	wire [4-1:0] node58278;
	wire [4-1:0] node58279;
	wire [4-1:0] node58280;
	wire [4-1:0] node58283;
	wire [4-1:0] node58286;
	wire [4-1:0] node58287;
	wire [4-1:0] node58290;
	wire [4-1:0] node58293;
	wire [4-1:0] node58294;
	wire [4-1:0] node58295;
	wire [4-1:0] node58296;
	wire [4-1:0] node58297;
	wire [4-1:0] node58298;
	wire [4-1:0] node58301;
	wire [4-1:0] node58304;
	wire [4-1:0] node58305;
	wire [4-1:0] node58308;
	wire [4-1:0] node58311;
	wire [4-1:0] node58312;
	wire [4-1:0] node58314;
	wire [4-1:0] node58318;
	wire [4-1:0] node58319;
	wire [4-1:0] node58320;
	wire [4-1:0] node58321;
	wire [4-1:0] node58324;
	wire [4-1:0] node58327;
	wire [4-1:0] node58328;
	wire [4-1:0] node58331;
	wire [4-1:0] node58334;
	wire [4-1:0] node58335;
	wire [4-1:0] node58339;
	wire [4-1:0] node58340;
	wire [4-1:0] node58342;
	wire [4-1:0] node58343;
	wire [4-1:0] node58346;
	wire [4-1:0] node58349;
	wire [4-1:0] node58350;
	wire [4-1:0] node58353;
	wire [4-1:0] node58356;
	wire [4-1:0] node58357;
	wire [4-1:0] node58358;
	wire [4-1:0] node58359;
	wire [4-1:0] node58360;
	wire [4-1:0] node58361;
	wire [4-1:0] node58362;
	wire [4-1:0] node58365;
	wire [4-1:0] node58368;
	wire [4-1:0] node58369;
	wire [4-1:0] node58372;
	wire [4-1:0] node58374;
	wire [4-1:0] node58377;
	wire [4-1:0] node58378;
	wire [4-1:0] node58379;
	wire [4-1:0] node58380;
	wire [4-1:0] node58385;
	wire [4-1:0] node58386;
	wire [4-1:0] node58387;
	wire [4-1:0] node58391;
	wire [4-1:0] node58392;
	wire [4-1:0] node58396;
	wire [4-1:0] node58397;
	wire [4-1:0] node58398;
	wire [4-1:0] node58399;
	wire [4-1:0] node58400;
	wire [4-1:0] node58403;
	wire [4-1:0] node58406;
	wire [4-1:0] node58408;
	wire [4-1:0] node58411;
	wire [4-1:0] node58413;
	wire [4-1:0] node58414;
	wire [4-1:0] node58417;
	wire [4-1:0] node58420;
	wire [4-1:0] node58421;
	wire [4-1:0] node58422;
	wire [4-1:0] node58423;
	wire [4-1:0] node58426;
	wire [4-1:0] node58429;
	wire [4-1:0] node58430;
	wire [4-1:0] node58434;
	wire [4-1:0] node58435;
	wire [4-1:0] node58438;
	wire [4-1:0] node58440;
	wire [4-1:0] node58443;
	wire [4-1:0] node58444;
	wire [4-1:0] node58445;
	wire [4-1:0] node58446;
	wire [4-1:0] node58447;
	wire [4-1:0] node58448;
	wire [4-1:0] node58451;
	wire [4-1:0] node58454;
	wire [4-1:0] node58455;
	wire [4-1:0] node58459;
	wire [4-1:0] node58460;
	wire [4-1:0] node58462;
	wire [4-1:0] node58466;
	wire [4-1:0] node58467;
	wire [4-1:0] node58468;
	wire [4-1:0] node58469;
	wire [4-1:0] node58473;
	wire [4-1:0] node58474;
	wire [4-1:0] node58477;
	wire [4-1:0] node58480;
	wire [4-1:0] node58481;
	wire [4-1:0] node58482;
	wire [4-1:0] node58485;
	wire [4-1:0] node58489;
	wire [4-1:0] node58490;
	wire [4-1:0] node58491;
	wire [4-1:0] node58492;
	wire [4-1:0] node58493;
	wire [4-1:0] node58497;
	wire [4-1:0] node58498;
	wire [4-1:0] node58502;
	wire [4-1:0] node58504;
	wire [4-1:0] node58507;
	wire [4-1:0] node58508;
	wire [4-1:0] node58509;
	wire [4-1:0] node58511;
	wire [4-1:0] node58514;
	wire [4-1:0] node58515;
	wire [4-1:0] node58518;
	wire [4-1:0] node58521;
	wire [4-1:0] node58524;
	wire [4-1:0] node58525;
	wire [4-1:0] node58526;
	wire [4-1:0] node58527;
	wire [4-1:0] node58528;
	wire [4-1:0] node58529;
	wire [4-1:0] node58531;
	wire [4-1:0] node58534;
	wire [4-1:0] node58536;
	wire [4-1:0] node58539;
	wire [4-1:0] node58540;
	wire [4-1:0] node58541;
	wire [4-1:0] node58545;
	wire [4-1:0] node58546;
	wire [4-1:0] node58549;
	wire [4-1:0] node58552;
	wire [4-1:0] node58553;
	wire [4-1:0] node58554;
	wire [4-1:0] node58555;
	wire [4-1:0] node58561;
	wire [4-1:0] node58562;
	wire [4-1:0] node58563;
	wire [4-1:0] node58564;
	wire [4-1:0] node58566;
	wire [4-1:0] node58570;
	wire [4-1:0] node58571;
	wire [4-1:0] node58572;
	wire [4-1:0] node58575;
	wire [4-1:0] node58579;
	wire [4-1:0] node58580;
	wire [4-1:0] node58581;
	wire [4-1:0] node58585;
	wire [4-1:0] node58586;
	wire [4-1:0] node58587;
	wire [4-1:0] node58591;
	wire [4-1:0] node58592;
	wire [4-1:0] node58596;
	wire [4-1:0] node58597;
	wire [4-1:0] node58598;
	wire [4-1:0] node58599;
	wire [4-1:0] node58600;
	wire [4-1:0] node58603;
	wire [4-1:0] node58606;
	wire [4-1:0] node58608;
	wire [4-1:0] node58611;
	wire [4-1:0] node58612;
	wire [4-1:0] node58615;
	wire [4-1:0] node58618;
	wire [4-1:0] node58619;
	wire [4-1:0] node58620;
	wire [4-1:0] node58621;
	wire [4-1:0] node58624;
	wire [4-1:0] node58627;
	wire [4-1:0] node58628;
	wire [4-1:0] node58631;
	wire [4-1:0] node58634;
	wire [4-1:0] node58635;
	wire [4-1:0] node58636;
	wire [4-1:0] node58640;
	wire [4-1:0] node58643;
	wire [4-1:0] node58644;
	wire [4-1:0] node58645;
	wire [4-1:0] node58646;
	wire [4-1:0] node58647;
	wire [4-1:0] node58648;
	wire [4-1:0] node58649;
	wire [4-1:0] node58651;
	wire [4-1:0] node58654;
	wire [4-1:0] node58655;
	wire [4-1:0] node58658;
	wire [4-1:0] node58661;
	wire [4-1:0] node58662;
	wire [4-1:0] node58663;
	wire [4-1:0] node58665;
	wire [4-1:0] node58668;
	wire [4-1:0] node58669;
	wire [4-1:0] node58673;
	wire [4-1:0] node58674;
	wire [4-1:0] node58678;
	wire [4-1:0] node58679;
	wire [4-1:0] node58680;
	wire [4-1:0] node58681;
	wire [4-1:0] node58684;
	wire [4-1:0] node58687;
	wire [4-1:0] node58688;
	wire [4-1:0] node58691;
	wire [4-1:0] node58694;
	wire [4-1:0] node58695;
	wire [4-1:0] node58698;
	wire [4-1:0] node58701;
	wire [4-1:0] node58702;
	wire [4-1:0] node58703;
	wire [4-1:0] node58704;
	wire [4-1:0] node58705;
	wire [4-1:0] node58708;
	wire [4-1:0] node58711;
	wire [4-1:0] node58712;
	wire [4-1:0] node58715;
	wire [4-1:0] node58718;
	wire [4-1:0] node58719;
	wire [4-1:0] node58720;
	wire [4-1:0] node58723;
	wire [4-1:0] node58727;
	wire [4-1:0] node58728;
	wire [4-1:0] node58730;
	wire [4-1:0] node58731;
	wire [4-1:0] node58732;
	wire [4-1:0] node58736;
	wire [4-1:0] node58738;
	wire [4-1:0] node58741;
	wire [4-1:0] node58742;
	wire [4-1:0] node58743;
	wire [4-1:0] node58746;
	wire [4-1:0] node58749;
	wire [4-1:0] node58750;
	wire [4-1:0] node58753;
	wire [4-1:0] node58756;
	wire [4-1:0] node58757;
	wire [4-1:0] node58758;
	wire [4-1:0] node58759;
	wire [4-1:0] node58760;
	wire [4-1:0] node58761;
	wire [4-1:0] node58764;
	wire [4-1:0] node58767;
	wire [4-1:0] node58768;
	wire [4-1:0] node58771;
	wire [4-1:0] node58774;
	wire [4-1:0] node58775;
	wire [4-1:0] node58776;
	wire [4-1:0] node58777;
	wire [4-1:0] node58781;
	wire [4-1:0] node58782;
	wire [4-1:0] node58785;
	wire [4-1:0] node58788;
	wire [4-1:0] node58789;
	wire [4-1:0] node58793;
	wire [4-1:0] node58794;
	wire [4-1:0] node58795;
	wire [4-1:0] node58796;
	wire [4-1:0] node58797;
	wire [4-1:0] node58800;
	wire [4-1:0] node58803;
	wire [4-1:0] node58805;
	wire [4-1:0] node58808;
	wire [4-1:0] node58809;
	wire [4-1:0] node58811;
	wire [4-1:0] node58815;
	wire [4-1:0] node58816;
	wire [4-1:0] node58817;
	wire [4-1:0] node58820;
	wire [4-1:0] node58823;
	wire [4-1:0] node58824;
	wire [4-1:0] node58828;
	wire [4-1:0] node58829;
	wire [4-1:0] node58830;
	wire [4-1:0] node58831;
	wire [4-1:0] node58832;
	wire [4-1:0] node58835;
	wire [4-1:0] node58836;
	wire [4-1:0] node58840;
	wire [4-1:0] node58841;
	wire [4-1:0] node58844;
	wire [4-1:0] node58847;
	wire [4-1:0] node58849;
	wire [4-1:0] node58850;
	wire [4-1:0] node58853;
	wire [4-1:0] node58856;
	wire [4-1:0] node58857;
	wire [4-1:0] node58858;
	wire [4-1:0] node58860;
	wire [4-1:0] node58861;
	wire [4-1:0] node58864;
	wire [4-1:0] node58867;
	wire [4-1:0] node58869;
	wire [4-1:0] node58870;
	wire [4-1:0] node58873;
	wire [4-1:0] node58876;
	wire [4-1:0] node58877;
	wire [4-1:0] node58878;
	wire [4-1:0] node58881;
	wire [4-1:0] node58884;
	wire [4-1:0] node58886;
	wire [4-1:0] node58889;
	wire [4-1:0] node58890;
	wire [4-1:0] node58891;
	wire [4-1:0] node58892;
	wire [4-1:0] node58893;
	wire [4-1:0] node58894;
	wire [4-1:0] node58895;
	wire [4-1:0] node58896;
	wire [4-1:0] node58900;
	wire [4-1:0] node58901;
	wire [4-1:0] node58904;
	wire [4-1:0] node58907;
	wire [4-1:0] node58908;
	wire [4-1:0] node58909;
	wire [4-1:0] node58912;
	wire [4-1:0] node58915;
	wire [4-1:0] node58916;
	wire [4-1:0] node58920;
	wire [4-1:0] node58921;
	wire [4-1:0] node58923;
	wire [4-1:0] node58924;
	wire [4-1:0] node58927;
	wire [4-1:0] node58930;
	wire [4-1:0] node58931;
	wire [4-1:0] node58934;
	wire [4-1:0] node58935;
	wire [4-1:0] node58939;
	wire [4-1:0] node58940;
	wire [4-1:0] node58941;
	wire [4-1:0] node58942;
	wire [4-1:0] node58943;
	wire [4-1:0] node58946;
	wire [4-1:0] node58949;
	wire [4-1:0] node58950;
	wire [4-1:0] node58954;
	wire [4-1:0] node58955;
	wire [4-1:0] node58956;
	wire [4-1:0] node58959;
	wire [4-1:0] node58962;
	wire [4-1:0] node58963;
	wire [4-1:0] node58966;
	wire [4-1:0] node58969;
	wire [4-1:0] node58970;
	wire [4-1:0] node58971;
	wire [4-1:0] node58975;
	wire [4-1:0] node58976;
	wire [4-1:0] node58979;
	wire [4-1:0] node58982;
	wire [4-1:0] node58983;
	wire [4-1:0] node58984;
	wire [4-1:0] node58985;
	wire [4-1:0] node58986;
	wire [4-1:0] node58990;
	wire [4-1:0] node58993;
	wire [4-1:0] node58994;
	wire [4-1:0] node58995;
	wire [4-1:0] node58999;
	wire [4-1:0] node59002;
	wire [4-1:0] node59003;
	wire [4-1:0] node59004;
	wire [4-1:0] node59006;
	wire [4-1:0] node59009;
	wire [4-1:0] node59010;
	wire [4-1:0] node59011;
	wire [4-1:0] node59015;
	wire [4-1:0] node59018;
	wire [4-1:0] node59019;
	wire [4-1:0] node59020;
	wire [4-1:0] node59023;
	wire [4-1:0] node59026;
	wire [4-1:0] node59027;
	wire [4-1:0] node59028;
	wire [4-1:0] node59031;
	wire [4-1:0] node59034;
	wire [4-1:0] node59036;
	wire [4-1:0] node59039;
	wire [4-1:0] node59040;
	wire [4-1:0] node59041;
	wire [4-1:0] node59042;
	wire [4-1:0] node59043;
	wire [4-1:0] node59045;
	wire [4-1:0] node59048;
	wire [4-1:0] node59049;
	wire [4-1:0] node59050;
	wire [4-1:0] node59054;
	wire [4-1:0] node59057;
	wire [4-1:0] node59058;
	wire [4-1:0] node59059;
	wire [4-1:0] node59060;
	wire [4-1:0] node59063;
	wire [4-1:0] node59066;
	wire [4-1:0] node59067;
	wire [4-1:0] node59070;
	wire [4-1:0] node59073;
	wire [4-1:0] node59074;
	wire [4-1:0] node59075;
	wire [4-1:0] node59079;
	wire [4-1:0] node59082;
	wire [4-1:0] node59083;
	wire [4-1:0] node59084;
	wire [4-1:0] node59085;
	wire [4-1:0] node59086;
	wire [4-1:0] node59090;
	wire [4-1:0] node59093;
	wire [4-1:0] node59095;
	wire [4-1:0] node59096;
	wire [4-1:0] node59100;
	wire [4-1:0] node59102;
	wire [4-1:0] node59103;
	wire [4-1:0] node59104;
	wire [4-1:0] node59108;
	wire [4-1:0] node59111;
	wire [4-1:0] node59112;
	wire [4-1:0] node59113;
	wire [4-1:0] node59114;
	wire [4-1:0] node59115;
	wire [4-1:0] node59118;
	wire [4-1:0] node59119;
	wire [4-1:0] node59123;
	wire [4-1:0] node59124;
	wire [4-1:0] node59125;
	wire [4-1:0] node59128;
	wire [4-1:0] node59132;
	wire [4-1:0] node59133;
	wire [4-1:0] node59134;
	wire [4-1:0] node59135;
	wire [4-1:0] node59138;
	wire [4-1:0] node59141;
	wire [4-1:0] node59142;
	wire [4-1:0] node59145;
	wire [4-1:0] node59148;
	wire [4-1:0] node59149;
	wire [4-1:0] node59152;
	wire [4-1:0] node59155;
	wire [4-1:0] node59156;
	wire [4-1:0] node59157;
	wire [4-1:0] node59158;
	wire [4-1:0] node59162;
	wire [4-1:0] node59163;
	wire [4-1:0] node59167;
	wire [4-1:0] node59168;
	wire [4-1:0] node59169;
	wire [4-1:0] node59173;
	wire [4-1:0] node59174;
	wire [4-1:0] node59178;
	wire [4-1:0] node59179;
	wire [4-1:0] node59180;
	wire [4-1:0] node59181;
	wire [4-1:0] node59182;
	wire [4-1:0] node59183;
	wire [4-1:0] node59184;
	wire [4-1:0] node59185;
	wire [4-1:0] node59186;
	wire [4-1:0] node59187;
	wire [4-1:0] node59190;
	wire [4-1:0] node59194;
	wire [4-1:0] node59195;
	wire [4-1:0] node59199;
	wire [4-1:0] node59200;
	wire [4-1:0] node59201;
	wire [4-1:0] node59202;
	wire [4-1:0] node59206;
	wire [4-1:0] node59209;
	wire [4-1:0] node59210;
	wire [4-1:0] node59213;
	wire [4-1:0] node59214;
	wire [4-1:0] node59218;
	wire [4-1:0] node59219;
	wire [4-1:0] node59220;
	wire [4-1:0] node59221;
	wire [4-1:0] node59224;
	wire [4-1:0] node59227;
	wire [4-1:0] node59228;
	wire [4-1:0] node59231;
	wire [4-1:0] node59234;
	wire [4-1:0] node59235;
	wire [4-1:0] node59236;
	wire [4-1:0] node59237;
	wire [4-1:0] node59240;
	wire [4-1:0] node59243;
	wire [4-1:0] node59244;
	wire [4-1:0] node59247;
	wire [4-1:0] node59250;
	wire [4-1:0] node59252;
	wire [4-1:0] node59255;
	wire [4-1:0] node59256;
	wire [4-1:0] node59257;
	wire [4-1:0] node59258;
	wire [4-1:0] node59260;
	wire [4-1:0] node59261;
	wire [4-1:0] node59264;
	wire [4-1:0] node59267;
	wire [4-1:0] node59268;
	wire [4-1:0] node59271;
	wire [4-1:0] node59274;
	wire [4-1:0] node59275;
	wire [4-1:0] node59276;
	wire [4-1:0] node59280;
	wire [4-1:0] node59282;
	wire [4-1:0] node59285;
	wire [4-1:0] node59286;
	wire [4-1:0] node59287;
	wire [4-1:0] node59289;
	wire [4-1:0] node59292;
	wire [4-1:0] node59293;
	wire [4-1:0] node59294;
	wire [4-1:0] node59299;
	wire [4-1:0] node59301;
	wire [4-1:0] node59302;
	wire [4-1:0] node59306;
	wire [4-1:0] node59307;
	wire [4-1:0] node59308;
	wire [4-1:0] node59309;
	wire [4-1:0] node59310;
	wire [4-1:0] node59311;
	wire [4-1:0] node59312;
	wire [4-1:0] node59315;
	wire [4-1:0] node59319;
	wire [4-1:0] node59320;
	wire [4-1:0] node59322;
	wire [4-1:0] node59325;
	wire [4-1:0] node59326;
	wire [4-1:0] node59329;
	wire [4-1:0] node59332;
	wire [4-1:0] node59333;
	wire [4-1:0] node59335;
	wire [4-1:0] node59338;
	wire [4-1:0] node59339;
	wire [4-1:0] node59342;
	wire [4-1:0] node59345;
	wire [4-1:0] node59346;
	wire [4-1:0] node59347;
	wire [4-1:0] node59348;
	wire [4-1:0] node59349;
	wire [4-1:0] node59353;
	wire [4-1:0] node59354;
	wire [4-1:0] node59357;
	wire [4-1:0] node59360;
	wire [4-1:0] node59361;
	wire [4-1:0] node59362;
	wire [4-1:0] node59366;
	wire [4-1:0] node59367;
	wire [4-1:0] node59370;
	wire [4-1:0] node59373;
	wire [4-1:0] node59374;
	wire [4-1:0] node59377;
	wire [4-1:0] node59378;
	wire [4-1:0] node59381;
	wire [4-1:0] node59384;
	wire [4-1:0] node59385;
	wire [4-1:0] node59386;
	wire [4-1:0] node59387;
	wire [4-1:0] node59388;
	wire [4-1:0] node59392;
	wire [4-1:0] node59393;
	wire [4-1:0] node59394;
	wire [4-1:0] node59397;
	wire [4-1:0] node59401;
	wire [4-1:0] node59402;
	wire [4-1:0] node59403;
	wire [4-1:0] node59406;
	wire [4-1:0] node59409;
	wire [4-1:0] node59410;
	wire [4-1:0] node59411;
	wire [4-1:0] node59414;
	wire [4-1:0] node59418;
	wire [4-1:0] node59419;
	wire [4-1:0] node59420;
	wire [4-1:0] node59422;
	wire [4-1:0] node59423;
	wire [4-1:0] node59426;
	wire [4-1:0] node59429;
	wire [4-1:0] node59431;
	wire [4-1:0] node59434;
	wire [4-1:0] node59435;
	wire [4-1:0] node59436;
	wire [4-1:0] node59438;
	wire [4-1:0] node59441;
	wire [4-1:0] node59442;
	wire [4-1:0] node59445;
	wire [4-1:0] node59448;
	wire [4-1:0] node59449;
	wire [4-1:0] node59450;
	wire [4-1:0] node59455;
	wire [4-1:0] node59456;
	wire [4-1:0] node59457;
	wire [4-1:0] node59458;
	wire [4-1:0] node59459;
	wire [4-1:0] node59460;
	wire [4-1:0] node59461;
	wire [4-1:0] node59463;
	wire [4-1:0] node59466;
	wire [4-1:0] node59467;
	wire [4-1:0] node59471;
	wire [4-1:0] node59472;
	wire [4-1:0] node59473;
	wire [4-1:0] node59476;
	wire [4-1:0] node59480;
	wire [4-1:0] node59481;
	wire [4-1:0] node59482;
	wire [4-1:0] node59485;
	wire [4-1:0] node59488;
	wire [4-1:0] node59490;
	wire [4-1:0] node59491;
	wire [4-1:0] node59494;
	wire [4-1:0] node59497;
	wire [4-1:0] node59498;
	wire [4-1:0] node59499;
	wire [4-1:0] node59502;
	wire [4-1:0] node59503;
	wire [4-1:0] node59506;
	wire [4-1:0] node59509;
	wire [4-1:0] node59510;
	wire [4-1:0] node59512;
	wire [4-1:0] node59515;
	wire [4-1:0] node59517;
	wire [4-1:0] node59520;
	wire [4-1:0] node59521;
	wire [4-1:0] node59522;
	wire [4-1:0] node59523;
	wire [4-1:0] node59524;
	wire [4-1:0] node59528;
	wire [4-1:0] node59529;
	wire [4-1:0] node59532;
	wire [4-1:0] node59534;
	wire [4-1:0] node59537;
	wire [4-1:0] node59538;
	wire [4-1:0] node59539;
	wire [4-1:0] node59540;
	wire [4-1:0] node59543;
	wire [4-1:0] node59547;
	wire [4-1:0] node59549;
	wire [4-1:0] node59552;
	wire [4-1:0] node59553;
	wire [4-1:0] node59555;
	wire [4-1:0] node59556;
	wire [4-1:0] node59559;
	wire [4-1:0] node59562;
	wire [4-1:0] node59563;
	wire [4-1:0] node59566;
	wire [4-1:0] node59569;
	wire [4-1:0] node59570;
	wire [4-1:0] node59571;
	wire [4-1:0] node59572;
	wire [4-1:0] node59573;
	wire [4-1:0] node59575;
	wire [4-1:0] node59576;
	wire [4-1:0] node59579;
	wire [4-1:0] node59582;
	wire [4-1:0] node59583;
	wire [4-1:0] node59585;
	wire [4-1:0] node59588;
	wire [4-1:0] node59590;
	wire [4-1:0] node59593;
	wire [4-1:0] node59594;
	wire [4-1:0] node59597;
	wire [4-1:0] node59598;
	wire [4-1:0] node59599;
	wire [4-1:0] node59603;
	wire [4-1:0] node59604;
	wire [4-1:0] node59608;
	wire [4-1:0] node59609;
	wire [4-1:0] node59610;
	wire [4-1:0] node59612;
	wire [4-1:0] node59615;
	wire [4-1:0] node59616;
	wire [4-1:0] node59619;
	wire [4-1:0] node59622;
	wire [4-1:0] node59623;
	wire [4-1:0] node59624;
	wire [4-1:0] node59627;
	wire [4-1:0] node59630;
	wire [4-1:0] node59631;
	wire [4-1:0] node59634;
	wire [4-1:0] node59637;
	wire [4-1:0] node59638;
	wire [4-1:0] node59639;
	wire [4-1:0] node59640;
	wire [4-1:0] node59642;
	wire [4-1:0] node59645;
	wire [4-1:0] node59646;
	wire [4-1:0] node59647;
	wire [4-1:0] node59651;
	wire [4-1:0] node59654;
	wire [4-1:0] node59655;
	wire [4-1:0] node59656;
	wire [4-1:0] node59657;
	wire [4-1:0] node59661;
	wire [4-1:0] node59662;
	wire [4-1:0] node59666;
	wire [4-1:0] node59668;
	wire [4-1:0] node59671;
	wire [4-1:0] node59672;
	wire [4-1:0] node59673;
	wire [4-1:0] node59674;
	wire [4-1:0] node59678;
	wire [4-1:0] node59679;
	wire [4-1:0] node59682;
	wire [4-1:0] node59685;
	wire [4-1:0] node59686;
	wire [4-1:0] node59687;
	wire [4-1:0] node59689;
	wire [4-1:0] node59692;
	wire [4-1:0] node59695;
	wire [4-1:0] node59697;
	wire [4-1:0] node59700;
	wire [4-1:0] node59701;
	wire [4-1:0] node59702;
	wire [4-1:0] node59703;
	wire [4-1:0] node59704;
	wire [4-1:0] node59705;
	wire [4-1:0] node59706;
	wire [4-1:0] node59707;
	wire [4-1:0] node59710;
	wire [4-1:0] node59713;
	wire [4-1:0] node59714;
	wire [4-1:0] node59717;
	wire [4-1:0] node59720;
	wire [4-1:0] node59721;
	wire [4-1:0] node59723;
	wire [4-1:0] node59726;
	wire [4-1:0] node59727;
	wire [4-1:0] node59730;
	wire [4-1:0] node59733;
	wire [4-1:0] node59734;
	wire [4-1:0] node59735;
	wire [4-1:0] node59736;
	wire [4-1:0] node59739;
	wire [4-1:0] node59742;
	wire [4-1:0] node59743;
	wire [4-1:0] node59744;
	wire [4-1:0] node59747;
	wire [4-1:0] node59751;
	wire [4-1:0] node59752;
	wire [4-1:0] node59756;
	wire [4-1:0] node59757;
	wire [4-1:0] node59758;
	wire [4-1:0] node59759;
	wire [4-1:0] node59760;
	wire [4-1:0] node59763;
	wire [4-1:0] node59767;
	wire [4-1:0] node59769;
	wire [4-1:0] node59770;
	wire [4-1:0] node59771;
	wire [4-1:0] node59774;
	wire [4-1:0] node59777;
	wire [4-1:0] node59779;
	wire [4-1:0] node59782;
	wire [4-1:0] node59783;
	wire [4-1:0] node59784;
	wire [4-1:0] node59785;
	wire [4-1:0] node59788;
	wire [4-1:0] node59791;
	wire [4-1:0] node59793;
	wire [4-1:0] node59796;
	wire [4-1:0] node59797;
	wire [4-1:0] node59800;
	wire [4-1:0] node59803;
	wire [4-1:0] node59804;
	wire [4-1:0] node59805;
	wire [4-1:0] node59806;
	wire [4-1:0] node59807;
	wire [4-1:0] node59810;
	wire [4-1:0] node59813;
	wire [4-1:0] node59814;
	wire [4-1:0] node59816;
	wire [4-1:0] node59819;
	wire [4-1:0] node59820;
	wire [4-1:0] node59823;
	wire [4-1:0] node59825;
	wire [4-1:0] node59828;
	wire [4-1:0] node59829;
	wire [4-1:0] node59830;
	wire [4-1:0] node59831;
	wire [4-1:0] node59832;
	wire [4-1:0] node59835;
	wire [4-1:0] node59839;
	wire [4-1:0] node59841;
	wire [4-1:0] node59843;
	wire [4-1:0] node59846;
	wire [4-1:0] node59847;
	wire [4-1:0] node59848;
	wire [4-1:0] node59852;
	wire [4-1:0] node59853;
	wire [4-1:0] node59856;
	wire [4-1:0] node59859;
	wire [4-1:0] node59860;
	wire [4-1:0] node59861;
	wire [4-1:0] node59862;
	wire [4-1:0] node59863;
	wire [4-1:0] node59864;
	wire [4-1:0] node59867;
	wire [4-1:0] node59870;
	wire [4-1:0] node59871;
	wire [4-1:0] node59874;
	wire [4-1:0] node59877;
	wire [4-1:0] node59878;
	wire [4-1:0] node59879;
	wire [4-1:0] node59882;
	wire [4-1:0] node59885;
	wire [4-1:0] node59886;
	wire [4-1:0] node59890;
	wire [4-1:0] node59891;
	wire [4-1:0] node59892;
	wire [4-1:0] node59895;
	wire [4-1:0] node59898;
	wire [4-1:0] node59899;
	wire [4-1:0] node59902;
	wire [4-1:0] node59905;
	wire [4-1:0] node59906;
	wire [4-1:0] node59907;
	wire [4-1:0] node59908;
	wire [4-1:0] node59909;
	wire [4-1:0] node59913;
	wire [4-1:0] node59914;
	wire [4-1:0] node59917;
	wire [4-1:0] node59920;
	wire [4-1:0] node59921;
	wire [4-1:0] node59922;
	wire [4-1:0] node59926;
	wire [4-1:0] node59927;
	wire [4-1:0] node59930;
	wire [4-1:0] node59933;
	wire [4-1:0] node59934;
	wire [4-1:0] node59935;
	wire [4-1:0] node59938;
	wire [4-1:0] node59941;
	wire [4-1:0] node59942;
	wire [4-1:0] node59945;
	wire [4-1:0] node59948;
	wire [4-1:0] node59949;
	wire [4-1:0] node59950;
	wire [4-1:0] node59951;
	wire [4-1:0] node59952;
	wire [4-1:0] node59953;
	wire [4-1:0] node59954;
	wire [4-1:0] node59958;
	wire [4-1:0] node59959;
	wire [4-1:0] node59963;
	wire [4-1:0] node59964;
	wire [4-1:0] node59965;
	wire [4-1:0] node59969;
	wire [4-1:0] node59970;
	wire [4-1:0] node59974;
	wire [4-1:0] node59975;
	wire [4-1:0] node59976;
	wire [4-1:0] node59977;
	wire [4-1:0] node59978;
	wire [4-1:0] node59981;
	wire [4-1:0] node59985;
	wire [4-1:0] node59986;
	wire [4-1:0] node59987;
	wire [4-1:0] node59991;
	wire [4-1:0] node59994;
	wire [4-1:0] node59995;
	wire [4-1:0] node59996;
	wire [4-1:0] node59999;
	wire [4-1:0] node60000;
	wire [4-1:0] node60004;
	wire [4-1:0] node60006;
	wire [4-1:0] node60009;
	wire [4-1:0] node60010;
	wire [4-1:0] node60011;
	wire [4-1:0] node60013;
	wire [4-1:0] node60014;
	wire [4-1:0] node60018;
	wire [4-1:0] node60019;
	wire [4-1:0] node60020;
	wire [4-1:0] node60024;
	wire [4-1:0] node60025;
	wire [4-1:0] node60029;
	wire [4-1:0] node60030;
	wire [4-1:0] node60031;
	wire [4-1:0] node60032;
	wire [4-1:0] node60035;
	wire [4-1:0] node60038;
	wire [4-1:0] node60039;
	wire [4-1:0] node60040;
	wire [4-1:0] node60044;
	wire [4-1:0] node60047;
	wire [4-1:0] node60048;
	wire [4-1:0] node60051;
	wire [4-1:0] node60054;
	wire [4-1:0] node60055;
	wire [4-1:0] node60056;
	wire [4-1:0] node60057;
	wire [4-1:0] node60058;
	wire [4-1:0] node60059;
	wire [4-1:0] node60063;
	wire [4-1:0] node60064;
	wire [4-1:0] node60068;
	wire [4-1:0] node60069;
	wire [4-1:0] node60070;
	wire [4-1:0] node60074;
	wire [4-1:0] node60075;
	wire [4-1:0] node60079;
	wire [4-1:0] node60080;
	wire [4-1:0] node60081;
	wire [4-1:0] node60082;
	wire [4-1:0] node60085;
	wire [4-1:0] node60088;
	wire [4-1:0] node60090;
	wire [4-1:0] node60093;
	wire [4-1:0] node60094;
	wire [4-1:0] node60097;
	wire [4-1:0] node60100;
	wire [4-1:0] node60101;
	wire [4-1:0] node60102;
	wire [4-1:0] node60103;
	wire [4-1:0] node60106;
	wire [4-1:0] node60107;
	wire [4-1:0] node60111;
	wire [4-1:0] node60112;
	wire [4-1:0] node60113;
	wire [4-1:0] node60117;
	wire [4-1:0] node60118;
	wire [4-1:0] node60122;
	wire [4-1:0] node60123;
	wire [4-1:0] node60124;
	wire [4-1:0] node60125;
	wire [4-1:0] node60129;
	wire [4-1:0] node60130;
	wire [4-1:0] node60134;
	wire [4-1:0] node60135;
	wire [4-1:0] node60138;
	wire [4-1:0] node60139;
	wire [4-1:0] node60143;
	wire [4-1:0] node60144;
	wire [4-1:0] node60145;
	wire [4-1:0] node60146;
	wire [4-1:0] node60147;
	wire [4-1:0] node60148;
	wire [4-1:0] node60149;
	wire [4-1:0] node60150;
	wire [4-1:0] node60151;
	wire [4-1:0] node60152;
	wire [4-1:0] node60155;
	wire [4-1:0] node60156;
	wire [4-1:0] node60160;
	wire [4-1:0] node60162;
	wire [4-1:0] node60163;
	wire [4-1:0] node60167;
	wire [4-1:0] node60168;
	wire [4-1:0] node60169;
	wire [4-1:0] node60170;
	wire [4-1:0] node60174;
	wire [4-1:0] node60175;
	wire [4-1:0] node60179;
	wire [4-1:0] node60181;
	wire [4-1:0] node60184;
	wire [4-1:0] node60185;
	wire [4-1:0] node60186;
	wire [4-1:0] node60187;
	wire [4-1:0] node60188;
	wire [4-1:0] node60193;
	wire [4-1:0] node60194;
	wire [4-1:0] node60195;
	wire [4-1:0] node60199;
	wire [4-1:0] node60200;
	wire [4-1:0] node60204;
	wire [4-1:0] node60205;
	wire [4-1:0] node60206;
	wire [4-1:0] node60207;
	wire [4-1:0] node60212;
	wire [4-1:0] node60213;
	wire [4-1:0] node60216;
	wire [4-1:0] node60217;
	wire [4-1:0] node60221;
	wire [4-1:0] node60222;
	wire [4-1:0] node60223;
	wire [4-1:0] node60224;
	wire [4-1:0] node60225;
	wire [4-1:0] node60227;
	wire [4-1:0] node60230;
	wire [4-1:0] node60231;
	wire [4-1:0] node60234;
	wire [4-1:0] node60237;
	wire [4-1:0] node60238;
	wire [4-1:0] node60240;
	wire [4-1:0] node60243;
	wire [4-1:0] node60244;
	wire [4-1:0] node60248;
	wire [4-1:0] node60249;
	wire [4-1:0] node60250;
	wire [4-1:0] node60251;
	wire [4-1:0] node60255;
	wire [4-1:0] node60258;
	wire [4-1:0] node60260;
	wire [4-1:0] node60263;
	wire [4-1:0] node60264;
	wire [4-1:0] node60265;
	wire [4-1:0] node60267;
	wire [4-1:0] node60268;
	wire [4-1:0] node60272;
	wire [4-1:0] node60273;
	wire [4-1:0] node60274;
	wire [4-1:0] node60278;
	wire [4-1:0] node60279;
	wire [4-1:0] node60283;
	wire [4-1:0] node60284;
	wire [4-1:0] node60285;
	wire [4-1:0] node60288;
	wire [4-1:0] node60289;
	wire [4-1:0] node60293;
	wire [4-1:0] node60294;
	wire [4-1:0] node60295;
	wire [4-1:0] node60299;
	wire [4-1:0] node60300;
	wire [4-1:0] node60304;
	wire [4-1:0] node60305;
	wire [4-1:0] node60306;
	wire [4-1:0] node60307;
	wire [4-1:0] node60308;
	wire [4-1:0] node60309;
	wire [4-1:0] node60310;
	wire [4-1:0] node60315;
	wire [4-1:0] node60316;
	wire [4-1:0] node60317;
	wire [4-1:0] node60321;
	wire [4-1:0] node60322;
	wire [4-1:0] node60326;
	wire [4-1:0] node60327;
	wire [4-1:0] node60328;
	wire [4-1:0] node60330;
	wire [4-1:0] node60333;
	wire [4-1:0] node60334;
	wire [4-1:0] node60337;
	wire [4-1:0] node60340;
	wire [4-1:0] node60342;
	wire [4-1:0] node60345;
	wire [4-1:0] node60346;
	wire [4-1:0] node60347;
	wire [4-1:0] node60350;
	wire [4-1:0] node60352;
	wire [4-1:0] node60355;
	wire [4-1:0] node60356;
	wire [4-1:0] node60357;
	wire [4-1:0] node60359;
	wire [4-1:0] node60362;
	wire [4-1:0] node60363;
	wire [4-1:0] node60366;
	wire [4-1:0] node60369;
	wire [4-1:0] node60370;
	wire [4-1:0] node60371;
	wire [4-1:0] node60374;
	wire [4-1:0] node60378;
	wire [4-1:0] node60379;
	wire [4-1:0] node60380;
	wire [4-1:0] node60381;
	wire [4-1:0] node60382;
	wire [4-1:0] node60383;
	wire [4-1:0] node60387;
	wire [4-1:0] node60388;
	wire [4-1:0] node60391;
	wire [4-1:0] node60394;
	wire [4-1:0] node60395;
	wire [4-1:0] node60398;
	wire [4-1:0] node60401;
	wire [4-1:0] node60402;
	wire [4-1:0] node60403;
	wire [4-1:0] node60404;
	wire [4-1:0] node60408;
	wire [4-1:0] node60411;
	wire [4-1:0] node60412;
	wire [4-1:0] node60413;
	wire [4-1:0] node60417;
	wire [4-1:0] node60418;
	wire [4-1:0] node60422;
	wire [4-1:0] node60423;
	wire [4-1:0] node60424;
	wire [4-1:0] node60427;
	wire [4-1:0] node60430;
	wire [4-1:0] node60431;
	wire [4-1:0] node60432;
	wire [4-1:0] node60433;
	wire [4-1:0] node60436;
	wire [4-1:0] node60440;
	wire [4-1:0] node60441;
	wire [4-1:0] node60444;
	wire [4-1:0] node60447;
	wire [4-1:0] node60448;
	wire [4-1:0] node60449;
	wire [4-1:0] node60450;
	wire [4-1:0] node60451;
	wire [4-1:0] node60452;
	wire [4-1:0] node60454;
	wire [4-1:0] node60456;
	wire [4-1:0] node60459;
	wire [4-1:0] node60460;
	wire [4-1:0] node60462;
	wire [4-1:0] node60465;
	wire [4-1:0] node60468;
	wire [4-1:0] node60469;
	wire [4-1:0] node60470;
	wire [4-1:0] node60471;
	wire [4-1:0] node60475;
	wire [4-1:0] node60477;
	wire [4-1:0] node60480;
	wire [4-1:0] node60482;
	wire [4-1:0] node60483;
	wire [4-1:0] node60486;
	wire [4-1:0] node60489;
	wire [4-1:0] node60490;
	wire [4-1:0] node60491;
	wire [4-1:0] node60493;
	wire [4-1:0] node60496;
	wire [4-1:0] node60498;
	wire [4-1:0] node60501;
	wire [4-1:0] node60502;
	wire [4-1:0] node60504;
	wire [4-1:0] node60507;
	wire [4-1:0] node60509;
	wire [4-1:0] node60512;
	wire [4-1:0] node60513;
	wire [4-1:0] node60514;
	wire [4-1:0] node60515;
	wire [4-1:0] node60516;
	wire [4-1:0] node60518;
	wire [4-1:0] node60521;
	wire [4-1:0] node60524;
	wire [4-1:0] node60525;
	wire [4-1:0] node60527;
	wire [4-1:0] node60530;
	wire [4-1:0] node60533;
	wire [4-1:0] node60534;
	wire [4-1:0] node60535;
	wire [4-1:0] node60536;
	wire [4-1:0] node60541;
	wire [4-1:0] node60542;
	wire [4-1:0] node60543;
	wire [4-1:0] node60547;
	wire [4-1:0] node60548;
	wire [4-1:0] node60552;
	wire [4-1:0] node60553;
	wire [4-1:0] node60554;
	wire [4-1:0] node60555;
	wire [4-1:0] node60559;
	wire [4-1:0] node60560;
	wire [4-1:0] node60564;
	wire [4-1:0] node60565;
	wire [4-1:0] node60566;
	wire [4-1:0] node60570;
	wire [4-1:0] node60571;
	wire [4-1:0] node60575;
	wire [4-1:0] node60576;
	wire [4-1:0] node60577;
	wire [4-1:0] node60578;
	wire [4-1:0] node60579;
	wire [4-1:0] node60581;
	wire [4-1:0] node60584;
	wire [4-1:0] node60586;
	wire [4-1:0] node60588;
	wire [4-1:0] node60591;
	wire [4-1:0] node60592;
	wire [4-1:0] node60594;
	wire [4-1:0] node60595;
	wire [4-1:0] node60600;
	wire [4-1:0] node60601;
	wire [4-1:0] node60602;
	wire [4-1:0] node60603;
	wire [4-1:0] node60605;
	wire [4-1:0] node60608;
	wire [4-1:0] node60609;
	wire [4-1:0] node60612;
	wire [4-1:0] node60616;
	wire [4-1:0] node60617;
	wire [4-1:0] node60618;
	wire [4-1:0] node60619;
	wire [4-1:0] node60622;
	wire [4-1:0] node60625;
	wire [4-1:0] node60626;
	wire [4-1:0] node60629;
	wire [4-1:0] node60632;
	wire [4-1:0] node60633;
	wire [4-1:0] node60637;
	wire [4-1:0] node60638;
	wire [4-1:0] node60639;
	wire [4-1:0] node60640;
	wire [4-1:0] node60643;
	wire [4-1:0] node60644;
	wire [4-1:0] node60645;
	wire [4-1:0] node60649;
	wire [4-1:0] node60650;
	wire [4-1:0] node60654;
	wire [4-1:0] node60655;
	wire [4-1:0] node60657;
	wire [4-1:0] node60660;
	wire [4-1:0] node60661;
	wire [4-1:0] node60662;
	wire [4-1:0] node60667;
	wire [4-1:0] node60668;
	wire [4-1:0] node60669;
	wire [4-1:0] node60670;
	wire [4-1:0] node60674;
	wire [4-1:0] node60675;
	wire [4-1:0] node60679;
	wire [4-1:0] node60680;
	wire [4-1:0] node60681;
	wire [4-1:0] node60685;
	wire [4-1:0] node60686;
	wire [4-1:0] node60690;
	wire [4-1:0] node60691;
	wire [4-1:0] node60692;
	wire [4-1:0] node60693;
	wire [4-1:0] node60694;
	wire [4-1:0] node60695;
	wire [4-1:0] node60696;
	wire [4-1:0] node60697;
	wire [4-1:0] node60700;
	wire [4-1:0] node60703;
	wire [4-1:0] node60704;
	wire [4-1:0] node60707;
	wire [4-1:0] node60710;
	wire [4-1:0] node60711;
	wire [4-1:0] node60712;
	wire [4-1:0] node60713;
	wire [4-1:0] node60716;
	wire [4-1:0] node60720;
	wire [4-1:0] node60721;
	wire [4-1:0] node60724;
	wire [4-1:0] node60727;
	wire [4-1:0] node60728;
	wire [4-1:0] node60729;
	wire [4-1:0] node60730;
	wire [4-1:0] node60733;
	wire [4-1:0] node60736;
	wire [4-1:0] node60738;
	wire [4-1:0] node60741;
	wire [4-1:0] node60742;
	wire [4-1:0] node60743;
	wire [4-1:0] node60746;
	wire [4-1:0] node60749;
	wire [4-1:0] node60750;
	wire [4-1:0] node60753;
	wire [4-1:0] node60756;
	wire [4-1:0] node60757;
	wire [4-1:0] node60758;
	wire [4-1:0] node60759;
	wire [4-1:0] node60760;
	wire [4-1:0] node60761;
	wire [4-1:0] node60764;
	wire [4-1:0] node60767;
	wire [4-1:0] node60769;
	wire [4-1:0] node60772;
	wire [4-1:0] node60773;
	wire [4-1:0] node60776;
	wire [4-1:0] node60779;
	wire [4-1:0] node60780;
	wire [4-1:0] node60781;
	wire [4-1:0] node60784;
	wire [4-1:0] node60787;
	wire [4-1:0] node60788;
	wire [4-1:0] node60791;
	wire [4-1:0] node60794;
	wire [4-1:0] node60795;
	wire [4-1:0] node60796;
	wire [4-1:0] node60797;
	wire [4-1:0] node60801;
	wire [4-1:0] node60802;
	wire [4-1:0] node60805;
	wire [4-1:0] node60808;
	wire [4-1:0] node60809;
	wire [4-1:0] node60810;
	wire [4-1:0] node60813;
	wire [4-1:0] node60816;
	wire [4-1:0] node60817;
	wire [4-1:0] node60820;
	wire [4-1:0] node60823;
	wire [4-1:0] node60824;
	wire [4-1:0] node60825;
	wire [4-1:0] node60826;
	wire [4-1:0] node60829;
	wire [4-1:0] node60832;
	wire [4-1:0] node60833;
	wire [4-1:0] node60834;
	wire [4-1:0] node60835;
	wire [4-1:0] node60838;
	wire [4-1:0] node60841;
	wire [4-1:0] node60842;
	wire [4-1:0] node60845;
	wire [4-1:0] node60848;
	wire [4-1:0] node60849;
	wire [4-1:0] node60850;
	wire [4-1:0] node60851;
	wire [4-1:0] node60854;
	wire [4-1:0] node60857;
	wire [4-1:0] node60858;
	wire [4-1:0] node60861;
	wire [4-1:0] node60864;
	wire [4-1:0] node60865;
	wire [4-1:0] node60868;
	wire [4-1:0] node60871;
	wire [4-1:0] node60872;
	wire [4-1:0] node60873;
	wire [4-1:0] node60874;
	wire [4-1:0] node60875;
	wire [4-1:0] node60876;
	wire [4-1:0] node60881;
	wire [4-1:0] node60882;
	wire [4-1:0] node60883;
	wire [4-1:0] node60886;
	wire [4-1:0] node60889;
	wire [4-1:0] node60890;
	wire [4-1:0] node60893;
	wire [4-1:0] node60896;
	wire [4-1:0] node60897;
	wire [4-1:0] node60900;
	wire [4-1:0] node60903;
	wire [4-1:0] node60904;
	wire [4-1:0] node60905;
	wire [4-1:0] node60906;
	wire [4-1:0] node60909;
	wire [4-1:0] node60913;
	wire [4-1:0] node60914;
	wire [4-1:0] node60917;
	wire [4-1:0] node60920;
	wire [4-1:0] node60921;
	wire [4-1:0] node60922;
	wire [4-1:0] node60923;
	wire [4-1:0] node60924;
	wire [4-1:0] node60926;
	wire [4-1:0] node60927;
	wire [4-1:0] node60931;
	wire [4-1:0] node60932;
	wire [4-1:0] node60933;
	wire [4-1:0] node60938;
	wire [4-1:0] node60939;
	wire [4-1:0] node60940;
	wire [4-1:0] node60944;
	wire [4-1:0] node60945;
	wire [4-1:0] node60949;
	wire [4-1:0] node60950;
	wire [4-1:0] node60951;
	wire [4-1:0] node60952;
	wire [4-1:0] node60953;
	wire [4-1:0] node60957;
	wire [4-1:0] node60958;
	wire [4-1:0] node60962;
	wire [4-1:0] node60963;
	wire [4-1:0] node60964;
	wire [4-1:0] node60968;
	wire [4-1:0] node60969;
	wire [4-1:0] node60973;
	wire [4-1:0] node60974;
	wire [4-1:0] node60975;
	wire [4-1:0] node60976;
	wire [4-1:0] node60978;
	wire [4-1:0] node60981;
	wire [4-1:0] node60983;
	wire [4-1:0] node60986;
	wire [4-1:0] node60987;
	wire [4-1:0] node60991;
	wire [4-1:0] node60992;
	wire [4-1:0] node60993;
	wire [4-1:0] node60994;
	wire [4-1:0] node60998;
	wire [4-1:0] node60999;
	wire [4-1:0] node61003;
	wire [4-1:0] node61004;
	wire [4-1:0] node61005;
	wire [4-1:0] node61009;
	wire [4-1:0] node61012;
	wire [4-1:0] node61013;
	wire [4-1:0] node61014;
	wire [4-1:0] node61015;
	wire [4-1:0] node61016;
	wire [4-1:0] node61017;
	wire [4-1:0] node61021;
	wire [4-1:0] node61022;
	wire [4-1:0] node61026;
	wire [4-1:0] node61027;
	wire [4-1:0] node61028;
	wire [4-1:0] node61032;
	wire [4-1:0] node61033;
	wire [4-1:0] node61037;
	wire [4-1:0] node61038;
	wire [4-1:0] node61039;
	wire [4-1:0] node61040;
	wire [4-1:0] node61041;
	wire [4-1:0] node61046;
	wire [4-1:0] node61047;
	wire [4-1:0] node61049;
	wire [4-1:0] node61052;
	wire [4-1:0] node61055;
	wire [4-1:0] node61056;
	wire [4-1:0] node61058;
	wire [4-1:0] node61059;
	wire [4-1:0] node61062;
	wire [4-1:0] node61065;
	wire [4-1:0] node61067;
	wire [4-1:0] node61068;
	wire [4-1:0] node61071;
	wire [4-1:0] node61074;
	wire [4-1:0] node61075;
	wire [4-1:0] node61076;
	wire [4-1:0] node61077;
	wire [4-1:0] node61079;
	wire [4-1:0] node61083;
	wire [4-1:0] node61085;
	wire [4-1:0] node61086;
	wire [4-1:0] node61090;
	wire [4-1:0] node61091;
	wire [4-1:0] node61092;
	wire [4-1:0] node61093;
	wire [4-1:0] node61097;
	wire [4-1:0] node61098;
	wire [4-1:0] node61102;
	wire [4-1:0] node61103;
	wire [4-1:0] node61104;
	wire [4-1:0] node61108;
	wire [4-1:0] node61109;
	wire [4-1:0] node61113;
	wire [4-1:0] node61114;
	wire [4-1:0] node61115;
	wire [4-1:0] node61116;
	wire [4-1:0] node61117;
	wire [4-1:0] node61118;
	wire [4-1:0] node61119;
	wire [4-1:0] node61120;
	wire [4-1:0] node61121;
	wire [4-1:0] node61124;
	wire [4-1:0] node61127;
	wire [4-1:0] node61128;
	wire [4-1:0] node61132;
	wire [4-1:0] node61133;
	wire [4-1:0] node61134;
	wire [4-1:0] node61136;
	wire [4-1:0] node61139;
	wire [4-1:0] node61142;
	wire [4-1:0] node61143;
	wire [4-1:0] node61146;
	wire [4-1:0] node61147;
	wire [4-1:0] node61151;
	wire [4-1:0] node61152;
	wire [4-1:0] node61153;
	wire [4-1:0] node61154;
	wire [4-1:0] node61155;
	wire [4-1:0] node61159;
	wire [4-1:0] node61160;
	wire [4-1:0] node61163;
	wire [4-1:0] node61166;
	wire [4-1:0] node61167;
	wire [4-1:0] node61169;
	wire [4-1:0] node61172;
	wire [4-1:0] node61173;
	wire [4-1:0] node61176;
	wire [4-1:0] node61179;
	wire [4-1:0] node61180;
	wire [4-1:0] node61181;
	wire [4-1:0] node61182;
	wire [4-1:0] node61185;
	wire [4-1:0] node61188;
	wire [4-1:0] node61190;
	wire [4-1:0] node61193;
	wire [4-1:0] node61194;
	wire [4-1:0] node61196;
	wire [4-1:0] node61200;
	wire [4-1:0] node61201;
	wire [4-1:0] node61202;
	wire [4-1:0] node61203;
	wire [4-1:0] node61204;
	wire [4-1:0] node61207;
	wire [4-1:0] node61210;
	wire [4-1:0] node61211;
	wire [4-1:0] node61213;
	wire [4-1:0] node61216;
	wire [4-1:0] node61217;
	wire [4-1:0] node61220;
	wire [4-1:0] node61223;
	wire [4-1:0] node61224;
	wire [4-1:0] node61225;
	wire [4-1:0] node61227;
	wire [4-1:0] node61230;
	wire [4-1:0] node61231;
	wire [4-1:0] node61234;
	wire [4-1:0] node61237;
	wire [4-1:0] node61239;
	wire [4-1:0] node61242;
	wire [4-1:0] node61243;
	wire [4-1:0] node61244;
	wire [4-1:0] node61245;
	wire [4-1:0] node61246;
	wire [4-1:0] node61249;
	wire [4-1:0] node61252;
	wire [4-1:0] node61253;
	wire [4-1:0] node61256;
	wire [4-1:0] node61259;
	wire [4-1:0] node61260;
	wire [4-1:0] node61261;
	wire [4-1:0] node61265;
	wire [4-1:0] node61266;
	wire [4-1:0] node61269;
	wire [4-1:0] node61272;
	wire [4-1:0] node61273;
	wire [4-1:0] node61274;
	wire [4-1:0] node61276;
	wire [4-1:0] node61279;
	wire [4-1:0] node61280;
	wire [4-1:0] node61283;
	wire [4-1:0] node61286;
	wire [4-1:0] node61288;
	wire [4-1:0] node61290;
	wire [4-1:0] node61293;
	wire [4-1:0] node61294;
	wire [4-1:0] node61295;
	wire [4-1:0] node61296;
	wire [4-1:0] node61297;
	wire [4-1:0] node61298;
	wire [4-1:0] node61300;
	wire [4-1:0] node61303;
	wire [4-1:0] node61304;
	wire [4-1:0] node61308;
	wire [4-1:0] node61311;
	wire [4-1:0] node61312;
	wire [4-1:0] node61313;
	wire [4-1:0] node61314;
	wire [4-1:0] node61317;
	wire [4-1:0] node61320;
	wire [4-1:0] node61321;
	wire [4-1:0] node61324;
	wire [4-1:0] node61327;
	wire [4-1:0] node61330;
	wire [4-1:0] node61331;
	wire [4-1:0] node61332;
	wire [4-1:0] node61334;
	wire [4-1:0] node61335;
	wire [4-1:0] node61338;
	wire [4-1:0] node61341;
	wire [4-1:0] node61343;
	wire [4-1:0] node61346;
	wire [4-1:0] node61347;
	wire [4-1:0] node61348;
	wire [4-1:0] node61350;
	wire [4-1:0] node61353;
	wire [4-1:0] node61354;
	wire [4-1:0] node61358;
	wire [4-1:0] node61359;
	wire [4-1:0] node61362;
	wire [4-1:0] node61365;
	wire [4-1:0] node61366;
	wire [4-1:0] node61367;
	wire [4-1:0] node61368;
	wire [4-1:0] node61369;
	wire [4-1:0] node61370;
	wire [4-1:0] node61374;
	wire [4-1:0] node61375;
	wire [4-1:0] node61378;
	wire [4-1:0] node61382;
	wire [4-1:0] node61383;
	wire [4-1:0] node61384;
	wire [4-1:0] node61386;
	wire [4-1:0] node61389;
	wire [4-1:0] node61392;
	wire [4-1:0] node61393;
	wire [4-1:0] node61396;
	wire [4-1:0] node61399;
	wire [4-1:0] node61400;
	wire [4-1:0] node61401;
	wire [4-1:0] node61402;
	wire [4-1:0] node61405;
	wire [4-1:0] node61407;
	wire [4-1:0] node61410;
	wire [4-1:0] node61411;
	wire [4-1:0] node61412;
	wire [4-1:0] node61416;
	wire [4-1:0] node61419;
	wire [4-1:0] node61420;
	wire [4-1:0] node61421;
	wire [4-1:0] node61423;
	wire [4-1:0] node61426;
	wire [4-1:0] node61427;
	wire [4-1:0] node61430;
	wire [4-1:0] node61433;
	wire [4-1:0] node61434;
	wire [4-1:0] node61438;
	wire [4-1:0] node61439;
	wire [4-1:0] node61440;
	wire [4-1:0] node61441;
	wire [4-1:0] node61442;
	wire [4-1:0] node61444;
	wire [4-1:0] node61445;
	wire [4-1:0] node61446;
	wire [4-1:0] node61451;
	wire [4-1:0] node61452;
	wire [4-1:0] node61453;
	wire [4-1:0] node61456;
	wire [4-1:0] node61457;
	wire [4-1:0] node61461;
	wire [4-1:0] node61462;
	wire [4-1:0] node61463;
	wire [4-1:0] node61467;
	wire [4-1:0] node61468;
	wire [4-1:0] node61472;
	wire [4-1:0] node61473;
	wire [4-1:0] node61474;
	wire [4-1:0] node61477;
	wire [4-1:0] node61478;
	wire [4-1:0] node61479;
	wire [4-1:0] node61484;
	wire [4-1:0] node61485;
	wire [4-1:0] node61486;
	wire [4-1:0] node61490;
	wire [4-1:0] node61491;
	wire [4-1:0] node61495;
	wire [4-1:0] node61496;
	wire [4-1:0] node61497;
	wire [4-1:0] node61498;
	wire [4-1:0] node61501;
	wire [4-1:0] node61502;
	wire [4-1:0] node61503;
	wire [4-1:0] node61507;
	wire [4-1:0] node61508;
	wire [4-1:0] node61512;
	wire [4-1:0] node61513;
	wire [4-1:0] node61514;
	wire [4-1:0] node61515;
	wire [4-1:0] node61519;
	wire [4-1:0] node61522;
	wire [4-1:0] node61523;
	wire [4-1:0] node61525;
	wire [4-1:0] node61528;
	wire [4-1:0] node61531;
	wire [4-1:0] node61532;
	wire [4-1:0] node61533;
	wire [4-1:0] node61534;
	wire [4-1:0] node61535;
	wire [4-1:0] node61540;
	wire [4-1:0] node61542;
	wire [4-1:0] node61543;
	wire [4-1:0] node61547;
	wire [4-1:0] node61548;
	wire [4-1:0] node61550;
	wire [4-1:0] node61553;
	wire [4-1:0] node61554;
	wire [4-1:0] node61555;
	wire [4-1:0] node61559;
	wire [4-1:0] node61562;
	wire [4-1:0] node61563;
	wire [4-1:0] node61564;
	wire [4-1:0] node61565;
	wire [4-1:0] node61566;
	wire [4-1:0] node61567;
	wire [4-1:0] node61568;
	wire [4-1:0] node61572;
	wire [4-1:0] node61575;
	wire [4-1:0] node61576;
	wire [4-1:0] node61580;
	wire [4-1:0] node61581;
	wire [4-1:0] node61582;
	wire [4-1:0] node61586;
	wire [4-1:0] node61587;
	wire [4-1:0] node61590;
	wire [4-1:0] node61593;
	wire [4-1:0] node61594;
	wire [4-1:0] node61595;
	wire [4-1:0] node61596;
	wire [4-1:0] node61597;
	wire [4-1:0] node61601;
	wire [4-1:0] node61604;
	wire [4-1:0] node61605;
	wire [4-1:0] node61606;
	wire [4-1:0] node61610;
	wire [4-1:0] node61611;
	wire [4-1:0] node61615;
	wire [4-1:0] node61616;
	wire [4-1:0] node61618;
	wire [4-1:0] node61621;
	wire [4-1:0] node61622;
	wire [4-1:0] node61623;
	wire [4-1:0] node61627;
	wire [4-1:0] node61628;
	wire [4-1:0] node61632;
	wire [4-1:0] node61633;
	wire [4-1:0] node61634;
	wire [4-1:0] node61635;
	wire [4-1:0] node61636;
	wire [4-1:0] node61637;
	wire [4-1:0] node61640;
	wire [4-1:0] node61644;
	wire [4-1:0] node61645;
	wire [4-1:0] node61648;
	wire [4-1:0] node61651;
	wire [4-1:0] node61652;
	wire [4-1:0] node61653;
	wire [4-1:0] node61654;
	wire [4-1:0] node61658;
	wire [4-1:0] node61659;
	wire [4-1:0] node61663;
	wire [4-1:0] node61664;
	wire [4-1:0] node61665;
	wire [4-1:0] node61670;
	wire [4-1:0] node61671;
	wire [4-1:0] node61672;
	wire [4-1:0] node61673;
	wire [4-1:0] node61676;
	wire [4-1:0] node61679;
	wire [4-1:0] node61680;
	wire [4-1:0] node61681;
	wire [4-1:0] node61686;
	wire [4-1:0] node61687;
	wire [4-1:0] node61689;
	wire [4-1:0] node61692;
	wire [4-1:0] node61693;
	wire [4-1:0] node61694;
	wire [4-1:0] node61698;
	wire [4-1:0] node61699;
	wire [4-1:0] node61703;
	wire [4-1:0] node61704;
	wire [4-1:0] node61705;
	wire [4-1:0] node61706;
	wire [4-1:0] node61707;
	wire [4-1:0] node61708;
	wire [4-1:0] node61709;
	wire [4-1:0] node61710;
	wire [4-1:0] node61713;
	wire [4-1:0] node61716;
	wire [4-1:0] node61717;
	wire [4-1:0] node61721;
	wire [4-1:0] node61722;
	wire [4-1:0] node61723;
	wire [4-1:0] node61726;
	wire [4-1:0] node61729;
	wire [4-1:0] node61730;
	wire [4-1:0] node61734;
	wire [4-1:0] node61735;
	wire [4-1:0] node61736;
	wire [4-1:0] node61737;
	wire [4-1:0] node61740;
	wire [4-1:0] node61743;
	wire [4-1:0] node61745;
	wire [4-1:0] node61747;
	wire [4-1:0] node61750;
	wire [4-1:0] node61751;
	wire [4-1:0] node61752;
	wire [4-1:0] node61755;
	wire [4-1:0] node61758;
	wire [4-1:0] node61759;
	wire [4-1:0] node61760;
	wire [4-1:0] node61763;
	wire [4-1:0] node61766;
	wire [4-1:0] node61767;
	wire [4-1:0] node61770;
	wire [4-1:0] node61773;
	wire [4-1:0] node61774;
	wire [4-1:0] node61775;
	wire [4-1:0] node61776;
	wire [4-1:0] node61777;
	wire [4-1:0] node61780;
	wire [4-1:0] node61783;
	wire [4-1:0] node61784;
	wire [4-1:0] node61785;
	wire [4-1:0] node61788;
	wire [4-1:0] node61792;
	wire [4-1:0] node61793;
	wire [4-1:0] node61794;
	wire [4-1:0] node61797;
	wire [4-1:0] node61800;
	wire [4-1:0] node61801;
	wire [4-1:0] node61804;
	wire [4-1:0] node61807;
	wire [4-1:0] node61808;
	wire [4-1:0] node61809;
	wire [4-1:0] node61810;
	wire [4-1:0] node61814;
	wire [4-1:0] node61815;
	wire [4-1:0] node61818;
	wire [4-1:0] node61821;
	wire [4-1:0] node61822;
	wire [4-1:0] node61823;
	wire [4-1:0] node61824;
	wire [4-1:0] node61827;
	wire [4-1:0] node61831;
	wire [4-1:0] node61832;
	wire [4-1:0] node61833;
	wire [4-1:0] node61836;
	wire [4-1:0] node61840;
	wire [4-1:0] node61841;
	wire [4-1:0] node61842;
	wire [4-1:0] node61843;
	wire [4-1:0] node61844;
	wire [4-1:0] node61845;
	wire [4-1:0] node61847;
	wire [4-1:0] node61850;
	wire [4-1:0] node61851;
	wire [4-1:0] node61854;
	wire [4-1:0] node61857;
	wire [4-1:0] node61858;
	wire [4-1:0] node61862;
	wire [4-1:0] node61863;
	wire [4-1:0] node61864;
	wire [4-1:0] node61867;
	wire [4-1:0] node61870;
	wire [4-1:0] node61871;
	wire [4-1:0] node61874;
	wire [4-1:0] node61877;
	wire [4-1:0] node61878;
	wire [4-1:0] node61879;
	wire [4-1:0] node61881;
	wire [4-1:0] node61882;
	wire [4-1:0] node61885;
	wire [4-1:0] node61888;
	wire [4-1:0] node61889;
	wire [4-1:0] node61892;
	wire [4-1:0] node61895;
	wire [4-1:0] node61896;
	wire [4-1:0] node61897;
	wire [4-1:0] node61901;
	wire [4-1:0] node61902;
	wire [4-1:0] node61905;
	wire [4-1:0] node61908;
	wire [4-1:0] node61909;
	wire [4-1:0] node61910;
	wire [4-1:0] node61911;
	wire [4-1:0] node61912;
	wire [4-1:0] node61915;
	wire [4-1:0] node61918;
	wire [4-1:0] node61919;
	wire [4-1:0] node61922;
	wire [4-1:0] node61925;
	wire [4-1:0] node61926;
	wire [4-1:0] node61927;
	wire [4-1:0] node61931;
	wire [4-1:0] node61934;
	wire [4-1:0] node61935;
	wire [4-1:0] node61936;
	wire [4-1:0] node61937;
	wire [4-1:0] node61940;
	wire [4-1:0] node61943;
	wire [4-1:0] node61945;
	wire [4-1:0] node61948;
	wire [4-1:0] node61949;
	wire [4-1:0] node61950;
	wire [4-1:0] node61953;
	wire [4-1:0] node61956;
	wire [4-1:0] node61957;
	wire [4-1:0] node61958;
	wire [4-1:0] node61961;
	wire [4-1:0] node61965;
	wire [4-1:0] node61966;
	wire [4-1:0] node61967;
	wire [4-1:0] node61968;
	wire [4-1:0] node61969;
	wire [4-1:0] node61970;
	wire [4-1:0] node61973;
	wire [4-1:0] node61976;
	wire [4-1:0] node61977;
	wire [4-1:0] node61980;
	wire [4-1:0] node61983;
	wire [4-1:0] node61984;
	wire [4-1:0] node61985;
	wire [4-1:0] node61989;
	wire [4-1:0] node61992;
	wire [4-1:0] node61993;
	wire [4-1:0] node61994;
	wire [4-1:0] node61995;
	wire [4-1:0] node61996;
	wire [4-1:0] node61997;
	wire [4-1:0] node62001;
	wire [4-1:0] node62002;
	wire [4-1:0] node62005;
	wire [4-1:0] node62008;
	wire [4-1:0] node62010;
	wire [4-1:0] node62013;
	wire [4-1:0] node62014;
	wire [4-1:0] node62017;
	wire [4-1:0] node62020;
	wire [4-1:0] node62021;
	wire [4-1:0] node62022;
	wire [4-1:0] node62026;
	wire [4-1:0] node62029;
	wire [4-1:0] node62030;
	wire [4-1:0] node62031;
	wire [4-1:0] node62032;
	wire [4-1:0] node62033;
	wire [4-1:0] node62034;
	wire [4-1:0] node62037;
	wire [4-1:0] node62040;
	wire [4-1:0] node62041;
	wire [4-1:0] node62044;
	wire [4-1:0] node62047;
	wire [4-1:0] node62048;
	wire [4-1:0] node62051;
	wire [4-1:0] node62054;
	wire [4-1:0] node62055;
	wire [4-1:0] node62056;
	wire [4-1:0] node62060;
	wire [4-1:0] node62063;
	wire [4-1:0] node62064;
	wire [4-1:0] node62065;
	wire [4-1:0] node62066;
	wire [4-1:0] node62068;
	wire [4-1:0] node62070;
	wire [4-1:0] node62073;
	wire [4-1:0] node62074;
	wire [4-1:0] node62075;
	wire [4-1:0] node62079;
	wire [4-1:0] node62080;
	wire [4-1:0] node62084;
	wire [4-1:0] node62085;
	wire [4-1:0] node62088;
	wire [4-1:0] node62091;
	wire [4-1:0] node62092;
	wire [4-1:0] node62093;
	wire [4-1:0] node62094;
	wire [4-1:0] node62098;
	wire [4-1:0] node62101;
	wire [4-1:0] node62102;
	wire [4-1:0] node62103;
	wire [4-1:0] node62105;
	wire [4-1:0] node62109;
	wire [4-1:0] node62110;
	wire [4-1:0] node62113;
	wire [4-1:0] node62116;
	wire [4-1:0] node62117;
	wire [4-1:0] node62118;
	wire [4-1:0] node62119;
	wire [4-1:0] node62120;
	wire [4-1:0] node62121;
	wire [4-1:0] node62122;
	wire [4-1:0] node62123;
	wire [4-1:0] node62124;
	wire [4-1:0] node62125;
	wire [4-1:0] node62126;
	wire [4-1:0] node62127;
	wire [4-1:0] node62132;
	wire [4-1:0] node62134;
	wire [4-1:0] node62136;
	wire [4-1:0] node62139;
	wire [4-1:0] node62140;
	wire [4-1:0] node62141;
	wire [4-1:0] node62144;
	wire [4-1:0] node62147;
	wire [4-1:0] node62148;
	wire [4-1:0] node62149;
	wire [4-1:0] node62152;
	wire [4-1:0] node62155;
	wire [4-1:0] node62156;
	wire [4-1:0] node62159;
	wire [4-1:0] node62162;
	wire [4-1:0] node62163;
	wire [4-1:0] node62164;
	wire [4-1:0] node62165;
	wire [4-1:0] node62166;
	wire [4-1:0] node62169;
	wire [4-1:0] node62172;
	wire [4-1:0] node62174;
	wire [4-1:0] node62177;
	wire [4-1:0] node62179;
	wire [4-1:0] node62181;
	wire [4-1:0] node62184;
	wire [4-1:0] node62185;
	wire [4-1:0] node62186;
	wire [4-1:0] node62190;
	wire [4-1:0] node62191;
	wire [4-1:0] node62192;
	wire [4-1:0] node62195;
	wire [4-1:0] node62198;
	wire [4-1:0] node62199;
	wire [4-1:0] node62203;
	wire [4-1:0] node62204;
	wire [4-1:0] node62205;
	wire [4-1:0] node62206;
	wire [4-1:0] node62208;
	wire [4-1:0] node62209;
	wire [4-1:0] node62212;
	wire [4-1:0] node62215;
	wire [4-1:0] node62216;
	wire [4-1:0] node62217;
	wire [4-1:0] node62221;
	wire [4-1:0] node62222;
	wire [4-1:0] node62225;
	wire [4-1:0] node62228;
	wire [4-1:0] node62229;
	wire [4-1:0] node62230;
	wire [4-1:0] node62231;
	wire [4-1:0] node62235;
	wire [4-1:0] node62237;
	wire [4-1:0] node62240;
	wire [4-1:0] node62242;
	wire [4-1:0] node62245;
	wire [4-1:0] node62246;
	wire [4-1:0] node62247;
	wire [4-1:0] node62248;
	wire [4-1:0] node62249;
	wire [4-1:0] node62252;
	wire [4-1:0] node62256;
	wire [4-1:0] node62257;
	wire [4-1:0] node62261;
	wire [4-1:0] node62262;
	wire [4-1:0] node62263;
	wire [4-1:0] node62264;
	wire [4-1:0] node62268;
	wire [4-1:0] node62269;
	wire [4-1:0] node62273;
	wire [4-1:0] node62275;
	wire [4-1:0] node62276;
	wire [4-1:0] node62279;
	wire [4-1:0] node62282;
	wire [4-1:0] node62283;
	wire [4-1:0] node62284;
	wire [4-1:0] node62285;
	wire [4-1:0] node62286;
	wire [4-1:0] node62287;
	wire [4-1:0] node62288;
	wire [4-1:0] node62291;
	wire [4-1:0] node62295;
	wire [4-1:0] node62296;
	wire [4-1:0] node62300;
	wire [4-1:0] node62301;
	wire [4-1:0] node62302;
	wire [4-1:0] node62303;
	wire [4-1:0] node62306;
	wire [4-1:0] node62309;
	wire [4-1:0] node62310;
	wire [4-1:0] node62313;
	wire [4-1:0] node62316;
	wire [4-1:0] node62317;
	wire [4-1:0] node62318;
	wire [4-1:0] node62321;
	wire [4-1:0] node62325;
	wire [4-1:0] node62326;
	wire [4-1:0] node62327;
	wire [4-1:0] node62328;
	wire [4-1:0] node62329;
	wire [4-1:0] node62333;
	wire [4-1:0] node62334;
	wire [4-1:0] node62337;
	wire [4-1:0] node62340;
	wire [4-1:0] node62341;
	wire [4-1:0] node62343;
	wire [4-1:0] node62347;
	wire [4-1:0] node62348;
	wire [4-1:0] node62349;
	wire [4-1:0] node62353;
	wire [4-1:0] node62354;
	wire [4-1:0] node62357;
	wire [4-1:0] node62360;
	wire [4-1:0] node62361;
	wire [4-1:0] node62362;
	wire [4-1:0] node62363;
	wire [4-1:0] node62364;
	wire [4-1:0] node62365;
	wire [4-1:0] node62368;
	wire [4-1:0] node62372;
	wire [4-1:0] node62373;
	wire [4-1:0] node62374;
	wire [4-1:0] node62379;
	wire [4-1:0] node62380;
	wire [4-1:0] node62381;
	wire [4-1:0] node62384;
	wire [4-1:0] node62387;
	wire [4-1:0] node62388;
	wire [4-1:0] node62392;
	wire [4-1:0] node62393;
	wire [4-1:0] node62394;
	wire [4-1:0] node62396;
	wire [4-1:0] node62398;
	wire [4-1:0] node62401;
	wire [4-1:0] node62402;
	wire [4-1:0] node62406;
	wire [4-1:0] node62407;
	wire [4-1:0] node62408;
	wire [4-1:0] node62411;
	wire [4-1:0] node62414;
	wire [4-1:0] node62415;
	wire [4-1:0] node62418;
	wire [4-1:0] node62421;
	wire [4-1:0] node62422;
	wire [4-1:0] node62423;
	wire [4-1:0] node62424;
	wire [4-1:0] node62425;
	wire [4-1:0] node62426;
	wire [4-1:0] node62427;
	wire [4-1:0] node62428;
	wire [4-1:0] node62431;
	wire [4-1:0] node62434;
	wire [4-1:0] node62436;
	wire [4-1:0] node62439;
	wire [4-1:0] node62440;
	wire [4-1:0] node62441;
	wire [4-1:0] node62444;
	wire [4-1:0] node62447;
	wire [4-1:0] node62449;
	wire [4-1:0] node62452;
	wire [4-1:0] node62453;
	wire [4-1:0] node62454;
	wire [4-1:0] node62455;
	wire [4-1:0] node62458;
	wire [4-1:0] node62461;
	wire [4-1:0] node62462;
	wire [4-1:0] node62465;
	wire [4-1:0] node62468;
	wire [4-1:0] node62469;
	wire [4-1:0] node62470;
	wire [4-1:0] node62473;
	wire [4-1:0] node62476;
	wire [4-1:0] node62477;
	wire [4-1:0] node62481;
	wire [4-1:0] node62482;
	wire [4-1:0] node62483;
	wire [4-1:0] node62484;
	wire [4-1:0] node62485;
	wire [4-1:0] node62489;
	wire [4-1:0] node62490;
	wire [4-1:0] node62493;
	wire [4-1:0] node62496;
	wire [4-1:0] node62497;
	wire [4-1:0] node62498;
	wire [4-1:0] node62502;
	wire [4-1:0] node62503;
	wire [4-1:0] node62507;
	wire [4-1:0] node62508;
	wire [4-1:0] node62509;
	wire [4-1:0] node62510;
	wire [4-1:0] node62513;
	wire [4-1:0] node62517;
	wire [4-1:0] node62518;
	wire [4-1:0] node62520;
	wire [4-1:0] node62523;
	wire [4-1:0] node62525;
	wire [4-1:0] node62528;
	wire [4-1:0] node62529;
	wire [4-1:0] node62530;
	wire [4-1:0] node62531;
	wire [4-1:0] node62532;
	wire [4-1:0] node62534;
	wire [4-1:0] node62537;
	wire [4-1:0] node62538;
	wire [4-1:0] node62541;
	wire [4-1:0] node62544;
	wire [4-1:0] node62545;
	wire [4-1:0] node62546;
	wire [4-1:0] node62549;
	wire [4-1:0] node62552;
	wire [4-1:0] node62553;
	wire [4-1:0] node62557;
	wire [4-1:0] node62558;
	wire [4-1:0] node62559;
	wire [4-1:0] node62560;
	wire [4-1:0] node62563;
	wire [4-1:0] node62567;
	wire [4-1:0] node62568;
	wire [4-1:0] node62571;
	wire [4-1:0] node62574;
	wire [4-1:0] node62575;
	wire [4-1:0] node62576;
	wire [4-1:0] node62577;
	wire [4-1:0] node62578;
	wire [4-1:0] node62583;
	wire [4-1:0] node62584;
	wire [4-1:0] node62585;
	wire [4-1:0] node62588;
	wire [4-1:0] node62591;
	wire [4-1:0] node62592;
	wire [4-1:0] node62596;
	wire [4-1:0] node62597;
	wire [4-1:0] node62598;
	wire [4-1:0] node62601;
	wire [4-1:0] node62604;
	wire [4-1:0] node62605;
	wire [4-1:0] node62608;
	wire [4-1:0] node62611;
	wire [4-1:0] node62612;
	wire [4-1:0] node62613;
	wire [4-1:0] node62614;
	wire [4-1:0] node62615;
	wire [4-1:0] node62616;
	wire [4-1:0] node62617;
	wire [4-1:0] node62620;
	wire [4-1:0] node62624;
	wire [4-1:0] node62625;
	wire [4-1:0] node62626;
	wire [4-1:0] node62630;
	wire [4-1:0] node62631;
	wire [4-1:0] node62635;
	wire [4-1:0] node62636;
	wire [4-1:0] node62637;
	wire [4-1:0] node62638;
	wire [4-1:0] node62641;
	wire [4-1:0] node62644;
	wire [4-1:0] node62645;
	wire [4-1:0] node62648;
	wire [4-1:0] node62651;
	wire [4-1:0] node62653;
	wire [4-1:0] node62656;
	wire [4-1:0] node62657;
	wire [4-1:0] node62658;
	wire [4-1:0] node62659;
	wire [4-1:0] node62660;
	wire [4-1:0] node62664;
	wire [4-1:0] node62665;
	wire [4-1:0] node62668;
	wire [4-1:0] node62671;
	wire [4-1:0] node62672;
	wire [4-1:0] node62675;
	wire [4-1:0] node62678;
	wire [4-1:0] node62679;
	wire [4-1:0] node62680;
	wire [4-1:0] node62681;
	wire [4-1:0] node62685;
	wire [4-1:0] node62687;
	wire [4-1:0] node62690;
	wire [4-1:0] node62692;
	wire [4-1:0] node62695;
	wire [4-1:0] node62696;
	wire [4-1:0] node62697;
	wire [4-1:0] node62698;
	wire [4-1:0] node62700;
	wire [4-1:0] node62701;
	wire [4-1:0] node62705;
	wire [4-1:0] node62706;
	wire [4-1:0] node62709;
	wire [4-1:0] node62712;
	wire [4-1:0] node62713;
	wire [4-1:0] node62714;
	wire [4-1:0] node62715;
	wire [4-1:0] node62719;
	wire [4-1:0] node62720;
	wire [4-1:0] node62723;
	wire [4-1:0] node62726;
	wire [4-1:0] node62727;
	wire [4-1:0] node62728;
	wire [4-1:0] node62731;
	wire [4-1:0] node62734;
	wire [4-1:0] node62736;
	wire [4-1:0] node62739;
	wire [4-1:0] node62740;
	wire [4-1:0] node62741;
	wire [4-1:0] node62743;
	wire [4-1:0] node62744;
	wire [4-1:0] node62747;
	wire [4-1:0] node62750;
	wire [4-1:0] node62751;
	wire [4-1:0] node62754;
	wire [4-1:0] node62757;
	wire [4-1:0] node62758;
	wire [4-1:0] node62761;
	wire [4-1:0] node62762;
	wire [4-1:0] node62763;
	wire [4-1:0] node62767;
	wire [4-1:0] node62769;
	wire [4-1:0] node62772;
	wire [4-1:0] node62773;
	wire [4-1:0] node62774;
	wire [4-1:0] node62775;
	wire [4-1:0] node62776;
	wire [4-1:0] node62777;
	wire [4-1:0] node62778;
	wire [4-1:0] node62780;
	wire [4-1:0] node62781;
	wire [4-1:0] node62784;
	wire [4-1:0] node62787;
	wire [4-1:0] node62788;
	wire [4-1:0] node62790;
	wire [4-1:0] node62793;
	wire [4-1:0] node62794;
	wire [4-1:0] node62798;
	wire [4-1:0] node62799;
	wire [4-1:0] node62800;
	wire [4-1:0] node62801;
	wire [4-1:0] node62804;
	wire [4-1:0] node62807;
	wire [4-1:0] node62808;
	wire [4-1:0] node62811;
	wire [4-1:0] node62814;
	wire [4-1:0] node62815;
	wire [4-1:0] node62816;
	wire [4-1:0] node62820;
	wire [4-1:0] node62821;
	wire [4-1:0] node62824;
	wire [4-1:0] node62827;
	wire [4-1:0] node62828;
	wire [4-1:0] node62829;
	wire [4-1:0] node62830;
	wire [4-1:0] node62832;
	wire [4-1:0] node62836;
	wire [4-1:0] node62837;
	wire [4-1:0] node62839;
	wire [4-1:0] node62842;
	wire [4-1:0] node62845;
	wire [4-1:0] node62846;
	wire [4-1:0] node62847;
	wire [4-1:0] node62848;
	wire [4-1:0] node62852;
	wire [4-1:0] node62854;
	wire [4-1:0] node62857;
	wire [4-1:0] node62858;
	wire [4-1:0] node62859;
	wire [4-1:0] node62862;
	wire [4-1:0] node62865;
	wire [4-1:0] node62866;
	wire [4-1:0] node62869;
	wire [4-1:0] node62872;
	wire [4-1:0] node62873;
	wire [4-1:0] node62874;
	wire [4-1:0] node62875;
	wire [4-1:0] node62876;
	wire [4-1:0] node62879;
	wire [4-1:0] node62882;
	wire [4-1:0] node62883;
	wire [4-1:0] node62886;
	wire [4-1:0] node62889;
	wire [4-1:0] node62890;
	wire [4-1:0] node62891;
	wire [4-1:0] node62892;
	wire [4-1:0] node62895;
	wire [4-1:0] node62898;
	wire [4-1:0] node62900;
	wire [4-1:0] node62903;
	wire [4-1:0] node62904;
	wire [4-1:0] node62905;
	wire [4-1:0] node62908;
	wire [4-1:0] node62911;
	wire [4-1:0] node62912;
	wire [4-1:0] node62915;
	wire [4-1:0] node62918;
	wire [4-1:0] node62919;
	wire [4-1:0] node62920;
	wire [4-1:0] node62921;
	wire [4-1:0] node62924;
	wire [4-1:0] node62927;
	wire [4-1:0] node62928;
	wire [4-1:0] node62929;
	wire [4-1:0] node62932;
	wire [4-1:0] node62936;
	wire [4-1:0] node62938;
	wire [4-1:0] node62939;
	wire [4-1:0] node62941;
	wire [4-1:0] node62944;
	wire [4-1:0] node62945;
	wire [4-1:0] node62949;
	wire [4-1:0] node62950;
	wire [4-1:0] node62951;
	wire [4-1:0] node62952;
	wire [4-1:0] node62953;
	wire [4-1:0] node62954;
	wire [4-1:0] node62956;
	wire [4-1:0] node62959;
	wire [4-1:0] node62960;
	wire [4-1:0] node62964;
	wire [4-1:0] node62965;
	wire [4-1:0] node62967;
	wire [4-1:0] node62970;
	wire [4-1:0] node62971;
	wire [4-1:0] node62975;
	wire [4-1:0] node62976;
	wire [4-1:0] node62977;
	wire [4-1:0] node62980;
	wire [4-1:0] node62983;
	wire [4-1:0] node62984;
	wire [4-1:0] node62987;
	wire [4-1:0] node62990;
	wire [4-1:0] node62991;
	wire [4-1:0] node62992;
	wire [4-1:0] node62993;
	wire [4-1:0] node62994;
	wire [4-1:0] node62998;
	wire [4-1:0] node62999;
	wire [4-1:0] node63003;
	wire [4-1:0] node63006;
	wire [4-1:0] node63007;
	wire [4-1:0] node63008;
	wire [4-1:0] node63011;
	wire [4-1:0] node63014;
	wire [4-1:0] node63016;
	wire [4-1:0] node63019;
	wire [4-1:0] node63020;
	wire [4-1:0] node63021;
	wire [4-1:0] node63022;
	wire [4-1:0] node63023;
	wire [4-1:0] node63025;
	wire [4-1:0] node63028;
	wire [4-1:0] node63029;
	wire [4-1:0] node63032;
	wire [4-1:0] node63035;
	wire [4-1:0] node63037;
	wire [4-1:0] node63040;
	wire [4-1:0] node63041;
	wire [4-1:0] node63042;
	wire [4-1:0] node63043;
	wire [4-1:0] node63047;
	wire [4-1:0] node63048;
	wire [4-1:0] node63051;
	wire [4-1:0] node63054;
	wire [4-1:0] node63055;
	wire [4-1:0] node63059;
	wire [4-1:0] node63060;
	wire [4-1:0] node63061;
	wire [4-1:0] node63063;
	wire [4-1:0] node63064;
	wire [4-1:0] node63067;
	wire [4-1:0] node63070;
	wire [4-1:0] node63071;
	wire [4-1:0] node63073;
	wire [4-1:0] node63076;
	wire [4-1:0] node63077;
	wire [4-1:0] node63080;
	wire [4-1:0] node63083;
	wire [4-1:0] node63084;
	wire [4-1:0] node63085;
	wire [4-1:0] node63087;
	wire [4-1:0] node63090;
	wire [4-1:0] node63091;
	wire [4-1:0] node63094;
	wire [4-1:0] node63097;
	wire [4-1:0] node63098;
	wire [4-1:0] node63099;
	wire [4-1:0] node63102;
	wire [4-1:0] node63106;
	wire [4-1:0] node63107;
	wire [4-1:0] node63108;
	wire [4-1:0] node63109;
	wire [4-1:0] node63110;
	wire [4-1:0] node63111;
	wire [4-1:0] node63112;
	wire [4-1:0] node63114;
	wire [4-1:0] node63118;
	wire [4-1:0] node63119;
	wire [4-1:0] node63120;
	wire [4-1:0] node63123;
	wire [4-1:0] node63126;
	wire [4-1:0] node63127;
	wire [4-1:0] node63130;
	wire [4-1:0] node63133;
	wire [4-1:0] node63134;
	wire [4-1:0] node63135;
	wire [4-1:0] node63136;
	wire [4-1:0] node63139;
	wire [4-1:0] node63142;
	wire [4-1:0] node63143;
	wire [4-1:0] node63147;
	wire [4-1:0] node63149;
	wire [4-1:0] node63152;
	wire [4-1:0] node63153;
	wire [4-1:0] node63154;
	wire [4-1:0] node63156;
	wire [4-1:0] node63157;
	wire [4-1:0] node63160;
	wire [4-1:0] node63163;
	wire [4-1:0] node63165;
	wire [4-1:0] node63168;
	wire [4-1:0] node63169;
	wire [4-1:0] node63170;
	wire [4-1:0] node63173;
	wire [4-1:0] node63176;
	wire [4-1:0] node63178;
	wire [4-1:0] node63181;
	wire [4-1:0] node63182;
	wire [4-1:0] node63183;
	wire [4-1:0] node63184;
	wire [4-1:0] node63185;
	wire [4-1:0] node63186;
	wire [4-1:0] node63189;
	wire [4-1:0] node63193;
	wire [4-1:0] node63195;
	wire [4-1:0] node63196;
	wire [4-1:0] node63200;
	wire [4-1:0] node63201;
	wire [4-1:0] node63202;
	wire [4-1:0] node63203;
	wire [4-1:0] node63206;
	wire [4-1:0] node63209;
	wire [4-1:0] node63210;
	wire [4-1:0] node63213;
	wire [4-1:0] node63216;
	wire [4-1:0] node63217;
	wire [4-1:0] node63220;
	wire [4-1:0] node63223;
	wire [4-1:0] node63224;
	wire [4-1:0] node63225;
	wire [4-1:0] node63226;
	wire [4-1:0] node63227;
	wire [4-1:0] node63230;
	wire [4-1:0] node63233;
	wire [4-1:0] node63235;
	wire [4-1:0] node63238;
	wire [4-1:0] node63239;
	wire [4-1:0] node63240;
	wire [4-1:0] node63243;
	wire [4-1:0] node63247;
	wire [4-1:0] node63248;
	wire [4-1:0] node63249;
	wire [4-1:0] node63252;
	wire [4-1:0] node63255;
	wire [4-1:0] node63256;
	wire [4-1:0] node63258;
	wire [4-1:0] node63261;
	wire [4-1:0] node63264;
	wire [4-1:0] node63265;
	wire [4-1:0] node63266;
	wire [4-1:0] node63267;
	wire [4-1:0] node63268;
	wire [4-1:0] node63269;
	wire [4-1:0] node63270;
	wire [4-1:0] node63273;
	wire [4-1:0] node63277;
	wire [4-1:0] node63279;
	wire [4-1:0] node63280;
	wire [4-1:0] node63283;
	wire [4-1:0] node63286;
	wire [4-1:0] node63287;
	wire [4-1:0] node63289;
	wire [4-1:0] node63290;
	wire [4-1:0] node63293;
	wire [4-1:0] node63296;
	wire [4-1:0] node63297;
	wire [4-1:0] node63299;
	wire [4-1:0] node63303;
	wire [4-1:0] node63304;
	wire [4-1:0] node63305;
	wire [4-1:0] node63306;
	wire [4-1:0] node63307;
	wire [4-1:0] node63310;
	wire [4-1:0] node63314;
	wire [4-1:0] node63315;
	wire [4-1:0] node63317;
	wire [4-1:0] node63320;
	wire [4-1:0] node63321;
	wire [4-1:0] node63324;
	wire [4-1:0] node63327;
	wire [4-1:0] node63328;
	wire [4-1:0] node63329;
	wire [4-1:0] node63332;
	wire [4-1:0] node63335;
	wire [4-1:0] node63336;
	wire [4-1:0] node63337;
	wire [4-1:0] node63341;
	wire [4-1:0] node63342;
	wire [4-1:0] node63345;
	wire [4-1:0] node63348;
	wire [4-1:0] node63349;
	wire [4-1:0] node63350;
	wire [4-1:0] node63351;
	wire [4-1:0] node63352;
	wire [4-1:0] node63353;
	wire [4-1:0] node63356;
	wire [4-1:0] node63359;
	wire [4-1:0] node63360;
	wire [4-1:0] node63363;
	wire [4-1:0] node63366;
	wire [4-1:0] node63367;
	wire [4-1:0] node63368;
	wire [4-1:0] node63371;
	wire [4-1:0] node63375;
	wire [4-1:0] node63376;
	wire [4-1:0] node63377;
	wire [4-1:0] node63380;
	wire [4-1:0] node63383;
	wire [4-1:0] node63384;
	wire [4-1:0] node63385;
	wire [4-1:0] node63388;
	wire [4-1:0] node63392;
	wire [4-1:0] node63393;
	wire [4-1:0] node63394;
	wire [4-1:0] node63396;
	wire [4-1:0] node63398;
	wire [4-1:0] node63401;
	wire [4-1:0] node63402;
	wire [4-1:0] node63404;
	wire [4-1:0] node63408;
	wire [4-1:0] node63409;
	wire [4-1:0] node63410;
	wire [4-1:0] node63411;
	wire [4-1:0] node63414;
	wire [4-1:0] node63417;
	wire [4-1:0] node63418;
	wire [4-1:0] node63422;
	wire [4-1:0] node63423;
	wire [4-1:0] node63426;
	wire [4-1:0] node63429;
	wire [4-1:0] node63430;
	wire [4-1:0] node63431;
	wire [4-1:0] node63432;
	wire [4-1:0] node63433;
	wire [4-1:0] node63434;
	wire [4-1:0] node63435;
	wire [4-1:0] node63436;
	wire [4-1:0] node63439;
	wire [4-1:0] node63440;
	wire [4-1:0] node63442;
	wire [4-1:0] node63445;
	wire [4-1:0] node63446;
	wire [4-1:0] node63449;
	wire [4-1:0] node63452;
	wire [4-1:0] node63453;
	wire [4-1:0] node63454;
	wire [4-1:0] node63456;
	wire [4-1:0] node63460;
	wire [4-1:0] node63461;
	wire [4-1:0] node63462;
	wire [4-1:0] node63465;
	wire [4-1:0] node63469;
	wire [4-1:0] node63470;
	wire [4-1:0] node63471;
	wire [4-1:0] node63472;
	wire [4-1:0] node63474;
	wire [4-1:0] node63477;
	wire [4-1:0] node63478;
	wire [4-1:0] node63482;
	wire [4-1:0] node63483;
	wire [4-1:0] node63484;
	wire [4-1:0] node63487;
	wire [4-1:0] node63490;
	wire [4-1:0] node63492;
	wire [4-1:0] node63495;
	wire [4-1:0] node63496;
	wire [4-1:0] node63497;
	wire [4-1:0] node63498;
	wire [4-1:0] node63501;
	wire [4-1:0] node63504;
	wire [4-1:0] node63505;
	wire [4-1:0] node63508;
	wire [4-1:0] node63511;
	wire [4-1:0] node63512;
	wire [4-1:0] node63513;
	wire [4-1:0] node63517;
	wire [4-1:0] node63519;
	wire [4-1:0] node63522;
	wire [4-1:0] node63523;
	wire [4-1:0] node63524;
	wire [4-1:0] node63525;
	wire [4-1:0] node63526;
	wire [4-1:0] node63527;
	wire [4-1:0] node63530;
	wire [4-1:0] node63533;
	wire [4-1:0] node63536;
	wire [4-1:0] node63537;
	wire [4-1:0] node63540;
	wire [4-1:0] node63542;
	wire [4-1:0] node63545;
	wire [4-1:0] node63546;
	wire [4-1:0] node63549;
	wire [4-1:0] node63550;
	wire [4-1:0] node63551;
	wire [4-1:0] node63555;
	wire [4-1:0] node63556;
	wire [4-1:0] node63560;
	wire [4-1:0] node63561;
	wire [4-1:0] node63562;
	wire [4-1:0] node63563;
	wire [4-1:0] node63564;
	wire [4-1:0] node63567;
	wire [4-1:0] node63571;
	wire [4-1:0] node63572;
	wire [4-1:0] node63575;
	wire [4-1:0] node63578;
	wire [4-1:0] node63579;
	wire [4-1:0] node63580;
	wire [4-1:0] node63582;
	wire [4-1:0] node63586;
	wire [4-1:0] node63587;
	wire [4-1:0] node63591;
	wire [4-1:0] node63592;
	wire [4-1:0] node63593;
	wire [4-1:0] node63594;
	wire [4-1:0] node63595;
	wire [4-1:0] node63596;
	wire [4-1:0] node63597;
	wire [4-1:0] node63601;
	wire [4-1:0] node63602;
	wire [4-1:0] node63606;
	wire [4-1:0] node63607;
	wire [4-1:0] node63609;
	wire [4-1:0] node63612;
	wire [4-1:0] node63614;
	wire [4-1:0] node63617;
	wire [4-1:0] node63618;
	wire [4-1:0] node63619;
	wire [4-1:0] node63622;
	wire [4-1:0] node63625;
	wire [4-1:0] node63626;
	wire [4-1:0] node63628;
	wire [4-1:0] node63631;
	wire [4-1:0] node63632;
	wire [4-1:0] node63636;
	wire [4-1:0] node63637;
	wire [4-1:0] node63638;
	wire [4-1:0] node63639;
	wire [4-1:0] node63640;
	wire [4-1:0] node63643;
	wire [4-1:0] node63646;
	wire [4-1:0] node63647;
	wire [4-1:0] node63650;
	wire [4-1:0] node63653;
	wire [4-1:0] node63654;
	wire [4-1:0] node63656;
	wire [4-1:0] node63659;
	wire [4-1:0] node63660;
	wire [4-1:0] node63664;
	wire [4-1:0] node63665;
	wire [4-1:0] node63666;
	wire [4-1:0] node63667;
	wire [4-1:0] node63670;
	wire [4-1:0] node63674;
	wire [4-1:0] node63675;
	wire [4-1:0] node63678;
	wire [4-1:0] node63681;
	wire [4-1:0] node63682;
	wire [4-1:0] node63683;
	wire [4-1:0] node63684;
	wire [4-1:0] node63685;
	wire [4-1:0] node63686;
	wire [4-1:0] node63689;
	wire [4-1:0] node63692;
	wire [4-1:0] node63693;
	wire [4-1:0] node63696;
	wire [4-1:0] node63699;
	wire [4-1:0] node63700;
	wire [4-1:0] node63702;
	wire [4-1:0] node63705;
	wire [4-1:0] node63707;
	wire [4-1:0] node63710;
	wire [4-1:0] node63711;
	wire [4-1:0] node63712;
	wire [4-1:0] node63715;
	wire [4-1:0] node63718;
	wire [4-1:0] node63719;
	wire [4-1:0] node63723;
	wire [4-1:0] node63724;
	wire [4-1:0] node63725;
	wire [4-1:0] node63726;
	wire [4-1:0] node63727;
	wire [4-1:0] node63730;
	wire [4-1:0] node63733;
	wire [4-1:0] node63735;
	wire [4-1:0] node63738;
	wire [4-1:0] node63740;
	wire [4-1:0] node63741;
	wire [4-1:0] node63744;
	wire [4-1:0] node63747;
	wire [4-1:0] node63748;
	wire [4-1:0] node63749;
	wire [4-1:0] node63753;
	wire [4-1:0] node63754;
	wire [4-1:0] node63757;
	wire [4-1:0] node63760;
	wire [4-1:0] node63761;
	wire [4-1:0] node63762;
	wire [4-1:0] node63763;
	wire [4-1:0] node63764;
	wire [4-1:0] node63765;
	wire [4-1:0] node63766;
	wire [4-1:0] node63767;
	wire [4-1:0] node63770;
	wire [4-1:0] node63774;
	wire [4-1:0] node63775;
	wire [4-1:0] node63777;
	wire [4-1:0] node63780;
	wire [4-1:0] node63781;
	wire [4-1:0] node63784;
	wire [4-1:0] node63787;
	wire [4-1:0] node63788;
	wire [4-1:0] node63789;
	wire [4-1:0] node63792;
	wire [4-1:0] node63795;
	wire [4-1:0] node63796;
	wire [4-1:0] node63799;
	wire [4-1:0] node63802;
	wire [4-1:0] node63803;
	wire [4-1:0] node63804;
	wire [4-1:0] node63805;
	wire [4-1:0] node63806;
	wire [4-1:0] node63809;
	wire [4-1:0] node63812;
	wire [4-1:0] node63813;
	wire [4-1:0] node63816;
	wire [4-1:0] node63819;
	wire [4-1:0] node63820;
	wire [4-1:0] node63821;
	wire [4-1:0] node63825;
	wire [4-1:0] node63827;
	wire [4-1:0] node63830;
	wire [4-1:0] node63831;
	wire [4-1:0] node63832;
	wire [4-1:0] node63835;
	wire [4-1:0] node63838;
	wire [4-1:0] node63839;
	wire [4-1:0] node63842;
	wire [4-1:0] node63845;
	wire [4-1:0] node63846;
	wire [4-1:0] node63847;
	wire [4-1:0] node63848;
	wire [4-1:0] node63850;
	wire [4-1:0] node63852;
	wire [4-1:0] node63855;
	wire [4-1:0] node63857;
	wire [4-1:0] node63858;
	wire [4-1:0] node63861;
	wire [4-1:0] node63864;
	wire [4-1:0] node63865;
	wire [4-1:0] node63866;
	wire [4-1:0] node63869;
	wire [4-1:0] node63872;
	wire [4-1:0] node63873;
	wire [4-1:0] node63876;
	wire [4-1:0] node63879;
	wire [4-1:0] node63880;
	wire [4-1:0] node63881;
	wire [4-1:0] node63882;
	wire [4-1:0] node63883;
	wire [4-1:0] node63887;
	wire [4-1:0] node63888;
	wire [4-1:0] node63892;
	wire [4-1:0] node63894;
	wire [4-1:0] node63895;
	wire [4-1:0] node63899;
	wire [4-1:0] node63900;
	wire [4-1:0] node63901;
	wire [4-1:0] node63902;
	wire [4-1:0] node63905;
	wire [4-1:0] node63908;
	wire [4-1:0] node63909;
	wire [4-1:0] node63913;
	wire [4-1:0] node63915;
	wire [4-1:0] node63916;
	wire [4-1:0] node63919;
	wire [4-1:0] node63922;
	wire [4-1:0] node63923;
	wire [4-1:0] node63924;
	wire [4-1:0] node63925;
	wire [4-1:0] node63926;
	wire [4-1:0] node63927;
	wire [4-1:0] node63928;
	wire [4-1:0] node63931;
	wire [4-1:0] node63935;
	wire [4-1:0] node63936;
	wire [4-1:0] node63940;
	wire [4-1:0] node63941;
	wire [4-1:0] node63942;
	wire [4-1:0] node63944;
	wire [4-1:0] node63948;
	wire [4-1:0] node63949;
	wire [4-1:0] node63950;
	wire [4-1:0] node63954;
	wire [4-1:0] node63956;
	wire [4-1:0] node63959;
	wire [4-1:0] node63960;
	wire [4-1:0] node63961;
	wire [4-1:0] node63962;
	wire [4-1:0] node63963;
	wire [4-1:0] node63966;
	wire [4-1:0] node63969;
	wire [4-1:0] node63970;
	wire [4-1:0] node63973;
	wire [4-1:0] node63976;
	wire [4-1:0] node63977;
	wire [4-1:0] node63978;
	wire [4-1:0] node63981;
	wire [4-1:0] node63984;
	wire [4-1:0] node63986;
	wire [4-1:0] node63989;
	wire [4-1:0] node63990;
	wire [4-1:0] node63991;
	wire [4-1:0] node63992;
	wire [4-1:0] node63996;
	wire [4-1:0] node63997;
	wire [4-1:0] node64000;
	wire [4-1:0] node64003;
	wire [4-1:0] node64004;
	wire [4-1:0] node64005;
	wire [4-1:0] node64010;
	wire [4-1:0] node64011;
	wire [4-1:0] node64012;
	wire [4-1:0] node64013;
	wire [4-1:0] node64015;
	wire [4-1:0] node64017;
	wire [4-1:0] node64020;
	wire [4-1:0] node64021;
	wire [4-1:0] node64022;
	wire [4-1:0] node64025;
	wire [4-1:0] node64028;
	wire [4-1:0] node64029;
	wire [4-1:0] node64033;
	wire [4-1:0] node64034;
	wire [4-1:0] node64035;
	wire [4-1:0] node64036;
	wire [4-1:0] node64039;
	wire [4-1:0] node64042;
	wire [4-1:0] node64043;
	wire [4-1:0] node64046;
	wire [4-1:0] node64049;
	wire [4-1:0] node64050;
	wire [4-1:0] node64051;
	wire [4-1:0] node64055;
	wire [4-1:0] node64056;
	wire [4-1:0] node64059;
	wire [4-1:0] node64062;
	wire [4-1:0] node64063;
	wire [4-1:0] node64064;
	wire [4-1:0] node64065;
	wire [4-1:0] node64068;
	wire [4-1:0] node64069;
	wire [4-1:0] node64072;
	wire [4-1:0] node64075;
	wire [4-1:0] node64076;
	wire [4-1:0] node64078;
	wire [4-1:0] node64081;
	wire [4-1:0] node64084;
	wire [4-1:0] node64085;
	wire [4-1:0] node64086;
	wire [4-1:0] node64087;
	wire [4-1:0] node64090;
	wire [4-1:0] node64093;
	wire [4-1:0] node64094;
	wire [4-1:0] node64097;
	wire [4-1:0] node64100;
	wire [4-1:0] node64101;
	wire [4-1:0] node64103;
	wire [4-1:0] node64106;
	wire [4-1:0] node64107;
	wire [4-1:0] node64111;
	wire [4-1:0] node64112;
	wire [4-1:0] node64113;
	wire [4-1:0] node64114;
	wire [4-1:0] node64115;
	wire [4-1:0] node64116;
	wire [4-1:0] node64117;
	wire [4-1:0] node64118;
	wire [4-1:0] node64120;
	wire [4-1:0] node64123;
	wire [4-1:0] node64125;
	wire [4-1:0] node64128;
	wire [4-1:0] node64129;
	wire [4-1:0] node64130;
	wire [4-1:0] node64134;
	wire [4-1:0] node64135;
	wire [4-1:0] node64138;
	wire [4-1:0] node64141;
	wire [4-1:0] node64142;
	wire [4-1:0] node64143;
	wire [4-1:0] node64144;
	wire [4-1:0] node64147;
	wire [4-1:0] node64150;
	wire [4-1:0] node64152;
	wire [4-1:0] node64155;
	wire [4-1:0] node64156;
	wire [4-1:0] node64159;
	wire [4-1:0] node64162;
	wire [4-1:0] node64163;
	wire [4-1:0] node64164;
	wire [4-1:0] node64165;
	wire [4-1:0] node64166;
	wire [4-1:0] node64170;
	wire [4-1:0] node64172;
	wire [4-1:0] node64175;
	wire [4-1:0] node64176;
	wire [4-1:0] node64177;
	wire [4-1:0] node64181;
	wire [4-1:0] node64182;
	wire [4-1:0] node64185;
	wire [4-1:0] node64188;
	wire [4-1:0] node64189;
	wire [4-1:0] node64190;
	wire [4-1:0] node64191;
	wire [4-1:0] node64194;
	wire [4-1:0] node64197;
	wire [4-1:0] node64198;
	wire [4-1:0] node64201;
	wire [4-1:0] node64204;
	wire [4-1:0] node64205;
	wire [4-1:0] node64209;
	wire [4-1:0] node64210;
	wire [4-1:0] node64211;
	wire [4-1:0] node64212;
	wire [4-1:0] node64214;
	wire [4-1:0] node64216;
	wire [4-1:0] node64219;
	wire [4-1:0] node64221;
	wire [4-1:0] node64222;
	wire [4-1:0] node64226;
	wire [4-1:0] node64227;
	wire [4-1:0] node64228;
	wire [4-1:0] node64229;
	wire [4-1:0] node64233;
	wire [4-1:0] node64234;
	wire [4-1:0] node64237;
	wire [4-1:0] node64240;
	wire [4-1:0] node64241;
	wire [4-1:0] node64242;
	wire [4-1:0] node64245;
	wire [4-1:0] node64248;
	wire [4-1:0] node64249;
	wire [4-1:0] node64253;
	wire [4-1:0] node64254;
	wire [4-1:0] node64255;
	wire [4-1:0] node64256;
	wire [4-1:0] node64257;
	wire [4-1:0] node64261;
	wire [4-1:0] node64262;
	wire [4-1:0] node64265;
	wire [4-1:0] node64268;
	wire [4-1:0] node64270;
	wire [4-1:0] node64272;
	wire [4-1:0] node64275;
	wire [4-1:0] node64276;
	wire [4-1:0] node64278;
	wire [4-1:0] node64281;
	wire [4-1:0] node64282;
	wire [4-1:0] node64286;
	wire [4-1:0] node64287;
	wire [4-1:0] node64288;
	wire [4-1:0] node64289;
	wire [4-1:0] node64290;
	wire [4-1:0] node64291;
	wire [4-1:0] node64292;
	wire [4-1:0] node64295;
	wire [4-1:0] node64298;
	wire [4-1:0] node64299;
	wire [4-1:0] node64303;
	wire [4-1:0] node64305;
	wire [4-1:0] node64306;
	wire [4-1:0] node64309;
	wire [4-1:0] node64312;
	wire [4-1:0] node64313;
	wire [4-1:0] node64314;
	wire [4-1:0] node64317;
	wire [4-1:0] node64320;
	wire [4-1:0] node64321;
	wire [4-1:0] node64325;
	wire [4-1:0] node64326;
	wire [4-1:0] node64327;
	wire [4-1:0] node64328;
	wire [4-1:0] node64329;
	wire [4-1:0] node64332;
	wire [4-1:0] node64335;
	wire [4-1:0] node64336;
	wire [4-1:0] node64340;
	wire [4-1:0] node64341;
	wire [4-1:0] node64342;
	wire [4-1:0] node64346;
	wire [4-1:0] node64347;
	wire [4-1:0] node64351;
	wire [4-1:0] node64352;
	wire [4-1:0] node64353;
	wire [4-1:0] node64354;
	wire [4-1:0] node64357;
	wire [4-1:0] node64361;
	wire [4-1:0] node64362;
	wire [4-1:0] node64363;
	wire [4-1:0] node64366;
	wire [4-1:0] node64370;
	wire [4-1:0] node64371;
	wire [4-1:0] node64372;
	wire [4-1:0] node64373;
	wire [4-1:0] node64375;
	wire [4-1:0] node64377;
	wire [4-1:0] node64380;
	wire [4-1:0] node64381;
	wire [4-1:0] node64383;
	wire [4-1:0] node64386;
	wire [4-1:0] node64388;
	wire [4-1:0] node64391;
	wire [4-1:0] node64392;
	wire [4-1:0] node64393;
	wire [4-1:0] node64396;
	wire [4-1:0] node64399;
	wire [4-1:0] node64400;
	wire [4-1:0] node64401;
	wire [4-1:0] node64404;
	wire [4-1:0] node64407;
	wire [4-1:0] node64409;
	wire [4-1:0] node64412;
	wire [4-1:0] node64413;
	wire [4-1:0] node64414;
	wire [4-1:0] node64416;
	wire [4-1:0] node64417;
	wire [4-1:0] node64420;
	wire [4-1:0] node64423;
	wire [4-1:0] node64424;
	wire [4-1:0] node64425;
	wire [4-1:0] node64428;
	wire [4-1:0] node64432;
	wire [4-1:0] node64433;
	wire [4-1:0] node64434;
	wire [4-1:0] node64435;
	wire [4-1:0] node64438;
	wire [4-1:0] node64442;
	wire [4-1:0] node64444;
	wire [4-1:0] node64446;
	wire [4-1:0] node64449;
	wire [4-1:0] node64450;
	wire [4-1:0] node64451;
	wire [4-1:0] node64452;
	wire [4-1:0] node64453;
	wire [4-1:0] node64454;
	wire [4-1:0] node64456;
	wire [4-1:0] node64457;
	wire [4-1:0] node64460;
	wire [4-1:0] node64463;
	wire [4-1:0] node64465;
	wire [4-1:0] node64468;
	wire [4-1:0] node64469;
	wire [4-1:0] node64470;
	wire [4-1:0] node64471;
	wire [4-1:0] node64475;
	wire [4-1:0] node64476;
	wire [4-1:0] node64479;
	wire [4-1:0] node64482;
	wire [4-1:0] node64483;
	wire [4-1:0] node64486;
	wire [4-1:0] node64489;
	wire [4-1:0] node64490;
	wire [4-1:0] node64491;
	wire [4-1:0] node64494;
	wire [4-1:0] node64496;
	wire [4-1:0] node64497;
	wire [4-1:0] node64500;
	wire [4-1:0] node64503;
	wire [4-1:0] node64504;
	wire [4-1:0] node64506;
	wire [4-1:0] node64507;
	wire [4-1:0] node64510;
	wire [4-1:0] node64513;
	wire [4-1:0] node64514;
	wire [4-1:0] node64516;
	wire [4-1:0] node64519;
	wire [4-1:0] node64520;
	wire [4-1:0] node64523;
	wire [4-1:0] node64526;
	wire [4-1:0] node64527;
	wire [4-1:0] node64528;
	wire [4-1:0] node64529;
	wire [4-1:0] node64532;
	wire [4-1:0] node64533;
	wire [4-1:0] node64534;
	wire [4-1:0] node64537;
	wire [4-1:0] node64540;
	wire [4-1:0] node64542;
	wire [4-1:0] node64545;
	wire [4-1:0] node64546;
	wire [4-1:0] node64547;
	wire [4-1:0] node64548;
	wire [4-1:0] node64551;
	wire [4-1:0] node64555;
	wire [4-1:0] node64556;
	wire [4-1:0] node64557;
	wire [4-1:0] node64560;
	wire [4-1:0] node64563;
	wire [4-1:0] node64564;
	wire [4-1:0] node64567;
	wire [4-1:0] node64570;
	wire [4-1:0] node64571;
	wire [4-1:0] node64572;
	wire [4-1:0] node64574;
	wire [4-1:0] node64576;
	wire [4-1:0] node64579;
	wire [4-1:0] node64581;
	wire [4-1:0] node64582;
	wire [4-1:0] node64585;
	wire [4-1:0] node64588;
	wire [4-1:0] node64589;
	wire [4-1:0] node64590;
	wire [4-1:0] node64591;
	wire [4-1:0] node64594;
	wire [4-1:0] node64597;
	wire [4-1:0] node64598;
	wire [4-1:0] node64601;
	wire [4-1:0] node64604;
	wire [4-1:0] node64605;
	wire [4-1:0] node64608;
	wire [4-1:0] node64611;
	wire [4-1:0] node64612;
	wire [4-1:0] node64613;
	wire [4-1:0] node64614;
	wire [4-1:0] node64615;
	wire [4-1:0] node64616;
	wire [4-1:0] node64617;
	wire [4-1:0] node64620;
	wire [4-1:0] node64623;
	wire [4-1:0] node64625;
	wire [4-1:0] node64628;
	wire [4-1:0] node64629;
	wire [4-1:0] node64632;
	wire [4-1:0] node64635;
	wire [4-1:0] node64636;
	wire [4-1:0] node64637;
	wire [4-1:0] node64638;
	wire [4-1:0] node64641;
	wire [4-1:0] node64644;
	wire [4-1:0] node64645;
	wire [4-1:0] node64648;
	wire [4-1:0] node64651;
	wire [4-1:0] node64652;
	wire [4-1:0] node64653;
	wire [4-1:0] node64656;
	wire [4-1:0] node64660;
	wire [4-1:0] node64661;
	wire [4-1:0] node64662;
	wire [4-1:0] node64663;
	wire [4-1:0] node64664;
	wire [4-1:0] node64668;
	wire [4-1:0] node64669;
	wire [4-1:0] node64673;
	wire [4-1:0] node64674;
	wire [4-1:0] node64675;
	wire [4-1:0] node64679;
	wire [4-1:0] node64680;
	wire [4-1:0] node64684;
	wire [4-1:0] node64685;
	wire [4-1:0] node64686;
	wire [4-1:0] node64687;
	wire [4-1:0] node64690;
	wire [4-1:0] node64693;
	wire [4-1:0] node64694;
	wire [4-1:0] node64697;
	wire [4-1:0] node64701;
	wire [4-1:0] node64702;
	wire [4-1:0] node64703;
	wire [4-1:0] node64704;
	wire [4-1:0] node64705;
	wire [4-1:0] node64706;
	wire [4-1:0] node64709;
	wire [4-1:0] node64713;
	wire [4-1:0] node64714;
	wire [4-1:0] node64715;
	wire [4-1:0] node64719;
	wire [4-1:0] node64720;
	wire [4-1:0] node64724;
	wire [4-1:0] node64725;
	wire [4-1:0] node64726;
	wire [4-1:0] node64727;
	wire [4-1:0] node64731;
	wire [4-1:0] node64732;
	wire [4-1:0] node64736;
	wire [4-1:0] node64737;
	wire [4-1:0] node64738;
	wire [4-1:0] node64742;
	wire [4-1:0] node64743;
	wire [4-1:0] node64747;
	wire [4-1:0] node64748;
	wire [4-1:0] node64749;
	wire [4-1:0] node64750;
	wire [4-1:0] node64751;
	wire [4-1:0] node64754;
	wire [4-1:0] node64757;
	wire [4-1:0] node64758;
	wire [4-1:0] node64762;
	wire [4-1:0] node64763;
	wire [4-1:0] node64766;
	wire [4-1:0] node64769;
	wire [4-1:0] node64770;
	wire [4-1:0] node64772;
	wire [4-1:0] node64773;
	wire [4-1:0] node64776;
	wire [4-1:0] node64779;
	wire [4-1:0] node64780;
	wire [4-1:0] node64783;
	wire [4-1:0] node64786;
	wire [4-1:0] node64787;
	wire [4-1:0] node64788;
	wire [4-1:0] node64789;
	wire [4-1:0] node64790;
	wire [4-1:0] node64791;
	wire [4-1:0] node64792;
	wire [4-1:0] node64793;
	wire [4-1:0] node64794;
	wire [4-1:0] node64795;
	wire [4-1:0] node64799;
	wire [4-1:0] node64801;
	wire [4-1:0] node64804;
	wire [4-1:0] node64806;
	wire [4-1:0] node64808;
	wire [4-1:0] node64811;
	wire [4-1:0] node64812;
	wire [4-1:0] node64813;
	wire [4-1:0] node64816;
	wire [4-1:0] node64819;
	wire [4-1:0] node64820;
	wire [4-1:0] node64821;
	wire [4-1:0] node64822;
	wire [4-1:0] node64825;
	wire [4-1:0] node64829;
	wire [4-1:0] node64830;
	wire [4-1:0] node64831;
	wire [4-1:0] node64834;
	wire [4-1:0] node64837;
	wire [4-1:0] node64838;
	wire [4-1:0] node64842;
	wire [4-1:0] node64843;
	wire [4-1:0] node64844;
	wire [4-1:0] node64845;
	wire [4-1:0] node64847;
	wire [4-1:0] node64849;
	wire [4-1:0] node64852;
	wire [4-1:0] node64854;
	wire [4-1:0] node64857;
	wire [4-1:0] node64858;
	wire [4-1:0] node64859;
	wire [4-1:0] node64862;
	wire [4-1:0] node64863;
	wire [4-1:0] node64867;
	wire [4-1:0] node64868;
	wire [4-1:0] node64872;
	wire [4-1:0] node64873;
	wire [4-1:0] node64874;
	wire [4-1:0] node64876;
	wire [4-1:0] node64879;
	wire [4-1:0] node64881;
	wire [4-1:0] node64884;
	wire [4-1:0] node64885;
	wire [4-1:0] node64887;
	wire [4-1:0] node64890;
	wire [4-1:0] node64892;
	wire [4-1:0] node64895;
	wire [4-1:0] node64896;
	wire [4-1:0] node64897;
	wire [4-1:0] node64898;
	wire [4-1:0] node64899;
	wire [4-1:0] node64902;
	wire [4-1:0] node64905;
	wire [4-1:0] node64906;
	wire [4-1:0] node64907;
	wire [4-1:0] node64911;
	wire [4-1:0] node64912;
	wire [4-1:0] node64915;
	wire [4-1:0] node64918;
	wire [4-1:0] node64919;
	wire [4-1:0] node64920;
	wire [4-1:0] node64923;
	wire [4-1:0] node64926;
	wire [4-1:0] node64927;
	wire [4-1:0] node64928;
	wire [4-1:0] node64929;
	wire [4-1:0] node64932;
	wire [4-1:0] node64936;
	wire [4-1:0] node64938;
	wire [4-1:0] node64941;
	wire [4-1:0] node64942;
	wire [4-1:0] node64943;
	wire [4-1:0] node64944;
	wire [4-1:0] node64945;
	wire [4-1:0] node64948;
	wire [4-1:0] node64951;
	wire [4-1:0] node64952;
	wire [4-1:0] node64955;
	wire [4-1:0] node64958;
	wire [4-1:0] node64959;
	wire [4-1:0] node64960;
	wire [4-1:0] node64963;
	wire [4-1:0] node64966;
	wire [4-1:0] node64967;
	wire [4-1:0] node64970;
	wire [4-1:0] node64973;
	wire [4-1:0] node64974;
	wire [4-1:0] node64975;
	wire [4-1:0] node64976;
	wire [4-1:0] node64979;
	wire [4-1:0] node64982;
	wire [4-1:0] node64984;
	wire [4-1:0] node64985;
	wire [4-1:0] node64988;
	wire [4-1:0] node64991;
	wire [4-1:0] node64992;
	wire [4-1:0] node64993;
	wire [4-1:0] node64996;
	wire [4-1:0] node64999;
	wire [4-1:0] node65000;
	wire [4-1:0] node65003;
	wire [4-1:0] node65006;
	wire [4-1:0] node65007;
	wire [4-1:0] node65008;
	wire [4-1:0] node65009;
	wire [4-1:0] node65010;
	wire [4-1:0] node65011;
	wire [4-1:0] node65013;
	wire [4-1:0] node65016;
	wire [4-1:0] node65017;
	wire [4-1:0] node65021;
	wire [4-1:0] node65022;
	wire [4-1:0] node65023;
	wire [4-1:0] node65026;
	wire [4-1:0] node65029;
	wire [4-1:0] node65030;
	wire [4-1:0] node65034;
	wire [4-1:0] node65035;
	wire [4-1:0] node65036;
	wire [4-1:0] node65039;
	wire [4-1:0] node65042;
	wire [4-1:0] node65043;
	wire [4-1:0] node65046;
	wire [4-1:0] node65047;
	wire [4-1:0] node65051;
	wire [4-1:0] node65052;
	wire [4-1:0] node65053;
	wire [4-1:0] node65054;
	wire [4-1:0] node65055;
	wire [4-1:0] node65058;
	wire [4-1:0] node65060;
	wire [4-1:0] node65063;
	wire [4-1:0] node65064;
	wire [4-1:0] node65065;
	wire [4-1:0] node65068;
	wire [4-1:0] node65071;
	wire [4-1:0] node65072;
	wire [4-1:0] node65075;
	wire [4-1:0] node65078;
	wire [4-1:0] node65079;
	wire [4-1:0] node65080;
	wire [4-1:0] node65083;
	wire [4-1:0] node65086;
	wire [4-1:0] node65087;
	wire [4-1:0] node65088;
	wire [4-1:0] node65091;
	wire [4-1:0] node65094;
	wire [4-1:0] node65095;
	wire [4-1:0] node65099;
	wire [4-1:0] node65100;
	wire [4-1:0] node65101;
	wire [4-1:0] node65103;
	wire [4-1:0] node65106;
	wire [4-1:0] node65107;
	wire [4-1:0] node65108;
	wire [4-1:0] node65112;
	wire [4-1:0] node65113;
	wire [4-1:0] node65116;
	wire [4-1:0] node65119;
	wire [4-1:0] node65120;
	wire [4-1:0] node65122;
	wire [4-1:0] node65125;
	wire [4-1:0] node65126;
	wire [4-1:0] node65129;
	wire [4-1:0] node65132;
	wire [4-1:0] node65133;
	wire [4-1:0] node65134;
	wire [4-1:0] node65135;
	wire [4-1:0] node65136;
	wire [4-1:0] node65137;
	wire [4-1:0] node65138;
	wire [4-1:0] node65141;
	wire [4-1:0] node65144;
	wire [4-1:0] node65145;
	wire [4-1:0] node65148;
	wire [4-1:0] node65151;
	wire [4-1:0] node65152;
	wire [4-1:0] node65155;
	wire [4-1:0] node65158;
	wire [4-1:0] node65159;
	wire [4-1:0] node65160;
	wire [4-1:0] node65163;
	wire [4-1:0] node65166;
	wire [4-1:0] node65167;
	wire [4-1:0] node65169;
	wire [4-1:0] node65172;
	wire [4-1:0] node65173;
	wire [4-1:0] node65176;
	wire [4-1:0] node65179;
	wire [4-1:0] node65180;
	wire [4-1:0] node65181;
	wire [4-1:0] node65182;
	wire [4-1:0] node65185;
	wire [4-1:0] node65188;
	wire [4-1:0] node65190;
	wire [4-1:0] node65193;
	wire [4-1:0] node65194;
	wire [4-1:0] node65195;
	wire [4-1:0] node65196;
	wire [4-1:0] node65199;
	wire [4-1:0] node65202;
	wire [4-1:0] node65204;
	wire [4-1:0] node65207;
	wire [4-1:0] node65208;
	wire [4-1:0] node65209;
	wire [4-1:0] node65212;
	wire [4-1:0] node65215;
	wire [4-1:0] node65217;
	wire [4-1:0] node65220;
	wire [4-1:0] node65221;
	wire [4-1:0] node65222;
	wire [4-1:0] node65223;
	wire [4-1:0] node65225;
	wire [4-1:0] node65226;
	wire [4-1:0] node65229;
	wire [4-1:0] node65232;
	wire [4-1:0] node65234;
	wire [4-1:0] node65236;
	wire [4-1:0] node65239;
	wire [4-1:0] node65240;
	wire [4-1:0] node65241;
	wire [4-1:0] node65244;
	wire [4-1:0] node65247;
	wire [4-1:0] node65248;
	wire [4-1:0] node65251;
	wire [4-1:0] node65254;
	wire [4-1:0] node65255;
	wire [4-1:0] node65256;
	wire [4-1:0] node65257;
	wire [4-1:0] node65261;
	wire [4-1:0] node65262;
	wire [4-1:0] node65265;
	wire [4-1:0] node65268;
	wire [4-1:0] node65269;
	wire [4-1:0] node65270;
	wire [4-1:0] node65273;
	wire [4-1:0] node65276;
	wire [4-1:0] node65277;
	wire [4-1:0] node65278;
	wire [4-1:0] node65281;
	wire [4-1:0] node65285;
	wire [4-1:0] node65286;
	wire [4-1:0] node65287;
	wire [4-1:0] node65288;
	wire [4-1:0] node65289;
	wire [4-1:0] node65290;
	wire [4-1:0] node65291;
	wire [4-1:0] node65294;
	wire [4-1:0] node65296;
	wire [4-1:0] node65299;
	wire [4-1:0] node65300;
	wire [4-1:0] node65302;
	wire [4-1:0] node65305;
	wire [4-1:0] node65308;
	wire [4-1:0] node65309;
	wire [4-1:0] node65310;
	wire [4-1:0] node65311;
	wire [4-1:0] node65315;
	wire [4-1:0] node65316;
	wire [4-1:0] node65320;
	wire [4-1:0] node65321;
	wire [4-1:0] node65322;
	wire [4-1:0] node65326;
	wire [4-1:0] node65329;
	wire [4-1:0] node65330;
	wire [4-1:0] node65331;
	wire [4-1:0] node65332;
	wire [4-1:0] node65333;
	wire [4-1:0] node65336;
	wire [4-1:0] node65339;
	wire [4-1:0] node65340;
	wire [4-1:0] node65343;
	wire [4-1:0] node65346;
	wire [4-1:0] node65347;
	wire [4-1:0] node65350;
	wire [4-1:0] node65353;
	wire [4-1:0] node65354;
	wire [4-1:0] node65355;
	wire [4-1:0] node65356;
	wire [4-1:0] node65359;
	wire [4-1:0] node65362;
	wire [4-1:0] node65363;
	wire [4-1:0] node65364;
	wire [4-1:0] node65367;
	wire [4-1:0] node65371;
	wire [4-1:0] node65372;
	wire [4-1:0] node65373;
	wire [4-1:0] node65377;
	wire [4-1:0] node65378;
	wire [4-1:0] node65381;
	wire [4-1:0] node65384;
	wire [4-1:0] node65385;
	wire [4-1:0] node65386;
	wire [4-1:0] node65387;
	wire [4-1:0] node65388;
	wire [4-1:0] node65391;
	wire [4-1:0] node65394;
	wire [4-1:0] node65395;
	wire [4-1:0] node65396;
	wire [4-1:0] node65399;
	wire [4-1:0] node65402;
	wire [4-1:0] node65403;
	wire [4-1:0] node65407;
	wire [4-1:0] node65408;
	wire [4-1:0] node65409;
	wire [4-1:0] node65410;
	wire [4-1:0] node65413;
	wire [4-1:0] node65416;
	wire [4-1:0] node65417;
	wire [4-1:0] node65418;
	wire [4-1:0] node65421;
	wire [4-1:0] node65424;
	wire [4-1:0] node65425;
	wire [4-1:0] node65429;
	wire [4-1:0] node65430;
	wire [4-1:0] node65431;
	wire [4-1:0] node65434;
	wire [4-1:0] node65437;
	wire [4-1:0] node65438;
	wire [4-1:0] node65441;
	wire [4-1:0] node65444;
	wire [4-1:0] node65445;
	wire [4-1:0] node65446;
	wire [4-1:0] node65447;
	wire [4-1:0] node65450;
	wire [4-1:0] node65453;
	wire [4-1:0] node65455;
	wire [4-1:0] node65458;
	wire [4-1:0] node65459;
	wire [4-1:0] node65460;
	wire [4-1:0] node65461;
	wire [4-1:0] node65462;
	wire [4-1:0] node65465;
	wire [4-1:0] node65468;
	wire [4-1:0] node65469;
	wire [4-1:0] node65472;
	wire [4-1:0] node65475;
	wire [4-1:0] node65476;
	wire [4-1:0] node65479;
	wire [4-1:0] node65482;
	wire [4-1:0] node65483;
	wire [4-1:0] node65484;
	wire [4-1:0] node65489;
	wire [4-1:0] node65490;
	wire [4-1:0] node65491;
	wire [4-1:0] node65492;
	wire [4-1:0] node65493;
	wire [4-1:0] node65494;
	wire [4-1:0] node65495;
	wire [4-1:0] node65496;
	wire [4-1:0] node65500;
	wire [4-1:0] node65502;
	wire [4-1:0] node65505;
	wire [4-1:0] node65506;
	wire [4-1:0] node65509;
	wire [4-1:0] node65512;
	wire [4-1:0] node65513;
	wire [4-1:0] node65514;
	wire [4-1:0] node65518;
	wire [4-1:0] node65519;
	wire [4-1:0] node65520;
	wire [4-1:0] node65523;
	wire [4-1:0] node65526;
	wire [4-1:0] node65527;
	wire [4-1:0] node65530;
	wire [4-1:0] node65533;
	wire [4-1:0] node65534;
	wire [4-1:0] node65535;
	wire [4-1:0] node65536;
	wire [4-1:0] node65537;
	wire [4-1:0] node65540;
	wire [4-1:0] node65543;
	wire [4-1:0] node65544;
	wire [4-1:0] node65548;
	wire [4-1:0] node65549;
	wire [4-1:0] node65552;
	wire [4-1:0] node65555;
	wire [4-1:0] node65556;
	wire [4-1:0] node65559;
	wire [4-1:0] node65562;
	wire [4-1:0] node65563;
	wire [4-1:0] node65564;
	wire [4-1:0] node65565;
	wire [4-1:0] node65566;
	wire [4-1:0] node65569;
	wire [4-1:0] node65572;
	wire [4-1:0] node65573;
	wire [4-1:0] node65576;
	wire [4-1:0] node65579;
	wire [4-1:0] node65580;
	wire [4-1:0] node65581;
	wire [4-1:0] node65585;
	wire [4-1:0] node65588;
	wire [4-1:0] node65589;
	wire [4-1:0] node65590;
	wire [4-1:0] node65591;
	wire [4-1:0] node65594;
	wire [4-1:0] node65597;
	wire [4-1:0] node65598;
	wire [4-1:0] node65601;
	wire [4-1:0] node65604;
	wire [4-1:0] node65605;
	wire [4-1:0] node65606;
	wire [4-1:0] node65610;
	wire [4-1:0] node65613;
	wire [4-1:0] node65614;
	wire [4-1:0] node65615;
	wire [4-1:0] node65616;
	wire [4-1:0] node65617;
	wire [4-1:0] node65618;
	wire [4-1:0] node65619;
	wire [4-1:0] node65622;
	wire [4-1:0] node65626;
	wire [4-1:0] node65627;
	wire [4-1:0] node65630;
	wire [4-1:0] node65633;
	wire [4-1:0] node65634;
	wire [4-1:0] node65635;
	wire [4-1:0] node65638;
	wire [4-1:0] node65641;
	wire [4-1:0] node65643;
	wire [4-1:0] node65645;
	wire [4-1:0] node65648;
	wire [4-1:0] node65649;
	wire [4-1:0] node65651;
	wire [4-1:0] node65652;
	wire [4-1:0] node65655;
	wire [4-1:0] node65658;
	wire [4-1:0] node65659;
	wire [4-1:0] node65660;
	wire [4-1:0] node65663;
	wire [4-1:0] node65666;
	wire [4-1:0] node65667;
	wire [4-1:0] node65670;
	wire [4-1:0] node65673;
	wire [4-1:0] node65674;
	wire [4-1:0] node65675;
	wire [4-1:0] node65676;
	wire [4-1:0] node65677;
	wire [4-1:0] node65678;
	wire [4-1:0] node65682;
	wire [4-1:0] node65683;
	wire [4-1:0] node65686;
	wire [4-1:0] node65689;
	wire [4-1:0] node65690;
	wire [4-1:0] node65692;
	wire [4-1:0] node65695;
	wire [4-1:0] node65696;
	wire [4-1:0] node65699;
	wire [4-1:0] node65702;
	wire [4-1:0] node65703;
	wire [4-1:0] node65704;
	wire [4-1:0] node65707;
	wire [4-1:0] node65710;
	wire [4-1:0] node65712;
	wire [4-1:0] node65715;
	wire [4-1:0] node65716;
	wire [4-1:0] node65717;
	wire [4-1:0] node65720;
	wire [4-1:0] node65723;
	wire [4-1:0] node65724;
	wire [4-1:0] node65725;
	wire [4-1:0] node65727;
	wire [4-1:0] node65730;
	wire [4-1:0] node65731;
	wire [4-1:0] node65735;
	wire [4-1:0] node65736;
	wire [4-1:0] node65740;
	wire [4-1:0] node65741;
	wire [4-1:0] node65742;
	wire [4-1:0] node65743;
	wire [4-1:0] node65744;
	wire [4-1:0] node65745;
	wire [4-1:0] node65746;
	wire [4-1:0] node65747;
	wire [4-1:0] node65748;
	wire [4-1:0] node65751;
	wire [4-1:0] node65754;
	wire [4-1:0] node65755;
	wire [4-1:0] node65759;
	wire [4-1:0] node65760;
	wire [4-1:0] node65763;
	wire [4-1:0] node65766;
	wire [4-1:0] node65767;
	wire [4-1:0] node65768;
	wire [4-1:0] node65769;
	wire [4-1:0] node65770;
	wire [4-1:0] node65773;
	wire [4-1:0] node65776;
	wire [4-1:0] node65778;
	wire [4-1:0] node65781;
	wire [4-1:0] node65782;
	wire [4-1:0] node65783;
	wire [4-1:0] node65786;
	wire [4-1:0] node65790;
	wire [4-1:0] node65791;
	wire [4-1:0] node65794;
	wire [4-1:0] node65797;
	wire [4-1:0] node65798;
	wire [4-1:0] node65799;
	wire [4-1:0] node65800;
	wire [4-1:0] node65803;
	wire [4-1:0] node65806;
	wire [4-1:0] node65807;
	wire [4-1:0] node65810;
	wire [4-1:0] node65813;
	wire [4-1:0] node65814;
	wire [4-1:0] node65815;
	wire [4-1:0] node65818;
	wire [4-1:0] node65821;
	wire [4-1:0] node65822;
	wire [4-1:0] node65825;
	wire [4-1:0] node65828;
	wire [4-1:0] node65829;
	wire [4-1:0] node65830;
	wire [4-1:0] node65831;
	wire [4-1:0] node65832;
	wire [4-1:0] node65833;
	wire [4-1:0] node65836;
	wire [4-1:0] node65839;
	wire [4-1:0] node65840;
	wire [4-1:0] node65843;
	wire [4-1:0] node65844;
	wire [4-1:0] node65848;
	wire [4-1:0] node65849;
	wire [4-1:0] node65852;
	wire [4-1:0] node65855;
	wire [4-1:0] node65856;
	wire [4-1:0] node65857;
	wire [4-1:0] node65858;
	wire [4-1:0] node65859;
	wire [4-1:0] node65863;
	wire [4-1:0] node65864;
	wire [4-1:0] node65867;
	wire [4-1:0] node65870;
	wire [4-1:0] node65871;
	wire [4-1:0] node65874;
	wire [4-1:0] node65877;
	wire [4-1:0] node65878;
	wire [4-1:0] node65879;
	wire [4-1:0] node65882;
	wire [4-1:0] node65885;
	wire [4-1:0] node65887;
	wire [4-1:0] node65890;
	wire [4-1:0] node65891;
	wire [4-1:0] node65892;
	wire [4-1:0] node65893;
	wire [4-1:0] node65895;
	wire [4-1:0] node65898;
	wire [4-1:0] node65899;
	wire [4-1:0] node65902;
	wire [4-1:0] node65905;
	wire [4-1:0] node65906;
	wire [4-1:0] node65907;
	wire [4-1:0] node65910;
	wire [4-1:0] node65913;
	wire [4-1:0] node65914;
	wire [4-1:0] node65917;
	wire [4-1:0] node65920;
	wire [4-1:0] node65921;
	wire [4-1:0] node65922;
	wire [4-1:0] node65923;
	wire [4-1:0] node65926;
	wire [4-1:0] node65929;
	wire [4-1:0] node65930;
	wire [4-1:0] node65933;
	wire [4-1:0] node65936;
	wire [4-1:0] node65938;
	wire [4-1:0] node65939;
	wire [4-1:0] node65942;
	wire [4-1:0] node65945;
	wire [4-1:0] node65946;
	wire [4-1:0] node65947;
	wire [4-1:0] node65948;
	wire [4-1:0] node65949;
	wire [4-1:0] node65952;
	wire [4-1:0] node65955;
	wire [4-1:0] node65956;
	wire [4-1:0] node65957;
	wire [4-1:0] node65958;
	wire [4-1:0] node65962;
	wire [4-1:0] node65963;
	wire [4-1:0] node65966;
	wire [4-1:0] node65969;
	wire [4-1:0] node65970;
	wire [4-1:0] node65971;
	wire [4-1:0] node65974;
	wire [4-1:0] node65977;
	wire [4-1:0] node65978;
	wire [4-1:0] node65981;
	wire [4-1:0] node65984;
	wire [4-1:0] node65985;
	wire [4-1:0] node65986;
	wire [4-1:0] node65987;
	wire [4-1:0] node65988;
	wire [4-1:0] node65991;
	wire [4-1:0] node65994;
	wire [4-1:0] node65995;
	wire [4-1:0] node65998;
	wire [4-1:0] node66001;
	wire [4-1:0] node66002;
	wire [4-1:0] node66003;
	wire [4-1:0] node66006;
	wire [4-1:0] node66009;
	wire [4-1:0] node66010;
	wire [4-1:0] node66014;
	wire [4-1:0] node66015;
	wire [4-1:0] node66016;
	wire [4-1:0] node66019;
	wire [4-1:0] node66022;
	wire [4-1:0] node66023;
	wire [4-1:0] node66026;
	wire [4-1:0] node66029;
	wire [4-1:0] node66030;
	wire [4-1:0] node66031;
	wire [4-1:0] node66032;
	wire [4-1:0] node66033;
	wire [4-1:0] node66034;
	wire [4-1:0] node66037;
	wire [4-1:0] node66040;
	wire [4-1:0] node66041;
	wire [4-1:0] node66044;
	wire [4-1:0] node66047;
	wire [4-1:0] node66048;
	wire [4-1:0] node66051;
	wire [4-1:0] node66054;
	wire [4-1:0] node66055;
	wire [4-1:0] node66056;
	wire [4-1:0] node66059;
	wire [4-1:0] node66062;
	wire [4-1:0] node66063;
	wire [4-1:0] node66066;
	wire [4-1:0] node66069;
	wire [4-1:0] node66070;
	wire [4-1:0] node66071;
	wire [4-1:0] node66072;
	wire [4-1:0] node66073;
	wire [4-1:0] node66076;
	wire [4-1:0] node66080;
	wire [4-1:0] node66081;
	wire [4-1:0] node66084;
	wire [4-1:0] node66087;
	wire [4-1:0] node66088;
	wire [4-1:0] node66089;
	wire [4-1:0] node66090;
	wire [4-1:0] node66093;
	wire [4-1:0] node66096;
	wire [4-1:0] node66097;
	wire [4-1:0] node66101;
	wire [4-1:0] node66102;
	wire [4-1:0] node66105;
	wire [4-1:0] node66108;
	wire [4-1:0] node66109;
	wire [4-1:0] node66110;
	wire [4-1:0] node66111;
	wire [4-1:0] node66112;
	wire [4-1:0] node66113;
	wire [4-1:0] node66114;
	wire [4-1:0] node66116;
	wire [4-1:0] node66119;
	wire [4-1:0] node66120;
	wire [4-1:0] node66121;
	wire [4-1:0] node66124;
	wire [4-1:0] node66127;
	wire [4-1:0] node66128;
	wire [4-1:0] node66132;
	wire [4-1:0] node66133;
	wire [4-1:0] node66134;
	wire [4-1:0] node66138;
	wire [4-1:0] node66141;
	wire [4-1:0] node66142;
	wire [4-1:0] node66143;
	wire [4-1:0] node66144;
	wire [4-1:0] node66147;
	wire [4-1:0] node66150;
	wire [4-1:0] node66151;
	wire [4-1:0] node66155;
	wire [4-1:0] node66156;
	wire [4-1:0] node66157;
	wire [4-1:0] node66161;
	wire [4-1:0] node66164;
	wire [4-1:0] node66165;
	wire [4-1:0] node66166;
	wire [4-1:0] node66167;
	wire [4-1:0] node66168;
	wire [4-1:0] node66170;
	wire [4-1:0] node66173;
	wire [4-1:0] node66174;
	wire [4-1:0] node66177;
	wire [4-1:0] node66180;
	wire [4-1:0] node66182;
	wire [4-1:0] node66185;
	wire [4-1:0] node66186;
	wire [4-1:0] node66187;
	wire [4-1:0] node66188;
	wire [4-1:0] node66191;
	wire [4-1:0] node66195;
	wire [4-1:0] node66196;
	wire [4-1:0] node66198;
	wire [4-1:0] node66201;
	wire [4-1:0] node66202;
	wire [4-1:0] node66206;
	wire [4-1:0] node66207;
	wire [4-1:0] node66208;
	wire [4-1:0] node66209;
	wire [4-1:0] node66210;
	wire [4-1:0] node66213;
	wire [4-1:0] node66216;
	wire [4-1:0] node66217;
	wire [4-1:0] node66220;
	wire [4-1:0] node66223;
	wire [4-1:0] node66224;
	wire [4-1:0] node66226;
	wire [4-1:0] node66229;
	wire [4-1:0] node66230;
	wire [4-1:0] node66233;
	wire [4-1:0] node66236;
	wire [4-1:0] node66237;
	wire [4-1:0] node66238;
	wire [4-1:0] node66239;
	wire [4-1:0] node66243;
	wire [4-1:0] node66244;
	wire [4-1:0] node66248;
	wire [4-1:0] node66250;
	wire [4-1:0] node66253;
	wire [4-1:0] node66254;
	wire [4-1:0] node66255;
	wire [4-1:0] node66256;
	wire [4-1:0] node66257;
	wire [4-1:0] node66261;
	wire [4-1:0] node66264;
	wire [4-1:0] node66265;
	wire [4-1:0] node66266;
	wire [4-1:0] node66270;
	wire [4-1:0] node66273;
	wire [4-1:0] node66274;
	wire [4-1:0] node66275;
	wire [4-1:0] node66276;
	wire [4-1:0] node66280;
	wire [4-1:0] node66283;
	wire [4-1:0] node66284;
	wire [4-1:0] node66285;
	wire [4-1:0] node66287;
	wire [4-1:0] node66290;
	wire [4-1:0] node66291;
	wire [4-1:0] node66294;
	wire [4-1:0] node66297;
	wire [4-1:0] node66298;
	wire [4-1:0] node66300;
	wire [4-1:0] node66303;
	wire [4-1:0] node66304;
	wire [4-1:0] node66308;
	wire [4-1:0] node66309;
	wire [4-1:0] node66310;
	wire [4-1:0] node66311;
	wire [4-1:0] node66312;
	wire [4-1:0] node66313;
	wire [4-1:0] node66316;
	wire [4-1:0] node66319;
	wire [4-1:0] node66320;
	wire [4-1:0] node66321;
	wire [4-1:0] node66324;
	wire [4-1:0] node66327;
	wire [4-1:0] node66329;
	wire [4-1:0] node66330;
	wire [4-1:0] node66334;
	wire [4-1:0] node66335;
	wire [4-1:0] node66336;
	wire [4-1:0] node66340;
	wire [4-1:0] node66343;
	wire [4-1:0] node66344;
	wire [4-1:0] node66345;
	wire [4-1:0] node66346;
	wire [4-1:0] node66349;
	wire [4-1:0] node66352;
	wire [4-1:0] node66353;
	wire [4-1:0] node66354;
	wire [4-1:0] node66357;
	wire [4-1:0] node66360;
	wire [4-1:0] node66362;
	wire [4-1:0] node66363;
	wire [4-1:0] node66366;
	wire [4-1:0] node66369;
	wire [4-1:0] node66370;
	wire [4-1:0] node66371;
	wire [4-1:0] node66375;
	wire [4-1:0] node66378;
	wire [4-1:0] node66379;
	wire [4-1:0] node66380;
	wire [4-1:0] node66381;
	wire [4-1:0] node66382;
	wire [4-1:0] node66383;
	wire [4-1:0] node66384;
	wire [4-1:0] node66387;
	wire [4-1:0] node66390;
	wire [4-1:0] node66391;
	wire [4-1:0] node66394;
	wire [4-1:0] node66397;
	wire [4-1:0] node66398;
	wire [4-1:0] node66399;
	wire [4-1:0] node66402;
	wire [4-1:0] node66405;
	wire [4-1:0] node66406;
	wire [4-1:0] node66409;
	wire [4-1:0] node66412;
	wire [4-1:0] node66413;
	wire [4-1:0] node66414;
	wire [4-1:0] node66416;
	wire [4-1:0] node66420;
	wire [4-1:0] node66421;
	wire [4-1:0] node66424;
	wire [4-1:0] node66427;
	wire [4-1:0] node66428;
	wire [4-1:0] node66429;
	wire [4-1:0] node66433;
	wire [4-1:0] node66434;
	wire [4-1:0] node66435;
	wire [4-1:0] node66436;
	wire [4-1:0] node66441;
	wire [4-1:0] node66442;
	wire [4-1:0] node66445;
	wire [4-1:0] node66448;
	wire [4-1:0] node66449;
	wire [4-1:0] node66450;
	wire [4-1:0] node66451;
	wire [4-1:0] node66452;
	wire [4-1:0] node66453;
	wire [4-1:0] node66456;
	wire [4-1:0] node66459;
	wire [4-1:0] node66460;
	wire [4-1:0] node66463;
	wire [4-1:0] node66466;
	wire [4-1:0] node66467;
	wire [4-1:0] node66470;
	wire [4-1:0] node66473;
	wire [4-1:0] node66474;
	wire [4-1:0] node66477;
	wire [4-1:0] node66480;
	wire [4-1:0] node66481;
	wire [4-1:0] node66482;
	wire [4-1:0] node66485;
	wire [4-1:0] node66488;
	wire [4-1:0] node66489;
	wire [4-1:0] node66492;

	assign outp = (inp[6]) ? node33430 : node1;
		assign node1 = (inp[11]) ? node16585 : node2;
			assign node2 = (inp[13]) ? node8630 : node3;
				assign node3 = (inp[1]) ? node4475 : node4;
					assign node4 = (inp[2]) ? node2430 : node5;
						assign node5 = (inp[7]) ? node1279 : node6;
							assign node6 = (inp[10]) ? node608 : node7;
								assign node7 = (inp[3]) ? node299 : node8;
									assign node8 = (inp[14]) ? node138 : node9;
										assign node9 = (inp[8]) ? node99 : node10;
											assign node10 = (inp[12]) ? node52 : node11;
												assign node11 = (inp[5]) ? node31 : node12;
													assign node12 = (inp[0]) ? node18 : node13;
														assign node13 = (inp[15]) ? node15 : 4'b1111;
															assign node15 = (inp[4]) ? 4'b1101 : 4'b1001;
														assign node18 = (inp[15]) ? node24 : node19;
															assign node19 = (inp[4]) ? node21 : 4'b1001;
																assign node21 = (inp[9]) ? 4'b1101 : 4'b1001;
															assign node24 = (inp[9]) ? node28 : node25;
																assign node25 = (inp[4]) ? 4'b1011 : 4'b1111;
																assign node28 = (inp[4]) ? 4'b1111 : 4'b1011;
													assign node31 = (inp[15]) ? node39 : node32;
														assign node32 = (inp[0]) ? node34 : 4'b1011;
															assign node34 = (inp[9]) ? node36 : 4'b1001;
																assign node36 = (inp[4]) ? 4'b1111 : 4'b1001;
														assign node39 = (inp[0]) ? node47 : node40;
															assign node40 = (inp[9]) ? node44 : node41;
																assign node41 = (inp[4]) ? 4'b1001 : 4'b1101;
																assign node44 = (inp[4]) ? 4'b1111 : 4'b1001;
															assign node47 = (inp[9]) ? 4'b1011 : node48;
																assign node48 = (inp[4]) ? 4'b1011 : 4'b1111;
												assign node52 = (inp[5]) ? node74 : node53;
													assign node53 = (inp[9]) ? node63 : node54;
														assign node54 = (inp[4]) ? 4'b1001 : node55;
															assign node55 = (inp[0]) ? node59 : node56;
																assign node56 = (inp[15]) ? 4'b1101 : 4'b1111;
																assign node59 = (inp[15]) ? 4'b1111 : 4'b1101;
														assign node63 = (inp[4]) ? node69 : node64;
															assign node64 = (inp[15]) ? node66 : 4'b1001;
																assign node66 = (inp[0]) ? 4'b1011 : 4'b1001;
															assign node69 = (inp[0]) ? node71 : 4'b1111;
																assign node71 = (inp[15]) ? 4'b1111 : 4'b1101;
													assign node74 = (inp[0]) ? node86 : node75;
														assign node75 = (inp[4]) ? node79 : node76;
															assign node76 = (inp[9]) ? 4'b1011 : 4'b1111;
															assign node79 = (inp[9]) ? node83 : node80;
																assign node80 = (inp[15]) ? 4'b1001 : 4'b1011;
																assign node83 = (inp[15]) ? 4'b1111 : 4'b1101;
														assign node86 = (inp[15]) ? node94 : node87;
															assign node87 = (inp[9]) ? node91 : node88;
																assign node88 = (inp[4]) ? 4'b1001 : 4'b1101;
																assign node91 = (inp[4]) ? 4'b1111 : 4'b1001;
															assign node94 = (inp[9]) ? 4'b1101 : node95;
																assign node95 = (inp[4]) ? 4'b1011 : 4'b1111;
											assign node99 = (inp[9]) ? node115 : node100;
												assign node100 = (inp[4]) ? node108 : node101;
													assign node101 = (inp[0]) ? node105 : node102;
														assign node102 = (inp[15]) ? 4'b1100 : 4'b1110;
														assign node105 = (inp[15]) ? 4'b1110 : 4'b1100;
													assign node108 = (inp[0]) ? node112 : node109;
														assign node109 = (inp[15]) ? 4'b1000 : 4'b1010;
														assign node112 = (inp[15]) ? 4'b1010 : 4'b1000;
												assign node115 = (inp[4]) ? node123 : node116;
													assign node116 = (inp[0]) ? node120 : node117;
														assign node117 = (inp[15]) ? 4'b1000 : 4'b1010;
														assign node120 = (inp[15]) ? 4'b1010 : 4'b1000;
													assign node123 = (inp[0]) ? node131 : node124;
														assign node124 = (inp[5]) ? node128 : node125;
															assign node125 = (inp[15]) ? 4'b1100 : 4'b1110;
															assign node128 = (inp[15]) ? 4'b1110 : 4'b1100;
														assign node131 = (inp[15]) ? node135 : node132;
															assign node132 = (inp[5]) ? 4'b1110 : 4'b1100;
															assign node135 = (inp[5]) ? 4'b1100 : 4'b1110;
										assign node138 = (inp[8]) ? node236 : node139;
											assign node139 = (inp[5]) ? node193 : node140;
												assign node140 = (inp[12]) ? node166 : node141;
													assign node141 = (inp[0]) ? node153 : node142;
														assign node142 = (inp[15]) ? node148 : node143;
															assign node143 = (inp[9]) ? 4'b1110 : node144;
																assign node144 = (inp[4]) ? 4'b1010 : 4'b1110;
															assign node148 = (inp[4]) ? node150 : 4'b1000;
																assign node150 = (inp[9]) ? 4'b1100 : 4'b1000;
														assign node153 = (inp[15]) ? node161 : node154;
															assign node154 = (inp[4]) ? node158 : node155;
																assign node155 = (inp[9]) ? 4'b1000 : 4'b1100;
																assign node158 = (inp[9]) ? 4'b1100 : 4'b1000;
															assign node161 = (inp[9]) ? node163 : 4'b1110;
																assign node163 = (inp[4]) ? 4'b1110 : 4'b1010;
													assign node166 = (inp[15]) ? node178 : node167;
														assign node167 = (inp[0]) ? node173 : node168;
															assign node168 = (inp[9]) ? node170 : 4'b1010;
																assign node170 = (inp[4]) ? 4'b1110 : 4'b1010;
															assign node173 = (inp[4]) ? 4'b1000 : node174;
																assign node174 = (inp[9]) ? 4'b1000 : 4'b1100;
														assign node178 = (inp[0]) ? node186 : node179;
															assign node179 = (inp[9]) ? node183 : node180;
																assign node180 = (inp[4]) ? 4'b1000 : 4'b1100;
																assign node183 = (inp[4]) ? 4'b1100 : 4'b1000;
															assign node186 = (inp[4]) ? node190 : node187;
																assign node187 = (inp[9]) ? 4'b1010 : 4'b1110;
																assign node190 = (inp[9]) ? 4'b1110 : 4'b1010;
												assign node193 = (inp[12]) ? node213 : node194;
													assign node194 = (inp[4]) ? node206 : node195;
														assign node195 = (inp[9]) ? node201 : node196;
															assign node196 = (inp[15]) ? 4'b1110 : node197;
																assign node197 = (inp[0]) ? 4'b1100 : 4'b1110;
															assign node201 = (inp[15]) ? node203 : 4'b1000;
																assign node203 = (inp[0]) ? 4'b1010 : 4'b1000;
														assign node206 = (inp[9]) ? node208 : 4'b1000;
															assign node208 = (inp[15]) ? 4'b1100 : node209;
																assign node209 = (inp[0]) ? 4'b1110 : 4'b1100;
													assign node213 = (inp[15]) ? node229 : node214;
														assign node214 = (inp[0]) ? node222 : node215;
															assign node215 = (inp[4]) ? node219 : node216;
																assign node216 = (inp[9]) ? 4'b1010 : 4'b1110;
																assign node219 = (inp[9]) ? 4'b1100 : 4'b1010;
															assign node222 = (inp[9]) ? node226 : node223;
																assign node223 = (inp[4]) ? 4'b1000 : 4'b1100;
																assign node226 = (inp[4]) ? 4'b1110 : 4'b1000;
														assign node229 = (inp[9]) ? 4'b1100 : node230;
															assign node230 = (inp[4]) ? 4'b1010 : node231;
																assign node231 = (inp[0]) ? 4'b1110 : 4'b1100;
											assign node236 = (inp[5]) ? node276 : node237;
												assign node237 = (inp[9]) ? node255 : node238;
													assign node238 = (inp[4]) ? node246 : node239;
														assign node239 = (inp[0]) ? node243 : node240;
															assign node240 = (inp[15]) ? 4'b1101 : 4'b1111;
															assign node243 = (inp[15]) ? 4'b1111 : 4'b1101;
														assign node246 = (inp[12]) ? 4'b1001 : node247;
															assign node247 = (inp[15]) ? node251 : node248;
																assign node248 = (inp[0]) ? 4'b1001 : 4'b1011;
																assign node251 = (inp[0]) ? 4'b1011 : 4'b1001;
													assign node255 = (inp[4]) ? node263 : node256;
														assign node256 = (inp[0]) ? node260 : node257;
															assign node257 = (inp[15]) ? 4'b1001 : 4'b1011;
															assign node260 = (inp[15]) ? 4'b1011 : 4'b1001;
														assign node263 = (inp[12]) ? node271 : node264;
															assign node264 = (inp[15]) ? node268 : node265;
																assign node265 = (inp[0]) ? 4'b1101 : 4'b1111;
																assign node268 = (inp[0]) ? 4'b1111 : 4'b1101;
															assign node271 = (inp[0]) ? node273 : 4'b1111;
																assign node273 = (inp[15]) ? 4'b1111 : 4'b1101;
												assign node276 = (inp[0]) ? node286 : node277;
													assign node277 = (inp[15]) ? 4'b1111 : node278;
														assign node278 = (inp[4]) ? node282 : node279;
															assign node279 = (inp[9]) ? 4'b1011 : 4'b1111;
															assign node282 = (inp[9]) ? 4'b1101 : 4'b1011;
													assign node286 = (inp[15]) ? node292 : node287;
														assign node287 = (inp[12]) ? 4'b1001 : node288;
															assign node288 = (inp[9]) ? 4'b1111 : 4'b1101;
														assign node292 = (inp[12]) ? node294 : 4'b1011;
															assign node294 = (inp[9]) ? 4'b1101 : node295;
																assign node295 = (inp[4]) ? 4'b1011 : 4'b1111;
									assign node299 = (inp[14]) ? node453 : node300;
										assign node300 = (inp[8]) ? node362 : node301;
											assign node301 = (inp[5]) ? node333 : node302;
												assign node302 = (inp[0]) ? node318 : node303;
													assign node303 = (inp[15]) ? node311 : node304;
														assign node304 = (inp[4]) ? node308 : node305;
															assign node305 = (inp[9]) ? 4'b1011 : 4'b1111;
															assign node308 = (inp[9]) ? 4'b1101 : 4'b1011;
														assign node311 = (inp[9]) ? node315 : node312;
															assign node312 = (inp[4]) ? 4'b1001 : 4'b1101;
															assign node315 = (inp[4]) ? 4'b1111 : 4'b1001;
													assign node318 = (inp[15]) ? node326 : node319;
														assign node319 = (inp[9]) ? node323 : node320;
															assign node320 = (inp[4]) ? 4'b1001 : 4'b1101;
															assign node323 = (inp[4]) ? 4'b1111 : 4'b1001;
														assign node326 = (inp[4]) ? node330 : node327;
															assign node327 = (inp[9]) ? 4'b1011 : 4'b1111;
															assign node330 = (inp[9]) ? 4'b1101 : 4'b1011;
												assign node333 = (inp[15]) ? node347 : node334;
													assign node334 = (inp[0]) ? node342 : node335;
														assign node335 = (inp[4]) ? node339 : node336;
															assign node336 = (inp[9]) ? 4'b1001 : 4'b1101;
															assign node339 = (inp[9]) ? 4'b1101 : 4'b1001;
														assign node342 = (inp[9]) ? node344 : 4'b1011;
															assign node344 = (inp[4]) ? 4'b1111 : 4'b1011;
													assign node347 = (inp[0]) ? node355 : node348;
														assign node348 = (inp[9]) ? node352 : node349;
															assign node349 = (inp[4]) ? 4'b1011 : 4'b1111;
															assign node352 = (inp[4]) ? 4'b1111 : 4'b1011;
														assign node355 = (inp[9]) ? node359 : node356;
															assign node356 = (inp[4]) ? 4'b1001 : 4'b1101;
															assign node359 = (inp[4]) ? 4'b1101 : 4'b1001;
											assign node362 = (inp[12]) ? node412 : node363;
												assign node363 = (inp[0]) ? node389 : node364;
													assign node364 = (inp[5]) ? node376 : node365;
														assign node365 = (inp[15]) ? node371 : node366;
															assign node366 = (inp[9]) ? 4'b1100 : node367;
																assign node367 = (inp[4]) ? 4'b1010 : 4'b1110;
															assign node371 = (inp[4]) ? 4'b1000 : node372;
																assign node372 = (inp[9]) ? 4'b1000 : 4'b1100;
														assign node376 = (inp[15]) ? node382 : node377;
															assign node377 = (inp[4]) ? node379 : 4'b1000;
																assign node379 = (inp[9]) ? 4'b1100 : 4'b1000;
															assign node382 = (inp[9]) ? node386 : node383;
																assign node383 = (inp[4]) ? 4'b1010 : 4'b1110;
																assign node386 = (inp[4]) ? 4'b1110 : 4'b1010;
													assign node389 = (inp[4]) ? node401 : node390;
														assign node390 = (inp[9]) ? node396 : node391;
															assign node391 = (inp[5]) ? 4'b1110 : node392;
																assign node392 = (inp[15]) ? 4'b1110 : 4'b1100;
															assign node396 = (inp[15]) ? 4'b1010 : node397;
																assign node397 = (inp[5]) ? 4'b1010 : 4'b1000;
														assign node401 = (inp[9]) ? node409 : node402;
															assign node402 = (inp[5]) ? node406 : node403;
																assign node403 = (inp[15]) ? 4'b1010 : 4'b1000;
																assign node406 = (inp[15]) ? 4'b1000 : 4'b1010;
															assign node409 = (inp[15]) ? 4'b1100 : 4'b1110;
												assign node412 = (inp[5]) ? node432 : node413;
													assign node413 = (inp[0]) ? node421 : node414;
														assign node414 = (inp[9]) ? node416 : 4'b1110;
															assign node416 = (inp[4]) ? 4'b1110 : node417;
																assign node417 = (inp[15]) ? 4'b1000 : 4'b1010;
														assign node421 = (inp[9]) ? node425 : node422;
															assign node422 = (inp[4]) ? 4'b1000 : 4'b1100;
															assign node425 = (inp[4]) ? node429 : node426;
																assign node426 = (inp[15]) ? 4'b1010 : 4'b1000;
																assign node429 = (inp[15]) ? 4'b1100 : 4'b1110;
													assign node432 = (inp[9]) ? node444 : node433;
														assign node433 = (inp[4]) ? node439 : node434;
															assign node434 = (inp[0]) ? 4'b1110 : node435;
																assign node435 = (inp[15]) ? 4'b1110 : 4'b1100;
															assign node439 = (inp[0]) ? node441 : 4'b1000;
																assign node441 = (inp[15]) ? 4'b1000 : 4'b1010;
														assign node444 = (inp[4]) ? node446 : 4'b1000;
															assign node446 = (inp[0]) ? node450 : node447;
																assign node447 = (inp[15]) ? 4'b1110 : 4'b1100;
																assign node450 = (inp[15]) ? 4'b1100 : 4'b1110;
										assign node453 = (inp[8]) ? node507 : node454;
											assign node454 = (inp[15]) ? node478 : node455;
												assign node455 = (inp[0]) ? node469 : node456;
													assign node456 = (inp[5]) ? node462 : node457;
														assign node457 = (inp[9]) ? 4'b1100 : node458;
															assign node458 = (inp[4]) ? 4'b1010 : 4'b1110;
														assign node462 = (inp[4]) ? node466 : node463;
															assign node463 = (inp[9]) ? 4'b1000 : 4'b1100;
															assign node466 = (inp[9]) ? 4'b1100 : 4'b1000;
													assign node469 = (inp[5]) ? node473 : node470;
														assign node470 = (inp[12]) ? 4'b1000 : 4'b1100;
														assign node473 = (inp[4]) ? 4'b1110 : node474;
															assign node474 = (inp[9]) ? 4'b1010 : 4'b1110;
												assign node478 = (inp[5]) ? node494 : node479;
													assign node479 = (inp[0]) ? node487 : node480;
														assign node480 = (inp[9]) ? node484 : node481;
															assign node481 = (inp[4]) ? 4'b1000 : 4'b1100;
															assign node484 = (inp[4]) ? 4'b1110 : 4'b1000;
														assign node487 = (inp[9]) ? node491 : node488;
															assign node488 = (inp[4]) ? 4'b1010 : 4'b1110;
															assign node491 = (inp[4]) ? 4'b1100 : 4'b1010;
													assign node494 = (inp[0]) ? node500 : node495;
														assign node495 = (inp[9]) ? node497 : 4'b1010;
															assign node497 = (inp[4]) ? 4'b1110 : 4'b1010;
														assign node500 = (inp[9]) ? node504 : node501;
															assign node501 = (inp[4]) ? 4'b1000 : 4'b1100;
															assign node504 = (inp[4]) ? 4'b1100 : 4'b1000;
											assign node507 = (inp[5]) ? node551 : node508;
												assign node508 = (inp[4]) ? node530 : node509;
													assign node509 = (inp[9]) ? node517 : node510;
														assign node510 = (inp[0]) ? node514 : node511;
															assign node511 = (inp[15]) ? 4'b1101 : 4'b1111;
															assign node514 = (inp[15]) ? 4'b1111 : 4'b1101;
														assign node517 = (inp[12]) ? node523 : node518;
															assign node518 = (inp[15]) ? node520 : 4'b1011;
																assign node520 = (inp[0]) ? 4'b1011 : 4'b1001;
															assign node523 = (inp[15]) ? node527 : node524;
																assign node524 = (inp[0]) ? 4'b1001 : 4'b1011;
																assign node527 = (inp[0]) ? 4'b1011 : 4'b1001;
													assign node530 = (inp[9]) ? node536 : node531;
														assign node531 = (inp[15]) ? 4'b1001 : node532;
															assign node532 = (inp[0]) ? 4'b1001 : 4'b1011;
														assign node536 = (inp[12]) ? node544 : node537;
															assign node537 = (inp[0]) ? node541 : node538;
																assign node538 = (inp[15]) ? 4'b1111 : 4'b1101;
																assign node541 = (inp[15]) ? 4'b1101 : 4'b1111;
															assign node544 = (inp[15]) ? node548 : node545;
																assign node545 = (inp[0]) ? 4'b1111 : 4'b1101;
																assign node548 = (inp[0]) ? 4'b1101 : 4'b1111;
												assign node551 = (inp[12]) ? node579 : node552;
													assign node552 = (inp[4]) ? node564 : node553;
														assign node553 = (inp[9]) ? node559 : node554;
															assign node554 = (inp[15]) ? 4'b1111 : node555;
																assign node555 = (inp[0]) ? 4'b1111 : 4'b1101;
															assign node559 = (inp[0]) ? node561 : 4'b1011;
																assign node561 = (inp[15]) ? 4'b1001 : 4'b1011;
														assign node564 = (inp[9]) ? node572 : node565;
															assign node565 = (inp[0]) ? node569 : node566;
																assign node566 = (inp[15]) ? 4'b1011 : 4'b1001;
																assign node569 = (inp[15]) ? 4'b1001 : 4'b1011;
															assign node572 = (inp[0]) ? node576 : node573;
																assign node573 = (inp[15]) ? 4'b1111 : 4'b1101;
																assign node576 = (inp[15]) ? 4'b1101 : 4'b1111;
													assign node579 = (inp[15]) ? node595 : node580;
														assign node580 = (inp[0]) ? node588 : node581;
															assign node581 = (inp[9]) ? node585 : node582;
																assign node582 = (inp[4]) ? 4'b1001 : 4'b1101;
																assign node585 = (inp[4]) ? 4'b1101 : 4'b1001;
															assign node588 = (inp[4]) ? node592 : node589;
																assign node589 = (inp[9]) ? 4'b1011 : 4'b1111;
																assign node592 = (inp[9]) ? 4'b1111 : 4'b1011;
														assign node595 = (inp[0]) ? node601 : node596;
															assign node596 = (inp[9]) ? 4'b1011 : node597;
																assign node597 = (inp[4]) ? 4'b1011 : 4'b1111;
															assign node601 = (inp[4]) ? node605 : node602;
																assign node602 = (inp[9]) ? 4'b1001 : 4'b1101;
																assign node605 = (inp[9]) ? 4'b1101 : 4'b1001;
								assign node608 = (inp[8]) ? node964 : node609;
									assign node609 = (inp[14]) ? node799 : node610;
										assign node610 = (inp[5]) ? node710 : node611;
											assign node611 = (inp[0]) ? node663 : node612;
												assign node612 = (inp[15]) ? node638 : node613;
													assign node613 = (inp[3]) ? node627 : node614;
														assign node614 = (inp[4]) ? node620 : node615;
															assign node615 = (inp[9]) ? node617 : 4'b1111;
																assign node617 = (inp[12]) ? 4'b1111 : 4'b1011;
															assign node620 = (inp[12]) ? node624 : node621;
																assign node621 = (inp[9]) ? 4'b1111 : 4'b1011;
																assign node624 = (inp[9]) ? 4'b1011 : 4'b1111;
														assign node627 = (inp[9]) ? node633 : node628;
															assign node628 = (inp[4]) ? 4'b1011 : node629;
																assign node629 = (inp[12]) ? 4'b1011 : 4'b1111;
															assign node633 = (inp[12]) ? node635 : 4'b1101;
																assign node635 = (inp[4]) ? 4'b1001 : 4'b1101;
													assign node638 = (inp[3]) ? node654 : node639;
														assign node639 = (inp[4]) ? node647 : node640;
															assign node640 = (inp[12]) ? node644 : node641;
																assign node641 = (inp[9]) ? 4'b1001 : 4'b1101;
																assign node644 = (inp[9]) ? 4'b1101 : 4'b1001;
															assign node647 = (inp[12]) ? node651 : node648;
																assign node648 = (inp[9]) ? 4'b1101 : 4'b1001;
																assign node651 = (inp[9]) ? 4'b1001 : 4'b1101;
														assign node654 = (inp[4]) ? node656 : 4'b1001;
															assign node656 = (inp[9]) ? node660 : node657;
																assign node657 = (inp[12]) ? 4'b1111 : 4'b1001;
																assign node660 = (inp[12]) ? 4'b1011 : 4'b1111;
												assign node663 = (inp[15]) ? node691 : node664;
													assign node664 = (inp[3]) ? node680 : node665;
														assign node665 = (inp[12]) ? node673 : node666;
															assign node666 = (inp[4]) ? node670 : node667;
																assign node667 = (inp[9]) ? 4'b1001 : 4'b1101;
																assign node670 = (inp[9]) ? 4'b1101 : 4'b1001;
															assign node673 = (inp[9]) ? node677 : node674;
																assign node674 = (inp[4]) ? 4'b1101 : 4'b1001;
																assign node677 = (inp[4]) ? 4'b1001 : 4'b1101;
														assign node680 = (inp[12]) ? node686 : node681;
															assign node681 = (inp[9]) ? 4'b1001 : node682;
																assign node682 = (inp[4]) ? 4'b1001 : 4'b1101;
															assign node686 = (inp[4]) ? 4'b1111 : node687;
																assign node687 = (inp[9]) ? 4'b1111 : 4'b1001;
													assign node691 = (inp[3]) ? node701 : node692;
														assign node692 = (inp[9]) ? node694 : 4'b1111;
															assign node694 = (inp[12]) ? node698 : node695;
																assign node695 = (inp[4]) ? 4'b1111 : 4'b1011;
																assign node698 = (inp[4]) ? 4'b1011 : 4'b1111;
														assign node701 = (inp[9]) ? 4'b1101 : node702;
															assign node702 = (inp[12]) ? node706 : node703;
																assign node703 = (inp[4]) ? 4'b1011 : 4'b1111;
																assign node706 = (inp[4]) ? 4'b1101 : 4'b1011;
											assign node710 = (inp[15]) ? node760 : node711;
												assign node711 = (inp[0]) ? node735 : node712;
													assign node712 = (inp[3]) ? node726 : node713;
														assign node713 = (inp[4]) ? node719 : node714;
															assign node714 = (inp[12]) ? 4'b1011 : node715;
																assign node715 = (inp[9]) ? 4'b1011 : 4'b1111;
															assign node719 = (inp[9]) ? node723 : node720;
																assign node720 = (inp[12]) ? 4'b1101 : 4'b1011;
																assign node723 = (inp[12]) ? 4'b1001 : 4'b1101;
														assign node726 = (inp[12]) ? node728 : 4'b1001;
															assign node728 = (inp[9]) ? node732 : node729;
																assign node729 = (inp[4]) ? 4'b1101 : 4'b1001;
																assign node732 = (inp[4]) ? 4'b1001 : 4'b1101;
													assign node735 = (inp[3]) ? node751 : node736;
														assign node736 = (inp[9]) ? node744 : node737;
															assign node737 = (inp[4]) ? node741 : node738;
																assign node738 = (inp[12]) ? 4'b1001 : 4'b1101;
																assign node741 = (inp[12]) ? 4'b1111 : 4'b1001;
															assign node744 = (inp[12]) ? node748 : node745;
																assign node745 = (inp[4]) ? 4'b1111 : 4'b1001;
																assign node748 = (inp[4]) ? 4'b1011 : 4'b1111;
														assign node751 = (inp[4]) ? node753 : 4'b1111;
															assign node753 = (inp[12]) ? node757 : node754;
																assign node754 = (inp[9]) ? 4'b1111 : 4'b1011;
																assign node757 = (inp[9]) ? 4'b1011 : 4'b1111;
												assign node760 = (inp[0]) ? node784 : node761;
													assign node761 = (inp[3]) ? node771 : node762;
														assign node762 = (inp[4]) ? 4'b1111 : node763;
															assign node763 = (inp[9]) ? node767 : node764;
																assign node764 = (inp[12]) ? 4'b1001 : 4'b1101;
																assign node767 = (inp[12]) ? 4'b1111 : 4'b1001;
														assign node771 = (inp[4]) ? node779 : node772;
															assign node772 = (inp[9]) ? node776 : node773;
																assign node773 = (inp[12]) ? 4'b1011 : 4'b1111;
																assign node776 = (inp[12]) ? 4'b1111 : 4'b1011;
															assign node779 = (inp[9]) ? node781 : 4'b1111;
																assign node781 = (inp[12]) ? 4'b1011 : 4'b1111;
													assign node784 = (inp[3]) ? node796 : node785;
														assign node785 = (inp[9]) ? node791 : node786;
															assign node786 = (inp[4]) ? 4'b1011 : node787;
																assign node787 = (inp[12]) ? 4'b1011 : 4'b1111;
															assign node791 = (inp[12]) ? node793 : 4'b1011;
																assign node793 = (inp[4]) ? 4'b1001 : 4'b1101;
														assign node796 = (inp[9]) ? 4'b1101 : 4'b1001;
										assign node799 = (inp[15]) ? node873 : node800;
											assign node800 = (inp[4]) ? node834 : node801;
												assign node801 = (inp[0]) ? node819 : node802;
													assign node802 = (inp[3]) ? node810 : node803;
														assign node803 = (inp[5]) ? node807 : node804;
															assign node804 = (inp[9]) ? 4'b1110 : 4'b1010;
															assign node807 = (inp[9]) ? 4'b1010 : 4'b1110;
														assign node810 = (inp[5]) ? node814 : node811;
															assign node811 = (inp[12]) ? 4'b1010 : 4'b1110;
															assign node814 = (inp[12]) ? 4'b1000 : node815;
																assign node815 = (inp[9]) ? 4'b1000 : 4'b1100;
													assign node819 = (inp[9]) ? node823 : node820;
														assign node820 = (inp[12]) ? 4'b1000 : 4'b1100;
														assign node823 = (inp[12]) ? node829 : node824;
															assign node824 = (inp[5]) ? node826 : 4'b1000;
																assign node826 = (inp[3]) ? 4'b1010 : 4'b1000;
															assign node829 = (inp[5]) ? 4'b1110 : node830;
																assign node830 = (inp[3]) ? 4'b1110 : 4'b1100;
												assign node834 = (inp[0]) ? node858 : node835;
													assign node835 = (inp[5]) ? node849 : node836;
														assign node836 = (inp[3]) ? node844 : node837;
															assign node837 = (inp[9]) ? node841 : node838;
																assign node838 = (inp[12]) ? 4'b1110 : 4'b1010;
																assign node841 = (inp[12]) ? 4'b1010 : 4'b1110;
															assign node844 = (inp[12]) ? 4'b1100 : node845;
																assign node845 = (inp[9]) ? 4'b1100 : 4'b1010;
														assign node849 = (inp[3]) ? 4'b1100 : node850;
															assign node850 = (inp[12]) ? node854 : node851;
																assign node851 = (inp[9]) ? 4'b1100 : 4'b1010;
																assign node854 = (inp[9]) ? 4'b1000 : 4'b1100;
													assign node858 = (inp[5]) ? node866 : node859;
														assign node859 = (inp[3]) ? node861 : 4'b1100;
															assign node861 = (inp[9]) ? node863 : 4'b1000;
																assign node863 = (inp[12]) ? 4'b1010 : 4'b1110;
														assign node866 = (inp[9]) ? node870 : node867;
															assign node867 = (inp[12]) ? 4'b1110 : 4'b1010;
															assign node870 = (inp[12]) ? 4'b1010 : 4'b1110;
											assign node873 = (inp[0]) ? node915 : node874;
												assign node874 = (inp[3]) ? node894 : node875;
													assign node875 = (inp[5]) ? node889 : node876;
														assign node876 = (inp[12]) ? node884 : node877;
															assign node877 = (inp[4]) ? node881 : node878;
																assign node878 = (inp[9]) ? 4'b1000 : 4'b1100;
																assign node881 = (inp[9]) ? 4'b1100 : 4'b1000;
															assign node884 = (inp[9]) ? node886 : 4'b1100;
																assign node886 = (inp[4]) ? 4'b1000 : 4'b1100;
														assign node889 = (inp[4]) ? node891 : 4'b1000;
															assign node891 = (inp[12]) ? 4'b1010 : 4'b1000;
													assign node894 = (inp[5]) ? node908 : node895;
														assign node895 = (inp[9]) ? node901 : node896;
															assign node896 = (inp[4]) ? 4'b1000 : node897;
																assign node897 = (inp[12]) ? 4'b1000 : 4'b1100;
															assign node901 = (inp[4]) ? node905 : node902;
																assign node902 = (inp[12]) ? 4'b1110 : 4'b1000;
																assign node905 = (inp[12]) ? 4'b1010 : 4'b1110;
														assign node908 = (inp[9]) ? node910 : 4'b1110;
															assign node910 = (inp[12]) ? node912 : 4'b1010;
																assign node912 = (inp[4]) ? 4'b1010 : 4'b1110;
												assign node915 = (inp[5]) ? node945 : node916;
													assign node916 = (inp[3]) ? node932 : node917;
														assign node917 = (inp[9]) ? node925 : node918;
															assign node918 = (inp[4]) ? node922 : node919;
																assign node919 = (inp[12]) ? 4'b1010 : 4'b1110;
																assign node922 = (inp[12]) ? 4'b1110 : 4'b1010;
															assign node925 = (inp[12]) ? node929 : node926;
																assign node926 = (inp[4]) ? 4'b1110 : 4'b1010;
																assign node929 = (inp[4]) ? 4'b1010 : 4'b1110;
														assign node932 = (inp[12]) ? node938 : node933;
															assign node933 = (inp[9]) ? 4'b1010 : node934;
																assign node934 = (inp[4]) ? 4'b1010 : 4'b1110;
															assign node938 = (inp[9]) ? node942 : node939;
																assign node939 = (inp[4]) ? 4'b1100 : 4'b1010;
																assign node942 = (inp[4]) ? 4'b1000 : 4'b1100;
													assign node945 = (inp[4]) ? node953 : node946;
														assign node946 = (inp[9]) ? node948 : 4'b1010;
															assign node948 = (inp[12]) ? 4'b1100 : node949;
																assign node949 = (inp[3]) ? 4'b1000 : 4'b1010;
														assign node953 = (inp[3]) ? node959 : node954;
															assign node954 = (inp[9]) ? node956 : 4'b1100;
																assign node956 = (inp[12]) ? 4'b1000 : 4'b1100;
															assign node959 = (inp[9]) ? node961 : 4'b1000;
																assign node961 = (inp[12]) ? 4'b1000 : 4'b1100;
									assign node964 = (inp[14]) ? node1106 : node965;
										assign node965 = (inp[9]) ? node1045 : node966;
											assign node966 = (inp[15]) ? node1012 : node967;
												assign node967 = (inp[0]) ? node991 : node968;
													assign node968 = (inp[5]) ? node982 : node969;
														assign node969 = (inp[3]) ? node977 : node970;
															assign node970 = (inp[4]) ? node974 : node971;
																assign node971 = (inp[12]) ? 4'b1010 : 4'b1110;
																assign node974 = (inp[12]) ? 4'b1110 : 4'b1010;
															assign node977 = (inp[12]) ? node979 : 4'b1010;
																assign node979 = (inp[4]) ? 4'b1100 : 4'b1010;
														assign node982 = (inp[3]) ? node988 : node983;
															assign node983 = (inp[4]) ? node985 : 4'b1010;
																assign node985 = (inp[12]) ? 4'b1100 : 4'b1010;
															assign node988 = (inp[12]) ? 4'b1000 : 4'b1100;
													assign node991 = (inp[3]) ? node1001 : node992;
														assign node992 = (inp[12]) ? node996 : node993;
															assign node993 = (inp[4]) ? 4'b1000 : 4'b1100;
															assign node996 = (inp[4]) ? node998 : 4'b1000;
																assign node998 = (inp[5]) ? 4'b1110 : 4'b1100;
														assign node1001 = (inp[5]) ? node1007 : node1002;
															assign node1002 = (inp[4]) ? 4'b1110 : node1003;
																assign node1003 = (inp[12]) ? 4'b1000 : 4'b1100;
															assign node1007 = (inp[4]) ? 4'b1010 : node1008;
																assign node1008 = (inp[12]) ? 4'b1010 : 4'b1110;
												assign node1012 = (inp[0]) ? node1030 : node1013;
													assign node1013 = (inp[3]) ? node1019 : node1014;
														assign node1014 = (inp[4]) ? node1016 : 4'b1000;
															assign node1016 = (inp[12]) ? 4'b1100 : 4'b1000;
														assign node1019 = (inp[5]) ? node1025 : node1020;
															assign node1020 = (inp[12]) ? node1022 : 4'b1000;
																assign node1022 = (inp[4]) ? 4'b1110 : 4'b1000;
															assign node1025 = (inp[4]) ? 4'b1010 : node1026;
																assign node1026 = (inp[12]) ? 4'b1010 : 4'b1110;
													assign node1030 = (inp[5]) ? node1038 : node1031;
														assign node1031 = (inp[12]) ? node1035 : node1032;
															assign node1032 = (inp[4]) ? 4'b1010 : 4'b1110;
															assign node1035 = (inp[4]) ? 4'b1110 : 4'b1010;
														assign node1038 = (inp[3]) ? 4'b1000 : node1039;
															assign node1039 = (inp[4]) ? 4'b1010 : node1040;
																assign node1040 = (inp[12]) ? 4'b1010 : 4'b1110;
											assign node1045 = (inp[12]) ? node1073 : node1046;
												assign node1046 = (inp[4]) ? node1060 : node1047;
													assign node1047 = (inp[15]) ? node1049 : 4'b1000;
														assign node1049 = (inp[0]) ? node1055 : node1050;
															assign node1050 = (inp[5]) ? node1052 : 4'b1000;
																assign node1052 = (inp[3]) ? 4'b1010 : 4'b1000;
															assign node1055 = (inp[5]) ? node1057 : 4'b1010;
																assign node1057 = (inp[3]) ? 4'b1000 : 4'b1010;
													assign node1060 = (inp[15]) ? node1068 : node1061;
														assign node1061 = (inp[0]) ? node1063 : 4'b1100;
															assign node1063 = (inp[3]) ? 4'b1110 : node1064;
																assign node1064 = (inp[5]) ? 4'b1110 : 4'b1100;
														assign node1068 = (inp[0]) ? 4'b1100 : node1069;
															assign node1069 = (inp[5]) ? 4'b1110 : 4'b1100;
												assign node1073 = (inp[4]) ? node1089 : node1074;
													assign node1074 = (inp[15]) ? node1080 : node1075;
														assign node1075 = (inp[0]) ? node1077 : 4'b1100;
															assign node1077 = (inp[3]) ? 4'b1110 : 4'b1100;
														assign node1080 = (inp[0]) ? node1086 : node1081;
															assign node1081 = (inp[5]) ? 4'b1110 : node1082;
																assign node1082 = (inp[3]) ? 4'b1110 : 4'b1100;
															assign node1086 = (inp[3]) ? 4'b1100 : 4'b1110;
													assign node1089 = (inp[15]) ? node1101 : node1090;
														assign node1090 = (inp[0]) ? node1096 : node1091;
															assign node1091 = (inp[5]) ? 4'b1000 : node1092;
																assign node1092 = (inp[3]) ? 4'b1000 : 4'b1010;
															assign node1096 = (inp[3]) ? 4'b1010 : node1097;
																assign node1097 = (inp[5]) ? 4'b1010 : 4'b1000;
														assign node1101 = (inp[0]) ? node1103 : 4'b1010;
															assign node1103 = (inp[5]) ? 4'b1000 : 4'b1010;
										assign node1106 = (inp[12]) ? node1194 : node1107;
											assign node1107 = (inp[3]) ? node1149 : node1108;
												assign node1108 = (inp[5]) ? node1128 : node1109;
													assign node1109 = (inp[0]) ? node1115 : node1110;
														assign node1110 = (inp[15]) ? node1112 : 4'b1111;
															assign node1112 = (inp[4]) ? 4'b1001 : 4'b1101;
														assign node1115 = (inp[15]) ? node1121 : node1116;
															assign node1116 = (inp[9]) ? node1118 : 4'b1001;
																assign node1118 = (inp[4]) ? 4'b1101 : 4'b1001;
															assign node1121 = (inp[4]) ? node1125 : node1122;
																assign node1122 = (inp[9]) ? 4'b1011 : 4'b1111;
																assign node1125 = (inp[9]) ? 4'b1111 : 4'b1011;
													assign node1128 = (inp[0]) ? node1140 : node1129;
														assign node1129 = (inp[15]) ? node1135 : node1130;
															assign node1130 = (inp[9]) ? node1132 : 4'b1011;
																assign node1132 = (inp[4]) ? 4'b1101 : 4'b1011;
															assign node1135 = (inp[9]) ? 4'b1001 : node1136;
																assign node1136 = (inp[4]) ? 4'b1001 : 4'b1101;
														assign node1140 = (inp[15]) ? node1146 : node1141;
															assign node1141 = (inp[9]) ? node1143 : 4'b1001;
																assign node1143 = (inp[4]) ? 4'b1111 : 4'b1001;
															assign node1146 = (inp[9]) ? 4'b1011 : 4'b1111;
												assign node1149 = (inp[9]) ? node1171 : node1150;
													assign node1150 = (inp[4]) ? node1164 : node1151;
														assign node1151 = (inp[5]) ? node1159 : node1152;
															assign node1152 = (inp[15]) ? node1156 : node1153;
																assign node1153 = (inp[0]) ? 4'b1101 : 4'b1111;
																assign node1156 = (inp[0]) ? 4'b1111 : 4'b1101;
															assign node1159 = (inp[0]) ? node1161 : 4'b1111;
																assign node1161 = (inp[15]) ? 4'b1101 : 4'b1111;
														assign node1164 = (inp[0]) ? node1168 : node1165;
															assign node1165 = (inp[15]) ? 4'b1001 : 4'b1011;
															assign node1168 = (inp[15]) ? 4'b1011 : 4'b1001;
													assign node1171 = (inp[4]) ? node1187 : node1172;
														assign node1172 = (inp[15]) ? node1180 : node1173;
															assign node1173 = (inp[0]) ? node1177 : node1174;
																assign node1174 = (inp[5]) ? 4'b1001 : 4'b1011;
																assign node1177 = (inp[5]) ? 4'b1011 : 4'b1001;
															assign node1180 = (inp[0]) ? node1184 : node1181;
																assign node1181 = (inp[5]) ? 4'b1011 : 4'b1001;
																assign node1184 = (inp[5]) ? 4'b1001 : 4'b1011;
														assign node1187 = (inp[15]) ? node1191 : node1188;
															assign node1188 = (inp[0]) ? 4'b1111 : 4'b1101;
															assign node1191 = (inp[0]) ? 4'b1101 : 4'b1111;
											assign node1194 = (inp[0]) ? node1238 : node1195;
												assign node1195 = (inp[15]) ? node1219 : node1196;
													assign node1196 = (inp[5]) ? node1210 : node1197;
														assign node1197 = (inp[3]) ? node1205 : node1198;
															assign node1198 = (inp[9]) ? node1202 : node1199;
																assign node1199 = (inp[4]) ? 4'b1111 : 4'b1011;
																assign node1202 = (inp[4]) ? 4'b1011 : 4'b1111;
															assign node1205 = (inp[4]) ? 4'b1101 : node1206;
																assign node1206 = (inp[9]) ? 4'b1101 : 4'b1011;
														assign node1210 = (inp[3]) ? 4'b1001 : node1211;
															assign node1211 = (inp[4]) ? node1215 : node1212;
																assign node1212 = (inp[9]) ? 4'b1101 : 4'b1011;
																assign node1215 = (inp[9]) ? 4'b1001 : 4'b1101;
													assign node1219 = (inp[4]) ? node1231 : node1220;
														assign node1220 = (inp[9]) ? node1226 : node1221;
															assign node1221 = (inp[5]) ? node1223 : 4'b1001;
																assign node1223 = (inp[3]) ? 4'b1011 : 4'b1001;
															assign node1226 = (inp[3]) ? 4'b1111 : node1227;
																assign node1227 = (inp[5]) ? 4'b1111 : 4'b1101;
														assign node1231 = (inp[9]) ? node1233 : 4'b1111;
															assign node1233 = (inp[5]) ? 4'b1011 : node1234;
																assign node1234 = (inp[3]) ? 4'b1011 : 4'b1001;
												assign node1238 = (inp[15]) ? node1262 : node1239;
													assign node1239 = (inp[3]) ? node1253 : node1240;
														assign node1240 = (inp[5]) ? node1248 : node1241;
															assign node1241 = (inp[4]) ? node1245 : node1242;
																assign node1242 = (inp[9]) ? 4'b1101 : 4'b1001;
																assign node1245 = (inp[9]) ? 4'b1001 : 4'b1101;
															assign node1248 = (inp[9]) ? node1250 : 4'b1001;
																assign node1250 = (inp[4]) ? 4'b1011 : 4'b1111;
														assign node1253 = (inp[5]) ? 4'b1011 : node1254;
															assign node1254 = (inp[4]) ? node1258 : node1255;
																assign node1255 = (inp[9]) ? 4'b1111 : 4'b1001;
																assign node1258 = (inp[9]) ? 4'b1011 : 4'b1111;
													assign node1262 = (inp[5]) ? node1270 : node1263;
														assign node1263 = (inp[4]) ? node1265 : 4'b1011;
															assign node1265 = (inp[9]) ? node1267 : 4'b1101;
																assign node1267 = (inp[3]) ? 4'b1001 : 4'b1011;
														assign node1270 = (inp[4]) ? node1276 : node1271;
															assign node1271 = (inp[9]) ? 4'b1101 : node1272;
																assign node1272 = (inp[3]) ? 4'b1001 : 4'b1011;
															assign node1276 = (inp[9]) ? 4'b1001 : 4'b1101;
							assign node1279 = (inp[8]) ? node1853 : node1280;
								assign node1280 = (inp[14]) ? node1548 : node1281;
									assign node1281 = (inp[9]) ? node1403 : node1282;
										assign node1282 = (inp[4]) ? node1336 : node1283;
											assign node1283 = (inp[10]) ? node1311 : node1284;
												assign node1284 = (inp[5]) ? node1296 : node1285;
													assign node1285 = (inp[12]) ? node1291 : node1286;
														assign node1286 = (inp[15]) ? node1288 : 4'b1110;
															assign node1288 = (inp[0]) ? 4'b1110 : 4'b1100;
														assign node1291 = (inp[15]) ? node1293 : 4'b1100;
															assign node1293 = (inp[0]) ? 4'b1110 : 4'b1100;
													assign node1296 = (inp[0]) ? node1304 : node1297;
														assign node1297 = (inp[3]) ? node1301 : node1298;
															assign node1298 = (inp[15]) ? 4'b1100 : 4'b1110;
															assign node1301 = (inp[15]) ? 4'b1110 : 4'b1100;
														assign node1304 = (inp[15]) ? node1308 : node1305;
															assign node1305 = (inp[3]) ? 4'b1110 : 4'b1100;
															assign node1308 = (inp[3]) ? 4'b1100 : 4'b1110;
												assign node1311 = (inp[12]) ? node1319 : node1312;
													assign node1312 = (inp[0]) ? node1316 : node1313;
														assign node1313 = (inp[15]) ? 4'b1100 : 4'b1110;
														assign node1316 = (inp[15]) ? 4'b1110 : 4'b1100;
													assign node1319 = (inp[15]) ? node1329 : node1320;
														assign node1320 = (inp[0]) ? node1324 : node1321;
															assign node1321 = (inp[5]) ? 4'b1000 : 4'b1010;
															assign node1324 = (inp[5]) ? node1326 : 4'b1000;
																assign node1326 = (inp[3]) ? 4'b1010 : 4'b1000;
														assign node1329 = (inp[0]) ? 4'b1010 : node1330;
															assign node1330 = (inp[3]) ? node1332 : 4'b1000;
																assign node1332 = (inp[5]) ? 4'b1010 : 4'b1000;
											assign node1336 = (inp[10]) ? node1358 : node1337;
												assign node1337 = (inp[15]) ? node1349 : node1338;
													assign node1338 = (inp[0]) ? node1344 : node1339;
														assign node1339 = (inp[3]) ? node1341 : 4'b1010;
															assign node1341 = (inp[5]) ? 4'b1000 : 4'b1010;
														assign node1344 = (inp[3]) ? node1346 : 4'b1000;
															assign node1346 = (inp[5]) ? 4'b1010 : 4'b1000;
													assign node1349 = (inp[0]) ? node1353 : node1350;
														assign node1350 = (inp[3]) ? 4'b1010 : 4'b1000;
														assign node1353 = (inp[3]) ? node1355 : 4'b1010;
															assign node1355 = (inp[5]) ? 4'b1000 : 4'b1010;
												assign node1358 = (inp[12]) ? node1374 : node1359;
													assign node1359 = (inp[5]) ? node1365 : node1360;
														assign node1360 = (inp[15]) ? node1362 : 4'b1000;
															assign node1362 = (inp[0]) ? 4'b1010 : 4'b1000;
														assign node1365 = (inp[15]) ? node1367 : 4'b1010;
															assign node1367 = (inp[3]) ? node1371 : node1368;
																assign node1368 = (inp[0]) ? 4'b1010 : 4'b1000;
																assign node1371 = (inp[0]) ? 4'b1000 : 4'b1010;
													assign node1374 = (inp[5]) ? node1388 : node1375;
														assign node1375 = (inp[0]) ? node1383 : node1376;
															assign node1376 = (inp[3]) ? node1380 : node1377;
																assign node1377 = (inp[15]) ? 4'b1100 : 4'b1110;
																assign node1380 = (inp[15]) ? 4'b1110 : 4'b1100;
															assign node1383 = (inp[15]) ? node1385 : 4'b1110;
																assign node1385 = (inp[3]) ? 4'b1100 : 4'b1110;
														assign node1388 = (inp[3]) ? node1396 : node1389;
															assign node1389 = (inp[15]) ? node1393 : node1390;
																assign node1390 = (inp[0]) ? 4'b1110 : 4'b1100;
																assign node1393 = (inp[0]) ? 4'b1100 : 4'b1110;
															assign node1396 = (inp[15]) ? node1400 : node1397;
																assign node1397 = (inp[0]) ? 4'b1110 : 4'b1100;
																assign node1400 = (inp[0]) ? 4'b1100 : 4'b1110;
										assign node1403 = (inp[4]) ? node1471 : node1404;
											assign node1404 = (inp[10]) ? node1440 : node1405;
												assign node1405 = (inp[3]) ? node1425 : node1406;
													assign node1406 = (inp[5]) ? node1416 : node1407;
														assign node1407 = (inp[12]) ? 4'b1010 : node1408;
															assign node1408 = (inp[15]) ? node1412 : node1409;
																assign node1409 = (inp[0]) ? 4'b1000 : 4'b1010;
																assign node1412 = (inp[0]) ? 4'b1010 : 4'b1000;
														assign node1416 = (inp[12]) ? node1418 : 4'b1010;
															assign node1418 = (inp[0]) ? node1422 : node1419;
																assign node1419 = (inp[15]) ? 4'b1000 : 4'b1010;
																assign node1422 = (inp[15]) ? 4'b1010 : 4'b1000;
													assign node1425 = (inp[0]) ? node1435 : node1426;
														assign node1426 = (inp[12]) ? node1428 : 4'b1000;
															assign node1428 = (inp[15]) ? node1432 : node1429;
																assign node1429 = (inp[5]) ? 4'b1000 : 4'b1010;
																assign node1432 = (inp[5]) ? 4'b1010 : 4'b1000;
														assign node1435 = (inp[5]) ? node1437 : 4'b1010;
															assign node1437 = (inp[15]) ? 4'b1000 : 4'b1010;
												assign node1440 = (inp[12]) ? node1456 : node1441;
													assign node1441 = (inp[15]) ? node1447 : node1442;
														assign node1442 = (inp[0]) ? node1444 : 4'b1010;
															assign node1444 = (inp[3]) ? 4'b1010 : 4'b1000;
														assign node1447 = (inp[3]) ? node1449 : 4'b1000;
															assign node1449 = (inp[5]) ? node1453 : node1450;
																assign node1450 = (inp[0]) ? 4'b1010 : 4'b1000;
																assign node1453 = (inp[0]) ? 4'b1000 : 4'b1010;
													assign node1456 = (inp[15]) ? node1468 : node1457;
														assign node1457 = (inp[0]) ? node1463 : node1458;
															assign node1458 = (inp[5]) ? 4'b1100 : node1459;
																assign node1459 = (inp[3]) ? 4'b1100 : 4'b1110;
															assign node1463 = (inp[5]) ? 4'b1110 : node1464;
																assign node1464 = (inp[3]) ? 4'b1110 : 4'b1100;
														assign node1468 = (inp[0]) ? 4'b1100 : 4'b1110;
											assign node1471 = (inp[12]) ? node1507 : node1472;
												assign node1472 = (inp[3]) ? node1486 : node1473;
													assign node1473 = (inp[15]) ? node1479 : node1474;
														assign node1474 = (inp[5]) ? 4'b1110 : node1475;
															assign node1475 = (inp[0]) ? 4'b1100 : 4'b1110;
														assign node1479 = (inp[5]) ? node1483 : node1480;
															assign node1480 = (inp[0]) ? 4'b1110 : 4'b1100;
															assign node1483 = (inp[0]) ? 4'b1100 : 4'b1110;
													assign node1486 = (inp[5]) ? node1494 : node1487;
														assign node1487 = (inp[15]) ? node1491 : node1488;
															assign node1488 = (inp[0]) ? 4'b1110 : 4'b1100;
															assign node1491 = (inp[0]) ? 4'b1100 : 4'b1110;
														assign node1494 = (inp[10]) ? node1502 : node1495;
															assign node1495 = (inp[0]) ? node1499 : node1496;
																assign node1496 = (inp[15]) ? 4'b1110 : 4'b1100;
																assign node1499 = (inp[15]) ? 4'b1100 : 4'b1110;
															assign node1502 = (inp[15]) ? node1504 : 4'b1100;
																assign node1504 = (inp[0]) ? 4'b1100 : 4'b1110;
												assign node1507 = (inp[10]) ? node1531 : node1508;
													assign node1508 = (inp[3]) ? node1518 : node1509;
														assign node1509 = (inp[5]) ? 4'b1110 : node1510;
															assign node1510 = (inp[15]) ? node1514 : node1511;
																assign node1511 = (inp[0]) ? 4'b1100 : 4'b1110;
																assign node1514 = (inp[0]) ? 4'b1110 : 4'b1100;
														assign node1518 = (inp[5]) ? node1526 : node1519;
															assign node1519 = (inp[15]) ? node1523 : node1520;
																assign node1520 = (inp[0]) ? 4'b1110 : 4'b1100;
																assign node1523 = (inp[0]) ? 4'b1100 : 4'b1110;
															assign node1526 = (inp[0]) ? node1528 : 4'b1100;
																assign node1528 = (inp[15]) ? 4'b1100 : 4'b1110;
													assign node1531 = (inp[5]) ? node1543 : node1532;
														assign node1532 = (inp[15]) ? node1538 : node1533;
															assign node1533 = (inp[0]) ? node1535 : 4'b1000;
																assign node1535 = (inp[3]) ? 4'b1010 : 4'b1000;
															assign node1538 = (inp[3]) ? node1540 : 4'b1010;
																assign node1540 = (inp[0]) ? 4'b1000 : 4'b1010;
														assign node1543 = (inp[15]) ? node1545 : 4'b1010;
															assign node1545 = (inp[0]) ? 4'b1000 : 4'b1010;
									assign node1548 = (inp[10]) ? node1674 : node1549;
										assign node1549 = (inp[3]) ? node1615 : node1550;
											assign node1550 = (inp[0]) ? node1580 : node1551;
												assign node1551 = (inp[15]) ? node1565 : node1552;
													assign node1552 = (inp[5]) ? node1558 : node1553;
														assign node1553 = (inp[4]) ? node1555 : 4'b1011;
															assign node1555 = (inp[9]) ? 4'b1111 : 4'b1011;
														assign node1558 = (inp[4]) ? node1562 : node1559;
															assign node1559 = (inp[9]) ? 4'b1011 : 4'b1111;
															assign node1562 = (inp[9]) ? 4'b1101 : 4'b1011;
													assign node1565 = (inp[5]) ? node1573 : node1566;
														assign node1566 = (inp[4]) ? node1570 : node1567;
															assign node1567 = (inp[9]) ? 4'b1001 : 4'b1101;
															assign node1570 = (inp[9]) ? 4'b1101 : 4'b1001;
														assign node1573 = (inp[9]) ? node1577 : node1574;
															assign node1574 = (inp[4]) ? 4'b1001 : 4'b1101;
															assign node1577 = (inp[4]) ? 4'b1111 : 4'b1001;
												assign node1580 = (inp[15]) ? node1596 : node1581;
													assign node1581 = (inp[5]) ? node1589 : node1582;
														assign node1582 = (inp[4]) ? node1586 : node1583;
															assign node1583 = (inp[9]) ? 4'b1001 : 4'b1101;
															assign node1586 = (inp[9]) ? 4'b1101 : 4'b1001;
														assign node1589 = (inp[9]) ? node1593 : node1590;
															assign node1590 = (inp[4]) ? 4'b1001 : 4'b1101;
															assign node1593 = (inp[4]) ? 4'b1111 : 4'b1001;
													assign node1596 = (inp[5]) ? node1610 : node1597;
														assign node1597 = (inp[12]) ? node1605 : node1598;
															assign node1598 = (inp[4]) ? node1602 : node1599;
																assign node1599 = (inp[9]) ? 4'b1011 : 4'b1111;
																assign node1602 = (inp[9]) ? 4'b1111 : 4'b1011;
															assign node1605 = (inp[9]) ? 4'b1111 : node1606;
																assign node1606 = (inp[4]) ? 4'b1011 : 4'b1111;
														assign node1610 = (inp[4]) ? node1612 : 4'b1011;
															assign node1612 = (inp[9]) ? 4'b1101 : 4'b1011;
											assign node1615 = (inp[9]) ? node1643 : node1616;
												assign node1616 = (inp[4]) ? node1630 : node1617;
													assign node1617 = (inp[0]) ? node1623 : node1618;
														assign node1618 = (inp[5]) ? 4'b1101 : node1619;
															assign node1619 = (inp[15]) ? 4'b1101 : 4'b1111;
														assign node1623 = (inp[15]) ? node1627 : node1624;
															assign node1624 = (inp[5]) ? 4'b1111 : 4'b1101;
															assign node1627 = (inp[5]) ? 4'b1101 : 4'b1111;
													assign node1630 = (inp[15]) ? node1638 : node1631;
														assign node1631 = (inp[5]) ? node1635 : node1632;
															assign node1632 = (inp[0]) ? 4'b1001 : 4'b1011;
															assign node1635 = (inp[0]) ? 4'b1011 : 4'b1001;
														assign node1638 = (inp[5]) ? node1640 : 4'b1011;
															assign node1640 = (inp[0]) ? 4'b1001 : 4'b1011;
												assign node1643 = (inp[4]) ? node1659 : node1644;
													assign node1644 = (inp[0]) ? node1646 : 4'b1011;
														assign node1646 = (inp[12]) ? node1654 : node1647;
															assign node1647 = (inp[15]) ? node1651 : node1648;
																assign node1648 = (inp[5]) ? 4'b1011 : 4'b1001;
																assign node1651 = (inp[5]) ? 4'b1001 : 4'b1011;
															assign node1654 = (inp[5]) ? node1656 : 4'b1011;
																assign node1656 = (inp[15]) ? 4'b1001 : 4'b1011;
													assign node1659 = (inp[5]) ? node1667 : node1660;
														assign node1660 = (inp[12]) ? node1662 : 4'b1111;
															assign node1662 = (inp[15]) ? node1664 : 4'b1101;
																assign node1664 = (inp[0]) ? 4'b1101 : 4'b1111;
														assign node1667 = (inp[12]) ? 4'b1111 : node1668;
															assign node1668 = (inp[15]) ? 4'b1111 : node1669;
																assign node1669 = (inp[0]) ? 4'b1111 : 4'b1101;
										assign node1674 = (inp[0]) ? node1762 : node1675;
											assign node1675 = (inp[4]) ? node1723 : node1676;
												assign node1676 = (inp[3]) ? node1696 : node1677;
													assign node1677 = (inp[15]) ? node1685 : node1678;
														assign node1678 = (inp[5]) ? node1682 : node1679;
															assign node1679 = (inp[12]) ? 4'b1111 : 4'b1011;
															assign node1682 = (inp[9]) ? 4'b1101 : 4'b1111;
														assign node1685 = (inp[5]) ? node1693 : node1686;
															assign node1686 = (inp[9]) ? node1690 : node1687;
																assign node1687 = (inp[12]) ? 4'b1001 : 4'b1101;
																assign node1690 = (inp[12]) ? 4'b1101 : 4'b1001;
															assign node1693 = (inp[12]) ? 4'b1111 : 4'b1101;
													assign node1696 = (inp[15]) ? node1710 : node1697;
														assign node1697 = (inp[5]) ? node1703 : node1698;
															assign node1698 = (inp[9]) ? 4'b1101 : node1699;
																assign node1699 = (inp[12]) ? 4'b1011 : 4'b1111;
															assign node1703 = (inp[12]) ? node1707 : node1704;
																assign node1704 = (inp[9]) ? 4'b1001 : 4'b1101;
																assign node1707 = (inp[9]) ? 4'b1101 : 4'b1001;
														assign node1710 = (inp[5]) ? node1716 : node1711;
															assign node1711 = (inp[12]) ? 4'b1111 : node1712;
																assign node1712 = (inp[9]) ? 4'b1001 : 4'b1101;
															assign node1716 = (inp[9]) ? node1720 : node1717;
																assign node1717 = (inp[12]) ? 4'b1011 : 4'b1111;
																assign node1720 = (inp[12]) ? 4'b1111 : 4'b1011;
												assign node1723 = (inp[15]) ? node1741 : node1724;
													assign node1724 = (inp[3]) ? node1734 : node1725;
														assign node1725 = (inp[12]) ? node1729 : node1726;
															assign node1726 = (inp[9]) ? 4'b1111 : 4'b1011;
															assign node1729 = (inp[5]) ? node1731 : 4'b1011;
																assign node1731 = (inp[9]) ? 4'b1001 : 4'b1101;
														assign node1734 = (inp[12]) ? node1738 : node1735;
															assign node1735 = (inp[9]) ? 4'b1101 : 4'b1001;
															assign node1738 = (inp[9]) ? 4'b1001 : 4'b1101;
													assign node1741 = (inp[3]) ? node1753 : node1742;
														assign node1742 = (inp[5]) ? node1748 : node1743;
															assign node1743 = (inp[12]) ? node1745 : 4'b1101;
																assign node1745 = (inp[9]) ? 4'b1001 : 4'b1101;
															assign node1748 = (inp[9]) ? node1750 : 4'b1001;
																assign node1750 = (inp[12]) ? 4'b1011 : 4'b1111;
														assign node1753 = (inp[12]) ? node1759 : node1754;
															assign node1754 = (inp[9]) ? 4'b1111 : node1755;
																assign node1755 = (inp[5]) ? 4'b1011 : 4'b1001;
															assign node1759 = (inp[9]) ? 4'b1011 : 4'b1111;
											assign node1762 = (inp[15]) ? node1800 : node1763;
												assign node1763 = (inp[5]) ? node1785 : node1764;
													assign node1764 = (inp[3]) ? node1774 : node1765;
														assign node1765 = (inp[4]) ? 4'b1101 : node1766;
															assign node1766 = (inp[9]) ? node1770 : node1767;
																assign node1767 = (inp[12]) ? 4'b1001 : 4'b1101;
																assign node1770 = (inp[12]) ? 4'b1101 : 4'b1001;
														assign node1774 = (inp[4]) ? node1780 : node1775;
															assign node1775 = (inp[9]) ? 4'b1111 : node1776;
																assign node1776 = (inp[12]) ? 4'b1001 : 4'b1101;
															assign node1780 = (inp[12]) ? node1782 : 4'b1111;
																assign node1782 = (inp[9]) ? 4'b1011 : 4'b1111;
													assign node1785 = (inp[4]) ? node1795 : node1786;
														assign node1786 = (inp[12]) ? node1792 : node1787;
															assign node1787 = (inp[3]) ? node1789 : 4'b1001;
																assign node1789 = (inp[9]) ? 4'b1011 : 4'b1111;
															assign node1792 = (inp[9]) ? 4'b1111 : 4'b1011;
														assign node1795 = (inp[12]) ? node1797 : 4'b1111;
															assign node1797 = (inp[9]) ? 4'b1011 : 4'b1111;
												assign node1800 = (inp[5]) ? node1830 : node1801;
													assign node1801 = (inp[3]) ? node1817 : node1802;
														assign node1802 = (inp[4]) ? node1810 : node1803;
															assign node1803 = (inp[9]) ? node1807 : node1804;
																assign node1804 = (inp[12]) ? 4'b1011 : 4'b1111;
																assign node1807 = (inp[12]) ? 4'b1111 : 4'b1011;
															assign node1810 = (inp[12]) ? node1814 : node1811;
																assign node1811 = (inp[9]) ? 4'b1111 : 4'b1011;
																assign node1814 = (inp[9]) ? 4'b1011 : 4'b1111;
														assign node1817 = (inp[9]) ? node1825 : node1818;
															assign node1818 = (inp[4]) ? node1822 : node1819;
																assign node1819 = (inp[12]) ? 4'b1011 : 4'b1111;
																assign node1822 = (inp[12]) ? 4'b1101 : 4'b1011;
															assign node1825 = (inp[12]) ? node1827 : 4'b1101;
																assign node1827 = (inp[4]) ? 4'b1001 : 4'b1101;
													assign node1830 = (inp[12]) ? node1840 : node1831;
														assign node1831 = (inp[4]) ? 4'b1101 : node1832;
															assign node1832 = (inp[3]) ? node1836 : node1833;
																assign node1833 = (inp[9]) ? 4'b1011 : 4'b1111;
																assign node1836 = (inp[9]) ? 4'b1001 : 4'b1101;
														assign node1840 = (inp[3]) ? node1846 : node1841;
															assign node1841 = (inp[9]) ? node1843 : 4'b1101;
																assign node1843 = (inp[4]) ? 4'b1001 : 4'b1101;
															assign node1846 = (inp[4]) ? node1850 : node1847;
																assign node1847 = (inp[9]) ? 4'b1101 : 4'b1001;
																assign node1850 = (inp[9]) ? 4'b1001 : 4'b1101;
								assign node1853 = (inp[14]) ? node2119 : node1854;
									assign node1854 = (inp[5]) ? node1966 : node1855;
										assign node1855 = (inp[9]) ? node1909 : node1856;
											assign node1856 = (inp[4]) ? node1876 : node1857;
												assign node1857 = (inp[10]) ? node1865 : node1858;
													assign node1858 = (inp[0]) ? node1862 : node1859;
														assign node1859 = (inp[15]) ? 4'b1101 : 4'b1111;
														assign node1862 = (inp[15]) ? 4'b1111 : 4'b1101;
													assign node1865 = (inp[12]) ? node1871 : node1866;
														assign node1866 = (inp[15]) ? 4'b1111 : node1867;
															assign node1867 = (inp[3]) ? 4'b1101 : 4'b1111;
														assign node1871 = (inp[0]) ? node1873 : 4'b1001;
															assign node1873 = (inp[15]) ? 4'b1011 : 4'b1001;
												assign node1876 = (inp[10]) ? node1884 : node1877;
													assign node1877 = (inp[15]) ? node1881 : node1878;
														assign node1878 = (inp[0]) ? 4'b1001 : 4'b1011;
														assign node1881 = (inp[0]) ? 4'b1011 : 4'b1001;
													assign node1884 = (inp[12]) ? node1894 : node1885;
														assign node1885 = (inp[3]) ? node1889 : node1886;
															assign node1886 = (inp[15]) ? 4'b1011 : 4'b1001;
															assign node1889 = (inp[15]) ? 4'b1001 : node1890;
																assign node1890 = (inp[0]) ? 4'b1001 : 4'b1011;
														assign node1894 = (inp[0]) ? node1902 : node1895;
															assign node1895 = (inp[15]) ? node1899 : node1896;
																assign node1896 = (inp[3]) ? 4'b1101 : 4'b1111;
																assign node1899 = (inp[3]) ? 4'b1111 : 4'b1101;
															assign node1902 = (inp[15]) ? node1906 : node1903;
																assign node1903 = (inp[3]) ? 4'b1111 : 4'b1101;
																assign node1906 = (inp[3]) ? 4'b1101 : 4'b1111;
											assign node1909 = (inp[4]) ? node1933 : node1910;
												assign node1910 = (inp[12]) ? node1918 : node1911;
													assign node1911 = (inp[15]) ? node1915 : node1912;
														assign node1912 = (inp[0]) ? 4'b1001 : 4'b1011;
														assign node1915 = (inp[0]) ? 4'b1011 : 4'b1001;
													assign node1918 = (inp[10]) ? node1924 : node1919;
														assign node1919 = (inp[0]) ? 4'b1001 : node1920;
															assign node1920 = (inp[15]) ? 4'b1001 : 4'b1011;
														assign node1924 = (inp[15]) ? node1926 : 4'b1101;
															assign node1926 = (inp[0]) ? node1930 : node1927;
																assign node1927 = (inp[3]) ? 4'b1111 : 4'b1101;
																assign node1930 = (inp[3]) ? 4'b1101 : 4'b1111;
												assign node1933 = (inp[10]) ? node1951 : node1934;
													assign node1934 = (inp[0]) ? 4'b1101 : node1935;
														assign node1935 = (inp[12]) ? node1943 : node1936;
															assign node1936 = (inp[15]) ? node1940 : node1937;
																assign node1937 = (inp[3]) ? 4'b1101 : 4'b1111;
																assign node1940 = (inp[3]) ? 4'b1111 : 4'b1101;
															assign node1943 = (inp[3]) ? node1947 : node1944;
																assign node1944 = (inp[15]) ? 4'b1101 : 4'b1111;
																assign node1947 = (inp[15]) ? 4'b1111 : 4'b1101;
													assign node1951 = (inp[12]) ? node1959 : node1952;
														assign node1952 = (inp[3]) ? node1954 : 4'b1101;
															assign node1954 = (inp[15]) ? 4'b1111 : node1955;
																assign node1955 = (inp[0]) ? 4'b1111 : 4'b1101;
														assign node1959 = (inp[0]) ? 4'b1011 : node1960;
															assign node1960 = (inp[15]) ? 4'b1001 : node1961;
																assign node1961 = (inp[3]) ? 4'b1001 : 4'b1011;
										assign node1966 = (inp[10]) ? node2040 : node1967;
											assign node1967 = (inp[0]) ? node1999 : node1968;
												assign node1968 = (inp[15]) ? node1984 : node1969;
													assign node1969 = (inp[3]) ? node1979 : node1970;
														assign node1970 = (inp[12]) ? node1974 : node1971;
															assign node1971 = (inp[9]) ? 4'b1101 : 4'b1111;
															assign node1974 = (inp[9]) ? 4'b1011 : node1975;
																assign node1975 = (inp[4]) ? 4'b1011 : 4'b1111;
														assign node1979 = (inp[4]) ? node1981 : 4'b1101;
															assign node1981 = (inp[9]) ? 4'b1101 : 4'b1001;
													assign node1984 = (inp[3]) ? node1992 : node1985;
														assign node1985 = (inp[12]) ? node1987 : 4'b1001;
															assign node1987 = (inp[4]) ? 4'b1111 : node1988;
																assign node1988 = (inp[9]) ? 4'b1001 : 4'b1101;
														assign node1992 = (inp[4]) ? node1996 : node1993;
															assign node1993 = (inp[9]) ? 4'b1011 : 4'b1111;
															assign node1996 = (inp[9]) ? 4'b1111 : 4'b1011;
												assign node1999 = (inp[15]) ? node2017 : node2000;
													assign node2000 = (inp[3]) ? node2008 : node2001;
														assign node2001 = (inp[4]) ? node2005 : node2002;
															assign node2002 = (inp[9]) ? 4'b1001 : 4'b1101;
															assign node2005 = (inp[9]) ? 4'b1111 : 4'b1001;
														assign node2008 = (inp[12]) ? 4'b1111 : node2009;
															assign node2009 = (inp[9]) ? node2013 : node2010;
																assign node2010 = (inp[4]) ? 4'b1011 : 4'b1111;
																assign node2013 = (inp[4]) ? 4'b1111 : 4'b1011;
													assign node2017 = (inp[3]) ? node2025 : node2018;
														assign node2018 = (inp[4]) ? node2022 : node2019;
															assign node2019 = (inp[9]) ? 4'b1011 : 4'b1111;
															assign node2022 = (inp[9]) ? 4'b1101 : 4'b1011;
														assign node2025 = (inp[12]) ? node2033 : node2026;
															assign node2026 = (inp[9]) ? node2030 : node2027;
																assign node2027 = (inp[4]) ? 4'b1001 : 4'b1101;
																assign node2030 = (inp[4]) ? 4'b1101 : 4'b1001;
															assign node2033 = (inp[4]) ? node2037 : node2034;
																assign node2034 = (inp[9]) ? 4'b1001 : 4'b1101;
																assign node2037 = (inp[9]) ? 4'b1101 : 4'b1001;
											assign node2040 = (inp[4]) ? node2090 : node2041;
												assign node2041 = (inp[3]) ? node2069 : node2042;
													assign node2042 = (inp[12]) ? node2058 : node2043;
														assign node2043 = (inp[9]) ? node2051 : node2044;
															assign node2044 = (inp[0]) ? node2048 : node2045;
																assign node2045 = (inp[15]) ? 4'b1101 : 4'b1111;
																assign node2048 = (inp[15]) ? 4'b1111 : 4'b1101;
															assign node2051 = (inp[0]) ? node2055 : node2052;
																assign node2052 = (inp[15]) ? 4'b1001 : 4'b1011;
																assign node2055 = (inp[15]) ? 4'b1011 : 4'b1001;
														assign node2058 = (inp[9]) ? node2064 : node2059;
															assign node2059 = (inp[15]) ? node2061 : 4'b1001;
																assign node2061 = (inp[0]) ? 4'b1011 : 4'b1001;
															assign node2064 = (inp[15]) ? node2066 : 4'b1101;
																assign node2066 = (inp[0]) ? 4'b1101 : 4'b1111;
													assign node2069 = (inp[15]) ? node2081 : node2070;
														assign node2070 = (inp[0]) ? node2076 : node2071;
															assign node2071 = (inp[9]) ? 4'b1001 : node2072;
																assign node2072 = (inp[12]) ? 4'b1001 : 4'b1101;
															assign node2076 = (inp[12]) ? node2078 : 4'b1011;
																assign node2078 = (inp[9]) ? 4'b1111 : 4'b1011;
														assign node2081 = (inp[0]) ? node2083 : 4'b1011;
															assign node2083 = (inp[9]) ? node2087 : node2084;
																assign node2084 = (inp[12]) ? 4'b1001 : 4'b1101;
																assign node2087 = (inp[12]) ? 4'b1101 : 4'b1001;
												assign node2090 = (inp[0]) ? node2106 : node2091;
													assign node2091 = (inp[15]) ? node2097 : node2092;
														assign node2092 = (inp[9]) ? 4'b1101 : node2093;
															assign node2093 = (inp[3]) ? 4'b1001 : 4'b1011;
														assign node2097 = (inp[12]) ? node2103 : node2098;
															assign node2098 = (inp[9]) ? 4'b1111 : node2099;
																assign node2099 = (inp[3]) ? 4'b1011 : 4'b1001;
															assign node2103 = (inp[9]) ? 4'b1011 : 4'b1111;
													assign node2106 = (inp[15]) ? node2114 : node2107;
														assign node2107 = (inp[12]) ? node2111 : node2108;
															assign node2108 = (inp[3]) ? 4'b1011 : 4'b1111;
															assign node2111 = (inp[9]) ? 4'b1011 : 4'b1111;
														assign node2114 = (inp[12]) ? node2116 : 4'b1011;
															assign node2116 = (inp[9]) ? 4'b1001 : 4'b1101;
									assign node2119 = (inp[12]) ? node2235 : node2120;
										assign node2120 = (inp[9]) ? node2162 : node2121;
											assign node2121 = (inp[4]) ? node2143 : node2122;
												assign node2122 = (inp[15]) ? node2134 : node2123;
													assign node2123 = (inp[0]) ? node2129 : node2124;
														assign node2124 = (inp[3]) ? node2126 : 4'b1110;
															assign node2126 = (inp[5]) ? 4'b1100 : 4'b1110;
														assign node2129 = (inp[3]) ? node2131 : 4'b1100;
															assign node2131 = (inp[5]) ? 4'b1110 : 4'b1100;
													assign node2134 = (inp[0]) ? node2140 : node2135;
														assign node2135 = (inp[3]) ? node2137 : 4'b1100;
															assign node2137 = (inp[5]) ? 4'b1110 : 4'b1100;
														assign node2140 = (inp[5]) ? 4'b1100 : 4'b1110;
												assign node2143 = (inp[3]) ? node2151 : node2144;
													assign node2144 = (inp[0]) ? node2148 : node2145;
														assign node2145 = (inp[15]) ? 4'b1000 : 4'b1010;
														assign node2148 = (inp[15]) ? 4'b1010 : 4'b1000;
													assign node2151 = (inp[5]) ? node2157 : node2152;
														assign node2152 = (inp[0]) ? 4'b1000 : node2153;
															assign node2153 = (inp[15]) ? 4'b1000 : 4'b1010;
														assign node2157 = (inp[0]) ? 4'b1010 : node2158;
															assign node2158 = (inp[15]) ? 4'b1010 : 4'b1000;
											assign node2162 = (inp[4]) ? node2196 : node2163;
												assign node2163 = (inp[5]) ? node2177 : node2164;
													assign node2164 = (inp[10]) ? node2170 : node2165;
														assign node2165 = (inp[15]) ? 4'b1000 : node2166;
															assign node2166 = (inp[0]) ? 4'b1000 : 4'b1010;
														assign node2170 = (inp[15]) ? node2174 : node2171;
															assign node2171 = (inp[0]) ? 4'b1000 : 4'b1010;
															assign node2174 = (inp[0]) ? 4'b1010 : 4'b1000;
													assign node2177 = (inp[0]) ? node2183 : node2178;
														assign node2178 = (inp[15]) ? 4'b1010 : node2179;
															assign node2179 = (inp[3]) ? 4'b1000 : 4'b1010;
														assign node2183 = (inp[10]) ? node2191 : node2184;
															assign node2184 = (inp[15]) ? node2188 : node2185;
																assign node2185 = (inp[3]) ? 4'b1010 : 4'b1000;
																assign node2188 = (inp[3]) ? 4'b1000 : 4'b1010;
															assign node2191 = (inp[3]) ? node2193 : 4'b1000;
																assign node2193 = (inp[15]) ? 4'b1000 : 4'b1010;
												assign node2196 = (inp[3]) ? node2214 : node2197;
													assign node2197 = (inp[5]) ? node2207 : node2198;
														assign node2198 = (inp[10]) ? node2202 : node2199;
															assign node2199 = (inp[0]) ? 4'b1110 : 4'b1100;
															assign node2202 = (inp[0]) ? 4'b1100 : node2203;
																assign node2203 = (inp[15]) ? 4'b1100 : 4'b1110;
														assign node2207 = (inp[0]) ? node2211 : node2208;
															assign node2208 = (inp[15]) ? 4'b1110 : 4'b1100;
															assign node2211 = (inp[15]) ? 4'b1100 : 4'b1110;
													assign node2214 = (inp[5]) ? node2230 : node2215;
														assign node2215 = (inp[10]) ? node2223 : node2216;
															assign node2216 = (inp[15]) ? node2220 : node2217;
																assign node2217 = (inp[0]) ? 4'b1110 : 4'b1100;
																assign node2220 = (inp[0]) ? 4'b1100 : 4'b1110;
															assign node2223 = (inp[15]) ? node2227 : node2224;
																assign node2224 = (inp[0]) ? 4'b1110 : 4'b1100;
																assign node2227 = (inp[0]) ? 4'b1100 : 4'b1110;
														assign node2230 = (inp[0]) ? node2232 : 4'b1100;
															assign node2232 = (inp[15]) ? 4'b1100 : 4'b1110;
										assign node2235 = (inp[0]) ? node2335 : node2236;
											assign node2236 = (inp[5]) ? node2294 : node2237;
												assign node2237 = (inp[15]) ? node2267 : node2238;
													assign node2238 = (inp[3]) ? node2254 : node2239;
														assign node2239 = (inp[9]) ? node2247 : node2240;
															assign node2240 = (inp[10]) ? node2244 : node2241;
																assign node2241 = (inp[4]) ? 4'b1010 : 4'b1110;
																assign node2244 = (inp[4]) ? 4'b1110 : 4'b1010;
															assign node2247 = (inp[10]) ? node2251 : node2248;
																assign node2248 = (inp[4]) ? 4'b1110 : 4'b1010;
																assign node2251 = (inp[4]) ? 4'b1010 : 4'b1110;
														assign node2254 = (inp[10]) ? node2260 : node2255;
															assign node2255 = (inp[9]) ? 4'b1010 : node2256;
																assign node2256 = (inp[4]) ? 4'b1010 : 4'b1110;
															assign node2260 = (inp[4]) ? node2264 : node2261;
																assign node2261 = (inp[9]) ? 4'b1100 : 4'b1010;
																assign node2264 = (inp[9]) ? 4'b1000 : 4'b1100;
													assign node2267 = (inp[3]) ? node2281 : node2268;
														assign node2268 = (inp[4]) ? node2276 : node2269;
															assign node2269 = (inp[10]) ? node2273 : node2270;
																assign node2270 = (inp[9]) ? 4'b1000 : 4'b1100;
																assign node2273 = (inp[9]) ? 4'b1100 : 4'b1000;
															assign node2276 = (inp[9]) ? node2278 : 4'b1100;
																assign node2278 = (inp[10]) ? 4'b1000 : 4'b1100;
														assign node2281 = (inp[10]) ? node2287 : node2282;
															assign node2282 = (inp[9]) ? node2284 : 4'b1000;
																assign node2284 = (inp[4]) ? 4'b1110 : 4'b1000;
															assign node2287 = (inp[4]) ? node2291 : node2288;
																assign node2288 = (inp[9]) ? 4'b1110 : 4'b1000;
																assign node2291 = (inp[9]) ? 4'b1010 : 4'b1110;
												assign node2294 = (inp[15]) ? node2312 : node2295;
													assign node2295 = (inp[3]) ? node2307 : node2296;
														assign node2296 = (inp[10]) ? node2302 : node2297;
															assign node2297 = (inp[9]) ? 4'b1010 : node2298;
																assign node2298 = (inp[4]) ? 4'b1010 : 4'b1110;
															assign node2302 = (inp[4]) ? 4'b1100 : node2303;
																assign node2303 = (inp[9]) ? 4'b1100 : 4'b1010;
														assign node2307 = (inp[4]) ? 4'b1100 : node2308;
															assign node2308 = (inp[9]) ? 4'b1100 : 4'b1000;
													assign node2312 = (inp[9]) ? node2324 : node2313;
														assign node2313 = (inp[3]) ? node2319 : node2314;
															assign node2314 = (inp[10]) ? 4'b1110 : node2315;
																assign node2315 = (inp[4]) ? 4'b1000 : 4'b1100;
															assign node2319 = (inp[4]) ? 4'b1110 : node2320;
																assign node2320 = (inp[10]) ? 4'b1010 : 4'b1110;
														assign node2324 = (inp[3]) ? node2330 : node2325;
															assign node2325 = (inp[4]) ? node2327 : 4'b1110;
																assign node2327 = (inp[10]) ? 4'b1010 : 4'b1110;
															assign node2330 = (inp[10]) ? 4'b1110 : node2331;
																assign node2331 = (inp[4]) ? 4'b1110 : 4'b1010;
											assign node2335 = (inp[15]) ? node2387 : node2336;
												assign node2336 = (inp[5]) ? node2364 : node2337;
													assign node2337 = (inp[3]) ? node2349 : node2338;
														assign node2338 = (inp[4]) ? node2344 : node2339;
															assign node2339 = (inp[9]) ? node2341 : 4'b1100;
																assign node2341 = (inp[10]) ? 4'b1100 : 4'b1000;
															assign node2344 = (inp[10]) ? 4'b1000 : node2345;
																assign node2345 = (inp[9]) ? 4'b1100 : 4'b1000;
														assign node2349 = (inp[4]) ? node2357 : node2350;
															assign node2350 = (inp[10]) ? node2354 : node2351;
																assign node2351 = (inp[9]) ? 4'b1000 : 4'b1100;
																assign node2354 = (inp[9]) ? 4'b1110 : 4'b1000;
															assign node2357 = (inp[10]) ? node2361 : node2358;
																assign node2358 = (inp[9]) ? 4'b1110 : 4'b1000;
																assign node2361 = (inp[9]) ? 4'b1010 : 4'b1110;
													assign node2364 = (inp[3]) ? node2378 : node2365;
														assign node2365 = (inp[4]) ? node2371 : node2366;
															assign node2366 = (inp[9]) ? node2368 : 4'b1000;
																assign node2368 = (inp[10]) ? 4'b1110 : 4'b1000;
															assign node2371 = (inp[9]) ? node2375 : node2372;
																assign node2372 = (inp[10]) ? 4'b1110 : 4'b1000;
																assign node2375 = (inp[10]) ? 4'b1010 : 4'b1110;
														assign node2378 = (inp[10]) ? 4'b1010 : node2379;
															assign node2379 = (inp[9]) ? node2383 : node2380;
																assign node2380 = (inp[4]) ? 4'b1010 : 4'b1110;
																assign node2383 = (inp[4]) ? 4'b1110 : 4'b1010;
												assign node2387 = (inp[3]) ? node2403 : node2388;
													assign node2388 = (inp[5]) ? node2400 : node2389;
														assign node2389 = (inp[9]) ? node2395 : node2390;
															assign node2390 = (inp[10]) ? 4'b1010 : node2391;
																assign node2391 = (inp[4]) ? 4'b1010 : 4'b1110;
															assign node2395 = (inp[10]) ? 4'b1110 : node2396;
																assign node2396 = (inp[4]) ? 4'b1110 : 4'b1010;
														assign node2400 = (inp[10]) ? 4'b1100 : 4'b1110;
													assign node2403 = (inp[5]) ? node2417 : node2404;
														assign node2404 = (inp[9]) ? node2412 : node2405;
															assign node2405 = (inp[10]) ? node2409 : node2406;
																assign node2406 = (inp[4]) ? 4'b1010 : 4'b1110;
																assign node2409 = (inp[4]) ? 4'b1100 : 4'b1010;
															assign node2412 = (inp[4]) ? node2414 : 4'b1100;
																assign node2414 = (inp[10]) ? 4'b1000 : 4'b1100;
														assign node2417 = (inp[10]) ? node2423 : node2418;
															assign node2418 = (inp[4]) ? node2420 : 4'b1000;
																assign node2420 = (inp[9]) ? 4'b1100 : 4'b1000;
															assign node2423 = (inp[9]) ? node2427 : node2424;
																assign node2424 = (inp[4]) ? 4'b1100 : 4'b1000;
																assign node2427 = (inp[4]) ? 4'b1000 : 4'b1100;
						assign node2430 = (inp[3]) ? node3490 : node2431;
							assign node2431 = (inp[4]) ? node2921 : node2432;
								assign node2432 = (inp[9]) ? node2686 : node2433;
									assign node2433 = (inp[12]) ? node2573 : node2434;
										assign node2434 = (inp[14]) ? node2522 : node2435;
											assign node2435 = (inp[5]) ? node2485 : node2436;
												assign node2436 = (inp[10]) ? node2464 : node2437;
													assign node2437 = (inp[15]) ? node2449 : node2438;
														assign node2438 = (inp[0]) ? node2444 : node2439;
															assign node2439 = (inp[7]) ? 4'b1111 : node2440;
																assign node2440 = (inp[8]) ? 4'b1111 : 4'b1110;
															assign node2444 = (inp[8]) ? 4'b1101 : node2445;
																assign node2445 = (inp[7]) ? 4'b1101 : 4'b1100;
														assign node2449 = (inp[0]) ? node2457 : node2450;
															assign node2450 = (inp[7]) ? node2454 : node2451;
																assign node2451 = (inp[8]) ? 4'b1101 : 4'b1100;
																assign node2454 = (inp[8]) ? 4'b1100 : 4'b1101;
															assign node2457 = (inp[7]) ? node2461 : node2458;
																assign node2458 = (inp[8]) ? 4'b1111 : 4'b1110;
																assign node2461 = (inp[8]) ? 4'b1110 : 4'b1111;
													assign node2464 = (inp[15]) ? node2476 : node2465;
														assign node2465 = (inp[0]) ? node2471 : node2466;
															assign node2466 = (inp[7]) ? node2468 : 4'b1110;
																assign node2468 = (inp[8]) ? 4'b1110 : 4'b1111;
															assign node2471 = (inp[8]) ? node2473 : 4'b1100;
																assign node2473 = (inp[7]) ? 4'b1100 : 4'b1101;
														assign node2476 = (inp[0]) ? 4'b1111 : node2477;
															assign node2477 = (inp[8]) ? node2481 : node2478;
																assign node2478 = (inp[7]) ? 4'b1101 : 4'b1100;
																assign node2481 = (inp[7]) ? 4'b1100 : 4'b1101;
												assign node2485 = (inp[7]) ? node2509 : node2486;
													assign node2486 = (inp[8]) ? node2494 : node2487;
														assign node2487 = (inp[10]) ? node2489 : 4'b1110;
															assign node2489 = (inp[0]) ? 4'b1100 : node2490;
																assign node2490 = (inp[15]) ? 4'b1100 : 4'b1110;
														assign node2494 = (inp[10]) ? node2502 : node2495;
															assign node2495 = (inp[0]) ? node2499 : node2496;
																assign node2496 = (inp[15]) ? 4'b1101 : 4'b1111;
																assign node2499 = (inp[15]) ? 4'b1111 : 4'b1101;
															assign node2502 = (inp[0]) ? node2506 : node2503;
																assign node2503 = (inp[15]) ? 4'b1101 : 4'b1111;
																assign node2506 = (inp[15]) ? 4'b1111 : 4'b1101;
													assign node2509 = (inp[8]) ? node2517 : node2510;
														assign node2510 = (inp[10]) ? node2512 : 4'b1101;
															assign node2512 = (inp[0]) ? 4'b1111 : node2513;
																assign node2513 = (inp[15]) ? 4'b1101 : 4'b1111;
														assign node2517 = (inp[15]) ? 4'b1110 : node2518;
															assign node2518 = (inp[0]) ? 4'b1100 : 4'b1110;
											assign node2522 = (inp[8]) ? node2548 : node2523;
												assign node2523 = (inp[7]) ? node2531 : node2524;
													assign node2524 = (inp[0]) ? node2528 : node2525;
														assign node2525 = (inp[15]) ? 4'b1100 : 4'b1110;
														assign node2528 = (inp[15]) ? 4'b1110 : 4'b1100;
													assign node2531 = (inp[5]) ? node2539 : node2532;
														assign node2532 = (inp[15]) ? node2536 : node2533;
															assign node2533 = (inp[0]) ? 4'b1101 : 4'b1111;
															assign node2536 = (inp[0]) ? 4'b1111 : 4'b1101;
														assign node2539 = (inp[10]) ? node2541 : 4'b1111;
															assign node2541 = (inp[0]) ? node2545 : node2542;
																assign node2542 = (inp[15]) ? 4'b1101 : 4'b1111;
																assign node2545 = (inp[15]) ? 4'b1111 : 4'b1101;
												assign node2548 = (inp[7]) ? node2556 : node2549;
													assign node2549 = (inp[10]) ? node2551 : 4'b1111;
														assign node2551 = (inp[0]) ? 4'b1101 : node2552;
															assign node2552 = (inp[15]) ? 4'b1101 : 4'b1111;
													assign node2556 = (inp[10]) ? node2566 : node2557;
														assign node2557 = (inp[5]) ? node2559 : 4'b1100;
															assign node2559 = (inp[15]) ? node2563 : node2560;
																assign node2560 = (inp[0]) ? 4'b1100 : 4'b1110;
																assign node2563 = (inp[0]) ? 4'b1110 : 4'b1100;
														assign node2566 = (inp[15]) ? node2570 : node2567;
															assign node2567 = (inp[0]) ? 4'b1100 : 4'b1110;
															assign node2570 = (inp[0]) ? 4'b1110 : 4'b1100;
										assign node2573 = (inp[10]) ? node2639 : node2574;
											assign node2574 = (inp[5]) ? node2610 : node2575;
												assign node2575 = (inp[7]) ? node2591 : node2576;
													assign node2576 = (inp[8]) ? node2584 : node2577;
														assign node2577 = (inp[0]) ? node2581 : node2578;
															assign node2578 = (inp[15]) ? 4'b1100 : 4'b1110;
															assign node2581 = (inp[15]) ? 4'b1110 : 4'b1100;
														assign node2584 = (inp[15]) ? node2588 : node2585;
															assign node2585 = (inp[0]) ? 4'b1101 : 4'b1111;
															assign node2588 = (inp[0]) ? 4'b1111 : 4'b1101;
													assign node2591 = (inp[8]) ? node2599 : node2592;
														assign node2592 = (inp[15]) ? node2596 : node2593;
															assign node2593 = (inp[0]) ? 4'b1101 : 4'b1111;
															assign node2596 = (inp[0]) ? 4'b1111 : 4'b1101;
														assign node2599 = (inp[14]) ? node2605 : node2600;
															assign node2600 = (inp[15]) ? node2602 : 4'b1100;
																assign node2602 = (inp[0]) ? 4'b1110 : 4'b1100;
															assign node2605 = (inp[0]) ? 4'b1110 : node2606;
																assign node2606 = (inp[15]) ? 4'b1100 : 4'b1110;
												assign node2610 = (inp[15]) ? node2624 : node2611;
													assign node2611 = (inp[0]) ? node2619 : node2612;
														assign node2612 = (inp[7]) ? node2616 : node2613;
															assign node2613 = (inp[8]) ? 4'b1111 : 4'b1110;
															assign node2616 = (inp[8]) ? 4'b1110 : 4'b1111;
														assign node2619 = (inp[7]) ? node2621 : 4'b1101;
															assign node2621 = (inp[8]) ? 4'b1100 : 4'b1101;
													assign node2624 = (inp[0]) ? node2632 : node2625;
														assign node2625 = (inp[8]) ? node2629 : node2626;
															assign node2626 = (inp[7]) ? 4'b1101 : 4'b1100;
															assign node2629 = (inp[7]) ? 4'b1100 : 4'b1101;
														assign node2632 = (inp[14]) ? 4'b1111 : node2633;
															assign node2633 = (inp[8]) ? 4'b1111 : node2634;
																assign node2634 = (inp[7]) ? 4'b1111 : 4'b1110;
											assign node2639 = (inp[8]) ? node2663 : node2640;
												assign node2640 = (inp[7]) ? node2648 : node2641;
													assign node2641 = (inp[0]) ? node2645 : node2642;
														assign node2642 = (inp[15]) ? 4'b1000 : 4'b1010;
														assign node2645 = (inp[15]) ? 4'b1010 : 4'b1000;
													assign node2648 = (inp[14]) ? node2656 : node2649;
														assign node2649 = (inp[0]) ? node2653 : node2650;
															assign node2650 = (inp[15]) ? 4'b1001 : 4'b1011;
															assign node2653 = (inp[15]) ? 4'b1011 : 4'b1001;
														assign node2656 = (inp[15]) ? node2660 : node2657;
															assign node2657 = (inp[0]) ? 4'b1001 : 4'b1011;
															assign node2660 = (inp[0]) ? 4'b1011 : 4'b1001;
												assign node2663 = (inp[7]) ? node2679 : node2664;
													assign node2664 = (inp[14]) ? node2672 : node2665;
														assign node2665 = (inp[15]) ? node2669 : node2666;
															assign node2666 = (inp[0]) ? 4'b1001 : 4'b1011;
															assign node2669 = (inp[0]) ? 4'b1011 : 4'b1001;
														assign node2672 = (inp[15]) ? node2676 : node2673;
															assign node2673 = (inp[0]) ? 4'b1001 : 4'b1011;
															assign node2676 = (inp[0]) ? 4'b1011 : 4'b1001;
													assign node2679 = (inp[0]) ? node2683 : node2680;
														assign node2680 = (inp[15]) ? 4'b1000 : 4'b1010;
														assign node2683 = (inp[15]) ? 4'b1010 : 4'b1000;
									assign node2686 = (inp[12]) ? node2788 : node2687;
										assign node2687 = (inp[7]) ? node2759 : node2688;
											assign node2688 = (inp[8]) ? node2718 : node2689;
												assign node2689 = (inp[10]) ? node2697 : node2690;
													assign node2690 = (inp[15]) ? node2694 : node2691;
														assign node2691 = (inp[0]) ? 4'b1000 : 4'b1010;
														assign node2694 = (inp[0]) ? 4'b1010 : 4'b1000;
													assign node2697 = (inp[14]) ? node2711 : node2698;
														assign node2698 = (inp[5]) ? node2706 : node2699;
															assign node2699 = (inp[0]) ? node2703 : node2700;
																assign node2700 = (inp[15]) ? 4'b1000 : 4'b1010;
																assign node2703 = (inp[15]) ? 4'b1010 : 4'b1000;
															assign node2706 = (inp[15]) ? 4'b1000 : node2707;
																assign node2707 = (inp[0]) ? 4'b1000 : 4'b1010;
														assign node2711 = (inp[0]) ? node2715 : node2712;
															assign node2712 = (inp[15]) ? 4'b1000 : 4'b1010;
															assign node2715 = (inp[15]) ? 4'b1010 : 4'b1000;
												assign node2718 = (inp[14]) ? node2740 : node2719;
													assign node2719 = (inp[10]) ? node2727 : node2720;
														assign node2720 = (inp[5]) ? 4'b1001 : node2721;
															assign node2721 = (inp[15]) ? node2723 : 4'b1001;
																assign node2723 = (inp[0]) ? 4'b1011 : 4'b1001;
														assign node2727 = (inp[5]) ? node2733 : node2728;
															assign node2728 = (inp[0]) ? 4'b1001 : node2729;
																assign node2729 = (inp[15]) ? 4'b1001 : 4'b1011;
															assign node2733 = (inp[15]) ? node2737 : node2734;
																assign node2734 = (inp[0]) ? 4'b1001 : 4'b1011;
																assign node2737 = (inp[0]) ? 4'b1011 : 4'b1001;
													assign node2740 = (inp[10]) ? node2752 : node2741;
														assign node2741 = (inp[5]) ? node2747 : node2742;
															assign node2742 = (inp[15]) ? node2744 : 4'b1001;
																assign node2744 = (inp[0]) ? 4'b1011 : 4'b1001;
															assign node2747 = (inp[15]) ? node2749 : 4'b1011;
																assign node2749 = (inp[0]) ? 4'b1011 : 4'b1001;
														assign node2752 = (inp[15]) ? node2756 : node2753;
															assign node2753 = (inp[0]) ? 4'b1001 : 4'b1011;
															assign node2756 = (inp[0]) ? 4'b1011 : 4'b1001;
											assign node2759 = (inp[8]) ? node2767 : node2760;
												assign node2760 = (inp[0]) ? node2764 : node2761;
													assign node2761 = (inp[15]) ? 4'b1001 : 4'b1011;
													assign node2764 = (inp[15]) ? 4'b1011 : 4'b1001;
												assign node2767 = (inp[10]) ? node2781 : node2768;
													assign node2768 = (inp[5]) ? node2774 : node2769;
														assign node2769 = (inp[15]) ? 4'b1000 : node2770;
															assign node2770 = (inp[0]) ? 4'b1000 : 4'b1010;
														assign node2774 = (inp[15]) ? node2778 : node2775;
															assign node2775 = (inp[0]) ? 4'b1000 : 4'b1010;
															assign node2778 = (inp[0]) ? 4'b1010 : 4'b1000;
													assign node2781 = (inp[15]) ? node2785 : node2782;
														assign node2782 = (inp[0]) ? 4'b1000 : 4'b1010;
														assign node2785 = (inp[0]) ? 4'b1010 : 4'b1000;
										assign node2788 = (inp[10]) ? node2856 : node2789;
											assign node2789 = (inp[14]) ? node2825 : node2790;
												assign node2790 = (inp[15]) ? node2812 : node2791;
													assign node2791 = (inp[0]) ? node2805 : node2792;
														assign node2792 = (inp[5]) ? node2798 : node2793;
															assign node2793 = (inp[7]) ? 4'b1011 : node2794;
																assign node2794 = (inp[8]) ? 4'b1011 : 4'b1010;
															assign node2798 = (inp[8]) ? node2802 : node2799;
																assign node2799 = (inp[7]) ? 4'b1011 : 4'b1010;
																assign node2802 = (inp[7]) ? 4'b1010 : 4'b1011;
														assign node2805 = (inp[8]) ? node2809 : node2806;
															assign node2806 = (inp[7]) ? 4'b1001 : 4'b1000;
															assign node2809 = (inp[7]) ? 4'b1000 : 4'b1001;
													assign node2812 = (inp[0]) ? node2820 : node2813;
														assign node2813 = (inp[7]) ? node2817 : node2814;
															assign node2814 = (inp[8]) ? 4'b1001 : 4'b1000;
															assign node2817 = (inp[8]) ? 4'b1000 : 4'b1001;
														assign node2820 = (inp[8]) ? node2822 : 4'b1011;
															assign node2822 = (inp[7]) ? 4'b1010 : 4'b1011;
												assign node2825 = (inp[8]) ? node2841 : node2826;
													assign node2826 = (inp[7]) ? node2834 : node2827;
														assign node2827 = (inp[15]) ? node2831 : node2828;
															assign node2828 = (inp[0]) ? 4'b1000 : 4'b1010;
															assign node2831 = (inp[0]) ? 4'b1010 : 4'b1000;
														assign node2834 = (inp[0]) ? node2838 : node2835;
															assign node2835 = (inp[15]) ? 4'b1001 : 4'b1011;
															assign node2838 = (inp[5]) ? 4'b1001 : 4'b1011;
													assign node2841 = (inp[7]) ? node2851 : node2842;
														assign node2842 = (inp[5]) ? node2844 : 4'b1011;
															assign node2844 = (inp[15]) ? node2848 : node2845;
																assign node2845 = (inp[0]) ? 4'b1001 : 4'b1011;
																assign node2848 = (inp[0]) ? 4'b1011 : 4'b1001;
														assign node2851 = (inp[5]) ? node2853 : 4'b1010;
															assign node2853 = (inp[15]) ? 4'b1010 : 4'b1000;
											assign node2856 = (inp[8]) ? node2892 : node2857;
												assign node2857 = (inp[7]) ? node2879 : node2858;
													assign node2858 = (inp[0]) ? node2872 : node2859;
														assign node2859 = (inp[14]) ? node2867 : node2860;
															assign node2860 = (inp[15]) ? node2864 : node2861;
																assign node2861 = (inp[5]) ? 4'b1100 : 4'b1110;
																assign node2864 = (inp[5]) ? 4'b1110 : 4'b1100;
															assign node2867 = (inp[5]) ? node2869 : 4'b1110;
																assign node2869 = (inp[15]) ? 4'b1110 : 4'b1100;
														assign node2872 = (inp[15]) ? node2876 : node2873;
															assign node2873 = (inp[5]) ? 4'b1110 : 4'b1100;
															assign node2876 = (inp[5]) ? 4'b1100 : 4'b1110;
													assign node2879 = (inp[0]) ? node2887 : node2880;
														assign node2880 = (inp[14]) ? node2882 : 4'b1101;
															assign node2882 = (inp[15]) ? node2884 : 4'b1101;
																assign node2884 = (inp[5]) ? 4'b1111 : 4'b1101;
														assign node2887 = (inp[15]) ? node2889 : 4'b1111;
															assign node2889 = (inp[5]) ? 4'b1101 : 4'b1111;
												assign node2892 = (inp[7]) ? node2908 : node2893;
													assign node2893 = (inp[5]) ? node2901 : node2894;
														assign node2894 = (inp[15]) ? node2898 : node2895;
															assign node2895 = (inp[0]) ? 4'b1101 : 4'b1111;
															assign node2898 = (inp[0]) ? 4'b1111 : 4'b1101;
														assign node2901 = (inp[0]) ? node2905 : node2902;
															assign node2902 = (inp[15]) ? 4'b1111 : 4'b1101;
															assign node2905 = (inp[15]) ? 4'b1101 : 4'b1111;
													assign node2908 = (inp[0]) ? node2914 : node2909;
														assign node2909 = (inp[5]) ? node2911 : 4'b1110;
															assign node2911 = (inp[14]) ? 4'b1110 : 4'b1100;
														assign node2914 = (inp[15]) ? node2918 : node2915;
															assign node2915 = (inp[5]) ? 4'b1110 : 4'b1100;
															assign node2918 = (inp[5]) ? 4'b1100 : 4'b1110;
								assign node2921 = (inp[9]) ? node3207 : node2922;
									assign node2922 = (inp[10]) ? node3064 : node2923;
										assign node2923 = (inp[5]) ? node2999 : node2924;
											assign node2924 = (inp[12]) ? node2958 : node2925;
												assign node2925 = (inp[7]) ? node2943 : node2926;
													assign node2926 = (inp[8]) ? node2934 : node2927;
														assign node2927 = (inp[15]) ? node2931 : node2928;
															assign node2928 = (inp[0]) ? 4'b1000 : 4'b1010;
															assign node2931 = (inp[0]) ? 4'b1010 : 4'b1000;
														assign node2934 = (inp[14]) ? node2936 : 4'b1001;
															assign node2936 = (inp[0]) ? node2940 : node2937;
																assign node2937 = (inp[15]) ? 4'b1001 : 4'b1011;
																assign node2940 = (inp[15]) ? 4'b1011 : 4'b1001;
													assign node2943 = (inp[8]) ? node2951 : node2944;
														assign node2944 = (inp[0]) ? node2948 : node2945;
															assign node2945 = (inp[15]) ? 4'b1001 : 4'b1011;
															assign node2948 = (inp[15]) ? 4'b1011 : 4'b1001;
														assign node2951 = (inp[14]) ? 4'b1010 : node2952;
															assign node2952 = (inp[0]) ? node2954 : 4'b1010;
																assign node2954 = (inp[15]) ? 4'b1010 : 4'b1000;
												assign node2958 = (inp[0]) ? node2978 : node2959;
													assign node2959 = (inp[15]) ? node2967 : node2960;
														assign node2960 = (inp[7]) ? node2964 : node2961;
															assign node2961 = (inp[8]) ? 4'b1011 : 4'b1010;
															assign node2964 = (inp[8]) ? 4'b1010 : 4'b1011;
														assign node2967 = (inp[14]) ? node2973 : node2968;
															assign node2968 = (inp[7]) ? node2970 : 4'b1001;
																assign node2970 = (inp[8]) ? 4'b1000 : 4'b1001;
															assign node2973 = (inp[8]) ? node2975 : 4'b1000;
																assign node2975 = (inp[7]) ? 4'b1000 : 4'b1001;
													assign node2978 = (inp[15]) ? node2986 : node2979;
														assign node2979 = (inp[8]) ? node2983 : node2980;
															assign node2980 = (inp[7]) ? 4'b1001 : 4'b1000;
															assign node2983 = (inp[7]) ? 4'b1000 : 4'b1001;
														assign node2986 = (inp[14]) ? node2994 : node2987;
															assign node2987 = (inp[7]) ? node2991 : node2988;
																assign node2988 = (inp[8]) ? 4'b1011 : 4'b1010;
																assign node2991 = (inp[8]) ? 4'b1010 : 4'b1011;
															assign node2994 = (inp[7]) ? 4'b1010 : node2995;
																assign node2995 = (inp[8]) ? 4'b1011 : 4'b1010;
											assign node2999 = (inp[7]) ? node3039 : node3000;
												assign node3000 = (inp[8]) ? node3016 : node3001;
													assign node3001 = (inp[12]) ? node3009 : node3002;
														assign node3002 = (inp[0]) ? node3006 : node3003;
															assign node3003 = (inp[15]) ? 4'b1000 : 4'b1010;
															assign node3006 = (inp[15]) ? 4'b1010 : 4'b1000;
														assign node3009 = (inp[15]) ? node3013 : node3010;
															assign node3010 = (inp[0]) ? 4'b1000 : 4'b1010;
															assign node3013 = (inp[14]) ? 4'b1000 : 4'b1010;
													assign node3016 = (inp[12]) ? node3024 : node3017;
														assign node3017 = (inp[15]) ? node3021 : node3018;
															assign node3018 = (inp[0]) ? 4'b1001 : 4'b1011;
															assign node3021 = (inp[0]) ? 4'b1011 : 4'b1001;
														assign node3024 = (inp[14]) ? node3032 : node3025;
															assign node3025 = (inp[15]) ? node3029 : node3026;
																assign node3026 = (inp[0]) ? 4'b1001 : 4'b1011;
																assign node3029 = (inp[0]) ? 4'b1011 : 4'b1001;
															assign node3032 = (inp[15]) ? node3036 : node3033;
																assign node3033 = (inp[0]) ? 4'b1001 : 4'b1011;
																assign node3036 = (inp[0]) ? 4'b1011 : 4'b1001;
												assign node3039 = (inp[8]) ? node3053 : node3040;
													assign node3040 = (inp[12]) ? node3048 : node3041;
														assign node3041 = (inp[0]) ? node3045 : node3042;
															assign node3042 = (inp[15]) ? 4'b1001 : 4'b1011;
															assign node3045 = (inp[15]) ? 4'b1011 : 4'b1001;
														assign node3048 = (inp[0]) ? 4'b1001 : node3049;
															assign node3049 = (inp[15]) ? 4'b1001 : 4'b1011;
													assign node3053 = (inp[14]) ? node3055 : 4'b1000;
														assign node3055 = (inp[12]) ? node3057 : 4'b1000;
															assign node3057 = (inp[15]) ? node3061 : node3058;
																assign node3058 = (inp[0]) ? 4'b1000 : 4'b1010;
																assign node3061 = (inp[0]) ? 4'b1010 : 4'b1000;
										assign node3064 = (inp[12]) ? node3132 : node3065;
											assign node3065 = (inp[0]) ? node3099 : node3066;
												assign node3066 = (inp[15]) ? node3074 : node3067;
													assign node3067 = (inp[7]) ? node3071 : node3068;
														assign node3068 = (inp[8]) ? 4'b1011 : 4'b1010;
														assign node3071 = (inp[8]) ? 4'b1010 : 4'b1011;
													assign node3074 = (inp[14]) ? node3090 : node3075;
														assign node3075 = (inp[5]) ? node3083 : node3076;
															assign node3076 = (inp[8]) ? node3080 : node3077;
																assign node3077 = (inp[7]) ? 4'b1001 : 4'b1000;
																assign node3080 = (inp[7]) ? 4'b1000 : 4'b1001;
															assign node3083 = (inp[8]) ? node3087 : node3084;
																assign node3084 = (inp[7]) ? 4'b1001 : 4'b1000;
																assign node3087 = (inp[7]) ? 4'b1000 : 4'b1001;
														assign node3090 = (inp[5]) ? 4'b1000 : node3091;
															assign node3091 = (inp[7]) ? node3095 : node3092;
																assign node3092 = (inp[8]) ? 4'b1001 : 4'b1000;
																assign node3095 = (inp[8]) ? 4'b1000 : 4'b1001;
												assign node3099 = (inp[15]) ? node3117 : node3100;
													assign node3100 = (inp[14]) ? node3106 : node3101;
														assign node3101 = (inp[8]) ? 4'b1000 : node3102;
															assign node3102 = (inp[7]) ? 4'b1001 : 4'b1000;
														assign node3106 = (inp[5]) ? node3112 : node3107;
															assign node3107 = (inp[8]) ? node3109 : 4'b1000;
																assign node3109 = (inp[7]) ? 4'b1000 : 4'b1001;
															assign node3112 = (inp[8]) ? node3114 : 4'b1001;
																assign node3114 = (inp[7]) ? 4'b1000 : 4'b1001;
													assign node3117 = (inp[5]) ? node3125 : node3118;
														assign node3118 = (inp[7]) ? node3122 : node3119;
															assign node3119 = (inp[8]) ? 4'b1011 : 4'b1010;
															assign node3122 = (inp[8]) ? 4'b1010 : 4'b1011;
														assign node3125 = (inp[8]) ? node3129 : node3126;
															assign node3126 = (inp[7]) ? 4'b1011 : 4'b1010;
															assign node3129 = (inp[7]) ? 4'b1010 : 4'b1011;
											assign node3132 = (inp[8]) ? node3168 : node3133;
												assign node3133 = (inp[7]) ? node3153 : node3134;
													assign node3134 = (inp[15]) ? node3140 : node3135;
														assign node3135 = (inp[14]) ? 4'b1110 : node3136;
															assign node3136 = (inp[0]) ? 4'b1110 : 4'b1100;
														assign node3140 = (inp[14]) ? node3146 : node3141;
															assign node3141 = (inp[5]) ? node3143 : 4'b1110;
																assign node3143 = (inp[0]) ? 4'b1100 : 4'b1110;
															assign node3146 = (inp[0]) ? node3150 : node3147;
																assign node3147 = (inp[5]) ? 4'b1110 : 4'b1100;
																assign node3150 = (inp[5]) ? 4'b1100 : 4'b1110;
													assign node3153 = (inp[0]) ? node3161 : node3154;
														assign node3154 = (inp[15]) ? node3158 : node3155;
															assign node3155 = (inp[5]) ? 4'b1101 : 4'b1111;
															assign node3158 = (inp[5]) ? 4'b1111 : 4'b1101;
														assign node3161 = (inp[5]) ? node3165 : node3162;
															assign node3162 = (inp[15]) ? 4'b1111 : 4'b1101;
															assign node3165 = (inp[15]) ? 4'b1101 : 4'b1111;
												assign node3168 = (inp[7]) ? node3192 : node3169;
													assign node3169 = (inp[14]) ? node3183 : node3170;
														assign node3170 = (inp[0]) ? node3178 : node3171;
															assign node3171 = (inp[5]) ? node3175 : node3172;
																assign node3172 = (inp[15]) ? 4'b1101 : 4'b1111;
																assign node3175 = (inp[15]) ? 4'b1111 : 4'b1101;
															assign node3178 = (inp[5]) ? 4'b1101 : node3179;
																assign node3179 = (inp[15]) ? 4'b1111 : 4'b1101;
														assign node3183 = (inp[5]) ? node3185 : 4'b1101;
															assign node3185 = (inp[15]) ? node3189 : node3186;
																assign node3186 = (inp[0]) ? 4'b1111 : 4'b1101;
																assign node3189 = (inp[0]) ? 4'b1101 : 4'b1111;
													assign node3192 = (inp[5]) ? node3200 : node3193;
														assign node3193 = (inp[0]) ? node3197 : node3194;
															assign node3194 = (inp[15]) ? 4'b1100 : 4'b1110;
															assign node3197 = (inp[15]) ? 4'b1110 : 4'b1100;
														assign node3200 = (inp[0]) ? node3204 : node3201;
															assign node3201 = (inp[15]) ? 4'b1110 : 4'b1100;
															assign node3204 = (inp[15]) ? 4'b1100 : 4'b1110;
									assign node3207 = (inp[12]) ? node3315 : node3208;
										assign node3208 = (inp[8]) ? node3260 : node3209;
											assign node3209 = (inp[7]) ? node3237 : node3210;
												assign node3210 = (inp[14]) ? node3224 : node3211;
													assign node3211 = (inp[15]) ? node3219 : node3212;
														assign node3212 = (inp[0]) ? node3216 : node3213;
															assign node3213 = (inp[5]) ? 4'b1100 : 4'b1110;
															assign node3216 = (inp[5]) ? 4'b1110 : 4'b1100;
														assign node3219 = (inp[0]) ? 4'b1110 : node3220;
															assign node3220 = (inp[5]) ? 4'b1110 : 4'b1100;
													assign node3224 = (inp[0]) ? node3232 : node3225;
														assign node3225 = (inp[15]) ? node3229 : node3226;
															assign node3226 = (inp[5]) ? 4'b1100 : 4'b1110;
															assign node3229 = (inp[5]) ? 4'b1110 : 4'b1100;
														assign node3232 = (inp[5]) ? node3234 : 4'b1100;
															assign node3234 = (inp[15]) ? 4'b1100 : 4'b1110;
												assign node3237 = (inp[0]) ? node3245 : node3238;
													assign node3238 = (inp[15]) ? node3242 : node3239;
														assign node3239 = (inp[5]) ? 4'b1101 : 4'b1111;
														assign node3242 = (inp[5]) ? 4'b1111 : 4'b1101;
													assign node3245 = (inp[14]) ? 4'b1111 : node3246;
														assign node3246 = (inp[10]) ? node3252 : node3247;
															assign node3247 = (inp[15]) ? node3249 : 4'b1111;
																assign node3249 = (inp[5]) ? 4'b1101 : 4'b1111;
															assign node3252 = (inp[15]) ? node3256 : node3253;
																assign node3253 = (inp[5]) ? 4'b1111 : 4'b1101;
																assign node3256 = (inp[5]) ? 4'b1101 : 4'b1111;
											assign node3260 = (inp[7]) ? node3292 : node3261;
												assign node3261 = (inp[5]) ? node3275 : node3262;
													assign node3262 = (inp[14]) ? node3268 : node3263;
														assign node3263 = (inp[0]) ? node3265 : 4'b1111;
															assign node3265 = (inp[15]) ? 4'b1111 : 4'b1101;
														assign node3268 = (inp[0]) ? node3272 : node3269;
															assign node3269 = (inp[15]) ? 4'b1101 : 4'b1111;
															assign node3272 = (inp[15]) ? 4'b1111 : 4'b1101;
													assign node3275 = (inp[14]) ? node3285 : node3276;
														assign node3276 = (inp[10]) ? 4'b1101 : node3277;
															assign node3277 = (inp[15]) ? node3281 : node3278;
																assign node3278 = (inp[0]) ? 4'b1111 : 4'b1101;
																assign node3281 = (inp[0]) ? 4'b1101 : 4'b1111;
														assign node3285 = (inp[15]) ? node3289 : node3286;
															assign node3286 = (inp[0]) ? 4'b1111 : 4'b1101;
															assign node3289 = (inp[0]) ? 4'b1101 : 4'b1111;
												assign node3292 = (inp[0]) ? node3308 : node3293;
													assign node3293 = (inp[14]) ? node3301 : node3294;
														assign node3294 = (inp[5]) ? node3298 : node3295;
															assign node3295 = (inp[15]) ? 4'b1100 : 4'b1110;
															assign node3298 = (inp[15]) ? 4'b1110 : 4'b1100;
														assign node3301 = (inp[15]) ? node3305 : node3302;
															assign node3302 = (inp[5]) ? 4'b1100 : 4'b1110;
															assign node3305 = (inp[5]) ? 4'b1110 : 4'b1100;
													assign node3308 = (inp[15]) ? node3312 : node3309;
														assign node3309 = (inp[5]) ? 4'b1110 : 4'b1100;
														assign node3312 = (inp[5]) ? 4'b1100 : 4'b1110;
										assign node3315 = (inp[10]) ? node3401 : node3316;
											assign node3316 = (inp[14]) ? node3352 : node3317;
												assign node3317 = (inp[8]) ? node3335 : node3318;
													assign node3318 = (inp[7]) ? node3330 : node3319;
														assign node3319 = (inp[0]) ? node3325 : node3320;
															assign node3320 = (inp[5]) ? 4'b1110 : node3321;
																assign node3321 = (inp[15]) ? 4'b1100 : 4'b1110;
															assign node3325 = (inp[15]) ? node3327 : 4'b1100;
																assign node3327 = (inp[5]) ? 4'b1100 : 4'b1110;
														assign node3330 = (inp[5]) ? node3332 : 4'b1101;
															assign node3332 = (inp[0]) ? 4'b1111 : 4'b1101;
													assign node3335 = (inp[7]) ? node3339 : node3336;
														assign node3336 = (inp[15]) ? 4'b1111 : 4'b1101;
														assign node3339 = (inp[5]) ? node3345 : node3340;
															assign node3340 = (inp[0]) ? node3342 : 4'b1110;
																assign node3342 = (inp[15]) ? 4'b1110 : 4'b1100;
															assign node3345 = (inp[15]) ? node3349 : node3346;
																assign node3346 = (inp[0]) ? 4'b1110 : 4'b1100;
																assign node3349 = (inp[0]) ? 4'b1100 : 4'b1110;
												assign node3352 = (inp[5]) ? node3372 : node3353;
													assign node3353 = (inp[7]) ? node3365 : node3354;
														assign node3354 = (inp[8]) ? node3360 : node3355;
															assign node3355 = (inp[0]) ? 4'b1110 : node3356;
																assign node3356 = (inp[15]) ? 4'b1100 : 4'b1110;
															assign node3360 = (inp[0]) ? node3362 : 4'b1101;
																assign node3362 = (inp[15]) ? 4'b1111 : 4'b1101;
														assign node3365 = (inp[8]) ? 4'b1110 : node3366;
															assign node3366 = (inp[0]) ? 4'b1101 : node3367;
																assign node3367 = (inp[15]) ? 4'b1101 : 4'b1111;
													assign node3372 = (inp[0]) ? node3388 : node3373;
														assign node3373 = (inp[15]) ? node3381 : node3374;
															assign node3374 = (inp[7]) ? node3378 : node3375;
																assign node3375 = (inp[8]) ? 4'b1101 : 4'b1100;
																assign node3378 = (inp[8]) ? 4'b1100 : 4'b1101;
															assign node3381 = (inp[7]) ? node3385 : node3382;
																assign node3382 = (inp[8]) ? 4'b1111 : 4'b1110;
																assign node3385 = (inp[8]) ? 4'b1110 : 4'b1111;
														assign node3388 = (inp[15]) ? node3396 : node3389;
															assign node3389 = (inp[8]) ? node3393 : node3390;
																assign node3390 = (inp[7]) ? 4'b1111 : 4'b1110;
																assign node3393 = (inp[7]) ? 4'b1110 : 4'b1111;
															assign node3396 = (inp[8]) ? node3398 : 4'b1100;
																assign node3398 = (inp[7]) ? 4'b1100 : 4'b1101;
											assign node3401 = (inp[15]) ? node3439 : node3402;
												assign node3402 = (inp[7]) ? node3418 : node3403;
													assign node3403 = (inp[8]) ? node3411 : node3404;
														assign node3404 = (inp[5]) ? node3408 : node3405;
															assign node3405 = (inp[0]) ? 4'b1000 : 4'b1010;
															assign node3408 = (inp[0]) ? 4'b1010 : 4'b1000;
														assign node3411 = (inp[0]) ? node3415 : node3412;
															assign node3412 = (inp[5]) ? 4'b1001 : 4'b1011;
															assign node3415 = (inp[5]) ? 4'b1011 : 4'b1001;
													assign node3418 = (inp[8]) ? node3432 : node3419;
														assign node3419 = (inp[14]) ? node3427 : node3420;
															assign node3420 = (inp[0]) ? node3424 : node3421;
																assign node3421 = (inp[5]) ? 4'b1001 : 4'b1011;
																assign node3424 = (inp[5]) ? 4'b1011 : 4'b1001;
															assign node3427 = (inp[5]) ? node3429 : 4'b1011;
																assign node3429 = (inp[0]) ? 4'b1011 : 4'b1001;
														assign node3432 = (inp[5]) ? node3436 : node3433;
															assign node3433 = (inp[0]) ? 4'b1000 : 4'b1010;
															assign node3436 = (inp[0]) ? 4'b1010 : 4'b1000;
												assign node3439 = (inp[14]) ? node3463 : node3440;
													assign node3440 = (inp[8]) ? node3454 : node3441;
														assign node3441 = (inp[7]) ? node3447 : node3442;
															assign node3442 = (inp[5]) ? node3444 : 4'b1010;
																assign node3444 = (inp[0]) ? 4'b1000 : 4'b1010;
															assign node3447 = (inp[5]) ? node3451 : node3448;
																assign node3448 = (inp[0]) ? 4'b1011 : 4'b1001;
																assign node3451 = (inp[0]) ? 4'b1001 : 4'b1011;
														assign node3454 = (inp[7]) ? node3460 : node3455;
															assign node3455 = (inp[5]) ? node3457 : 4'b1001;
																assign node3457 = (inp[0]) ? 4'b1001 : 4'b1011;
															assign node3460 = (inp[0]) ? 4'b1010 : 4'b1000;
													assign node3463 = (inp[8]) ? node3475 : node3464;
														assign node3464 = (inp[7]) ? node3470 : node3465;
															assign node3465 = (inp[5]) ? node3467 : 4'b1000;
																assign node3467 = (inp[0]) ? 4'b1000 : 4'b1010;
															assign node3470 = (inp[5]) ? 4'b1001 : node3471;
																assign node3471 = (inp[0]) ? 4'b1011 : 4'b1001;
														assign node3475 = (inp[7]) ? node3483 : node3476;
															assign node3476 = (inp[5]) ? node3480 : node3477;
																assign node3477 = (inp[0]) ? 4'b1011 : 4'b1001;
																assign node3480 = (inp[0]) ? 4'b1001 : 4'b1011;
															assign node3483 = (inp[5]) ? node3487 : node3484;
																assign node3484 = (inp[0]) ? 4'b1010 : 4'b1000;
																assign node3487 = (inp[0]) ? 4'b1000 : 4'b1010;
							assign node3490 = (inp[8]) ? node4008 : node3491;
								assign node3491 = (inp[7]) ? node3713 : node3492;
									assign node3492 = (inp[4]) ? node3644 : node3493;
										assign node3493 = (inp[9]) ? node3561 : node3494;
											assign node3494 = (inp[12]) ? node3524 : node3495;
												assign node3495 = (inp[0]) ? node3517 : node3496;
													assign node3496 = (inp[14]) ? node3510 : node3497;
														assign node3497 = (inp[10]) ? node3503 : node3498;
															assign node3498 = (inp[15]) ? node3500 : 4'b1100;
																assign node3500 = (inp[5]) ? 4'b1110 : 4'b1100;
															assign node3503 = (inp[5]) ? node3507 : node3504;
																assign node3504 = (inp[15]) ? 4'b1100 : 4'b1110;
																assign node3507 = (inp[15]) ? 4'b1110 : 4'b1100;
														assign node3510 = (inp[15]) ? node3514 : node3511;
															assign node3511 = (inp[5]) ? 4'b1100 : 4'b1110;
															assign node3514 = (inp[5]) ? 4'b1110 : 4'b1100;
													assign node3517 = (inp[15]) ? node3521 : node3518;
														assign node3518 = (inp[5]) ? 4'b1110 : 4'b1100;
														assign node3521 = (inp[5]) ? 4'b1100 : 4'b1110;
												assign node3524 = (inp[10]) ? node3548 : node3525;
													assign node3525 = (inp[0]) ? node3535 : node3526;
														assign node3526 = (inp[14]) ? node3532 : node3527;
															assign node3527 = (inp[5]) ? 4'b1110 : node3528;
																assign node3528 = (inp[15]) ? 4'b1100 : 4'b1110;
															assign node3532 = (inp[15]) ? 4'b1110 : 4'b1100;
														assign node3535 = (inp[14]) ? node3543 : node3536;
															assign node3536 = (inp[5]) ? node3540 : node3537;
																assign node3537 = (inp[15]) ? 4'b1110 : 4'b1100;
																assign node3540 = (inp[15]) ? 4'b1100 : 4'b1110;
															assign node3543 = (inp[15]) ? node3545 : 4'b1100;
																assign node3545 = (inp[5]) ? 4'b1100 : 4'b1110;
													assign node3548 = (inp[15]) ? node3554 : node3549;
														assign node3549 = (inp[0]) ? 4'b1000 : node3550;
															assign node3550 = (inp[5]) ? 4'b1000 : 4'b1010;
														assign node3554 = (inp[0]) ? node3558 : node3555;
															assign node3555 = (inp[5]) ? 4'b1010 : 4'b1000;
															assign node3558 = (inp[5]) ? 4'b1000 : 4'b1010;
											assign node3561 = (inp[12]) ? node3615 : node3562;
												assign node3562 = (inp[15]) ? node3592 : node3563;
													assign node3563 = (inp[14]) ? node3579 : node3564;
														assign node3564 = (inp[10]) ? node3572 : node3565;
															assign node3565 = (inp[0]) ? node3569 : node3566;
																assign node3566 = (inp[5]) ? 4'b1000 : 4'b1010;
																assign node3569 = (inp[5]) ? 4'b1010 : 4'b1000;
															assign node3572 = (inp[0]) ? node3576 : node3573;
																assign node3573 = (inp[5]) ? 4'b1000 : 4'b1010;
																assign node3576 = (inp[5]) ? 4'b1010 : 4'b1000;
														assign node3579 = (inp[10]) ? node3587 : node3580;
															assign node3580 = (inp[5]) ? node3584 : node3581;
																assign node3581 = (inp[0]) ? 4'b1000 : 4'b1010;
																assign node3584 = (inp[0]) ? 4'b1010 : 4'b1000;
															assign node3587 = (inp[0]) ? node3589 : 4'b1010;
																assign node3589 = (inp[5]) ? 4'b1010 : 4'b1000;
													assign node3592 = (inp[14]) ? node3608 : node3593;
														assign node3593 = (inp[10]) ? node3601 : node3594;
															assign node3594 = (inp[5]) ? node3598 : node3595;
																assign node3595 = (inp[0]) ? 4'b1010 : 4'b1000;
																assign node3598 = (inp[0]) ? 4'b1000 : 4'b1010;
															assign node3601 = (inp[5]) ? node3605 : node3602;
																assign node3602 = (inp[0]) ? 4'b1010 : 4'b1000;
																assign node3605 = (inp[0]) ? 4'b1000 : 4'b1010;
														assign node3608 = (inp[5]) ? node3612 : node3609;
															assign node3609 = (inp[0]) ? 4'b1010 : 4'b1000;
															assign node3612 = (inp[0]) ? 4'b1000 : 4'b1010;
												assign node3615 = (inp[10]) ? node3637 : node3616;
													assign node3616 = (inp[14]) ? node3630 : node3617;
														assign node3617 = (inp[15]) ? node3625 : node3618;
															assign node3618 = (inp[0]) ? node3622 : node3619;
																assign node3619 = (inp[5]) ? 4'b1000 : 4'b1010;
																assign node3622 = (inp[5]) ? 4'b1010 : 4'b1000;
															assign node3625 = (inp[5]) ? node3627 : 4'b1000;
																assign node3627 = (inp[0]) ? 4'b1000 : 4'b1010;
														assign node3630 = (inp[0]) ? 4'b1010 : node3631;
															assign node3631 = (inp[15]) ? 4'b1010 : node3632;
																assign node3632 = (inp[5]) ? 4'b1000 : 4'b1010;
													assign node3637 = (inp[15]) ? node3641 : node3638;
														assign node3638 = (inp[0]) ? 4'b1110 : 4'b1100;
														assign node3641 = (inp[0]) ? 4'b1100 : 4'b1110;
										assign node3644 = (inp[9]) ? node3682 : node3645;
											assign node3645 = (inp[10]) ? node3661 : node3646;
												assign node3646 = (inp[15]) ? node3654 : node3647;
													assign node3647 = (inp[5]) ? node3651 : node3648;
														assign node3648 = (inp[0]) ? 4'b1000 : 4'b1010;
														assign node3651 = (inp[0]) ? 4'b1010 : 4'b1000;
													assign node3654 = (inp[5]) ? node3658 : node3655;
														assign node3655 = (inp[0]) ? 4'b1010 : 4'b1000;
														assign node3658 = (inp[0]) ? 4'b1000 : 4'b1010;
												assign node3661 = (inp[12]) ? node3675 : node3662;
													assign node3662 = (inp[0]) ? node3668 : node3663;
														assign node3663 = (inp[5]) ? node3665 : 4'b1000;
															assign node3665 = (inp[14]) ? 4'b1010 : 4'b1000;
														assign node3668 = (inp[5]) ? node3672 : node3669;
															assign node3669 = (inp[15]) ? 4'b1010 : 4'b1000;
															assign node3672 = (inp[15]) ? 4'b1000 : 4'b1010;
													assign node3675 = (inp[0]) ? node3679 : node3676;
														assign node3676 = (inp[15]) ? 4'b1110 : 4'b1100;
														assign node3679 = (inp[15]) ? 4'b1100 : 4'b1110;
											assign node3682 = (inp[10]) ? node3698 : node3683;
												assign node3683 = (inp[14]) ? node3691 : node3684;
													assign node3684 = (inp[15]) ? node3688 : node3685;
														assign node3685 = (inp[0]) ? 4'b1110 : 4'b1100;
														assign node3688 = (inp[0]) ? 4'b1100 : 4'b1110;
													assign node3691 = (inp[15]) ? node3695 : node3692;
														assign node3692 = (inp[0]) ? 4'b1110 : 4'b1100;
														assign node3695 = (inp[0]) ? 4'b1100 : 4'b1110;
												assign node3698 = (inp[12]) ? node3706 : node3699;
													assign node3699 = (inp[0]) ? node3703 : node3700;
														assign node3700 = (inp[15]) ? 4'b1110 : 4'b1100;
														assign node3703 = (inp[15]) ? 4'b1100 : 4'b1110;
													assign node3706 = (inp[15]) ? node3710 : node3707;
														assign node3707 = (inp[0]) ? 4'b1010 : 4'b1000;
														assign node3710 = (inp[0]) ? 4'b1000 : 4'b1010;
									assign node3713 = (inp[14]) ? node3851 : node3714;
										assign node3714 = (inp[0]) ? node3782 : node3715;
											assign node3715 = (inp[15]) ? node3747 : node3716;
												assign node3716 = (inp[5]) ? node3730 : node3717;
													assign node3717 = (inp[9]) ? node3721 : node3718;
														assign node3718 = (inp[10]) ? 4'b1011 : 4'b1111;
														assign node3721 = (inp[12]) ? node3723 : 4'b1011;
															assign node3723 = (inp[10]) ? node3727 : node3724;
																assign node3724 = (inp[4]) ? 4'b1101 : 4'b1011;
																assign node3727 = (inp[4]) ? 4'b1001 : 4'b1101;
													assign node3730 = (inp[9]) ? node3736 : node3731;
														assign node3731 = (inp[12]) ? 4'b1101 : node3732;
															assign node3732 = (inp[4]) ? 4'b1001 : 4'b1101;
														assign node3736 = (inp[4]) ? node3742 : node3737;
															assign node3737 = (inp[10]) ? node3739 : 4'b1001;
																assign node3739 = (inp[12]) ? 4'b1101 : 4'b1001;
															assign node3742 = (inp[10]) ? node3744 : 4'b1101;
																assign node3744 = (inp[12]) ? 4'b1001 : 4'b1101;
												assign node3747 = (inp[5]) ? node3765 : node3748;
													assign node3748 = (inp[4]) ? node3760 : node3749;
														assign node3749 = (inp[9]) ? node3755 : node3750;
															assign node3750 = (inp[12]) ? node3752 : 4'b1101;
																assign node3752 = (inp[10]) ? 4'b1001 : 4'b1101;
															assign node3755 = (inp[12]) ? node3757 : 4'b1001;
																assign node3757 = (inp[10]) ? 4'b1111 : 4'b1001;
														assign node3760 = (inp[9]) ? node3762 : 4'b1001;
															assign node3762 = (inp[12]) ? 4'b1011 : 4'b1111;
													assign node3765 = (inp[10]) ? node3769 : node3766;
														assign node3766 = (inp[4]) ? 4'b1111 : 4'b1011;
														assign node3769 = (inp[12]) ? node3777 : node3770;
															assign node3770 = (inp[9]) ? node3774 : node3771;
																assign node3771 = (inp[4]) ? 4'b1011 : 4'b1111;
																assign node3774 = (inp[4]) ? 4'b1111 : 4'b1011;
															assign node3777 = (inp[4]) ? 4'b1011 : node3778;
																assign node3778 = (inp[9]) ? 4'b1111 : 4'b1011;
											assign node3782 = (inp[15]) ? node3814 : node3783;
												assign node3783 = (inp[5]) ? node3801 : node3784;
													assign node3784 = (inp[9]) ? node3794 : node3785;
														assign node3785 = (inp[4]) ? node3789 : node3786;
															assign node3786 = (inp[10]) ? 4'b1001 : 4'b1101;
															assign node3789 = (inp[12]) ? node3791 : 4'b1001;
																assign node3791 = (inp[10]) ? 4'b1111 : 4'b1001;
														assign node3794 = (inp[4]) ? node3796 : 4'b1001;
															assign node3796 = (inp[12]) ? node3798 : 4'b1111;
																assign node3798 = (inp[10]) ? 4'b1011 : 4'b1111;
													assign node3801 = (inp[9]) ? 4'b1011 : node3802;
														assign node3802 = (inp[4]) ? node3808 : node3803;
															assign node3803 = (inp[12]) ? node3805 : 4'b1111;
																assign node3805 = (inp[10]) ? 4'b1011 : 4'b1111;
															assign node3808 = (inp[10]) ? node3810 : 4'b1011;
																assign node3810 = (inp[12]) ? 4'b1111 : 4'b1011;
												assign node3814 = (inp[5]) ? node3834 : node3815;
													assign node3815 = (inp[12]) ? node3821 : node3816;
														assign node3816 = (inp[4]) ? 4'b1011 : node3817;
															assign node3817 = (inp[9]) ? 4'b1011 : 4'b1111;
														assign node3821 = (inp[4]) ? node3829 : node3822;
															assign node3822 = (inp[10]) ? node3826 : node3823;
																assign node3823 = (inp[9]) ? 4'b1011 : 4'b1111;
																assign node3826 = (inp[9]) ? 4'b1101 : 4'b1011;
															assign node3829 = (inp[9]) ? 4'b1101 : node3830;
																assign node3830 = (inp[10]) ? 4'b1101 : 4'b1011;
													assign node3834 = (inp[4]) ? node3840 : node3835;
														assign node3835 = (inp[9]) ? 4'b1001 : node3836;
															assign node3836 = (inp[12]) ? 4'b1001 : 4'b1101;
														assign node3840 = (inp[9]) ? node3846 : node3841;
															assign node3841 = (inp[10]) ? node3843 : 4'b1001;
																assign node3843 = (inp[12]) ? 4'b1101 : 4'b1001;
															assign node3846 = (inp[12]) ? node3848 : 4'b1101;
																assign node3848 = (inp[10]) ? 4'b1001 : 4'b1101;
										assign node3851 = (inp[5]) ? node3925 : node3852;
											assign node3852 = (inp[15]) ? node3896 : node3853;
												assign node3853 = (inp[0]) ? node3873 : node3854;
													assign node3854 = (inp[4]) ? node3866 : node3855;
														assign node3855 = (inp[9]) ? node3861 : node3856;
															assign node3856 = (inp[12]) ? node3858 : 4'b1111;
																assign node3858 = (inp[10]) ? 4'b1011 : 4'b1111;
															assign node3861 = (inp[10]) ? node3863 : 4'b1011;
																assign node3863 = (inp[12]) ? 4'b1101 : 4'b1011;
														assign node3866 = (inp[9]) ? 4'b1101 : node3867;
															assign node3867 = (inp[12]) ? node3869 : 4'b1011;
																assign node3869 = (inp[10]) ? 4'b1101 : 4'b1011;
													assign node3873 = (inp[4]) ? node3885 : node3874;
														assign node3874 = (inp[9]) ? node3880 : node3875;
															assign node3875 = (inp[10]) ? node3877 : 4'b1101;
																assign node3877 = (inp[12]) ? 4'b1001 : 4'b1101;
															assign node3880 = (inp[12]) ? node3882 : 4'b1001;
																assign node3882 = (inp[10]) ? 4'b1111 : 4'b1001;
														assign node3885 = (inp[9]) ? node3891 : node3886;
															assign node3886 = (inp[10]) ? node3888 : 4'b1001;
																assign node3888 = (inp[12]) ? 4'b1111 : 4'b1001;
															assign node3891 = (inp[10]) ? node3893 : 4'b1111;
																assign node3893 = (inp[12]) ? 4'b1011 : 4'b1111;
												assign node3896 = (inp[0]) ? node3908 : node3897;
													assign node3897 = (inp[4]) ? node3903 : node3898;
														assign node3898 = (inp[9]) ? 4'b1001 : node3899;
															assign node3899 = (inp[12]) ? 4'b1001 : 4'b1101;
														assign node3903 = (inp[9]) ? node3905 : 4'b1001;
															assign node3905 = (inp[12]) ? 4'b1011 : 4'b1111;
													assign node3908 = (inp[9]) ? node3920 : node3909;
														assign node3909 = (inp[4]) ? node3915 : node3910;
															assign node3910 = (inp[10]) ? node3912 : 4'b1111;
																assign node3912 = (inp[12]) ? 4'b1011 : 4'b1111;
															assign node3915 = (inp[12]) ? node3917 : 4'b1011;
																assign node3917 = (inp[10]) ? 4'b1101 : 4'b1011;
														assign node3920 = (inp[4]) ? 4'b1101 : node3921;
															assign node3921 = (inp[10]) ? 4'b1101 : 4'b1011;
											assign node3925 = (inp[9]) ? node3973 : node3926;
												assign node3926 = (inp[4]) ? node3952 : node3927;
													assign node3927 = (inp[12]) ? node3943 : node3928;
														assign node3928 = (inp[10]) ? node3936 : node3929;
															assign node3929 = (inp[0]) ? node3933 : node3930;
																assign node3930 = (inp[15]) ? 4'b1111 : 4'b1101;
																assign node3933 = (inp[15]) ? 4'b1101 : 4'b1111;
															assign node3936 = (inp[15]) ? node3940 : node3937;
																assign node3937 = (inp[0]) ? 4'b1111 : 4'b1101;
																assign node3940 = (inp[0]) ? 4'b1101 : 4'b1111;
														assign node3943 = (inp[10]) ? 4'b1001 : node3944;
															assign node3944 = (inp[15]) ? node3948 : node3945;
																assign node3945 = (inp[0]) ? 4'b1111 : 4'b1101;
																assign node3948 = (inp[0]) ? 4'b1101 : 4'b1111;
													assign node3952 = (inp[10]) ? node3964 : node3953;
														assign node3953 = (inp[12]) ? node3959 : node3954;
															assign node3954 = (inp[15]) ? 4'b1011 : node3955;
																assign node3955 = (inp[0]) ? 4'b1011 : 4'b1001;
															assign node3959 = (inp[15]) ? node3961 : 4'b1001;
																assign node3961 = (inp[0]) ? 4'b1001 : 4'b1011;
														assign node3964 = (inp[12]) ? node3968 : node3965;
															assign node3965 = (inp[15]) ? 4'b1001 : 4'b1011;
															assign node3968 = (inp[15]) ? node3970 : 4'b1101;
																assign node3970 = (inp[0]) ? 4'b1101 : 4'b1111;
												assign node3973 = (inp[4]) ? node3993 : node3974;
													assign node3974 = (inp[10]) ? node3982 : node3975;
														assign node3975 = (inp[15]) ? node3979 : node3976;
															assign node3976 = (inp[0]) ? 4'b1011 : 4'b1001;
															assign node3979 = (inp[0]) ? 4'b1001 : 4'b1011;
														assign node3982 = (inp[12]) ? node3988 : node3983;
															assign node3983 = (inp[0]) ? 4'b1011 : node3984;
																assign node3984 = (inp[15]) ? 4'b1011 : 4'b1001;
															assign node3988 = (inp[0]) ? 4'b1111 : node3989;
																assign node3989 = (inp[15]) ? 4'b1111 : 4'b1101;
													assign node3993 = (inp[10]) ? node4001 : node3994;
														assign node3994 = (inp[0]) ? node3998 : node3995;
															assign node3995 = (inp[15]) ? 4'b1111 : 4'b1101;
															assign node3998 = (inp[15]) ? 4'b1101 : 4'b1111;
														assign node4001 = (inp[12]) ? node4003 : 4'b1101;
															assign node4003 = (inp[15]) ? 4'b1001 : node4004;
																assign node4004 = (inp[0]) ? 4'b1011 : 4'b1001;
								assign node4008 = (inp[7]) ? node4256 : node4009;
									assign node4009 = (inp[10]) ? node4095 : node4010;
										assign node4010 = (inp[15]) ? node4054 : node4011;
											assign node4011 = (inp[0]) ? node4031 : node4012;
												assign node4012 = (inp[5]) ? node4020 : node4013;
													assign node4013 = (inp[4]) ? node4017 : node4014;
														assign node4014 = (inp[9]) ? 4'b1011 : 4'b1111;
														assign node4017 = (inp[9]) ? 4'b1101 : 4'b1011;
													assign node4020 = (inp[14]) ? node4026 : node4021;
														assign node4021 = (inp[9]) ? node4023 : 4'b1101;
															assign node4023 = (inp[4]) ? 4'b1101 : 4'b1001;
														assign node4026 = (inp[9]) ? 4'b1101 : node4027;
															assign node4027 = (inp[4]) ? 4'b1001 : 4'b1101;
												assign node4031 = (inp[5]) ? node4039 : node4032;
													assign node4032 = (inp[4]) ? node4036 : node4033;
														assign node4033 = (inp[9]) ? 4'b1001 : 4'b1101;
														assign node4036 = (inp[9]) ? 4'b1111 : 4'b1001;
													assign node4039 = (inp[12]) ? node4049 : node4040;
														assign node4040 = (inp[14]) ? node4044 : node4041;
															assign node4041 = (inp[4]) ? 4'b1111 : 4'b1011;
															assign node4044 = (inp[4]) ? 4'b1011 : node4045;
																assign node4045 = (inp[9]) ? 4'b1011 : 4'b1111;
														assign node4049 = (inp[9]) ? 4'b1111 : node4050;
															assign node4050 = (inp[14]) ? 4'b1111 : 4'b1011;
											assign node4054 = (inp[0]) ? node4072 : node4055;
												assign node4055 = (inp[5]) ? node4063 : node4056;
													assign node4056 = (inp[4]) ? node4060 : node4057;
														assign node4057 = (inp[9]) ? 4'b1001 : 4'b1101;
														assign node4060 = (inp[9]) ? 4'b1111 : 4'b1001;
													assign node4063 = (inp[12]) ? 4'b1011 : node4064;
														assign node4064 = (inp[4]) ? node4068 : node4065;
															assign node4065 = (inp[9]) ? 4'b1011 : 4'b1111;
															assign node4068 = (inp[9]) ? 4'b1111 : 4'b1011;
												assign node4072 = (inp[5]) ? node4080 : node4073;
													assign node4073 = (inp[4]) ? node4077 : node4074;
														assign node4074 = (inp[9]) ? 4'b1011 : 4'b1111;
														assign node4077 = (inp[9]) ? 4'b1101 : 4'b1011;
													assign node4080 = (inp[14]) ? node4086 : node4081;
														assign node4081 = (inp[9]) ? 4'b1101 : node4082;
															assign node4082 = (inp[4]) ? 4'b1001 : 4'b1101;
														assign node4086 = (inp[12]) ? 4'b1001 : node4087;
															assign node4087 = (inp[9]) ? node4091 : node4088;
																assign node4088 = (inp[4]) ? 4'b1001 : 4'b1101;
																assign node4091 = (inp[4]) ? 4'b1101 : 4'b1001;
										assign node4095 = (inp[5]) ? node4185 : node4096;
											assign node4096 = (inp[14]) ? node4136 : node4097;
												assign node4097 = (inp[0]) ? node4113 : node4098;
													assign node4098 = (inp[15]) ? node4104 : node4099;
														assign node4099 = (inp[9]) ? 4'b1011 : node4100;
															assign node4100 = (inp[12]) ? 4'b1011 : 4'b1111;
														assign node4104 = (inp[12]) ? node4108 : node4105;
															assign node4105 = (inp[4]) ? 4'b1111 : 4'b1101;
															assign node4108 = (inp[9]) ? node4110 : 4'b1111;
																assign node4110 = (inp[4]) ? 4'b1011 : 4'b1111;
													assign node4113 = (inp[15]) ? node4125 : node4114;
														assign node4114 = (inp[9]) ? node4120 : node4115;
															assign node4115 = (inp[4]) ? 4'b1111 : node4116;
																assign node4116 = (inp[12]) ? 4'b1001 : 4'b1101;
															assign node4120 = (inp[4]) ? node4122 : 4'b1111;
																assign node4122 = (inp[12]) ? 4'b1011 : 4'b1111;
														assign node4125 = (inp[9]) ? node4129 : node4126;
															assign node4126 = (inp[4]) ? 4'b1011 : 4'b1111;
															assign node4129 = (inp[12]) ? node4133 : node4130;
																assign node4130 = (inp[4]) ? 4'b1101 : 4'b1011;
																assign node4133 = (inp[4]) ? 4'b1001 : 4'b1101;
												assign node4136 = (inp[9]) ? node4158 : node4137;
													assign node4137 = (inp[4]) ? node4145 : node4138;
														assign node4138 = (inp[12]) ? 4'b1011 : node4139;
															assign node4139 = (inp[15]) ? 4'b1111 : node4140;
																assign node4140 = (inp[0]) ? 4'b1101 : 4'b1111;
														assign node4145 = (inp[12]) ? node4151 : node4146;
															assign node4146 = (inp[15]) ? node4148 : 4'b1011;
																assign node4148 = (inp[0]) ? 4'b1011 : 4'b1001;
															assign node4151 = (inp[0]) ? node4155 : node4152;
																assign node4152 = (inp[15]) ? 4'b1111 : 4'b1101;
																assign node4155 = (inp[15]) ? 4'b1101 : 4'b1111;
													assign node4158 = (inp[0]) ? node4172 : node4159;
														assign node4159 = (inp[15]) ? node4167 : node4160;
															assign node4160 = (inp[12]) ? node4164 : node4161;
																assign node4161 = (inp[4]) ? 4'b1101 : 4'b1011;
																assign node4164 = (inp[4]) ? 4'b1001 : 4'b1101;
															assign node4167 = (inp[12]) ? node4169 : 4'b1001;
																assign node4169 = (inp[4]) ? 4'b1011 : 4'b1111;
														assign node4172 = (inp[15]) ? node4178 : node4173;
															assign node4173 = (inp[12]) ? node4175 : 4'b1111;
																assign node4175 = (inp[4]) ? 4'b1011 : 4'b1111;
															assign node4178 = (inp[4]) ? node4182 : node4179;
																assign node4179 = (inp[12]) ? 4'b1101 : 4'b1011;
																assign node4182 = (inp[12]) ? 4'b1001 : 4'b1101;
											assign node4185 = (inp[15]) ? node4225 : node4186;
												assign node4186 = (inp[0]) ? node4208 : node4187;
													assign node4187 = (inp[12]) ? node4197 : node4188;
														assign node4188 = (inp[14]) ? 4'b1101 : node4189;
															assign node4189 = (inp[9]) ? node4193 : node4190;
																assign node4190 = (inp[4]) ? 4'b1001 : 4'b1101;
																assign node4193 = (inp[4]) ? 4'b1101 : 4'b1001;
														assign node4197 = (inp[14]) ? node4203 : node4198;
															assign node4198 = (inp[4]) ? node4200 : 4'b1101;
																assign node4200 = (inp[9]) ? 4'b1001 : 4'b1101;
															assign node4203 = (inp[4]) ? 4'b1001 : node4204;
																assign node4204 = (inp[9]) ? 4'b1101 : 4'b1001;
													assign node4208 = (inp[14]) ? node4218 : node4209;
														assign node4209 = (inp[9]) ? node4211 : 4'b1111;
															assign node4211 = (inp[12]) ? node4215 : node4212;
																assign node4212 = (inp[4]) ? 4'b1111 : 4'b1011;
																assign node4215 = (inp[4]) ? 4'b1011 : 4'b1111;
														assign node4218 = (inp[4]) ? node4222 : node4219;
															assign node4219 = (inp[12]) ? 4'b1011 : 4'b1111;
															assign node4222 = (inp[12]) ? 4'b1111 : 4'b1011;
												assign node4225 = (inp[0]) ? node4241 : node4226;
													assign node4226 = (inp[4]) ? node4234 : node4227;
														assign node4227 = (inp[9]) ? node4231 : node4228;
															assign node4228 = (inp[12]) ? 4'b1011 : 4'b1111;
															assign node4231 = (inp[12]) ? 4'b1111 : 4'b1011;
														assign node4234 = (inp[12]) ? node4238 : node4235;
															assign node4235 = (inp[9]) ? 4'b1111 : 4'b1011;
															assign node4238 = (inp[9]) ? 4'b1011 : 4'b1111;
													assign node4241 = (inp[9]) ? node4251 : node4242;
														assign node4242 = (inp[14]) ? node4246 : node4243;
															assign node4243 = (inp[12]) ? 4'b1001 : 4'b1101;
															assign node4246 = (inp[12]) ? node4248 : 4'b1001;
																assign node4248 = (inp[4]) ? 4'b1101 : 4'b1001;
														assign node4251 = (inp[12]) ? node4253 : 4'b1001;
															assign node4253 = (inp[4]) ? 4'b1001 : 4'b1101;
									assign node4256 = (inp[0]) ? node4362 : node4257;
										assign node4257 = (inp[15]) ? node4321 : node4258;
											assign node4258 = (inp[5]) ? node4284 : node4259;
												assign node4259 = (inp[9]) ? node4273 : node4260;
													assign node4260 = (inp[4]) ? node4268 : node4261;
														assign node4261 = (inp[14]) ? 4'b1110 : node4262;
															assign node4262 = (inp[10]) ? node4264 : 4'b1110;
																assign node4264 = (inp[12]) ? 4'b1010 : 4'b1110;
														assign node4268 = (inp[12]) ? node4270 : 4'b1010;
															assign node4270 = (inp[10]) ? 4'b1100 : 4'b1010;
													assign node4273 = (inp[4]) ? node4279 : node4274;
														assign node4274 = (inp[12]) ? node4276 : 4'b1010;
															assign node4276 = (inp[10]) ? 4'b1100 : 4'b1010;
														assign node4279 = (inp[12]) ? node4281 : 4'b1100;
															assign node4281 = (inp[10]) ? 4'b1000 : 4'b1100;
												assign node4284 = (inp[10]) ? node4306 : node4285;
													assign node4285 = (inp[12]) ? node4299 : node4286;
														assign node4286 = (inp[14]) ? node4292 : node4287;
															assign node4287 = (inp[9]) ? node4289 : 4'b1100;
																assign node4289 = (inp[4]) ? 4'b1100 : 4'b1000;
															assign node4292 = (inp[4]) ? node4296 : node4293;
																assign node4293 = (inp[9]) ? 4'b1000 : 4'b1100;
																assign node4296 = (inp[9]) ? 4'b1100 : 4'b1000;
														assign node4299 = (inp[4]) ? node4303 : node4300;
															assign node4300 = (inp[9]) ? 4'b1000 : 4'b1100;
															assign node4303 = (inp[9]) ? 4'b1100 : 4'b1000;
													assign node4306 = (inp[9]) ? node4314 : node4307;
														assign node4307 = (inp[4]) ? node4311 : node4308;
															assign node4308 = (inp[12]) ? 4'b1000 : 4'b1100;
															assign node4311 = (inp[12]) ? 4'b1100 : 4'b1000;
														assign node4314 = (inp[12]) ? node4318 : node4315;
															assign node4315 = (inp[4]) ? 4'b1100 : 4'b1000;
															assign node4318 = (inp[4]) ? 4'b1000 : 4'b1100;
											assign node4321 = (inp[5]) ? node4339 : node4322;
												assign node4322 = (inp[4]) ? node4334 : node4323;
													assign node4323 = (inp[9]) ? node4329 : node4324;
														assign node4324 = (inp[10]) ? node4326 : 4'b1100;
															assign node4326 = (inp[12]) ? 4'b1000 : 4'b1100;
														assign node4329 = (inp[10]) ? node4331 : 4'b1000;
															assign node4331 = (inp[14]) ? 4'b1110 : 4'b1000;
													assign node4334 = (inp[9]) ? 4'b1110 : node4335;
														assign node4335 = (inp[12]) ? 4'b1110 : 4'b1000;
												assign node4339 = (inp[9]) ? node4351 : node4340;
													assign node4340 = (inp[4]) ? node4346 : node4341;
														assign node4341 = (inp[10]) ? node4343 : 4'b1110;
															assign node4343 = (inp[12]) ? 4'b1010 : 4'b1110;
														assign node4346 = (inp[12]) ? node4348 : 4'b1010;
															assign node4348 = (inp[14]) ? 4'b1010 : 4'b1110;
													assign node4351 = (inp[4]) ? node4357 : node4352;
														assign node4352 = (inp[10]) ? node4354 : 4'b1010;
															assign node4354 = (inp[12]) ? 4'b1110 : 4'b1010;
														assign node4357 = (inp[12]) ? node4359 : 4'b1110;
															assign node4359 = (inp[10]) ? 4'b1010 : 4'b1110;
										assign node4362 = (inp[15]) ? node4426 : node4363;
											assign node4363 = (inp[5]) ? node4387 : node4364;
												assign node4364 = (inp[9]) ? node4376 : node4365;
													assign node4365 = (inp[4]) ? node4371 : node4366;
														assign node4366 = (inp[12]) ? node4368 : 4'b1100;
															assign node4368 = (inp[10]) ? 4'b1000 : 4'b1100;
														assign node4371 = (inp[12]) ? node4373 : 4'b1000;
															assign node4373 = (inp[10]) ? 4'b1110 : 4'b1000;
													assign node4376 = (inp[4]) ? node4382 : node4377;
														assign node4377 = (inp[10]) ? node4379 : 4'b1000;
															assign node4379 = (inp[12]) ? 4'b1110 : 4'b1000;
														assign node4382 = (inp[10]) ? node4384 : 4'b1110;
															assign node4384 = (inp[12]) ? 4'b1010 : 4'b1110;
												assign node4387 = (inp[12]) ? node4403 : node4388;
													assign node4388 = (inp[10]) ? node4396 : node4389;
														assign node4389 = (inp[9]) ? node4393 : node4390;
															assign node4390 = (inp[4]) ? 4'b1010 : 4'b1110;
															assign node4393 = (inp[4]) ? 4'b1110 : 4'b1010;
														assign node4396 = (inp[4]) ? node4400 : node4397;
															assign node4397 = (inp[9]) ? 4'b1010 : 4'b1110;
															assign node4400 = (inp[9]) ? 4'b1110 : 4'b1010;
													assign node4403 = (inp[10]) ? node4411 : node4404;
														assign node4404 = (inp[14]) ? 4'b1010 : node4405;
															assign node4405 = (inp[4]) ? 4'b1010 : node4406;
																assign node4406 = (inp[9]) ? 4'b1010 : 4'b1110;
														assign node4411 = (inp[14]) ? node4419 : node4412;
															assign node4412 = (inp[9]) ? node4416 : node4413;
																assign node4413 = (inp[4]) ? 4'b1110 : 4'b1010;
																assign node4416 = (inp[4]) ? 4'b1010 : 4'b1110;
															assign node4419 = (inp[9]) ? node4423 : node4420;
																assign node4420 = (inp[4]) ? 4'b1110 : 4'b1010;
																assign node4423 = (inp[4]) ? 4'b1010 : 4'b1110;
											assign node4426 = (inp[5]) ? node4448 : node4427;
												assign node4427 = (inp[4]) ? node4437 : node4428;
													assign node4428 = (inp[9]) ? node4432 : node4429;
														assign node4429 = (inp[10]) ? 4'b1010 : 4'b1110;
														assign node4432 = (inp[12]) ? node4434 : 4'b1010;
															assign node4434 = (inp[10]) ? 4'b1100 : 4'b1010;
													assign node4437 = (inp[9]) ? node4443 : node4438;
														assign node4438 = (inp[10]) ? node4440 : 4'b1010;
															assign node4440 = (inp[12]) ? 4'b1100 : 4'b1010;
														assign node4443 = (inp[12]) ? node4445 : 4'b1100;
															assign node4445 = (inp[10]) ? 4'b1000 : 4'b1100;
												assign node4448 = (inp[10]) ? node4462 : node4449;
													assign node4449 = (inp[14]) ? node4457 : node4450;
														assign node4450 = (inp[4]) ? node4454 : node4451;
															assign node4451 = (inp[9]) ? 4'b1000 : 4'b1100;
															assign node4454 = (inp[9]) ? 4'b1100 : 4'b1000;
														assign node4457 = (inp[9]) ? node4459 : 4'b1000;
															assign node4459 = (inp[4]) ? 4'b1100 : 4'b1000;
													assign node4462 = (inp[12]) ? node4470 : node4463;
														assign node4463 = (inp[9]) ? node4467 : node4464;
															assign node4464 = (inp[4]) ? 4'b1000 : 4'b1100;
															assign node4467 = (inp[4]) ? 4'b1100 : 4'b1000;
														assign node4470 = (inp[4]) ? 4'b1100 : node4471;
															assign node4471 = (inp[9]) ? 4'b1100 : 4'b1000;
					assign node4475 = (inp[8]) ? node6481 : node4476;
						assign node4476 = (inp[7]) ? node5504 : node4477;
							assign node4477 = (inp[2]) ? node5001 : node4478;
								assign node4478 = (inp[14]) ? node4764 : node4479;
									assign node4479 = (inp[15]) ? node4619 : node4480;
										assign node4480 = (inp[0]) ? node4538 : node4481;
											assign node4481 = (inp[5]) ? node4509 : node4482;
												assign node4482 = (inp[4]) ? node4494 : node4483;
													assign node4483 = (inp[9]) ? node4489 : node4484;
														assign node4484 = (inp[10]) ? node4486 : 4'b1111;
															assign node4486 = (inp[12]) ? 4'b1011 : 4'b1111;
														assign node4489 = (inp[12]) ? node4491 : 4'b1011;
															assign node4491 = (inp[10]) ? 4'b1111 : 4'b1011;
													assign node4494 = (inp[3]) ? node4502 : node4495;
														assign node4495 = (inp[9]) ? 4'b1111 : node4496;
															assign node4496 = (inp[10]) ? node4498 : 4'b1011;
																assign node4498 = (inp[12]) ? 4'b1111 : 4'b1011;
														assign node4502 = (inp[9]) ? node4506 : node4503;
															assign node4503 = (inp[10]) ? 4'b1101 : 4'b1011;
															assign node4506 = (inp[10]) ? 4'b1001 : 4'b1101;
												assign node4509 = (inp[3]) ? node4523 : node4510;
													assign node4510 = (inp[9]) ? node4518 : node4511;
														assign node4511 = (inp[4]) ? node4513 : 4'b1111;
															assign node4513 = (inp[12]) ? node4515 : 4'b1011;
																assign node4515 = (inp[10]) ? 4'b1101 : 4'b1011;
														assign node4518 = (inp[4]) ? 4'b1101 : node4519;
															assign node4519 = (inp[12]) ? 4'b1101 : 4'b1011;
													assign node4523 = (inp[4]) ? node4533 : node4524;
														assign node4524 = (inp[9]) ? node4530 : node4525;
															assign node4525 = (inp[12]) ? node4527 : 4'b1101;
																assign node4527 = (inp[10]) ? 4'b1001 : 4'b1101;
															assign node4530 = (inp[12]) ? 4'b1101 : 4'b1001;
														assign node4533 = (inp[12]) ? 4'b1001 : node4534;
															assign node4534 = (inp[9]) ? 4'b1101 : 4'b1001;
											assign node4538 = (inp[3]) ? node4588 : node4539;
												assign node4539 = (inp[5]) ? node4571 : node4540;
													assign node4540 = (inp[12]) ? node4556 : node4541;
														assign node4541 = (inp[10]) ? node4549 : node4542;
															assign node4542 = (inp[9]) ? node4546 : node4543;
																assign node4543 = (inp[4]) ? 4'b1001 : 4'b1101;
																assign node4546 = (inp[4]) ? 4'b1101 : 4'b1001;
															assign node4549 = (inp[4]) ? node4553 : node4550;
																assign node4550 = (inp[9]) ? 4'b1001 : 4'b1101;
																assign node4553 = (inp[9]) ? 4'b1101 : 4'b1001;
														assign node4556 = (inp[10]) ? node4564 : node4557;
															assign node4557 = (inp[4]) ? node4561 : node4558;
																assign node4558 = (inp[9]) ? 4'b1001 : 4'b1101;
																assign node4561 = (inp[9]) ? 4'b1101 : 4'b1001;
															assign node4564 = (inp[9]) ? node4568 : node4565;
																assign node4565 = (inp[4]) ? 4'b1101 : 4'b1001;
																assign node4568 = (inp[4]) ? 4'b1001 : 4'b1101;
													assign node4571 = (inp[9]) ? node4583 : node4572;
														assign node4572 = (inp[4]) ? node4578 : node4573;
															assign node4573 = (inp[12]) ? node4575 : 4'b1101;
																assign node4575 = (inp[10]) ? 4'b1001 : 4'b1101;
															assign node4578 = (inp[10]) ? node4580 : 4'b1001;
																assign node4580 = (inp[12]) ? 4'b1111 : 4'b1001;
														assign node4583 = (inp[4]) ? 4'b1111 : node4584;
															assign node4584 = (inp[12]) ? 4'b1111 : 4'b1001;
												assign node4588 = (inp[5]) ? node4608 : node4589;
													assign node4589 = (inp[9]) ? node4599 : node4590;
														assign node4590 = (inp[4]) ? node4596 : node4591;
															assign node4591 = (inp[10]) ? node4593 : 4'b1101;
																assign node4593 = (inp[12]) ? 4'b1001 : 4'b1101;
															assign node4596 = (inp[12]) ? 4'b1111 : 4'b1001;
														assign node4599 = (inp[10]) ? node4603 : node4600;
															assign node4600 = (inp[4]) ? 4'b1111 : 4'b1001;
															assign node4603 = (inp[12]) ? node4605 : 4'b1111;
																assign node4605 = (inp[4]) ? 4'b1011 : 4'b1111;
													assign node4608 = (inp[4]) ? node4614 : node4609;
														assign node4609 = (inp[9]) ? 4'b1011 : node4610;
															assign node4610 = (inp[10]) ? 4'b1011 : 4'b1111;
														assign node4614 = (inp[9]) ? 4'b1111 : node4615;
															assign node4615 = (inp[10]) ? 4'b1111 : 4'b1011;
										assign node4619 = (inp[0]) ? node4689 : node4620;
											assign node4620 = (inp[5]) ? node4654 : node4621;
												assign node4621 = (inp[3]) ? node4639 : node4622;
													assign node4622 = (inp[4]) ? node4634 : node4623;
														assign node4623 = (inp[9]) ? node4629 : node4624;
															assign node4624 = (inp[12]) ? node4626 : 4'b1101;
																assign node4626 = (inp[10]) ? 4'b1001 : 4'b1101;
															assign node4629 = (inp[10]) ? node4631 : 4'b1001;
																assign node4631 = (inp[12]) ? 4'b1101 : 4'b1001;
														assign node4634 = (inp[9]) ? 4'b1101 : node4635;
															assign node4635 = (inp[12]) ? 4'b1101 : 4'b1001;
													assign node4639 = (inp[9]) ? node4643 : node4640;
														assign node4640 = (inp[4]) ? 4'b1001 : 4'b1101;
														assign node4643 = (inp[4]) ? node4649 : node4644;
															assign node4644 = (inp[10]) ? node4646 : 4'b1001;
																assign node4646 = (inp[12]) ? 4'b1111 : 4'b1001;
															assign node4649 = (inp[12]) ? node4651 : 4'b1111;
																assign node4651 = (inp[10]) ? 4'b1011 : 4'b1111;
												assign node4654 = (inp[3]) ? node4674 : node4655;
													assign node4655 = (inp[4]) ? node4665 : node4656;
														assign node4656 = (inp[10]) ? node4658 : 4'b1001;
															assign node4658 = (inp[9]) ? node4662 : node4659;
																assign node4659 = (inp[12]) ? 4'b1001 : 4'b1101;
																assign node4662 = (inp[12]) ? 4'b1111 : 4'b1001;
														assign node4665 = (inp[9]) ? node4671 : node4666;
															assign node4666 = (inp[12]) ? node4668 : 4'b1001;
																assign node4668 = (inp[10]) ? 4'b1111 : 4'b1001;
															assign node4671 = (inp[12]) ? 4'b1011 : 4'b1111;
													assign node4674 = (inp[9]) ? node4682 : node4675;
														assign node4675 = (inp[4]) ? node4677 : 4'b1111;
															assign node4677 = (inp[12]) ? node4679 : 4'b1011;
																assign node4679 = (inp[10]) ? 4'b1111 : 4'b1011;
														assign node4682 = (inp[4]) ? node4684 : 4'b1011;
															assign node4684 = (inp[12]) ? node4686 : 4'b1111;
																assign node4686 = (inp[10]) ? 4'b1011 : 4'b1111;
											assign node4689 = (inp[3]) ? node4733 : node4690;
												assign node4690 = (inp[5]) ? node4710 : node4691;
													assign node4691 = (inp[9]) ? node4701 : node4692;
														assign node4692 = (inp[4]) ? node4696 : node4693;
															assign node4693 = (inp[12]) ? 4'b1011 : 4'b1111;
															assign node4696 = (inp[12]) ? node4698 : 4'b1011;
																assign node4698 = (inp[10]) ? 4'b1111 : 4'b1011;
														assign node4701 = (inp[4]) ? node4707 : node4702;
															assign node4702 = (inp[12]) ? node4704 : 4'b1011;
																assign node4704 = (inp[10]) ? 4'b1111 : 4'b1011;
															assign node4707 = (inp[10]) ? 4'b1011 : 4'b1111;
													assign node4710 = (inp[9]) ? node4722 : node4711;
														assign node4711 = (inp[4]) ? node4717 : node4712;
															assign node4712 = (inp[10]) ? node4714 : 4'b1111;
																assign node4714 = (inp[12]) ? 4'b1011 : 4'b1111;
															assign node4717 = (inp[12]) ? node4719 : 4'b1011;
																assign node4719 = (inp[10]) ? 4'b1101 : 4'b1011;
														assign node4722 = (inp[4]) ? node4728 : node4723;
															assign node4723 = (inp[12]) ? node4725 : 4'b1011;
																assign node4725 = (inp[10]) ? 4'b1101 : 4'b1011;
															assign node4728 = (inp[12]) ? node4730 : 4'b1101;
																assign node4730 = (inp[10]) ? 4'b1001 : 4'b1101;
												assign node4733 = (inp[5]) ? node4749 : node4734;
													assign node4734 = (inp[4]) ? node4740 : node4735;
														assign node4735 = (inp[12]) ? 4'b1011 : node4736;
															assign node4736 = (inp[9]) ? 4'b1011 : 4'b1111;
														assign node4740 = (inp[10]) ? node4744 : node4741;
															assign node4741 = (inp[9]) ? 4'b1101 : 4'b1011;
															assign node4744 = (inp[9]) ? node4746 : 4'b1101;
																assign node4746 = (inp[12]) ? 4'b1001 : 4'b1101;
													assign node4749 = (inp[4]) ? node4757 : node4750;
														assign node4750 = (inp[9]) ? node4752 : 4'b1101;
															assign node4752 = (inp[12]) ? node4754 : 4'b1001;
																assign node4754 = (inp[10]) ? 4'b1101 : 4'b1001;
														assign node4757 = (inp[9]) ? node4759 : 4'b1001;
															assign node4759 = (inp[10]) ? node4761 : 4'b1101;
																assign node4761 = (inp[12]) ? 4'b1001 : 4'b1101;
									assign node4764 = (inp[4]) ? node4888 : node4765;
										assign node4765 = (inp[9]) ? node4833 : node4766;
											assign node4766 = (inp[10]) ? node4804 : node4767;
												assign node4767 = (inp[12]) ? node4785 : node4768;
													assign node4768 = (inp[15]) ? node4778 : node4769;
														assign node4769 = (inp[0]) ? node4773 : node4770;
															assign node4770 = (inp[3]) ? 4'b1100 : 4'b1110;
															assign node4773 = (inp[3]) ? node4775 : 4'b1100;
																assign node4775 = (inp[5]) ? 4'b1110 : 4'b1100;
														assign node4778 = (inp[0]) ? 4'b1110 : node4779;
															assign node4779 = (inp[3]) ? node4781 : 4'b1100;
																assign node4781 = (inp[5]) ? 4'b1110 : 4'b1100;
													assign node4785 = (inp[5]) ? node4791 : node4786;
														assign node4786 = (inp[0]) ? 4'b1110 : node4787;
															assign node4787 = (inp[15]) ? 4'b1100 : 4'b1110;
														assign node4791 = (inp[3]) ? node4799 : node4792;
															assign node4792 = (inp[15]) ? node4796 : node4793;
																assign node4793 = (inp[0]) ? 4'b1100 : 4'b1110;
																assign node4796 = (inp[0]) ? 4'b1110 : 4'b1100;
															assign node4799 = (inp[0]) ? node4801 : 4'b1110;
																assign node4801 = (inp[15]) ? 4'b1100 : 4'b1110;
												assign node4804 = (inp[12]) ? node4822 : node4805;
													assign node4805 = (inp[5]) ? node4811 : node4806;
														assign node4806 = (inp[15]) ? node4808 : 4'b1110;
															assign node4808 = (inp[0]) ? 4'b1110 : 4'b1100;
														assign node4811 = (inp[15]) ? node4817 : node4812;
															assign node4812 = (inp[3]) ? 4'b1100 : node4813;
																assign node4813 = (inp[0]) ? 4'b1100 : 4'b1110;
															assign node4817 = (inp[0]) ? 4'b1110 : node4818;
																assign node4818 = (inp[3]) ? 4'b1110 : 4'b1100;
													assign node4822 = (inp[0]) ? node4830 : node4823;
														assign node4823 = (inp[15]) ? node4827 : node4824;
															assign node4824 = (inp[3]) ? 4'b1000 : 4'b1010;
															assign node4827 = (inp[5]) ? 4'b1010 : 4'b1000;
														assign node4830 = (inp[15]) ? 4'b1010 : 4'b1000;
											assign node4833 = (inp[12]) ? node4861 : node4834;
												assign node4834 = (inp[3]) ? node4842 : node4835;
													assign node4835 = (inp[0]) ? node4839 : node4836;
														assign node4836 = (inp[15]) ? 4'b1000 : 4'b1010;
														assign node4839 = (inp[15]) ? 4'b1010 : 4'b1000;
													assign node4842 = (inp[0]) ? node4854 : node4843;
														assign node4843 = (inp[10]) ? node4849 : node4844;
															assign node4844 = (inp[15]) ? node4846 : 4'b1000;
																assign node4846 = (inp[5]) ? 4'b1010 : 4'b1000;
															assign node4849 = (inp[15]) ? 4'b1000 : node4850;
																assign node4850 = (inp[5]) ? 4'b1000 : 4'b1010;
														assign node4854 = (inp[15]) ? node4858 : node4855;
															assign node4855 = (inp[5]) ? 4'b1010 : 4'b1000;
															assign node4858 = (inp[5]) ? 4'b1000 : 4'b1010;
												assign node4861 = (inp[10]) ? node4877 : node4862;
													assign node4862 = (inp[5]) ? node4868 : node4863;
														assign node4863 = (inp[15]) ? node4865 : 4'b1000;
															assign node4865 = (inp[0]) ? 4'b1010 : 4'b1000;
														assign node4868 = (inp[0]) ? 4'b1010 : node4869;
															assign node4869 = (inp[3]) ? node4873 : node4870;
																assign node4870 = (inp[15]) ? 4'b1000 : 4'b1010;
																assign node4873 = (inp[15]) ? 4'b1010 : 4'b1000;
													assign node4877 = (inp[15]) ? node4883 : node4878;
														assign node4878 = (inp[0]) ? node4880 : 4'b1100;
															assign node4880 = (inp[3]) ? 4'b1110 : 4'b1100;
														assign node4883 = (inp[0]) ? node4885 : 4'b1110;
															assign node4885 = (inp[3]) ? 4'b1100 : 4'b1110;
										assign node4888 = (inp[9]) ? node4950 : node4889;
											assign node4889 = (inp[10]) ? node4913 : node4890;
												assign node4890 = (inp[15]) ? node4902 : node4891;
													assign node4891 = (inp[0]) ? node4897 : node4892;
														assign node4892 = (inp[5]) ? node4894 : 4'b1010;
															assign node4894 = (inp[3]) ? 4'b1000 : 4'b1010;
														assign node4897 = (inp[5]) ? node4899 : 4'b1000;
															assign node4899 = (inp[3]) ? 4'b1010 : 4'b1000;
													assign node4902 = (inp[0]) ? node4908 : node4903;
														assign node4903 = (inp[5]) ? node4905 : 4'b1000;
															assign node4905 = (inp[3]) ? 4'b1010 : 4'b1000;
														assign node4908 = (inp[5]) ? node4910 : 4'b1010;
															assign node4910 = (inp[3]) ? 4'b1000 : 4'b1010;
												assign node4913 = (inp[12]) ? node4929 : node4914;
													assign node4914 = (inp[0]) ? node4920 : node4915;
														assign node4915 = (inp[3]) ? node4917 : 4'b1000;
															assign node4917 = (inp[15]) ? 4'b1010 : 4'b1000;
														assign node4920 = (inp[15]) ? node4924 : node4921;
															assign node4921 = (inp[3]) ? 4'b1010 : 4'b1000;
															assign node4924 = (inp[5]) ? node4926 : 4'b1010;
																assign node4926 = (inp[3]) ? 4'b1000 : 4'b1010;
													assign node4929 = (inp[5]) ? node4943 : node4930;
														assign node4930 = (inp[15]) ? node4938 : node4931;
															assign node4931 = (inp[0]) ? node4935 : node4932;
																assign node4932 = (inp[3]) ? 4'b1100 : 4'b1110;
																assign node4935 = (inp[3]) ? 4'b1110 : 4'b1100;
															assign node4938 = (inp[3]) ? 4'b1110 : node4939;
																assign node4939 = (inp[0]) ? 4'b1110 : 4'b1100;
														assign node4943 = (inp[0]) ? node4947 : node4944;
															assign node4944 = (inp[3]) ? 4'b1100 : 4'b1110;
															assign node4947 = (inp[15]) ? 4'b1100 : 4'b1110;
											assign node4950 = (inp[12]) ? node4972 : node4951;
												assign node4951 = (inp[15]) ? node4963 : node4952;
													assign node4952 = (inp[0]) ? node4958 : node4953;
														assign node4953 = (inp[5]) ? 4'b1100 : node4954;
															assign node4954 = (inp[3]) ? 4'b1100 : 4'b1110;
														assign node4958 = (inp[3]) ? 4'b1110 : node4959;
															assign node4959 = (inp[5]) ? 4'b1110 : 4'b1100;
													assign node4963 = (inp[0]) ? node4967 : node4964;
														assign node4964 = (inp[3]) ? 4'b1110 : 4'b1100;
														assign node4967 = (inp[5]) ? 4'b1100 : node4968;
															assign node4968 = (inp[3]) ? 4'b1100 : 4'b1110;
												assign node4972 = (inp[10]) ? node4990 : node4973;
													assign node4973 = (inp[3]) ? node4977 : node4974;
														assign node4974 = (inp[0]) ? 4'b1100 : 4'b1110;
														assign node4977 = (inp[5]) ? node4985 : node4978;
															assign node4978 = (inp[15]) ? node4982 : node4979;
																assign node4979 = (inp[0]) ? 4'b1110 : 4'b1100;
																assign node4982 = (inp[0]) ? 4'b1100 : 4'b1110;
															assign node4985 = (inp[0]) ? 4'b1110 : node4986;
																assign node4986 = (inp[15]) ? 4'b1110 : 4'b1100;
													assign node4990 = (inp[15]) ? node4996 : node4991;
														assign node4991 = (inp[0]) ? node4993 : 4'b1000;
															assign node4993 = (inp[3]) ? 4'b1010 : 4'b1000;
														assign node4996 = (inp[0]) ? node4998 : 4'b1010;
															assign node4998 = (inp[3]) ? 4'b1000 : 4'b1010;
								assign node5001 = (inp[12]) ? node5253 : node5002;
									assign node5002 = (inp[14]) ? node5108 : node5003;
										assign node5003 = (inp[4]) ? node5039 : node5004;
											assign node5004 = (inp[9]) ? node5022 : node5005;
												assign node5005 = (inp[15]) ? node5015 : node5006;
													assign node5006 = (inp[0]) ? node5010 : node5007;
														assign node5007 = (inp[5]) ? 4'b1100 : 4'b1110;
														assign node5010 = (inp[5]) ? node5012 : 4'b1100;
															assign node5012 = (inp[3]) ? 4'b1110 : 4'b1100;
													assign node5015 = (inp[0]) ? node5017 : 4'b1100;
														assign node5017 = (inp[10]) ? node5019 : 4'b1110;
															assign node5019 = (inp[3]) ? 4'b1100 : 4'b1110;
												assign node5022 = (inp[15]) ? node5028 : node5023;
													assign node5023 = (inp[10]) ? node5025 : 4'b1000;
														assign node5025 = (inp[3]) ? 4'b1000 : 4'b1010;
													assign node5028 = (inp[0]) ? node5034 : node5029;
														assign node5029 = (inp[5]) ? node5031 : 4'b1000;
															assign node5031 = (inp[3]) ? 4'b1010 : 4'b1000;
														assign node5034 = (inp[5]) ? node5036 : 4'b1010;
															assign node5036 = (inp[3]) ? 4'b1000 : 4'b1010;
											assign node5039 = (inp[9]) ? node5079 : node5040;
												assign node5040 = (inp[5]) ? node5062 : node5041;
													assign node5041 = (inp[3]) ? node5055 : node5042;
														assign node5042 = (inp[10]) ? node5048 : node5043;
															assign node5043 = (inp[0]) ? node5045 : 4'b1000;
																assign node5045 = (inp[15]) ? 4'b1010 : 4'b1000;
															assign node5048 = (inp[0]) ? node5052 : node5049;
																assign node5049 = (inp[15]) ? 4'b1000 : 4'b1010;
																assign node5052 = (inp[15]) ? 4'b1010 : 4'b1000;
														assign node5055 = (inp[15]) ? node5059 : node5056;
															assign node5056 = (inp[0]) ? 4'b1000 : 4'b1010;
															assign node5059 = (inp[0]) ? 4'b1010 : 4'b1000;
													assign node5062 = (inp[15]) ? node5070 : node5063;
														assign node5063 = (inp[0]) ? node5067 : node5064;
															assign node5064 = (inp[3]) ? 4'b1000 : 4'b1010;
															assign node5067 = (inp[3]) ? 4'b1010 : 4'b1000;
														assign node5070 = (inp[10]) ? node5074 : node5071;
															assign node5071 = (inp[3]) ? 4'b1000 : 4'b1010;
															assign node5074 = (inp[0]) ? 4'b1000 : node5075;
																assign node5075 = (inp[3]) ? 4'b1010 : 4'b1000;
												assign node5079 = (inp[5]) ? node5089 : node5080;
													assign node5080 = (inp[15]) ? node5082 : 4'b1100;
														assign node5082 = (inp[3]) ? node5086 : node5083;
															assign node5083 = (inp[0]) ? 4'b1110 : 4'b1100;
															assign node5086 = (inp[0]) ? 4'b1100 : 4'b1110;
													assign node5089 = (inp[10]) ? node5099 : node5090;
														assign node5090 = (inp[3]) ? node5092 : 4'b1100;
															assign node5092 = (inp[15]) ? node5096 : node5093;
																assign node5093 = (inp[0]) ? 4'b1110 : 4'b1100;
																assign node5096 = (inp[0]) ? 4'b1100 : 4'b1110;
														assign node5099 = (inp[3]) ? node5101 : 4'b1110;
															assign node5101 = (inp[0]) ? node5105 : node5102;
																assign node5102 = (inp[15]) ? 4'b1110 : 4'b1100;
																assign node5105 = (inp[15]) ? 4'b1100 : 4'b1110;
										assign node5108 = (inp[5]) ? node5192 : node5109;
											assign node5109 = (inp[3]) ? node5151 : node5110;
												assign node5110 = (inp[10]) ? node5130 : node5111;
													assign node5111 = (inp[15]) ? node5125 : node5112;
														assign node5112 = (inp[0]) ? node5120 : node5113;
															assign node5113 = (inp[4]) ? node5117 : node5114;
																assign node5114 = (inp[9]) ? 4'b1010 : 4'b1110;
																assign node5117 = (inp[9]) ? 4'b1110 : 4'b1010;
															assign node5120 = (inp[9]) ? node5122 : 4'b1000;
																assign node5122 = (inp[4]) ? 4'b1100 : 4'b1000;
														assign node5125 = (inp[0]) ? 4'b1110 : node5126;
															assign node5126 = (inp[4]) ? 4'b1100 : 4'b1000;
													assign node5130 = (inp[9]) ? node5144 : node5131;
														assign node5131 = (inp[4]) ? node5139 : node5132;
															assign node5132 = (inp[15]) ? node5136 : node5133;
																assign node5133 = (inp[0]) ? 4'b1100 : 4'b1110;
																assign node5136 = (inp[0]) ? 4'b1110 : 4'b1100;
															assign node5139 = (inp[15]) ? node5141 : 4'b1000;
																assign node5141 = (inp[0]) ? 4'b1010 : 4'b1000;
														assign node5144 = (inp[4]) ? 4'b1110 : node5145;
															assign node5145 = (inp[15]) ? node5147 : 4'b1000;
																assign node5147 = (inp[0]) ? 4'b1010 : 4'b1000;
												assign node5151 = (inp[4]) ? node5173 : node5152;
													assign node5152 = (inp[9]) ? node5166 : node5153;
														assign node5153 = (inp[10]) ? node5161 : node5154;
															assign node5154 = (inp[0]) ? node5158 : node5155;
																assign node5155 = (inp[15]) ? 4'b1100 : 4'b1110;
																assign node5158 = (inp[15]) ? 4'b1110 : 4'b1100;
															assign node5161 = (inp[0]) ? 4'b1110 : node5162;
																assign node5162 = (inp[15]) ? 4'b1100 : 4'b1110;
														assign node5166 = (inp[0]) ? node5170 : node5167;
															assign node5167 = (inp[10]) ? 4'b1010 : 4'b1000;
															assign node5170 = (inp[10]) ? 4'b1000 : 4'b1010;
													assign node5173 = (inp[9]) ? node5185 : node5174;
														assign node5174 = (inp[10]) ? node5180 : node5175;
															assign node5175 = (inp[0]) ? 4'b1000 : node5176;
																assign node5176 = (inp[15]) ? 4'b1000 : 4'b1010;
															assign node5180 = (inp[15]) ? node5182 : 4'b1000;
																assign node5182 = (inp[0]) ? 4'b1010 : 4'b1000;
														assign node5185 = (inp[15]) ? node5189 : node5186;
															assign node5186 = (inp[0]) ? 4'b1110 : 4'b1100;
															assign node5189 = (inp[0]) ? 4'b1100 : 4'b1110;
											assign node5192 = (inp[3]) ? node5226 : node5193;
												assign node5193 = (inp[15]) ? node5211 : node5194;
													assign node5194 = (inp[0]) ? node5206 : node5195;
														assign node5195 = (inp[10]) ? node5201 : node5196;
															assign node5196 = (inp[9]) ? 4'b1010 : node5197;
																assign node5197 = (inp[4]) ? 4'b1010 : 4'b1110;
															assign node5201 = (inp[9]) ? node5203 : 4'b1010;
																assign node5203 = (inp[4]) ? 4'b1100 : 4'b1010;
														assign node5206 = (inp[4]) ? 4'b1000 : node5207;
															assign node5207 = (inp[9]) ? 4'b1000 : 4'b1100;
													assign node5211 = (inp[0]) ? node5219 : node5212;
														assign node5212 = (inp[9]) ? node5216 : node5213;
															assign node5213 = (inp[4]) ? 4'b1000 : 4'b1100;
															assign node5216 = (inp[4]) ? 4'b1110 : 4'b1000;
														assign node5219 = (inp[9]) ? node5223 : node5220;
															assign node5220 = (inp[4]) ? 4'b1010 : 4'b1110;
															assign node5223 = (inp[4]) ? 4'b1100 : 4'b1010;
												assign node5226 = (inp[0]) ? node5240 : node5227;
													assign node5227 = (inp[15]) ? node5235 : node5228;
														assign node5228 = (inp[4]) ? node5232 : node5229;
															assign node5229 = (inp[9]) ? 4'b1000 : 4'b1100;
															assign node5232 = (inp[9]) ? 4'b1100 : 4'b1000;
														assign node5235 = (inp[4]) ? 4'b1110 : node5236;
															assign node5236 = (inp[9]) ? 4'b1010 : 4'b1110;
													assign node5240 = (inp[15]) ? node5248 : node5241;
														assign node5241 = (inp[4]) ? node5245 : node5242;
															assign node5242 = (inp[9]) ? 4'b1010 : 4'b1110;
															assign node5245 = (inp[9]) ? 4'b1110 : 4'b1010;
														assign node5248 = (inp[9]) ? node5250 : 4'b1000;
															assign node5250 = (inp[4]) ? 4'b1100 : 4'b1000;
									assign node5253 = (inp[15]) ? node5383 : node5254;
										assign node5254 = (inp[5]) ? node5310 : node5255;
											assign node5255 = (inp[0]) ? node5287 : node5256;
												assign node5256 = (inp[3]) ? node5272 : node5257;
													assign node5257 = (inp[4]) ? node5265 : node5258;
														assign node5258 = (inp[9]) ? node5262 : node5259;
															assign node5259 = (inp[10]) ? 4'b1010 : 4'b1110;
															assign node5262 = (inp[10]) ? 4'b1110 : 4'b1010;
														assign node5265 = (inp[10]) ? node5269 : node5266;
															assign node5266 = (inp[9]) ? 4'b1110 : 4'b1010;
															assign node5269 = (inp[9]) ? 4'b1010 : 4'b1110;
													assign node5272 = (inp[10]) ? node5280 : node5273;
														assign node5273 = (inp[4]) ? node5277 : node5274;
															assign node5274 = (inp[14]) ? 4'b1010 : 4'b1110;
															assign node5277 = (inp[14]) ? 4'b1100 : 4'b1010;
														assign node5280 = (inp[14]) ? 4'b1100 : node5281;
															assign node5281 = (inp[4]) ? node5283 : 4'b1100;
																assign node5283 = (inp[9]) ? 4'b1000 : 4'b1100;
												assign node5287 = (inp[3]) ? node5297 : node5288;
													assign node5288 = (inp[9]) ? node5290 : 4'b1100;
														assign node5290 = (inp[10]) ? node5294 : node5291;
															assign node5291 = (inp[4]) ? 4'b1100 : 4'b1000;
															assign node5294 = (inp[4]) ? 4'b1000 : 4'b1100;
													assign node5297 = (inp[4]) ? node5305 : node5298;
														assign node5298 = (inp[10]) ? node5302 : node5299;
															assign node5299 = (inp[9]) ? 4'b1000 : 4'b1100;
															assign node5302 = (inp[9]) ? 4'b1110 : 4'b1000;
														assign node5305 = (inp[14]) ? 4'b1110 : node5306;
															assign node5306 = (inp[9]) ? 4'b1010 : 4'b1110;
											assign node5310 = (inp[0]) ? node5344 : node5311;
												assign node5311 = (inp[3]) ? node5325 : node5312;
													assign node5312 = (inp[10]) ? node5320 : node5313;
														assign node5313 = (inp[4]) ? node5317 : node5314;
															assign node5314 = (inp[9]) ? 4'b1010 : 4'b1110;
															assign node5317 = (inp[9]) ? 4'b1100 : 4'b1010;
														assign node5320 = (inp[9]) ? node5322 : 4'b1100;
															assign node5322 = (inp[4]) ? 4'b1000 : 4'b1100;
													assign node5325 = (inp[4]) ? node5339 : node5326;
														assign node5326 = (inp[14]) ? node5334 : node5327;
															assign node5327 = (inp[9]) ? node5331 : node5328;
																assign node5328 = (inp[10]) ? 4'b1000 : 4'b1100;
																assign node5331 = (inp[10]) ? 4'b1100 : 4'b1000;
															assign node5334 = (inp[9]) ? node5336 : 4'b1100;
																assign node5336 = (inp[10]) ? 4'b1100 : 4'b1000;
														assign node5339 = (inp[10]) ? 4'b1000 : node5340;
															assign node5340 = (inp[9]) ? 4'b1100 : 4'b1000;
												assign node5344 = (inp[3]) ? node5360 : node5345;
													assign node5345 = (inp[4]) ? node5353 : node5346;
														assign node5346 = (inp[10]) ? node5350 : node5347;
															assign node5347 = (inp[9]) ? 4'b1000 : 4'b1100;
															assign node5350 = (inp[9]) ? 4'b1110 : 4'b1000;
														assign node5353 = (inp[14]) ? node5355 : 4'b1110;
															assign node5355 = (inp[9]) ? node5357 : 4'b1000;
																assign node5357 = (inp[10]) ? 4'b1010 : 4'b1110;
													assign node5360 = (inp[14]) ? node5374 : node5361;
														assign node5361 = (inp[4]) ? node5367 : node5362;
															assign node5362 = (inp[9]) ? 4'b1010 : node5363;
																assign node5363 = (inp[10]) ? 4'b1010 : 4'b1110;
															assign node5367 = (inp[10]) ? node5371 : node5368;
																assign node5368 = (inp[9]) ? 4'b1110 : 4'b1010;
																assign node5371 = (inp[9]) ? 4'b1010 : 4'b1110;
														assign node5374 = (inp[4]) ? node5376 : 4'b1110;
															assign node5376 = (inp[9]) ? node5380 : node5377;
																assign node5377 = (inp[10]) ? 4'b1110 : 4'b1010;
																assign node5380 = (inp[10]) ? 4'b1010 : 4'b1110;
										assign node5383 = (inp[9]) ? node5451 : node5384;
											assign node5384 = (inp[0]) ? node5416 : node5385;
												assign node5385 = (inp[5]) ? node5395 : node5386;
													assign node5386 = (inp[4]) ? node5390 : node5387;
														assign node5387 = (inp[10]) ? 4'b1000 : 4'b1100;
														assign node5390 = (inp[10]) ? node5392 : 4'b1000;
															assign node5392 = (inp[3]) ? 4'b1110 : 4'b1100;
													assign node5395 = (inp[3]) ? node5403 : node5396;
														assign node5396 = (inp[10]) ? node5400 : node5397;
															assign node5397 = (inp[4]) ? 4'b1000 : 4'b1100;
															assign node5400 = (inp[4]) ? 4'b1110 : 4'b1000;
														assign node5403 = (inp[14]) ? node5411 : node5404;
															assign node5404 = (inp[4]) ? node5408 : node5405;
																assign node5405 = (inp[10]) ? 4'b1010 : 4'b1110;
																assign node5408 = (inp[10]) ? 4'b1110 : 4'b1010;
															assign node5411 = (inp[10]) ? node5413 : 4'b1110;
																assign node5413 = (inp[4]) ? 4'b1110 : 4'b1010;
												assign node5416 = (inp[5]) ? node5436 : node5417;
													assign node5417 = (inp[3]) ? node5425 : node5418;
														assign node5418 = (inp[4]) ? node5422 : node5419;
															assign node5419 = (inp[10]) ? 4'b1010 : 4'b1110;
															assign node5422 = (inp[10]) ? 4'b1110 : 4'b1010;
														assign node5425 = (inp[14]) ? node5431 : node5426;
															assign node5426 = (inp[10]) ? node5428 : 4'b1010;
																assign node5428 = (inp[4]) ? 4'b1100 : 4'b1010;
															assign node5431 = (inp[10]) ? 4'b1010 : node5432;
																assign node5432 = (inp[4]) ? 4'b1010 : 4'b1110;
													assign node5436 = (inp[3]) ? node5444 : node5437;
														assign node5437 = (inp[10]) ? node5441 : node5438;
															assign node5438 = (inp[4]) ? 4'b1010 : 4'b1110;
															assign node5441 = (inp[4]) ? 4'b1100 : 4'b1010;
														assign node5444 = (inp[4]) ? node5448 : node5445;
															assign node5445 = (inp[10]) ? 4'b1000 : 4'b1100;
															assign node5448 = (inp[10]) ? 4'b1100 : 4'b1000;
											assign node5451 = (inp[0]) ? node5481 : node5452;
												assign node5452 = (inp[5]) ? node5474 : node5453;
													assign node5453 = (inp[3]) ? node5467 : node5454;
														assign node5454 = (inp[14]) ? node5462 : node5455;
															assign node5455 = (inp[10]) ? node5459 : node5456;
																assign node5456 = (inp[4]) ? 4'b1100 : 4'b1000;
																assign node5459 = (inp[4]) ? 4'b1000 : 4'b1100;
															assign node5462 = (inp[10]) ? 4'b1000 : node5463;
																assign node5463 = (inp[4]) ? 4'b1100 : 4'b1000;
														assign node5467 = (inp[4]) ? node5471 : node5468;
															assign node5468 = (inp[10]) ? 4'b1110 : 4'b1000;
															assign node5471 = (inp[10]) ? 4'b1010 : 4'b1110;
													assign node5474 = (inp[4]) ? node5478 : node5475;
														assign node5475 = (inp[10]) ? 4'b1110 : 4'b1010;
														assign node5478 = (inp[10]) ? 4'b1010 : 4'b1110;
												assign node5481 = (inp[5]) ? node5495 : node5482;
													assign node5482 = (inp[3]) ? node5490 : node5483;
														assign node5483 = (inp[10]) ? node5487 : node5484;
															assign node5484 = (inp[4]) ? 4'b1110 : 4'b1010;
															assign node5487 = (inp[4]) ? 4'b1010 : 4'b1110;
														assign node5490 = (inp[4]) ? 4'b1100 : node5491;
															assign node5491 = (inp[10]) ? 4'b1100 : 4'b1010;
													assign node5495 = (inp[4]) ? node5501 : node5496;
														assign node5496 = (inp[10]) ? 4'b1100 : node5497;
															assign node5497 = (inp[3]) ? 4'b1000 : 4'b1010;
														assign node5501 = (inp[10]) ? 4'b1000 : 4'b1100;
							assign node5504 = (inp[14]) ? node6038 : node5505;
								assign node5505 = (inp[2]) ? node5753 : node5506;
									assign node5506 = (inp[9]) ? node5632 : node5507;
										assign node5507 = (inp[4]) ? node5579 : node5508;
											assign node5508 = (inp[10]) ? node5544 : node5509;
												assign node5509 = (inp[5]) ? node5525 : node5510;
													assign node5510 = (inp[3]) ? node5518 : node5511;
														assign node5511 = (inp[15]) ? node5515 : node5512;
															assign node5512 = (inp[0]) ? 4'b1100 : 4'b1110;
															assign node5515 = (inp[0]) ? 4'b1110 : 4'b1100;
														assign node5518 = (inp[15]) ? node5522 : node5519;
															assign node5519 = (inp[0]) ? 4'b1100 : 4'b1110;
															assign node5522 = (inp[0]) ? 4'b1110 : 4'b1100;
													assign node5525 = (inp[15]) ? node5537 : node5526;
														assign node5526 = (inp[12]) ? node5532 : node5527;
															assign node5527 = (inp[3]) ? node5529 : 4'b1100;
																assign node5529 = (inp[0]) ? 4'b1110 : 4'b1100;
															assign node5532 = (inp[3]) ? node5534 : 4'b1110;
																assign node5534 = (inp[0]) ? 4'b1110 : 4'b1100;
														assign node5537 = (inp[12]) ? 4'b1100 : node5538;
															assign node5538 = (inp[0]) ? 4'b1100 : node5539;
																assign node5539 = (inp[3]) ? 4'b1110 : 4'b1100;
												assign node5544 = (inp[12]) ? node5556 : node5545;
													assign node5545 = (inp[15]) ? node5551 : node5546;
														assign node5546 = (inp[0]) ? 4'b1100 : node5547;
															assign node5547 = (inp[5]) ? 4'b1100 : 4'b1110;
														assign node5551 = (inp[0]) ? 4'b1110 : node5552;
															assign node5552 = (inp[3]) ? 4'b1110 : 4'b1100;
													assign node5556 = (inp[5]) ? node5564 : node5557;
														assign node5557 = (inp[15]) ? node5561 : node5558;
															assign node5558 = (inp[0]) ? 4'b1000 : 4'b1010;
															assign node5561 = (inp[0]) ? 4'b1010 : 4'b1000;
														assign node5564 = (inp[3]) ? node5572 : node5565;
															assign node5565 = (inp[15]) ? node5569 : node5566;
																assign node5566 = (inp[0]) ? 4'b1000 : 4'b1010;
																assign node5569 = (inp[0]) ? 4'b1010 : 4'b1000;
															assign node5572 = (inp[15]) ? node5576 : node5573;
																assign node5573 = (inp[0]) ? 4'b1010 : 4'b1000;
																assign node5576 = (inp[0]) ? 4'b1000 : 4'b1010;
											assign node5579 = (inp[12]) ? node5603 : node5580;
												assign node5580 = (inp[0]) ? node5592 : node5581;
													assign node5581 = (inp[15]) ? node5587 : node5582;
														assign node5582 = (inp[3]) ? node5584 : 4'b1010;
															assign node5584 = (inp[5]) ? 4'b1000 : 4'b1010;
														assign node5587 = (inp[3]) ? node5589 : 4'b1000;
															assign node5589 = (inp[5]) ? 4'b1010 : 4'b1000;
													assign node5592 = (inp[15]) ? node5598 : node5593;
														assign node5593 = (inp[3]) ? node5595 : 4'b1000;
															assign node5595 = (inp[5]) ? 4'b1010 : 4'b1000;
														assign node5598 = (inp[3]) ? node5600 : 4'b1010;
															assign node5600 = (inp[5]) ? 4'b1000 : 4'b1010;
												assign node5603 = (inp[10]) ? node5621 : node5604;
													assign node5604 = (inp[15]) ? node5614 : node5605;
														assign node5605 = (inp[3]) ? node5607 : 4'b1000;
															assign node5607 = (inp[5]) ? node5611 : node5608;
																assign node5608 = (inp[0]) ? 4'b1000 : 4'b1010;
																assign node5611 = (inp[0]) ? 4'b1010 : 4'b1000;
														assign node5614 = (inp[0]) ? node5618 : node5615;
															assign node5615 = (inp[3]) ? 4'b1010 : 4'b1000;
															assign node5618 = (inp[3]) ? 4'b1000 : 4'b1010;
													assign node5621 = (inp[15]) ? node5629 : node5622;
														assign node5622 = (inp[0]) ? 4'b1110 : node5623;
															assign node5623 = (inp[3]) ? 4'b1100 : node5624;
																assign node5624 = (inp[5]) ? 4'b1100 : 4'b1110;
														assign node5629 = (inp[0]) ? 4'b1100 : 4'b1110;
										assign node5632 = (inp[4]) ? node5698 : node5633;
											assign node5633 = (inp[10]) ? node5665 : node5634;
												assign node5634 = (inp[3]) ? node5650 : node5635;
													assign node5635 = (inp[5]) ? node5643 : node5636;
														assign node5636 = (inp[0]) ? node5640 : node5637;
															assign node5637 = (inp[15]) ? 4'b1000 : 4'b1010;
															assign node5640 = (inp[15]) ? 4'b1010 : 4'b1000;
														assign node5643 = (inp[15]) ? node5647 : node5644;
															assign node5644 = (inp[0]) ? 4'b1000 : 4'b1010;
															assign node5647 = (inp[0]) ? 4'b1010 : 4'b1000;
													assign node5650 = (inp[12]) ? node5652 : 4'b1010;
														assign node5652 = (inp[5]) ? node5660 : node5653;
															assign node5653 = (inp[0]) ? node5657 : node5654;
																assign node5654 = (inp[15]) ? 4'b1000 : 4'b1010;
																assign node5657 = (inp[15]) ? 4'b1010 : 4'b1000;
															assign node5660 = (inp[15]) ? 4'b1010 : node5661;
																assign node5661 = (inp[0]) ? 4'b1010 : 4'b1000;
												assign node5665 = (inp[12]) ? node5681 : node5666;
													assign node5666 = (inp[5]) ? node5674 : node5667;
														assign node5667 = (inp[0]) ? node5671 : node5668;
															assign node5668 = (inp[15]) ? 4'b1000 : 4'b1010;
															assign node5671 = (inp[15]) ? 4'b1010 : 4'b1000;
														assign node5674 = (inp[3]) ? node5676 : 4'b1000;
															assign node5676 = (inp[15]) ? 4'b1000 : node5677;
																assign node5677 = (inp[0]) ? 4'b1010 : 4'b1000;
													assign node5681 = (inp[3]) ? node5691 : node5682;
														assign node5682 = (inp[0]) ? 4'b1100 : node5683;
															assign node5683 = (inp[15]) ? node5687 : node5684;
																assign node5684 = (inp[5]) ? 4'b1100 : 4'b1110;
																assign node5687 = (inp[5]) ? 4'b1110 : 4'b1100;
														assign node5691 = (inp[15]) ? node5695 : node5692;
															assign node5692 = (inp[0]) ? 4'b1110 : 4'b1100;
															assign node5695 = (inp[0]) ? 4'b1100 : 4'b1110;
											assign node5698 = (inp[12]) ? node5722 : node5699;
												assign node5699 = (inp[0]) ? node5711 : node5700;
													assign node5700 = (inp[15]) ? node5706 : node5701;
														assign node5701 = (inp[3]) ? 4'b1100 : node5702;
															assign node5702 = (inp[5]) ? 4'b1100 : 4'b1110;
														assign node5706 = (inp[3]) ? 4'b1110 : node5707;
															assign node5707 = (inp[5]) ? 4'b1110 : 4'b1100;
													assign node5711 = (inp[15]) ? node5717 : node5712;
														assign node5712 = (inp[5]) ? 4'b1110 : node5713;
															assign node5713 = (inp[3]) ? 4'b1110 : 4'b1100;
														assign node5717 = (inp[5]) ? 4'b1100 : node5718;
															assign node5718 = (inp[3]) ? 4'b1100 : 4'b1110;
												assign node5722 = (inp[10]) ? node5742 : node5723;
													assign node5723 = (inp[0]) ? node5735 : node5724;
														assign node5724 = (inp[15]) ? node5730 : node5725;
															assign node5725 = (inp[3]) ? 4'b1100 : node5726;
																assign node5726 = (inp[5]) ? 4'b1100 : 4'b1110;
															assign node5730 = (inp[3]) ? 4'b1110 : node5731;
																assign node5731 = (inp[5]) ? 4'b1110 : 4'b1100;
														assign node5735 = (inp[15]) ? 4'b1100 : node5736;
															assign node5736 = (inp[5]) ? 4'b1110 : node5737;
																assign node5737 = (inp[3]) ? 4'b1110 : 4'b1100;
													assign node5742 = (inp[5]) ? node5748 : node5743;
														assign node5743 = (inp[15]) ? node5745 : 4'b1000;
															assign node5745 = (inp[3]) ? 4'b1010 : 4'b1000;
														assign node5748 = (inp[15]) ? node5750 : 4'b1010;
															assign node5750 = (inp[0]) ? 4'b1000 : 4'b1010;
									assign node5753 = (inp[10]) ? node5881 : node5754;
										assign node5754 = (inp[3]) ? node5808 : node5755;
											assign node5755 = (inp[4]) ? node5771 : node5756;
												assign node5756 = (inp[9]) ? node5764 : node5757;
													assign node5757 = (inp[0]) ? node5761 : node5758;
														assign node5758 = (inp[15]) ? 4'b0101 : 4'b0111;
														assign node5761 = (inp[15]) ? 4'b0111 : 4'b0101;
													assign node5764 = (inp[15]) ? node5768 : node5765;
														assign node5765 = (inp[0]) ? 4'b0001 : 4'b0011;
														assign node5768 = (inp[0]) ? 4'b0011 : 4'b0001;
												assign node5771 = (inp[9]) ? node5785 : node5772;
													assign node5772 = (inp[12]) ? node5778 : node5773;
														assign node5773 = (inp[5]) ? node5775 : 4'b0001;
															assign node5775 = (inp[15]) ? 4'b0011 : 4'b0001;
														assign node5778 = (inp[0]) ? node5782 : node5779;
															assign node5779 = (inp[15]) ? 4'b0001 : 4'b0011;
															assign node5782 = (inp[15]) ? 4'b0011 : 4'b0001;
													assign node5785 = (inp[5]) ? node5801 : node5786;
														assign node5786 = (inp[12]) ? node5794 : node5787;
															assign node5787 = (inp[0]) ? node5791 : node5788;
																assign node5788 = (inp[15]) ? 4'b0101 : 4'b0111;
																assign node5791 = (inp[15]) ? 4'b0111 : 4'b0101;
															assign node5794 = (inp[0]) ? node5798 : node5795;
																assign node5795 = (inp[15]) ? 4'b0101 : 4'b0111;
																assign node5798 = (inp[15]) ? 4'b0111 : 4'b0101;
														assign node5801 = (inp[0]) ? node5805 : node5802;
															assign node5802 = (inp[15]) ? 4'b0111 : 4'b0101;
															assign node5805 = (inp[15]) ? 4'b0101 : 4'b0111;
											assign node5808 = (inp[15]) ? node5842 : node5809;
												assign node5809 = (inp[0]) ? node5825 : node5810;
													assign node5810 = (inp[5]) ? node5818 : node5811;
														assign node5811 = (inp[9]) ? node5815 : node5812;
															assign node5812 = (inp[4]) ? 4'b0011 : 4'b0111;
															assign node5815 = (inp[4]) ? 4'b0101 : 4'b0011;
														assign node5818 = (inp[4]) ? node5822 : node5819;
															assign node5819 = (inp[9]) ? 4'b0001 : 4'b0101;
															assign node5822 = (inp[9]) ? 4'b0101 : 4'b0001;
													assign node5825 = (inp[5]) ? node5833 : node5826;
														assign node5826 = (inp[9]) ? node5830 : node5827;
															assign node5827 = (inp[4]) ? 4'b0001 : 4'b0101;
															assign node5830 = (inp[4]) ? 4'b0111 : 4'b0001;
														assign node5833 = (inp[12]) ? 4'b0011 : node5834;
															assign node5834 = (inp[4]) ? node5838 : node5835;
																assign node5835 = (inp[9]) ? 4'b0011 : 4'b0111;
																assign node5838 = (inp[9]) ? 4'b0111 : 4'b0011;
												assign node5842 = (inp[12]) ? node5860 : node5843;
													assign node5843 = (inp[4]) ? node5857 : node5844;
														assign node5844 = (inp[9]) ? node5852 : node5845;
															assign node5845 = (inp[0]) ? node5849 : node5846;
																assign node5846 = (inp[5]) ? 4'b0111 : 4'b0101;
																assign node5849 = (inp[5]) ? 4'b0101 : 4'b0111;
															assign node5852 = (inp[5]) ? 4'b0001 : node5853;
																assign node5853 = (inp[0]) ? 4'b0011 : 4'b0001;
														assign node5857 = (inp[9]) ? 4'b0101 : 4'b0001;
													assign node5860 = (inp[4]) ? node5874 : node5861;
														assign node5861 = (inp[9]) ? node5867 : node5862;
															assign node5862 = (inp[0]) ? node5864 : 4'b0101;
																assign node5864 = (inp[5]) ? 4'b0101 : 4'b0111;
															assign node5867 = (inp[0]) ? node5871 : node5868;
																assign node5868 = (inp[5]) ? 4'b0011 : 4'b0001;
																assign node5871 = (inp[5]) ? 4'b0001 : 4'b0011;
														assign node5874 = (inp[9]) ? node5878 : node5875;
															assign node5875 = (inp[0]) ? 4'b0011 : 4'b0001;
															assign node5878 = (inp[0]) ? 4'b0101 : 4'b0111;
										assign node5881 = (inp[12]) ? node5947 : node5882;
											assign node5882 = (inp[0]) ? node5914 : node5883;
												assign node5883 = (inp[15]) ? node5897 : node5884;
													assign node5884 = (inp[5]) ? node5890 : node5885;
														assign node5885 = (inp[4]) ? 4'b0011 : node5886;
															assign node5886 = (inp[9]) ? 4'b0011 : 4'b0111;
														assign node5890 = (inp[4]) ? node5892 : 4'b0011;
															assign node5892 = (inp[9]) ? 4'b0101 : node5893;
																assign node5893 = (inp[3]) ? 4'b0001 : 4'b0011;
													assign node5897 = (inp[5]) ? node5903 : node5898;
														assign node5898 = (inp[9]) ? 4'b0001 : node5899;
															assign node5899 = (inp[4]) ? 4'b0001 : 4'b0101;
														assign node5903 = (inp[3]) ? node5909 : node5904;
															assign node5904 = (inp[9]) ? 4'b0111 : node5905;
																assign node5905 = (inp[4]) ? 4'b0001 : 4'b0101;
															assign node5909 = (inp[9]) ? node5911 : 4'b0011;
																assign node5911 = (inp[4]) ? 4'b0111 : 4'b0011;
												assign node5914 = (inp[15]) ? node5934 : node5915;
													assign node5915 = (inp[3]) ? node5923 : node5916;
														assign node5916 = (inp[9]) ? node5920 : node5917;
															assign node5917 = (inp[4]) ? 4'b0001 : 4'b0101;
															assign node5920 = (inp[4]) ? 4'b0101 : 4'b0001;
														assign node5923 = (inp[5]) ? node5929 : node5924;
															assign node5924 = (inp[4]) ? node5926 : 4'b0001;
																assign node5926 = (inp[9]) ? 4'b0111 : 4'b0001;
															assign node5929 = (inp[9]) ? 4'b0111 : node5930;
																assign node5930 = (inp[4]) ? 4'b0011 : 4'b0111;
													assign node5934 = (inp[3]) ? node5942 : node5935;
														assign node5935 = (inp[4]) ? node5939 : node5936;
															assign node5936 = (inp[9]) ? 4'b0011 : 4'b0111;
															assign node5939 = (inp[9]) ? 4'b0111 : 4'b0011;
														assign node5942 = (inp[4]) ? node5944 : 4'b0011;
															assign node5944 = (inp[9]) ? 4'b0101 : 4'b0001;
											assign node5947 = (inp[5]) ? node5999 : node5948;
												assign node5948 = (inp[15]) ? node5968 : node5949;
													assign node5949 = (inp[3]) ? node5955 : node5950;
														assign node5950 = (inp[4]) ? node5952 : 4'b0011;
															assign node5952 = (inp[9]) ? 4'b0011 : 4'b0111;
														assign node5955 = (inp[0]) ? node5961 : node5956;
															assign node5956 = (inp[9]) ? node5958 : 4'b0011;
																assign node5958 = (inp[4]) ? 4'b0001 : 4'b0101;
															assign node5961 = (inp[4]) ? node5965 : node5962;
																assign node5962 = (inp[9]) ? 4'b0111 : 4'b0001;
																assign node5965 = (inp[9]) ? 4'b0011 : 4'b0111;
													assign node5968 = (inp[0]) ? node5984 : node5969;
														assign node5969 = (inp[3]) ? node5977 : node5970;
															assign node5970 = (inp[9]) ? node5974 : node5971;
																assign node5971 = (inp[4]) ? 4'b0101 : 4'b0001;
																assign node5974 = (inp[4]) ? 4'b0001 : 4'b0101;
															assign node5977 = (inp[9]) ? node5981 : node5978;
																assign node5978 = (inp[4]) ? 4'b0111 : 4'b0001;
																assign node5981 = (inp[4]) ? 4'b0011 : 4'b0111;
														assign node5984 = (inp[3]) ? node5992 : node5985;
															assign node5985 = (inp[9]) ? node5989 : node5986;
																assign node5986 = (inp[4]) ? 4'b0111 : 4'b0011;
																assign node5989 = (inp[4]) ? 4'b0011 : 4'b0111;
															assign node5992 = (inp[9]) ? node5996 : node5993;
																assign node5993 = (inp[4]) ? 4'b0101 : 4'b0011;
																assign node5996 = (inp[4]) ? 4'b0001 : 4'b0101;
												assign node5999 = (inp[0]) ? node6021 : node6000;
													assign node6000 = (inp[15]) ? node6008 : node6001;
														assign node6001 = (inp[9]) ? node6005 : node6002;
															assign node6002 = (inp[4]) ? 4'b0101 : 4'b0011;
															assign node6005 = (inp[4]) ? 4'b0001 : 4'b0101;
														assign node6008 = (inp[3]) ? node6014 : node6009;
															assign node6009 = (inp[4]) ? 4'b0111 : node6010;
																assign node6010 = (inp[9]) ? 4'b0111 : 4'b0001;
															assign node6014 = (inp[4]) ? node6018 : node6015;
																assign node6015 = (inp[9]) ? 4'b0111 : 4'b0011;
																assign node6018 = (inp[9]) ? 4'b0011 : 4'b0111;
													assign node6021 = (inp[15]) ? node6029 : node6022;
														assign node6022 = (inp[9]) ? node6026 : node6023;
															assign node6023 = (inp[4]) ? 4'b0111 : 4'b0001;
															assign node6026 = (inp[4]) ? 4'b0011 : 4'b0111;
														assign node6029 = (inp[4]) ? node6035 : node6030;
															assign node6030 = (inp[3]) ? node6032 : 4'b0011;
																assign node6032 = (inp[9]) ? 4'b0101 : 4'b0001;
															assign node6035 = (inp[9]) ? 4'b0001 : 4'b0101;
								assign node6038 = (inp[0]) ? node6250 : node6039;
									assign node6039 = (inp[15]) ? node6147 : node6040;
										assign node6040 = (inp[3]) ? node6100 : node6041;
											assign node6041 = (inp[5]) ? node6077 : node6042;
												assign node6042 = (inp[2]) ? node6062 : node6043;
													assign node6043 = (inp[12]) ? node6057 : node6044;
														assign node6044 = (inp[10]) ? node6050 : node6045;
															assign node6045 = (inp[4]) ? node6047 : 4'b0011;
																assign node6047 = (inp[9]) ? 4'b0111 : 4'b0011;
															assign node6050 = (inp[9]) ? node6054 : node6051;
																assign node6051 = (inp[4]) ? 4'b0011 : 4'b0111;
																assign node6054 = (inp[4]) ? 4'b0111 : 4'b0011;
														assign node6057 = (inp[10]) ? 4'b0111 : node6058;
															assign node6058 = (inp[9]) ? 4'b0111 : 4'b0011;
													assign node6062 = (inp[10]) ? node6068 : node6063;
														assign node6063 = (inp[4]) ? 4'b0111 : node6064;
															assign node6064 = (inp[9]) ? 4'b0011 : 4'b0111;
														assign node6068 = (inp[4]) ? node6070 : 4'b0111;
															assign node6070 = (inp[9]) ? node6074 : node6071;
																assign node6071 = (inp[12]) ? 4'b0111 : 4'b0011;
																assign node6074 = (inp[12]) ? 4'b0011 : 4'b0111;
												assign node6077 = (inp[9]) ? node6089 : node6078;
													assign node6078 = (inp[4]) ? node6084 : node6079;
														assign node6079 = (inp[10]) ? node6081 : 4'b0111;
															assign node6081 = (inp[12]) ? 4'b0011 : 4'b0111;
														assign node6084 = (inp[12]) ? node6086 : 4'b0011;
															assign node6086 = (inp[10]) ? 4'b0101 : 4'b0011;
													assign node6089 = (inp[4]) ? node6095 : node6090;
														assign node6090 = (inp[12]) ? node6092 : 4'b0011;
															assign node6092 = (inp[10]) ? 4'b0101 : 4'b0011;
														assign node6095 = (inp[12]) ? node6097 : 4'b0101;
															assign node6097 = (inp[10]) ? 4'b0001 : 4'b0101;
											assign node6100 = (inp[5]) ? node6124 : node6101;
												assign node6101 = (inp[9]) ? node6113 : node6102;
													assign node6102 = (inp[4]) ? node6108 : node6103;
														assign node6103 = (inp[10]) ? node6105 : 4'b0111;
															assign node6105 = (inp[12]) ? 4'b0011 : 4'b0111;
														assign node6108 = (inp[12]) ? node6110 : 4'b0011;
															assign node6110 = (inp[10]) ? 4'b0101 : 4'b0011;
													assign node6113 = (inp[4]) ? node6119 : node6114;
														assign node6114 = (inp[12]) ? node6116 : 4'b0011;
															assign node6116 = (inp[10]) ? 4'b0101 : 4'b0011;
														assign node6119 = (inp[12]) ? node6121 : 4'b0101;
															assign node6121 = (inp[10]) ? 4'b0001 : 4'b0101;
												assign node6124 = (inp[4]) ? node6136 : node6125;
													assign node6125 = (inp[9]) ? node6133 : node6126;
														assign node6126 = (inp[2]) ? node6128 : 4'b0101;
															assign node6128 = (inp[12]) ? node6130 : 4'b0101;
																assign node6130 = (inp[10]) ? 4'b0001 : 4'b0101;
														assign node6133 = (inp[10]) ? 4'b0101 : 4'b0001;
													assign node6136 = (inp[9]) ? node6142 : node6137;
														assign node6137 = (inp[12]) ? node6139 : 4'b0001;
															assign node6139 = (inp[10]) ? 4'b0101 : 4'b0001;
														assign node6142 = (inp[10]) ? node6144 : 4'b0101;
															assign node6144 = (inp[12]) ? 4'b0001 : 4'b0101;
										assign node6147 = (inp[3]) ? node6207 : node6148;
											assign node6148 = (inp[5]) ? node6184 : node6149;
												assign node6149 = (inp[10]) ? node6163 : node6150;
													assign node6150 = (inp[2]) ? node6156 : node6151;
														assign node6151 = (inp[4]) ? node6153 : 4'b0101;
															assign node6153 = (inp[9]) ? 4'b0101 : 4'b0001;
														assign node6156 = (inp[9]) ? node6160 : node6157;
															assign node6157 = (inp[4]) ? 4'b0001 : 4'b0101;
															assign node6160 = (inp[4]) ? 4'b0101 : 4'b0001;
													assign node6163 = (inp[2]) ? node6169 : node6164;
														assign node6164 = (inp[12]) ? node6166 : 4'b0001;
															assign node6166 = (inp[9]) ? 4'b0101 : 4'b0001;
														assign node6169 = (inp[9]) ? node6177 : node6170;
															assign node6170 = (inp[4]) ? node6174 : node6171;
																assign node6171 = (inp[12]) ? 4'b0001 : 4'b0101;
																assign node6174 = (inp[12]) ? 4'b0101 : 4'b0001;
															assign node6177 = (inp[4]) ? node6181 : node6178;
																assign node6178 = (inp[12]) ? 4'b0101 : 4'b0001;
																assign node6181 = (inp[12]) ? 4'b0001 : 4'b0101;
												assign node6184 = (inp[4]) ? node6196 : node6185;
													assign node6185 = (inp[9]) ? node6191 : node6186;
														assign node6186 = (inp[10]) ? node6188 : 4'b0101;
															assign node6188 = (inp[12]) ? 4'b0001 : 4'b0101;
														assign node6191 = (inp[10]) ? node6193 : 4'b0001;
															assign node6193 = (inp[12]) ? 4'b0111 : 4'b0001;
													assign node6196 = (inp[9]) ? node6202 : node6197;
														assign node6197 = (inp[10]) ? node6199 : 4'b0001;
															assign node6199 = (inp[12]) ? 4'b0111 : 4'b0001;
														assign node6202 = (inp[12]) ? node6204 : 4'b0111;
															assign node6204 = (inp[10]) ? 4'b0011 : 4'b0111;
											assign node6207 = (inp[5]) ? node6233 : node6208;
												assign node6208 = (inp[9]) ? node6222 : node6209;
													assign node6209 = (inp[4]) ? node6215 : node6210;
														assign node6210 = (inp[12]) ? node6212 : 4'b0101;
															assign node6212 = (inp[10]) ? 4'b0001 : 4'b0101;
														assign node6215 = (inp[2]) ? 4'b0001 : node6216;
															assign node6216 = (inp[12]) ? node6218 : 4'b0001;
																assign node6218 = (inp[10]) ? 4'b0111 : 4'b0001;
													assign node6222 = (inp[4]) ? node6228 : node6223;
														assign node6223 = (inp[10]) ? node6225 : 4'b0001;
															assign node6225 = (inp[12]) ? 4'b0111 : 4'b0001;
														assign node6228 = (inp[10]) ? node6230 : 4'b0111;
															assign node6230 = (inp[12]) ? 4'b0011 : 4'b0111;
												assign node6233 = (inp[12]) ? node6241 : node6234;
													assign node6234 = (inp[4]) ? node6238 : node6235;
														assign node6235 = (inp[9]) ? 4'b0011 : 4'b0111;
														assign node6238 = (inp[9]) ? 4'b0111 : 4'b0011;
													assign node6241 = (inp[4]) ? 4'b0111 : node6242;
														assign node6242 = (inp[10]) ? node6246 : node6243;
															assign node6243 = (inp[9]) ? 4'b0011 : 4'b0111;
															assign node6246 = (inp[9]) ? 4'b0111 : 4'b0011;
									assign node6250 = (inp[15]) ? node6372 : node6251;
										assign node6251 = (inp[5]) ? node6301 : node6252;
											assign node6252 = (inp[3]) ? node6280 : node6253;
												assign node6253 = (inp[10]) ? node6261 : node6254;
													assign node6254 = (inp[9]) ? node6258 : node6255;
														assign node6255 = (inp[4]) ? 4'b0001 : 4'b0101;
														assign node6258 = (inp[4]) ? 4'b0101 : 4'b0001;
													assign node6261 = (inp[12]) ? node6269 : node6262;
														assign node6262 = (inp[4]) ? node6266 : node6263;
															assign node6263 = (inp[9]) ? 4'b0001 : 4'b0101;
															assign node6266 = (inp[9]) ? 4'b0101 : 4'b0001;
														assign node6269 = (inp[2]) ? node6275 : node6270;
															assign node6270 = (inp[4]) ? 4'b0101 : node6271;
																assign node6271 = (inp[9]) ? 4'b0101 : 4'b0001;
															assign node6275 = (inp[9]) ? node6277 : 4'b0101;
																assign node6277 = (inp[4]) ? 4'b0001 : 4'b0101;
												assign node6280 = (inp[4]) ? node6290 : node6281;
													assign node6281 = (inp[9]) ? node6285 : node6282;
														assign node6282 = (inp[12]) ? 4'b0001 : 4'b0101;
														assign node6285 = (inp[12]) ? node6287 : 4'b0001;
															assign node6287 = (inp[10]) ? 4'b0111 : 4'b0001;
													assign node6290 = (inp[9]) ? node6296 : node6291;
														assign node6291 = (inp[12]) ? node6293 : 4'b0001;
															assign node6293 = (inp[10]) ? 4'b0111 : 4'b0001;
														assign node6296 = (inp[10]) ? node6298 : 4'b0111;
															assign node6298 = (inp[12]) ? 4'b0011 : 4'b0111;
											assign node6301 = (inp[3]) ? node6329 : node6302;
												assign node6302 = (inp[4]) ? node6314 : node6303;
													assign node6303 = (inp[9]) ? node6309 : node6304;
														assign node6304 = (inp[10]) ? node6306 : 4'b0101;
															assign node6306 = (inp[12]) ? 4'b0001 : 4'b0101;
														assign node6309 = (inp[12]) ? node6311 : 4'b0001;
															assign node6311 = (inp[10]) ? 4'b0111 : 4'b0001;
													assign node6314 = (inp[2]) ? node6322 : node6315;
														assign node6315 = (inp[9]) ? node6319 : node6316;
															assign node6316 = (inp[10]) ? 4'b0111 : 4'b0001;
															assign node6319 = (inp[12]) ? 4'b0011 : 4'b0111;
														assign node6322 = (inp[10]) ? node6324 : 4'b0111;
															assign node6324 = (inp[9]) ? node6326 : 4'b0111;
																assign node6326 = (inp[12]) ? 4'b0011 : 4'b0111;
												assign node6329 = (inp[2]) ? node6353 : node6330;
													assign node6330 = (inp[10]) ? node6338 : node6331;
														assign node6331 = (inp[9]) ? node6335 : node6332;
															assign node6332 = (inp[4]) ? 4'b0011 : 4'b0111;
															assign node6335 = (inp[4]) ? 4'b0111 : 4'b0011;
														assign node6338 = (inp[12]) ? node6346 : node6339;
															assign node6339 = (inp[9]) ? node6343 : node6340;
																assign node6340 = (inp[4]) ? 4'b0011 : 4'b0111;
																assign node6343 = (inp[4]) ? 4'b0111 : 4'b0011;
															assign node6346 = (inp[4]) ? node6350 : node6347;
																assign node6347 = (inp[9]) ? 4'b0111 : 4'b0011;
																assign node6350 = (inp[9]) ? 4'b0011 : 4'b0111;
													assign node6353 = (inp[9]) ? node6363 : node6354;
														assign node6354 = (inp[4]) ? node6358 : node6355;
															assign node6355 = (inp[10]) ? 4'b0011 : 4'b0111;
															assign node6358 = (inp[10]) ? node6360 : 4'b0011;
																assign node6360 = (inp[12]) ? 4'b0111 : 4'b0011;
														assign node6363 = (inp[10]) ? node6365 : 4'b0011;
															assign node6365 = (inp[12]) ? node6369 : node6366;
																assign node6366 = (inp[4]) ? 4'b0111 : 4'b0011;
																assign node6369 = (inp[4]) ? 4'b0011 : 4'b0111;
										assign node6372 = (inp[5]) ? node6422 : node6373;
											assign node6373 = (inp[3]) ? node6397 : node6374;
												assign node6374 = (inp[12]) ? node6382 : node6375;
													assign node6375 = (inp[9]) ? node6379 : node6376;
														assign node6376 = (inp[4]) ? 4'b0011 : 4'b0111;
														assign node6379 = (inp[4]) ? 4'b0111 : 4'b0011;
													assign node6382 = (inp[4]) ? node6392 : node6383;
														assign node6383 = (inp[2]) ? 4'b0111 : node6384;
															assign node6384 = (inp[9]) ? node6388 : node6385;
																assign node6385 = (inp[10]) ? 4'b0011 : 4'b0111;
																assign node6388 = (inp[10]) ? 4'b0111 : 4'b0011;
														assign node6392 = (inp[10]) ? 4'b0011 : node6393;
															assign node6393 = (inp[9]) ? 4'b0111 : 4'b0011;
												assign node6397 = (inp[9]) ? node6409 : node6398;
													assign node6398 = (inp[4]) ? node6404 : node6399;
														assign node6399 = (inp[10]) ? node6401 : 4'b0111;
															assign node6401 = (inp[12]) ? 4'b0011 : 4'b0111;
														assign node6404 = (inp[12]) ? node6406 : 4'b0011;
															assign node6406 = (inp[10]) ? 4'b0101 : 4'b0011;
													assign node6409 = (inp[4]) ? node6415 : node6410;
														assign node6410 = (inp[12]) ? node6412 : 4'b0011;
															assign node6412 = (inp[10]) ? 4'b0101 : 4'b0011;
														assign node6415 = (inp[2]) ? 4'b0101 : node6416;
															assign node6416 = (inp[12]) ? node6418 : 4'b0101;
																assign node6418 = (inp[10]) ? 4'b0001 : 4'b0101;
											assign node6422 = (inp[3]) ? node6442 : node6423;
												assign node6423 = (inp[4]) ? node6435 : node6424;
													assign node6424 = (inp[9]) ? node6430 : node6425;
														assign node6425 = (inp[12]) ? node6427 : 4'b0111;
															assign node6427 = (inp[10]) ? 4'b0011 : 4'b0111;
														assign node6430 = (inp[10]) ? node6432 : 4'b0011;
															assign node6432 = (inp[12]) ? 4'b0101 : 4'b0011;
													assign node6435 = (inp[9]) ? node6437 : 4'b0011;
														assign node6437 = (inp[12]) ? node6439 : 4'b0101;
															assign node6439 = (inp[10]) ? 4'b0001 : 4'b0101;
												assign node6442 = (inp[10]) ? node6460 : node6443;
													assign node6443 = (inp[2]) ? node6451 : node6444;
														assign node6444 = (inp[9]) ? node6448 : node6445;
															assign node6445 = (inp[4]) ? 4'b0001 : 4'b0101;
															assign node6448 = (inp[4]) ? 4'b0101 : 4'b0001;
														assign node6451 = (inp[12]) ? node6455 : node6452;
															assign node6452 = (inp[9]) ? 4'b0101 : 4'b0001;
															assign node6455 = (inp[9]) ? 4'b0001 : node6456;
																assign node6456 = (inp[4]) ? 4'b0001 : 4'b0101;
													assign node6460 = (inp[2]) ? node6466 : node6461;
														assign node6461 = (inp[4]) ? 4'b0101 : node6462;
															assign node6462 = (inp[12]) ? 4'b0101 : 4'b0001;
														assign node6466 = (inp[12]) ? node6474 : node6467;
															assign node6467 = (inp[9]) ? node6471 : node6468;
																assign node6468 = (inp[4]) ? 4'b0001 : 4'b0101;
																assign node6471 = (inp[4]) ? 4'b0101 : 4'b0001;
															assign node6474 = (inp[4]) ? node6478 : node6475;
																assign node6475 = (inp[9]) ? 4'b0101 : 4'b0001;
																assign node6478 = (inp[9]) ? 4'b0001 : 4'b0101;
						assign node6481 = (inp[7]) ? node7595 : node6482;
							assign node6482 = (inp[14]) ? node7040 : node6483;
								assign node6483 = (inp[2]) ? node6793 : node6484;
									assign node6484 = (inp[12]) ? node6614 : node6485;
										assign node6485 = (inp[4]) ? node6549 : node6486;
											assign node6486 = (inp[9]) ? node6512 : node6487;
												assign node6487 = (inp[3]) ? node6495 : node6488;
													assign node6488 = (inp[15]) ? node6492 : node6489;
														assign node6489 = (inp[0]) ? 4'b1100 : 4'b1110;
														assign node6492 = (inp[0]) ? 4'b1110 : 4'b1100;
													assign node6495 = (inp[5]) ? node6505 : node6496;
														assign node6496 = (inp[10]) ? node6500 : node6497;
															assign node6497 = (inp[15]) ? 4'b1110 : 4'b1100;
															assign node6500 = (inp[15]) ? 4'b1100 : node6501;
																assign node6501 = (inp[0]) ? 4'b1100 : 4'b1110;
														assign node6505 = (inp[15]) ? node6509 : node6506;
															assign node6506 = (inp[0]) ? 4'b1110 : 4'b1100;
															assign node6509 = (inp[0]) ? 4'b1100 : 4'b1110;
												assign node6512 = (inp[10]) ? node6528 : node6513;
													assign node6513 = (inp[15]) ? node6519 : node6514;
														assign node6514 = (inp[0]) ? 4'b1000 : node6515;
															assign node6515 = (inp[3]) ? 4'b1000 : 4'b1010;
														assign node6519 = (inp[5]) ? node6523 : node6520;
															assign node6520 = (inp[0]) ? 4'b1010 : 4'b1000;
															assign node6523 = (inp[0]) ? 4'b1000 : node6524;
																assign node6524 = (inp[3]) ? 4'b1010 : 4'b1000;
													assign node6528 = (inp[5]) ? node6534 : node6529;
														assign node6529 = (inp[0]) ? node6531 : 4'b1010;
															assign node6531 = (inp[15]) ? 4'b1010 : 4'b1000;
														assign node6534 = (inp[0]) ? node6542 : node6535;
															assign node6535 = (inp[3]) ? node6539 : node6536;
																assign node6536 = (inp[15]) ? 4'b1000 : 4'b1010;
																assign node6539 = (inp[15]) ? 4'b1010 : 4'b1000;
															assign node6542 = (inp[15]) ? node6546 : node6543;
																assign node6543 = (inp[3]) ? 4'b1010 : 4'b1000;
																assign node6546 = (inp[3]) ? 4'b1000 : 4'b1010;
											assign node6549 = (inp[9]) ? node6591 : node6550;
												assign node6550 = (inp[10]) ? node6574 : node6551;
													assign node6551 = (inp[5]) ? node6559 : node6552;
														assign node6552 = (inp[15]) ? node6556 : node6553;
															assign node6553 = (inp[0]) ? 4'b1000 : 4'b1010;
															assign node6556 = (inp[0]) ? 4'b1010 : 4'b1000;
														assign node6559 = (inp[3]) ? node6567 : node6560;
															assign node6560 = (inp[15]) ? node6564 : node6561;
																assign node6561 = (inp[0]) ? 4'b1000 : 4'b1010;
																assign node6564 = (inp[0]) ? 4'b1010 : 4'b1000;
															assign node6567 = (inp[15]) ? node6571 : node6568;
																assign node6568 = (inp[0]) ? 4'b1010 : 4'b1000;
																assign node6571 = (inp[0]) ? 4'b1000 : 4'b1010;
													assign node6574 = (inp[0]) ? node6580 : node6575;
														assign node6575 = (inp[5]) ? 4'b1000 : node6576;
															assign node6576 = (inp[3]) ? 4'b1010 : 4'b1000;
														assign node6580 = (inp[15]) ? node6586 : node6581;
															assign node6581 = (inp[5]) ? node6583 : 4'b1000;
																assign node6583 = (inp[3]) ? 4'b1010 : 4'b1000;
															assign node6586 = (inp[3]) ? node6588 : 4'b1010;
																assign node6588 = (inp[5]) ? 4'b1000 : 4'b1010;
												assign node6591 = (inp[3]) ? node6607 : node6592;
													assign node6592 = (inp[15]) ? node6600 : node6593;
														assign node6593 = (inp[5]) ? node6597 : node6594;
															assign node6594 = (inp[0]) ? 4'b1100 : 4'b1110;
															assign node6597 = (inp[0]) ? 4'b1110 : 4'b1100;
														assign node6600 = (inp[0]) ? node6604 : node6601;
															assign node6601 = (inp[5]) ? 4'b1110 : 4'b1100;
															assign node6604 = (inp[5]) ? 4'b1100 : 4'b1110;
													assign node6607 = (inp[0]) ? node6611 : node6608;
														assign node6608 = (inp[15]) ? 4'b1110 : 4'b1100;
														assign node6611 = (inp[15]) ? 4'b1100 : 4'b1110;
										assign node6614 = (inp[15]) ? node6700 : node6615;
											assign node6615 = (inp[4]) ? node6657 : node6616;
												assign node6616 = (inp[5]) ? node6626 : node6617;
													assign node6617 = (inp[0]) ? node6619 : 4'b1110;
														assign node6619 = (inp[10]) ? node6623 : node6620;
															assign node6620 = (inp[9]) ? 4'b1000 : 4'b1100;
															assign node6623 = (inp[9]) ? 4'b1100 : 4'b1000;
													assign node6626 = (inp[0]) ? node6642 : node6627;
														assign node6627 = (inp[3]) ? node6635 : node6628;
															assign node6628 = (inp[10]) ? node6632 : node6629;
																assign node6629 = (inp[9]) ? 4'b1010 : 4'b1110;
																assign node6632 = (inp[9]) ? 4'b1100 : 4'b1010;
															assign node6635 = (inp[10]) ? node6639 : node6636;
																assign node6636 = (inp[9]) ? 4'b1000 : 4'b1100;
																assign node6639 = (inp[9]) ? 4'b1100 : 4'b1000;
														assign node6642 = (inp[3]) ? node6650 : node6643;
															assign node6643 = (inp[10]) ? node6647 : node6644;
																assign node6644 = (inp[9]) ? 4'b1000 : 4'b1100;
																assign node6647 = (inp[9]) ? 4'b1110 : 4'b1000;
															assign node6650 = (inp[9]) ? node6654 : node6651;
																assign node6651 = (inp[10]) ? 4'b1010 : 4'b1110;
																assign node6654 = (inp[10]) ? 4'b1110 : 4'b1010;
												assign node6657 = (inp[0]) ? node6675 : node6658;
													assign node6658 = (inp[5]) ? node6670 : node6659;
														assign node6659 = (inp[3]) ? node6665 : node6660;
															assign node6660 = (inp[9]) ? 4'b1110 : node6661;
																assign node6661 = (inp[10]) ? 4'b1110 : 4'b1010;
															assign node6665 = (inp[9]) ? node6667 : 4'b1010;
																assign node6667 = (inp[10]) ? 4'b1000 : 4'b1100;
														assign node6670 = (inp[10]) ? 4'b1100 : node6671;
															assign node6671 = (inp[9]) ? 4'b1100 : 4'b1000;
													assign node6675 = (inp[3]) ? node6687 : node6676;
														assign node6676 = (inp[5]) ? node6682 : node6677;
															assign node6677 = (inp[10]) ? node6679 : 4'b1100;
																assign node6679 = (inp[9]) ? 4'b1000 : 4'b1100;
															assign node6682 = (inp[9]) ? 4'b1110 : node6683;
																assign node6683 = (inp[10]) ? 4'b1110 : 4'b1000;
														assign node6687 = (inp[5]) ? node6693 : node6688;
															assign node6688 = (inp[10]) ? node6690 : 4'b1110;
																assign node6690 = (inp[9]) ? 4'b1010 : 4'b1110;
															assign node6693 = (inp[10]) ? node6697 : node6694;
																assign node6694 = (inp[9]) ? 4'b1110 : 4'b1010;
																assign node6697 = (inp[9]) ? 4'b1010 : 4'b1110;
											assign node6700 = (inp[3]) ? node6744 : node6701;
												assign node6701 = (inp[0]) ? node6729 : node6702;
													assign node6702 = (inp[5]) ? node6716 : node6703;
														assign node6703 = (inp[9]) ? node6709 : node6704;
															assign node6704 = (inp[10]) ? node6706 : 4'b1000;
																assign node6706 = (inp[4]) ? 4'b1100 : 4'b1000;
															assign node6709 = (inp[4]) ? node6713 : node6710;
																assign node6710 = (inp[10]) ? 4'b1100 : 4'b1000;
																assign node6713 = (inp[10]) ? 4'b1000 : 4'b1100;
														assign node6716 = (inp[9]) ? node6724 : node6717;
															assign node6717 = (inp[4]) ? node6721 : node6718;
																assign node6718 = (inp[10]) ? 4'b1000 : 4'b1100;
																assign node6721 = (inp[10]) ? 4'b1110 : 4'b1000;
															assign node6724 = (inp[4]) ? node6726 : 4'b1110;
																assign node6726 = (inp[10]) ? 4'b1010 : 4'b1110;
													assign node6729 = (inp[9]) ? node6737 : node6730;
														assign node6730 = (inp[4]) ? node6734 : node6731;
															assign node6731 = (inp[10]) ? 4'b1010 : 4'b1110;
															assign node6734 = (inp[10]) ? 4'b1110 : 4'b1010;
														assign node6737 = (inp[5]) ? node6739 : 4'b1010;
															assign node6739 = (inp[10]) ? node6741 : 4'b1010;
																assign node6741 = (inp[4]) ? 4'b1000 : 4'b1100;
												assign node6744 = (inp[0]) ? node6772 : node6745;
													assign node6745 = (inp[5]) ? node6757 : node6746;
														assign node6746 = (inp[10]) ? node6752 : node6747;
															assign node6747 = (inp[9]) ? node6749 : 4'b1000;
																assign node6749 = (inp[4]) ? 4'b1110 : 4'b1000;
															assign node6752 = (inp[9]) ? 4'b1110 : node6753;
																assign node6753 = (inp[4]) ? 4'b1110 : 4'b1000;
														assign node6757 = (inp[10]) ? node6765 : node6758;
															assign node6758 = (inp[4]) ? node6762 : node6759;
																assign node6759 = (inp[9]) ? 4'b1010 : 4'b1110;
																assign node6762 = (inp[9]) ? 4'b1110 : 4'b1010;
															assign node6765 = (inp[9]) ? node6769 : node6766;
																assign node6766 = (inp[4]) ? 4'b1110 : 4'b1010;
																assign node6769 = (inp[4]) ? 4'b1010 : 4'b1110;
													assign node6772 = (inp[5]) ? node6782 : node6773;
														assign node6773 = (inp[9]) ? 4'b1100 : node6774;
															assign node6774 = (inp[4]) ? node6778 : node6775;
																assign node6775 = (inp[10]) ? 4'b1010 : 4'b1110;
																assign node6778 = (inp[10]) ? 4'b1100 : 4'b1010;
														assign node6782 = (inp[10]) ? node6788 : node6783;
															assign node6783 = (inp[4]) ? 4'b1000 : node6784;
																assign node6784 = (inp[9]) ? 4'b1000 : 4'b1100;
															assign node6788 = (inp[9]) ? 4'b1100 : node6789;
																assign node6789 = (inp[4]) ? 4'b1100 : 4'b1000;
									assign node6793 = (inp[9]) ? node6925 : node6794;
										assign node6794 = (inp[4]) ? node6858 : node6795;
											assign node6795 = (inp[10]) ? node6817 : node6796;
												assign node6796 = (inp[15]) ? node6806 : node6797;
													assign node6797 = (inp[0]) ? node6801 : node6798;
														assign node6798 = (inp[3]) ? 4'b0101 : 4'b0111;
														assign node6801 = (inp[3]) ? node6803 : 4'b0101;
															assign node6803 = (inp[5]) ? 4'b0111 : 4'b0101;
													assign node6806 = (inp[0]) ? node6812 : node6807;
														assign node6807 = (inp[5]) ? node6809 : 4'b0101;
															assign node6809 = (inp[3]) ? 4'b0111 : 4'b0101;
														assign node6812 = (inp[3]) ? node6814 : 4'b0111;
															assign node6814 = (inp[5]) ? 4'b0101 : 4'b0111;
												assign node6817 = (inp[12]) ? node6837 : node6818;
													assign node6818 = (inp[3]) ? node6828 : node6819;
														assign node6819 = (inp[5]) ? node6825 : node6820;
															assign node6820 = (inp[15]) ? node6822 : 4'b0111;
																assign node6822 = (inp[0]) ? 4'b0111 : 4'b0101;
															assign node6825 = (inp[15]) ? 4'b0111 : 4'b0101;
														assign node6828 = (inp[5]) ? node6830 : 4'b0101;
															assign node6830 = (inp[15]) ? node6834 : node6831;
																assign node6831 = (inp[0]) ? 4'b0111 : 4'b0101;
																assign node6834 = (inp[0]) ? 4'b0101 : 4'b0111;
													assign node6837 = (inp[3]) ? node6845 : node6838;
														assign node6838 = (inp[0]) ? node6842 : node6839;
															assign node6839 = (inp[15]) ? 4'b0001 : 4'b0011;
															assign node6842 = (inp[15]) ? 4'b0011 : 4'b0001;
														assign node6845 = (inp[15]) ? node6851 : node6846;
															assign node6846 = (inp[5]) ? 4'b0001 : node6847;
																assign node6847 = (inp[0]) ? 4'b0001 : 4'b0011;
															assign node6851 = (inp[0]) ? node6855 : node6852;
																assign node6852 = (inp[5]) ? 4'b0011 : 4'b0001;
																assign node6855 = (inp[5]) ? 4'b0001 : 4'b0011;
											assign node6858 = (inp[12]) ? node6896 : node6859;
												assign node6859 = (inp[5]) ? node6873 : node6860;
													assign node6860 = (inp[3]) ? node6866 : node6861;
														assign node6861 = (inp[0]) ? node6863 : 4'b0011;
															assign node6863 = (inp[15]) ? 4'b0011 : 4'b0001;
														assign node6866 = (inp[15]) ? node6870 : node6867;
															assign node6867 = (inp[0]) ? 4'b0001 : 4'b0011;
															assign node6870 = (inp[0]) ? 4'b0011 : 4'b0001;
													assign node6873 = (inp[10]) ? node6887 : node6874;
														assign node6874 = (inp[15]) ? node6880 : node6875;
															assign node6875 = (inp[0]) ? 4'b0011 : node6876;
																assign node6876 = (inp[3]) ? 4'b0001 : 4'b0011;
															assign node6880 = (inp[0]) ? node6884 : node6881;
																assign node6881 = (inp[3]) ? 4'b0011 : 4'b0001;
																assign node6884 = (inp[3]) ? 4'b0001 : 4'b0011;
														assign node6887 = (inp[3]) ? node6889 : 4'b0001;
															assign node6889 = (inp[15]) ? node6893 : node6890;
																assign node6890 = (inp[0]) ? 4'b0011 : 4'b0001;
																assign node6893 = (inp[0]) ? 4'b0001 : 4'b0011;
												assign node6896 = (inp[10]) ? node6910 : node6897;
													assign node6897 = (inp[3]) ? node6903 : node6898;
														assign node6898 = (inp[0]) ? 4'b0001 : node6899;
															assign node6899 = (inp[15]) ? 4'b0001 : 4'b0011;
														assign node6903 = (inp[0]) ? node6907 : node6904;
															assign node6904 = (inp[5]) ? 4'b0011 : 4'b0001;
															assign node6907 = (inp[5]) ? 4'b0001 : 4'b0011;
													assign node6910 = (inp[5]) ? node6918 : node6911;
														assign node6911 = (inp[3]) ? node6913 : 4'b0111;
															assign node6913 = (inp[15]) ? 4'b0101 : node6914;
																assign node6914 = (inp[0]) ? 4'b0111 : 4'b0101;
														assign node6918 = (inp[15]) ? node6922 : node6919;
															assign node6919 = (inp[0]) ? 4'b0111 : 4'b0101;
															assign node6922 = (inp[0]) ? 4'b0101 : 4'b0111;
										assign node6925 = (inp[4]) ? node6985 : node6926;
											assign node6926 = (inp[10]) ? node6948 : node6927;
												assign node6927 = (inp[15]) ? node6939 : node6928;
													assign node6928 = (inp[0]) ? node6934 : node6929;
														assign node6929 = (inp[5]) ? node6931 : 4'b0011;
															assign node6931 = (inp[3]) ? 4'b0001 : 4'b0011;
														assign node6934 = (inp[3]) ? node6936 : 4'b0001;
															assign node6936 = (inp[5]) ? 4'b0011 : 4'b0001;
													assign node6939 = (inp[0]) ? node6945 : node6940;
														assign node6940 = (inp[5]) ? node6942 : 4'b0001;
															assign node6942 = (inp[3]) ? 4'b0011 : 4'b0001;
														assign node6945 = (inp[3]) ? 4'b0001 : 4'b0011;
												assign node6948 = (inp[12]) ? node6964 : node6949;
													assign node6949 = (inp[15]) ? node6957 : node6950;
														assign node6950 = (inp[0]) ? node6954 : node6951;
															assign node6951 = (inp[3]) ? 4'b0001 : 4'b0011;
															assign node6954 = (inp[5]) ? 4'b0011 : 4'b0001;
														assign node6957 = (inp[5]) ? node6959 : 4'b0011;
															assign node6959 = (inp[3]) ? node6961 : 4'b0011;
																assign node6961 = (inp[0]) ? 4'b0001 : 4'b0011;
													assign node6964 = (inp[5]) ? node6980 : node6965;
														assign node6965 = (inp[15]) ? node6973 : node6966;
															assign node6966 = (inp[3]) ? node6970 : node6967;
																assign node6967 = (inp[0]) ? 4'b0101 : 4'b0111;
																assign node6970 = (inp[0]) ? 4'b0111 : 4'b0101;
															assign node6973 = (inp[3]) ? node6977 : node6974;
																assign node6974 = (inp[0]) ? 4'b0111 : 4'b0101;
																assign node6977 = (inp[0]) ? 4'b0101 : 4'b0111;
														assign node6980 = (inp[0]) ? node6982 : 4'b0101;
															assign node6982 = (inp[15]) ? 4'b0101 : 4'b0111;
											assign node6985 = (inp[10]) ? node7013 : node6986;
												assign node6986 = (inp[3]) ? node7006 : node6987;
													assign node6987 = (inp[0]) ? node6995 : node6988;
														assign node6988 = (inp[15]) ? node6992 : node6989;
															assign node6989 = (inp[5]) ? 4'b0101 : 4'b0111;
															assign node6992 = (inp[5]) ? 4'b0111 : 4'b0101;
														assign node6995 = (inp[12]) ? node7001 : node6996;
															assign node6996 = (inp[15]) ? node6998 : 4'b0101;
																assign node6998 = (inp[5]) ? 4'b0101 : 4'b0111;
															assign node7001 = (inp[5]) ? node7003 : 4'b0101;
																assign node7003 = (inp[15]) ? 4'b0101 : 4'b0111;
													assign node7006 = (inp[15]) ? node7010 : node7007;
														assign node7007 = (inp[0]) ? 4'b0111 : 4'b0101;
														assign node7010 = (inp[0]) ? 4'b0101 : 4'b0111;
												assign node7013 = (inp[12]) ? node7025 : node7014;
													assign node7014 = (inp[0]) ? node7022 : node7015;
														assign node7015 = (inp[15]) ? node7019 : node7016;
															assign node7016 = (inp[5]) ? 4'b0101 : 4'b0111;
															assign node7019 = (inp[5]) ? 4'b0111 : 4'b0101;
														assign node7022 = (inp[15]) ? 4'b0101 : 4'b0111;
													assign node7025 = (inp[5]) ? node7035 : node7026;
														assign node7026 = (inp[0]) ? 4'b0011 : node7027;
															assign node7027 = (inp[3]) ? node7031 : node7028;
																assign node7028 = (inp[15]) ? 4'b0001 : 4'b0011;
																assign node7031 = (inp[15]) ? 4'b0011 : 4'b0001;
														assign node7035 = (inp[0]) ? 4'b0001 : node7036;
															assign node7036 = (inp[3]) ? 4'b0001 : 4'b0011;
								assign node7040 = (inp[10]) ? node7248 : node7041;
									assign node7041 = (inp[12]) ? node7149 : node7042;
										assign node7042 = (inp[4]) ? node7092 : node7043;
											assign node7043 = (inp[9]) ? node7059 : node7044;
												assign node7044 = (inp[0]) ? node7052 : node7045;
													assign node7045 = (inp[15]) ? 4'b0101 : node7046;
														assign node7046 = (inp[3]) ? node7048 : 4'b0111;
															assign node7048 = (inp[5]) ? 4'b0101 : 4'b0111;
													assign node7052 = (inp[15]) ? 4'b0111 : node7053;
														assign node7053 = (inp[5]) ? node7055 : 4'b0101;
															assign node7055 = (inp[3]) ? 4'b0111 : 4'b0101;
												assign node7059 = (inp[2]) ? node7077 : node7060;
													assign node7060 = (inp[0]) ? node7072 : node7061;
														assign node7061 = (inp[15]) ? node7067 : node7062;
															assign node7062 = (inp[5]) ? node7064 : 4'b0011;
																assign node7064 = (inp[3]) ? 4'b0001 : 4'b0011;
															assign node7067 = (inp[5]) ? node7069 : 4'b0001;
																assign node7069 = (inp[3]) ? 4'b0011 : 4'b0001;
														assign node7072 = (inp[3]) ? 4'b0011 : node7073;
															assign node7073 = (inp[15]) ? 4'b0011 : 4'b0001;
													assign node7077 = (inp[15]) ? node7083 : node7078;
														assign node7078 = (inp[0]) ? 4'b0001 : node7079;
															assign node7079 = (inp[5]) ? 4'b0001 : 4'b0011;
														assign node7083 = (inp[0]) ? node7087 : node7084;
															assign node7084 = (inp[3]) ? 4'b0011 : 4'b0001;
															assign node7087 = (inp[3]) ? node7089 : 4'b0011;
																assign node7089 = (inp[5]) ? 4'b0001 : 4'b0011;
											assign node7092 = (inp[9]) ? node7116 : node7093;
												assign node7093 = (inp[0]) ? node7105 : node7094;
													assign node7094 = (inp[15]) ? node7100 : node7095;
														assign node7095 = (inp[3]) ? node7097 : 4'b0011;
															assign node7097 = (inp[5]) ? 4'b0001 : 4'b0011;
														assign node7100 = (inp[5]) ? node7102 : 4'b0001;
															assign node7102 = (inp[3]) ? 4'b0011 : 4'b0001;
													assign node7105 = (inp[15]) ? node7111 : node7106;
														assign node7106 = (inp[5]) ? node7108 : 4'b0001;
															assign node7108 = (inp[2]) ? 4'b0001 : 4'b0011;
														assign node7111 = (inp[3]) ? node7113 : 4'b0011;
															assign node7113 = (inp[5]) ? 4'b0001 : 4'b0011;
												assign node7116 = (inp[2]) ? node7130 : node7117;
													assign node7117 = (inp[15]) ? node7123 : node7118;
														assign node7118 = (inp[0]) ? node7120 : 4'b0101;
															assign node7120 = (inp[5]) ? 4'b0111 : 4'b0101;
														assign node7123 = (inp[0]) ? 4'b0101 : node7124;
															assign node7124 = (inp[3]) ? 4'b0111 : node7125;
																assign node7125 = (inp[5]) ? 4'b0111 : 4'b0101;
													assign node7130 = (inp[15]) ? node7140 : node7131;
														assign node7131 = (inp[0]) ? node7135 : node7132;
															assign node7132 = (inp[5]) ? 4'b0101 : 4'b0111;
															assign node7135 = (inp[5]) ? 4'b0111 : node7136;
																assign node7136 = (inp[3]) ? 4'b0111 : 4'b0101;
														assign node7140 = (inp[3]) ? 4'b0101 : node7141;
															assign node7141 = (inp[0]) ? node7145 : node7142;
																assign node7142 = (inp[5]) ? 4'b0111 : 4'b0101;
																assign node7145 = (inp[5]) ? 4'b0101 : 4'b0111;
										assign node7149 = (inp[0]) ? node7193 : node7150;
											assign node7150 = (inp[15]) ? node7172 : node7151;
												assign node7151 = (inp[3]) ? node7159 : node7152;
													assign node7152 = (inp[9]) ? node7156 : node7153;
														assign node7153 = (inp[4]) ? 4'b0011 : 4'b0111;
														assign node7156 = (inp[4]) ? 4'b0111 : 4'b0011;
													assign node7159 = (inp[5]) ? node7165 : node7160;
														assign node7160 = (inp[9]) ? node7162 : 4'b0011;
															assign node7162 = (inp[4]) ? 4'b0101 : 4'b0011;
														assign node7165 = (inp[9]) ? node7169 : node7166;
															assign node7166 = (inp[4]) ? 4'b0001 : 4'b0101;
															assign node7169 = (inp[4]) ? 4'b0101 : 4'b0001;
												assign node7172 = (inp[5]) ? node7178 : node7173;
													assign node7173 = (inp[4]) ? 4'b0001 : node7174;
														assign node7174 = (inp[9]) ? 4'b0001 : 4'b0101;
													assign node7178 = (inp[3]) ? node7186 : node7179;
														assign node7179 = (inp[9]) ? node7183 : node7180;
															assign node7180 = (inp[4]) ? 4'b0001 : 4'b0101;
															assign node7183 = (inp[4]) ? 4'b0111 : 4'b0001;
														assign node7186 = (inp[9]) ? node7190 : node7187;
															assign node7187 = (inp[4]) ? 4'b0011 : 4'b0111;
															assign node7190 = (inp[4]) ? 4'b0111 : 4'b0011;
											assign node7193 = (inp[15]) ? node7217 : node7194;
												assign node7194 = (inp[3]) ? node7204 : node7195;
													assign node7195 = (inp[4]) ? node7199 : node7196;
														assign node7196 = (inp[9]) ? 4'b0001 : 4'b0101;
														assign node7199 = (inp[9]) ? node7201 : 4'b0001;
															assign node7201 = (inp[5]) ? 4'b0111 : 4'b0101;
													assign node7204 = (inp[5]) ? node7212 : node7205;
														assign node7205 = (inp[9]) ? node7209 : node7206;
															assign node7206 = (inp[4]) ? 4'b0001 : 4'b0101;
															assign node7209 = (inp[4]) ? 4'b0111 : 4'b0001;
														assign node7212 = (inp[9]) ? node7214 : 4'b0011;
															assign node7214 = (inp[4]) ? 4'b0111 : 4'b0011;
												assign node7217 = (inp[5]) ? node7233 : node7218;
													assign node7218 = (inp[3]) ? node7226 : node7219;
														assign node7219 = (inp[9]) ? node7223 : node7220;
															assign node7220 = (inp[4]) ? 4'b0011 : 4'b0111;
															assign node7223 = (inp[4]) ? 4'b0111 : 4'b0011;
														assign node7226 = (inp[9]) ? node7230 : node7227;
															assign node7227 = (inp[4]) ? 4'b0011 : 4'b0111;
															assign node7230 = (inp[4]) ? 4'b0101 : 4'b0011;
													assign node7233 = (inp[3]) ? node7241 : node7234;
														assign node7234 = (inp[9]) ? node7238 : node7235;
															assign node7235 = (inp[4]) ? 4'b0011 : 4'b0111;
															assign node7238 = (inp[4]) ? 4'b0101 : 4'b0011;
														assign node7241 = (inp[2]) ? node7243 : 4'b0101;
															assign node7243 = (inp[4]) ? node7245 : 4'b0001;
																assign node7245 = (inp[9]) ? 4'b0101 : 4'b0001;
									assign node7248 = (inp[12]) ? node7420 : node7249;
										assign node7249 = (inp[2]) ? node7333 : node7250;
											assign node7250 = (inp[3]) ? node7290 : node7251;
												assign node7251 = (inp[9]) ? node7271 : node7252;
													assign node7252 = (inp[4]) ? node7260 : node7253;
														assign node7253 = (inp[0]) ? node7257 : node7254;
															assign node7254 = (inp[15]) ? 4'b0101 : 4'b0111;
															assign node7257 = (inp[15]) ? 4'b0111 : 4'b0101;
														assign node7260 = (inp[5]) ? node7266 : node7261;
															assign node7261 = (inp[0]) ? 4'b0011 : node7262;
																assign node7262 = (inp[15]) ? 4'b0001 : 4'b0011;
															assign node7266 = (inp[0]) ? node7268 : 4'b0001;
																assign node7268 = (inp[15]) ? 4'b0011 : 4'b0001;
													assign node7271 = (inp[4]) ? node7279 : node7272;
														assign node7272 = (inp[0]) ? node7276 : node7273;
															assign node7273 = (inp[15]) ? 4'b0001 : 4'b0011;
															assign node7276 = (inp[15]) ? 4'b0011 : 4'b0001;
														assign node7279 = (inp[5]) ? node7285 : node7280;
															assign node7280 = (inp[0]) ? node7282 : 4'b0101;
																assign node7282 = (inp[15]) ? 4'b0111 : 4'b0101;
															assign node7285 = (inp[0]) ? node7287 : 4'b0111;
																assign node7287 = (inp[15]) ? 4'b0101 : 4'b0111;
												assign node7290 = (inp[15]) ? node7306 : node7291;
													assign node7291 = (inp[5]) ? node7297 : node7292;
														assign node7292 = (inp[0]) ? node7294 : 4'b0011;
															assign node7294 = (inp[4]) ? 4'b0001 : 4'b0101;
														assign node7297 = (inp[0]) ? node7303 : node7298;
															assign node7298 = (inp[4]) ? 4'b0101 : node7299;
																assign node7299 = (inp[9]) ? 4'b0001 : 4'b0101;
															assign node7303 = (inp[4]) ? 4'b0011 : 4'b0111;
													assign node7306 = (inp[0]) ? node7318 : node7307;
														assign node7307 = (inp[5]) ? node7313 : node7308;
															assign node7308 = (inp[9]) ? 4'b0111 : node7309;
																assign node7309 = (inp[4]) ? 4'b0001 : 4'b0101;
															assign node7313 = (inp[4]) ? 4'b0111 : node7314;
																assign node7314 = (inp[9]) ? 4'b0011 : 4'b0111;
														assign node7318 = (inp[5]) ? node7326 : node7319;
															assign node7319 = (inp[4]) ? node7323 : node7320;
																assign node7320 = (inp[9]) ? 4'b0011 : 4'b0111;
																assign node7323 = (inp[9]) ? 4'b0101 : 4'b0011;
															assign node7326 = (inp[9]) ? node7330 : node7327;
																assign node7327 = (inp[4]) ? 4'b0001 : 4'b0101;
																assign node7330 = (inp[4]) ? 4'b0101 : 4'b0001;
											assign node7333 = (inp[0]) ? node7381 : node7334;
												assign node7334 = (inp[15]) ? node7358 : node7335;
													assign node7335 = (inp[3]) ? node7345 : node7336;
														assign node7336 = (inp[9]) ? node7340 : node7337;
															assign node7337 = (inp[4]) ? 4'b0011 : 4'b0111;
															assign node7340 = (inp[4]) ? node7342 : 4'b0011;
																assign node7342 = (inp[5]) ? 4'b0101 : 4'b0111;
														assign node7345 = (inp[5]) ? node7353 : node7346;
															assign node7346 = (inp[9]) ? node7350 : node7347;
																assign node7347 = (inp[4]) ? 4'b0011 : 4'b0111;
																assign node7350 = (inp[4]) ? 4'b0101 : 4'b0011;
															assign node7353 = (inp[9]) ? 4'b0001 : node7354;
																assign node7354 = (inp[4]) ? 4'b0001 : 4'b0101;
													assign node7358 = (inp[3]) ? node7366 : node7359;
														assign node7359 = (inp[4]) ? node7363 : node7360;
															assign node7360 = (inp[5]) ? 4'b0101 : 4'b0001;
															assign node7363 = (inp[9]) ? 4'b0101 : 4'b0001;
														assign node7366 = (inp[5]) ? node7374 : node7367;
															assign node7367 = (inp[4]) ? node7371 : node7368;
																assign node7368 = (inp[9]) ? 4'b0001 : 4'b0101;
																assign node7371 = (inp[9]) ? 4'b0111 : 4'b0001;
															assign node7374 = (inp[9]) ? node7378 : node7375;
																assign node7375 = (inp[4]) ? 4'b0011 : 4'b0111;
																assign node7378 = (inp[4]) ? 4'b0111 : 4'b0011;
												assign node7381 = (inp[15]) ? node7405 : node7382;
													assign node7382 = (inp[3]) ? node7392 : node7383;
														assign node7383 = (inp[5]) ? node7385 : 4'b0101;
															assign node7385 = (inp[4]) ? node7389 : node7386;
																assign node7386 = (inp[9]) ? 4'b0001 : 4'b0101;
																assign node7389 = (inp[9]) ? 4'b0111 : 4'b0001;
														assign node7392 = (inp[5]) ? node7398 : node7393;
															assign node7393 = (inp[9]) ? 4'b0111 : node7394;
																assign node7394 = (inp[4]) ? 4'b0001 : 4'b0101;
															assign node7398 = (inp[4]) ? node7402 : node7399;
																assign node7399 = (inp[9]) ? 4'b0011 : 4'b0111;
																assign node7402 = (inp[9]) ? 4'b0111 : 4'b0011;
													assign node7405 = (inp[9]) ? node7409 : node7406;
														assign node7406 = (inp[4]) ? 4'b0011 : 4'b0111;
														assign node7409 = (inp[4]) ? node7415 : node7410;
															assign node7410 = (inp[5]) ? node7412 : 4'b0011;
																assign node7412 = (inp[3]) ? 4'b0001 : 4'b0011;
															assign node7415 = (inp[5]) ? 4'b0101 : node7416;
																assign node7416 = (inp[3]) ? 4'b0101 : 4'b0111;
										assign node7420 = (inp[2]) ? node7508 : node7421;
											assign node7421 = (inp[3]) ? node7469 : node7422;
												assign node7422 = (inp[9]) ? node7438 : node7423;
													assign node7423 = (inp[4]) ? node7431 : node7424;
														assign node7424 = (inp[0]) ? node7428 : node7425;
															assign node7425 = (inp[15]) ? 4'b0001 : 4'b0011;
															assign node7428 = (inp[15]) ? 4'b0011 : 4'b0001;
														assign node7431 = (inp[5]) ? 4'b0111 : node7432;
															assign node7432 = (inp[0]) ? 4'b0101 : node7433;
																assign node7433 = (inp[15]) ? 4'b0101 : 4'b0111;
													assign node7438 = (inp[4]) ? node7454 : node7439;
														assign node7439 = (inp[15]) ? node7447 : node7440;
															assign node7440 = (inp[0]) ? node7444 : node7441;
																assign node7441 = (inp[5]) ? 4'b0101 : 4'b0111;
																assign node7444 = (inp[5]) ? 4'b0111 : 4'b0101;
															assign node7447 = (inp[0]) ? node7451 : node7448;
																assign node7448 = (inp[5]) ? 4'b0111 : 4'b0101;
																assign node7451 = (inp[5]) ? 4'b0101 : 4'b0111;
														assign node7454 = (inp[15]) ? node7462 : node7455;
															assign node7455 = (inp[0]) ? node7459 : node7456;
																assign node7456 = (inp[5]) ? 4'b0001 : 4'b0011;
																assign node7459 = (inp[5]) ? 4'b0011 : 4'b0001;
															assign node7462 = (inp[5]) ? node7466 : node7463;
																assign node7463 = (inp[0]) ? 4'b0011 : 4'b0001;
																assign node7466 = (inp[0]) ? 4'b0001 : 4'b0011;
												assign node7469 = (inp[4]) ? node7491 : node7470;
													assign node7470 = (inp[9]) ? node7486 : node7471;
														assign node7471 = (inp[15]) ? node7479 : node7472;
															assign node7472 = (inp[5]) ? node7476 : node7473;
																assign node7473 = (inp[0]) ? 4'b0001 : 4'b0011;
																assign node7476 = (inp[0]) ? 4'b0011 : 4'b0001;
															assign node7479 = (inp[5]) ? node7483 : node7480;
																assign node7480 = (inp[0]) ? 4'b0011 : 4'b0001;
																assign node7483 = (inp[0]) ? 4'b0001 : 4'b0011;
														assign node7486 = (inp[0]) ? 4'b0111 : node7487;
															assign node7487 = (inp[15]) ? 4'b0111 : 4'b0101;
													assign node7491 = (inp[9]) ? node7497 : node7492;
														assign node7492 = (inp[0]) ? node7494 : 4'b0111;
															assign node7494 = (inp[15]) ? 4'b0101 : 4'b0111;
														assign node7497 = (inp[5]) ? node7503 : node7498;
															assign node7498 = (inp[0]) ? 4'b0011 : node7499;
																assign node7499 = (inp[15]) ? 4'b0011 : 4'b0001;
															assign node7503 = (inp[15]) ? node7505 : 4'b0011;
																assign node7505 = (inp[0]) ? 4'b0001 : 4'b0011;
											assign node7508 = (inp[0]) ? node7552 : node7509;
												assign node7509 = (inp[15]) ? node7527 : node7510;
													assign node7510 = (inp[5]) ? node7518 : node7511;
														assign node7511 = (inp[3]) ? node7513 : 4'b0011;
															assign node7513 = (inp[9]) ? 4'b0101 : node7514;
																assign node7514 = (inp[4]) ? 4'b0101 : 4'b0011;
														assign node7518 = (inp[4]) ? node7524 : node7519;
															assign node7519 = (inp[9]) ? 4'b0101 : node7520;
																assign node7520 = (inp[3]) ? 4'b0001 : 4'b0011;
															assign node7524 = (inp[9]) ? 4'b0001 : 4'b0101;
													assign node7527 = (inp[5]) ? node7543 : node7528;
														assign node7528 = (inp[3]) ? node7536 : node7529;
															assign node7529 = (inp[4]) ? node7533 : node7530;
																assign node7530 = (inp[9]) ? 4'b0101 : 4'b0001;
																assign node7533 = (inp[9]) ? 4'b0001 : 4'b0101;
															assign node7536 = (inp[9]) ? node7540 : node7537;
																assign node7537 = (inp[4]) ? 4'b0111 : 4'b0001;
																assign node7540 = (inp[4]) ? 4'b0011 : 4'b0111;
														assign node7543 = (inp[3]) ? node7545 : 4'b0111;
															assign node7545 = (inp[9]) ? node7549 : node7546;
																assign node7546 = (inp[4]) ? 4'b0111 : 4'b0011;
																assign node7549 = (inp[4]) ? 4'b0011 : 4'b0111;
												assign node7552 = (inp[15]) ? node7574 : node7553;
													assign node7553 = (inp[5]) ? node7565 : node7554;
														assign node7554 = (inp[3]) ? node7558 : node7555;
															assign node7555 = (inp[4]) ? 4'b0001 : 4'b0101;
															assign node7558 = (inp[9]) ? node7562 : node7559;
																assign node7559 = (inp[4]) ? 4'b0111 : 4'b0001;
																assign node7562 = (inp[4]) ? 4'b0011 : 4'b0111;
														assign node7565 = (inp[9]) ? node7571 : node7566;
															assign node7566 = (inp[4]) ? 4'b0111 : node7567;
																assign node7567 = (inp[3]) ? 4'b0011 : 4'b0001;
															assign node7571 = (inp[4]) ? 4'b0011 : 4'b0111;
													assign node7574 = (inp[3]) ? node7586 : node7575;
														assign node7575 = (inp[5]) ? node7583 : node7576;
															assign node7576 = (inp[4]) ? node7580 : node7577;
																assign node7577 = (inp[9]) ? 4'b0111 : 4'b0011;
																assign node7580 = (inp[9]) ? 4'b0011 : 4'b0111;
															assign node7583 = (inp[9]) ? 4'b0001 : 4'b0011;
														assign node7586 = (inp[9]) ? node7592 : node7587;
															assign node7587 = (inp[4]) ? 4'b0101 : node7588;
																assign node7588 = (inp[5]) ? 4'b0001 : 4'b0011;
															assign node7592 = (inp[4]) ? 4'b0001 : 4'b0101;
							assign node7595 = (inp[2]) ? node8135 : node7596;
								assign node7596 = (inp[14]) ? node7892 : node7597;
									assign node7597 = (inp[15]) ? node7737 : node7598;
										assign node7598 = (inp[0]) ? node7674 : node7599;
											assign node7599 = (inp[5]) ? node7641 : node7600;
												assign node7600 = (inp[3]) ? node7624 : node7601;
													assign node7601 = (inp[9]) ? node7613 : node7602;
														assign node7602 = (inp[4]) ? node7608 : node7603;
															assign node7603 = (inp[12]) ? node7605 : 4'b0111;
																assign node7605 = (inp[10]) ? 4'b0011 : 4'b0111;
															assign node7608 = (inp[12]) ? node7610 : 4'b0011;
																assign node7610 = (inp[10]) ? 4'b0111 : 4'b0011;
														assign node7613 = (inp[4]) ? node7619 : node7614;
															assign node7614 = (inp[10]) ? node7616 : 4'b0011;
																assign node7616 = (inp[12]) ? 4'b0111 : 4'b0011;
															assign node7619 = (inp[10]) ? node7621 : 4'b0111;
																assign node7621 = (inp[12]) ? 4'b0011 : 4'b0111;
													assign node7624 = (inp[9]) ? node7632 : node7625;
														assign node7625 = (inp[4]) ? 4'b0011 : node7626;
															assign node7626 = (inp[12]) ? node7628 : 4'b0111;
																assign node7628 = (inp[10]) ? 4'b0011 : 4'b0111;
														assign node7632 = (inp[4]) ? node7638 : node7633;
															assign node7633 = (inp[12]) ? node7635 : 4'b0011;
																assign node7635 = (inp[10]) ? 4'b0101 : 4'b0011;
															assign node7638 = (inp[10]) ? 4'b0001 : 4'b0101;
												assign node7641 = (inp[3]) ? node7659 : node7642;
													assign node7642 = (inp[4]) ? node7650 : node7643;
														assign node7643 = (inp[9]) ? 4'b0011 : node7644;
															assign node7644 = (inp[12]) ? node7646 : 4'b0111;
																assign node7646 = (inp[10]) ? 4'b0011 : 4'b0111;
														assign node7650 = (inp[9]) ? node7656 : node7651;
															assign node7651 = (inp[10]) ? node7653 : 4'b0011;
																assign node7653 = (inp[12]) ? 4'b0101 : 4'b0011;
															assign node7656 = (inp[10]) ? 4'b0001 : 4'b0101;
													assign node7659 = (inp[12]) ? node7665 : node7660;
														assign node7660 = (inp[4]) ? node7662 : 4'b0101;
															assign node7662 = (inp[9]) ? 4'b0101 : 4'b0001;
														assign node7665 = (inp[4]) ? 4'b0001 : node7666;
															assign node7666 = (inp[10]) ? node7670 : node7667;
																assign node7667 = (inp[9]) ? 4'b0001 : 4'b0101;
																assign node7670 = (inp[9]) ? 4'b0101 : 4'b0001;
											assign node7674 = (inp[5]) ? node7700 : node7675;
												assign node7675 = (inp[4]) ? node7689 : node7676;
													assign node7676 = (inp[9]) ? node7682 : node7677;
														assign node7677 = (inp[12]) ? node7679 : 4'b0101;
															assign node7679 = (inp[10]) ? 4'b0001 : 4'b0101;
														assign node7682 = (inp[12]) ? node7684 : 4'b0001;
															assign node7684 = (inp[10]) ? node7686 : 4'b0001;
																assign node7686 = (inp[3]) ? 4'b0111 : 4'b0101;
													assign node7689 = (inp[12]) ? node7691 : 4'b0111;
														assign node7691 = (inp[3]) ? node7697 : node7692;
															assign node7692 = (inp[9]) ? node7694 : 4'b0101;
																assign node7694 = (inp[10]) ? 4'b0001 : 4'b0101;
															assign node7697 = (inp[10]) ? 4'b0111 : 4'b0001;
												assign node7700 = (inp[3]) ? node7716 : node7701;
													assign node7701 = (inp[9]) ? node7709 : node7702;
														assign node7702 = (inp[10]) ? node7704 : 4'b0001;
															assign node7704 = (inp[4]) ? 4'b0111 : node7705;
																assign node7705 = (inp[12]) ? 4'b0001 : 4'b0101;
														assign node7709 = (inp[4]) ? 4'b0111 : node7710;
															assign node7710 = (inp[10]) ? node7712 : 4'b0001;
																assign node7712 = (inp[12]) ? 4'b0111 : 4'b0001;
													assign node7716 = (inp[10]) ? node7722 : node7717;
														assign node7717 = (inp[4]) ? node7719 : 4'b0111;
															assign node7719 = (inp[9]) ? 4'b0111 : 4'b0011;
														assign node7722 = (inp[4]) ? node7730 : node7723;
															assign node7723 = (inp[12]) ? node7727 : node7724;
																assign node7724 = (inp[9]) ? 4'b0011 : 4'b0111;
																assign node7727 = (inp[9]) ? 4'b0111 : 4'b0011;
															assign node7730 = (inp[12]) ? node7734 : node7731;
																assign node7731 = (inp[9]) ? 4'b0111 : 4'b0011;
																assign node7734 = (inp[9]) ? 4'b0011 : 4'b0111;
										assign node7737 = (inp[5]) ? node7819 : node7738;
											assign node7738 = (inp[0]) ? node7776 : node7739;
												assign node7739 = (inp[3]) ? node7759 : node7740;
													assign node7740 = (inp[10]) ? node7748 : node7741;
														assign node7741 = (inp[12]) ? node7743 : 4'b0001;
															assign node7743 = (inp[4]) ? 4'b0101 : node7744;
																assign node7744 = (inp[9]) ? 4'b0001 : 4'b0101;
														assign node7748 = (inp[12]) ? node7754 : node7749;
															assign node7749 = (inp[4]) ? node7751 : 4'b0101;
																assign node7751 = (inp[9]) ? 4'b0101 : 4'b0001;
															assign node7754 = (inp[9]) ? 4'b0001 : node7755;
																assign node7755 = (inp[4]) ? 4'b0101 : 4'b0001;
													assign node7759 = (inp[12]) ? node7765 : node7760;
														assign node7760 = (inp[9]) ? 4'b0001 : node7761;
															assign node7761 = (inp[4]) ? 4'b0001 : 4'b0101;
														assign node7765 = (inp[4]) ? node7771 : node7766;
															assign node7766 = (inp[9]) ? 4'b0111 : node7767;
																assign node7767 = (inp[10]) ? 4'b0001 : 4'b0101;
															assign node7771 = (inp[9]) ? node7773 : 4'b0111;
																assign node7773 = (inp[10]) ? 4'b0011 : 4'b0111;
												assign node7776 = (inp[3]) ? node7802 : node7777;
													assign node7777 = (inp[10]) ? node7787 : node7778;
														assign node7778 = (inp[12]) ? 4'b0011 : node7779;
															assign node7779 = (inp[9]) ? node7783 : node7780;
																assign node7780 = (inp[4]) ? 4'b0011 : 4'b0111;
																assign node7783 = (inp[4]) ? 4'b0111 : 4'b0011;
														assign node7787 = (inp[12]) ? node7795 : node7788;
															assign node7788 = (inp[4]) ? node7792 : node7789;
																assign node7789 = (inp[9]) ? 4'b0011 : 4'b0111;
																assign node7792 = (inp[9]) ? 4'b0111 : 4'b0011;
															assign node7795 = (inp[4]) ? node7799 : node7796;
																assign node7796 = (inp[9]) ? 4'b0111 : 4'b0011;
																assign node7799 = (inp[9]) ? 4'b0011 : 4'b0111;
													assign node7802 = (inp[4]) ? node7812 : node7803;
														assign node7803 = (inp[9]) ? node7807 : node7804;
															assign node7804 = (inp[12]) ? 4'b0011 : 4'b0111;
															assign node7807 = (inp[10]) ? node7809 : 4'b0011;
																assign node7809 = (inp[12]) ? 4'b0101 : 4'b0011;
														assign node7812 = (inp[9]) ? 4'b0101 : node7813;
															assign node7813 = (inp[12]) ? node7815 : 4'b0011;
																assign node7815 = (inp[10]) ? 4'b0101 : 4'b0011;
											assign node7819 = (inp[0]) ? node7855 : node7820;
												assign node7820 = (inp[3]) ? node7836 : node7821;
													assign node7821 = (inp[9]) ? node7827 : node7822;
														assign node7822 = (inp[4]) ? 4'b0001 : node7823;
															assign node7823 = (inp[10]) ? 4'b0001 : 4'b0101;
														assign node7827 = (inp[4]) ? node7831 : node7828;
															assign node7828 = (inp[10]) ? 4'b0111 : 4'b0001;
															assign node7831 = (inp[10]) ? node7833 : 4'b0111;
																assign node7833 = (inp[12]) ? 4'b0011 : 4'b0111;
													assign node7836 = (inp[9]) ? node7846 : node7837;
														assign node7837 = (inp[12]) ? node7839 : 4'b0011;
															assign node7839 = (inp[4]) ? node7843 : node7840;
																assign node7840 = (inp[10]) ? 4'b0011 : 4'b0111;
																assign node7843 = (inp[10]) ? 4'b0111 : 4'b0011;
														assign node7846 = (inp[4]) ? node7852 : node7847;
															assign node7847 = (inp[10]) ? node7849 : 4'b0011;
																assign node7849 = (inp[12]) ? 4'b0111 : 4'b0011;
															assign node7852 = (inp[12]) ? 4'b0011 : 4'b0111;
												assign node7855 = (inp[3]) ? node7873 : node7856;
													assign node7856 = (inp[4]) ? node7866 : node7857;
														assign node7857 = (inp[9]) ? node7863 : node7858;
															assign node7858 = (inp[12]) ? node7860 : 4'b0111;
																assign node7860 = (inp[10]) ? 4'b0011 : 4'b0111;
															assign node7863 = (inp[10]) ? 4'b0101 : 4'b0011;
														assign node7866 = (inp[9]) ? node7870 : node7867;
															assign node7867 = (inp[10]) ? 4'b0101 : 4'b0011;
															assign node7870 = (inp[10]) ? 4'b0001 : 4'b0101;
													assign node7873 = (inp[4]) ? node7885 : node7874;
														assign node7874 = (inp[9]) ? node7880 : node7875;
															assign node7875 = (inp[10]) ? node7877 : 4'b0101;
																assign node7877 = (inp[12]) ? 4'b0001 : 4'b0101;
															assign node7880 = (inp[10]) ? node7882 : 4'b0001;
																assign node7882 = (inp[12]) ? 4'b0101 : 4'b0001;
														assign node7885 = (inp[9]) ? node7887 : 4'b0001;
															assign node7887 = (inp[12]) ? node7889 : 4'b0101;
																assign node7889 = (inp[10]) ? 4'b0001 : 4'b0101;
									assign node7892 = (inp[9]) ? node8010 : node7893;
										assign node7893 = (inp[4]) ? node7947 : node7894;
											assign node7894 = (inp[10]) ? node7916 : node7895;
												assign node7895 = (inp[0]) ? node7907 : node7896;
													assign node7896 = (inp[15]) ? node7902 : node7897;
														assign node7897 = (inp[3]) ? node7899 : 4'b0110;
															assign node7899 = (inp[5]) ? 4'b0100 : 4'b0110;
														assign node7902 = (inp[5]) ? node7904 : 4'b0100;
															assign node7904 = (inp[3]) ? 4'b0110 : 4'b0100;
													assign node7907 = (inp[15]) ? node7911 : node7908;
														assign node7908 = (inp[5]) ? 4'b0110 : 4'b0100;
														assign node7911 = (inp[5]) ? node7913 : 4'b0110;
															assign node7913 = (inp[3]) ? 4'b0100 : 4'b0110;
												assign node7916 = (inp[12]) ? node7928 : node7917;
													assign node7917 = (inp[5]) ? node7923 : node7918;
														assign node7918 = (inp[0]) ? 4'b0110 : node7919;
															assign node7919 = (inp[15]) ? 4'b0100 : 4'b0110;
														assign node7923 = (inp[15]) ? 4'b0100 : node7924;
															assign node7924 = (inp[3]) ? 4'b0110 : 4'b0100;
													assign node7928 = (inp[3]) ? node7934 : node7929;
														assign node7929 = (inp[15]) ? node7931 : 4'b0000;
															assign node7931 = (inp[0]) ? 4'b0010 : 4'b0000;
														assign node7934 = (inp[15]) ? node7940 : node7935;
															assign node7935 = (inp[5]) ? 4'b0010 : node7936;
																assign node7936 = (inp[0]) ? 4'b0000 : 4'b0010;
															assign node7940 = (inp[5]) ? node7944 : node7941;
																assign node7941 = (inp[0]) ? 4'b0010 : 4'b0000;
																assign node7944 = (inp[0]) ? 4'b0000 : 4'b0010;
											assign node7947 = (inp[12]) ? node7971 : node7948;
												assign node7948 = (inp[0]) ? node7960 : node7949;
													assign node7949 = (inp[15]) ? node7955 : node7950;
														assign node7950 = (inp[5]) ? node7952 : 4'b0010;
															assign node7952 = (inp[3]) ? 4'b0000 : 4'b0010;
														assign node7955 = (inp[5]) ? node7957 : 4'b0000;
															assign node7957 = (inp[3]) ? 4'b0010 : 4'b0000;
													assign node7960 = (inp[15]) ? node7966 : node7961;
														assign node7961 = (inp[3]) ? node7963 : 4'b0000;
															assign node7963 = (inp[5]) ? 4'b0010 : 4'b0000;
														assign node7966 = (inp[5]) ? node7968 : 4'b0010;
															assign node7968 = (inp[3]) ? 4'b0000 : 4'b0010;
												assign node7971 = (inp[10]) ? node7993 : node7972;
													assign node7972 = (inp[5]) ? node7980 : node7973;
														assign node7973 = (inp[15]) ? node7977 : node7974;
															assign node7974 = (inp[0]) ? 4'b0000 : 4'b0010;
															assign node7977 = (inp[0]) ? 4'b0010 : 4'b0000;
														assign node7980 = (inp[3]) ? node7986 : node7981;
															assign node7981 = (inp[0]) ? node7983 : 4'b0000;
																assign node7983 = (inp[15]) ? 4'b0010 : 4'b0000;
															assign node7986 = (inp[15]) ? node7990 : node7987;
																assign node7987 = (inp[0]) ? 4'b0010 : 4'b0000;
																assign node7990 = (inp[0]) ? 4'b0000 : 4'b0010;
													assign node7993 = (inp[5]) ? node8005 : node7994;
														assign node7994 = (inp[0]) ? node8000 : node7995;
															assign node7995 = (inp[15]) ? 4'b0110 : node7996;
																assign node7996 = (inp[3]) ? 4'b0100 : 4'b0110;
															assign node8000 = (inp[15]) ? 4'b0100 : node8001;
																assign node8001 = (inp[3]) ? 4'b0110 : 4'b0100;
														assign node8005 = (inp[15]) ? 4'b0110 : node8006;
															assign node8006 = (inp[0]) ? 4'b0110 : 4'b0100;
										assign node8010 = (inp[4]) ? node8064 : node8011;
											assign node8011 = (inp[12]) ? node8035 : node8012;
												assign node8012 = (inp[5]) ? node8020 : node8013;
													assign node8013 = (inp[15]) ? node8017 : node8014;
														assign node8014 = (inp[0]) ? 4'b0000 : 4'b0010;
														assign node8017 = (inp[0]) ? 4'b0010 : 4'b0000;
													assign node8020 = (inp[15]) ? node8028 : node8021;
														assign node8021 = (inp[0]) ? node8025 : node8022;
															assign node8022 = (inp[3]) ? 4'b0000 : 4'b0010;
															assign node8025 = (inp[10]) ? 4'b0000 : 4'b0010;
														assign node8028 = (inp[3]) ? node8032 : node8029;
															assign node8029 = (inp[0]) ? 4'b0010 : 4'b0000;
															assign node8032 = (inp[0]) ? 4'b0000 : 4'b0010;
												assign node8035 = (inp[10]) ? node8051 : node8036;
													assign node8036 = (inp[5]) ? node8044 : node8037;
														assign node8037 = (inp[0]) ? node8041 : node8038;
															assign node8038 = (inp[15]) ? 4'b0000 : 4'b0010;
															assign node8041 = (inp[15]) ? 4'b0010 : 4'b0000;
														assign node8044 = (inp[0]) ? node8046 : 4'b0010;
															assign node8046 = (inp[3]) ? node8048 : 4'b0010;
																assign node8048 = (inp[15]) ? 4'b0000 : 4'b0010;
													assign node8051 = (inp[15]) ? node8059 : node8052;
														assign node8052 = (inp[0]) ? 4'b0110 : node8053;
															assign node8053 = (inp[5]) ? 4'b0100 : node8054;
																assign node8054 = (inp[3]) ? 4'b0100 : 4'b0110;
														assign node8059 = (inp[0]) ? 4'b0100 : node8060;
															assign node8060 = (inp[3]) ? 4'b0110 : 4'b0100;
											assign node8064 = (inp[12]) ? node8098 : node8065;
												assign node8065 = (inp[3]) ? node8083 : node8066;
													assign node8066 = (inp[10]) ? node8072 : node8067;
														assign node8067 = (inp[5]) ? node8069 : 4'b0110;
															assign node8069 = (inp[0]) ? 4'b0110 : 4'b0100;
														assign node8072 = (inp[5]) ? node8078 : node8073;
															assign node8073 = (inp[15]) ? 4'b0100 : node8074;
																assign node8074 = (inp[0]) ? 4'b0100 : 4'b0110;
															assign node8078 = (inp[15]) ? 4'b0110 : node8079;
																assign node8079 = (inp[0]) ? 4'b0110 : 4'b0100;
													assign node8083 = (inp[10]) ? node8091 : node8084;
														assign node8084 = (inp[0]) ? node8088 : node8085;
															assign node8085 = (inp[15]) ? 4'b0110 : 4'b0100;
															assign node8088 = (inp[15]) ? 4'b0100 : 4'b0110;
														assign node8091 = (inp[15]) ? node8095 : node8092;
															assign node8092 = (inp[0]) ? 4'b0110 : 4'b0100;
															assign node8095 = (inp[0]) ? 4'b0100 : 4'b0110;
												assign node8098 = (inp[10]) ? node8120 : node8099;
													assign node8099 = (inp[5]) ? node8111 : node8100;
														assign node8100 = (inp[3]) ? node8106 : node8101;
															assign node8101 = (inp[15]) ? 4'b0100 : node8102;
																assign node8102 = (inp[0]) ? 4'b0100 : 4'b0110;
															assign node8106 = (inp[15]) ? 4'b0110 : node8107;
																assign node8107 = (inp[0]) ? 4'b0110 : 4'b0100;
														assign node8111 = (inp[3]) ? node8117 : node8112;
															assign node8112 = (inp[15]) ? 4'b0110 : node8113;
																assign node8113 = (inp[0]) ? 4'b0110 : 4'b0100;
															assign node8117 = (inp[15]) ? 4'b0100 : 4'b0110;
													assign node8120 = (inp[15]) ? node8128 : node8121;
														assign node8121 = (inp[0]) ? node8125 : node8122;
															assign node8122 = (inp[3]) ? 4'b0000 : 4'b0010;
															assign node8125 = (inp[3]) ? 4'b0010 : 4'b0000;
														assign node8128 = (inp[5]) ? 4'b0010 : node8129;
															assign node8129 = (inp[3]) ? 4'b0010 : node8130;
																assign node8130 = (inp[0]) ? 4'b0010 : 4'b0000;
								assign node8135 = (inp[3]) ? node8421 : node8136;
									assign node8136 = (inp[10]) ? node8262 : node8137;
										assign node8137 = (inp[12]) ? node8179 : node8138;
											assign node8138 = (inp[0]) ? node8158 : node8139;
												assign node8139 = (inp[15]) ? node8149 : node8140;
													assign node8140 = (inp[9]) ? node8144 : node8141;
														assign node8141 = (inp[4]) ? 4'b0010 : 4'b0110;
														assign node8144 = (inp[4]) ? node8146 : 4'b0010;
															assign node8146 = (inp[5]) ? 4'b0100 : 4'b0110;
													assign node8149 = (inp[9]) ? node8153 : node8150;
														assign node8150 = (inp[4]) ? 4'b0000 : 4'b0100;
														assign node8153 = (inp[5]) ? 4'b0110 : node8154;
															assign node8154 = (inp[4]) ? 4'b0100 : 4'b0000;
												assign node8158 = (inp[15]) ? node8172 : node8159;
													assign node8159 = (inp[5]) ? node8165 : node8160;
														assign node8160 = (inp[9]) ? node8162 : 4'b0000;
															assign node8162 = (inp[4]) ? 4'b0100 : 4'b0000;
														assign node8165 = (inp[9]) ? node8169 : node8166;
															assign node8166 = (inp[4]) ? 4'b0000 : 4'b0100;
															assign node8169 = (inp[4]) ? 4'b0110 : 4'b0000;
													assign node8172 = (inp[4]) ? node8176 : node8173;
														assign node8173 = (inp[9]) ? 4'b0010 : 4'b0110;
														assign node8176 = (inp[9]) ? 4'b0110 : 4'b0010;
											assign node8179 = (inp[14]) ? node8221 : node8180;
												assign node8180 = (inp[15]) ? node8198 : node8181;
													assign node8181 = (inp[0]) ? node8189 : node8182;
														assign node8182 = (inp[5]) ? node8186 : node8183;
															assign node8183 = (inp[9]) ? 4'b0110 : 4'b0010;
															assign node8186 = (inp[4]) ? 4'b0100 : 4'b0110;
														assign node8189 = (inp[4]) ? node8193 : node8190;
															assign node8190 = (inp[9]) ? 4'b0000 : 4'b0100;
															assign node8193 = (inp[9]) ? node8195 : 4'b0000;
																assign node8195 = (inp[5]) ? 4'b0110 : 4'b0100;
													assign node8198 = (inp[0]) ? node8214 : node8199;
														assign node8199 = (inp[5]) ? node8207 : node8200;
															assign node8200 = (inp[4]) ? node8204 : node8201;
																assign node8201 = (inp[9]) ? 4'b0000 : 4'b0100;
																assign node8204 = (inp[9]) ? 4'b0100 : 4'b0000;
															assign node8207 = (inp[9]) ? node8211 : node8208;
																assign node8208 = (inp[4]) ? 4'b0000 : 4'b0100;
																assign node8211 = (inp[4]) ? 4'b0110 : 4'b0000;
														assign node8214 = (inp[9]) ? node8218 : node8215;
															assign node8215 = (inp[4]) ? 4'b0010 : 4'b0110;
															assign node8218 = (inp[4]) ? 4'b0100 : 4'b0010;
												assign node8221 = (inp[15]) ? node8245 : node8222;
													assign node8222 = (inp[0]) ? node8232 : node8223;
														assign node8223 = (inp[4]) ? node8227 : node8224;
															assign node8224 = (inp[9]) ? 4'b0010 : 4'b0110;
															assign node8227 = (inp[9]) ? node8229 : 4'b0010;
																assign node8229 = (inp[5]) ? 4'b0100 : 4'b0110;
														assign node8232 = (inp[5]) ? node8240 : node8233;
															assign node8233 = (inp[4]) ? node8237 : node8234;
																assign node8234 = (inp[9]) ? 4'b0000 : 4'b0100;
																assign node8237 = (inp[9]) ? 4'b0100 : 4'b0000;
															assign node8240 = (inp[9]) ? node8242 : 4'b0000;
																assign node8242 = (inp[4]) ? 4'b0110 : 4'b0000;
													assign node8245 = (inp[0]) ? node8253 : node8246;
														assign node8246 = (inp[4]) ? node8250 : node8247;
															assign node8247 = (inp[9]) ? 4'b0000 : 4'b0100;
															assign node8250 = (inp[5]) ? 4'b0110 : 4'b0000;
														assign node8253 = (inp[5]) ? node8259 : node8254;
															assign node8254 = (inp[9]) ? node8256 : 4'b0110;
																assign node8256 = (inp[4]) ? 4'b0110 : 4'b0010;
															assign node8259 = (inp[9]) ? 4'b0100 : 4'b0110;
										assign node8262 = (inp[5]) ? node8336 : node8263;
											assign node8263 = (inp[4]) ? node8305 : node8264;
												assign node8264 = (inp[12]) ? node8284 : node8265;
													assign node8265 = (inp[9]) ? node8277 : node8266;
														assign node8266 = (inp[14]) ? node8272 : node8267;
															assign node8267 = (inp[15]) ? 4'b0110 : node8268;
																assign node8268 = (inp[0]) ? 4'b0100 : 4'b0110;
															assign node8272 = (inp[0]) ? 4'b0110 : node8273;
																assign node8273 = (inp[15]) ? 4'b0100 : 4'b0110;
														assign node8277 = (inp[15]) ? node8281 : node8278;
															assign node8278 = (inp[0]) ? 4'b0000 : 4'b0010;
															assign node8281 = (inp[0]) ? 4'b0010 : 4'b0000;
													assign node8284 = (inp[9]) ? node8298 : node8285;
														assign node8285 = (inp[14]) ? node8293 : node8286;
															assign node8286 = (inp[0]) ? node8290 : node8287;
																assign node8287 = (inp[15]) ? 4'b0000 : 4'b0010;
																assign node8290 = (inp[15]) ? 4'b0010 : 4'b0000;
															assign node8293 = (inp[0]) ? node8295 : 4'b0000;
																assign node8295 = (inp[15]) ? 4'b0010 : 4'b0000;
														assign node8298 = (inp[15]) ? node8302 : node8299;
															assign node8299 = (inp[0]) ? 4'b0100 : 4'b0110;
															assign node8302 = (inp[0]) ? 4'b0110 : 4'b0100;
												assign node8305 = (inp[9]) ? node8321 : node8306;
													assign node8306 = (inp[12]) ? node8314 : node8307;
														assign node8307 = (inp[0]) ? node8311 : node8308;
															assign node8308 = (inp[15]) ? 4'b0000 : 4'b0010;
															assign node8311 = (inp[15]) ? 4'b0010 : 4'b0000;
														assign node8314 = (inp[15]) ? node8318 : node8315;
															assign node8315 = (inp[0]) ? 4'b0100 : 4'b0110;
															assign node8318 = (inp[0]) ? 4'b0110 : 4'b0100;
													assign node8321 = (inp[12]) ? node8329 : node8322;
														assign node8322 = (inp[15]) ? node8326 : node8323;
															assign node8323 = (inp[0]) ? 4'b0100 : 4'b0110;
															assign node8326 = (inp[0]) ? 4'b0110 : 4'b0100;
														assign node8329 = (inp[0]) ? node8333 : node8330;
															assign node8330 = (inp[15]) ? 4'b0000 : 4'b0010;
															assign node8333 = (inp[15]) ? 4'b0010 : 4'b0000;
											assign node8336 = (inp[9]) ? node8376 : node8337;
												assign node8337 = (inp[12]) ? node8355 : node8338;
													assign node8338 = (inp[4]) ? node8346 : node8339;
														assign node8339 = (inp[15]) ? node8343 : node8340;
															assign node8340 = (inp[0]) ? 4'b0100 : 4'b0110;
															assign node8343 = (inp[0]) ? 4'b0110 : 4'b0100;
														assign node8346 = (inp[14]) ? node8352 : node8347;
															assign node8347 = (inp[0]) ? 4'b0010 : node8348;
																assign node8348 = (inp[15]) ? 4'b0000 : 4'b0010;
															assign node8352 = (inp[15]) ? 4'b0010 : 4'b0000;
													assign node8355 = (inp[4]) ? node8363 : node8356;
														assign node8356 = (inp[14]) ? 4'b0010 : node8357;
															assign node8357 = (inp[15]) ? node8359 : 4'b0010;
																assign node8359 = (inp[0]) ? 4'b0010 : 4'b0000;
														assign node8363 = (inp[14]) ? node8371 : node8364;
															assign node8364 = (inp[0]) ? node8368 : node8365;
																assign node8365 = (inp[15]) ? 4'b0110 : 4'b0100;
																assign node8368 = (inp[15]) ? 4'b0100 : 4'b0110;
															assign node8371 = (inp[0]) ? node8373 : 4'b0110;
																assign node8373 = (inp[15]) ? 4'b0100 : 4'b0110;
												assign node8376 = (inp[14]) ? node8404 : node8377;
													assign node8377 = (inp[15]) ? node8391 : node8378;
														assign node8378 = (inp[0]) ? node8384 : node8379;
															assign node8379 = (inp[4]) ? node8381 : 4'b0100;
																assign node8381 = (inp[12]) ? 4'b0000 : 4'b0100;
															assign node8384 = (inp[12]) ? node8388 : node8385;
																assign node8385 = (inp[4]) ? 4'b0110 : 4'b0000;
																assign node8388 = (inp[4]) ? 4'b0010 : 4'b0110;
														assign node8391 = (inp[0]) ? node8399 : node8392;
															assign node8392 = (inp[4]) ? node8396 : node8393;
																assign node8393 = (inp[12]) ? 4'b0110 : 4'b0000;
																assign node8396 = (inp[12]) ? 4'b0010 : 4'b0110;
															assign node8399 = (inp[4]) ? 4'b0100 : node8400;
																assign node8400 = (inp[12]) ? 4'b0100 : 4'b0010;
													assign node8404 = (inp[0]) ? node8414 : node8405;
														assign node8405 = (inp[15]) ? 4'b0010 : node8406;
															assign node8406 = (inp[4]) ? node8410 : node8407;
																assign node8407 = (inp[12]) ? 4'b0100 : 4'b0010;
																assign node8410 = (inp[12]) ? 4'b0000 : 4'b0100;
														assign node8414 = (inp[12]) ? node8418 : node8415;
															assign node8415 = (inp[4]) ? 4'b0100 : 4'b0000;
															assign node8418 = (inp[15]) ? 4'b0100 : 4'b0110;
									assign node8421 = (inp[10]) ? node8507 : node8422;
										assign node8422 = (inp[0]) ? node8462 : node8423;
											assign node8423 = (inp[15]) ? node8447 : node8424;
												assign node8424 = (inp[5]) ? node8440 : node8425;
													assign node8425 = (inp[12]) ? node8433 : node8426;
														assign node8426 = (inp[4]) ? node8430 : node8427;
															assign node8427 = (inp[9]) ? 4'b0010 : 4'b0110;
															assign node8430 = (inp[9]) ? 4'b0100 : 4'b0010;
														assign node8433 = (inp[14]) ? node8435 : 4'b0010;
															assign node8435 = (inp[9]) ? 4'b0010 : node8436;
																assign node8436 = (inp[4]) ? 4'b0010 : 4'b0110;
													assign node8440 = (inp[4]) ? node8444 : node8441;
														assign node8441 = (inp[9]) ? 4'b0000 : 4'b0100;
														assign node8444 = (inp[9]) ? 4'b0100 : 4'b0000;
												assign node8447 = (inp[5]) ? node8455 : node8448;
													assign node8448 = (inp[9]) ? node8452 : node8449;
														assign node8449 = (inp[4]) ? 4'b0000 : 4'b0100;
														assign node8452 = (inp[4]) ? 4'b0110 : 4'b0000;
													assign node8455 = (inp[9]) ? node8459 : node8456;
														assign node8456 = (inp[4]) ? 4'b0010 : 4'b0110;
														assign node8459 = (inp[4]) ? 4'b0110 : 4'b0010;
											assign node8462 = (inp[15]) ? node8484 : node8463;
												assign node8463 = (inp[5]) ? node8471 : node8464;
													assign node8464 = (inp[4]) ? node8468 : node8465;
														assign node8465 = (inp[9]) ? 4'b0000 : 4'b0100;
														assign node8468 = (inp[9]) ? 4'b0110 : 4'b0000;
													assign node8471 = (inp[12]) ? node8479 : node8472;
														assign node8472 = (inp[4]) ? node8476 : node8473;
															assign node8473 = (inp[9]) ? 4'b0010 : 4'b0110;
															assign node8476 = (inp[9]) ? 4'b0110 : 4'b0010;
														assign node8479 = (inp[4]) ? 4'b0010 : node8480;
															assign node8480 = (inp[9]) ? 4'b0010 : 4'b0110;
												assign node8484 = (inp[5]) ? node8492 : node8485;
													assign node8485 = (inp[9]) ? node8489 : node8486;
														assign node8486 = (inp[4]) ? 4'b0010 : 4'b0110;
														assign node8489 = (inp[4]) ? 4'b0100 : 4'b0010;
													assign node8492 = (inp[12]) ? node8498 : node8493;
														assign node8493 = (inp[4]) ? 4'b0000 : node8494;
															assign node8494 = (inp[9]) ? 4'b0000 : 4'b0100;
														assign node8498 = (inp[14]) ? node8500 : 4'b0100;
															assign node8500 = (inp[4]) ? node8504 : node8501;
																assign node8501 = (inp[9]) ? 4'b0000 : 4'b0100;
																assign node8504 = (inp[9]) ? 4'b0100 : 4'b0000;
										assign node8507 = (inp[12]) ? node8573 : node8508;
											assign node8508 = (inp[15]) ? node8540 : node8509;
												assign node8509 = (inp[0]) ? node8525 : node8510;
													assign node8510 = (inp[5]) ? node8518 : node8511;
														assign node8511 = (inp[9]) ? node8515 : node8512;
															assign node8512 = (inp[4]) ? 4'b0010 : 4'b0110;
															assign node8515 = (inp[4]) ? 4'b0100 : 4'b0010;
														assign node8518 = (inp[9]) ? node8522 : node8519;
															assign node8519 = (inp[4]) ? 4'b0000 : 4'b0100;
															assign node8522 = (inp[4]) ? 4'b0100 : 4'b0000;
													assign node8525 = (inp[5]) ? node8533 : node8526;
														assign node8526 = (inp[4]) ? node8530 : node8527;
															assign node8527 = (inp[9]) ? 4'b0000 : 4'b0100;
															assign node8530 = (inp[9]) ? 4'b0110 : 4'b0000;
														assign node8533 = (inp[4]) ? node8537 : node8534;
															assign node8534 = (inp[9]) ? 4'b0010 : 4'b0110;
															assign node8537 = (inp[9]) ? 4'b0110 : 4'b0010;
												assign node8540 = (inp[0]) ? node8556 : node8541;
													assign node8541 = (inp[5]) ? node8549 : node8542;
														assign node8542 = (inp[4]) ? node8546 : node8543;
															assign node8543 = (inp[9]) ? 4'b0000 : 4'b0100;
															assign node8546 = (inp[9]) ? 4'b0110 : 4'b0000;
														assign node8549 = (inp[4]) ? node8553 : node8550;
															assign node8550 = (inp[9]) ? 4'b0010 : 4'b0110;
															assign node8553 = (inp[9]) ? 4'b0110 : 4'b0010;
													assign node8556 = (inp[5]) ? node8566 : node8557;
														assign node8557 = (inp[14]) ? node8559 : 4'b0010;
															assign node8559 = (inp[9]) ? node8563 : node8560;
																assign node8560 = (inp[4]) ? 4'b0010 : 4'b0110;
																assign node8563 = (inp[4]) ? 4'b0100 : 4'b0010;
														assign node8566 = (inp[9]) ? node8570 : node8567;
															assign node8567 = (inp[4]) ? 4'b0000 : 4'b0100;
															assign node8570 = (inp[4]) ? 4'b0100 : 4'b0000;
											assign node8573 = (inp[4]) ? node8595 : node8574;
												assign node8574 = (inp[9]) ? node8588 : node8575;
													assign node8575 = (inp[5]) ? node8583 : node8576;
														assign node8576 = (inp[15]) ? node8580 : node8577;
															assign node8577 = (inp[0]) ? 4'b0000 : 4'b0010;
															assign node8580 = (inp[0]) ? 4'b0010 : 4'b0000;
														assign node8583 = (inp[0]) ? 4'b0000 : node8584;
															assign node8584 = (inp[15]) ? 4'b0010 : 4'b0000;
													assign node8588 = (inp[15]) ? node8592 : node8589;
														assign node8589 = (inp[0]) ? 4'b0110 : 4'b0100;
														assign node8592 = (inp[0]) ? 4'b0100 : 4'b0110;
												assign node8595 = (inp[9]) ? node8611 : node8596;
													assign node8596 = (inp[14]) ? node8602 : node8597;
														assign node8597 = (inp[5]) ? 4'b0110 : node8598;
															assign node8598 = (inp[0]) ? 4'b0100 : 4'b0110;
														assign node8602 = (inp[5]) ? 4'b0100 : node8603;
															assign node8603 = (inp[0]) ? node8607 : node8604;
																assign node8604 = (inp[15]) ? 4'b0110 : 4'b0100;
																assign node8607 = (inp[15]) ? 4'b0100 : 4'b0110;
													assign node8611 = (inp[14]) ? node8619 : node8612;
														assign node8612 = (inp[0]) ? node8616 : node8613;
															assign node8613 = (inp[15]) ? 4'b0010 : 4'b0000;
															assign node8616 = (inp[15]) ? 4'b0000 : 4'b0010;
														assign node8619 = (inp[5]) ? node8625 : node8620;
															assign node8620 = (inp[0]) ? 4'b0000 : node8621;
																assign node8621 = (inp[15]) ? 4'b0010 : 4'b0000;
															assign node8625 = (inp[15]) ? 4'b0000 : node8626;
																assign node8626 = (inp[0]) ? 4'b0010 : 4'b0000;
				assign node8630 = (inp[1]) ? node12452 : node8631;
					assign node8631 = (inp[7]) ? node10527 : node8632;
						assign node8632 = (inp[8]) ? node9564 : node8633;
							assign node8633 = (inp[2]) ? node9203 : node8634;
								assign node8634 = (inp[14]) ? node8924 : node8635;
									assign node8635 = (inp[12]) ? node8781 : node8636;
										assign node8636 = (inp[10]) ? node8712 : node8637;
											assign node8637 = (inp[3]) ? node8669 : node8638;
												assign node8638 = (inp[4]) ? node8650 : node8639;
													assign node8639 = (inp[9]) ? node8645 : node8640;
														assign node8640 = (inp[5]) ? 4'b1111 : node8641;
															assign node8641 = (inp[15]) ? 4'b1111 : 4'b1101;
														assign node8645 = (inp[0]) ? node8647 : 4'b1011;
															assign node8647 = (inp[15]) ? 4'b1011 : 4'b1001;
													assign node8650 = (inp[9]) ? node8656 : node8651;
														assign node8651 = (inp[0]) ? node8653 : 4'b1001;
															assign node8653 = (inp[15]) ? 4'b1011 : 4'b1001;
														assign node8656 = (inp[15]) ? node8662 : node8657;
															assign node8657 = (inp[5]) ? node8659 : 4'b1101;
																assign node8659 = (inp[0]) ? 4'b1111 : 4'b1101;
															assign node8662 = (inp[5]) ? node8666 : node8663;
																assign node8663 = (inp[0]) ? 4'b1111 : 4'b1101;
																assign node8666 = (inp[0]) ? 4'b1101 : 4'b1111;
												assign node8669 = (inp[15]) ? node8691 : node8670;
													assign node8670 = (inp[0]) ? node8678 : node8671;
														assign node8671 = (inp[5]) ? 4'b1001 : node8672;
															assign node8672 = (inp[9]) ? 4'b1011 : node8673;
																assign node8673 = (inp[4]) ? 4'b1011 : 4'b1111;
														assign node8678 = (inp[5]) ? node8684 : node8679;
															assign node8679 = (inp[4]) ? node8681 : 4'b1001;
																assign node8681 = (inp[9]) ? 4'b1111 : 4'b1001;
															assign node8684 = (inp[4]) ? node8688 : node8685;
																assign node8685 = (inp[9]) ? 4'b1011 : 4'b1111;
																assign node8688 = (inp[9]) ? 4'b1111 : 4'b1011;
													assign node8691 = (inp[0]) ? node8705 : node8692;
														assign node8692 = (inp[5]) ? node8698 : node8693;
															assign node8693 = (inp[9]) ? 4'b1001 : node8694;
																assign node8694 = (inp[4]) ? 4'b1001 : 4'b1101;
															assign node8698 = (inp[9]) ? node8702 : node8699;
																assign node8699 = (inp[4]) ? 4'b1011 : 4'b1111;
																assign node8702 = (inp[4]) ? 4'b1111 : 4'b1011;
														assign node8705 = (inp[5]) ? 4'b1001 : node8706;
															assign node8706 = (inp[9]) ? 4'b1011 : node8707;
																assign node8707 = (inp[4]) ? 4'b1011 : 4'b1111;
											assign node8712 = (inp[4]) ? node8744 : node8713;
												assign node8713 = (inp[9]) ? node8729 : node8714;
													assign node8714 = (inp[15]) ? node8722 : node8715;
														assign node8715 = (inp[0]) ? node8717 : 4'b1111;
															assign node8717 = (inp[3]) ? node8719 : 4'b1101;
																assign node8719 = (inp[5]) ? 4'b1111 : 4'b1101;
														assign node8722 = (inp[0]) ? node8724 : 4'b1101;
															assign node8724 = (inp[3]) ? node8726 : 4'b1111;
																assign node8726 = (inp[5]) ? 4'b1101 : 4'b1111;
													assign node8729 = (inp[0]) ? node8737 : node8730;
														assign node8730 = (inp[15]) ? node8734 : node8731;
															assign node8731 = (inp[3]) ? 4'b1001 : 4'b1011;
															assign node8734 = (inp[3]) ? 4'b1011 : 4'b1001;
														assign node8737 = (inp[5]) ? node8739 : 4'b1001;
															assign node8739 = (inp[3]) ? node8741 : 4'b1001;
																assign node8741 = (inp[15]) ? 4'b1001 : 4'b1011;
												assign node8744 = (inp[9]) ? node8756 : node8745;
													assign node8745 = (inp[0]) ? node8747 : 4'b1011;
														assign node8747 = (inp[15]) ? node8751 : node8748;
															assign node8748 = (inp[3]) ? 4'b1011 : 4'b1001;
															assign node8751 = (inp[5]) ? node8753 : 4'b1011;
																assign node8753 = (inp[3]) ? 4'b1001 : 4'b1011;
													assign node8756 = (inp[3]) ? node8766 : node8757;
														assign node8757 = (inp[15]) ? 4'b1111 : node8758;
															assign node8758 = (inp[0]) ? node8762 : node8759;
																assign node8759 = (inp[5]) ? 4'b1101 : 4'b1111;
																assign node8762 = (inp[5]) ? 4'b1111 : 4'b1101;
														assign node8766 = (inp[5]) ? node8774 : node8767;
															assign node8767 = (inp[15]) ? node8771 : node8768;
																assign node8768 = (inp[0]) ? 4'b1111 : 4'b1101;
																assign node8771 = (inp[0]) ? 4'b1101 : 4'b1111;
															assign node8774 = (inp[0]) ? node8778 : node8775;
																assign node8775 = (inp[15]) ? 4'b1111 : 4'b1101;
																assign node8778 = (inp[15]) ? 4'b1101 : 4'b1111;
										assign node8781 = (inp[3]) ? node8843 : node8782;
											assign node8782 = (inp[15]) ? node8814 : node8783;
												assign node8783 = (inp[0]) ? node8801 : node8784;
													assign node8784 = (inp[5]) ? node8790 : node8785;
														assign node8785 = (inp[4]) ? node8787 : 4'b1111;
															assign node8787 = (inp[9]) ? 4'b1111 : 4'b1011;
														assign node8790 = (inp[4]) ? node8796 : node8791;
															assign node8791 = (inp[9]) ? node8793 : 4'b1011;
																assign node8793 = (inp[10]) ? 4'b1101 : 4'b1011;
															assign node8796 = (inp[10]) ? node8798 : 4'b1101;
																assign node8798 = (inp[9]) ? 4'b1001 : 4'b1101;
													assign node8801 = (inp[9]) ? node8809 : node8802;
														assign node8802 = (inp[10]) ? node8806 : node8803;
															assign node8803 = (inp[4]) ? 4'b1001 : 4'b1101;
															assign node8806 = (inp[4]) ? 4'b1111 : 4'b1001;
														assign node8809 = (inp[10]) ? node8811 : 4'b1001;
															assign node8811 = (inp[5]) ? 4'b1011 : 4'b1001;
												assign node8814 = (inp[0]) ? node8828 : node8815;
													assign node8815 = (inp[9]) ? node8821 : node8816;
														assign node8816 = (inp[4]) ? 4'b1001 : node8817;
															assign node8817 = (inp[10]) ? 4'b1001 : 4'b1101;
														assign node8821 = (inp[4]) ? 4'b1111 : node8822;
															assign node8822 = (inp[10]) ? node8824 : 4'b1001;
																assign node8824 = (inp[5]) ? 4'b1111 : 4'b1101;
													assign node8828 = (inp[5]) ? node8836 : node8829;
														assign node8829 = (inp[9]) ? node8831 : 4'b1111;
															assign node8831 = (inp[4]) ? 4'b1011 : node8832;
																assign node8832 = (inp[10]) ? 4'b1111 : 4'b1011;
														assign node8836 = (inp[4]) ? node8838 : 4'b1011;
															assign node8838 = (inp[9]) ? 4'b1101 : node8839;
																assign node8839 = (inp[10]) ? 4'b1101 : 4'b1011;
											assign node8843 = (inp[15]) ? node8875 : node8844;
												assign node8844 = (inp[0]) ? node8856 : node8845;
													assign node8845 = (inp[10]) ? node8847 : 4'b1011;
														assign node8847 = (inp[4]) ? node8853 : node8848;
															assign node8848 = (inp[9]) ? 4'b1101 : node8849;
																assign node8849 = (inp[5]) ? 4'b1001 : 4'b1011;
															assign node8853 = (inp[9]) ? 4'b1001 : 4'b1101;
													assign node8856 = (inp[10]) ? node8868 : node8857;
														assign node8857 = (inp[5]) ? node8865 : node8858;
															assign node8858 = (inp[9]) ? node8862 : node8859;
																assign node8859 = (inp[4]) ? 4'b1001 : 4'b1101;
																assign node8862 = (inp[4]) ? 4'b1111 : 4'b1001;
															assign node8865 = (inp[4]) ? 4'b1111 : 4'b1011;
														assign node8868 = (inp[9]) ? node8872 : node8869;
															assign node8869 = (inp[4]) ? 4'b1111 : 4'b1011;
															assign node8872 = (inp[4]) ? 4'b1011 : 4'b1111;
												assign node8875 = (inp[0]) ? node8897 : node8876;
													assign node8876 = (inp[5]) ? node8888 : node8877;
														assign node8877 = (inp[9]) ? node8883 : node8878;
															assign node8878 = (inp[10]) ? 4'b1001 : node8879;
																assign node8879 = (inp[4]) ? 4'b1001 : 4'b1101;
															assign node8883 = (inp[4]) ? node8885 : 4'b1001;
																assign node8885 = (inp[10]) ? 4'b1011 : 4'b1111;
														assign node8888 = (inp[9]) ? 4'b1111 : node8889;
															assign node8889 = (inp[4]) ? node8893 : node8890;
																assign node8890 = (inp[10]) ? 4'b1011 : 4'b1111;
																assign node8893 = (inp[10]) ? 4'b1111 : 4'b1011;
													assign node8897 = (inp[5]) ? node8909 : node8898;
														assign node8898 = (inp[10]) ? node8904 : node8899;
															assign node8899 = (inp[4]) ? node8901 : 4'b1011;
																assign node8901 = (inp[9]) ? 4'b1101 : 4'b1011;
															assign node8904 = (inp[9]) ? 4'b1101 : node8905;
																assign node8905 = (inp[4]) ? 4'b1101 : 4'b1011;
														assign node8909 = (inp[9]) ? node8917 : node8910;
															assign node8910 = (inp[10]) ? node8914 : node8911;
																assign node8911 = (inp[4]) ? 4'b1001 : 4'b1101;
																assign node8914 = (inp[4]) ? 4'b1101 : 4'b1001;
															assign node8917 = (inp[10]) ? node8921 : node8918;
																assign node8918 = (inp[4]) ? 4'b1101 : 4'b1001;
																assign node8921 = (inp[4]) ? 4'b1001 : 4'b1101;
									assign node8924 = (inp[10]) ? node9056 : node8925;
										assign node8925 = (inp[15]) ? node9017 : node8926;
											assign node8926 = (inp[0]) ? node8972 : node8927;
												assign node8927 = (inp[3]) ? node8951 : node8928;
													assign node8928 = (inp[12]) ? node8942 : node8929;
														assign node8929 = (inp[5]) ? node8937 : node8930;
															assign node8930 = (inp[4]) ? node8934 : node8931;
																assign node8931 = (inp[9]) ? 4'b1010 : 4'b1110;
																assign node8934 = (inp[9]) ? 4'b1110 : 4'b1010;
															assign node8937 = (inp[4]) ? 4'b1010 : node8938;
																assign node8938 = (inp[9]) ? 4'b1010 : 4'b1110;
														assign node8942 = (inp[9]) ? node8946 : node8943;
															assign node8943 = (inp[4]) ? 4'b1010 : 4'b1110;
															assign node8946 = (inp[4]) ? node8948 : 4'b1010;
																assign node8948 = (inp[5]) ? 4'b1100 : 4'b1110;
													assign node8951 = (inp[5]) ? node8959 : node8952;
														assign node8952 = (inp[4]) ? node8956 : node8953;
															assign node8953 = (inp[9]) ? 4'b1010 : 4'b1110;
															assign node8956 = (inp[9]) ? 4'b1100 : 4'b1010;
														assign node8959 = (inp[12]) ? node8965 : node8960;
															assign node8960 = (inp[4]) ? node8962 : 4'b1100;
																assign node8962 = (inp[9]) ? 4'b1100 : 4'b1000;
															assign node8965 = (inp[4]) ? node8969 : node8966;
																assign node8966 = (inp[9]) ? 4'b1000 : 4'b1100;
																assign node8969 = (inp[9]) ? 4'b1100 : 4'b1000;
												assign node8972 = (inp[5]) ? node8996 : node8973;
													assign node8973 = (inp[3]) ? node8989 : node8974;
														assign node8974 = (inp[12]) ? node8982 : node8975;
															assign node8975 = (inp[4]) ? node8979 : node8976;
																assign node8976 = (inp[9]) ? 4'b1000 : 4'b1100;
																assign node8979 = (inp[9]) ? 4'b1100 : 4'b1000;
															assign node8982 = (inp[9]) ? node8986 : node8983;
																assign node8983 = (inp[4]) ? 4'b1000 : 4'b1100;
																assign node8986 = (inp[4]) ? 4'b1100 : 4'b1000;
														assign node8989 = (inp[9]) ? node8993 : node8990;
															assign node8990 = (inp[4]) ? 4'b1000 : 4'b1100;
															assign node8993 = (inp[4]) ? 4'b1110 : 4'b1000;
													assign node8996 = (inp[3]) ? node9004 : node8997;
														assign node8997 = (inp[4]) ? node9001 : node8998;
															assign node8998 = (inp[9]) ? 4'b1000 : 4'b1100;
															assign node9001 = (inp[9]) ? 4'b1110 : 4'b1000;
														assign node9004 = (inp[12]) ? node9010 : node9005;
															assign node9005 = (inp[9]) ? node9007 : 4'b1110;
																assign node9007 = (inp[4]) ? 4'b1110 : 4'b1010;
															assign node9010 = (inp[4]) ? node9014 : node9011;
																assign node9011 = (inp[9]) ? 4'b1010 : 4'b1110;
																assign node9014 = (inp[9]) ? 4'b1110 : 4'b1010;
											assign node9017 = (inp[0]) ? node9037 : node9018;
												assign node9018 = (inp[3]) ? node9024 : node9019;
													assign node9019 = (inp[9]) ? 4'b1000 : node9020;
														assign node9020 = (inp[4]) ? 4'b1000 : 4'b1100;
													assign node9024 = (inp[5]) ? node9030 : node9025;
														assign node9025 = (inp[9]) ? 4'b1110 : node9026;
															assign node9026 = (inp[4]) ? 4'b1000 : 4'b1100;
														assign node9030 = (inp[4]) ? node9034 : node9031;
															assign node9031 = (inp[9]) ? 4'b1010 : 4'b1110;
															assign node9034 = (inp[9]) ? 4'b1110 : 4'b1010;
												assign node9037 = (inp[4]) ? node9045 : node9038;
													assign node9038 = (inp[9]) ? 4'b1010 : node9039;
														assign node9039 = (inp[5]) ? node9041 : 4'b1110;
															assign node9041 = (inp[3]) ? 4'b1100 : 4'b1110;
													assign node9045 = (inp[9]) ? node9051 : node9046;
														assign node9046 = (inp[3]) ? node9048 : 4'b1010;
															assign node9048 = (inp[5]) ? 4'b1000 : 4'b1010;
														assign node9051 = (inp[5]) ? 4'b1100 : node9052;
															assign node9052 = (inp[3]) ? 4'b1100 : 4'b1110;
										assign node9056 = (inp[4]) ? node9136 : node9057;
											assign node9057 = (inp[12]) ? node9097 : node9058;
												assign node9058 = (inp[9]) ? node9074 : node9059;
													assign node9059 = (inp[5]) ? node9065 : node9060;
														assign node9060 = (inp[3]) ? 4'b1110 : node9061;
															assign node9061 = (inp[0]) ? 4'b1110 : 4'b1100;
														assign node9065 = (inp[15]) ? 4'b1100 : node9066;
															assign node9066 = (inp[0]) ? node9070 : node9067;
																assign node9067 = (inp[3]) ? 4'b1100 : 4'b1110;
																assign node9070 = (inp[3]) ? 4'b1110 : 4'b1100;
													assign node9074 = (inp[15]) ? node9086 : node9075;
														assign node9075 = (inp[0]) ? node9081 : node9076;
															assign node9076 = (inp[5]) ? node9078 : 4'b1010;
																assign node9078 = (inp[3]) ? 4'b1000 : 4'b1010;
															assign node9081 = (inp[3]) ? node9083 : 4'b1000;
																assign node9083 = (inp[5]) ? 4'b1010 : 4'b1000;
														assign node9086 = (inp[0]) ? node9092 : node9087;
															assign node9087 = (inp[3]) ? node9089 : 4'b1000;
																assign node9089 = (inp[5]) ? 4'b1010 : 4'b1000;
															assign node9092 = (inp[3]) ? node9094 : 4'b1010;
																assign node9094 = (inp[5]) ? 4'b1000 : 4'b1010;
												assign node9097 = (inp[9]) ? node9119 : node9098;
													assign node9098 = (inp[3]) ? node9108 : node9099;
														assign node9099 = (inp[5]) ? node9101 : 4'b1010;
															assign node9101 = (inp[15]) ? node9105 : node9102;
																assign node9102 = (inp[0]) ? 4'b1000 : 4'b1010;
																assign node9105 = (inp[0]) ? 4'b1010 : 4'b1000;
														assign node9108 = (inp[5]) ? node9114 : node9109;
															assign node9109 = (inp[0]) ? node9111 : 4'b1000;
																assign node9111 = (inp[15]) ? 4'b1010 : 4'b1000;
															assign node9114 = (inp[15]) ? node9116 : 4'b1010;
																assign node9116 = (inp[0]) ? 4'b1000 : 4'b1010;
													assign node9119 = (inp[0]) ? node9127 : node9120;
														assign node9120 = (inp[15]) ? node9124 : node9121;
															assign node9121 = (inp[3]) ? 4'b1100 : 4'b1110;
															assign node9124 = (inp[3]) ? 4'b1110 : 4'b1100;
														assign node9127 = (inp[15]) ? node9133 : node9128;
															assign node9128 = (inp[3]) ? 4'b1110 : node9129;
																assign node9129 = (inp[5]) ? 4'b1110 : 4'b1100;
															assign node9133 = (inp[3]) ? 4'b1100 : 4'b1110;
											assign node9136 = (inp[5]) ? node9172 : node9137;
												assign node9137 = (inp[15]) ? node9155 : node9138;
													assign node9138 = (inp[9]) ? node9144 : node9139;
														assign node9139 = (inp[12]) ? 4'b1110 : node9140;
															assign node9140 = (inp[0]) ? 4'b1000 : 4'b1010;
														assign node9144 = (inp[12]) ? node9150 : node9145;
															assign node9145 = (inp[0]) ? 4'b1100 : node9146;
																assign node9146 = (inp[3]) ? 4'b1100 : 4'b1110;
															assign node9150 = (inp[0]) ? node9152 : 4'b1000;
																assign node9152 = (inp[3]) ? 4'b1010 : 4'b1000;
													assign node9155 = (inp[3]) ? node9163 : node9156;
														assign node9156 = (inp[0]) ? node9158 : 4'b1100;
															assign node9158 = (inp[9]) ? 4'b1110 : node9159;
																assign node9159 = (inp[12]) ? 4'b1110 : 4'b1010;
														assign node9163 = (inp[0]) ? node9167 : node9164;
															assign node9164 = (inp[9]) ? 4'b1110 : 4'b1000;
															assign node9167 = (inp[9]) ? node9169 : 4'b1100;
																assign node9169 = (inp[12]) ? 4'b1000 : 4'b1100;
												assign node9172 = (inp[15]) ? node9192 : node9173;
													assign node9173 = (inp[0]) ? node9185 : node9174;
														assign node9174 = (inp[3]) ? node9180 : node9175;
															assign node9175 = (inp[9]) ? node9177 : 4'b1100;
																assign node9177 = (inp[12]) ? 4'b1000 : 4'b1100;
															assign node9180 = (inp[12]) ? 4'b1100 : node9181;
																assign node9181 = (inp[9]) ? 4'b1100 : 4'b1000;
														assign node9185 = (inp[9]) ? node9189 : node9186;
															assign node9186 = (inp[12]) ? 4'b1110 : 4'b1010;
															assign node9189 = (inp[12]) ? 4'b1010 : 4'b1110;
													assign node9192 = (inp[0]) ? node9194 : 4'b1010;
														assign node9194 = (inp[9]) ? node9200 : node9195;
															assign node9195 = (inp[12]) ? 4'b1100 : node9196;
																assign node9196 = (inp[3]) ? 4'b1000 : 4'b1010;
															assign node9200 = (inp[12]) ? 4'b1000 : 4'b1100;
								assign node9203 = (inp[9]) ? node9383 : node9204;
									assign node9204 = (inp[4]) ? node9286 : node9205;
										assign node9205 = (inp[10]) ? node9229 : node9206;
											assign node9206 = (inp[15]) ? node9218 : node9207;
												assign node9207 = (inp[0]) ? node9213 : node9208;
													assign node9208 = (inp[5]) ? node9210 : 4'b1110;
														assign node9210 = (inp[3]) ? 4'b1100 : 4'b1110;
													assign node9213 = (inp[3]) ? node9215 : 4'b1100;
														assign node9215 = (inp[5]) ? 4'b1110 : 4'b1100;
												assign node9218 = (inp[0]) ? node9224 : node9219;
													assign node9219 = (inp[5]) ? node9221 : 4'b1100;
														assign node9221 = (inp[3]) ? 4'b1110 : 4'b1100;
													assign node9224 = (inp[5]) ? node9226 : 4'b1110;
														assign node9226 = (inp[3]) ? 4'b1100 : 4'b1110;
											assign node9229 = (inp[12]) ? node9263 : node9230;
												assign node9230 = (inp[5]) ? node9238 : node9231;
													assign node9231 = (inp[0]) ? node9235 : node9232;
														assign node9232 = (inp[15]) ? 4'b1100 : 4'b1110;
														assign node9235 = (inp[15]) ? 4'b1110 : 4'b1100;
													assign node9238 = (inp[0]) ? node9248 : node9239;
														assign node9239 = (inp[14]) ? node9245 : node9240;
															assign node9240 = (inp[3]) ? node9242 : 4'b1110;
																assign node9242 = (inp[15]) ? 4'b1110 : 4'b1100;
															assign node9245 = (inp[3]) ? 4'b1110 : 4'b1100;
														assign node9248 = (inp[14]) ? node9256 : node9249;
															assign node9249 = (inp[15]) ? node9253 : node9250;
																assign node9250 = (inp[3]) ? 4'b1110 : 4'b1100;
																assign node9253 = (inp[3]) ? 4'b1100 : 4'b1110;
															assign node9256 = (inp[15]) ? node9260 : node9257;
																assign node9257 = (inp[3]) ? 4'b1110 : 4'b1100;
																assign node9260 = (inp[3]) ? 4'b1100 : 4'b1110;
												assign node9263 = (inp[3]) ? node9273 : node9264;
													assign node9264 = (inp[14]) ? 4'b1010 : node9265;
														assign node9265 = (inp[0]) ? node9269 : node9266;
															assign node9266 = (inp[15]) ? 4'b1000 : 4'b1010;
															assign node9269 = (inp[15]) ? 4'b1010 : 4'b1000;
													assign node9273 = (inp[15]) ? node9283 : node9274;
														assign node9274 = (inp[14]) ? node9276 : 4'b1010;
															assign node9276 = (inp[5]) ? node9280 : node9277;
																assign node9277 = (inp[0]) ? 4'b1000 : 4'b1010;
																assign node9280 = (inp[0]) ? 4'b1010 : 4'b1000;
														assign node9283 = (inp[5]) ? 4'b1010 : 4'b1000;
										assign node9286 = (inp[10]) ? node9326 : node9287;
											assign node9287 = (inp[3]) ? node9295 : node9288;
												assign node9288 = (inp[0]) ? node9292 : node9289;
													assign node9289 = (inp[15]) ? 4'b1000 : 4'b1010;
													assign node9292 = (inp[15]) ? 4'b1010 : 4'b1000;
												assign node9295 = (inp[12]) ? node9307 : node9296;
													assign node9296 = (inp[5]) ? node9302 : node9297;
														assign node9297 = (inp[0]) ? node9299 : 4'b1000;
															assign node9299 = (inp[15]) ? 4'b1010 : 4'b1000;
														assign node9302 = (inp[0]) ? 4'b1010 : node9303;
															assign node9303 = (inp[15]) ? 4'b1010 : 4'b1000;
													assign node9307 = (inp[0]) ? node9321 : node9308;
														assign node9308 = (inp[14]) ? node9316 : node9309;
															assign node9309 = (inp[15]) ? node9313 : node9310;
																assign node9310 = (inp[5]) ? 4'b1000 : 4'b1010;
																assign node9313 = (inp[5]) ? 4'b1010 : 4'b1000;
															assign node9316 = (inp[15]) ? node9318 : 4'b1010;
																assign node9318 = (inp[5]) ? 4'b1010 : 4'b1000;
														assign node9321 = (inp[5]) ? 4'b1000 : node9322;
															assign node9322 = (inp[15]) ? 4'b1010 : 4'b1000;
											assign node9326 = (inp[12]) ? node9352 : node9327;
												assign node9327 = (inp[5]) ? node9335 : node9328;
													assign node9328 = (inp[0]) ? node9332 : node9329;
														assign node9329 = (inp[15]) ? 4'b1000 : 4'b1010;
														assign node9332 = (inp[15]) ? 4'b1010 : 4'b1000;
													assign node9335 = (inp[0]) ? node9343 : node9336;
														assign node9336 = (inp[14]) ? 4'b1010 : node9337;
															assign node9337 = (inp[3]) ? node9339 : 4'b1000;
																assign node9339 = (inp[15]) ? 4'b1010 : 4'b1000;
														assign node9343 = (inp[14]) ? 4'b1000 : node9344;
															assign node9344 = (inp[3]) ? node9348 : node9345;
																assign node9345 = (inp[15]) ? 4'b1010 : 4'b1000;
																assign node9348 = (inp[15]) ? 4'b1000 : 4'b1010;
												assign node9352 = (inp[5]) ? node9376 : node9353;
													assign node9353 = (inp[15]) ? node9361 : node9354;
														assign node9354 = (inp[0]) ? node9358 : node9355;
															assign node9355 = (inp[3]) ? 4'b1100 : 4'b1110;
															assign node9358 = (inp[3]) ? 4'b1110 : 4'b1100;
														assign node9361 = (inp[14]) ? node9369 : node9362;
															assign node9362 = (inp[0]) ? node9366 : node9363;
																assign node9363 = (inp[3]) ? 4'b1110 : 4'b1100;
																assign node9366 = (inp[3]) ? 4'b1100 : 4'b1110;
															assign node9369 = (inp[0]) ? node9373 : node9370;
																assign node9370 = (inp[3]) ? 4'b1110 : 4'b1100;
																assign node9373 = (inp[3]) ? 4'b1100 : 4'b1110;
													assign node9376 = (inp[15]) ? node9380 : node9377;
														assign node9377 = (inp[0]) ? 4'b1110 : 4'b1100;
														assign node9380 = (inp[0]) ? 4'b1100 : 4'b1110;
									assign node9383 = (inp[4]) ? node9475 : node9384;
										assign node9384 = (inp[10]) ? node9418 : node9385;
											assign node9385 = (inp[5]) ? node9393 : node9386;
												assign node9386 = (inp[15]) ? node9390 : node9387;
													assign node9387 = (inp[0]) ? 4'b1000 : 4'b1010;
													assign node9390 = (inp[0]) ? 4'b1010 : 4'b1000;
												assign node9393 = (inp[14]) ? node9409 : node9394;
													assign node9394 = (inp[0]) ? node9402 : node9395;
														assign node9395 = (inp[15]) ? node9399 : node9396;
															assign node9396 = (inp[3]) ? 4'b1000 : 4'b1010;
															assign node9399 = (inp[3]) ? 4'b1010 : 4'b1000;
														assign node9402 = (inp[3]) ? node9406 : node9403;
															assign node9403 = (inp[15]) ? 4'b1010 : 4'b1000;
															assign node9406 = (inp[15]) ? 4'b1000 : 4'b1010;
													assign node9409 = (inp[0]) ? node9411 : 4'b1000;
														assign node9411 = (inp[15]) ? node9415 : node9412;
															assign node9412 = (inp[3]) ? 4'b1010 : 4'b1000;
															assign node9415 = (inp[3]) ? 4'b1000 : 4'b1010;
											assign node9418 = (inp[12]) ? node9446 : node9419;
												assign node9419 = (inp[14]) ? node9435 : node9420;
													assign node9420 = (inp[0]) ? node9432 : node9421;
														assign node9421 = (inp[15]) ? node9427 : node9422;
															assign node9422 = (inp[3]) ? node9424 : 4'b1010;
																assign node9424 = (inp[5]) ? 4'b1000 : 4'b1010;
															assign node9427 = (inp[3]) ? node9429 : 4'b1000;
																assign node9429 = (inp[5]) ? 4'b1010 : 4'b1000;
														assign node9432 = (inp[15]) ? 4'b1010 : 4'b1000;
													assign node9435 = (inp[0]) ? node9437 : 4'b1010;
														assign node9437 = (inp[15]) ? node9441 : node9438;
															assign node9438 = (inp[5]) ? 4'b1010 : 4'b1000;
															assign node9441 = (inp[3]) ? node9443 : 4'b1010;
																assign node9443 = (inp[5]) ? 4'b1000 : 4'b1010;
												assign node9446 = (inp[3]) ? node9462 : node9447;
													assign node9447 = (inp[5]) ? node9455 : node9448;
														assign node9448 = (inp[0]) ? node9452 : node9449;
															assign node9449 = (inp[15]) ? 4'b1100 : 4'b1110;
															assign node9452 = (inp[15]) ? 4'b1110 : 4'b1100;
														assign node9455 = (inp[0]) ? node9459 : node9456;
															assign node9456 = (inp[15]) ? 4'b1110 : 4'b1100;
															assign node9459 = (inp[15]) ? 4'b1100 : 4'b1110;
													assign node9462 = (inp[14]) ? node9470 : node9463;
														assign node9463 = (inp[0]) ? node9467 : node9464;
															assign node9464 = (inp[15]) ? 4'b1110 : 4'b1100;
															assign node9467 = (inp[15]) ? 4'b1100 : 4'b1110;
														assign node9470 = (inp[15]) ? 4'b1110 : node9471;
															assign node9471 = (inp[5]) ? 4'b1110 : 4'b1100;
										assign node9475 = (inp[12]) ? node9523 : node9476;
											assign node9476 = (inp[10]) ? node9500 : node9477;
												assign node9477 = (inp[5]) ? node9493 : node9478;
													assign node9478 = (inp[15]) ? node9486 : node9479;
														assign node9479 = (inp[0]) ? node9483 : node9480;
															assign node9480 = (inp[3]) ? 4'b1100 : 4'b1110;
															assign node9483 = (inp[3]) ? 4'b1110 : 4'b1100;
														assign node9486 = (inp[0]) ? node9490 : node9487;
															assign node9487 = (inp[3]) ? 4'b1110 : 4'b1100;
															assign node9490 = (inp[3]) ? 4'b1100 : 4'b1110;
													assign node9493 = (inp[15]) ? node9497 : node9494;
														assign node9494 = (inp[0]) ? 4'b1110 : 4'b1100;
														assign node9497 = (inp[0]) ? 4'b1100 : 4'b1110;
												assign node9500 = (inp[5]) ? node9516 : node9501;
													assign node9501 = (inp[3]) ? node9503 : 4'b1110;
														assign node9503 = (inp[14]) ? node9509 : node9504;
															assign node9504 = (inp[15]) ? node9506 : 4'b1110;
																assign node9506 = (inp[0]) ? 4'b1100 : 4'b1110;
															assign node9509 = (inp[0]) ? node9513 : node9510;
																assign node9510 = (inp[15]) ? 4'b1110 : 4'b1100;
																assign node9513 = (inp[15]) ? 4'b1100 : 4'b1110;
													assign node9516 = (inp[0]) ? node9520 : node9517;
														assign node9517 = (inp[15]) ? 4'b1110 : 4'b1100;
														assign node9520 = (inp[15]) ? 4'b1100 : 4'b1110;
											assign node9523 = (inp[10]) ? node9545 : node9524;
												assign node9524 = (inp[15]) ? node9534 : node9525;
													assign node9525 = (inp[3]) ? 4'b1100 : node9526;
														assign node9526 = (inp[5]) ? node9530 : node9527;
															assign node9527 = (inp[0]) ? 4'b1100 : 4'b1110;
															assign node9530 = (inp[0]) ? 4'b1110 : 4'b1100;
													assign node9534 = (inp[0]) ? node9540 : node9535;
														assign node9535 = (inp[5]) ? 4'b1110 : node9536;
															assign node9536 = (inp[3]) ? 4'b1110 : 4'b1100;
														assign node9540 = (inp[3]) ? 4'b1100 : node9541;
															assign node9541 = (inp[5]) ? 4'b1100 : 4'b1110;
												assign node9545 = (inp[0]) ? node9557 : node9546;
													assign node9546 = (inp[15]) ? node9552 : node9547;
														assign node9547 = (inp[3]) ? 4'b1000 : node9548;
															assign node9548 = (inp[5]) ? 4'b1000 : 4'b1010;
														assign node9552 = (inp[3]) ? 4'b1010 : node9553;
															assign node9553 = (inp[5]) ? 4'b1010 : 4'b1000;
													assign node9557 = (inp[15]) ? node9559 : 4'b1010;
														assign node9559 = (inp[3]) ? 4'b1000 : node9560;
															assign node9560 = (inp[5]) ? 4'b1000 : 4'b1010;
							assign node9564 = (inp[14]) ? node10124 : node9565;
								assign node9565 = (inp[2]) ? node9827 : node9566;
									assign node9566 = (inp[12]) ? node9672 : node9567;
										assign node9567 = (inp[0]) ? node9619 : node9568;
											assign node9568 = (inp[15]) ? node9594 : node9569;
												assign node9569 = (inp[5]) ? node9579 : node9570;
													assign node9570 = (inp[9]) ? node9574 : node9571;
														assign node9571 = (inp[4]) ? 4'b1010 : 4'b1110;
														assign node9574 = (inp[4]) ? node9576 : 4'b1010;
															assign node9576 = (inp[3]) ? 4'b1100 : 4'b1110;
													assign node9579 = (inp[3]) ? node9587 : node9580;
														assign node9580 = (inp[9]) ? node9584 : node9581;
															assign node9581 = (inp[4]) ? 4'b1010 : 4'b1110;
															assign node9584 = (inp[4]) ? 4'b1100 : 4'b1010;
														assign node9587 = (inp[4]) ? node9591 : node9588;
															assign node9588 = (inp[9]) ? 4'b1000 : 4'b1100;
															assign node9591 = (inp[9]) ? 4'b1100 : 4'b1000;
												assign node9594 = (inp[5]) ? node9604 : node9595;
													assign node9595 = (inp[9]) ? node9599 : node9596;
														assign node9596 = (inp[4]) ? 4'b1000 : 4'b1100;
														assign node9599 = (inp[4]) ? node9601 : 4'b1000;
															assign node9601 = (inp[3]) ? 4'b1110 : 4'b1100;
													assign node9604 = (inp[3]) ? node9612 : node9605;
														assign node9605 = (inp[9]) ? node9609 : node9606;
															assign node9606 = (inp[4]) ? 4'b1000 : 4'b1100;
															assign node9609 = (inp[4]) ? 4'b1110 : 4'b1000;
														assign node9612 = (inp[9]) ? node9616 : node9613;
															assign node9613 = (inp[4]) ? 4'b1010 : 4'b1110;
															assign node9616 = (inp[4]) ? 4'b1110 : 4'b1010;
											assign node9619 = (inp[15]) ? node9647 : node9620;
												assign node9620 = (inp[5]) ? node9630 : node9621;
													assign node9621 = (inp[9]) ? node9625 : node9622;
														assign node9622 = (inp[4]) ? 4'b1000 : 4'b1100;
														assign node9625 = (inp[4]) ? node9627 : 4'b1000;
															assign node9627 = (inp[3]) ? 4'b1110 : 4'b1100;
													assign node9630 = (inp[3]) ? node9638 : node9631;
														assign node9631 = (inp[4]) ? node9635 : node9632;
															assign node9632 = (inp[9]) ? 4'b1000 : 4'b1100;
															assign node9635 = (inp[9]) ? 4'b1110 : 4'b1000;
														assign node9638 = (inp[10]) ? node9640 : 4'b1110;
															assign node9640 = (inp[9]) ? node9644 : node9641;
																assign node9641 = (inp[4]) ? 4'b1010 : 4'b1110;
																assign node9644 = (inp[4]) ? 4'b1110 : 4'b1010;
												assign node9647 = (inp[3]) ? node9657 : node9648;
													assign node9648 = (inp[9]) ? node9652 : node9649;
														assign node9649 = (inp[4]) ? 4'b1010 : 4'b1110;
														assign node9652 = (inp[4]) ? node9654 : 4'b1010;
															assign node9654 = (inp[5]) ? 4'b1100 : 4'b1110;
													assign node9657 = (inp[5]) ? node9665 : node9658;
														assign node9658 = (inp[4]) ? node9662 : node9659;
															assign node9659 = (inp[9]) ? 4'b1010 : 4'b1110;
															assign node9662 = (inp[9]) ? 4'b1100 : 4'b1010;
														assign node9665 = (inp[9]) ? node9669 : node9666;
															assign node9666 = (inp[4]) ? 4'b1000 : 4'b1100;
															assign node9669 = (inp[4]) ? 4'b1100 : 4'b1000;
										assign node9672 = (inp[5]) ? node9750 : node9673;
											assign node9673 = (inp[10]) ? node9705 : node9674;
												assign node9674 = (inp[4]) ? node9692 : node9675;
													assign node9675 = (inp[9]) ? node9687 : node9676;
														assign node9676 = (inp[3]) ? node9682 : node9677;
															assign node9677 = (inp[15]) ? 4'b1110 : node9678;
																assign node9678 = (inp[0]) ? 4'b1100 : 4'b1110;
															assign node9682 = (inp[0]) ? node9684 : 4'b1100;
																assign node9684 = (inp[15]) ? 4'b1110 : 4'b1100;
														assign node9687 = (inp[15]) ? node9689 : 4'b1010;
															assign node9689 = (inp[0]) ? 4'b1010 : 4'b1000;
													assign node9692 = (inp[9]) ? node9698 : node9693;
														assign node9693 = (inp[15]) ? node9695 : 4'b1000;
															assign node9695 = (inp[0]) ? 4'b1010 : 4'b1000;
														assign node9698 = (inp[3]) ? node9700 : 4'b1100;
															assign node9700 = (inp[0]) ? 4'b1110 : node9701;
																assign node9701 = (inp[15]) ? 4'b1110 : 4'b1100;
												assign node9705 = (inp[3]) ? node9723 : node9706;
													assign node9706 = (inp[9]) ? node9720 : node9707;
														assign node9707 = (inp[4]) ? node9715 : node9708;
															assign node9708 = (inp[0]) ? node9712 : node9709;
																assign node9709 = (inp[15]) ? 4'b1000 : 4'b1010;
																assign node9712 = (inp[15]) ? 4'b1010 : 4'b1000;
															assign node9715 = (inp[0]) ? node9717 : 4'b1110;
																assign node9717 = (inp[15]) ? 4'b1110 : 4'b1100;
														assign node9720 = (inp[4]) ? 4'b1010 : 4'b1110;
													assign node9723 = (inp[4]) ? node9735 : node9724;
														assign node9724 = (inp[9]) ? node9728 : node9725;
															assign node9725 = (inp[15]) ? 4'b1000 : 4'b1010;
															assign node9728 = (inp[15]) ? node9732 : node9729;
																assign node9729 = (inp[0]) ? 4'b1110 : 4'b1100;
																assign node9732 = (inp[0]) ? 4'b1100 : 4'b1110;
														assign node9735 = (inp[9]) ? node9743 : node9736;
															assign node9736 = (inp[0]) ? node9740 : node9737;
																assign node9737 = (inp[15]) ? 4'b1110 : 4'b1100;
																assign node9740 = (inp[15]) ? 4'b1100 : 4'b1110;
															assign node9743 = (inp[0]) ? node9747 : node9744;
																assign node9744 = (inp[15]) ? 4'b1010 : 4'b1000;
																assign node9747 = (inp[15]) ? 4'b1000 : 4'b1010;
											assign node9750 = (inp[0]) ? node9800 : node9751;
												assign node9751 = (inp[15]) ? node9773 : node9752;
													assign node9752 = (inp[3]) ? node9760 : node9753;
														assign node9753 = (inp[9]) ? 4'b1100 : node9754;
															assign node9754 = (inp[4]) ? 4'b1010 : node9755;
																assign node9755 = (inp[10]) ? 4'b1010 : 4'b1110;
														assign node9760 = (inp[4]) ? node9768 : node9761;
															assign node9761 = (inp[10]) ? node9765 : node9762;
																assign node9762 = (inp[9]) ? 4'b1000 : 4'b1100;
																assign node9765 = (inp[9]) ? 4'b1100 : 4'b1000;
															assign node9768 = (inp[9]) ? node9770 : 4'b1100;
																assign node9770 = (inp[10]) ? 4'b1000 : 4'b1100;
													assign node9773 = (inp[3]) ? node9787 : node9774;
														assign node9774 = (inp[9]) ? node9782 : node9775;
															assign node9775 = (inp[10]) ? node9779 : node9776;
																assign node9776 = (inp[4]) ? 4'b1000 : 4'b1100;
																assign node9779 = (inp[4]) ? 4'b1110 : 4'b1000;
															assign node9782 = (inp[10]) ? node9784 : 4'b1110;
																assign node9784 = (inp[4]) ? 4'b1010 : 4'b1110;
														assign node9787 = (inp[9]) ? node9793 : node9788;
															assign node9788 = (inp[4]) ? node9790 : 4'b1110;
																assign node9790 = (inp[10]) ? 4'b1110 : 4'b1010;
															assign node9793 = (inp[4]) ? node9797 : node9794;
																assign node9794 = (inp[10]) ? 4'b1110 : 4'b1010;
																assign node9797 = (inp[10]) ? 4'b1010 : 4'b1110;
												assign node9800 = (inp[15]) ? node9822 : node9801;
													assign node9801 = (inp[3]) ? node9809 : node9802;
														assign node9802 = (inp[4]) ? node9804 : 4'b1110;
															assign node9804 = (inp[9]) ? node9806 : 4'b1110;
																assign node9806 = (inp[10]) ? 4'b1010 : 4'b1110;
														assign node9809 = (inp[10]) ? node9815 : node9810;
															assign node9810 = (inp[9]) ? 4'b1010 : node9811;
																assign node9811 = (inp[4]) ? 4'b1010 : 4'b1110;
															assign node9815 = (inp[9]) ? node9819 : node9816;
																assign node9816 = (inp[4]) ? 4'b1110 : 4'b1010;
																assign node9819 = (inp[4]) ? 4'b1010 : 4'b1110;
													assign node9822 = (inp[4]) ? 4'b1100 : node9823;
														assign node9823 = (inp[3]) ? 4'b1000 : 4'b1010;
									assign node9827 = (inp[3]) ? node9963 : node9828;
										assign node9828 = (inp[15]) ? node9904 : node9829;
											assign node9829 = (inp[0]) ? node9875 : node9830;
												assign node9830 = (inp[5]) ? node9854 : node9831;
													assign node9831 = (inp[9]) ? node9843 : node9832;
														assign node9832 = (inp[4]) ? node9838 : node9833;
															assign node9833 = (inp[10]) ? node9835 : 4'b0111;
																assign node9835 = (inp[12]) ? 4'b0011 : 4'b0111;
															assign node9838 = (inp[10]) ? node9840 : 4'b0011;
																assign node9840 = (inp[12]) ? 4'b0111 : 4'b0011;
														assign node9843 = (inp[4]) ? node9849 : node9844;
															assign node9844 = (inp[12]) ? node9846 : 4'b0011;
																assign node9846 = (inp[10]) ? 4'b0111 : 4'b0011;
															assign node9849 = (inp[10]) ? node9851 : 4'b0111;
																assign node9851 = (inp[12]) ? 4'b0011 : 4'b0111;
													assign node9854 = (inp[9]) ? node9866 : node9855;
														assign node9855 = (inp[4]) ? node9861 : node9856;
															assign node9856 = (inp[12]) ? node9858 : 4'b0111;
																assign node9858 = (inp[10]) ? 4'b0011 : 4'b0111;
															assign node9861 = (inp[10]) ? node9863 : 4'b0011;
																assign node9863 = (inp[12]) ? 4'b0101 : 4'b0011;
														assign node9866 = (inp[10]) ? node9868 : 4'b0011;
															assign node9868 = (inp[4]) ? node9872 : node9869;
																assign node9869 = (inp[12]) ? 4'b0101 : 4'b0011;
																assign node9872 = (inp[12]) ? 4'b0001 : 4'b0101;
												assign node9875 = (inp[5]) ? node9891 : node9876;
													assign node9876 = (inp[9]) ? node9884 : node9877;
														assign node9877 = (inp[4]) ? 4'b0001 : node9878;
															assign node9878 = (inp[12]) ? node9880 : 4'b0101;
																assign node9880 = (inp[10]) ? 4'b0001 : 4'b0101;
														assign node9884 = (inp[4]) ? node9888 : node9885;
															assign node9885 = (inp[10]) ? 4'b0101 : 4'b0001;
															assign node9888 = (inp[10]) ? 4'b0001 : 4'b0101;
													assign node9891 = (inp[12]) ? node9899 : node9892;
														assign node9892 = (inp[4]) ? node9896 : node9893;
															assign node9893 = (inp[9]) ? 4'b0001 : 4'b0101;
															assign node9896 = (inp[9]) ? 4'b0111 : 4'b0001;
														assign node9899 = (inp[10]) ? node9901 : 4'b0111;
															assign node9901 = (inp[4]) ? 4'b0011 : 4'b0111;
											assign node9904 = (inp[0]) ? node9936 : node9905;
												assign node9905 = (inp[5]) ? node9921 : node9906;
													assign node9906 = (inp[4]) ? node9916 : node9907;
														assign node9907 = (inp[9]) ? node9911 : node9908;
															assign node9908 = (inp[10]) ? 4'b0001 : 4'b0101;
															assign node9911 = (inp[12]) ? node9913 : 4'b0001;
																assign node9913 = (inp[10]) ? 4'b0101 : 4'b0001;
														assign node9916 = (inp[9]) ? 4'b0101 : node9917;
															assign node9917 = (inp[10]) ? 4'b0101 : 4'b0001;
													assign node9921 = (inp[9]) ? node9929 : node9922;
														assign node9922 = (inp[12]) ? node9924 : 4'b0001;
															assign node9924 = (inp[4]) ? 4'b0111 : node9925;
																assign node9925 = (inp[10]) ? 4'b0001 : 4'b0101;
														assign node9929 = (inp[12]) ? node9931 : 4'b0111;
															assign node9931 = (inp[4]) ? node9933 : 4'b0111;
																assign node9933 = (inp[10]) ? 4'b0011 : 4'b0111;
												assign node9936 = (inp[5]) ? node9946 : node9937;
													assign node9937 = (inp[10]) ? 4'b0111 : node9938;
														assign node9938 = (inp[9]) ? node9942 : node9939;
															assign node9939 = (inp[4]) ? 4'b0011 : 4'b0111;
															assign node9942 = (inp[4]) ? 4'b0111 : 4'b0011;
													assign node9946 = (inp[4]) ? node9956 : node9947;
														assign node9947 = (inp[9]) ? node9953 : node9948;
															assign node9948 = (inp[12]) ? node9950 : 4'b0111;
																assign node9950 = (inp[10]) ? 4'b0011 : 4'b0111;
															assign node9953 = (inp[12]) ? 4'b0101 : 4'b0011;
														assign node9956 = (inp[12]) ? node9958 : 4'b0101;
															assign node9958 = (inp[10]) ? node9960 : 4'b0011;
																assign node9960 = (inp[9]) ? 4'b0001 : 4'b0101;
										assign node9963 = (inp[0]) ? node10055 : node9964;
											assign node9964 = (inp[15]) ? node10012 : node9965;
												assign node9965 = (inp[5]) ? node9985 : node9966;
													assign node9966 = (inp[12]) ? node9972 : node9967;
														assign node9967 = (inp[4]) ? 4'b0011 : node9968;
															assign node9968 = (inp[9]) ? 4'b0011 : 4'b0111;
														assign node9972 = (inp[4]) ? node9980 : node9973;
															assign node9973 = (inp[9]) ? node9977 : node9974;
																assign node9974 = (inp[10]) ? 4'b0011 : 4'b0111;
																assign node9977 = (inp[10]) ? 4'b0101 : 4'b0011;
															assign node9980 = (inp[10]) ? node9982 : 4'b0101;
																assign node9982 = (inp[9]) ? 4'b0001 : 4'b0101;
													assign node9985 = (inp[10]) ? node9999 : node9986;
														assign node9986 = (inp[12]) ? node9992 : node9987;
															assign node9987 = (inp[9]) ? 4'b0101 : node9988;
																assign node9988 = (inp[4]) ? 4'b0001 : 4'b0101;
															assign node9992 = (inp[4]) ? node9996 : node9993;
																assign node9993 = (inp[9]) ? 4'b0001 : 4'b0101;
																assign node9996 = (inp[9]) ? 4'b0101 : 4'b0001;
														assign node9999 = (inp[4]) ? node10007 : node10000;
															assign node10000 = (inp[12]) ? node10004 : node10001;
																assign node10001 = (inp[9]) ? 4'b0001 : 4'b0101;
																assign node10004 = (inp[9]) ? 4'b0101 : 4'b0001;
															assign node10007 = (inp[9]) ? 4'b0001 : node10008;
																assign node10008 = (inp[12]) ? 4'b0101 : 4'b0001;
												assign node10012 = (inp[5]) ? node10030 : node10013;
													assign node10013 = (inp[10]) ? node10019 : node10014;
														assign node10014 = (inp[12]) ? 4'b0001 : node10015;
															assign node10015 = (inp[9]) ? 4'b0001 : 4'b0101;
														assign node10019 = (inp[9]) ? node10027 : node10020;
															assign node10020 = (inp[12]) ? node10024 : node10021;
																assign node10021 = (inp[4]) ? 4'b0001 : 4'b0101;
																assign node10024 = (inp[4]) ? 4'b0111 : 4'b0001;
															assign node10027 = (inp[4]) ? 4'b0011 : 4'b0111;
													assign node10030 = (inp[10]) ? node10040 : node10031;
														assign node10031 = (inp[12]) ? 4'b0111 : node10032;
															assign node10032 = (inp[4]) ? node10036 : node10033;
																assign node10033 = (inp[9]) ? 4'b0011 : 4'b0111;
																assign node10036 = (inp[9]) ? 4'b0111 : 4'b0011;
														assign node10040 = (inp[12]) ? node10048 : node10041;
															assign node10041 = (inp[9]) ? node10045 : node10042;
																assign node10042 = (inp[4]) ? 4'b0011 : 4'b0111;
																assign node10045 = (inp[4]) ? 4'b0111 : 4'b0011;
															assign node10048 = (inp[9]) ? node10052 : node10049;
																assign node10049 = (inp[4]) ? 4'b0111 : 4'b0011;
																assign node10052 = (inp[4]) ? 4'b0011 : 4'b0111;
											assign node10055 = (inp[15]) ? node10087 : node10056;
												assign node10056 = (inp[5]) ? node10074 : node10057;
													assign node10057 = (inp[4]) ? node10069 : node10058;
														assign node10058 = (inp[9]) ? node10064 : node10059;
															assign node10059 = (inp[10]) ? node10061 : 4'b0101;
																assign node10061 = (inp[12]) ? 4'b0001 : 4'b0101;
															assign node10064 = (inp[10]) ? node10066 : 4'b0001;
																assign node10066 = (inp[12]) ? 4'b0111 : 4'b0001;
														assign node10069 = (inp[9]) ? 4'b0111 : node10070;
															assign node10070 = (inp[10]) ? 4'b0111 : 4'b0001;
													assign node10074 = (inp[4]) ? node10082 : node10075;
														assign node10075 = (inp[9]) ? node10077 : 4'b0111;
															assign node10077 = (inp[10]) ? node10079 : 4'b0011;
																assign node10079 = (inp[12]) ? 4'b0111 : 4'b0011;
														assign node10082 = (inp[10]) ? 4'b0111 : node10083;
															assign node10083 = (inp[9]) ? 4'b0111 : 4'b0011;
												assign node10087 = (inp[5]) ? node10101 : node10088;
													assign node10088 = (inp[4]) ? node10094 : node10089;
														assign node10089 = (inp[9]) ? 4'b0011 : node10090;
															assign node10090 = (inp[10]) ? 4'b0011 : 4'b0111;
														assign node10094 = (inp[9]) ? 4'b0101 : node10095;
															assign node10095 = (inp[10]) ? node10097 : 4'b0011;
																assign node10097 = (inp[12]) ? 4'b0101 : 4'b0011;
													assign node10101 = (inp[10]) ? node10109 : node10102;
														assign node10102 = (inp[9]) ? node10106 : node10103;
															assign node10103 = (inp[4]) ? 4'b0001 : 4'b0101;
															assign node10106 = (inp[4]) ? 4'b0101 : 4'b0001;
														assign node10109 = (inp[12]) ? node10117 : node10110;
															assign node10110 = (inp[9]) ? node10114 : node10111;
																assign node10111 = (inp[4]) ? 4'b0001 : 4'b0101;
																assign node10114 = (inp[4]) ? 4'b0101 : 4'b0001;
															assign node10117 = (inp[4]) ? node10121 : node10118;
																assign node10118 = (inp[9]) ? 4'b0101 : 4'b0001;
																assign node10121 = (inp[9]) ? 4'b0001 : 4'b0101;
								assign node10124 = (inp[4]) ? node10332 : node10125;
									assign node10125 = (inp[9]) ? node10263 : node10126;
										assign node10126 = (inp[12]) ? node10194 : node10127;
											assign node10127 = (inp[2]) ? node10171 : node10128;
												assign node10128 = (inp[10]) ? node10150 : node10129;
													assign node10129 = (inp[5]) ? node10137 : node10130;
														assign node10130 = (inp[15]) ? node10134 : node10131;
															assign node10131 = (inp[0]) ? 4'b0101 : 4'b0111;
															assign node10134 = (inp[0]) ? 4'b0111 : 4'b0101;
														assign node10137 = (inp[15]) ? node10145 : node10138;
															assign node10138 = (inp[3]) ? node10142 : node10139;
																assign node10139 = (inp[0]) ? 4'b0101 : 4'b0111;
																assign node10142 = (inp[0]) ? 4'b0111 : 4'b0101;
															assign node10145 = (inp[0]) ? node10147 : 4'b0111;
																assign node10147 = (inp[3]) ? 4'b0101 : 4'b0111;
													assign node10150 = (inp[15]) ? node10162 : node10151;
														assign node10151 = (inp[0]) ? node10157 : node10152;
															assign node10152 = (inp[3]) ? node10154 : 4'b0111;
																assign node10154 = (inp[5]) ? 4'b0101 : 4'b0111;
															assign node10157 = (inp[3]) ? node10159 : 4'b0101;
																assign node10159 = (inp[5]) ? 4'b0111 : 4'b0101;
														assign node10162 = (inp[0]) ? node10168 : node10163;
															assign node10163 = (inp[5]) ? node10165 : 4'b0101;
																assign node10165 = (inp[3]) ? 4'b0111 : 4'b0101;
															assign node10168 = (inp[3]) ? 4'b0101 : 4'b0111;
												assign node10171 = (inp[15]) ? node10183 : node10172;
													assign node10172 = (inp[0]) ? node10178 : node10173;
														assign node10173 = (inp[3]) ? node10175 : 4'b0111;
															assign node10175 = (inp[5]) ? 4'b0101 : 4'b0111;
														assign node10178 = (inp[3]) ? node10180 : 4'b0101;
															assign node10180 = (inp[5]) ? 4'b0111 : 4'b0101;
													assign node10183 = (inp[0]) ? node10189 : node10184;
														assign node10184 = (inp[3]) ? node10186 : 4'b0101;
															assign node10186 = (inp[5]) ? 4'b0111 : 4'b0101;
														assign node10189 = (inp[5]) ? node10191 : 4'b0111;
															assign node10191 = (inp[3]) ? 4'b0101 : 4'b0111;
											assign node10194 = (inp[10]) ? node10234 : node10195;
												assign node10195 = (inp[3]) ? node10211 : node10196;
													assign node10196 = (inp[5]) ? node10198 : 4'b0101;
														assign node10198 = (inp[2]) ? node10204 : node10199;
															assign node10199 = (inp[15]) ? node10201 : 4'b0101;
																assign node10201 = (inp[0]) ? 4'b0111 : 4'b0101;
															assign node10204 = (inp[15]) ? node10208 : node10205;
																assign node10205 = (inp[0]) ? 4'b0101 : 4'b0111;
																assign node10208 = (inp[0]) ? 4'b0111 : 4'b0101;
													assign node10211 = (inp[0]) ? node10219 : node10212;
														assign node10212 = (inp[5]) ? node10216 : node10213;
															assign node10213 = (inp[15]) ? 4'b0101 : 4'b0111;
															assign node10216 = (inp[15]) ? 4'b0111 : 4'b0101;
														assign node10219 = (inp[2]) ? node10227 : node10220;
															assign node10220 = (inp[15]) ? node10224 : node10221;
																assign node10221 = (inp[5]) ? 4'b0111 : 4'b0101;
																assign node10224 = (inp[5]) ? 4'b0101 : 4'b0111;
															assign node10227 = (inp[15]) ? node10231 : node10228;
																assign node10228 = (inp[5]) ? 4'b0111 : 4'b0101;
																assign node10231 = (inp[5]) ? 4'b0101 : 4'b0111;
												assign node10234 = (inp[3]) ? node10242 : node10235;
													assign node10235 = (inp[0]) ? node10239 : node10236;
														assign node10236 = (inp[15]) ? 4'b0001 : 4'b0011;
														assign node10239 = (inp[15]) ? 4'b0011 : 4'b0001;
													assign node10242 = (inp[15]) ? node10248 : node10243;
														assign node10243 = (inp[0]) ? node10245 : 4'b0011;
															assign node10245 = (inp[5]) ? 4'b0011 : 4'b0001;
														assign node10248 = (inp[2]) ? node10256 : node10249;
															assign node10249 = (inp[0]) ? node10253 : node10250;
																assign node10250 = (inp[5]) ? 4'b0011 : 4'b0001;
																assign node10253 = (inp[5]) ? 4'b0001 : 4'b0011;
															assign node10256 = (inp[0]) ? node10260 : node10257;
																assign node10257 = (inp[5]) ? 4'b0011 : 4'b0001;
																assign node10260 = (inp[5]) ? 4'b0001 : 4'b0011;
										assign node10263 = (inp[10]) ? node10287 : node10264;
											assign node10264 = (inp[0]) ? node10276 : node10265;
												assign node10265 = (inp[15]) ? node10271 : node10266;
													assign node10266 = (inp[3]) ? node10268 : 4'b0011;
														assign node10268 = (inp[5]) ? 4'b0001 : 4'b0011;
													assign node10271 = (inp[3]) ? node10273 : 4'b0001;
														assign node10273 = (inp[5]) ? 4'b0011 : 4'b0001;
												assign node10276 = (inp[15]) ? node10282 : node10277;
													assign node10277 = (inp[5]) ? node10279 : 4'b0001;
														assign node10279 = (inp[3]) ? 4'b0011 : 4'b0001;
													assign node10282 = (inp[3]) ? node10284 : 4'b0011;
														assign node10284 = (inp[5]) ? 4'b0001 : 4'b0011;
											assign node10287 = (inp[12]) ? node10309 : node10288;
												assign node10288 = (inp[15]) ? node10300 : node10289;
													assign node10289 = (inp[0]) ? node10295 : node10290;
														assign node10290 = (inp[5]) ? node10292 : 4'b0011;
															assign node10292 = (inp[3]) ? 4'b0001 : 4'b0011;
														assign node10295 = (inp[3]) ? node10297 : 4'b0001;
															assign node10297 = (inp[5]) ? 4'b0011 : 4'b0001;
													assign node10300 = (inp[0]) ? node10306 : node10301;
														assign node10301 = (inp[5]) ? node10303 : 4'b0001;
															assign node10303 = (inp[3]) ? 4'b0011 : 4'b0001;
														assign node10306 = (inp[5]) ? 4'b0001 : 4'b0011;
												assign node10309 = (inp[15]) ? node10321 : node10310;
													assign node10310 = (inp[0]) ? node10316 : node10311;
														assign node10311 = (inp[3]) ? 4'b0101 : node10312;
															assign node10312 = (inp[5]) ? 4'b0101 : 4'b0111;
														assign node10316 = (inp[3]) ? 4'b0111 : node10317;
															assign node10317 = (inp[5]) ? 4'b0111 : 4'b0101;
													assign node10321 = (inp[0]) ? node10327 : node10322;
														assign node10322 = (inp[5]) ? 4'b0111 : node10323;
															assign node10323 = (inp[3]) ? 4'b0111 : 4'b0101;
														assign node10327 = (inp[2]) ? node10329 : 4'b0101;
															assign node10329 = (inp[3]) ? 4'b0101 : 4'b0111;
									assign node10332 = (inp[9]) ? node10424 : node10333;
										assign node10333 = (inp[10]) ? node10369 : node10334;
											assign node10334 = (inp[3]) ? node10350 : node10335;
												assign node10335 = (inp[12]) ? node10343 : node10336;
													assign node10336 = (inp[0]) ? node10340 : node10337;
														assign node10337 = (inp[15]) ? 4'b0001 : 4'b0011;
														assign node10340 = (inp[15]) ? 4'b0011 : 4'b0001;
													assign node10343 = (inp[15]) ? node10347 : node10344;
														assign node10344 = (inp[0]) ? 4'b0001 : 4'b0011;
														assign node10347 = (inp[0]) ? 4'b0011 : 4'b0001;
												assign node10350 = (inp[15]) ? node10362 : node10351;
													assign node10351 = (inp[2]) ? node10357 : node10352;
														assign node10352 = (inp[5]) ? 4'b0011 : node10353;
															assign node10353 = (inp[0]) ? 4'b0001 : 4'b0011;
														assign node10357 = (inp[0]) ? 4'b0011 : node10358;
															assign node10358 = (inp[5]) ? 4'b0001 : 4'b0011;
													assign node10362 = (inp[0]) ? node10366 : node10363;
														assign node10363 = (inp[5]) ? 4'b0011 : 4'b0001;
														assign node10366 = (inp[5]) ? 4'b0001 : 4'b0011;
											assign node10369 = (inp[12]) ? node10403 : node10370;
												assign node10370 = (inp[2]) ? node10386 : node10371;
													assign node10371 = (inp[15]) ? node10379 : node10372;
														assign node10372 = (inp[0]) ? 4'b0001 : node10373;
															assign node10373 = (inp[5]) ? node10375 : 4'b0011;
																assign node10375 = (inp[3]) ? 4'b0001 : 4'b0011;
														assign node10379 = (inp[0]) ? node10381 : 4'b0001;
															assign node10381 = (inp[5]) ? node10383 : 4'b0011;
																assign node10383 = (inp[3]) ? 4'b0001 : 4'b0011;
													assign node10386 = (inp[15]) ? node10398 : node10387;
														assign node10387 = (inp[0]) ? node10393 : node10388;
															assign node10388 = (inp[5]) ? node10390 : 4'b0011;
																assign node10390 = (inp[3]) ? 4'b0001 : 4'b0011;
															assign node10393 = (inp[3]) ? node10395 : 4'b0001;
																assign node10395 = (inp[5]) ? 4'b0011 : 4'b0001;
														assign node10398 = (inp[0]) ? 4'b0011 : node10399;
															assign node10399 = (inp[3]) ? 4'b0011 : 4'b0001;
												assign node10403 = (inp[0]) ? node10415 : node10404;
													assign node10404 = (inp[15]) ? node10410 : node10405;
														assign node10405 = (inp[5]) ? 4'b0101 : node10406;
															assign node10406 = (inp[3]) ? 4'b0101 : 4'b0111;
														assign node10410 = (inp[3]) ? 4'b0111 : node10411;
															assign node10411 = (inp[2]) ? 4'b0111 : 4'b0101;
													assign node10415 = (inp[15]) ? node10419 : node10416;
														assign node10416 = (inp[5]) ? 4'b0111 : 4'b0101;
														assign node10419 = (inp[5]) ? 4'b0101 : node10420;
															assign node10420 = (inp[3]) ? 4'b0101 : 4'b0111;
										assign node10424 = (inp[10]) ? node10474 : node10425;
											assign node10425 = (inp[12]) ? node10455 : node10426;
												assign node10426 = (inp[5]) ? node10438 : node10427;
													assign node10427 = (inp[3]) ? node10433 : node10428;
														assign node10428 = (inp[15]) ? 4'b0101 : node10429;
															assign node10429 = (inp[0]) ? 4'b0101 : 4'b0111;
														assign node10433 = (inp[15]) ? 4'b0111 : node10434;
															assign node10434 = (inp[0]) ? 4'b0111 : 4'b0101;
													assign node10438 = (inp[3]) ? node10444 : node10439;
														assign node10439 = (inp[15]) ? 4'b0111 : node10440;
															assign node10440 = (inp[0]) ? 4'b0111 : 4'b0101;
														assign node10444 = (inp[2]) ? node10450 : node10445;
															assign node10445 = (inp[0]) ? 4'b0101 : node10446;
																assign node10446 = (inp[15]) ? 4'b0111 : 4'b0101;
															assign node10450 = (inp[0]) ? node10452 : 4'b0101;
																assign node10452 = (inp[15]) ? 4'b0101 : 4'b0111;
												assign node10455 = (inp[15]) ? node10465 : node10456;
													assign node10456 = (inp[0]) ? node10460 : node10457;
														assign node10457 = (inp[5]) ? 4'b0101 : 4'b0111;
														assign node10460 = (inp[5]) ? 4'b0111 : node10461;
															assign node10461 = (inp[3]) ? 4'b0111 : 4'b0101;
													assign node10465 = (inp[0]) ? node10471 : node10466;
														assign node10466 = (inp[3]) ? 4'b0111 : node10467;
															assign node10467 = (inp[5]) ? 4'b0111 : 4'b0101;
														assign node10471 = (inp[3]) ? 4'b0101 : 4'b0111;
											assign node10474 = (inp[12]) ? node10498 : node10475;
												assign node10475 = (inp[15]) ? node10487 : node10476;
													assign node10476 = (inp[0]) ? node10482 : node10477;
														assign node10477 = (inp[3]) ? 4'b0101 : node10478;
															assign node10478 = (inp[5]) ? 4'b0101 : 4'b0111;
														assign node10482 = (inp[3]) ? 4'b0111 : node10483;
															assign node10483 = (inp[2]) ? 4'b0101 : 4'b0111;
													assign node10487 = (inp[0]) ? node10493 : node10488;
														assign node10488 = (inp[5]) ? 4'b0111 : node10489;
															assign node10489 = (inp[3]) ? 4'b0111 : 4'b0101;
														assign node10493 = (inp[5]) ? 4'b0101 : node10494;
															assign node10494 = (inp[3]) ? 4'b0101 : 4'b0111;
												assign node10498 = (inp[2]) ? node10516 : node10499;
													assign node10499 = (inp[5]) ? node10509 : node10500;
														assign node10500 = (inp[15]) ? 4'b0001 : node10501;
															assign node10501 = (inp[3]) ? node10505 : node10502;
																assign node10502 = (inp[0]) ? 4'b0001 : 4'b0011;
																assign node10505 = (inp[0]) ? 4'b0011 : 4'b0001;
														assign node10509 = (inp[15]) ? node10513 : node10510;
															assign node10510 = (inp[0]) ? 4'b0011 : 4'b0001;
															assign node10513 = (inp[0]) ? 4'b0001 : 4'b0011;
													assign node10516 = (inp[0]) ? node10518 : 4'b0011;
														assign node10518 = (inp[3]) ? node10524 : node10519;
															assign node10519 = (inp[15]) ? node10521 : 4'b0001;
																assign node10521 = (inp[5]) ? 4'b0001 : 4'b0011;
															assign node10524 = (inp[15]) ? 4'b0001 : 4'b0011;
						assign node10527 = (inp[8]) ? node11607 : node10528;
							assign node10528 = (inp[14]) ? node11096 : node10529;
								assign node10529 = (inp[2]) ? node10793 : node10530;
									assign node10530 = (inp[4]) ? node10652 : node10531;
										assign node10531 = (inp[9]) ? node10595 : node10532;
											assign node10532 = (inp[12]) ? node10560 : node10533;
												assign node10533 = (inp[10]) ? node10547 : node10534;
													assign node10534 = (inp[15]) ? node10542 : node10535;
														assign node10535 = (inp[0]) ? node10539 : node10536;
															assign node10536 = (inp[3]) ? 4'b1100 : 4'b1110;
															assign node10539 = (inp[3]) ? 4'b1110 : 4'b1100;
														assign node10542 = (inp[3]) ? 4'b1110 : node10543;
															assign node10543 = (inp[0]) ? 4'b1110 : 4'b1100;
													assign node10547 = (inp[5]) ? node10555 : node10548;
														assign node10548 = (inp[15]) ? node10552 : node10549;
															assign node10549 = (inp[0]) ? 4'b1100 : 4'b1110;
															assign node10552 = (inp[0]) ? 4'b1110 : 4'b1100;
														assign node10555 = (inp[3]) ? node10557 : 4'b1100;
															assign node10557 = (inp[15]) ? 4'b1100 : 4'b1110;
												assign node10560 = (inp[10]) ? node10574 : node10561;
													assign node10561 = (inp[5]) ? node10563 : 4'b1110;
														assign node10563 = (inp[0]) ? node10569 : node10564;
															assign node10564 = (inp[3]) ? 4'b1100 : node10565;
																assign node10565 = (inp[15]) ? 4'b1100 : 4'b1110;
															assign node10569 = (inp[3]) ? 4'b1110 : node10570;
																assign node10570 = (inp[15]) ? 4'b1110 : 4'b1100;
													assign node10574 = (inp[5]) ? node10582 : node10575;
														assign node10575 = (inp[15]) ? node10579 : node10576;
															assign node10576 = (inp[0]) ? 4'b1000 : 4'b1010;
															assign node10579 = (inp[0]) ? 4'b1010 : 4'b1000;
														assign node10582 = (inp[0]) ? node10590 : node10583;
															assign node10583 = (inp[15]) ? node10587 : node10584;
																assign node10584 = (inp[3]) ? 4'b1000 : 4'b1010;
																assign node10587 = (inp[3]) ? 4'b1010 : 4'b1000;
															assign node10590 = (inp[15]) ? 4'b1000 : node10591;
																assign node10591 = (inp[3]) ? 4'b1010 : 4'b1000;
											assign node10595 = (inp[12]) ? node10619 : node10596;
												assign node10596 = (inp[0]) ? node10608 : node10597;
													assign node10597 = (inp[15]) ? node10603 : node10598;
														assign node10598 = (inp[5]) ? node10600 : 4'b1010;
															assign node10600 = (inp[3]) ? 4'b1000 : 4'b1010;
														assign node10603 = (inp[5]) ? node10605 : 4'b1000;
															assign node10605 = (inp[3]) ? 4'b1010 : 4'b1000;
													assign node10608 = (inp[15]) ? node10614 : node10609;
														assign node10609 = (inp[5]) ? node10611 : 4'b1000;
															assign node10611 = (inp[3]) ? 4'b1010 : 4'b1000;
														assign node10614 = (inp[5]) ? node10616 : 4'b1010;
															assign node10616 = (inp[3]) ? 4'b1000 : 4'b1010;
												assign node10619 = (inp[10]) ? node10639 : node10620;
													assign node10620 = (inp[0]) ? node10630 : node10621;
														assign node10621 = (inp[5]) ? node10623 : 4'b1010;
															assign node10623 = (inp[15]) ? node10627 : node10624;
																assign node10624 = (inp[3]) ? 4'b1000 : 4'b1010;
																assign node10627 = (inp[3]) ? 4'b1010 : 4'b1000;
														assign node10630 = (inp[3]) ? node10632 : 4'b1000;
															assign node10632 = (inp[5]) ? node10636 : node10633;
																assign node10633 = (inp[15]) ? 4'b1010 : 4'b1000;
																assign node10636 = (inp[15]) ? 4'b1000 : 4'b1010;
													assign node10639 = (inp[15]) ? node10647 : node10640;
														assign node10640 = (inp[0]) ? 4'b1110 : node10641;
															assign node10641 = (inp[3]) ? 4'b1100 : node10642;
																assign node10642 = (inp[5]) ? 4'b1100 : 4'b1110;
														assign node10647 = (inp[0]) ? 4'b1100 : node10648;
															assign node10648 = (inp[5]) ? 4'b1110 : 4'b1100;
										assign node10652 = (inp[9]) ? node10732 : node10653;
											assign node10653 = (inp[12]) ? node10693 : node10654;
												assign node10654 = (inp[3]) ? node10676 : node10655;
													assign node10655 = (inp[5]) ? node10667 : node10656;
														assign node10656 = (inp[10]) ? node10662 : node10657;
															assign node10657 = (inp[15]) ? node10659 : 4'b1010;
																assign node10659 = (inp[0]) ? 4'b1010 : 4'b1000;
															assign node10662 = (inp[15]) ? 4'b1010 : node10663;
																assign node10663 = (inp[0]) ? 4'b1000 : 4'b1010;
														assign node10667 = (inp[10]) ? node10671 : node10668;
															assign node10668 = (inp[15]) ? 4'b1000 : 4'b1010;
															assign node10671 = (inp[15]) ? node10673 : 4'b1000;
																assign node10673 = (inp[0]) ? 4'b1010 : 4'b1000;
													assign node10676 = (inp[5]) ? node10684 : node10677;
														assign node10677 = (inp[0]) ? node10681 : node10678;
															assign node10678 = (inp[15]) ? 4'b1000 : 4'b1010;
															assign node10681 = (inp[15]) ? 4'b1010 : 4'b1000;
														assign node10684 = (inp[10]) ? node10688 : node10685;
															assign node10685 = (inp[15]) ? 4'b1010 : 4'b1000;
															assign node10688 = (inp[0]) ? node10690 : 4'b1010;
																assign node10690 = (inp[15]) ? 4'b1000 : 4'b1010;
												assign node10693 = (inp[10]) ? node10711 : node10694;
													assign node10694 = (inp[5]) ? node10702 : node10695;
														assign node10695 = (inp[15]) ? node10699 : node10696;
															assign node10696 = (inp[0]) ? 4'b1000 : 4'b1010;
															assign node10699 = (inp[0]) ? 4'b1010 : 4'b1000;
														assign node10702 = (inp[15]) ? node10704 : 4'b1000;
															assign node10704 = (inp[3]) ? node10708 : node10705;
																assign node10705 = (inp[0]) ? 4'b1010 : 4'b1000;
																assign node10708 = (inp[0]) ? 4'b1000 : 4'b1010;
													assign node10711 = (inp[5]) ? node10725 : node10712;
														assign node10712 = (inp[15]) ? node10718 : node10713;
															assign node10713 = (inp[0]) ? node10715 : 4'b1110;
																assign node10715 = (inp[3]) ? 4'b1110 : 4'b1100;
															assign node10718 = (inp[0]) ? node10722 : node10719;
																assign node10719 = (inp[3]) ? 4'b1110 : 4'b1100;
																assign node10722 = (inp[3]) ? 4'b1100 : 4'b1110;
														assign node10725 = (inp[0]) ? node10729 : node10726;
															assign node10726 = (inp[15]) ? 4'b1110 : 4'b1100;
															assign node10729 = (inp[15]) ? 4'b1100 : 4'b1110;
											assign node10732 = (inp[12]) ? node10754 : node10733;
												assign node10733 = (inp[0]) ? node10743 : node10734;
													assign node10734 = (inp[15]) ? node10738 : node10735;
														assign node10735 = (inp[5]) ? 4'b1100 : 4'b1110;
														assign node10738 = (inp[5]) ? 4'b1110 : node10739;
															assign node10739 = (inp[3]) ? 4'b1110 : 4'b1100;
													assign node10743 = (inp[15]) ? node10749 : node10744;
														assign node10744 = (inp[5]) ? 4'b1110 : node10745;
															assign node10745 = (inp[3]) ? 4'b1110 : 4'b1100;
														assign node10749 = (inp[3]) ? 4'b1100 : node10750;
															assign node10750 = (inp[5]) ? 4'b1100 : 4'b1110;
												assign node10754 = (inp[10]) ? node10774 : node10755;
													assign node10755 = (inp[0]) ? node10765 : node10756;
														assign node10756 = (inp[3]) ? node10762 : node10757;
															assign node10757 = (inp[15]) ? 4'b1100 : node10758;
																assign node10758 = (inp[5]) ? 4'b1100 : 4'b1110;
															assign node10762 = (inp[15]) ? 4'b1110 : 4'b1100;
														assign node10765 = (inp[3]) ? node10771 : node10766;
															assign node10766 = (inp[15]) ? 4'b1110 : node10767;
																assign node10767 = (inp[5]) ? 4'b1110 : 4'b1100;
															assign node10771 = (inp[15]) ? 4'b1100 : 4'b1110;
													assign node10774 = (inp[0]) ? node10786 : node10775;
														assign node10775 = (inp[15]) ? node10781 : node10776;
															assign node10776 = (inp[5]) ? 4'b1000 : node10777;
																assign node10777 = (inp[3]) ? 4'b1000 : 4'b1010;
															assign node10781 = (inp[5]) ? 4'b1010 : node10782;
																assign node10782 = (inp[3]) ? 4'b1010 : 4'b1000;
														assign node10786 = (inp[15]) ? node10788 : 4'b1010;
															assign node10788 = (inp[3]) ? 4'b1000 : node10789;
																assign node10789 = (inp[5]) ? 4'b1000 : 4'b1010;
									assign node10793 = (inp[12]) ? node10933 : node10794;
										assign node10794 = (inp[5]) ? node10860 : node10795;
											assign node10795 = (inp[4]) ? node10819 : node10796;
												assign node10796 = (inp[9]) ? node10812 : node10797;
													assign node10797 = (inp[3]) ? node10803 : node10798;
														assign node10798 = (inp[0]) ? 4'b0101 : node10799;
															assign node10799 = (inp[15]) ? 4'b0101 : 4'b0111;
														assign node10803 = (inp[10]) ? 4'b0111 : node10804;
															assign node10804 = (inp[0]) ? node10808 : node10805;
																assign node10805 = (inp[15]) ? 4'b0101 : 4'b0111;
																assign node10808 = (inp[15]) ? 4'b0111 : 4'b0101;
													assign node10812 = (inp[15]) ? node10816 : node10813;
														assign node10813 = (inp[0]) ? 4'b0001 : 4'b0011;
														assign node10816 = (inp[0]) ? 4'b0011 : 4'b0001;
												assign node10819 = (inp[9]) ? node10833 : node10820;
													assign node10820 = (inp[3]) ? node10828 : node10821;
														assign node10821 = (inp[0]) ? node10825 : node10822;
															assign node10822 = (inp[15]) ? 4'b0001 : 4'b0011;
															assign node10825 = (inp[15]) ? 4'b0011 : 4'b0001;
														assign node10828 = (inp[0]) ? node10830 : 4'b0001;
															assign node10830 = (inp[15]) ? 4'b0011 : 4'b0001;
													assign node10833 = (inp[10]) ? node10847 : node10834;
														assign node10834 = (inp[3]) ? node10842 : node10835;
															assign node10835 = (inp[15]) ? node10839 : node10836;
																assign node10836 = (inp[0]) ? 4'b0101 : 4'b0111;
																assign node10839 = (inp[0]) ? 4'b0111 : 4'b0101;
															assign node10842 = (inp[15]) ? 4'b0111 : node10843;
																assign node10843 = (inp[0]) ? 4'b0111 : 4'b0101;
														assign node10847 = (inp[3]) ? node10855 : node10848;
															assign node10848 = (inp[15]) ? node10852 : node10849;
																assign node10849 = (inp[0]) ? 4'b0101 : 4'b0111;
																assign node10852 = (inp[0]) ? 4'b0111 : 4'b0101;
															assign node10855 = (inp[0]) ? 4'b0101 : node10856;
																assign node10856 = (inp[15]) ? 4'b0111 : 4'b0101;
											assign node10860 = (inp[15]) ? node10896 : node10861;
												assign node10861 = (inp[0]) ? node10877 : node10862;
													assign node10862 = (inp[3]) ? node10870 : node10863;
														assign node10863 = (inp[4]) ? node10867 : node10864;
															assign node10864 = (inp[9]) ? 4'b0011 : 4'b0111;
															assign node10867 = (inp[9]) ? 4'b0101 : 4'b0011;
														assign node10870 = (inp[4]) ? node10874 : node10871;
															assign node10871 = (inp[9]) ? 4'b0001 : 4'b0101;
															assign node10874 = (inp[9]) ? 4'b0101 : 4'b0001;
													assign node10877 = (inp[3]) ? node10885 : node10878;
														assign node10878 = (inp[4]) ? node10882 : node10879;
															assign node10879 = (inp[9]) ? 4'b0001 : 4'b0101;
															assign node10882 = (inp[10]) ? 4'b0111 : 4'b0001;
														assign node10885 = (inp[10]) ? node10891 : node10886;
															assign node10886 = (inp[9]) ? 4'b0011 : node10887;
																assign node10887 = (inp[4]) ? 4'b0011 : 4'b0111;
															assign node10891 = (inp[4]) ? 4'b0111 : node10892;
																assign node10892 = (inp[9]) ? 4'b0011 : 4'b0111;
												assign node10896 = (inp[0]) ? node10920 : node10897;
													assign node10897 = (inp[3]) ? node10905 : node10898;
														assign node10898 = (inp[4]) ? node10902 : node10899;
															assign node10899 = (inp[9]) ? 4'b0001 : 4'b0101;
															assign node10902 = (inp[9]) ? 4'b0111 : 4'b0001;
														assign node10905 = (inp[10]) ? node10913 : node10906;
															assign node10906 = (inp[4]) ? node10910 : node10907;
																assign node10907 = (inp[9]) ? 4'b0011 : 4'b0111;
																assign node10910 = (inp[9]) ? 4'b0111 : 4'b0011;
															assign node10913 = (inp[4]) ? node10917 : node10914;
																assign node10914 = (inp[9]) ? 4'b0011 : 4'b0111;
																assign node10917 = (inp[9]) ? 4'b0111 : 4'b0011;
													assign node10920 = (inp[3]) ? node10928 : node10921;
														assign node10921 = (inp[9]) ? node10925 : node10922;
															assign node10922 = (inp[4]) ? 4'b0011 : 4'b0111;
															assign node10925 = (inp[4]) ? 4'b0101 : 4'b0011;
														assign node10928 = (inp[4]) ? node10930 : 4'b0101;
															assign node10930 = (inp[9]) ? 4'b0101 : 4'b0001;
										assign node10933 = (inp[5]) ? node11013 : node10934;
											assign node10934 = (inp[10]) ? node10968 : node10935;
												assign node10935 = (inp[9]) ? node10955 : node10936;
													assign node10936 = (inp[4]) ? node10942 : node10937;
														assign node10937 = (inp[0]) ? node10939 : 4'b0111;
															assign node10939 = (inp[15]) ? 4'b0111 : 4'b0101;
														assign node10942 = (inp[3]) ? node10950 : node10943;
															assign node10943 = (inp[0]) ? node10947 : node10944;
																assign node10944 = (inp[15]) ? 4'b0001 : 4'b0011;
																assign node10947 = (inp[15]) ? 4'b0011 : 4'b0001;
															assign node10950 = (inp[15]) ? 4'b0001 : node10951;
																assign node10951 = (inp[0]) ? 4'b0001 : 4'b0011;
													assign node10955 = (inp[4]) ? node10961 : node10956;
														assign node10956 = (inp[15]) ? 4'b0001 : node10957;
															assign node10957 = (inp[0]) ? 4'b0001 : 4'b0011;
														assign node10961 = (inp[0]) ? 4'b0111 : node10962;
															assign node10962 = (inp[15]) ? node10964 : 4'b0101;
																assign node10964 = (inp[3]) ? 4'b0111 : 4'b0101;
												assign node10968 = (inp[4]) ? node10990 : node10969;
													assign node10969 = (inp[9]) ? node10981 : node10970;
														assign node10970 = (inp[3]) ? node10976 : node10971;
															assign node10971 = (inp[0]) ? 4'b0001 : node10972;
																assign node10972 = (inp[15]) ? 4'b0001 : 4'b0011;
															assign node10976 = (inp[0]) ? 4'b0011 : node10977;
																assign node10977 = (inp[15]) ? 4'b0001 : 4'b0011;
														assign node10981 = (inp[15]) ? 4'b0111 : node10982;
															assign node10982 = (inp[3]) ? node10986 : node10983;
																assign node10983 = (inp[0]) ? 4'b0101 : 4'b0111;
																assign node10986 = (inp[0]) ? 4'b0111 : 4'b0101;
													assign node10990 = (inp[9]) ? node11006 : node10991;
														assign node10991 = (inp[3]) ? node10999 : node10992;
															assign node10992 = (inp[15]) ? node10996 : node10993;
																assign node10993 = (inp[0]) ? 4'b0101 : 4'b0111;
																assign node10996 = (inp[0]) ? 4'b0111 : 4'b0101;
															assign node10999 = (inp[0]) ? node11003 : node11000;
																assign node11000 = (inp[15]) ? 4'b0111 : 4'b0101;
																assign node11003 = (inp[15]) ? 4'b0101 : 4'b0111;
														assign node11006 = (inp[15]) ? node11008 : 4'b0001;
															assign node11008 = (inp[3]) ? node11010 : 4'b0011;
																assign node11010 = (inp[0]) ? 4'b0001 : 4'b0011;
											assign node11013 = (inp[9]) ? node11067 : node11014;
												assign node11014 = (inp[4]) ? node11040 : node11015;
													assign node11015 = (inp[10]) ? node11025 : node11016;
														assign node11016 = (inp[15]) ? 4'b0101 : node11017;
															assign node11017 = (inp[3]) ? node11021 : node11018;
																assign node11018 = (inp[0]) ? 4'b0101 : 4'b0111;
																assign node11021 = (inp[0]) ? 4'b0111 : 4'b0101;
														assign node11025 = (inp[15]) ? node11033 : node11026;
															assign node11026 = (inp[3]) ? node11030 : node11027;
																assign node11027 = (inp[0]) ? 4'b0001 : 4'b0011;
																assign node11030 = (inp[0]) ? 4'b0011 : 4'b0001;
															assign node11033 = (inp[3]) ? node11037 : node11034;
																assign node11034 = (inp[0]) ? 4'b0011 : 4'b0001;
																assign node11037 = (inp[0]) ? 4'b0001 : 4'b0011;
													assign node11040 = (inp[10]) ? node11054 : node11041;
														assign node11041 = (inp[15]) ? node11049 : node11042;
															assign node11042 = (inp[3]) ? node11046 : node11043;
																assign node11043 = (inp[0]) ? 4'b0001 : 4'b0011;
																assign node11046 = (inp[0]) ? 4'b0011 : 4'b0001;
															assign node11049 = (inp[0]) ? 4'b0011 : node11050;
																assign node11050 = (inp[3]) ? 4'b0011 : 4'b0001;
														assign node11054 = (inp[3]) ? node11060 : node11055;
															assign node11055 = (inp[0]) ? node11057 : 4'b0111;
																assign node11057 = (inp[15]) ? 4'b0101 : 4'b0111;
															assign node11060 = (inp[0]) ? node11064 : node11061;
																assign node11061 = (inp[15]) ? 4'b0111 : 4'b0101;
																assign node11064 = (inp[15]) ? 4'b0101 : 4'b0111;
												assign node11067 = (inp[3]) ? node11083 : node11068;
													assign node11068 = (inp[10]) ? node11076 : node11069;
														assign node11069 = (inp[4]) ? node11071 : 4'b0011;
															assign node11071 = (inp[15]) ? 4'b0111 : node11072;
																assign node11072 = (inp[0]) ? 4'b0111 : 4'b0101;
														assign node11076 = (inp[4]) ? node11078 : 4'b0101;
															assign node11078 = (inp[0]) ? 4'b0011 : node11079;
																assign node11079 = (inp[15]) ? 4'b0011 : 4'b0001;
													assign node11083 = (inp[15]) ? node11087 : node11084;
														assign node11084 = (inp[0]) ? 4'b0011 : 4'b0001;
														assign node11087 = (inp[0]) ? node11091 : node11088;
															assign node11088 = (inp[4]) ? 4'b0011 : 4'b0111;
															assign node11091 = (inp[4]) ? 4'b0001 : node11092;
																assign node11092 = (inp[10]) ? 4'b0101 : 4'b0001;
								assign node11096 = (inp[12]) ? node11316 : node11097;
									assign node11097 = (inp[2]) ? node11203 : node11098;
										assign node11098 = (inp[0]) ? node11150 : node11099;
											assign node11099 = (inp[15]) ? node11125 : node11100;
												assign node11100 = (inp[5]) ? node11110 : node11101;
													assign node11101 = (inp[9]) ? node11105 : node11102;
														assign node11102 = (inp[4]) ? 4'b0011 : 4'b0111;
														assign node11105 = (inp[4]) ? node11107 : 4'b0011;
															assign node11107 = (inp[3]) ? 4'b0101 : 4'b0111;
													assign node11110 = (inp[3]) ? node11118 : node11111;
														assign node11111 = (inp[4]) ? node11115 : node11112;
															assign node11112 = (inp[9]) ? 4'b0011 : 4'b0111;
															assign node11115 = (inp[9]) ? 4'b0101 : 4'b0011;
														assign node11118 = (inp[4]) ? node11122 : node11119;
															assign node11119 = (inp[9]) ? 4'b0001 : 4'b0101;
															assign node11122 = (inp[9]) ? 4'b0101 : 4'b0001;
												assign node11125 = (inp[5]) ? node11135 : node11126;
													assign node11126 = (inp[4]) ? node11130 : node11127;
														assign node11127 = (inp[9]) ? 4'b0001 : 4'b0101;
														assign node11130 = (inp[9]) ? node11132 : 4'b0001;
															assign node11132 = (inp[3]) ? 4'b0111 : 4'b0101;
													assign node11135 = (inp[3]) ? node11143 : node11136;
														assign node11136 = (inp[4]) ? node11140 : node11137;
															assign node11137 = (inp[9]) ? 4'b0001 : 4'b0101;
															assign node11140 = (inp[9]) ? 4'b0111 : 4'b0001;
														assign node11143 = (inp[4]) ? node11147 : node11144;
															assign node11144 = (inp[9]) ? 4'b0011 : 4'b0111;
															assign node11147 = (inp[9]) ? 4'b0111 : 4'b0011;
											assign node11150 = (inp[15]) ? node11176 : node11151;
												assign node11151 = (inp[5]) ? node11161 : node11152;
													assign node11152 = (inp[9]) ? node11156 : node11153;
														assign node11153 = (inp[4]) ? 4'b0001 : 4'b0101;
														assign node11156 = (inp[4]) ? node11158 : 4'b0001;
															assign node11158 = (inp[3]) ? 4'b0111 : 4'b0101;
													assign node11161 = (inp[3]) ? node11169 : node11162;
														assign node11162 = (inp[9]) ? node11166 : node11163;
															assign node11163 = (inp[4]) ? 4'b0001 : 4'b0101;
															assign node11166 = (inp[4]) ? 4'b0111 : 4'b0001;
														assign node11169 = (inp[4]) ? node11173 : node11170;
															assign node11170 = (inp[9]) ? 4'b0011 : 4'b0111;
															assign node11173 = (inp[9]) ? 4'b0111 : 4'b0011;
												assign node11176 = (inp[5]) ? node11186 : node11177;
													assign node11177 = (inp[9]) ? node11181 : node11178;
														assign node11178 = (inp[4]) ? 4'b0011 : 4'b0111;
														assign node11181 = (inp[4]) ? node11183 : 4'b0011;
															assign node11183 = (inp[3]) ? 4'b0101 : 4'b0111;
													assign node11186 = (inp[3]) ? node11194 : node11187;
														assign node11187 = (inp[9]) ? node11191 : node11188;
															assign node11188 = (inp[4]) ? 4'b0011 : 4'b0111;
															assign node11191 = (inp[4]) ? 4'b0101 : 4'b0011;
														assign node11194 = (inp[10]) ? 4'b0101 : node11195;
															assign node11195 = (inp[4]) ? node11199 : node11196;
																assign node11196 = (inp[9]) ? 4'b0001 : 4'b0101;
																assign node11199 = (inp[9]) ? 4'b0101 : 4'b0001;
										assign node11203 = (inp[0]) ? node11267 : node11204;
											assign node11204 = (inp[15]) ? node11236 : node11205;
												assign node11205 = (inp[5]) ? node11215 : node11206;
													assign node11206 = (inp[4]) ? node11210 : node11207;
														assign node11207 = (inp[9]) ? 4'b0011 : 4'b0111;
														assign node11210 = (inp[3]) ? 4'b0101 : node11211;
															assign node11211 = (inp[10]) ? 4'b0111 : 4'b0011;
													assign node11215 = (inp[3]) ? node11223 : node11216;
														assign node11216 = (inp[9]) ? node11220 : node11217;
															assign node11217 = (inp[4]) ? 4'b0011 : 4'b0111;
															assign node11220 = (inp[4]) ? 4'b0101 : 4'b0011;
														assign node11223 = (inp[10]) ? node11229 : node11224;
															assign node11224 = (inp[9]) ? 4'b0001 : node11225;
																assign node11225 = (inp[4]) ? 4'b0001 : 4'b0101;
															assign node11229 = (inp[9]) ? node11233 : node11230;
																assign node11230 = (inp[4]) ? 4'b0001 : 4'b0101;
																assign node11233 = (inp[4]) ? 4'b0101 : 4'b0001;
												assign node11236 = (inp[5]) ? node11252 : node11237;
													assign node11237 = (inp[10]) ? node11247 : node11238;
														assign node11238 = (inp[4]) ? node11242 : node11239;
															assign node11239 = (inp[9]) ? 4'b0001 : 4'b0101;
															assign node11242 = (inp[9]) ? node11244 : 4'b0001;
																assign node11244 = (inp[3]) ? 4'b0111 : 4'b0101;
														assign node11247 = (inp[4]) ? node11249 : 4'b0001;
															assign node11249 = (inp[9]) ? 4'b0111 : 4'b0001;
													assign node11252 = (inp[3]) ? node11260 : node11253;
														assign node11253 = (inp[4]) ? node11257 : node11254;
															assign node11254 = (inp[9]) ? 4'b0001 : 4'b0101;
															assign node11257 = (inp[9]) ? 4'b0111 : 4'b0001;
														assign node11260 = (inp[10]) ? 4'b0111 : node11261;
															assign node11261 = (inp[4]) ? 4'b0011 : node11262;
																assign node11262 = (inp[9]) ? 4'b0011 : 4'b0111;
											assign node11267 = (inp[15]) ? node11297 : node11268;
												assign node11268 = (inp[5]) ? node11284 : node11269;
													assign node11269 = (inp[10]) ? node11277 : node11270;
														assign node11270 = (inp[9]) ? node11274 : node11271;
															assign node11271 = (inp[4]) ? 4'b0001 : 4'b0101;
															assign node11274 = (inp[4]) ? 4'b0101 : 4'b0001;
														assign node11277 = (inp[3]) ? node11281 : node11278;
															assign node11278 = (inp[4]) ? 4'b0101 : 4'b0001;
															assign node11281 = (inp[4]) ? 4'b0111 : 4'b0101;
													assign node11284 = (inp[3]) ? node11290 : node11285;
														assign node11285 = (inp[9]) ? 4'b0111 : node11286;
															assign node11286 = (inp[4]) ? 4'b0001 : 4'b0101;
														assign node11290 = (inp[9]) ? node11294 : node11291;
															assign node11291 = (inp[4]) ? 4'b0011 : 4'b0111;
															assign node11294 = (inp[4]) ? 4'b0111 : 4'b0011;
												assign node11297 = (inp[4]) ? node11305 : node11298;
													assign node11298 = (inp[9]) ? 4'b0011 : node11299;
														assign node11299 = (inp[5]) ? node11301 : 4'b0111;
															assign node11301 = (inp[3]) ? 4'b0101 : 4'b0111;
													assign node11305 = (inp[9]) ? node11311 : node11306;
														assign node11306 = (inp[3]) ? node11308 : 4'b0011;
															assign node11308 = (inp[5]) ? 4'b0001 : 4'b0011;
														assign node11311 = (inp[5]) ? 4'b0101 : node11312;
															assign node11312 = (inp[3]) ? 4'b0101 : 4'b0111;
									assign node11316 = (inp[10]) ? node11494 : node11317;
										assign node11317 = (inp[2]) ? node11399 : node11318;
											assign node11318 = (inp[0]) ? node11368 : node11319;
												assign node11319 = (inp[3]) ? node11347 : node11320;
													assign node11320 = (inp[15]) ? node11336 : node11321;
														assign node11321 = (inp[5]) ? node11329 : node11322;
															assign node11322 = (inp[9]) ? node11326 : node11323;
																assign node11323 = (inp[4]) ? 4'b0011 : 4'b0111;
																assign node11326 = (inp[4]) ? 4'b0111 : 4'b0011;
															assign node11329 = (inp[4]) ? node11333 : node11330;
																assign node11330 = (inp[9]) ? 4'b0011 : 4'b0111;
																assign node11333 = (inp[9]) ? 4'b0101 : 4'b0011;
														assign node11336 = (inp[5]) ? node11342 : node11337;
															assign node11337 = (inp[4]) ? node11339 : 4'b0001;
																assign node11339 = (inp[9]) ? 4'b0101 : 4'b0001;
															assign node11342 = (inp[4]) ? 4'b0111 : node11343;
																assign node11343 = (inp[9]) ? 4'b0001 : 4'b0101;
													assign node11347 = (inp[15]) ? node11359 : node11348;
														assign node11348 = (inp[5]) ? node11352 : node11349;
															assign node11349 = (inp[4]) ? 4'b0101 : 4'b0111;
															assign node11352 = (inp[9]) ? node11356 : node11353;
																assign node11353 = (inp[4]) ? 4'b0001 : 4'b0101;
																assign node11356 = (inp[4]) ? 4'b0101 : 4'b0001;
														assign node11359 = (inp[4]) ? node11365 : node11360;
															assign node11360 = (inp[5]) ? 4'b0011 : node11361;
																assign node11361 = (inp[9]) ? 4'b0001 : 4'b0101;
															assign node11365 = (inp[9]) ? 4'b0111 : 4'b0011;
												assign node11368 = (inp[15]) ? node11390 : node11369;
													assign node11369 = (inp[5]) ? node11377 : node11370;
														assign node11370 = (inp[3]) ? 4'b0001 : node11371;
															assign node11371 = (inp[9]) ? 4'b0001 : node11372;
																assign node11372 = (inp[4]) ? 4'b0001 : 4'b0101;
														assign node11377 = (inp[3]) ? node11385 : node11378;
															assign node11378 = (inp[4]) ? node11382 : node11379;
																assign node11379 = (inp[9]) ? 4'b0001 : 4'b0101;
																assign node11382 = (inp[9]) ? 4'b0111 : 4'b0001;
															assign node11385 = (inp[9]) ? node11387 : 4'b0111;
																assign node11387 = (inp[4]) ? 4'b0111 : 4'b0011;
													assign node11390 = (inp[4]) ? node11394 : node11391;
														assign node11391 = (inp[9]) ? 4'b0011 : 4'b0111;
														assign node11394 = (inp[9]) ? 4'b0101 : node11395;
															assign node11395 = (inp[5]) ? 4'b0001 : 4'b0011;
											assign node11399 = (inp[0]) ? node11447 : node11400;
												assign node11400 = (inp[15]) ? node11422 : node11401;
													assign node11401 = (inp[3]) ? node11409 : node11402;
														assign node11402 = (inp[4]) ? node11406 : node11403;
															assign node11403 = (inp[9]) ? 4'b0011 : 4'b0111;
															assign node11406 = (inp[9]) ? 4'b0101 : 4'b0011;
														assign node11409 = (inp[5]) ? node11415 : node11410;
															assign node11410 = (inp[9]) ? node11412 : 4'b0011;
																assign node11412 = (inp[4]) ? 4'b0101 : 4'b0011;
															assign node11415 = (inp[4]) ? node11419 : node11416;
																assign node11416 = (inp[9]) ? 4'b0001 : 4'b0101;
																assign node11419 = (inp[9]) ? 4'b0101 : 4'b0001;
													assign node11422 = (inp[3]) ? node11436 : node11423;
														assign node11423 = (inp[5]) ? node11431 : node11424;
															assign node11424 = (inp[9]) ? node11428 : node11425;
																assign node11425 = (inp[4]) ? 4'b0001 : 4'b0101;
																assign node11428 = (inp[4]) ? 4'b0101 : 4'b0001;
															assign node11431 = (inp[9]) ? 4'b0001 : node11432;
																assign node11432 = (inp[4]) ? 4'b0001 : 4'b0101;
														assign node11436 = (inp[5]) ? node11444 : node11437;
															assign node11437 = (inp[4]) ? node11441 : node11438;
																assign node11438 = (inp[9]) ? 4'b0001 : 4'b0101;
																assign node11441 = (inp[9]) ? 4'b0111 : 4'b0001;
															assign node11444 = (inp[9]) ? 4'b0111 : 4'b0011;
												assign node11447 = (inp[15]) ? node11473 : node11448;
													assign node11448 = (inp[5]) ? node11458 : node11449;
														assign node11449 = (inp[9]) ? node11453 : node11450;
															assign node11450 = (inp[4]) ? 4'b0001 : 4'b0101;
															assign node11453 = (inp[4]) ? node11455 : 4'b0001;
																assign node11455 = (inp[3]) ? 4'b0111 : 4'b0101;
														assign node11458 = (inp[3]) ? node11466 : node11459;
															assign node11459 = (inp[9]) ? node11463 : node11460;
																assign node11460 = (inp[4]) ? 4'b0001 : 4'b0101;
																assign node11463 = (inp[4]) ? 4'b0111 : 4'b0001;
															assign node11466 = (inp[4]) ? node11470 : node11467;
																assign node11467 = (inp[9]) ? 4'b0011 : 4'b0111;
																assign node11470 = (inp[9]) ? 4'b0111 : 4'b0011;
													assign node11473 = (inp[3]) ? node11481 : node11474;
														assign node11474 = (inp[4]) ? node11478 : node11475;
															assign node11475 = (inp[9]) ? 4'b0011 : 4'b0111;
															assign node11478 = (inp[5]) ? 4'b0101 : 4'b0011;
														assign node11481 = (inp[5]) ? node11487 : node11482;
															assign node11482 = (inp[9]) ? 4'b0101 : node11483;
																assign node11483 = (inp[4]) ? 4'b0011 : 4'b0111;
															assign node11487 = (inp[4]) ? node11491 : node11488;
																assign node11488 = (inp[9]) ? 4'b0001 : 4'b0101;
																assign node11491 = (inp[9]) ? 4'b0101 : 4'b0001;
										assign node11494 = (inp[9]) ? node11548 : node11495;
											assign node11495 = (inp[4]) ? node11525 : node11496;
												assign node11496 = (inp[3]) ? node11510 : node11497;
													assign node11497 = (inp[2]) ? node11503 : node11498;
														assign node11498 = (inp[0]) ? 4'b0011 : node11499;
															assign node11499 = (inp[15]) ? 4'b0001 : 4'b0011;
														assign node11503 = (inp[15]) ? node11507 : node11504;
															assign node11504 = (inp[0]) ? 4'b0001 : 4'b0011;
															assign node11507 = (inp[0]) ? 4'b0011 : 4'b0001;
													assign node11510 = (inp[5]) ? node11518 : node11511;
														assign node11511 = (inp[15]) ? node11515 : node11512;
															assign node11512 = (inp[0]) ? 4'b0001 : 4'b0011;
															assign node11515 = (inp[0]) ? 4'b0011 : 4'b0001;
														assign node11518 = (inp[0]) ? node11522 : node11519;
															assign node11519 = (inp[15]) ? 4'b0011 : 4'b0001;
															assign node11522 = (inp[15]) ? 4'b0001 : 4'b0011;
												assign node11525 = (inp[0]) ? node11537 : node11526;
													assign node11526 = (inp[15]) ? node11532 : node11527;
														assign node11527 = (inp[5]) ? 4'b0101 : node11528;
															assign node11528 = (inp[3]) ? 4'b0101 : 4'b0111;
														assign node11532 = (inp[5]) ? 4'b0111 : node11533;
															assign node11533 = (inp[3]) ? 4'b0111 : 4'b0101;
													assign node11537 = (inp[15]) ? node11543 : node11538;
														assign node11538 = (inp[5]) ? 4'b0111 : node11539;
															assign node11539 = (inp[3]) ? 4'b0111 : 4'b0101;
														assign node11543 = (inp[2]) ? 4'b0101 : node11544;
															assign node11544 = (inp[5]) ? 4'b0101 : 4'b0111;
											assign node11548 = (inp[4]) ? node11572 : node11549;
												assign node11549 = (inp[0]) ? node11561 : node11550;
													assign node11550 = (inp[5]) ? node11558 : node11551;
														assign node11551 = (inp[15]) ? node11555 : node11552;
															assign node11552 = (inp[3]) ? 4'b0101 : 4'b0111;
															assign node11555 = (inp[3]) ? 4'b0111 : 4'b0101;
														assign node11558 = (inp[15]) ? 4'b0111 : 4'b0101;
													assign node11561 = (inp[15]) ? node11567 : node11562;
														assign node11562 = (inp[5]) ? 4'b0111 : node11563;
															assign node11563 = (inp[3]) ? 4'b0111 : 4'b0101;
														assign node11567 = (inp[5]) ? 4'b0101 : node11568;
															assign node11568 = (inp[3]) ? 4'b0101 : 4'b0111;
												assign node11572 = (inp[5]) ? node11588 : node11573;
													assign node11573 = (inp[3]) ? node11581 : node11574;
														assign node11574 = (inp[0]) ? node11578 : node11575;
															assign node11575 = (inp[15]) ? 4'b0001 : 4'b0011;
															assign node11578 = (inp[15]) ? 4'b0011 : 4'b0001;
														assign node11581 = (inp[0]) ? node11585 : node11582;
															assign node11582 = (inp[15]) ? 4'b0011 : 4'b0001;
															assign node11585 = (inp[15]) ? 4'b0001 : 4'b0011;
													assign node11588 = (inp[3]) ? node11596 : node11589;
														assign node11589 = (inp[15]) ? node11593 : node11590;
															assign node11590 = (inp[0]) ? 4'b0011 : 4'b0001;
															assign node11593 = (inp[0]) ? 4'b0001 : 4'b0011;
														assign node11596 = (inp[2]) ? node11602 : node11597;
															assign node11597 = (inp[0]) ? node11599 : 4'b0011;
																assign node11599 = (inp[15]) ? 4'b0001 : 4'b0011;
															assign node11602 = (inp[0]) ? 4'b0011 : node11603;
																assign node11603 = (inp[15]) ? 4'b0011 : 4'b0001;
							assign node11607 = (inp[2]) ? node12087 : node11608;
								assign node11608 = (inp[14]) ? node11814 : node11609;
									assign node11609 = (inp[4]) ? node11711 : node11610;
										assign node11610 = (inp[9]) ? node11664 : node11611;
											assign node11611 = (inp[12]) ? node11633 : node11612;
												assign node11612 = (inp[15]) ? node11624 : node11613;
													assign node11613 = (inp[0]) ? node11619 : node11614;
														assign node11614 = (inp[3]) ? node11616 : 4'b0111;
															assign node11616 = (inp[5]) ? 4'b0101 : 4'b0111;
														assign node11619 = (inp[5]) ? node11621 : 4'b0101;
															assign node11621 = (inp[3]) ? 4'b0111 : 4'b0101;
													assign node11624 = (inp[0]) ? node11630 : node11625;
														assign node11625 = (inp[5]) ? node11627 : 4'b0101;
															assign node11627 = (inp[3]) ? 4'b0111 : 4'b0101;
														assign node11630 = (inp[10]) ? 4'b0101 : 4'b0111;
												assign node11633 = (inp[10]) ? node11651 : node11634;
													assign node11634 = (inp[15]) ? node11646 : node11635;
														assign node11635 = (inp[0]) ? node11641 : node11636;
															assign node11636 = (inp[5]) ? node11638 : 4'b0111;
																assign node11638 = (inp[3]) ? 4'b0101 : 4'b0111;
															assign node11641 = (inp[5]) ? node11643 : 4'b0101;
																assign node11643 = (inp[3]) ? 4'b0111 : 4'b0101;
														assign node11646 = (inp[0]) ? 4'b0111 : node11647;
															assign node11647 = (inp[5]) ? 4'b0111 : 4'b0101;
													assign node11651 = (inp[3]) ? node11659 : node11652;
														assign node11652 = (inp[0]) ? node11656 : node11653;
															assign node11653 = (inp[15]) ? 4'b0001 : 4'b0011;
															assign node11656 = (inp[15]) ? 4'b0011 : 4'b0001;
														assign node11659 = (inp[15]) ? node11661 : 4'b0001;
															assign node11661 = (inp[5]) ? 4'b0001 : 4'b0011;
											assign node11664 = (inp[10]) ? node11688 : node11665;
												assign node11665 = (inp[15]) ? node11677 : node11666;
													assign node11666 = (inp[0]) ? node11672 : node11667;
														assign node11667 = (inp[3]) ? node11669 : 4'b0011;
															assign node11669 = (inp[5]) ? 4'b0001 : 4'b0011;
														assign node11672 = (inp[3]) ? node11674 : 4'b0001;
															assign node11674 = (inp[5]) ? 4'b0011 : 4'b0001;
													assign node11677 = (inp[0]) ? node11683 : node11678;
														assign node11678 = (inp[5]) ? node11680 : 4'b0001;
															assign node11680 = (inp[3]) ? 4'b0011 : 4'b0001;
														assign node11683 = (inp[5]) ? node11685 : 4'b0011;
															assign node11685 = (inp[3]) ? 4'b0001 : 4'b0011;
												assign node11688 = (inp[12]) ? node11702 : node11689;
													assign node11689 = (inp[0]) ? node11697 : node11690;
														assign node11690 = (inp[15]) ? 4'b0001 : node11691;
															assign node11691 = (inp[3]) ? node11693 : 4'b0011;
																assign node11693 = (inp[5]) ? 4'b0001 : 4'b0011;
														assign node11697 = (inp[15]) ? node11699 : 4'b0001;
															assign node11699 = (inp[5]) ? 4'b0001 : 4'b0011;
													assign node11702 = (inp[0]) ? node11706 : node11703;
														assign node11703 = (inp[15]) ? 4'b0111 : 4'b0101;
														assign node11706 = (inp[3]) ? node11708 : 4'b0101;
															assign node11708 = (inp[15]) ? 4'b0101 : 4'b0111;
										assign node11711 = (inp[9]) ? node11761 : node11712;
											assign node11712 = (inp[12]) ? node11730 : node11713;
												assign node11713 = (inp[15]) ? node11725 : node11714;
													assign node11714 = (inp[0]) ? node11720 : node11715;
														assign node11715 = (inp[5]) ? node11717 : 4'b0011;
															assign node11717 = (inp[3]) ? 4'b0001 : 4'b0011;
														assign node11720 = (inp[3]) ? node11722 : 4'b0001;
															assign node11722 = (inp[5]) ? 4'b0011 : 4'b0001;
													assign node11725 = (inp[0]) ? 4'b0011 : node11726;
														assign node11726 = (inp[3]) ? 4'b0011 : 4'b0001;
												assign node11730 = (inp[10]) ? node11742 : node11731;
													assign node11731 = (inp[15]) ? node11733 : 4'b0001;
														assign node11733 = (inp[0]) ? node11739 : node11734;
															assign node11734 = (inp[3]) ? node11736 : 4'b0001;
																assign node11736 = (inp[5]) ? 4'b0011 : 4'b0001;
															assign node11739 = (inp[5]) ? 4'b0001 : 4'b0011;
													assign node11742 = (inp[15]) ? node11750 : node11743;
														assign node11743 = (inp[0]) ? 4'b0111 : node11744;
															assign node11744 = (inp[5]) ? 4'b0101 : node11745;
																assign node11745 = (inp[3]) ? 4'b0101 : 4'b0111;
														assign node11750 = (inp[0]) ? node11756 : node11751;
															assign node11751 = (inp[3]) ? 4'b0111 : node11752;
																assign node11752 = (inp[5]) ? 4'b0111 : 4'b0101;
															assign node11756 = (inp[5]) ? 4'b0101 : node11757;
																assign node11757 = (inp[3]) ? 4'b0101 : 4'b0111;
											assign node11761 = (inp[12]) ? node11785 : node11762;
												assign node11762 = (inp[15]) ? node11774 : node11763;
													assign node11763 = (inp[0]) ? node11769 : node11764;
														assign node11764 = (inp[3]) ? 4'b0101 : node11765;
															assign node11765 = (inp[10]) ? 4'b0101 : 4'b0111;
														assign node11769 = (inp[5]) ? 4'b0111 : node11770;
															assign node11770 = (inp[3]) ? 4'b0111 : 4'b0101;
													assign node11774 = (inp[0]) ? node11780 : node11775;
														assign node11775 = (inp[5]) ? 4'b0111 : node11776;
															assign node11776 = (inp[3]) ? 4'b0111 : 4'b0101;
														assign node11780 = (inp[5]) ? 4'b0101 : node11781;
															assign node11781 = (inp[3]) ? 4'b0101 : 4'b0111;
												assign node11785 = (inp[10]) ? node11799 : node11786;
													assign node11786 = (inp[15]) ? node11794 : node11787;
														assign node11787 = (inp[0]) ? 4'b0111 : node11788;
															assign node11788 = (inp[5]) ? 4'b0101 : node11789;
																assign node11789 = (inp[3]) ? 4'b0101 : 4'b0111;
														assign node11794 = (inp[0]) ? 4'b0101 : node11795;
															assign node11795 = (inp[3]) ? 4'b0111 : 4'b0101;
													assign node11799 = (inp[0]) ? node11809 : node11800;
														assign node11800 = (inp[15]) ? node11806 : node11801;
															assign node11801 = (inp[3]) ? 4'b0001 : node11802;
																assign node11802 = (inp[5]) ? 4'b0001 : 4'b0011;
															assign node11806 = (inp[5]) ? 4'b0011 : 4'b0001;
														assign node11809 = (inp[15]) ? node11811 : 4'b0011;
															assign node11811 = (inp[5]) ? 4'b0001 : 4'b0011;
									assign node11814 = (inp[15]) ? node11960 : node11815;
										assign node11815 = (inp[5]) ? node11879 : node11816;
											assign node11816 = (inp[0]) ? node11848 : node11817;
												assign node11817 = (inp[3]) ? node11827 : node11818;
													assign node11818 = (inp[10]) ? node11820 : 4'b0010;
														assign node11820 = (inp[12]) ? node11822 : 4'b0110;
															assign node11822 = (inp[4]) ? node11824 : 4'b0010;
																assign node11824 = (inp[9]) ? 4'b0010 : 4'b0110;
													assign node11827 = (inp[4]) ? node11839 : node11828;
														assign node11828 = (inp[9]) ? node11834 : node11829;
															assign node11829 = (inp[12]) ? node11831 : 4'b0110;
																assign node11831 = (inp[10]) ? 4'b0010 : 4'b0110;
															assign node11834 = (inp[12]) ? node11836 : 4'b0010;
																assign node11836 = (inp[10]) ? 4'b0100 : 4'b0010;
														assign node11839 = (inp[9]) ? node11845 : node11840;
															assign node11840 = (inp[10]) ? node11842 : 4'b0010;
																assign node11842 = (inp[12]) ? 4'b0100 : 4'b0010;
															assign node11845 = (inp[10]) ? 4'b0000 : 4'b0100;
												assign node11848 = (inp[3]) ? node11858 : node11849;
													assign node11849 = (inp[12]) ? 4'b0000 : node11850;
														assign node11850 = (inp[9]) ? node11854 : node11851;
															assign node11851 = (inp[4]) ? 4'b0000 : 4'b0100;
															assign node11854 = (inp[4]) ? 4'b0100 : 4'b0000;
													assign node11858 = (inp[9]) ? node11870 : node11859;
														assign node11859 = (inp[4]) ? node11865 : node11860;
															assign node11860 = (inp[10]) ? node11862 : 4'b0100;
																assign node11862 = (inp[12]) ? 4'b0000 : 4'b0100;
															assign node11865 = (inp[10]) ? node11867 : 4'b0000;
																assign node11867 = (inp[12]) ? 4'b0110 : 4'b0000;
														assign node11870 = (inp[4]) ? node11876 : node11871;
															assign node11871 = (inp[12]) ? node11873 : 4'b0000;
																assign node11873 = (inp[10]) ? 4'b0110 : 4'b0000;
															assign node11876 = (inp[10]) ? 4'b0010 : 4'b0110;
											assign node11879 = (inp[0]) ? node11919 : node11880;
												assign node11880 = (inp[3]) ? node11898 : node11881;
													assign node11881 = (inp[9]) ? node11891 : node11882;
														assign node11882 = (inp[4]) ? node11886 : node11883;
															assign node11883 = (inp[12]) ? 4'b0010 : 4'b0110;
															assign node11886 = (inp[10]) ? node11888 : 4'b0010;
																assign node11888 = (inp[12]) ? 4'b0100 : 4'b0010;
														assign node11891 = (inp[4]) ? node11895 : node11892;
															assign node11892 = (inp[12]) ? 4'b0100 : 4'b0010;
															assign node11895 = (inp[12]) ? 4'b0000 : 4'b0100;
													assign node11898 = (inp[12]) ? node11906 : node11899;
														assign node11899 = (inp[9]) ? node11903 : node11900;
															assign node11900 = (inp[4]) ? 4'b0000 : 4'b0100;
															assign node11903 = (inp[4]) ? 4'b0100 : 4'b0000;
														assign node11906 = (inp[4]) ? node11912 : node11907;
															assign node11907 = (inp[9]) ? node11909 : 4'b0100;
																assign node11909 = (inp[10]) ? 4'b0100 : 4'b0000;
															assign node11912 = (inp[9]) ? node11916 : node11913;
																assign node11913 = (inp[10]) ? 4'b0100 : 4'b0000;
																assign node11916 = (inp[10]) ? 4'b0000 : 4'b0100;
												assign node11919 = (inp[3]) ? node11939 : node11920;
													assign node11920 = (inp[4]) ? node11930 : node11921;
														assign node11921 = (inp[10]) ? node11923 : 4'b0000;
															assign node11923 = (inp[12]) ? node11927 : node11924;
																assign node11924 = (inp[9]) ? 4'b0000 : 4'b0100;
																assign node11927 = (inp[9]) ? 4'b0110 : 4'b0000;
														assign node11930 = (inp[9]) ? node11934 : node11931;
															assign node11931 = (inp[10]) ? 4'b0110 : 4'b0000;
															assign node11934 = (inp[12]) ? node11936 : 4'b0110;
																assign node11936 = (inp[10]) ? 4'b0010 : 4'b0110;
													assign node11939 = (inp[4]) ? node11949 : node11940;
														assign node11940 = (inp[9]) ? node11946 : node11941;
															assign node11941 = (inp[10]) ? node11943 : 4'b0110;
																assign node11943 = (inp[12]) ? 4'b0010 : 4'b0110;
															assign node11946 = (inp[12]) ? 4'b0110 : 4'b0010;
														assign node11949 = (inp[9]) ? node11955 : node11950;
															assign node11950 = (inp[10]) ? node11952 : 4'b0010;
																assign node11952 = (inp[12]) ? 4'b0110 : 4'b0010;
															assign node11955 = (inp[12]) ? node11957 : 4'b0110;
																assign node11957 = (inp[10]) ? 4'b0010 : 4'b0110;
										assign node11960 = (inp[0]) ? node12030 : node11961;
											assign node11961 = (inp[5]) ? node12001 : node11962;
												assign node11962 = (inp[3]) ? node11980 : node11963;
													assign node11963 = (inp[9]) ? node11971 : node11964;
														assign node11964 = (inp[12]) ? node11968 : node11965;
															assign node11965 = (inp[4]) ? 4'b0000 : 4'b0100;
															assign node11968 = (inp[4]) ? 4'b0100 : 4'b0000;
														assign node11971 = (inp[12]) ? node11973 : 4'b0100;
															assign node11973 = (inp[10]) ? node11977 : node11974;
																assign node11974 = (inp[4]) ? 4'b0100 : 4'b0000;
																assign node11977 = (inp[4]) ? 4'b0000 : 4'b0100;
													assign node11980 = (inp[9]) ? node11992 : node11981;
														assign node11981 = (inp[4]) ? node11987 : node11982;
															assign node11982 = (inp[10]) ? node11984 : 4'b0100;
																assign node11984 = (inp[12]) ? 4'b0000 : 4'b0100;
															assign node11987 = (inp[10]) ? node11989 : 4'b0000;
																assign node11989 = (inp[12]) ? 4'b0110 : 4'b0000;
														assign node11992 = (inp[12]) ? node11994 : 4'b0110;
															assign node11994 = (inp[4]) ? node11998 : node11995;
																assign node11995 = (inp[10]) ? 4'b0110 : 4'b0000;
																assign node11998 = (inp[10]) ? 4'b0010 : 4'b0110;
												assign node12001 = (inp[3]) ? node12015 : node12002;
													assign node12002 = (inp[9]) ? node12010 : node12003;
														assign node12003 = (inp[10]) ? node12007 : node12004;
															assign node12004 = (inp[4]) ? 4'b0000 : 4'b0100;
															assign node12007 = (inp[4]) ? 4'b0110 : 4'b0000;
														assign node12010 = (inp[4]) ? 4'b0110 : node12011;
															assign node12011 = (inp[12]) ? 4'b0110 : 4'b0000;
													assign node12015 = (inp[10]) ? node12023 : node12016;
														assign node12016 = (inp[4]) ? node12020 : node12017;
															assign node12017 = (inp[9]) ? 4'b0010 : 4'b0110;
															assign node12020 = (inp[9]) ? 4'b0110 : 4'b0010;
														assign node12023 = (inp[4]) ? node12027 : node12024;
															assign node12024 = (inp[12]) ? 4'b0110 : 4'b0010;
															assign node12027 = (inp[12]) ? 4'b0010 : 4'b0110;
											assign node12030 = (inp[5]) ? node12056 : node12031;
												assign node12031 = (inp[4]) ? node12043 : node12032;
													assign node12032 = (inp[9]) ? node12038 : node12033;
														assign node12033 = (inp[12]) ? node12035 : 4'b0110;
															assign node12035 = (inp[10]) ? 4'b0010 : 4'b0110;
														assign node12038 = (inp[12]) ? node12040 : 4'b0010;
															assign node12040 = (inp[10]) ? 4'b0110 : 4'b0010;
													assign node12043 = (inp[9]) ? node12049 : node12044;
														assign node12044 = (inp[12]) ? node12046 : 4'b0010;
															assign node12046 = (inp[10]) ? 4'b0110 : 4'b0010;
														assign node12049 = (inp[3]) ? 4'b0100 : node12050;
															assign node12050 = (inp[12]) ? node12052 : 4'b0110;
																assign node12052 = (inp[10]) ? 4'b0010 : 4'b0110;
												assign node12056 = (inp[3]) ? node12072 : node12057;
													assign node12057 = (inp[9]) ? node12065 : node12058;
														assign node12058 = (inp[4]) ? node12060 : 4'b0110;
															assign node12060 = (inp[12]) ? node12062 : 4'b0010;
																assign node12062 = (inp[10]) ? 4'b0100 : 4'b0010;
														assign node12065 = (inp[4]) ? node12069 : node12066;
															assign node12066 = (inp[12]) ? 4'b0100 : 4'b0010;
															assign node12069 = (inp[12]) ? 4'b0000 : 4'b0100;
													assign node12072 = (inp[9]) ? node12078 : node12073;
														assign node12073 = (inp[4]) ? 4'b0000 : node12074;
															assign node12074 = (inp[12]) ? 4'b0000 : 4'b0100;
														assign node12078 = (inp[12]) ? node12082 : node12079;
															assign node12079 = (inp[4]) ? 4'b0100 : 4'b0000;
															assign node12082 = (inp[4]) ? node12084 : 4'b0100;
																assign node12084 = (inp[10]) ? 4'b0000 : 4'b0100;
								assign node12087 = (inp[9]) ? node12265 : node12088;
									assign node12088 = (inp[4]) ? node12166 : node12089;
										assign node12089 = (inp[12]) ? node12113 : node12090;
											assign node12090 = (inp[15]) ? node12102 : node12091;
												assign node12091 = (inp[0]) ? node12097 : node12092;
													assign node12092 = (inp[3]) ? node12094 : 4'b0110;
														assign node12094 = (inp[5]) ? 4'b0100 : 4'b0110;
													assign node12097 = (inp[5]) ? node12099 : 4'b0100;
														assign node12099 = (inp[3]) ? 4'b0110 : 4'b0100;
												assign node12102 = (inp[0]) ? node12108 : node12103;
													assign node12103 = (inp[3]) ? node12105 : 4'b0100;
														assign node12105 = (inp[5]) ? 4'b0110 : 4'b0100;
													assign node12108 = (inp[5]) ? node12110 : 4'b0110;
														assign node12110 = (inp[3]) ? 4'b0100 : 4'b0110;
											assign node12113 = (inp[10]) ? node12137 : node12114;
												assign node12114 = (inp[0]) ? node12126 : node12115;
													assign node12115 = (inp[15]) ? node12121 : node12116;
														assign node12116 = (inp[5]) ? node12118 : 4'b0110;
															assign node12118 = (inp[3]) ? 4'b0100 : 4'b0110;
														assign node12121 = (inp[3]) ? node12123 : 4'b0100;
															assign node12123 = (inp[5]) ? 4'b0110 : 4'b0100;
													assign node12126 = (inp[15]) ? node12132 : node12127;
														assign node12127 = (inp[5]) ? node12129 : 4'b0100;
															assign node12129 = (inp[3]) ? 4'b0110 : 4'b0100;
														assign node12132 = (inp[5]) ? node12134 : 4'b0110;
															assign node12134 = (inp[3]) ? 4'b0100 : 4'b0110;
												assign node12137 = (inp[3]) ? node12153 : node12138;
													assign node12138 = (inp[5]) ? node12148 : node12139;
														assign node12139 = (inp[14]) ? 4'b0000 : node12140;
															assign node12140 = (inp[0]) ? node12144 : node12141;
																assign node12141 = (inp[15]) ? 4'b0000 : 4'b0010;
																assign node12144 = (inp[15]) ? 4'b0010 : 4'b0000;
														assign node12148 = (inp[0]) ? node12150 : 4'b0000;
															assign node12150 = (inp[15]) ? 4'b0010 : 4'b0000;
													assign node12153 = (inp[15]) ? node12161 : node12154;
														assign node12154 = (inp[0]) ? node12158 : node12155;
															assign node12155 = (inp[5]) ? 4'b0000 : 4'b0010;
															assign node12158 = (inp[5]) ? 4'b0010 : 4'b0000;
														assign node12161 = (inp[0]) ? 4'b0000 : node12162;
															assign node12162 = (inp[5]) ? 4'b0010 : 4'b0000;
										assign node12166 = (inp[12]) ? node12190 : node12167;
											assign node12167 = (inp[0]) ? node12179 : node12168;
												assign node12168 = (inp[15]) ? node12174 : node12169;
													assign node12169 = (inp[3]) ? node12171 : 4'b0010;
														assign node12171 = (inp[5]) ? 4'b0000 : 4'b0010;
													assign node12174 = (inp[3]) ? node12176 : 4'b0000;
														assign node12176 = (inp[5]) ? 4'b0010 : 4'b0000;
												assign node12179 = (inp[15]) ? node12185 : node12180;
													assign node12180 = (inp[5]) ? node12182 : 4'b0000;
														assign node12182 = (inp[3]) ? 4'b0010 : 4'b0000;
													assign node12185 = (inp[5]) ? node12187 : 4'b0010;
														assign node12187 = (inp[3]) ? 4'b0000 : 4'b0010;
											assign node12190 = (inp[10]) ? node12228 : node12191;
												assign node12191 = (inp[5]) ? node12213 : node12192;
													assign node12192 = (inp[14]) ? node12206 : node12193;
														assign node12193 = (inp[3]) ? node12201 : node12194;
															assign node12194 = (inp[15]) ? node12198 : node12195;
																assign node12195 = (inp[0]) ? 4'b0000 : 4'b0010;
																assign node12198 = (inp[0]) ? 4'b0010 : 4'b0000;
															assign node12201 = (inp[15]) ? 4'b0000 : node12202;
																assign node12202 = (inp[0]) ? 4'b0000 : 4'b0010;
														assign node12206 = (inp[3]) ? 4'b0010 : node12207;
															assign node12207 = (inp[15]) ? 4'b0010 : node12208;
																assign node12208 = (inp[0]) ? 4'b0000 : 4'b0010;
													assign node12213 = (inp[3]) ? node12221 : node12214;
														assign node12214 = (inp[14]) ? node12218 : node12215;
															assign node12215 = (inp[0]) ? 4'b0000 : 4'b0010;
															assign node12218 = (inp[0]) ? 4'b0010 : 4'b0000;
														assign node12221 = (inp[14]) ? 4'b0000 : node12222;
															assign node12222 = (inp[15]) ? 4'b0000 : node12223;
																assign node12223 = (inp[0]) ? 4'b0010 : 4'b0000;
												assign node12228 = (inp[5]) ? node12244 : node12229;
													assign node12229 = (inp[15]) ? node12237 : node12230;
														assign node12230 = (inp[0]) ? node12234 : node12231;
															assign node12231 = (inp[3]) ? 4'b0100 : 4'b0110;
															assign node12234 = (inp[3]) ? 4'b0110 : 4'b0100;
														assign node12237 = (inp[3]) ? node12241 : node12238;
															assign node12238 = (inp[0]) ? 4'b0110 : 4'b0100;
															assign node12241 = (inp[0]) ? 4'b0100 : 4'b0110;
													assign node12244 = (inp[3]) ? node12260 : node12245;
														assign node12245 = (inp[14]) ? node12253 : node12246;
															assign node12246 = (inp[0]) ? node12250 : node12247;
																assign node12247 = (inp[15]) ? 4'b0110 : 4'b0100;
																assign node12250 = (inp[15]) ? 4'b0100 : 4'b0110;
															assign node12253 = (inp[15]) ? node12257 : node12254;
																assign node12254 = (inp[0]) ? 4'b0110 : 4'b0100;
																assign node12257 = (inp[0]) ? 4'b0100 : 4'b0110;
														assign node12260 = (inp[15]) ? node12262 : 4'b0110;
															assign node12262 = (inp[0]) ? 4'b0100 : 4'b0110;
									assign node12265 = (inp[4]) ? node12379 : node12266;
										assign node12266 = (inp[12]) ? node12306 : node12267;
											assign node12267 = (inp[3]) ? node12275 : node12268;
												assign node12268 = (inp[0]) ? node12272 : node12269;
													assign node12269 = (inp[15]) ? 4'b0000 : 4'b0010;
													assign node12272 = (inp[15]) ? 4'b0010 : 4'b0000;
												assign node12275 = (inp[15]) ? node12299 : node12276;
													assign node12276 = (inp[10]) ? node12284 : node12277;
														assign node12277 = (inp[0]) ? node12281 : node12278;
															assign node12278 = (inp[5]) ? 4'b0000 : 4'b0010;
															assign node12281 = (inp[5]) ? 4'b0010 : 4'b0000;
														assign node12284 = (inp[14]) ? node12292 : node12285;
															assign node12285 = (inp[5]) ? node12289 : node12286;
																assign node12286 = (inp[0]) ? 4'b0000 : 4'b0010;
																assign node12289 = (inp[0]) ? 4'b0010 : 4'b0000;
															assign node12292 = (inp[0]) ? node12296 : node12293;
																assign node12293 = (inp[5]) ? 4'b0000 : 4'b0010;
																assign node12296 = (inp[5]) ? 4'b0010 : 4'b0000;
													assign node12299 = (inp[0]) ? node12303 : node12300;
														assign node12300 = (inp[5]) ? 4'b0010 : 4'b0000;
														assign node12303 = (inp[5]) ? 4'b0000 : 4'b0010;
											assign node12306 = (inp[10]) ? node12352 : node12307;
												assign node12307 = (inp[14]) ? node12325 : node12308;
													assign node12308 = (inp[5]) ? node12314 : node12309;
														assign node12309 = (inp[0]) ? 4'b0010 : node12310;
															assign node12310 = (inp[15]) ? 4'b0000 : 4'b0010;
														assign node12314 = (inp[0]) ? node12320 : node12315;
															assign node12315 = (inp[3]) ? 4'b0010 : node12316;
																assign node12316 = (inp[15]) ? 4'b0000 : 4'b0010;
															assign node12320 = (inp[3]) ? 4'b0000 : node12321;
																assign node12321 = (inp[15]) ? 4'b0010 : 4'b0000;
													assign node12325 = (inp[5]) ? node12339 : node12326;
														assign node12326 = (inp[3]) ? node12334 : node12327;
															assign node12327 = (inp[0]) ? node12331 : node12328;
																assign node12328 = (inp[15]) ? 4'b0000 : 4'b0010;
																assign node12331 = (inp[15]) ? 4'b0010 : 4'b0000;
															assign node12334 = (inp[0]) ? node12336 : 4'b0000;
																assign node12336 = (inp[15]) ? 4'b0010 : 4'b0000;
														assign node12339 = (inp[3]) ? node12347 : node12340;
															assign node12340 = (inp[15]) ? node12344 : node12341;
																assign node12341 = (inp[0]) ? 4'b0000 : 4'b0010;
																assign node12344 = (inp[0]) ? 4'b0010 : 4'b0000;
															assign node12347 = (inp[15]) ? node12349 : 4'b0010;
																assign node12349 = (inp[0]) ? 4'b0000 : 4'b0010;
												assign node12352 = (inp[5]) ? node12372 : node12353;
													assign node12353 = (inp[3]) ? node12367 : node12354;
														assign node12354 = (inp[14]) ? node12362 : node12355;
															assign node12355 = (inp[0]) ? node12359 : node12356;
																assign node12356 = (inp[15]) ? 4'b0100 : 4'b0110;
																assign node12359 = (inp[15]) ? 4'b0110 : 4'b0100;
															assign node12362 = (inp[15]) ? node12364 : 4'b0100;
																assign node12364 = (inp[0]) ? 4'b0110 : 4'b0100;
														assign node12367 = (inp[15]) ? 4'b0100 : node12368;
															assign node12368 = (inp[0]) ? 4'b0110 : 4'b0100;
													assign node12372 = (inp[0]) ? node12376 : node12373;
														assign node12373 = (inp[15]) ? 4'b0110 : 4'b0100;
														assign node12376 = (inp[15]) ? 4'b0100 : 4'b0110;
										assign node12379 = (inp[12]) ? node12403 : node12380;
											assign node12380 = (inp[0]) ? node12392 : node12381;
												assign node12381 = (inp[15]) ? node12387 : node12382;
													assign node12382 = (inp[3]) ? 4'b0100 : node12383;
														assign node12383 = (inp[5]) ? 4'b0100 : 4'b0110;
													assign node12387 = (inp[5]) ? 4'b0110 : node12388;
														assign node12388 = (inp[3]) ? 4'b0110 : 4'b0100;
												assign node12392 = (inp[15]) ? node12398 : node12393;
													assign node12393 = (inp[5]) ? 4'b0110 : node12394;
														assign node12394 = (inp[3]) ? 4'b0110 : 4'b0100;
													assign node12398 = (inp[5]) ? 4'b0100 : node12399;
														assign node12399 = (inp[3]) ? 4'b0100 : 4'b0110;
											assign node12403 = (inp[10]) ? node12425 : node12404;
												assign node12404 = (inp[3]) ? node12418 : node12405;
													assign node12405 = (inp[0]) ? node12413 : node12406;
														assign node12406 = (inp[15]) ? node12410 : node12407;
															assign node12407 = (inp[5]) ? 4'b0100 : 4'b0110;
															assign node12410 = (inp[5]) ? 4'b0110 : 4'b0100;
														assign node12413 = (inp[14]) ? 4'b0110 : node12414;
															assign node12414 = (inp[15]) ? 4'b0100 : 4'b0110;
													assign node12418 = (inp[15]) ? node12422 : node12419;
														assign node12419 = (inp[0]) ? 4'b0110 : 4'b0100;
														assign node12422 = (inp[0]) ? 4'b0100 : 4'b0110;
												assign node12425 = (inp[3]) ? node12445 : node12426;
													assign node12426 = (inp[0]) ? node12434 : node12427;
														assign node12427 = (inp[14]) ? node12431 : node12428;
															assign node12428 = (inp[5]) ? 4'b0010 : 4'b0000;
															assign node12431 = (inp[5]) ? 4'b0000 : 4'b0010;
														assign node12434 = (inp[14]) ? node12440 : node12435;
															assign node12435 = (inp[15]) ? 4'b0000 : node12436;
																assign node12436 = (inp[5]) ? 4'b0010 : 4'b0000;
															assign node12440 = (inp[5]) ? 4'b0000 : node12441;
																assign node12441 = (inp[15]) ? 4'b0010 : 4'b0000;
													assign node12445 = (inp[15]) ? node12449 : node12446;
														assign node12446 = (inp[0]) ? 4'b0010 : 4'b0000;
														assign node12449 = (inp[0]) ? 4'b0000 : 4'b0010;
					assign node12452 = (inp[9]) ? node14496 : node12453;
						assign node12453 = (inp[4]) ? node13397 : node12454;
							assign node12454 = (inp[12]) ? node12838 : node12455;
								assign node12455 = (inp[14]) ? node12675 : node12456;
									assign node12456 = (inp[8]) ? node12574 : node12457;
										assign node12457 = (inp[15]) ? node12511 : node12458;
											assign node12458 = (inp[0]) ? node12484 : node12459;
												assign node12459 = (inp[5]) ? node12467 : node12460;
													assign node12460 = (inp[7]) ? node12464 : node12461;
														assign node12461 = (inp[2]) ? 4'b0110 : 4'b0111;
														assign node12464 = (inp[2]) ? 4'b0111 : 4'b0110;
													assign node12467 = (inp[3]) ? node12477 : node12468;
														assign node12468 = (inp[10]) ? node12470 : 4'b0111;
															assign node12470 = (inp[2]) ? node12474 : node12471;
																assign node12471 = (inp[7]) ? 4'b0110 : 4'b0111;
																assign node12474 = (inp[7]) ? 4'b0111 : 4'b0110;
														assign node12477 = (inp[2]) ? node12481 : node12478;
															assign node12478 = (inp[7]) ? 4'b0100 : 4'b0101;
															assign node12481 = (inp[7]) ? 4'b0101 : 4'b0100;
												assign node12484 = (inp[3]) ? node12498 : node12485;
													assign node12485 = (inp[5]) ? node12493 : node12486;
														assign node12486 = (inp[10]) ? node12488 : 4'b0100;
															assign node12488 = (inp[2]) ? 4'b0101 : node12489;
																assign node12489 = (inp[7]) ? 4'b0100 : 4'b0101;
														assign node12493 = (inp[7]) ? node12495 : 4'b0101;
															assign node12495 = (inp[2]) ? 4'b0101 : 4'b0100;
													assign node12498 = (inp[5]) ? node12504 : node12499;
														assign node12499 = (inp[2]) ? node12501 : 4'b0101;
															assign node12501 = (inp[7]) ? 4'b0101 : 4'b0100;
														assign node12504 = (inp[7]) ? node12508 : node12505;
															assign node12505 = (inp[2]) ? 4'b0110 : 4'b0111;
															assign node12508 = (inp[2]) ? 4'b0111 : 4'b0110;
											assign node12511 = (inp[0]) ? node12545 : node12512;
												assign node12512 = (inp[5]) ? node12528 : node12513;
													assign node12513 = (inp[3]) ? node12521 : node12514;
														assign node12514 = (inp[7]) ? node12518 : node12515;
															assign node12515 = (inp[2]) ? 4'b0100 : 4'b0101;
															assign node12518 = (inp[2]) ? 4'b0101 : 4'b0100;
														assign node12521 = (inp[2]) ? node12525 : node12522;
															assign node12522 = (inp[7]) ? 4'b0100 : 4'b0101;
															assign node12525 = (inp[7]) ? 4'b0101 : 4'b0100;
													assign node12528 = (inp[3]) ? node12536 : node12529;
														assign node12529 = (inp[7]) ? node12533 : node12530;
															assign node12530 = (inp[2]) ? 4'b0100 : 4'b0101;
															assign node12533 = (inp[2]) ? 4'b0101 : 4'b0100;
														assign node12536 = (inp[10]) ? 4'b0111 : node12537;
															assign node12537 = (inp[2]) ? node12541 : node12538;
																assign node12538 = (inp[7]) ? 4'b0110 : 4'b0111;
																assign node12541 = (inp[7]) ? 4'b0111 : 4'b0110;
												assign node12545 = (inp[3]) ? node12561 : node12546;
													assign node12546 = (inp[5]) ? node12554 : node12547;
														assign node12547 = (inp[2]) ? node12551 : node12548;
															assign node12548 = (inp[7]) ? 4'b0110 : 4'b0111;
															assign node12551 = (inp[7]) ? 4'b0111 : 4'b0110;
														assign node12554 = (inp[7]) ? node12558 : node12555;
															assign node12555 = (inp[2]) ? 4'b0110 : 4'b0111;
															assign node12558 = (inp[2]) ? 4'b0111 : 4'b0110;
													assign node12561 = (inp[5]) ? node12567 : node12562;
														assign node12562 = (inp[7]) ? node12564 : 4'b0111;
															assign node12564 = (inp[2]) ? 4'b0111 : 4'b0110;
														assign node12567 = (inp[2]) ? node12571 : node12568;
															assign node12568 = (inp[7]) ? 4'b0100 : 4'b0101;
															assign node12571 = (inp[7]) ? 4'b0101 : 4'b0100;
										assign node12574 = (inp[2]) ? node12634 : node12575;
											assign node12575 = (inp[7]) ? node12599 : node12576;
												assign node12576 = (inp[0]) ? node12588 : node12577;
													assign node12577 = (inp[15]) ? node12583 : node12578;
														assign node12578 = (inp[3]) ? node12580 : 4'b0110;
															assign node12580 = (inp[5]) ? 4'b0100 : 4'b0110;
														assign node12583 = (inp[5]) ? node12585 : 4'b0100;
															assign node12585 = (inp[3]) ? 4'b0110 : 4'b0100;
													assign node12588 = (inp[15]) ? node12594 : node12589;
														assign node12589 = (inp[10]) ? 4'b0100 : node12590;
															assign node12590 = (inp[3]) ? 4'b0110 : 4'b0100;
														assign node12594 = (inp[3]) ? node12596 : 4'b0110;
															assign node12596 = (inp[5]) ? 4'b0100 : 4'b0110;
												assign node12599 = (inp[5]) ? node12623 : node12600;
													assign node12600 = (inp[10]) ? node12610 : node12601;
														assign node12601 = (inp[3]) ? 4'b0101 : node12602;
															assign node12602 = (inp[15]) ? node12606 : node12603;
																assign node12603 = (inp[0]) ? 4'b0101 : 4'b0111;
																assign node12606 = (inp[0]) ? 4'b0111 : 4'b0101;
														assign node12610 = (inp[3]) ? node12616 : node12611;
															assign node12611 = (inp[15]) ? node12613 : 4'b0101;
																assign node12613 = (inp[0]) ? 4'b0111 : 4'b0101;
															assign node12616 = (inp[15]) ? node12620 : node12617;
																assign node12617 = (inp[0]) ? 4'b0101 : 4'b0111;
																assign node12620 = (inp[0]) ? 4'b0111 : 4'b0101;
													assign node12623 = (inp[15]) ? 4'b0101 : node12624;
														assign node12624 = (inp[10]) ? node12626 : 4'b0101;
															assign node12626 = (inp[3]) ? node12630 : node12627;
																assign node12627 = (inp[0]) ? 4'b0101 : 4'b0111;
																assign node12630 = (inp[0]) ? 4'b0111 : 4'b0101;
											assign node12634 = (inp[7]) ? node12656 : node12635;
												assign node12635 = (inp[15]) ? node12645 : node12636;
													assign node12636 = (inp[0]) ? node12640 : node12637;
														assign node12637 = (inp[3]) ? 4'b0101 : 4'b0111;
														assign node12640 = (inp[3]) ? node12642 : 4'b0101;
															assign node12642 = (inp[5]) ? 4'b0111 : 4'b0101;
													assign node12645 = (inp[0]) ? node12651 : node12646;
														assign node12646 = (inp[5]) ? node12648 : 4'b0101;
															assign node12648 = (inp[3]) ? 4'b0111 : 4'b0101;
														assign node12651 = (inp[5]) ? node12653 : 4'b0111;
															assign node12653 = (inp[3]) ? 4'b0101 : 4'b0111;
												assign node12656 = (inp[15]) ? node12664 : node12657;
													assign node12657 = (inp[0]) ? node12659 : 4'b0110;
														assign node12659 = (inp[3]) ? node12661 : 4'b0100;
															assign node12661 = (inp[5]) ? 4'b0110 : 4'b0100;
													assign node12664 = (inp[0]) ? node12670 : node12665;
														assign node12665 = (inp[3]) ? node12667 : 4'b0100;
															assign node12667 = (inp[5]) ? 4'b0110 : 4'b0100;
														assign node12670 = (inp[5]) ? node12672 : 4'b0110;
															assign node12672 = (inp[10]) ? 4'b0100 : 4'b0110;
									assign node12675 = (inp[15]) ? node12747 : node12676;
										assign node12676 = (inp[0]) ? node12716 : node12677;
											assign node12677 = (inp[5]) ? node12685 : node12678;
												assign node12678 = (inp[7]) ? node12682 : node12679;
													assign node12679 = (inp[8]) ? 4'b0111 : 4'b0110;
													assign node12682 = (inp[8]) ? 4'b0110 : 4'b0111;
												assign node12685 = (inp[3]) ? node12693 : node12686;
													assign node12686 = (inp[8]) ? node12690 : node12687;
														assign node12687 = (inp[7]) ? 4'b0111 : 4'b0110;
														assign node12690 = (inp[7]) ? 4'b0110 : 4'b0111;
													assign node12693 = (inp[2]) ? node12705 : node12694;
														assign node12694 = (inp[10]) ? node12700 : node12695;
															assign node12695 = (inp[7]) ? 4'b0100 : node12696;
																assign node12696 = (inp[8]) ? 4'b0101 : 4'b0100;
															assign node12700 = (inp[7]) ? node12702 : 4'b0100;
																assign node12702 = (inp[8]) ? 4'b0100 : 4'b0101;
														assign node12705 = (inp[10]) ? node12711 : node12706;
															assign node12706 = (inp[8]) ? node12708 : 4'b0101;
																assign node12708 = (inp[7]) ? 4'b0100 : 4'b0101;
															assign node12711 = (inp[7]) ? 4'b0100 : node12712;
																assign node12712 = (inp[8]) ? 4'b0101 : 4'b0100;
											assign node12716 = (inp[3]) ? node12732 : node12717;
												assign node12717 = (inp[2]) ? node12725 : node12718;
													assign node12718 = (inp[7]) ? node12722 : node12719;
														assign node12719 = (inp[8]) ? 4'b0101 : 4'b0100;
														assign node12722 = (inp[8]) ? 4'b0100 : 4'b0101;
													assign node12725 = (inp[7]) ? node12729 : node12726;
														assign node12726 = (inp[8]) ? 4'b0101 : 4'b0100;
														assign node12729 = (inp[8]) ? 4'b0100 : 4'b0101;
												assign node12732 = (inp[5]) ? node12740 : node12733;
													assign node12733 = (inp[7]) ? node12737 : node12734;
														assign node12734 = (inp[8]) ? 4'b0101 : 4'b0100;
														assign node12737 = (inp[8]) ? 4'b0100 : 4'b0101;
													assign node12740 = (inp[8]) ? node12744 : node12741;
														assign node12741 = (inp[7]) ? 4'b0111 : 4'b0110;
														assign node12744 = (inp[7]) ? 4'b0110 : 4'b0111;
										assign node12747 = (inp[0]) ? node12799 : node12748;
											assign node12748 = (inp[5]) ? node12784 : node12749;
												assign node12749 = (inp[2]) ? node12767 : node12750;
													assign node12750 = (inp[3]) ? node12760 : node12751;
														assign node12751 = (inp[10]) ? node12755 : node12752;
															assign node12752 = (inp[8]) ? 4'b0100 : 4'b0101;
															assign node12755 = (inp[7]) ? 4'b0100 : node12756;
																assign node12756 = (inp[8]) ? 4'b0101 : 4'b0100;
														assign node12760 = (inp[8]) ? node12764 : node12761;
															assign node12761 = (inp[7]) ? 4'b0101 : 4'b0100;
															assign node12764 = (inp[7]) ? 4'b0100 : 4'b0101;
													assign node12767 = (inp[10]) ? node12777 : node12768;
														assign node12768 = (inp[3]) ? node12770 : 4'b0101;
															assign node12770 = (inp[8]) ? node12774 : node12771;
																assign node12771 = (inp[7]) ? 4'b0101 : 4'b0100;
																assign node12774 = (inp[7]) ? 4'b0100 : 4'b0101;
														assign node12777 = (inp[8]) ? node12781 : node12778;
															assign node12778 = (inp[7]) ? 4'b0101 : 4'b0100;
															assign node12781 = (inp[7]) ? 4'b0100 : 4'b0101;
												assign node12784 = (inp[3]) ? node12792 : node12785;
													assign node12785 = (inp[8]) ? node12789 : node12786;
														assign node12786 = (inp[7]) ? 4'b0101 : 4'b0100;
														assign node12789 = (inp[7]) ? 4'b0100 : 4'b0101;
													assign node12792 = (inp[8]) ? node12796 : node12793;
														assign node12793 = (inp[7]) ? 4'b0111 : 4'b0110;
														assign node12796 = (inp[7]) ? 4'b0110 : 4'b0111;
											assign node12799 = (inp[5]) ? node12807 : node12800;
												assign node12800 = (inp[7]) ? node12804 : node12801;
													assign node12801 = (inp[8]) ? 4'b0111 : 4'b0110;
													assign node12804 = (inp[8]) ? 4'b0110 : 4'b0111;
												assign node12807 = (inp[3]) ? node12823 : node12808;
													assign node12808 = (inp[10]) ? node12818 : node12809;
														assign node12809 = (inp[2]) ? 4'b0110 : node12810;
															assign node12810 = (inp[8]) ? node12814 : node12811;
																assign node12811 = (inp[7]) ? 4'b0111 : 4'b0110;
																assign node12814 = (inp[7]) ? 4'b0110 : 4'b0111;
														assign node12818 = (inp[8]) ? node12820 : 4'b0111;
															assign node12820 = (inp[7]) ? 4'b0110 : 4'b0111;
													assign node12823 = (inp[10]) ? node12831 : node12824;
														assign node12824 = (inp[7]) ? node12828 : node12825;
															assign node12825 = (inp[8]) ? 4'b0101 : 4'b0100;
															assign node12828 = (inp[8]) ? 4'b0100 : 4'b0101;
														assign node12831 = (inp[2]) ? 4'b0101 : node12832;
															assign node12832 = (inp[7]) ? node12834 : 4'b0101;
																assign node12834 = (inp[8]) ? 4'b0100 : 4'b0101;
								assign node12838 = (inp[10]) ? node13092 : node12839;
									assign node12839 = (inp[2]) ? node12981 : node12840;
										assign node12840 = (inp[5]) ? node12906 : node12841;
											assign node12841 = (inp[8]) ? node12877 : node12842;
												assign node12842 = (inp[15]) ? node12858 : node12843;
													assign node12843 = (inp[0]) ? node12851 : node12844;
														assign node12844 = (inp[7]) ? node12848 : node12845;
															assign node12845 = (inp[14]) ? 4'b0110 : 4'b0111;
															assign node12848 = (inp[14]) ? 4'b0111 : 4'b0110;
														assign node12851 = (inp[7]) ? node12855 : node12852;
															assign node12852 = (inp[14]) ? 4'b0100 : 4'b0101;
															assign node12855 = (inp[14]) ? 4'b0101 : 4'b0100;
													assign node12858 = (inp[0]) ? node12870 : node12859;
														assign node12859 = (inp[3]) ? node12865 : node12860;
															assign node12860 = (inp[7]) ? 4'b0101 : node12861;
																assign node12861 = (inp[14]) ? 4'b0100 : 4'b0101;
															assign node12865 = (inp[14]) ? 4'b0101 : node12866;
																assign node12866 = (inp[7]) ? 4'b0100 : 4'b0101;
														assign node12870 = (inp[14]) ? node12874 : node12871;
															assign node12871 = (inp[7]) ? 4'b0110 : 4'b0111;
															assign node12874 = (inp[7]) ? 4'b0111 : 4'b0110;
												assign node12877 = (inp[15]) ? node12891 : node12878;
													assign node12878 = (inp[0]) ? node12884 : node12879;
														assign node12879 = (inp[7]) ? node12881 : 4'b0110;
															assign node12881 = (inp[14]) ? 4'b0110 : 4'b0111;
														assign node12884 = (inp[14]) ? node12888 : node12885;
															assign node12885 = (inp[7]) ? 4'b0101 : 4'b0100;
															assign node12888 = (inp[7]) ? 4'b0100 : 4'b0101;
													assign node12891 = (inp[0]) ? node12899 : node12892;
														assign node12892 = (inp[14]) ? node12896 : node12893;
															assign node12893 = (inp[7]) ? 4'b0101 : 4'b0100;
															assign node12896 = (inp[7]) ? 4'b0100 : 4'b0101;
														assign node12899 = (inp[7]) ? node12903 : node12900;
															assign node12900 = (inp[14]) ? 4'b0111 : 4'b0110;
															assign node12903 = (inp[14]) ? 4'b0110 : 4'b0111;
											assign node12906 = (inp[8]) ? node12940 : node12907;
												assign node12907 = (inp[3]) ? node12923 : node12908;
													assign node12908 = (inp[14]) ? node12920 : node12909;
														assign node12909 = (inp[7]) ? node12917 : node12910;
															assign node12910 = (inp[15]) ? node12914 : node12911;
																assign node12911 = (inp[0]) ? 4'b0101 : 4'b0111;
																assign node12914 = (inp[0]) ? 4'b0111 : 4'b0101;
															assign node12917 = (inp[0]) ? 4'b0110 : 4'b0100;
														assign node12920 = (inp[7]) ? 4'b0101 : 4'b0100;
													assign node12923 = (inp[14]) ? node12933 : node12924;
														assign node12924 = (inp[7]) ? node12926 : 4'b0101;
															assign node12926 = (inp[0]) ? node12930 : node12927;
																assign node12927 = (inp[15]) ? 4'b0110 : 4'b0100;
																assign node12930 = (inp[15]) ? 4'b0100 : 4'b0110;
														assign node12933 = (inp[7]) ? node12935 : 4'b0110;
															assign node12935 = (inp[15]) ? node12937 : 4'b0111;
																assign node12937 = (inp[0]) ? 4'b0101 : 4'b0111;
												assign node12940 = (inp[0]) ? node12960 : node12941;
													assign node12941 = (inp[14]) ? node12951 : node12942;
														assign node12942 = (inp[7]) ? node12944 : 4'b0110;
															assign node12944 = (inp[15]) ? node12948 : node12945;
																assign node12945 = (inp[3]) ? 4'b0101 : 4'b0111;
																assign node12948 = (inp[3]) ? 4'b0111 : 4'b0101;
														assign node12951 = (inp[7]) ? 4'b0110 : node12952;
															assign node12952 = (inp[3]) ? node12956 : node12953;
																assign node12953 = (inp[15]) ? 4'b0101 : 4'b0111;
																assign node12956 = (inp[15]) ? 4'b0111 : 4'b0101;
													assign node12960 = (inp[14]) ? node12974 : node12961;
														assign node12961 = (inp[7]) ? node12967 : node12962;
															assign node12962 = (inp[3]) ? node12964 : 4'b0110;
																assign node12964 = (inp[15]) ? 4'b0100 : 4'b0110;
															assign node12967 = (inp[3]) ? node12971 : node12968;
																assign node12968 = (inp[15]) ? 4'b0111 : 4'b0101;
																assign node12971 = (inp[15]) ? 4'b0101 : 4'b0111;
														assign node12974 = (inp[7]) ? 4'b0100 : node12975;
															assign node12975 = (inp[15]) ? 4'b0101 : node12976;
																assign node12976 = (inp[3]) ? 4'b0111 : 4'b0101;
										assign node12981 = (inp[7]) ? node13037 : node12982;
											assign node12982 = (inp[8]) ? node13004 : node12983;
												assign node12983 = (inp[0]) ? node12993 : node12984;
													assign node12984 = (inp[15]) ? node12988 : node12985;
														assign node12985 = (inp[5]) ? 4'b0100 : 4'b0110;
														assign node12988 = (inp[5]) ? node12990 : 4'b0100;
															assign node12990 = (inp[3]) ? 4'b0110 : 4'b0100;
													assign node12993 = (inp[15]) ? node12999 : node12994;
														assign node12994 = (inp[3]) ? node12996 : 4'b0100;
															assign node12996 = (inp[5]) ? 4'b0110 : 4'b0100;
														assign node12999 = (inp[3]) ? node13001 : 4'b0110;
															assign node13001 = (inp[14]) ? 4'b0100 : 4'b0110;
												assign node13004 = (inp[3]) ? node13018 : node13005;
													assign node13005 = (inp[14]) ? node13013 : node13006;
														assign node13006 = (inp[0]) ? node13010 : node13007;
															assign node13007 = (inp[15]) ? 4'b0101 : 4'b0111;
															assign node13010 = (inp[15]) ? 4'b0111 : 4'b0101;
														assign node13013 = (inp[0]) ? node13015 : 4'b0101;
															assign node13015 = (inp[15]) ? 4'b0111 : 4'b0101;
													assign node13018 = (inp[14]) ? node13032 : node13019;
														assign node13019 = (inp[5]) ? node13027 : node13020;
															assign node13020 = (inp[0]) ? node13024 : node13021;
																assign node13021 = (inp[15]) ? 4'b0101 : 4'b0111;
																assign node13024 = (inp[15]) ? 4'b0111 : 4'b0101;
															assign node13027 = (inp[15]) ? node13029 : 4'b0101;
																assign node13029 = (inp[0]) ? 4'b0101 : 4'b0111;
														assign node13032 = (inp[0]) ? 4'b0111 : node13033;
															assign node13033 = (inp[5]) ? 4'b0101 : 4'b0111;
											assign node13037 = (inp[8]) ? node13055 : node13038;
												assign node13038 = (inp[0]) ? node13044 : node13039;
													assign node13039 = (inp[15]) ? node13041 : 4'b0111;
														assign node13041 = (inp[5]) ? 4'b0111 : 4'b0101;
													assign node13044 = (inp[15]) ? node13050 : node13045;
														assign node13045 = (inp[5]) ? node13047 : 4'b0101;
															assign node13047 = (inp[3]) ? 4'b0111 : 4'b0101;
														assign node13050 = (inp[3]) ? node13052 : 4'b0111;
															assign node13052 = (inp[5]) ? 4'b0101 : 4'b0111;
												assign node13055 = (inp[14]) ? node13075 : node13056;
													assign node13056 = (inp[3]) ? node13062 : node13057;
														assign node13057 = (inp[0]) ? node13059 : 4'b0100;
															assign node13059 = (inp[15]) ? 4'b0110 : 4'b0100;
														assign node13062 = (inp[0]) ? node13070 : node13063;
															assign node13063 = (inp[15]) ? node13067 : node13064;
																assign node13064 = (inp[5]) ? 4'b0100 : 4'b0110;
																assign node13067 = (inp[5]) ? 4'b0110 : 4'b0100;
															assign node13070 = (inp[5]) ? node13072 : 4'b0100;
																assign node13072 = (inp[15]) ? 4'b0100 : 4'b0110;
													assign node13075 = (inp[5]) ? node13083 : node13076;
														assign node13076 = (inp[15]) ? node13080 : node13077;
															assign node13077 = (inp[0]) ? 4'b0100 : 4'b0110;
															assign node13080 = (inp[0]) ? 4'b0110 : 4'b0100;
														assign node13083 = (inp[0]) ? 4'b0100 : node13084;
															assign node13084 = (inp[15]) ? node13088 : node13085;
																assign node13085 = (inp[3]) ? 4'b0100 : 4'b0110;
																assign node13088 = (inp[3]) ? 4'b0110 : 4'b0100;
									assign node13092 = (inp[5]) ? node13254 : node13093;
										assign node13093 = (inp[3]) ? node13171 : node13094;
											assign node13094 = (inp[8]) ? node13128 : node13095;
												assign node13095 = (inp[7]) ? node13111 : node13096;
													assign node13096 = (inp[14]) ? node13106 : node13097;
														assign node13097 = (inp[2]) ? 4'b0000 : node13098;
															assign node13098 = (inp[15]) ? node13102 : node13099;
																assign node13099 = (inp[0]) ? 4'b0001 : 4'b0011;
																assign node13102 = (inp[0]) ? 4'b0011 : 4'b0001;
														assign node13106 = (inp[15]) ? node13108 : 4'b0000;
															assign node13108 = (inp[0]) ? 4'b0010 : 4'b0000;
													assign node13111 = (inp[14]) ? node13121 : node13112;
														assign node13112 = (inp[2]) ? node13114 : 4'b0010;
															assign node13114 = (inp[0]) ? node13118 : node13115;
																assign node13115 = (inp[15]) ? 4'b0001 : 4'b0011;
																assign node13118 = (inp[15]) ? 4'b0011 : 4'b0001;
														assign node13121 = (inp[15]) ? node13125 : node13122;
															assign node13122 = (inp[0]) ? 4'b0001 : 4'b0011;
															assign node13125 = (inp[0]) ? 4'b0011 : 4'b0001;
												assign node13128 = (inp[7]) ? node13148 : node13129;
													assign node13129 = (inp[2]) ? node13141 : node13130;
														assign node13130 = (inp[14]) ? node13134 : node13131;
															assign node13131 = (inp[15]) ? 4'b0010 : 4'b0000;
															assign node13134 = (inp[15]) ? node13138 : node13135;
																assign node13135 = (inp[0]) ? 4'b0001 : 4'b0011;
																assign node13138 = (inp[0]) ? 4'b0011 : 4'b0001;
														assign node13141 = (inp[15]) ? node13145 : node13142;
															assign node13142 = (inp[0]) ? 4'b0001 : 4'b0011;
															assign node13145 = (inp[0]) ? 4'b0011 : 4'b0001;
													assign node13148 = (inp[2]) ? node13158 : node13149;
														assign node13149 = (inp[14]) ? node13151 : 4'b0001;
															assign node13151 = (inp[0]) ? node13155 : node13152;
																assign node13152 = (inp[15]) ? 4'b0000 : 4'b0010;
																assign node13155 = (inp[15]) ? 4'b0010 : 4'b0000;
														assign node13158 = (inp[14]) ? node13164 : node13159;
															assign node13159 = (inp[15]) ? node13161 : 4'b0010;
																assign node13161 = (inp[0]) ? 4'b0010 : 4'b0000;
															assign node13164 = (inp[0]) ? node13168 : node13165;
																assign node13165 = (inp[15]) ? 4'b0000 : 4'b0010;
																assign node13168 = (inp[15]) ? 4'b0010 : 4'b0000;
											assign node13171 = (inp[14]) ? node13223 : node13172;
												assign node13172 = (inp[8]) ? node13200 : node13173;
													assign node13173 = (inp[15]) ? node13187 : node13174;
														assign node13174 = (inp[0]) ? node13182 : node13175;
															assign node13175 = (inp[7]) ? node13179 : node13176;
																assign node13176 = (inp[2]) ? 4'b0010 : 4'b0011;
																assign node13179 = (inp[2]) ? 4'b0011 : 4'b0010;
															assign node13182 = (inp[7]) ? 4'b0000 : node13183;
																assign node13183 = (inp[2]) ? 4'b0000 : 4'b0001;
														assign node13187 = (inp[0]) ? node13195 : node13188;
															assign node13188 = (inp[2]) ? node13192 : node13189;
																assign node13189 = (inp[7]) ? 4'b0000 : 4'b0001;
																assign node13192 = (inp[7]) ? 4'b0001 : 4'b0000;
															assign node13195 = (inp[2]) ? node13197 : 4'b0011;
																assign node13197 = (inp[7]) ? 4'b0011 : 4'b0010;
													assign node13200 = (inp[15]) ? node13210 : node13201;
														assign node13201 = (inp[0]) ? node13205 : node13202;
															assign node13202 = (inp[2]) ? 4'b0011 : 4'b0010;
															assign node13205 = (inp[2]) ? node13207 : 4'b0001;
																assign node13207 = (inp[7]) ? 4'b0000 : 4'b0001;
														assign node13210 = (inp[0]) ? node13218 : node13211;
															assign node13211 = (inp[7]) ? node13215 : node13212;
																assign node13212 = (inp[2]) ? 4'b0001 : 4'b0000;
																assign node13215 = (inp[2]) ? 4'b0000 : 4'b0001;
															assign node13218 = (inp[7]) ? node13220 : 4'b0010;
																assign node13220 = (inp[2]) ? 4'b0010 : 4'b0011;
												assign node13223 = (inp[8]) ? node13239 : node13224;
													assign node13224 = (inp[7]) ? node13232 : node13225;
														assign node13225 = (inp[0]) ? node13229 : node13226;
															assign node13226 = (inp[15]) ? 4'b0000 : 4'b0010;
															assign node13229 = (inp[15]) ? 4'b0010 : 4'b0000;
														assign node13232 = (inp[0]) ? node13236 : node13233;
															assign node13233 = (inp[15]) ? 4'b0001 : 4'b0011;
															assign node13236 = (inp[15]) ? 4'b0011 : 4'b0001;
													assign node13239 = (inp[7]) ? node13245 : node13240;
														assign node13240 = (inp[15]) ? 4'b0011 : node13241;
															assign node13241 = (inp[0]) ? 4'b0001 : 4'b0011;
														assign node13245 = (inp[2]) ? node13251 : node13246;
															assign node13246 = (inp[15]) ? node13248 : 4'b0010;
																assign node13248 = (inp[0]) ? 4'b0010 : 4'b0000;
															assign node13251 = (inp[0]) ? 4'b0000 : 4'b0010;
										assign node13254 = (inp[7]) ? node13330 : node13255;
											assign node13255 = (inp[8]) ? node13289 : node13256;
												assign node13256 = (inp[2]) ? node13272 : node13257;
													assign node13257 = (inp[14]) ? node13265 : node13258;
														assign node13258 = (inp[15]) ? 4'b0011 : node13259;
															assign node13259 = (inp[3]) ? 4'b0011 : node13260;
																assign node13260 = (inp[0]) ? 4'b0001 : 4'b0011;
														assign node13265 = (inp[0]) ? node13267 : 4'b0000;
															assign node13267 = (inp[15]) ? 4'b0010 : node13268;
																assign node13268 = (inp[3]) ? 4'b0010 : 4'b0000;
													assign node13272 = (inp[3]) ? node13282 : node13273;
														assign node13273 = (inp[14]) ? node13277 : node13274;
															assign node13274 = (inp[15]) ? 4'b0000 : 4'b0010;
															assign node13277 = (inp[0]) ? node13279 : 4'b0010;
																assign node13279 = (inp[15]) ? 4'b0010 : 4'b0000;
														assign node13282 = (inp[15]) ? node13286 : node13283;
															assign node13283 = (inp[0]) ? 4'b0010 : 4'b0000;
															assign node13286 = (inp[0]) ? 4'b0000 : 4'b0010;
												assign node13289 = (inp[14]) ? node13311 : node13290;
													assign node13290 = (inp[2]) ? node13306 : node13291;
														assign node13291 = (inp[15]) ? node13299 : node13292;
															assign node13292 = (inp[3]) ? node13296 : node13293;
																assign node13293 = (inp[0]) ? 4'b0000 : 4'b0010;
																assign node13296 = (inp[0]) ? 4'b0010 : 4'b0000;
															assign node13299 = (inp[0]) ? node13303 : node13300;
																assign node13300 = (inp[3]) ? 4'b0010 : 4'b0000;
																assign node13303 = (inp[3]) ? 4'b0000 : 4'b0010;
														assign node13306 = (inp[0]) ? 4'b0011 : node13307;
															assign node13307 = (inp[15]) ? 4'b0001 : 4'b0011;
													assign node13311 = (inp[2]) ? node13321 : node13312;
														assign node13312 = (inp[0]) ? 4'b0011 : node13313;
															assign node13313 = (inp[15]) ? node13317 : node13314;
																assign node13314 = (inp[3]) ? 4'b0001 : 4'b0011;
																assign node13317 = (inp[3]) ? 4'b0011 : 4'b0001;
														assign node13321 = (inp[0]) ? 4'b0001 : node13322;
															assign node13322 = (inp[3]) ? node13326 : node13323;
																assign node13323 = (inp[15]) ? 4'b0001 : 4'b0011;
																assign node13326 = (inp[15]) ? 4'b0011 : 4'b0001;
											assign node13330 = (inp[8]) ? node13358 : node13331;
												assign node13331 = (inp[2]) ? node13349 : node13332;
													assign node13332 = (inp[14]) ? node13342 : node13333;
														assign node13333 = (inp[15]) ? 4'b0000 : node13334;
															assign node13334 = (inp[3]) ? node13338 : node13335;
																assign node13335 = (inp[0]) ? 4'b0000 : 4'b0010;
																assign node13338 = (inp[0]) ? 4'b0010 : 4'b0000;
														assign node13342 = (inp[15]) ? 4'b0011 : node13343;
															assign node13343 = (inp[0]) ? node13345 : 4'b0001;
																assign node13345 = (inp[3]) ? 4'b0011 : 4'b0001;
													assign node13349 = (inp[15]) ? 4'b0001 : node13350;
														assign node13350 = (inp[3]) ? node13354 : node13351;
															assign node13351 = (inp[0]) ? 4'b0001 : 4'b0011;
															assign node13354 = (inp[0]) ? 4'b0011 : 4'b0001;
												assign node13358 = (inp[2]) ? node13382 : node13359;
													assign node13359 = (inp[14]) ? node13371 : node13360;
														assign node13360 = (inp[15]) ? node13366 : node13361;
															assign node13361 = (inp[3]) ? node13363 : 4'b0001;
																assign node13363 = (inp[0]) ? 4'b0011 : 4'b0001;
															assign node13366 = (inp[0]) ? node13368 : 4'b0011;
																assign node13368 = (inp[3]) ? 4'b0001 : 4'b0011;
														assign node13371 = (inp[0]) ? node13377 : node13372;
															assign node13372 = (inp[3]) ? node13374 : 4'b0000;
																assign node13374 = (inp[15]) ? 4'b0010 : 4'b0000;
															assign node13377 = (inp[3]) ? node13379 : 4'b0010;
																assign node13379 = (inp[15]) ? 4'b0000 : 4'b0010;
													assign node13382 = (inp[0]) ? node13390 : node13383;
														assign node13383 = (inp[15]) ? node13387 : node13384;
															assign node13384 = (inp[3]) ? 4'b0000 : 4'b0010;
															assign node13387 = (inp[3]) ? 4'b0010 : 4'b0000;
														assign node13390 = (inp[3]) ? node13394 : node13391;
															assign node13391 = (inp[15]) ? 4'b0010 : 4'b0000;
															assign node13394 = (inp[15]) ? 4'b0000 : 4'b0010;
							assign node13397 = (inp[10]) ? node13897 : node13398;
								assign node13398 = (inp[2]) ? node13668 : node13399;
									assign node13399 = (inp[3]) ? node13515 : node13400;
										assign node13400 = (inp[15]) ? node13468 : node13401;
											assign node13401 = (inp[0]) ? node13429 : node13402;
												assign node13402 = (inp[12]) ? node13416 : node13403;
													assign node13403 = (inp[14]) ? node13411 : node13404;
														assign node13404 = (inp[7]) ? node13408 : node13405;
															assign node13405 = (inp[8]) ? 4'b0010 : 4'b0011;
															assign node13408 = (inp[8]) ? 4'b0011 : 4'b0010;
														assign node13411 = (inp[8]) ? node13413 : 4'b0010;
															assign node13413 = (inp[7]) ? 4'b0010 : 4'b0011;
													assign node13416 = (inp[8]) ? node13422 : node13417;
														assign node13417 = (inp[7]) ? node13419 : 4'b0011;
															assign node13419 = (inp[14]) ? 4'b0011 : 4'b0010;
														assign node13422 = (inp[7]) ? node13426 : node13423;
															assign node13423 = (inp[14]) ? 4'b0011 : 4'b0010;
															assign node13426 = (inp[14]) ? 4'b0010 : 4'b0011;
												assign node13429 = (inp[7]) ? node13451 : node13430;
													assign node13430 = (inp[5]) ? node13444 : node13431;
														assign node13431 = (inp[12]) ? node13439 : node13432;
															assign node13432 = (inp[8]) ? node13436 : node13433;
																assign node13433 = (inp[14]) ? 4'b0000 : 4'b0001;
																assign node13436 = (inp[14]) ? 4'b0001 : 4'b0000;
															assign node13439 = (inp[8]) ? 4'b0000 : node13440;
																assign node13440 = (inp[14]) ? 4'b0000 : 4'b0001;
														assign node13444 = (inp[12]) ? node13446 : 4'b0000;
															assign node13446 = (inp[14]) ? node13448 : 4'b0000;
																assign node13448 = (inp[8]) ? 4'b0001 : 4'b0000;
													assign node13451 = (inp[12]) ? node13459 : node13452;
														assign node13452 = (inp[14]) ? node13456 : node13453;
															assign node13453 = (inp[8]) ? 4'b0001 : 4'b0000;
															assign node13456 = (inp[8]) ? 4'b0000 : 4'b0001;
														assign node13459 = (inp[5]) ? 4'b0000 : node13460;
															assign node13460 = (inp[8]) ? node13464 : node13461;
																assign node13461 = (inp[14]) ? 4'b0001 : 4'b0000;
																assign node13464 = (inp[14]) ? 4'b0000 : 4'b0001;
											assign node13468 = (inp[0]) ? node13482 : node13469;
												assign node13469 = (inp[14]) ? node13475 : node13470;
													assign node13470 = (inp[7]) ? 4'b0000 : node13471;
														assign node13471 = (inp[8]) ? 4'b0000 : 4'b0001;
													assign node13475 = (inp[12]) ? 4'b0001 : node13476;
														assign node13476 = (inp[8]) ? node13478 : 4'b0000;
															assign node13478 = (inp[7]) ? 4'b0000 : 4'b0001;
												assign node13482 = (inp[5]) ? node13496 : node13483;
													assign node13483 = (inp[7]) ? node13491 : node13484;
														assign node13484 = (inp[14]) ? node13488 : node13485;
															assign node13485 = (inp[8]) ? 4'b0010 : 4'b0011;
															assign node13488 = (inp[8]) ? 4'b0011 : 4'b0010;
														assign node13491 = (inp[14]) ? 4'b0010 : node13492;
															assign node13492 = (inp[8]) ? 4'b0011 : 4'b0010;
													assign node13496 = (inp[8]) ? node13508 : node13497;
														assign node13497 = (inp[12]) ? node13503 : node13498;
															assign node13498 = (inp[14]) ? 4'b0011 : node13499;
																assign node13499 = (inp[7]) ? 4'b0010 : 4'b0011;
															assign node13503 = (inp[14]) ? node13505 : 4'b0010;
																assign node13505 = (inp[7]) ? 4'b0011 : 4'b0010;
														assign node13508 = (inp[14]) ? node13512 : node13509;
															assign node13509 = (inp[7]) ? 4'b0011 : 4'b0010;
															assign node13512 = (inp[7]) ? 4'b0010 : 4'b0011;
										assign node13515 = (inp[14]) ? node13601 : node13516;
											assign node13516 = (inp[0]) ? node13560 : node13517;
												assign node13517 = (inp[7]) ? node13539 : node13518;
													assign node13518 = (inp[8]) ? node13534 : node13519;
														assign node13519 = (inp[12]) ? node13527 : node13520;
															assign node13520 = (inp[5]) ? node13524 : node13521;
																assign node13521 = (inp[15]) ? 4'b0001 : 4'b0011;
																assign node13524 = (inp[15]) ? 4'b0011 : 4'b0001;
															assign node13527 = (inp[15]) ? node13531 : node13528;
																assign node13528 = (inp[5]) ? 4'b0001 : 4'b0011;
																assign node13531 = (inp[5]) ? 4'b0011 : 4'b0001;
														assign node13534 = (inp[12]) ? node13536 : 4'b0010;
															assign node13536 = (inp[15]) ? 4'b0010 : 4'b0000;
													assign node13539 = (inp[8]) ? node13553 : node13540;
														assign node13540 = (inp[12]) ? node13546 : node13541;
															assign node13541 = (inp[5]) ? 4'b0000 : node13542;
																assign node13542 = (inp[15]) ? 4'b0000 : 4'b0010;
															assign node13546 = (inp[15]) ? node13550 : node13547;
																assign node13547 = (inp[5]) ? 4'b0000 : 4'b0010;
																assign node13550 = (inp[5]) ? 4'b0010 : 4'b0000;
														assign node13553 = (inp[5]) ? node13557 : node13554;
															assign node13554 = (inp[15]) ? 4'b0001 : 4'b0011;
															assign node13557 = (inp[15]) ? 4'b0011 : 4'b0001;
												assign node13560 = (inp[5]) ? node13576 : node13561;
													assign node13561 = (inp[15]) ? node13569 : node13562;
														assign node13562 = (inp[8]) ? node13566 : node13563;
															assign node13563 = (inp[7]) ? 4'b0000 : 4'b0001;
															assign node13566 = (inp[7]) ? 4'b0001 : 4'b0000;
														assign node13569 = (inp[8]) ? node13573 : node13570;
															assign node13570 = (inp[12]) ? 4'b0011 : 4'b0010;
															assign node13573 = (inp[7]) ? 4'b0011 : 4'b0010;
													assign node13576 = (inp[15]) ? node13588 : node13577;
														assign node13577 = (inp[12]) ? node13583 : node13578;
															assign node13578 = (inp[8]) ? 4'b0011 : node13579;
																assign node13579 = (inp[7]) ? 4'b0010 : 4'b0011;
															assign node13583 = (inp[7]) ? 4'b0011 : node13584;
																assign node13584 = (inp[8]) ? 4'b0010 : 4'b0011;
														assign node13588 = (inp[12]) ? node13594 : node13589;
															assign node13589 = (inp[7]) ? 4'b0001 : node13590;
																assign node13590 = (inp[8]) ? 4'b0000 : 4'b0001;
															assign node13594 = (inp[7]) ? node13598 : node13595;
																assign node13595 = (inp[8]) ? 4'b0000 : 4'b0001;
																assign node13598 = (inp[8]) ? 4'b0001 : 4'b0000;
											assign node13601 = (inp[7]) ? node13637 : node13602;
												assign node13602 = (inp[8]) ? node13618 : node13603;
													assign node13603 = (inp[5]) ? node13611 : node13604;
														assign node13604 = (inp[15]) ? node13608 : node13605;
															assign node13605 = (inp[0]) ? 4'b0000 : 4'b0010;
															assign node13608 = (inp[0]) ? 4'b0010 : 4'b0000;
														assign node13611 = (inp[15]) ? node13615 : node13612;
															assign node13612 = (inp[0]) ? 4'b0010 : 4'b0000;
															assign node13615 = (inp[0]) ? 4'b0000 : 4'b0010;
													assign node13618 = (inp[12]) ? node13630 : node13619;
														assign node13619 = (inp[15]) ? node13625 : node13620;
															assign node13620 = (inp[5]) ? 4'b0011 : node13621;
																assign node13621 = (inp[0]) ? 4'b0001 : 4'b0011;
															assign node13625 = (inp[5]) ? node13627 : 4'b0001;
																assign node13627 = (inp[0]) ? 4'b0001 : 4'b0011;
														assign node13630 = (inp[0]) ? 4'b0011 : node13631;
															assign node13631 = (inp[15]) ? 4'b0011 : node13632;
																assign node13632 = (inp[5]) ? 4'b0001 : 4'b0011;
												assign node13637 = (inp[8]) ? node13653 : node13638;
													assign node13638 = (inp[0]) ? node13646 : node13639;
														assign node13639 = (inp[5]) ? node13643 : node13640;
															assign node13640 = (inp[15]) ? 4'b0001 : 4'b0011;
															assign node13643 = (inp[15]) ? 4'b0011 : 4'b0001;
														assign node13646 = (inp[5]) ? node13650 : node13647;
															assign node13647 = (inp[15]) ? 4'b0011 : 4'b0001;
															assign node13650 = (inp[15]) ? 4'b0001 : 4'b0011;
													assign node13653 = (inp[5]) ? node13661 : node13654;
														assign node13654 = (inp[0]) ? node13658 : node13655;
															assign node13655 = (inp[15]) ? 4'b0000 : 4'b0010;
															assign node13658 = (inp[15]) ? 4'b0010 : 4'b0000;
														assign node13661 = (inp[0]) ? node13665 : node13662;
															assign node13662 = (inp[15]) ? 4'b0010 : 4'b0000;
															assign node13665 = (inp[15]) ? 4'b0000 : 4'b0010;
									assign node13668 = (inp[15]) ? node13782 : node13669;
										assign node13669 = (inp[0]) ? node13747 : node13670;
											assign node13670 = (inp[5]) ? node13710 : node13671;
												assign node13671 = (inp[3]) ? node13685 : node13672;
													assign node13672 = (inp[14]) ? node13678 : node13673;
														assign node13673 = (inp[7]) ? 4'b0010 : node13674;
															assign node13674 = (inp[8]) ? 4'b0011 : 4'b0010;
														assign node13678 = (inp[7]) ? node13682 : node13679;
															assign node13679 = (inp[8]) ? 4'b0011 : 4'b0010;
															assign node13682 = (inp[8]) ? 4'b0010 : 4'b0011;
													assign node13685 = (inp[12]) ? node13701 : node13686;
														assign node13686 = (inp[14]) ? node13694 : node13687;
															assign node13687 = (inp[8]) ? node13691 : node13688;
																assign node13688 = (inp[7]) ? 4'b0011 : 4'b0010;
																assign node13691 = (inp[7]) ? 4'b0010 : 4'b0011;
															assign node13694 = (inp[8]) ? node13698 : node13695;
																assign node13695 = (inp[7]) ? 4'b0011 : 4'b0010;
																assign node13698 = (inp[7]) ? 4'b0010 : 4'b0011;
														assign node13701 = (inp[14]) ? node13703 : 4'b0011;
															assign node13703 = (inp[8]) ? node13707 : node13704;
																assign node13704 = (inp[7]) ? 4'b0011 : 4'b0010;
																assign node13707 = (inp[7]) ? 4'b0010 : 4'b0011;
												assign node13710 = (inp[3]) ? node13724 : node13711;
													assign node13711 = (inp[12]) ? node13717 : node13712;
														assign node13712 = (inp[8]) ? 4'b0010 : node13713;
															assign node13713 = (inp[7]) ? 4'b0011 : 4'b0010;
														assign node13717 = (inp[8]) ? node13721 : node13718;
															assign node13718 = (inp[7]) ? 4'b0011 : 4'b0010;
															assign node13721 = (inp[7]) ? 4'b0010 : 4'b0011;
													assign node13724 = (inp[14]) ? node13740 : node13725;
														assign node13725 = (inp[12]) ? node13733 : node13726;
															assign node13726 = (inp[7]) ? node13730 : node13727;
																assign node13727 = (inp[8]) ? 4'b0001 : 4'b0000;
																assign node13730 = (inp[8]) ? 4'b0000 : 4'b0001;
															assign node13733 = (inp[7]) ? node13737 : node13734;
																assign node13734 = (inp[8]) ? 4'b0001 : 4'b0000;
																assign node13737 = (inp[8]) ? 4'b0000 : 4'b0001;
														assign node13740 = (inp[8]) ? node13744 : node13741;
															assign node13741 = (inp[7]) ? 4'b0001 : 4'b0000;
															assign node13744 = (inp[7]) ? 4'b0000 : 4'b0001;
											assign node13747 = (inp[5]) ? node13755 : node13748;
												assign node13748 = (inp[7]) ? node13752 : node13749;
													assign node13749 = (inp[8]) ? 4'b0001 : 4'b0000;
													assign node13752 = (inp[8]) ? 4'b0000 : 4'b0001;
												assign node13755 = (inp[3]) ? node13775 : node13756;
													assign node13756 = (inp[14]) ? node13762 : node13757;
														assign node13757 = (inp[12]) ? 4'b0001 : node13758;
															assign node13758 = (inp[8]) ? 4'b0001 : 4'b0000;
														assign node13762 = (inp[12]) ? node13768 : node13763;
															assign node13763 = (inp[8]) ? node13765 : 4'b0001;
																assign node13765 = (inp[7]) ? 4'b0000 : 4'b0001;
															assign node13768 = (inp[8]) ? node13772 : node13769;
																assign node13769 = (inp[7]) ? 4'b0001 : 4'b0000;
																assign node13772 = (inp[7]) ? 4'b0000 : 4'b0001;
													assign node13775 = (inp[8]) ? node13779 : node13776;
														assign node13776 = (inp[7]) ? 4'b0011 : 4'b0010;
														assign node13779 = (inp[7]) ? 4'b0010 : 4'b0011;
										assign node13782 = (inp[0]) ? node13816 : node13783;
											assign node13783 = (inp[5]) ? node13791 : node13784;
												assign node13784 = (inp[7]) ? node13788 : node13785;
													assign node13785 = (inp[8]) ? 4'b0001 : 4'b0000;
													assign node13788 = (inp[8]) ? 4'b0000 : 4'b0001;
												assign node13791 = (inp[3]) ? node13807 : node13792;
													assign node13792 = (inp[12]) ? node13800 : node13793;
														assign node13793 = (inp[7]) ? node13797 : node13794;
															assign node13794 = (inp[8]) ? 4'b0001 : 4'b0000;
															assign node13797 = (inp[8]) ? 4'b0000 : 4'b0001;
														assign node13800 = (inp[14]) ? node13802 : 4'b0001;
															assign node13802 = (inp[8]) ? node13804 : 4'b0001;
																assign node13804 = (inp[7]) ? 4'b0000 : 4'b0001;
													assign node13807 = (inp[12]) ? node13809 : 4'b0011;
														assign node13809 = (inp[8]) ? node13813 : node13810;
															assign node13810 = (inp[7]) ? 4'b0011 : 4'b0010;
															assign node13813 = (inp[7]) ? 4'b0010 : 4'b0011;
											assign node13816 = (inp[3]) ? node13862 : node13817;
												assign node13817 = (inp[12]) ? node13839 : node13818;
													assign node13818 = (inp[14]) ? node13832 : node13819;
														assign node13819 = (inp[5]) ? node13825 : node13820;
															assign node13820 = (inp[7]) ? 4'b0011 : node13821;
																assign node13821 = (inp[8]) ? 4'b0011 : 4'b0010;
															assign node13825 = (inp[8]) ? node13829 : node13826;
																assign node13826 = (inp[7]) ? 4'b0011 : 4'b0010;
																assign node13829 = (inp[7]) ? 4'b0010 : 4'b0011;
														assign node13832 = (inp[8]) ? node13836 : node13833;
															assign node13833 = (inp[7]) ? 4'b0011 : 4'b0010;
															assign node13836 = (inp[7]) ? 4'b0010 : 4'b0011;
													assign node13839 = (inp[14]) ? node13855 : node13840;
														assign node13840 = (inp[5]) ? node13848 : node13841;
															assign node13841 = (inp[7]) ? node13845 : node13842;
																assign node13842 = (inp[8]) ? 4'b0011 : 4'b0010;
																assign node13845 = (inp[8]) ? 4'b0010 : 4'b0011;
															assign node13848 = (inp[7]) ? node13852 : node13849;
																assign node13849 = (inp[8]) ? 4'b0011 : 4'b0010;
																assign node13852 = (inp[8]) ? 4'b0010 : 4'b0011;
														assign node13855 = (inp[8]) ? node13859 : node13856;
															assign node13856 = (inp[7]) ? 4'b0011 : 4'b0010;
															assign node13859 = (inp[5]) ? 4'b0010 : 4'b0011;
												assign node13862 = (inp[5]) ? node13876 : node13863;
													assign node13863 = (inp[12]) ? node13869 : node13864;
														assign node13864 = (inp[8]) ? 4'b0011 : node13865;
															assign node13865 = (inp[7]) ? 4'b0011 : 4'b0010;
														assign node13869 = (inp[8]) ? node13873 : node13870;
															assign node13870 = (inp[7]) ? 4'b0011 : 4'b0010;
															assign node13873 = (inp[7]) ? 4'b0010 : 4'b0011;
													assign node13876 = (inp[14]) ? node13884 : node13877;
														assign node13877 = (inp[8]) ? node13881 : node13878;
															assign node13878 = (inp[7]) ? 4'b0001 : 4'b0000;
															assign node13881 = (inp[7]) ? 4'b0000 : 4'b0001;
														assign node13884 = (inp[12]) ? node13890 : node13885;
															assign node13885 = (inp[7]) ? 4'b0001 : node13886;
																assign node13886 = (inp[8]) ? 4'b0001 : 4'b0000;
															assign node13890 = (inp[8]) ? node13894 : node13891;
																assign node13891 = (inp[7]) ? 4'b0001 : 4'b0000;
																assign node13894 = (inp[7]) ? 4'b0000 : 4'b0001;
								assign node13897 = (inp[12]) ? node14215 : node13898;
									assign node13898 = (inp[14]) ? node14072 : node13899;
										assign node13899 = (inp[0]) ? node13981 : node13900;
											assign node13900 = (inp[15]) ? node13944 : node13901;
												assign node13901 = (inp[3]) ? node13923 : node13902;
													assign node13902 = (inp[7]) ? node13910 : node13903;
														assign node13903 = (inp[8]) ? node13907 : node13904;
															assign node13904 = (inp[2]) ? 4'b0010 : 4'b0011;
															assign node13907 = (inp[2]) ? 4'b0011 : 4'b0010;
														assign node13910 = (inp[5]) ? node13916 : node13911;
															assign node13911 = (inp[8]) ? node13913 : 4'b0010;
																assign node13913 = (inp[2]) ? 4'b0010 : 4'b0011;
															assign node13916 = (inp[8]) ? node13920 : node13917;
																assign node13917 = (inp[2]) ? 4'b0011 : 4'b0010;
																assign node13920 = (inp[2]) ? 4'b0010 : 4'b0011;
													assign node13923 = (inp[5]) ? node13929 : node13924;
														assign node13924 = (inp[7]) ? node13926 : 4'b0010;
															assign node13926 = (inp[2]) ? 4'b0011 : 4'b0010;
														assign node13929 = (inp[8]) ? node13937 : node13930;
															assign node13930 = (inp[2]) ? node13934 : node13931;
																assign node13931 = (inp[7]) ? 4'b0000 : 4'b0001;
																assign node13934 = (inp[7]) ? 4'b0001 : 4'b0000;
															assign node13937 = (inp[2]) ? node13941 : node13938;
																assign node13938 = (inp[7]) ? 4'b0001 : 4'b0000;
																assign node13941 = (inp[7]) ? 4'b0000 : 4'b0001;
												assign node13944 = (inp[5]) ? node13962 : node13945;
													assign node13945 = (inp[2]) ? node13955 : node13946;
														assign node13946 = (inp[3]) ? node13952 : node13947;
															assign node13947 = (inp[8]) ? node13949 : 4'b0000;
																assign node13949 = (inp[7]) ? 4'b0001 : 4'b0000;
															assign node13952 = (inp[8]) ? 4'b0000 : 4'b0001;
														assign node13955 = (inp[8]) ? node13959 : node13956;
															assign node13956 = (inp[7]) ? 4'b0001 : 4'b0000;
															assign node13959 = (inp[7]) ? 4'b0000 : 4'b0001;
													assign node13962 = (inp[3]) ? node13974 : node13963;
														assign node13963 = (inp[2]) ? node13969 : node13964;
															assign node13964 = (inp[7]) ? 4'b0000 : node13965;
																assign node13965 = (inp[8]) ? 4'b0000 : 4'b0001;
															assign node13969 = (inp[7]) ? node13971 : 4'b0001;
																assign node13971 = (inp[8]) ? 4'b0000 : 4'b0001;
														assign node13974 = (inp[7]) ? 4'b0011 : node13975;
															assign node13975 = (inp[8]) ? 4'b0011 : node13976;
																assign node13976 = (inp[2]) ? 4'b0010 : 4'b0011;
											assign node13981 = (inp[15]) ? node14033 : node13982;
												assign node13982 = (inp[5]) ? node14006 : node13983;
													assign node13983 = (inp[7]) ? node13999 : node13984;
														assign node13984 = (inp[3]) ? node13992 : node13985;
															assign node13985 = (inp[2]) ? node13989 : node13986;
																assign node13986 = (inp[8]) ? 4'b0000 : 4'b0001;
																assign node13989 = (inp[8]) ? 4'b0001 : 4'b0000;
															assign node13992 = (inp[2]) ? node13996 : node13993;
																assign node13993 = (inp[8]) ? 4'b0000 : 4'b0001;
																assign node13996 = (inp[8]) ? 4'b0001 : 4'b0000;
														assign node13999 = (inp[2]) ? node14003 : node14000;
															assign node14000 = (inp[8]) ? 4'b0001 : 4'b0000;
															assign node14003 = (inp[8]) ? 4'b0000 : 4'b0001;
													assign node14006 = (inp[3]) ? node14020 : node14007;
														assign node14007 = (inp[7]) ? node14015 : node14008;
															assign node14008 = (inp[2]) ? node14012 : node14009;
																assign node14009 = (inp[8]) ? 4'b0000 : 4'b0001;
																assign node14012 = (inp[8]) ? 4'b0001 : 4'b0000;
															assign node14015 = (inp[8]) ? 4'b0001 : node14016;
																assign node14016 = (inp[2]) ? 4'b0001 : 4'b0000;
														assign node14020 = (inp[2]) ? node14028 : node14021;
															assign node14021 = (inp[7]) ? node14025 : node14022;
																assign node14022 = (inp[8]) ? 4'b0010 : 4'b0011;
																assign node14025 = (inp[8]) ? 4'b0011 : 4'b0010;
															assign node14028 = (inp[7]) ? 4'b0011 : node14029;
																assign node14029 = (inp[8]) ? 4'b0011 : 4'b0010;
												assign node14033 = (inp[5]) ? node14053 : node14034;
													assign node14034 = (inp[2]) ? node14042 : node14035;
														assign node14035 = (inp[8]) ? node14039 : node14036;
															assign node14036 = (inp[7]) ? 4'b0010 : 4'b0011;
															assign node14039 = (inp[7]) ? 4'b0011 : 4'b0010;
														assign node14042 = (inp[3]) ? node14048 : node14043;
															assign node14043 = (inp[8]) ? 4'b0011 : node14044;
																assign node14044 = (inp[7]) ? 4'b0011 : 4'b0010;
															assign node14048 = (inp[7]) ? node14050 : 4'b0011;
																assign node14050 = (inp[8]) ? 4'b0010 : 4'b0011;
													assign node14053 = (inp[3]) ? node14059 : node14054;
														assign node14054 = (inp[2]) ? node14056 : 4'b0011;
															assign node14056 = (inp[7]) ? 4'b0010 : 4'b0011;
														assign node14059 = (inp[8]) ? node14065 : node14060;
															assign node14060 = (inp[2]) ? node14062 : 4'b0001;
																assign node14062 = (inp[7]) ? 4'b0001 : 4'b0000;
															assign node14065 = (inp[2]) ? node14069 : node14066;
																assign node14066 = (inp[7]) ? 4'b0001 : 4'b0000;
																assign node14069 = (inp[7]) ? 4'b0000 : 4'b0001;
										assign node14072 = (inp[3]) ? node14118 : node14073;
											assign node14073 = (inp[7]) ? node14089 : node14074;
												assign node14074 = (inp[8]) ? node14082 : node14075;
													assign node14075 = (inp[0]) ? node14079 : node14076;
														assign node14076 = (inp[15]) ? 4'b0000 : 4'b0010;
														assign node14079 = (inp[15]) ? 4'b0010 : 4'b0000;
													assign node14082 = (inp[15]) ? node14086 : node14083;
														assign node14083 = (inp[0]) ? 4'b0001 : 4'b0011;
														assign node14086 = (inp[0]) ? 4'b0011 : 4'b0001;
												assign node14089 = (inp[8]) ? node14111 : node14090;
													assign node14090 = (inp[5]) ? node14104 : node14091;
														assign node14091 = (inp[2]) ? node14099 : node14092;
															assign node14092 = (inp[15]) ? node14096 : node14093;
																assign node14093 = (inp[0]) ? 4'b0001 : 4'b0011;
																assign node14096 = (inp[0]) ? 4'b0011 : 4'b0001;
															assign node14099 = (inp[15]) ? node14101 : 4'b0011;
																assign node14101 = (inp[0]) ? 4'b0011 : 4'b0001;
														assign node14104 = (inp[15]) ? node14108 : node14105;
															assign node14105 = (inp[0]) ? 4'b0001 : 4'b0011;
															assign node14108 = (inp[0]) ? 4'b0011 : 4'b0001;
													assign node14111 = (inp[0]) ? node14115 : node14112;
														assign node14112 = (inp[15]) ? 4'b0000 : 4'b0010;
														assign node14115 = (inp[15]) ? 4'b0010 : 4'b0000;
											assign node14118 = (inp[2]) ? node14160 : node14119;
												assign node14119 = (inp[0]) ? node14139 : node14120;
													assign node14120 = (inp[8]) ? node14128 : node14121;
														assign node14121 = (inp[7]) ? 4'b0011 : node14122;
															assign node14122 = (inp[15]) ? node14124 : 4'b0010;
																assign node14124 = (inp[5]) ? 4'b0010 : 4'b0000;
														assign node14128 = (inp[7]) ? node14134 : node14129;
															assign node14129 = (inp[5]) ? 4'b0011 : node14130;
																assign node14130 = (inp[15]) ? 4'b0001 : 4'b0011;
															assign node14134 = (inp[15]) ? node14136 : 4'b0000;
																assign node14136 = (inp[5]) ? 4'b0010 : 4'b0000;
													assign node14139 = (inp[5]) ? node14149 : node14140;
														assign node14140 = (inp[15]) ? node14142 : 4'b0001;
															assign node14142 = (inp[7]) ? node14146 : node14143;
																assign node14143 = (inp[8]) ? 4'b0011 : 4'b0010;
																assign node14146 = (inp[8]) ? 4'b0010 : 4'b0011;
														assign node14149 = (inp[15]) ? node14153 : node14150;
															assign node14150 = (inp[8]) ? 4'b0010 : 4'b0011;
															assign node14153 = (inp[8]) ? node14157 : node14154;
																assign node14154 = (inp[7]) ? 4'b0001 : 4'b0000;
																assign node14157 = (inp[7]) ? 4'b0000 : 4'b0001;
												assign node14160 = (inp[8]) ? node14184 : node14161;
													assign node14161 = (inp[7]) ? node14175 : node14162;
														assign node14162 = (inp[5]) ? node14170 : node14163;
															assign node14163 = (inp[0]) ? node14167 : node14164;
																assign node14164 = (inp[15]) ? 4'b0000 : 4'b0010;
																assign node14167 = (inp[15]) ? 4'b0010 : 4'b0000;
															assign node14170 = (inp[0]) ? node14172 : 4'b0000;
																assign node14172 = (inp[15]) ? 4'b0000 : 4'b0010;
														assign node14175 = (inp[15]) ? node14177 : 4'b0001;
															assign node14177 = (inp[5]) ? node14181 : node14178;
																assign node14178 = (inp[0]) ? 4'b0011 : 4'b0001;
																assign node14181 = (inp[0]) ? 4'b0001 : 4'b0011;
													assign node14184 = (inp[7]) ? node14200 : node14185;
														assign node14185 = (inp[0]) ? node14193 : node14186;
															assign node14186 = (inp[5]) ? node14190 : node14187;
																assign node14187 = (inp[15]) ? 4'b0001 : 4'b0011;
																assign node14190 = (inp[15]) ? 4'b0011 : 4'b0001;
															assign node14193 = (inp[5]) ? node14197 : node14194;
																assign node14194 = (inp[15]) ? 4'b0011 : 4'b0001;
																assign node14197 = (inp[15]) ? 4'b0001 : 4'b0011;
														assign node14200 = (inp[5]) ? node14208 : node14201;
															assign node14201 = (inp[0]) ? node14205 : node14202;
																assign node14202 = (inp[15]) ? 4'b0000 : 4'b0010;
																assign node14205 = (inp[15]) ? 4'b0010 : 4'b0000;
															assign node14208 = (inp[0]) ? node14212 : node14209;
																assign node14209 = (inp[15]) ? 4'b0010 : 4'b0000;
																assign node14212 = (inp[15]) ? 4'b0000 : 4'b0010;
									assign node14215 = (inp[5]) ? node14387 : node14216;
										assign node14216 = (inp[14]) ? node14308 : node14217;
											assign node14217 = (inp[15]) ? node14263 : node14218;
												assign node14218 = (inp[8]) ? node14238 : node14219;
													assign node14219 = (inp[2]) ? node14229 : node14220;
														assign node14220 = (inp[7]) ? node14224 : node14221;
															assign node14221 = (inp[3]) ? 4'b0101 : 4'b0111;
															assign node14224 = (inp[3]) ? node14226 : 4'b0100;
																assign node14226 = (inp[0]) ? 4'b0110 : 4'b0100;
														assign node14229 = (inp[7]) ? node14235 : node14230;
															assign node14230 = (inp[0]) ? 4'b0100 : node14231;
																assign node14231 = (inp[3]) ? 4'b0100 : 4'b0110;
															assign node14235 = (inp[3]) ? 4'b0111 : 4'b0101;
													assign node14238 = (inp[3]) ? node14248 : node14239;
														assign node14239 = (inp[0]) ? 4'b0100 : node14240;
															assign node14240 = (inp[7]) ? node14244 : node14241;
																assign node14241 = (inp[2]) ? 4'b0111 : 4'b0110;
																assign node14244 = (inp[2]) ? 4'b0110 : 4'b0111;
														assign node14248 = (inp[0]) ? node14256 : node14249;
															assign node14249 = (inp[7]) ? node14253 : node14250;
																assign node14250 = (inp[2]) ? 4'b0101 : 4'b0100;
																assign node14253 = (inp[2]) ? 4'b0100 : 4'b0101;
															assign node14256 = (inp[7]) ? node14260 : node14257;
																assign node14257 = (inp[2]) ? 4'b0111 : 4'b0110;
																assign node14260 = (inp[2]) ? 4'b0110 : 4'b0111;
												assign node14263 = (inp[0]) ? node14281 : node14264;
													assign node14264 = (inp[3]) ? node14272 : node14265;
														assign node14265 = (inp[7]) ? node14267 : 4'b0101;
															assign node14267 = (inp[8]) ? node14269 : 4'b0101;
																assign node14269 = (inp[2]) ? 4'b0100 : 4'b0101;
														assign node14272 = (inp[8]) ? node14274 : 4'b0111;
															assign node14274 = (inp[7]) ? node14278 : node14275;
																assign node14275 = (inp[2]) ? 4'b0111 : 4'b0110;
																assign node14278 = (inp[2]) ? 4'b0110 : 4'b0111;
													assign node14281 = (inp[3]) ? node14297 : node14282;
														assign node14282 = (inp[7]) ? node14290 : node14283;
															assign node14283 = (inp[8]) ? node14287 : node14284;
																assign node14284 = (inp[2]) ? 4'b0110 : 4'b0111;
																assign node14287 = (inp[2]) ? 4'b0111 : 4'b0110;
															assign node14290 = (inp[2]) ? node14294 : node14291;
																assign node14291 = (inp[8]) ? 4'b0111 : 4'b0110;
																assign node14294 = (inp[8]) ? 4'b0110 : 4'b0111;
														assign node14297 = (inp[8]) ? node14303 : node14298;
															assign node14298 = (inp[7]) ? node14300 : 4'b0100;
																assign node14300 = (inp[2]) ? 4'b0101 : 4'b0100;
															assign node14303 = (inp[2]) ? node14305 : 4'b0101;
																assign node14305 = (inp[7]) ? 4'b0100 : 4'b0101;
											assign node14308 = (inp[7]) ? node14346 : node14309;
												assign node14309 = (inp[8]) ? node14319 : node14310;
													assign node14310 = (inp[0]) ? node14312 : 4'b0100;
														assign node14312 = (inp[3]) ? node14316 : node14313;
															assign node14313 = (inp[15]) ? 4'b0110 : 4'b0100;
															assign node14316 = (inp[15]) ? 4'b0100 : 4'b0110;
													assign node14319 = (inp[15]) ? node14333 : node14320;
														assign node14320 = (inp[2]) ? node14328 : node14321;
															assign node14321 = (inp[0]) ? node14325 : node14322;
																assign node14322 = (inp[3]) ? 4'b0101 : 4'b0111;
																assign node14325 = (inp[3]) ? 4'b0111 : 4'b0101;
															assign node14328 = (inp[3]) ? node14330 : 4'b0101;
																assign node14330 = (inp[0]) ? 4'b0111 : 4'b0101;
														assign node14333 = (inp[2]) ? node14339 : node14334;
															assign node14334 = (inp[0]) ? node14336 : 4'b0111;
																assign node14336 = (inp[3]) ? 4'b0101 : 4'b0111;
															assign node14339 = (inp[3]) ? node14343 : node14340;
																assign node14340 = (inp[0]) ? 4'b0111 : 4'b0101;
																assign node14343 = (inp[0]) ? 4'b0101 : 4'b0111;
												assign node14346 = (inp[8]) ? node14376 : node14347;
													assign node14347 = (inp[2]) ? node14363 : node14348;
														assign node14348 = (inp[3]) ? node14356 : node14349;
															assign node14349 = (inp[0]) ? node14353 : node14350;
																assign node14350 = (inp[15]) ? 4'b0101 : 4'b0111;
																assign node14353 = (inp[15]) ? 4'b0111 : 4'b0101;
															assign node14356 = (inp[15]) ? node14360 : node14357;
																assign node14357 = (inp[0]) ? 4'b0111 : 4'b0101;
																assign node14360 = (inp[0]) ? 4'b0101 : 4'b0111;
														assign node14363 = (inp[15]) ? node14369 : node14364;
															assign node14364 = (inp[3]) ? node14366 : 4'b0101;
																assign node14366 = (inp[0]) ? 4'b0111 : 4'b0101;
															assign node14369 = (inp[0]) ? node14373 : node14370;
																assign node14370 = (inp[3]) ? 4'b0111 : 4'b0101;
																assign node14373 = (inp[3]) ? 4'b0101 : 4'b0111;
													assign node14376 = (inp[15]) ? node14382 : node14377;
														assign node14377 = (inp[2]) ? node14379 : 4'b0110;
															assign node14379 = (inp[0]) ? 4'b0110 : 4'b0100;
														assign node14382 = (inp[2]) ? node14384 : 4'b0100;
															assign node14384 = (inp[3]) ? 4'b0110 : 4'b0100;
										assign node14387 = (inp[7]) ? node14437 : node14388;
											assign node14388 = (inp[8]) ? node14414 : node14389;
												assign node14389 = (inp[14]) ? node14399 : node14390;
													assign node14390 = (inp[2]) ? 4'b0110 : node14391;
														assign node14391 = (inp[15]) ? node14395 : node14392;
															assign node14392 = (inp[0]) ? 4'b0111 : 4'b0101;
															assign node14395 = (inp[0]) ? 4'b0101 : 4'b0111;
													assign node14399 = (inp[2]) ? node14407 : node14400;
														assign node14400 = (inp[15]) ? node14404 : node14401;
															assign node14401 = (inp[0]) ? 4'b0110 : 4'b0100;
															assign node14404 = (inp[0]) ? 4'b0100 : 4'b0110;
														assign node14407 = (inp[0]) ? node14411 : node14408;
															assign node14408 = (inp[15]) ? 4'b0110 : 4'b0100;
															assign node14411 = (inp[15]) ? 4'b0100 : 4'b0110;
												assign node14414 = (inp[2]) ? node14430 : node14415;
													assign node14415 = (inp[14]) ? node14421 : node14416;
														assign node14416 = (inp[15]) ? node14418 : 4'b0110;
															assign node14418 = (inp[0]) ? 4'b0100 : 4'b0110;
														assign node14421 = (inp[3]) ? node14423 : 4'b0111;
															assign node14423 = (inp[15]) ? node14427 : node14424;
																assign node14424 = (inp[0]) ? 4'b0111 : 4'b0101;
																assign node14427 = (inp[0]) ? 4'b0101 : 4'b0111;
													assign node14430 = (inp[0]) ? node14434 : node14431;
														assign node14431 = (inp[15]) ? 4'b0111 : 4'b0101;
														assign node14434 = (inp[15]) ? 4'b0101 : 4'b0111;
											assign node14437 = (inp[8]) ? node14463 : node14438;
												assign node14438 = (inp[14]) ? node14456 : node14439;
													assign node14439 = (inp[2]) ? node14451 : node14440;
														assign node14440 = (inp[3]) ? node14446 : node14441;
															assign node14441 = (inp[15]) ? node14443 : 4'b0100;
																assign node14443 = (inp[0]) ? 4'b0100 : 4'b0110;
															assign node14446 = (inp[15]) ? 4'b0110 : node14447;
																assign node14447 = (inp[0]) ? 4'b0110 : 4'b0100;
														assign node14451 = (inp[0]) ? 4'b0111 : node14452;
															assign node14452 = (inp[15]) ? 4'b0111 : 4'b0101;
													assign node14456 = (inp[15]) ? node14460 : node14457;
														assign node14457 = (inp[0]) ? 4'b0111 : 4'b0101;
														assign node14460 = (inp[0]) ? 4'b0101 : 4'b0111;
												assign node14463 = (inp[2]) ? node14481 : node14464;
													assign node14464 = (inp[14]) ? node14472 : node14465;
														assign node14465 = (inp[0]) ? node14469 : node14466;
															assign node14466 = (inp[15]) ? 4'b0111 : 4'b0101;
															assign node14469 = (inp[15]) ? 4'b0101 : 4'b0111;
														assign node14472 = (inp[3]) ? node14474 : 4'b0110;
															assign node14474 = (inp[15]) ? node14478 : node14475;
																assign node14475 = (inp[0]) ? 4'b0110 : 4'b0100;
																assign node14478 = (inp[0]) ? 4'b0100 : 4'b0110;
													assign node14481 = (inp[14]) ? node14489 : node14482;
														assign node14482 = (inp[0]) ? node14486 : node14483;
															assign node14483 = (inp[15]) ? 4'b0110 : 4'b0100;
															assign node14486 = (inp[15]) ? 4'b0100 : 4'b0110;
														assign node14489 = (inp[15]) ? node14493 : node14490;
															assign node14490 = (inp[0]) ? 4'b0110 : 4'b0100;
															assign node14493 = (inp[0]) ? 4'b0100 : 4'b0110;
						assign node14496 = (inp[4]) ? node15438 : node14497;
							assign node14497 = (inp[12]) ? node14963 : node14498;
								assign node14498 = (inp[14]) ? node14794 : node14499;
									assign node14499 = (inp[3]) ? node14663 : node14500;
										assign node14500 = (inp[10]) ? node14582 : node14501;
											assign node14501 = (inp[7]) ? node14543 : node14502;
												assign node14502 = (inp[5]) ? node14520 : node14503;
													assign node14503 = (inp[0]) ? node14511 : node14504;
														assign node14504 = (inp[15]) ? 4'b0000 : node14505;
															assign node14505 = (inp[2]) ? 4'b0010 : node14506;
																assign node14506 = (inp[8]) ? 4'b0010 : 4'b0011;
														assign node14511 = (inp[15]) ? node14513 : 4'b0001;
															assign node14513 = (inp[2]) ? node14517 : node14514;
																assign node14514 = (inp[8]) ? 4'b0010 : 4'b0011;
																assign node14517 = (inp[8]) ? 4'b0011 : 4'b0010;
													assign node14520 = (inp[0]) ? node14534 : node14521;
														assign node14521 = (inp[15]) ? node14529 : node14522;
															assign node14522 = (inp[2]) ? node14526 : node14523;
																assign node14523 = (inp[8]) ? 4'b0010 : 4'b0011;
																assign node14526 = (inp[8]) ? 4'b0011 : 4'b0010;
															assign node14529 = (inp[8]) ? node14531 : 4'b0001;
																assign node14531 = (inp[2]) ? 4'b0001 : 4'b0000;
														assign node14534 = (inp[15]) ? node14536 : 4'b0000;
															assign node14536 = (inp[2]) ? node14540 : node14537;
																assign node14537 = (inp[8]) ? 4'b0010 : 4'b0011;
																assign node14540 = (inp[8]) ? 4'b0011 : 4'b0010;
												assign node14543 = (inp[5]) ? node14565 : node14544;
													assign node14544 = (inp[8]) ? node14552 : node14545;
														assign node14545 = (inp[2]) ? node14547 : 4'b0010;
															assign node14547 = (inp[0]) ? 4'b0011 : node14548;
																assign node14548 = (inp[15]) ? 4'b0001 : 4'b0011;
														assign node14552 = (inp[2]) ? node14560 : node14553;
															assign node14553 = (inp[15]) ? node14557 : node14554;
																assign node14554 = (inp[0]) ? 4'b0001 : 4'b0011;
																assign node14557 = (inp[0]) ? 4'b0011 : 4'b0001;
															assign node14560 = (inp[15]) ? 4'b0010 : node14561;
																assign node14561 = (inp[0]) ? 4'b0000 : 4'b0010;
													assign node14565 = (inp[8]) ? node14579 : node14566;
														assign node14566 = (inp[2]) ? node14572 : node14567;
															assign node14567 = (inp[15]) ? node14569 : 4'b0010;
																assign node14569 = (inp[0]) ? 4'b0010 : 4'b0000;
															assign node14572 = (inp[0]) ? node14576 : node14573;
																assign node14573 = (inp[15]) ? 4'b0001 : 4'b0011;
																assign node14576 = (inp[15]) ? 4'b0011 : 4'b0001;
														assign node14579 = (inp[2]) ? 4'b0010 : 4'b0011;
											assign node14582 = (inp[2]) ? node14622 : node14583;
												assign node14583 = (inp[15]) ? node14603 : node14584;
													assign node14584 = (inp[0]) ? node14592 : node14585;
														assign node14585 = (inp[8]) ? node14589 : node14586;
															assign node14586 = (inp[7]) ? 4'b0010 : 4'b0011;
															assign node14589 = (inp[7]) ? 4'b0011 : 4'b0010;
														assign node14592 = (inp[5]) ? node14598 : node14593;
															assign node14593 = (inp[8]) ? 4'b0000 : node14594;
																assign node14594 = (inp[7]) ? 4'b0000 : 4'b0001;
															assign node14598 = (inp[8]) ? 4'b0001 : node14599;
																assign node14599 = (inp[7]) ? 4'b0000 : 4'b0001;
													assign node14603 = (inp[0]) ? node14615 : node14604;
														assign node14604 = (inp[5]) ? node14610 : node14605;
															assign node14605 = (inp[8]) ? node14607 : 4'b0001;
																assign node14607 = (inp[7]) ? 4'b0001 : 4'b0000;
															assign node14610 = (inp[8]) ? node14612 : 4'b0000;
																assign node14612 = (inp[7]) ? 4'b0001 : 4'b0000;
														assign node14615 = (inp[8]) ? node14619 : node14616;
															assign node14616 = (inp[7]) ? 4'b0010 : 4'b0011;
															assign node14619 = (inp[7]) ? 4'b0011 : 4'b0010;
												assign node14622 = (inp[8]) ? node14648 : node14623;
													assign node14623 = (inp[7]) ? node14637 : node14624;
														assign node14624 = (inp[5]) ? node14632 : node14625;
															assign node14625 = (inp[0]) ? node14629 : node14626;
																assign node14626 = (inp[15]) ? 4'b0000 : 4'b0010;
																assign node14629 = (inp[15]) ? 4'b0010 : 4'b0000;
															assign node14632 = (inp[0]) ? 4'b0010 : node14633;
																assign node14633 = (inp[15]) ? 4'b0000 : 4'b0010;
														assign node14637 = (inp[5]) ? node14643 : node14638;
															assign node14638 = (inp[15]) ? 4'b0011 : node14639;
																assign node14639 = (inp[0]) ? 4'b0001 : 4'b0011;
															assign node14643 = (inp[0]) ? 4'b0011 : node14644;
																assign node14644 = (inp[15]) ? 4'b0001 : 4'b0011;
													assign node14648 = (inp[7]) ? node14656 : node14649;
														assign node14649 = (inp[5]) ? 4'b0001 : node14650;
															assign node14650 = (inp[0]) ? 4'b0011 : node14651;
																assign node14651 = (inp[15]) ? 4'b0001 : 4'b0011;
														assign node14656 = (inp[0]) ? node14660 : node14657;
															assign node14657 = (inp[15]) ? 4'b0000 : 4'b0010;
															assign node14660 = (inp[15]) ? 4'b0010 : 4'b0000;
										assign node14663 = (inp[2]) ? node14721 : node14664;
											assign node14664 = (inp[5]) ? node14692 : node14665;
												assign node14665 = (inp[15]) ? node14681 : node14666;
													assign node14666 = (inp[0]) ? node14674 : node14667;
														assign node14667 = (inp[8]) ? node14671 : node14668;
															assign node14668 = (inp[7]) ? 4'b0010 : 4'b0011;
															assign node14671 = (inp[7]) ? 4'b0011 : 4'b0010;
														assign node14674 = (inp[10]) ? node14676 : 4'b0000;
															assign node14676 = (inp[8]) ? 4'b0001 : node14677;
																assign node14677 = (inp[7]) ? 4'b0000 : 4'b0001;
													assign node14681 = (inp[0]) ? node14687 : node14682;
														assign node14682 = (inp[10]) ? node14684 : 4'b0001;
															assign node14684 = (inp[7]) ? 4'b0000 : 4'b0001;
														assign node14687 = (inp[7]) ? node14689 : 4'b0011;
															assign node14689 = (inp[8]) ? 4'b0011 : 4'b0010;
												assign node14692 = (inp[0]) ? node14708 : node14693;
													assign node14693 = (inp[15]) ? node14701 : node14694;
														assign node14694 = (inp[7]) ? node14698 : node14695;
															assign node14695 = (inp[8]) ? 4'b0000 : 4'b0001;
															assign node14698 = (inp[8]) ? 4'b0001 : 4'b0000;
														assign node14701 = (inp[10]) ? node14703 : 4'b0011;
															assign node14703 = (inp[7]) ? node14705 : 4'b0010;
																assign node14705 = (inp[8]) ? 4'b0011 : 4'b0010;
													assign node14708 = (inp[15]) ? node14716 : node14709;
														assign node14709 = (inp[7]) ? node14713 : node14710;
															assign node14710 = (inp[8]) ? 4'b0010 : 4'b0011;
															assign node14713 = (inp[8]) ? 4'b0011 : 4'b0010;
														assign node14716 = (inp[7]) ? node14718 : 4'b0000;
															assign node14718 = (inp[8]) ? 4'b0001 : 4'b0000;
											assign node14721 = (inp[15]) ? node14751 : node14722;
												assign node14722 = (inp[7]) ? node14732 : node14723;
													assign node14723 = (inp[8]) ? node14725 : 4'b0000;
														assign node14725 = (inp[5]) ? node14729 : node14726;
															assign node14726 = (inp[0]) ? 4'b0001 : 4'b0011;
															assign node14729 = (inp[0]) ? 4'b0011 : 4'b0001;
													assign node14732 = (inp[8]) ? node14744 : node14733;
														assign node14733 = (inp[10]) ? node14739 : node14734;
															assign node14734 = (inp[0]) ? 4'b0001 : node14735;
																assign node14735 = (inp[5]) ? 4'b0001 : 4'b0011;
															assign node14739 = (inp[5]) ? 4'b0011 : node14740;
																assign node14740 = (inp[0]) ? 4'b0001 : 4'b0011;
														assign node14744 = (inp[10]) ? 4'b0000 : node14745;
															assign node14745 = (inp[0]) ? 4'b0010 : node14746;
																assign node14746 = (inp[5]) ? 4'b0000 : 4'b0010;
												assign node14751 = (inp[8]) ? node14773 : node14752;
													assign node14752 = (inp[7]) ? node14762 : node14753;
														assign node14753 = (inp[10]) ? 4'b0000 : node14754;
															assign node14754 = (inp[0]) ? node14758 : node14755;
																assign node14755 = (inp[5]) ? 4'b0010 : 4'b0000;
																assign node14758 = (inp[5]) ? 4'b0000 : 4'b0010;
														assign node14762 = (inp[10]) ? node14768 : node14763;
															assign node14763 = (inp[5]) ? 4'b0011 : node14764;
																assign node14764 = (inp[0]) ? 4'b0011 : 4'b0001;
															assign node14768 = (inp[0]) ? node14770 : 4'b0001;
																assign node14770 = (inp[5]) ? 4'b0001 : 4'b0011;
													assign node14773 = (inp[7]) ? node14781 : node14774;
														assign node14774 = (inp[0]) ? node14778 : node14775;
															assign node14775 = (inp[5]) ? 4'b0011 : 4'b0001;
															assign node14778 = (inp[5]) ? 4'b0001 : 4'b0011;
														assign node14781 = (inp[10]) ? node14789 : node14782;
															assign node14782 = (inp[0]) ? node14786 : node14783;
																assign node14783 = (inp[5]) ? 4'b0010 : 4'b0000;
																assign node14786 = (inp[5]) ? 4'b0000 : 4'b0010;
															assign node14789 = (inp[0]) ? 4'b0010 : node14790;
																assign node14790 = (inp[5]) ? 4'b0010 : 4'b0000;
									assign node14794 = (inp[7]) ? node14882 : node14795;
										assign node14795 = (inp[8]) ? node14859 : node14796;
											assign node14796 = (inp[5]) ? node14824 : node14797;
												assign node14797 = (inp[3]) ? node14805 : node14798;
													assign node14798 = (inp[0]) ? node14802 : node14799;
														assign node14799 = (inp[15]) ? 4'b0000 : 4'b0010;
														assign node14802 = (inp[15]) ? 4'b0010 : 4'b0000;
													assign node14805 = (inp[2]) ? node14811 : node14806;
														assign node14806 = (inp[0]) ? 4'b0010 : node14807;
															assign node14807 = (inp[15]) ? 4'b0000 : 4'b0010;
														assign node14811 = (inp[10]) ? node14819 : node14812;
															assign node14812 = (inp[0]) ? node14816 : node14813;
																assign node14813 = (inp[15]) ? 4'b0000 : 4'b0010;
																assign node14816 = (inp[15]) ? 4'b0010 : 4'b0000;
															assign node14819 = (inp[15]) ? 4'b0010 : node14820;
																assign node14820 = (inp[0]) ? 4'b0000 : 4'b0010;
												assign node14824 = (inp[3]) ? node14854 : node14825;
													assign node14825 = (inp[10]) ? node14839 : node14826;
														assign node14826 = (inp[2]) ? node14834 : node14827;
															assign node14827 = (inp[0]) ? node14831 : node14828;
																assign node14828 = (inp[15]) ? 4'b0000 : 4'b0010;
																assign node14831 = (inp[15]) ? 4'b0010 : 4'b0000;
															assign node14834 = (inp[0]) ? node14836 : 4'b0000;
																assign node14836 = (inp[15]) ? 4'b0010 : 4'b0000;
														assign node14839 = (inp[2]) ? node14847 : node14840;
															assign node14840 = (inp[15]) ? node14844 : node14841;
																assign node14841 = (inp[0]) ? 4'b0000 : 4'b0010;
																assign node14844 = (inp[0]) ? 4'b0010 : 4'b0000;
															assign node14847 = (inp[0]) ? node14851 : node14848;
																assign node14848 = (inp[15]) ? 4'b0000 : 4'b0010;
																assign node14851 = (inp[15]) ? 4'b0010 : 4'b0000;
													assign node14854 = (inp[0]) ? 4'b0000 : node14855;
														assign node14855 = (inp[15]) ? 4'b0010 : 4'b0000;
											assign node14859 = (inp[0]) ? node14871 : node14860;
												assign node14860 = (inp[15]) ? node14866 : node14861;
													assign node14861 = (inp[5]) ? node14863 : 4'b0011;
														assign node14863 = (inp[3]) ? 4'b0001 : 4'b0011;
													assign node14866 = (inp[3]) ? node14868 : 4'b0001;
														assign node14868 = (inp[5]) ? 4'b0011 : 4'b0001;
												assign node14871 = (inp[15]) ? node14877 : node14872;
													assign node14872 = (inp[3]) ? node14874 : 4'b0001;
														assign node14874 = (inp[5]) ? 4'b0011 : 4'b0001;
													assign node14877 = (inp[5]) ? node14879 : 4'b0011;
														assign node14879 = (inp[3]) ? 4'b0001 : 4'b0011;
										assign node14882 = (inp[8]) ? node14918 : node14883;
											assign node14883 = (inp[10]) ? node14901 : node14884;
												assign node14884 = (inp[15]) ? node14896 : node14885;
													assign node14885 = (inp[0]) ? node14891 : node14886;
														assign node14886 = (inp[5]) ? node14888 : 4'b0011;
															assign node14888 = (inp[3]) ? 4'b0001 : 4'b0011;
														assign node14891 = (inp[3]) ? node14893 : 4'b0001;
															assign node14893 = (inp[5]) ? 4'b0011 : 4'b0001;
													assign node14896 = (inp[0]) ? 4'b0011 : node14897;
														assign node14897 = (inp[3]) ? 4'b0011 : 4'b0001;
												assign node14901 = (inp[15]) ? node14907 : node14902;
													assign node14902 = (inp[0]) ? node14904 : 4'b0011;
														assign node14904 = (inp[5]) ? 4'b0011 : 4'b0001;
													assign node14907 = (inp[0]) ? node14913 : node14908;
														assign node14908 = (inp[5]) ? node14910 : 4'b0001;
															assign node14910 = (inp[3]) ? 4'b0011 : 4'b0001;
														assign node14913 = (inp[3]) ? node14915 : 4'b0011;
															assign node14915 = (inp[5]) ? 4'b0001 : 4'b0011;
											assign node14918 = (inp[2]) ? node14942 : node14919;
												assign node14919 = (inp[0]) ? node14931 : node14920;
													assign node14920 = (inp[15]) ? node14926 : node14921;
														assign node14921 = (inp[3]) ? node14923 : 4'b0010;
															assign node14923 = (inp[5]) ? 4'b0000 : 4'b0010;
														assign node14926 = (inp[3]) ? node14928 : 4'b0000;
															assign node14928 = (inp[5]) ? 4'b0010 : 4'b0000;
													assign node14931 = (inp[15]) ? node14937 : node14932;
														assign node14932 = (inp[5]) ? node14934 : 4'b0000;
															assign node14934 = (inp[3]) ? 4'b0010 : 4'b0000;
														assign node14937 = (inp[3]) ? node14939 : 4'b0010;
															assign node14939 = (inp[5]) ? 4'b0000 : 4'b0010;
												assign node14942 = (inp[3]) ? node14950 : node14943;
													assign node14943 = (inp[0]) ? node14947 : node14944;
														assign node14944 = (inp[15]) ? 4'b0000 : 4'b0010;
														assign node14947 = (inp[15]) ? 4'b0010 : 4'b0000;
													assign node14950 = (inp[0]) ? node14956 : node14951;
														assign node14951 = (inp[15]) ? node14953 : 4'b0000;
															assign node14953 = (inp[5]) ? 4'b0010 : 4'b0000;
														assign node14956 = (inp[15]) ? node14960 : node14957;
															assign node14957 = (inp[5]) ? 4'b0010 : 4'b0000;
															assign node14960 = (inp[5]) ? 4'b0000 : 4'b0010;
								assign node14963 = (inp[10]) ? node15187 : node14964;
									assign node14964 = (inp[0]) ? node15064 : node14965;
										assign node14965 = (inp[15]) ? node15021 : node14966;
											assign node14966 = (inp[3]) ? node14990 : node14967;
												assign node14967 = (inp[14]) ? node14983 : node14968;
													assign node14968 = (inp[2]) ? node14976 : node14969;
														assign node14969 = (inp[7]) ? node14973 : node14970;
															assign node14970 = (inp[8]) ? 4'b0010 : 4'b0011;
															assign node14973 = (inp[8]) ? 4'b0011 : 4'b0010;
														assign node14976 = (inp[7]) ? node14980 : node14977;
															assign node14977 = (inp[8]) ? 4'b0011 : 4'b0010;
															assign node14980 = (inp[8]) ? 4'b0010 : 4'b0011;
													assign node14983 = (inp[7]) ? node14987 : node14984;
														assign node14984 = (inp[8]) ? 4'b0011 : 4'b0010;
														assign node14987 = (inp[8]) ? 4'b0010 : 4'b0011;
												assign node14990 = (inp[5]) ? node15002 : node14991;
													assign node14991 = (inp[7]) ? node14997 : node14992;
														assign node14992 = (inp[8]) ? 4'b0011 : node14993;
															assign node14993 = (inp[2]) ? 4'b0010 : 4'b0011;
														assign node14997 = (inp[8]) ? 4'b0010 : node14998;
															assign node14998 = (inp[14]) ? 4'b0011 : 4'b0010;
													assign node15002 = (inp[14]) ? node15012 : node15003;
														assign node15003 = (inp[8]) ? 4'b0000 : node15004;
															assign node15004 = (inp[7]) ? node15008 : node15005;
																assign node15005 = (inp[2]) ? 4'b0000 : 4'b0001;
																assign node15008 = (inp[2]) ? 4'b0001 : 4'b0000;
														assign node15012 = (inp[2]) ? 4'b0001 : node15013;
															assign node15013 = (inp[8]) ? node15017 : node15014;
																assign node15014 = (inp[7]) ? 4'b0001 : 4'b0000;
																assign node15017 = (inp[7]) ? 4'b0000 : 4'b0001;
											assign node15021 = (inp[5]) ? node15047 : node15022;
												assign node15022 = (inp[14]) ? node15040 : node15023;
													assign node15023 = (inp[7]) ? node15033 : node15024;
														assign node15024 = (inp[3]) ? node15026 : 4'b0000;
															assign node15026 = (inp[2]) ? node15030 : node15027;
																assign node15027 = (inp[8]) ? 4'b0000 : 4'b0001;
																assign node15030 = (inp[8]) ? 4'b0001 : 4'b0000;
														assign node15033 = (inp[2]) ? node15037 : node15034;
															assign node15034 = (inp[8]) ? 4'b0001 : 4'b0000;
															assign node15037 = (inp[8]) ? 4'b0000 : 4'b0001;
													assign node15040 = (inp[7]) ? node15044 : node15041;
														assign node15041 = (inp[8]) ? 4'b0001 : 4'b0000;
														assign node15044 = (inp[8]) ? 4'b0000 : 4'b0001;
												assign node15047 = (inp[3]) ? node15051 : node15048;
													assign node15048 = (inp[8]) ? 4'b0000 : 4'b0001;
													assign node15051 = (inp[7]) ? 4'b0010 : node15052;
														assign node15052 = (inp[8]) ? node15058 : node15053;
															assign node15053 = (inp[2]) ? 4'b0010 : node15054;
																assign node15054 = (inp[14]) ? 4'b0010 : 4'b0011;
															assign node15058 = (inp[2]) ? 4'b0011 : node15059;
																assign node15059 = (inp[14]) ? 4'b0011 : 4'b0010;
										assign node15064 = (inp[15]) ? node15144 : node15065;
											assign node15065 = (inp[3]) ? node15105 : node15066;
												assign node15066 = (inp[14]) ? node15098 : node15067;
													assign node15067 = (inp[8]) ? node15083 : node15068;
														assign node15068 = (inp[5]) ? node15076 : node15069;
															assign node15069 = (inp[2]) ? node15073 : node15070;
																assign node15070 = (inp[7]) ? 4'b0000 : 4'b0001;
																assign node15073 = (inp[7]) ? 4'b0001 : 4'b0000;
															assign node15076 = (inp[7]) ? node15080 : node15077;
																assign node15077 = (inp[2]) ? 4'b0000 : 4'b0001;
																assign node15080 = (inp[2]) ? 4'b0001 : 4'b0000;
														assign node15083 = (inp[5]) ? node15091 : node15084;
															assign node15084 = (inp[7]) ? node15088 : node15085;
																assign node15085 = (inp[2]) ? 4'b0001 : 4'b0000;
																assign node15088 = (inp[2]) ? 4'b0000 : 4'b0001;
															assign node15091 = (inp[7]) ? node15095 : node15092;
																assign node15092 = (inp[2]) ? 4'b0001 : 4'b0000;
																assign node15095 = (inp[2]) ? 4'b0000 : 4'b0001;
													assign node15098 = (inp[7]) ? node15102 : node15099;
														assign node15099 = (inp[8]) ? 4'b0001 : 4'b0000;
														assign node15102 = (inp[8]) ? 4'b0000 : 4'b0001;
												assign node15105 = (inp[5]) ? node15125 : node15106;
													assign node15106 = (inp[14]) ? node15120 : node15107;
														assign node15107 = (inp[2]) ? node15113 : node15108;
															assign node15108 = (inp[7]) ? 4'b0001 : node15109;
																assign node15109 = (inp[8]) ? 4'b0000 : 4'b0001;
															assign node15113 = (inp[8]) ? node15117 : node15114;
																assign node15114 = (inp[7]) ? 4'b0001 : 4'b0000;
																assign node15117 = (inp[7]) ? 4'b0000 : 4'b0001;
														assign node15120 = (inp[7]) ? node15122 : 4'b0000;
															assign node15122 = (inp[8]) ? 4'b0000 : 4'b0001;
													assign node15125 = (inp[7]) ? node15133 : node15126;
														assign node15126 = (inp[8]) ? node15128 : 4'b0010;
															assign node15128 = (inp[2]) ? 4'b0011 : node15129;
																assign node15129 = (inp[14]) ? 4'b0011 : 4'b0010;
														assign node15133 = (inp[8]) ? node15139 : node15134;
															assign node15134 = (inp[2]) ? 4'b0011 : node15135;
																assign node15135 = (inp[14]) ? 4'b0011 : 4'b0010;
															assign node15139 = (inp[14]) ? 4'b0010 : node15140;
																assign node15140 = (inp[2]) ? 4'b0010 : 4'b0011;
											assign node15144 = (inp[5]) ? node15160 : node15145;
												assign node15145 = (inp[7]) ? node15153 : node15146;
													assign node15146 = (inp[8]) ? node15148 : 4'b0010;
														assign node15148 = (inp[14]) ? 4'b0011 : node15149;
															assign node15149 = (inp[2]) ? 4'b0011 : 4'b0010;
													assign node15153 = (inp[8]) ? node15155 : 4'b0011;
														assign node15155 = (inp[2]) ? 4'b0010 : node15156;
															assign node15156 = (inp[14]) ? 4'b0010 : 4'b0011;
												assign node15160 = (inp[3]) ? node15174 : node15161;
													assign node15161 = (inp[14]) ? 4'b0010 : node15162;
														assign node15162 = (inp[8]) ? node15168 : node15163;
															assign node15163 = (inp[7]) ? node15165 : 4'b0010;
																assign node15165 = (inp[2]) ? 4'b0011 : 4'b0010;
															assign node15168 = (inp[7]) ? node15170 : 4'b0011;
																assign node15170 = (inp[2]) ? 4'b0010 : 4'b0011;
													assign node15174 = (inp[7]) ? node15182 : node15175;
														assign node15175 = (inp[8]) ? node15179 : node15176;
															assign node15176 = (inp[2]) ? 4'b0000 : 4'b0001;
															assign node15179 = (inp[2]) ? 4'b0001 : 4'b0000;
														assign node15182 = (inp[14]) ? node15184 : 4'b0001;
															assign node15184 = (inp[2]) ? 4'b0001 : 4'b0000;
									assign node15187 = (inp[7]) ? node15317 : node15188;
										assign node15188 = (inp[8]) ? node15260 : node15189;
											assign node15189 = (inp[2]) ? node15221 : node15190;
												assign node15190 = (inp[14]) ? node15202 : node15191;
													assign node15191 = (inp[3]) ? node15197 : node15192;
														assign node15192 = (inp[0]) ? 4'b0111 : node15193;
															assign node15193 = (inp[15]) ? 4'b0111 : 4'b0101;
														assign node15197 = (inp[0]) ? 4'b0101 : node15198;
															assign node15198 = (inp[15]) ? 4'b0111 : 4'b0101;
													assign node15202 = (inp[0]) ? node15214 : node15203;
														assign node15203 = (inp[15]) ? node15209 : node15204;
															assign node15204 = (inp[5]) ? 4'b0100 : node15205;
																assign node15205 = (inp[3]) ? 4'b0100 : 4'b0110;
															assign node15209 = (inp[3]) ? 4'b0110 : node15210;
																assign node15210 = (inp[5]) ? 4'b0110 : 4'b0100;
														assign node15214 = (inp[15]) ? 4'b0100 : node15215;
															assign node15215 = (inp[5]) ? 4'b0110 : node15216;
																assign node15216 = (inp[3]) ? 4'b0110 : 4'b0100;
												assign node15221 = (inp[3]) ? node15245 : node15222;
													assign node15222 = (inp[14]) ? node15236 : node15223;
														assign node15223 = (inp[15]) ? node15229 : node15224;
															assign node15224 = (inp[5]) ? 4'b0110 : node15225;
																assign node15225 = (inp[0]) ? 4'b0100 : 4'b0110;
															assign node15229 = (inp[0]) ? node15233 : node15230;
																assign node15230 = (inp[5]) ? 4'b0110 : 4'b0100;
																assign node15233 = (inp[5]) ? 4'b0100 : 4'b0110;
														assign node15236 = (inp[15]) ? 4'b0110 : node15237;
															assign node15237 = (inp[0]) ? node15241 : node15238;
																assign node15238 = (inp[5]) ? 4'b0100 : 4'b0110;
																assign node15241 = (inp[5]) ? 4'b0110 : 4'b0100;
													assign node15245 = (inp[5]) ? node15253 : node15246;
														assign node15246 = (inp[0]) ? node15250 : node15247;
															assign node15247 = (inp[15]) ? 4'b0110 : 4'b0100;
															assign node15250 = (inp[15]) ? 4'b0100 : 4'b0110;
														assign node15253 = (inp[15]) ? node15257 : node15254;
															assign node15254 = (inp[0]) ? 4'b0110 : 4'b0100;
															assign node15257 = (inp[0]) ? 4'b0100 : 4'b0110;
											assign node15260 = (inp[14]) ? node15298 : node15261;
												assign node15261 = (inp[2]) ? node15285 : node15262;
													assign node15262 = (inp[3]) ? node15276 : node15263;
														assign node15263 = (inp[0]) ? node15269 : node15264;
															assign node15264 = (inp[15]) ? 4'b0110 : node15265;
																assign node15265 = (inp[5]) ? 4'b0100 : 4'b0110;
															assign node15269 = (inp[15]) ? node15273 : node15270;
																assign node15270 = (inp[5]) ? 4'b0110 : 4'b0100;
																assign node15273 = (inp[5]) ? 4'b0100 : 4'b0110;
														assign node15276 = (inp[5]) ? node15282 : node15277;
															assign node15277 = (inp[15]) ? node15279 : 4'b0100;
																assign node15279 = (inp[0]) ? 4'b0100 : 4'b0110;
															assign node15282 = (inp[15]) ? 4'b0100 : 4'b0110;
													assign node15285 = (inp[0]) ? node15291 : node15286;
														assign node15286 = (inp[15]) ? node15288 : 4'b0101;
															assign node15288 = (inp[3]) ? 4'b0111 : 4'b0101;
														assign node15291 = (inp[15]) ? node15293 : 4'b0111;
															assign node15293 = (inp[5]) ? 4'b0101 : node15294;
																assign node15294 = (inp[3]) ? 4'b0101 : 4'b0111;
												assign node15298 = (inp[15]) ? node15310 : node15299;
													assign node15299 = (inp[0]) ? node15305 : node15300;
														assign node15300 = (inp[3]) ? 4'b0101 : node15301;
															assign node15301 = (inp[5]) ? 4'b0101 : 4'b0111;
														assign node15305 = (inp[3]) ? 4'b0111 : node15306;
															assign node15306 = (inp[5]) ? 4'b0111 : 4'b0101;
													assign node15310 = (inp[0]) ? node15312 : 4'b0111;
														assign node15312 = (inp[3]) ? 4'b0101 : node15313;
															assign node15313 = (inp[5]) ? 4'b0101 : 4'b0111;
										assign node15317 = (inp[8]) ? node15379 : node15318;
											assign node15318 = (inp[14]) ? node15352 : node15319;
												assign node15319 = (inp[2]) ? node15335 : node15320;
													assign node15320 = (inp[3]) ? node15328 : node15321;
														assign node15321 = (inp[15]) ? 4'b0110 : node15322;
															assign node15322 = (inp[5]) ? node15324 : 4'b0110;
																assign node15324 = (inp[0]) ? 4'b0110 : 4'b0100;
														assign node15328 = (inp[15]) ? node15332 : node15329;
															assign node15329 = (inp[0]) ? 4'b0110 : 4'b0100;
															assign node15332 = (inp[0]) ? 4'b0100 : 4'b0110;
													assign node15335 = (inp[15]) ? node15347 : node15336;
														assign node15336 = (inp[0]) ? node15342 : node15337;
															assign node15337 = (inp[3]) ? 4'b0101 : node15338;
																assign node15338 = (inp[5]) ? 4'b0101 : 4'b0111;
															assign node15342 = (inp[3]) ? 4'b0111 : node15343;
																assign node15343 = (inp[5]) ? 4'b0111 : 4'b0101;
														assign node15347 = (inp[0]) ? 4'b0101 : node15348;
															assign node15348 = (inp[3]) ? 4'b0111 : 4'b0101;
												assign node15352 = (inp[3]) ? node15372 : node15353;
													assign node15353 = (inp[5]) ? node15363 : node15354;
														assign node15354 = (inp[2]) ? node15356 : 4'b0101;
															assign node15356 = (inp[15]) ? node15360 : node15357;
																assign node15357 = (inp[0]) ? 4'b0101 : 4'b0111;
																assign node15360 = (inp[0]) ? 4'b0111 : 4'b0101;
														assign node15363 = (inp[2]) ? 4'b0111 : node15364;
															assign node15364 = (inp[15]) ? node15368 : node15365;
																assign node15365 = (inp[0]) ? 4'b0111 : 4'b0101;
																assign node15368 = (inp[0]) ? 4'b0101 : 4'b0111;
													assign node15372 = (inp[15]) ? node15376 : node15373;
														assign node15373 = (inp[0]) ? 4'b0111 : 4'b0101;
														assign node15376 = (inp[0]) ? 4'b0101 : 4'b0111;
											assign node15379 = (inp[2]) ? node15415 : node15380;
												assign node15380 = (inp[14]) ? node15402 : node15381;
													assign node15381 = (inp[5]) ? node15395 : node15382;
														assign node15382 = (inp[3]) ? node15390 : node15383;
															assign node15383 = (inp[15]) ? node15387 : node15384;
																assign node15384 = (inp[0]) ? 4'b0101 : 4'b0111;
																assign node15387 = (inp[0]) ? 4'b0111 : 4'b0101;
															assign node15390 = (inp[0]) ? node15392 : 4'b0101;
																assign node15392 = (inp[15]) ? 4'b0101 : 4'b0111;
														assign node15395 = (inp[0]) ? node15399 : node15396;
															assign node15396 = (inp[15]) ? 4'b0111 : 4'b0101;
															assign node15399 = (inp[15]) ? 4'b0101 : 4'b0111;
													assign node15402 = (inp[5]) ? node15410 : node15403;
														assign node15403 = (inp[3]) ? node15405 : 4'b0110;
															assign node15405 = (inp[15]) ? 4'b0100 : node15406;
																assign node15406 = (inp[0]) ? 4'b0110 : 4'b0100;
														assign node15410 = (inp[0]) ? 4'b0100 : node15411;
															assign node15411 = (inp[15]) ? 4'b0110 : 4'b0100;
												assign node15415 = (inp[15]) ? node15427 : node15416;
													assign node15416 = (inp[0]) ? node15422 : node15417;
														assign node15417 = (inp[3]) ? 4'b0100 : node15418;
															assign node15418 = (inp[5]) ? 4'b0100 : 4'b0110;
														assign node15422 = (inp[3]) ? 4'b0110 : node15423;
															assign node15423 = (inp[5]) ? 4'b0110 : 4'b0100;
													assign node15427 = (inp[0]) ? node15433 : node15428;
														assign node15428 = (inp[3]) ? 4'b0110 : node15429;
															assign node15429 = (inp[5]) ? 4'b0110 : 4'b0100;
														assign node15433 = (inp[5]) ? 4'b0100 : node15434;
															assign node15434 = (inp[3]) ? 4'b0100 : 4'b0110;
							assign node15438 = (inp[12]) ? node16050 : node15439;
								assign node15439 = (inp[2]) ? node15777 : node15440;
									assign node15440 = (inp[5]) ? node15636 : node15441;
										assign node15441 = (inp[14]) ? node15541 : node15442;
											assign node15442 = (inp[0]) ? node15492 : node15443;
												assign node15443 = (inp[10]) ? node15469 : node15444;
													assign node15444 = (inp[15]) ? node15456 : node15445;
														assign node15445 = (inp[3]) ? node15453 : node15446;
															assign node15446 = (inp[8]) ? node15450 : node15447;
																assign node15447 = (inp[7]) ? 4'b0110 : 4'b0111;
																assign node15450 = (inp[7]) ? 4'b0111 : 4'b0110;
															assign node15453 = (inp[8]) ? 4'b0100 : 4'b0101;
														assign node15456 = (inp[3]) ? node15462 : node15457;
															assign node15457 = (inp[7]) ? node15459 : 4'b0100;
																assign node15459 = (inp[8]) ? 4'b0101 : 4'b0100;
															assign node15462 = (inp[7]) ? node15466 : node15463;
																assign node15463 = (inp[8]) ? 4'b0110 : 4'b0111;
																assign node15466 = (inp[8]) ? 4'b0111 : 4'b0110;
													assign node15469 = (inp[3]) ? node15479 : node15470;
														assign node15470 = (inp[15]) ? node15474 : node15471;
															assign node15471 = (inp[8]) ? 4'b0111 : 4'b0110;
															assign node15474 = (inp[8]) ? node15476 : 4'b0101;
																assign node15476 = (inp[7]) ? 4'b0101 : 4'b0100;
														assign node15479 = (inp[15]) ? node15487 : node15480;
															assign node15480 = (inp[7]) ? node15484 : node15481;
																assign node15481 = (inp[8]) ? 4'b0100 : 4'b0101;
																assign node15484 = (inp[8]) ? 4'b0101 : 4'b0100;
															assign node15487 = (inp[8]) ? 4'b0110 : node15488;
																assign node15488 = (inp[7]) ? 4'b0110 : 4'b0111;
												assign node15492 = (inp[10]) ? node15518 : node15493;
													assign node15493 = (inp[3]) ? node15503 : node15494;
														assign node15494 = (inp[15]) ? 4'b0111 : node15495;
															assign node15495 = (inp[8]) ? node15499 : node15496;
																assign node15496 = (inp[7]) ? 4'b0100 : 4'b0101;
																assign node15499 = (inp[7]) ? 4'b0101 : 4'b0100;
														assign node15503 = (inp[15]) ? node15511 : node15504;
															assign node15504 = (inp[8]) ? node15508 : node15505;
																assign node15505 = (inp[7]) ? 4'b0110 : 4'b0111;
																assign node15508 = (inp[7]) ? 4'b0111 : 4'b0110;
															assign node15511 = (inp[7]) ? node15515 : node15512;
																assign node15512 = (inp[8]) ? 4'b0100 : 4'b0101;
																assign node15515 = (inp[8]) ? 4'b0101 : 4'b0100;
													assign node15518 = (inp[8]) ? node15534 : node15519;
														assign node15519 = (inp[7]) ? node15527 : node15520;
															assign node15520 = (inp[3]) ? node15524 : node15521;
																assign node15521 = (inp[15]) ? 4'b0111 : 4'b0101;
																assign node15524 = (inp[15]) ? 4'b0101 : 4'b0111;
															assign node15527 = (inp[15]) ? node15531 : node15528;
																assign node15528 = (inp[3]) ? 4'b0110 : 4'b0100;
																assign node15531 = (inp[3]) ? 4'b0100 : 4'b0110;
														assign node15534 = (inp[7]) ? node15536 : 4'b0110;
															assign node15536 = (inp[3]) ? node15538 : 4'b0111;
																assign node15538 = (inp[15]) ? 4'b0101 : 4'b0111;
											assign node15541 = (inp[10]) ? node15593 : node15542;
												assign node15542 = (inp[7]) ? node15570 : node15543;
													assign node15543 = (inp[8]) ? node15557 : node15544;
														assign node15544 = (inp[15]) ? node15550 : node15545;
															assign node15545 = (inp[0]) ? 4'b0110 : node15546;
																assign node15546 = (inp[3]) ? 4'b0100 : 4'b0110;
															assign node15550 = (inp[0]) ? node15554 : node15551;
																assign node15551 = (inp[3]) ? 4'b0110 : 4'b0100;
																assign node15554 = (inp[3]) ? 4'b0100 : 4'b0110;
														assign node15557 = (inp[0]) ? node15563 : node15558;
															assign node15558 = (inp[15]) ? node15560 : 4'b0111;
																assign node15560 = (inp[3]) ? 4'b0111 : 4'b0101;
															assign node15563 = (inp[15]) ? node15567 : node15564;
																assign node15564 = (inp[3]) ? 4'b0111 : 4'b0101;
																assign node15567 = (inp[3]) ? 4'b0101 : 4'b0111;
													assign node15570 = (inp[8]) ? node15578 : node15571;
														assign node15571 = (inp[0]) ? 4'b0101 : node15572;
															assign node15572 = (inp[3]) ? node15574 : 4'b0111;
																assign node15574 = (inp[15]) ? 4'b0111 : 4'b0101;
														assign node15578 = (inp[15]) ? node15586 : node15579;
															assign node15579 = (inp[3]) ? node15583 : node15580;
																assign node15580 = (inp[0]) ? 4'b0100 : 4'b0110;
																assign node15583 = (inp[0]) ? 4'b0110 : 4'b0100;
															assign node15586 = (inp[0]) ? node15590 : node15587;
																assign node15587 = (inp[3]) ? 4'b0110 : 4'b0100;
																assign node15590 = (inp[3]) ? 4'b0100 : 4'b0110;
												assign node15593 = (inp[3]) ? node15613 : node15594;
													assign node15594 = (inp[7]) ? node15606 : node15595;
														assign node15595 = (inp[8]) ? node15599 : node15596;
															assign node15596 = (inp[15]) ? 4'b0100 : 4'b0110;
															assign node15599 = (inp[15]) ? node15603 : node15600;
																assign node15600 = (inp[0]) ? 4'b0101 : 4'b0111;
																assign node15603 = (inp[0]) ? 4'b0111 : 4'b0101;
														assign node15606 = (inp[8]) ? node15608 : 4'b0111;
															assign node15608 = (inp[15]) ? node15610 : 4'b0110;
																assign node15610 = (inp[0]) ? 4'b0110 : 4'b0100;
													assign node15613 = (inp[0]) ? node15627 : node15614;
														assign node15614 = (inp[15]) ? node15620 : node15615;
															assign node15615 = (inp[8]) ? 4'b0100 : node15616;
																assign node15616 = (inp[7]) ? 4'b0101 : 4'b0100;
															assign node15620 = (inp[8]) ? node15624 : node15621;
																assign node15621 = (inp[7]) ? 4'b0111 : 4'b0110;
																assign node15624 = (inp[7]) ? 4'b0110 : 4'b0111;
														assign node15627 = (inp[15]) ? 4'b0100 : node15628;
															assign node15628 = (inp[7]) ? node15632 : node15629;
																assign node15629 = (inp[8]) ? 4'b0111 : 4'b0110;
																assign node15632 = (inp[8]) ? 4'b0110 : 4'b0111;
										assign node15636 = (inp[14]) ? node15702 : node15637;
											assign node15637 = (inp[3]) ? node15673 : node15638;
												assign node15638 = (inp[15]) ? node15658 : node15639;
													assign node15639 = (inp[0]) ? node15643 : node15640;
														assign node15640 = (inp[7]) ? 4'b0101 : 4'b0100;
														assign node15643 = (inp[10]) ? node15651 : node15644;
															assign node15644 = (inp[8]) ? node15648 : node15645;
																assign node15645 = (inp[7]) ? 4'b0110 : 4'b0111;
																assign node15648 = (inp[7]) ? 4'b0111 : 4'b0110;
															assign node15651 = (inp[7]) ? node15655 : node15652;
																assign node15652 = (inp[8]) ? 4'b0110 : 4'b0111;
																assign node15655 = (inp[8]) ? 4'b0111 : 4'b0110;
													assign node15658 = (inp[0]) ? node15666 : node15659;
														assign node15659 = (inp[8]) ? node15663 : node15660;
															assign node15660 = (inp[7]) ? 4'b0110 : 4'b0111;
															assign node15663 = (inp[7]) ? 4'b0111 : 4'b0110;
														assign node15666 = (inp[10]) ? node15668 : 4'b0100;
															assign node15668 = (inp[8]) ? 4'b0101 : node15669;
																assign node15669 = (inp[7]) ? 4'b0100 : 4'b0101;
												assign node15673 = (inp[7]) ? node15689 : node15674;
													assign node15674 = (inp[8]) ? node15682 : node15675;
														assign node15675 = (inp[10]) ? node15677 : 4'b0101;
															assign node15677 = (inp[0]) ? node15679 : 4'b0111;
																assign node15679 = (inp[15]) ? 4'b0101 : 4'b0111;
														assign node15682 = (inp[15]) ? node15686 : node15683;
															assign node15683 = (inp[0]) ? 4'b0110 : 4'b0100;
															assign node15686 = (inp[0]) ? 4'b0100 : 4'b0110;
													assign node15689 = (inp[8]) ? node15695 : node15690;
														assign node15690 = (inp[0]) ? node15692 : 4'b0110;
															assign node15692 = (inp[10]) ? 4'b0100 : 4'b0110;
														assign node15695 = (inp[0]) ? node15699 : node15696;
															assign node15696 = (inp[15]) ? 4'b0111 : 4'b0101;
															assign node15699 = (inp[15]) ? 4'b0101 : 4'b0111;
											assign node15702 = (inp[3]) ? node15748 : node15703;
												assign node15703 = (inp[15]) ? node15725 : node15704;
													assign node15704 = (inp[0]) ? node15718 : node15705;
														assign node15705 = (inp[10]) ? node15711 : node15706;
															assign node15706 = (inp[7]) ? 4'b0100 : node15707;
																assign node15707 = (inp[8]) ? 4'b0101 : 4'b0100;
															assign node15711 = (inp[7]) ? node15715 : node15712;
																assign node15712 = (inp[8]) ? 4'b0101 : 4'b0100;
																assign node15715 = (inp[8]) ? 4'b0100 : 4'b0101;
														assign node15718 = (inp[10]) ? 4'b0111 : node15719;
															assign node15719 = (inp[7]) ? 4'b0110 : node15720;
																assign node15720 = (inp[8]) ? 4'b0111 : 4'b0110;
													assign node15725 = (inp[0]) ? node15739 : node15726;
														assign node15726 = (inp[10]) ? node15734 : node15727;
															assign node15727 = (inp[8]) ? node15731 : node15728;
																assign node15728 = (inp[7]) ? 4'b0111 : 4'b0110;
																assign node15731 = (inp[7]) ? 4'b0110 : 4'b0111;
															assign node15734 = (inp[8]) ? 4'b0111 : node15735;
																assign node15735 = (inp[7]) ? 4'b0111 : 4'b0110;
														assign node15739 = (inp[10]) ? 4'b0100 : node15740;
															assign node15740 = (inp[7]) ? node15744 : node15741;
																assign node15741 = (inp[8]) ? 4'b0101 : 4'b0100;
																assign node15744 = (inp[8]) ? 4'b0100 : 4'b0101;
												assign node15748 = (inp[8]) ? node15762 : node15749;
													assign node15749 = (inp[7]) ? node15755 : node15750;
														assign node15750 = (inp[15]) ? 4'b0110 : node15751;
															assign node15751 = (inp[0]) ? 4'b0110 : 4'b0100;
														assign node15755 = (inp[0]) ? node15759 : node15756;
															assign node15756 = (inp[15]) ? 4'b0111 : 4'b0101;
															assign node15759 = (inp[15]) ? 4'b0101 : 4'b0111;
													assign node15762 = (inp[7]) ? node15770 : node15763;
														assign node15763 = (inp[15]) ? node15767 : node15764;
															assign node15764 = (inp[0]) ? 4'b0111 : 4'b0101;
															assign node15767 = (inp[0]) ? 4'b0101 : 4'b0111;
														assign node15770 = (inp[0]) ? node15774 : node15771;
															assign node15771 = (inp[15]) ? 4'b0110 : 4'b0100;
															assign node15774 = (inp[15]) ? 4'b0100 : 4'b0110;
									assign node15777 = (inp[10]) ? node15891 : node15778;
										assign node15778 = (inp[8]) ? node15840 : node15779;
											assign node15779 = (inp[7]) ? node15807 : node15780;
												assign node15780 = (inp[5]) ? node15792 : node15781;
													assign node15781 = (inp[0]) ? 4'b0100 : node15782;
														assign node15782 = (inp[14]) ? node15788 : node15783;
															assign node15783 = (inp[15]) ? node15785 : 4'b0100;
																assign node15785 = (inp[3]) ? 4'b0110 : 4'b0100;
															assign node15788 = (inp[3]) ? 4'b0100 : 4'b0110;
													assign node15792 = (inp[14]) ? node15800 : node15793;
														assign node15793 = (inp[15]) ? node15797 : node15794;
															assign node15794 = (inp[0]) ? 4'b0110 : 4'b0100;
															assign node15797 = (inp[0]) ? 4'b0100 : 4'b0110;
														assign node15800 = (inp[0]) ? node15804 : node15801;
															assign node15801 = (inp[15]) ? 4'b0110 : 4'b0100;
															assign node15804 = (inp[15]) ? 4'b0100 : 4'b0110;
												assign node15807 = (inp[3]) ? node15817 : node15808;
													assign node15808 = (inp[0]) ? 4'b0111 : node15809;
														assign node15809 = (inp[15]) ? node15813 : node15810;
															assign node15810 = (inp[5]) ? 4'b0101 : 4'b0111;
															assign node15813 = (inp[5]) ? 4'b0111 : 4'b0101;
													assign node15817 = (inp[14]) ? node15825 : node15818;
														assign node15818 = (inp[0]) ? node15822 : node15819;
															assign node15819 = (inp[15]) ? 4'b0111 : 4'b0101;
															assign node15822 = (inp[15]) ? 4'b0101 : 4'b0111;
														assign node15825 = (inp[5]) ? node15833 : node15826;
															assign node15826 = (inp[15]) ? node15830 : node15827;
																assign node15827 = (inp[0]) ? 4'b0111 : 4'b0101;
																assign node15830 = (inp[0]) ? 4'b0101 : 4'b0111;
															assign node15833 = (inp[0]) ? node15837 : node15834;
																assign node15834 = (inp[15]) ? 4'b0111 : 4'b0101;
																assign node15837 = (inp[15]) ? 4'b0101 : 4'b0111;
											assign node15840 = (inp[7]) ? node15872 : node15841;
												assign node15841 = (inp[14]) ? node15857 : node15842;
													assign node15842 = (inp[5]) ? node15852 : node15843;
														assign node15843 = (inp[3]) ? node15845 : 4'b0101;
															assign node15845 = (inp[15]) ? node15849 : node15846;
																assign node15846 = (inp[0]) ? 4'b0111 : 4'b0101;
																assign node15849 = (inp[0]) ? 4'b0101 : 4'b0111;
														assign node15852 = (inp[0]) ? 4'b0111 : node15853;
															assign node15853 = (inp[15]) ? 4'b0111 : 4'b0101;
													assign node15857 = (inp[0]) ? node15867 : node15858;
														assign node15858 = (inp[15]) ? node15862 : node15859;
															assign node15859 = (inp[5]) ? 4'b0101 : 4'b0111;
															assign node15862 = (inp[5]) ? 4'b0111 : node15863;
																assign node15863 = (inp[3]) ? 4'b0111 : 4'b0101;
														assign node15867 = (inp[15]) ? node15869 : 4'b0111;
															assign node15869 = (inp[5]) ? 4'b0101 : 4'b0111;
												assign node15872 = (inp[15]) ? node15880 : node15873;
													assign node15873 = (inp[0]) ? 4'b0110 : node15874;
														assign node15874 = (inp[3]) ? 4'b0100 : node15875;
															assign node15875 = (inp[5]) ? 4'b0100 : 4'b0110;
													assign node15880 = (inp[0]) ? node15886 : node15881;
														assign node15881 = (inp[3]) ? 4'b0110 : node15882;
															assign node15882 = (inp[5]) ? 4'b0110 : 4'b0100;
														assign node15886 = (inp[5]) ? 4'b0100 : node15887;
															assign node15887 = (inp[3]) ? 4'b0100 : 4'b0110;
										assign node15891 = (inp[14]) ? node15971 : node15892;
											assign node15892 = (inp[3]) ? node15934 : node15893;
												assign node15893 = (inp[7]) ? node15915 : node15894;
													assign node15894 = (inp[8]) ? node15906 : node15895;
														assign node15895 = (inp[5]) ? node15901 : node15896;
															assign node15896 = (inp[15]) ? node15898 : 4'b0110;
																assign node15898 = (inp[0]) ? 4'b0110 : 4'b0100;
															assign node15901 = (inp[0]) ? 4'b0100 : node15902;
																assign node15902 = (inp[15]) ? 4'b0110 : 4'b0100;
														assign node15906 = (inp[15]) ? 4'b0111 : node15907;
															assign node15907 = (inp[5]) ? node15911 : node15908;
																assign node15908 = (inp[0]) ? 4'b0101 : 4'b0111;
																assign node15911 = (inp[0]) ? 4'b0111 : 4'b0101;
													assign node15915 = (inp[8]) ? node15921 : node15916;
														assign node15916 = (inp[15]) ? node15918 : 4'b0111;
															assign node15918 = (inp[5]) ? 4'b0111 : 4'b0101;
														assign node15921 = (inp[15]) ? node15929 : node15922;
															assign node15922 = (inp[0]) ? node15926 : node15923;
																assign node15923 = (inp[5]) ? 4'b0100 : 4'b0110;
																assign node15926 = (inp[5]) ? 4'b0110 : 4'b0100;
															assign node15929 = (inp[5]) ? 4'b0110 : node15930;
																assign node15930 = (inp[0]) ? 4'b0110 : 4'b0100;
												assign node15934 = (inp[15]) ? node15948 : node15935;
													assign node15935 = (inp[0]) ? node15943 : node15936;
														assign node15936 = (inp[7]) ? node15940 : node15937;
															assign node15937 = (inp[8]) ? 4'b0101 : 4'b0100;
															assign node15940 = (inp[8]) ? 4'b0100 : 4'b0101;
														assign node15943 = (inp[5]) ? 4'b0110 : node15944;
															assign node15944 = (inp[7]) ? 4'b0111 : 4'b0110;
													assign node15948 = (inp[0]) ? node15956 : node15949;
														assign node15949 = (inp[8]) ? node15953 : node15950;
															assign node15950 = (inp[5]) ? 4'b0111 : 4'b0110;
															assign node15953 = (inp[7]) ? 4'b0110 : 4'b0111;
														assign node15956 = (inp[5]) ? node15964 : node15957;
															assign node15957 = (inp[7]) ? node15961 : node15958;
																assign node15958 = (inp[8]) ? 4'b0101 : 4'b0100;
																assign node15961 = (inp[8]) ? 4'b0100 : 4'b0101;
															assign node15964 = (inp[7]) ? node15968 : node15965;
																assign node15965 = (inp[8]) ? 4'b0101 : 4'b0100;
																assign node15968 = (inp[8]) ? 4'b0100 : 4'b0101;
											assign node15971 = (inp[0]) ? node16005 : node15972;
												assign node15972 = (inp[15]) ? node15988 : node15973;
													assign node15973 = (inp[3]) ? node15981 : node15974;
														assign node15974 = (inp[5]) ? node15976 : 4'b0110;
															assign node15976 = (inp[8]) ? 4'b0100 : node15977;
																assign node15977 = (inp[7]) ? 4'b0101 : 4'b0100;
														assign node15981 = (inp[7]) ? node15985 : node15982;
															assign node15982 = (inp[8]) ? 4'b0101 : 4'b0100;
															assign node15985 = (inp[8]) ? 4'b0100 : 4'b0101;
													assign node15988 = (inp[3]) ? node16000 : node15989;
														assign node15989 = (inp[5]) ? node15997 : node15990;
															assign node15990 = (inp[7]) ? node15994 : node15991;
																assign node15991 = (inp[8]) ? 4'b0101 : 4'b0100;
																assign node15994 = (inp[8]) ? 4'b0100 : 4'b0101;
															assign node15997 = (inp[8]) ? 4'b0111 : 4'b0110;
														assign node16000 = (inp[8]) ? node16002 : 4'b0110;
															assign node16002 = (inp[7]) ? 4'b0110 : 4'b0111;
												assign node16005 = (inp[15]) ? node16033 : node16006;
													assign node16006 = (inp[5]) ? node16020 : node16007;
														assign node16007 = (inp[3]) ? node16015 : node16008;
															assign node16008 = (inp[7]) ? node16012 : node16009;
																assign node16009 = (inp[8]) ? 4'b0101 : 4'b0100;
																assign node16012 = (inp[8]) ? 4'b0100 : 4'b0101;
															assign node16015 = (inp[7]) ? node16017 : 4'b0111;
																assign node16017 = (inp[8]) ? 4'b0110 : 4'b0111;
														assign node16020 = (inp[3]) ? node16028 : node16021;
															assign node16021 = (inp[8]) ? node16025 : node16022;
																assign node16022 = (inp[7]) ? 4'b0111 : 4'b0110;
																assign node16025 = (inp[7]) ? 4'b0110 : 4'b0111;
															assign node16028 = (inp[7]) ? node16030 : 4'b0110;
																assign node16030 = (inp[8]) ? 4'b0110 : 4'b0111;
													assign node16033 = (inp[3]) ? node16043 : node16034;
														assign node16034 = (inp[5]) ? node16038 : node16035;
															assign node16035 = (inp[8]) ? 4'b0110 : 4'b0111;
															assign node16038 = (inp[7]) ? 4'b0101 : node16039;
																assign node16039 = (inp[8]) ? 4'b0101 : 4'b0100;
														assign node16043 = (inp[8]) ? node16047 : node16044;
															assign node16044 = (inp[7]) ? 4'b0101 : 4'b0100;
															assign node16047 = (inp[7]) ? 4'b0100 : 4'b0101;
								assign node16050 = (inp[10]) ? node16288 : node16051;
									assign node16051 = (inp[0]) ? node16155 : node16052;
										assign node16052 = (inp[15]) ? node16104 : node16053;
											assign node16053 = (inp[5]) ? node16081 : node16054;
												assign node16054 = (inp[3]) ? node16072 : node16055;
													assign node16055 = (inp[8]) ? node16067 : node16056;
														assign node16056 = (inp[7]) ? node16062 : node16057;
															assign node16057 = (inp[14]) ? 4'b0110 : node16058;
																assign node16058 = (inp[2]) ? 4'b0110 : 4'b0111;
															assign node16062 = (inp[14]) ? 4'b0111 : node16063;
																assign node16063 = (inp[2]) ? 4'b0111 : 4'b0110;
														assign node16067 = (inp[14]) ? 4'b0111 : node16068;
															assign node16068 = (inp[2]) ? 4'b0111 : 4'b0110;
													assign node16072 = (inp[8]) ? node16074 : 4'b0101;
														assign node16074 = (inp[7]) ? 4'b0100 : node16075;
															assign node16075 = (inp[14]) ? 4'b0101 : node16076;
																assign node16076 = (inp[2]) ? 4'b0101 : 4'b0100;
												assign node16081 = (inp[8]) ? node16093 : node16082;
													assign node16082 = (inp[7]) ? node16088 : node16083;
														assign node16083 = (inp[2]) ? 4'b0100 : node16084;
															assign node16084 = (inp[14]) ? 4'b0100 : 4'b0101;
														assign node16088 = (inp[14]) ? 4'b0101 : node16089;
															assign node16089 = (inp[2]) ? 4'b0101 : 4'b0100;
													assign node16093 = (inp[7]) ? node16099 : node16094;
														assign node16094 = (inp[14]) ? 4'b0101 : node16095;
															assign node16095 = (inp[2]) ? 4'b0101 : 4'b0100;
														assign node16099 = (inp[2]) ? 4'b0100 : node16100;
															assign node16100 = (inp[14]) ? 4'b0100 : 4'b0101;
											assign node16104 = (inp[5]) ? node16132 : node16105;
												assign node16105 = (inp[3]) ? node16119 : node16106;
													assign node16106 = (inp[2]) ? node16112 : node16107;
														assign node16107 = (inp[7]) ? 4'b0101 : node16108;
															assign node16108 = (inp[14]) ? 4'b0100 : 4'b0101;
														assign node16112 = (inp[8]) ? node16116 : node16113;
															assign node16113 = (inp[7]) ? 4'b0101 : 4'b0100;
															assign node16116 = (inp[7]) ? 4'b0100 : 4'b0101;
													assign node16119 = (inp[8]) ? node16127 : node16120;
														assign node16120 = (inp[7]) ? 4'b0111 : node16121;
															assign node16121 = (inp[2]) ? 4'b0110 : node16122;
																assign node16122 = (inp[14]) ? 4'b0110 : 4'b0111;
														assign node16127 = (inp[7]) ? 4'b0110 : node16128;
															assign node16128 = (inp[14]) ? 4'b0111 : 4'b0110;
												assign node16132 = (inp[8]) ? node16144 : node16133;
													assign node16133 = (inp[7]) ? node16139 : node16134;
														assign node16134 = (inp[14]) ? 4'b0110 : node16135;
															assign node16135 = (inp[2]) ? 4'b0110 : 4'b0111;
														assign node16139 = (inp[2]) ? 4'b0111 : node16140;
															assign node16140 = (inp[14]) ? 4'b0111 : 4'b0110;
													assign node16144 = (inp[7]) ? node16150 : node16145;
														assign node16145 = (inp[2]) ? 4'b0111 : node16146;
															assign node16146 = (inp[14]) ? 4'b0111 : 4'b0110;
														assign node16150 = (inp[2]) ? 4'b0110 : node16151;
															assign node16151 = (inp[14]) ? 4'b0110 : 4'b0111;
										assign node16155 = (inp[15]) ? node16223 : node16156;
											assign node16156 = (inp[5]) ? node16196 : node16157;
												assign node16157 = (inp[3]) ? node16179 : node16158;
													assign node16158 = (inp[2]) ? node16174 : node16159;
														assign node16159 = (inp[14]) ? node16167 : node16160;
															assign node16160 = (inp[7]) ? node16164 : node16161;
																assign node16161 = (inp[8]) ? 4'b0100 : 4'b0101;
																assign node16164 = (inp[8]) ? 4'b0101 : 4'b0100;
															assign node16167 = (inp[7]) ? node16171 : node16168;
																assign node16168 = (inp[8]) ? 4'b0101 : 4'b0100;
																assign node16171 = (inp[8]) ? 4'b0100 : 4'b0101;
														assign node16174 = (inp[14]) ? 4'b0100 : node16175;
															assign node16175 = (inp[7]) ? 4'b0101 : 4'b0100;
													assign node16179 = (inp[14]) ? node16187 : node16180;
														assign node16180 = (inp[8]) ? 4'b0111 : node16181;
															assign node16181 = (inp[2]) ? 4'b0110 : node16182;
																assign node16182 = (inp[7]) ? 4'b0110 : 4'b0111;
														assign node16187 = (inp[2]) ? node16189 : 4'b0110;
															assign node16189 = (inp[7]) ? node16193 : node16190;
																assign node16190 = (inp[8]) ? 4'b0111 : 4'b0110;
																assign node16193 = (inp[8]) ? 4'b0110 : 4'b0111;
												assign node16196 = (inp[14]) ? node16210 : node16197;
													assign node16197 = (inp[8]) ? node16203 : node16198;
														assign node16198 = (inp[2]) ? 4'b0110 : node16199;
															assign node16199 = (inp[7]) ? 4'b0110 : 4'b0111;
														assign node16203 = (inp[2]) ? node16207 : node16204;
															assign node16204 = (inp[7]) ? 4'b0111 : 4'b0110;
															assign node16207 = (inp[7]) ? 4'b0110 : 4'b0111;
													assign node16210 = (inp[2]) ? node16216 : node16211;
														assign node16211 = (inp[7]) ? node16213 : 4'b0110;
															assign node16213 = (inp[8]) ? 4'b0110 : 4'b0111;
														assign node16216 = (inp[7]) ? node16220 : node16217;
															assign node16217 = (inp[8]) ? 4'b0111 : 4'b0110;
															assign node16220 = (inp[8]) ? 4'b0110 : 4'b0111;
											assign node16223 = (inp[3]) ? node16247 : node16224;
												assign node16224 = (inp[5]) ? node16238 : node16225;
													assign node16225 = (inp[14]) ? node16231 : node16226;
														assign node16226 = (inp[2]) ? node16228 : 4'b0110;
															assign node16228 = (inp[8]) ? 4'b0111 : 4'b0110;
														assign node16231 = (inp[8]) ? node16235 : node16232;
															assign node16232 = (inp[7]) ? 4'b0111 : 4'b0110;
															assign node16235 = (inp[7]) ? 4'b0110 : 4'b0111;
													assign node16238 = (inp[8]) ? node16240 : 4'b0101;
														assign node16240 = (inp[7]) ? node16242 : 4'b0101;
															assign node16242 = (inp[14]) ? 4'b0100 : node16243;
																assign node16243 = (inp[2]) ? 4'b0100 : 4'b0101;
												assign node16247 = (inp[5]) ? node16275 : node16248;
													assign node16248 = (inp[14]) ? node16262 : node16249;
														assign node16249 = (inp[7]) ? node16255 : node16250;
															assign node16250 = (inp[8]) ? node16252 : 4'b0101;
																assign node16252 = (inp[2]) ? 4'b0101 : 4'b0100;
															assign node16255 = (inp[8]) ? node16259 : node16256;
																assign node16256 = (inp[2]) ? 4'b0101 : 4'b0100;
																assign node16259 = (inp[2]) ? 4'b0100 : 4'b0101;
														assign node16262 = (inp[2]) ? node16270 : node16263;
															assign node16263 = (inp[8]) ? node16267 : node16264;
																assign node16264 = (inp[7]) ? 4'b0101 : 4'b0100;
																assign node16267 = (inp[7]) ? 4'b0100 : 4'b0101;
															assign node16270 = (inp[7]) ? node16272 : 4'b0100;
																assign node16272 = (inp[8]) ? 4'b0100 : 4'b0101;
													assign node16275 = (inp[14]) ? node16277 : 4'b0100;
														assign node16277 = (inp[2]) ? node16283 : node16278;
															assign node16278 = (inp[7]) ? node16280 : 4'b0101;
																assign node16280 = (inp[8]) ? 4'b0100 : 4'b0101;
															assign node16283 = (inp[8]) ? node16285 : 4'b0100;
																assign node16285 = (inp[7]) ? 4'b0100 : 4'b0101;
									assign node16288 = (inp[8]) ? node16446 : node16289;
										assign node16289 = (inp[7]) ? node16365 : node16290;
											assign node16290 = (inp[2]) ? node16326 : node16291;
												assign node16291 = (inp[14]) ? node16309 : node16292;
													assign node16292 = (inp[0]) ? node16298 : node16293;
														assign node16293 = (inp[3]) ? node16295 : 4'b0011;
															assign node16295 = (inp[15]) ? 4'b0011 : 4'b0001;
														assign node16298 = (inp[15]) ? node16304 : node16299;
															assign node16299 = (inp[5]) ? 4'b0011 : node16300;
																assign node16300 = (inp[3]) ? 4'b0011 : 4'b0001;
															assign node16304 = (inp[3]) ? 4'b0001 : node16305;
																assign node16305 = (inp[5]) ? 4'b0001 : 4'b0011;
													assign node16309 = (inp[5]) ? node16319 : node16310;
														assign node16310 = (inp[3]) ? node16312 : 4'b0010;
															assign node16312 = (inp[0]) ? node16316 : node16313;
																assign node16313 = (inp[15]) ? 4'b0010 : 4'b0000;
																assign node16316 = (inp[15]) ? 4'b0000 : 4'b0010;
														assign node16319 = (inp[3]) ? 4'b0010 : node16320;
															assign node16320 = (inp[0]) ? node16322 : 4'b0000;
																assign node16322 = (inp[15]) ? 4'b0000 : 4'b0010;
												assign node16326 = (inp[14]) ? node16350 : node16327;
													assign node16327 = (inp[5]) ? node16335 : node16328;
														assign node16328 = (inp[15]) ? node16330 : 4'b0000;
															assign node16330 = (inp[3]) ? node16332 : 4'b0000;
																assign node16332 = (inp[0]) ? 4'b0000 : 4'b0010;
														assign node16335 = (inp[3]) ? node16343 : node16336;
															assign node16336 = (inp[15]) ? node16340 : node16337;
																assign node16337 = (inp[0]) ? 4'b0010 : 4'b0000;
																assign node16340 = (inp[0]) ? 4'b0000 : 4'b0010;
															assign node16343 = (inp[15]) ? node16347 : node16344;
																assign node16344 = (inp[0]) ? 4'b0010 : 4'b0000;
																assign node16347 = (inp[0]) ? 4'b0000 : 4'b0010;
													assign node16350 = (inp[3]) ? node16358 : node16351;
														assign node16351 = (inp[15]) ? node16353 : 4'b0010;
															assign node16353 = (inp[5]) ? node16355 : 4'b0010;
																assign node16355 = (inp[0]) ? 4'b0000 : 4'b0010;
														assign node16358 = (inp[0]) ? node16362 : node16359;
															assign node16359 = (inp[15]) ? 4'b0010 : 4'b0000;
															assign node16362 = (inp[15]) ? 4'b0000 : 4'b0010;
											assign node16365 = (inp[2]) ? node16405 : node16366;
												assign node16366 = (inp[14]) ? node16384 : node16367;
													assign node16367 = (inp[0]) ? node16375 : node16368;
														assign node16368 = (inp[15]) ? node16372 : node16369;
															assign node16369 = (inp[5]) ? 4'b0000 : 4'b0010;
															assign node16372 = (inp[5]) ? 4'b0010 : 4'b0000;
														assign node16375 = (inp[5]) ? 4'b0000 : node16376;
															assign node16376 = (inp[3]) ? node16380 : node16377;
																assign node16377 = (inp[15]) ? 4'b0010 : 4'b0000;
																assign node16380 = (inp[15]) ? 4'b0000 : 4'b0010;
													assign node16384 = (inp[0]) ? node16396 : node16385;
														assign node16385 = (inp[15]) ? node16391 : node16386;
															assign node16386 = (inp[5]) ? 4'b0001 : node16387;
																assign node16387 = (inp[3]) ? 4'b0001 : 4'b0011;
															assign node16391 = (inp[3]) ? 4'b0011 : node16392;
																assign node16392 = (inp[5]) ? 4'b0011 : 4'b0001;
														assign node16396 = (inp[15]) ? node16402 : node16397;
															assign node16397 = (inp[3]) ? 4'b0011 : node16398;
																assign node16398 = (inp[5]) ? 4'b0011 : 4'b0001;
															assign node16402 = (inp[3]) ? 4'b0001 : 4'b0011;
												assign node16405 = (inp[14]) ? node16427 : node16406;
													assign node16406 = (inp[15]) ? node16418 : node16407;
														assign node16407 = (inp[0]) ? node16413 : node16408;
															assign node16408 = (inp[5]) ? 4'b0001 : node16409;
																assign node16409 = (inp[3]) ? 4'b0001 : 4'b0011;
															assign node16413 = (inp[3]) ? 4'b0011 : node16414;
																assign node16414 = (inp[5]) ? 4'b0011 : 4'b0001;
														assign node16418 = (inp[0]) ? node16422 : node16419;
															assign node16419 = (inp[5]) ? 4'b0011 : 4'b0001;
															assign node16422 = (inp[5]) ? 4'b0001 : node16423;
																assign node16423 = (inp[3]) ? 4'b0001 : 4'b0011;
													assign node16427 = (inp[0]) ? node16437 : node16428;
														assign node16428 = (inp[3]) ? node16434 : node16429;
															assign node16429 = (inp[15]) ? node16431 : 4'b0011;
																assign node16431 = (inp[5]) ? 4'b0011 : 4'b0001;
															assign node16434 = (inp[15]) ? 4'b0011 : 4'b0001;
														assign node16437 = (inp[15]) ? node16443 : node16438;
															assign node16438 = (inp[3]) ? 4'b0011 : node16439;
																assign node16439 = (inp[5]) ? 4'b0011 : 4'b0001;
															assign node16443 = (inp[5]) ? 4'b0001 : 4'b0011;
										assign node16446 = (inp[7]) ? node16518 : node16447;
											assign node16447 = (inp[14]) ? node16481 : node16448;
												assign node16448 = (inp[2]) ? node16466 : node16449;
													assign node16449 = (inp[3]) ? node16459 : node16450;
														assign node16450 = (inp[5]) ? node16452 : 4'b0000;
															assign node16452 = (inp[0]) ? node16456 : node16453;
																assign node16453 = (inp[15]) ? 4'b0010 : 4'b0000;
																assign node16456 = (inp[15]) ? 4'b0000 : 4'b0010;
														assign node16459 = (inp[0]) ? node16463 : node16460;
															assign node16460 = (inp[15]) ? 4'b0010 : 4'b0000;
															assign node16463 = (inp[15]) ? 4'b0000 : 4'b0010;
													assign node16466 = (inp[15]) ? node16476 : node16467;
														assign node16467 = (inp[5]) ? node16473 : node16468;
															assign node16468 = (inp[0]) ? 4'b0001 : node16469;
																assign node16469 = (inp[3]) ? 4'b0001 : 4'b0011;
															assign node16473 = (inp[0]) ? 4'b0011 : 4'b0001;
														assign node16476 = (inp[0]) ? 4'b0001 : node16477;
															assign node16477 = (inp[5]) ? 4'b0011 : 4'b0001;
												assign node16481 = (inp[2]) ? node16505 : node16482;
													assign node16482 = (inp[0]) ? node16494 : node16483;
														assign node16483 = (inp[15]) ? node16489 : node16484;
															assign node16484 = (inp[5]) ? 4'b0001 : node16485;
																assign node16485 = (inp[3]) ? 4'b0001 : 4'b0011;
															assign node16489 = (inp[3]) ? 4'b0011 : node16490;
																assign node16490 = (inp[5]) ? 4'b0011 : 4'b0001;
														assign node16494 = (inp[15]) ? node16500 : node16495;
															assign node16495 = (inp[3]) ? 4'b0011 : node16496;
																assign node16496 = (inp[5]) ? 4'b0011 : 4'b0001;
															assign node16500 = (inp[5]) ? 4'b0001 : node16501;
																assign node16501 = (inp[3]) ? 4'b0001 : 4'b0011;
													assign node16505 = (inp[15]) ? node16513 : node16506;
														assign node16506 = (inp[0]) ? node16510 : node16507;
															assign node16507 = (inp[3]) ? 4'b0001 : 4'b0011;
															assign node16510 = (inp[3]) ? 4'b0011 : 4'b0001;
														assign node16513 = (inp[0]) ? 4'b0001 : node16514;
															assign node16514 = (inp[3]) ? 4'b0011 : 4'b0001;
											assign node16518 = (inp[14]) ? node16556 : node16519;
												assign node16519 = (inp[2]) ? node16543 : node16520;
													assign node16520 = (inp[15]) ? node16532 : node16521;
														assign node16521 = (inp[0]) ? node16527 : node16522;
															assign node16522 = (inp[5]) ? 4'b0001 : node16523;
																assign node16523 = (inp[3]) ? 4'b0001 : 4'b0011;
															assign node16527 = (inp[5]) ? 4'b0011 : node16528;
																assign node16528 = (inp[3]) ? 4'b0011 : 4'b0001;
														assign node16532 = (inp[0]) ? node16538 : node16533;
															assign node16533 = (inp[3]) ? 4'b0011 : node16534;
																assign node16534 = (inp[5]) ? 4'b0011 : 4'b0001;
															assign node16538 = (inp[5]) ? 4'b0001 : node16539;
																assign node16539 = (inp[3]) ? 4'b0001 : 4'b0011;
													assign node16543 = (inp[0]) ? node16549 : node16544;
														assign node16544 = (inp[15]) ? node16546 : 4'b0000;
															assign node16546 = (inp[5]) ? 4'b0010 : 4'b0000;
														assign node16549 = (inp[15]) ? 4'b0000 : node16550;
															assign node16550 = (inp[5]) ? 4'b0010 : node16551;
																assign node16551 = (inp[3]) ? 4'b0010 : 4'b0000;
												assign node16556 = (inp[2]) ? node16572 : node16557;
													assign node16557 = (inp[15]) ? node16567 : node16558;
														assign node16558 = (inp[0]) ? node16564 : node16559;
															assign node16559 = (inp[3]) ? 4'b0000 : node16560;
																assign node16560 = (inp[5]) ? 4'b0000 : 4'b0010;
															assign node16564 = (inp[5]) ? 4'b0010 : 4'b0000;
														assign node16567 = (inp[0]) ? 4'b0000 : node16568;
															assign node16568 = (inp[3]) ? 4'b0010 : 4'b0000;
													assign node16572 = (inp[3]) ? node16578 : node16573;
														assign node16573 = (inp[0]) ? node16575 : 4'b0010;
															assign node16575 = (inp[15]) ? 4'b0010 : 4'b0000;
														assign node16578 = (inp[15]) ? node16582 : node16579;
															assign node16579 = (inp[0]) ? 4'b0010 : 4'b0000;
															assign node16582 = (inp[0]) ? 4'b0000 : 4'b0010;
			assign node16585 = (inp[13]) ? node24785 : node16586;
				assign node16586 = (inp[1]) ? node20854 : node16587;
					assign node16587 = (inp[0]) ? node18677 : node16588;
						assign node16588 = (inp[15]) ? node17604 : node16589;
							assign node16589 = (inp[5]) ? node17139 : node16590;
								assign node16590 = (inp[3]) ? node16870 : node16591;
									assign node16591 = (inp[12]) ? node16711 : node16592;
										assign node16592 = (inp[8]) ? node16642 : node16593;
											assign node16593 = (inp[7]) ? node16617 : node16594;
												assign node16594 = (inp[2]) ? node16610 : node16595;
													assign node16595 = (inp[14]) ? node16603 : node16596;
														assign node16596 = (inp[9]) ? node16600 : node16597;
															assign node16597 = (inp[4]) ? 4'b0011 : 4'b0111;
															assign node16600 = (inp[4]) ? 4'b0111 : 4'b0011;
														assign node16603 = (inp[4]) ? node16607 : node16604;
															assign node16604 = (inp[9]) ? 4'b0010 : 4'b0110;
															assign node16607 = (inp[9]) ? 4'b0110 : 4'b0010;
													assign node16610 = (inp[4]) ? node16614 : node16611;
														assign node16611 = (inp[9]) ? 4'b0010 : 4'b0110;
														assign node16614 = (inp[9]) ? 4'b0110 : 4'b0010;
												assign node16617 = (inp[14]) ? node16627 : node16618;
													assign node16618 = (inp[2]) ? node16622 : node16619;
														assign node16619 = (inp[10]) ? 4'b0010 : 4'b0110;
														assign node16622 = (inp[9]) ? node16624 : 4'b0111;
															assign node16624 = (inp[4]) ? 4'b0111 : 4'b0011;
													assign node16627 = (inp[10]) ? node16635 : node16628;
														assign node16628 = (inp[9]) ? node16632 : node16629;
															assign node16629 = (inp[4]) ? 4'b0011 : 4'b0111;
															assign node16632 = (inp[4]) ? 4'b0111 : 4'b0011;
														assign node16635 = (inp[9]) ? node16639 : node16636;
															assign node16636 = (inp[4]) ? 4'b0011 : 4'b0111;
															assign node16639 = (inp[4]) ? 4'b0111 : 4'b0011;
											assign node16642 = (inp[7]) ? node16670 : node16643;
												assign node16643 = (inp[2]) ? node16657 : node16644;
													assign node16644 = (inp[14]) ? node16652 : node16645;
														assign node16645 = (inp[4]) ? node16649 : node16646;
															assign node16646 = (inp[9]) ? 4'b0010 : 4'b0110;
															assign node16649 = (inp[9]) ? 4'b0110 : 4'b0010;
														assign node16652 = (inp[4]) ? node16654 : 4'b0011;
															assign node16654 = (inp[9]) ? 4'b0111 : 4'b0011;
													assign node16657 = (inp[10]) ? node16663 : node16658;
														assign node16658 = (inp[9]) ? node16660 : 4'b0111;
															assign node16660 = (inp[4]) ? 4'b0111 : 4'b0011;
														assign node16663 = (inp[4]) ? node16667 : node16664;
															assign node16664 = (inp[9]) ? 4'b0011 : 4'b0111;
															assign node16667 = (inp[9]) ? 4'b0111 : 4'b0011;
												assign node16670 = (inp[14]) ? node16688 : node16671;
													assign node16671 = (inp[2]) ? node16679 : node16672;
														assign node16672 = (inp[10]) ? node16674 : 4'b0011;
															assign node16674 = (inp[9]) ? 4'b0111 : node16675;
																assign node16675 = (inp[4]) ? 4'b0011 : 4'b0111;
														assign node16679 = (inp[10]) ? 4'b0110 : node16680;
															assign node16680 = (inp[4]) ? node16684 : node16681;
																assign node16681 = (inp[9]) ? 4'b0010 : 4'b0110;
																assign node16684 = (inp[9]) ? 4'b0110 : 4'b0010;
													assign node16688 = (inp[2]) ? node16704 : node16689;
														assign node16689 = (inp[10]) ? node16697 : node16690;
															assign node16690 = (inp[4]) ? node16694 : node16691;
																assign node16691 = (inp[9]) ? 4'b0010 : 4'b0110;
																assign node16694 = (inp[9]) ? 4'b0110 : 4'b0010;
															assign node16697 = (inp[9]) ? node16701 : node16698;
																assign node16698 = (inp[4]) ? 4'b0010 : 4'b0110;
																assign node16701 = (inp[4]) ? 4'b0110 : 4'b0010;
														assign node16704 = (inp[4]) ? node16708 : node16705;
															assign node16705 = (inp[9]) ? 4'b0010 : 4'b0110;
															assign node16708 = (inp[9]) ? 4'b0110 : 4'b0010;
										assign node16711 = (inp[7]) ? node16787 : node16712;
											assign node16712 = (inp[8]) ? node16748 : node16713;
												assign node16713 = (inp[14]) ? node16733 : node16714;
													assign node16714 = (inp[2]) ? node16722 : node16715;
														assign node16715 = (inp[9]) ? node16717 : 4'b0011;
															assign node16717 = (inp[10]) ? node16719 : 4'b0011;
																assign node16719 = (inp[4]) ? 4'b0011 : 4'b0111;
														assign node16722 = (inp[10]) ? node16728 : node16723;
															assign node16723 = (inp[4]) ? node16725 : 4'b0010;
																assign node16725 = (inp[9]) ? 4'b0110 : 4'b0010;
															assign node16728 = (inp[4]) ? node16730 : 4'b0110;
																assign node16730 = (inp[9]) ? 4'b0010 : 4'b0110;
													assign node16733 = (inp[9]) ? node16741 : node16734;
														assign node16734 = (inp[4]) ? node16738 : node16735;
															assign node16735 = (inp[10]) ? 4'b0010 : 4'b0110;
															assign node16738 = (inp[10]) ? 4'b0110 : 4'b0010;
														assign node16741 = (inp[4]) ? node16745 : node16742;
															assign node16742 = (inp[10]) ? 4'b0110 : 4'b0010;
															assign node16745 = (inp[2]) ? 4'b0110 : 4'b0010;
												assign node16748 = (inp[14]) ? node16764 : node16749;
													assign node16749 = (inp[2]) ? node16757 : node16750;
														assign node16750 = (inp[10]) ? 4'b0010 : node16751;
															assign node16751 = (inp[4]) ? 4'b0010 : node16752;
																assign node16752 = (inp[9]) ? 4'b0010 : 4'b0110;
														assign node16757 = (inp[10]) ? node16759 : 4'b0011;
															assign node16759 = (inp[4]) ? node16761 : 4'b0111;
																assign node16761 = (inp[9]) ? 4'b0011 : 4'b0111;
													assign node16764 = (inp[2]) ? node16778 : node16765;
														assign node16765 = (inp[4]) ? node16771 : node16766;
															assign node16766 = (inp[10]) ? node16768 : 4'b0111;
																assign node16768 = (inp[9]) ? 4'b0111 : 4'b0011;
															assign node16771 = (inp[10]) ? node16775 : node16772;
																assign node16772 = (inp[9]) ? 4'b0111 : 4'b0011;
																assign node16775 = (inp[9]) ? 4'b0011 : 4'b0111;
														assign node16778 = (inp[10]) ? 4'b0011 : node16779;
															assign node16779 = (inp[4]) ? node16783 : node16780;
																assign node16780 = (inp[9]) ? 4'b0011 : 4'b0111;
																assign node16783 = (inp[9]) ? 4'b0111 : 4'b0011;
											assign node16787 = (inp[8]) ? node16825 : node16788;
												assign node16788 = (inp[14]) ? node16810 : node16789;
													assign node16789 = (inp[2]) ? node16803 : node16790;
														assign node16790 = (inp[9]) ? node16798 : node16791;
															assign node16791 = (inp[10]) ? node16795 : node16792;
																assign node16792 = (inp[4]) ? 4'b0010 : 4'b0110;
																assign node16795 = (inp[4]) ? 4'b0110 : 4'b0010;
															assign node16798 = (inp[4]) ? node16800 : 4'b0010;
																assign node16800 = (inp[10]) ? 4'b0010 : 4'b0110;
														assign node16803 = (inp[10]) ? 4'b0111 : node16804;
															assign node16804 = (inp[4]) ? 4'b0011 : node16805;
																assign node16805 = (inp[9]) ? 4'b0011 : 4'b0111;
													assign node16810 = (inp[10]) ? node16818 : node16811;
														assign node16811 = (inp[9]) ? node16815 : node16812;
															assign node16812 = (inp[4]) ? 4'b0011 : 4'b0111;
															assign node16815 = (inp[4]) ? 4'b0111 : 4'b0011;
														assign node16818 = (inp[9]) ? node16822 : node16819;
															assign node16819 = (inp[4]) ? 4'b0111 : 4'b0011;
															assign node16822 = (inp[4]) ? 4'b0011 : 4'b0111;
												assign node16825 = (inp[14]) ? node16845 : node16826;
													assign node16826 = (inp[2]) ? node16838 : node16827;
														assign node16827 = (inp[10]) ? node16833 : node16828;
															assign node16828 = (inp[9]) ? 4'b0111 : node16829;
																assign node16829 = (inp[4]) ? 4'b0011 : 4'b0111;
															assign node16833 = (inp[9]) ? node16835 : 4'b0011;
																assign node16835 = (inp[4]) ? 4'b0011 : 4'b0111;
														assign node16838 = (inp[10]) ? 4'b0110 : node16839;
															assign node16839 = (inp[4]) ? node16841 : 4'b0010;
																assign node16841 = (inp[9]) ? 4'b0110 : 4'b0010;
													assign node16845 = (inp[2]) ? node16855 : node16846;
														assign node16846 = (inp[9]) ? node16848 : 4'b0010;
															assign node16848 = (inp[4]) ? node16852 : node16849;
																assign node16849 = (inp[10]) ? 4'b0110 : 4'b0010;
																assign node16852 = (inp[10]) ? 4'b0010 : 4'b0110;
														assign node16855 = (inp[10]) ? node16863 : node16856;
															assign node16856 = (inp[4]) ? node16860 : node16857;
																assign node16857 = (inp[9]) ? 4'b0010 : 4'b0110;
																assign node16860 = (inp[9]) ? 4'b0110 : 4'b0010;
															assign node16863 = (inp[4]) ? node16867 : node16864;
																assign node16864 = (inp[9]) ? 4'b0110 : 4'b0010;
																assign node16867 = (inp[9]) ? 4'b0010 : 4'b0110;
									assign node16870 = (inp[4]) ? node16986 : node16871;
										assign node16871 = (inp[9]) ? node16923 : node16872;
											assign node16872 = (inp[12]) ? node16894 : node16873;
												assign node16873 = (inp[8]) ? node16887 : node16874;
													assign node16874 = (inp[7]) ? node16882 : node16875;
														assign node16875 = (inp[10]) ? 4'b0110 : node16876;
															assign node16876 = (inp[14]) ? 4'b0110 : node16877;
																assign node16877 = (inp[2]) ? 4'b0110 : 4'b0111;
														assign node16882 = (inp[2]) ? 4'b0111 : node16883;
															assign node16883 = (inp[14]) ? 4'b0111 : 4'b0110;
													assign node16887 = (inp[7]) ? 4'b0110 : node16888;
														assign node16888 = (inp[2]) ? 4'b0111 : node16889;
															assign node16889 = (inp[14]) ? 4'b0111 : 4'b0110;
												assign node16894 = (inp[10]) ? node16912 : node16895;
													assign node16895 = (inp[7]) ? node16907 : node16896;
														assign node16896 = (inp[8]) ? node16902 : node16897;
															assign node16897 = (inp[14]) ? 4'b0110 : node16898;
																assign node16898 = (inp[2]) ? 4'b0110 : 4'b0111;
															assign node16902 = (inp[14]) ? 4'b0111 : node16903;
																assign node16903 = (inp[2]) ? 4'b0111 : 4'b0110;
														assign node16907 = (inp[8]) ? 4'b0110 : node16908;
															assign node16908 = (inp[14]) ? 4'b0111 : 4'b0110;
													assign node16912 = (inp[8]) ? node16920 : node16913;
														assign node16913 = (inp[7]) ? node16915 : 4'b0010;
															assign node16915 = (inp[2]) ? 4'b0011 : node16916;
																assign node16916 = (inp[14]) ? 4'b0011 : 4'b0010;
														assign node16920 = (inp[7]) ? 4'b0010 : 4'b0011;
											assign node16923 = (inp[10]) ? node16951 : node16924;
												assign node16924 = (inp[14]) ? node16944 : node16925;
													assign node16925 = (inp[8]) ? node16933 : node16926;
														assign node16926 = (inp[7]) ? node16930 : node16927;
															assign node16927 = (inp[2]) ? 4'b0010 : 4'b0011;
															assign node16930 = (inp[2]) ? 4'b0011 : 4'b0010;
														assign node16933 = (inp[12]) ? node16939 : node16934;
															assign node16934 = (inp[7]) ? node16936 : 4'b0011;
																assign node16936 = (inp[2]) ? 4'b0010 : 4'b0011;
															assign node16939 = (inp[2]) ? 4'b0011 : node16940;
																assign node16940 = (inp[7]) ? 4'b0011 : 4'b0010;
													assign node16944 = (inp[8]) ? node16948 : node16945;
														assign node16945 = (inp[7]) ? 4'b0011 : 4'b0010;
														assign node16948 = (inp[7]) ? 4'b0010 : 4'b0011;
												assign node16951 = (inp[12]) ? node16969 : node16952;
													assign node16952 = (inp[8]) ? node16960 : node16953;
														assign node16953 = (inp[7]) ? node16955 : 4'b0010;
															assign node16955 = (inp[2]) ? 4'b0011 : node16956;
																assign node16956 = (inp[14]) ? 4'b0011 : 4'b0010;
														assign node16960 = (inp[7]) ? node16966 : node16961;
															assign node16961 = (inp[14]) ? 4'b0011 : node16962;
																assign node16962 = (inp[2]) ? 4'b0011 : 4'b0010;
															assign node16966 = (inp[2]) ? 4'b0010 : 4'b0011;
													assign node16969 = (inp[14]) ? node16981 : node16970;
														assign node16970 = (inp[8]) ? node16976 : node16971;
															assign node16971 = (inp[7]) ? node16973 : 4'b0101;
																assign node16973 = (inp[2]) ? 4'b0101 : 4'b0100;
															assign node16976 = (inp[2]) ? 4'b0100 : node16977;
																assign node16977 = (inp[7]) ? 4'b0101 : 4'b0100;
														assign node16981 = (inp[8]) ? 4'b0101 : node16982;
															assign node16982 = (inp[7]) ? 4'b0101 : 4'b0100;
										assign node16986 = (inp[9]) ? node17052 : node16987;
											assign node16987 = (inp[10]) ? node17025 : node16988;
												assign node16988 = (inp[2]) ? node17010 : node16989;
													assign node16989 = (inp[7]) ? node16995 : node16990;
														assign node16990 = (inp[14]) ? node16992 : 4'b0010;
															assign node16992 = (inp[12]) ? 4'b0010 : 4'b0011;
														assign node16995 = (inp[12]) ? node17003 : node16996;
															assign node16996 = (inp[8]) ? node17000 : node16997;
																assign node16997 = (inp[14]) ? 4'b0011 : 4'b0010;
																assign node17000 = (inp[14]) ? 4'b0010 : 4'b0011;
															assign node17003 = (inp[8]) ? node17007 : node17004;
																assign node17004 = (inp[14]) ? 4'b0011 : 4'b0010;
																assign node17007 = (inp[14]) ? 4'b0010 : 4'b0011;
													assign node17010 = (inp[14]) ? node17018 : node17011;
														assign node17011 = (inp[8]) ? node17015 : node17012;
															assign node17012 = (inp[7]) ? 4'b0011 : 4'b0010;
															assign node17015 = (inp[7]) ? 4'b0010 : 4'b0011;
														assign node17018 = (inp[7]) ? node17022 : node17019;
															assign node17019 = (inp[8]) ? 4'b0011 : 4'b0010;
															assign node17022 = (inp[8]) ? 4'b0010 : 4'b0011;
												assign node17025 = (inp[12]) ? node17039 : node17026;
													assign node17026 = (inp[2]) ? node17034 : node17027;
														assign node17027 = (inp[7]) ? 4'b0011 : node17028;
															assign node17028 = (inp[14]) ? node17030 : 4'b0010;
																assign node17030 = (inp[8]) ? 4'b0011 : 4'b0010;
														assign node17034 = (inp[8]) ? node17036 : 4'b0011;
															assign node17036 = (inp[7]) ? 4'b0010 : 4'b0011;
													assign node17039 = (inp[14]) ? node17047 : node17040;
														assign node17040 = (inp[8]) ? node17042 : 4'b0101;
															assign node17042 = (inp[7]) ? node17044 : 4'b0100;
																assign node17044 = (inp[2]) ? 4'b0100 : 4'b0101;
														assign node17047 = (inp[8]) ? node17049 : 4'b0100;
															assign node17049 = (inp[7]) ? 4'b0100 : 4'b0101;
											assign node17052 = (inp[12]) ? node17090 : node17053;
												assign node17053 = (inp[2]) ? node17075 : node17054;
													assign node17054 = (inp[10]) ? node17060 : node17055;
														assign node17055 = (inp[14]) ? 4'b0101 : node17056;
															assign node17056 = (inp[7]) ? 4'b0100 : 4'b0101;
														assign node17060 = (inp[7]) ? node17068 : node17061;
															assign node17061 = (inp[8]) ? node17065 : node17062;
																assign node17062 = (inp[14]) ? 4'b0100 : 4'b0101;
																assign node17065 = (inp[14]) ? 4'b0101 : 4'b0100;
															assign node17068 = (inp[14]) ? node17072 : node17069;
																assign node17069 = (inp[8]) ? 4'b0101 : 4'b0100;
																assign node17072 = (inp[8]) ? 4'b0100 : 4'b0101;
													assign node17075 = (inp[10]) ? node17083 : node17076;
														assign node17076 = (inp[8]) ? node17080 : node17077;
															assign node17077 = (inp[7]) ? 4'b0101 : 4'b0100;
															assign node17080 = (inp[7]) ? 4'b0100 : 4'b0101;
														assign node17083 = (inp[8]) ? node17087 : node17084;
															assign node17084 = (inp[7]) ? 4'b0101 : 4'b0100;
															assign node17087 = (inp[7]) ? 4'b0100 : 4'b0101;
												assign node17090 = (inp[10]) ? node17114 : node17091;
													assign node17091 = (inp[2]) ? node17107 : node17092;
														assign node17092 = (inp[14]) ? node17100 : node17093;
															assign node17093 = (inp[7]) ? node17097 : node17094;
																assign node17094 = (inp[8]) ? 4'b0100 : 4'b0101;
																assign node17097 = (inp[8]) ? 4'b0101 : 4'b0100;
															assign node17100 = (inp[8]) ? node17104 : node17101;
																assign node17101 = (inp[7]) ? 4'b0101 : 4'b0100;
																assign node17104 = (inp[7]) ? 4'b0100 : 4'b0101;
														assign node17107 = (inp[7]) ? node17111 : node17108;
															assign node17108 = (inp[8]) ? 4'b0101 : 4'b0100;
															assign node17111 = (inp[8]) ? 4'b0100 : 4'b0101;
													assign node17114 = (inp[14]) ? node17130 : node17115;
														assign node17115 = (inp[2]) ? node17123 : node17116;
															assign node17116 = (inp[8]) ? node17120 : node17117;
																assign node17117 = (inp[7]) ? 4'b0000 : 4'b0001;
																assign node17120 = (inp[7]) ? 4'b0001 : 4'b0000;
															assign node17123 = (inp[7]) ? node17127 : node17124;
																assign node17124 = (inp[8]) ? 4'b0001 : 4'b0000;
																assign node17127 = (inp[8]) ? 4'b0000 : 4'b0001;
														assign node17130 = (inp[2]) ? node17134 : node17131;
															assign node17131 = (inp[7]) ? 4'b0000 : 4'b0001;
															assign node17134 = (inp[8]) ? 4'b0000 : node17135;
																assign node17135 = (inp[7]) ? 4'b0001 : 4'b0000;
								assign node17139 = (inp[3]) ? node17369 : node17140;
									assign node17140 = (inp[4]) ? node17256 : node17141;
										assign node17141 = (inp[9]) ? node17195 : node17142;
											assign node17142 = (inp[10]) ? node17162 : node17143;
												assign node17143 = (inp[8]) ? node17157 : node17144;
													assign node17144 = (inp[7]) ? node17152 : node17145;
														assign node17145 = (inp[12]) ? 4'b0110 : node17146;
															assign node17146 = (inp[2]) ? 4'b0110 : node17147;
																assign node17147 = (inp[14]) ? 4'b0110 : 4'b0111;
														assign node17152 = (inp[2]) ? 4'b0111 : node17153;
															assign node17153 = (inp[14]) ? 4'b0111 : 4'b0110;
													assign node17157 = (inp[7]) ? node17159 : 4'b0111;
														assign node17159 = (inp[14]) ? 4'b0110 : 4'b0111;
												assign node17162 = (inp[12]) ? node17178 : node17163;
													assign node17163 = (inp[14]) ? node17171 : node17164;
														assign node17164 = (inp[2]) ? node17166 : 4'b0111;
															assign node17166 = (inp[8]) ? 4'b0110 : node17167;
																assign node17167 = (inp[7]) ? 4'b0111 : 4'b0110;
														assign node17171 = (inp[8]) ? node17175 : node17172;
															assign node17172 = (inp[7]) ? 4'b0111 : 4'b0110;
															assign node17175 = (inp[7]) ? 4'b0110 : 4'b0111;
													assign node17178 = (inp[2]) ? node17188 : node17179;
														assign node17179 = (inp[8]) ? node17181 : 4'b0010;
															assign node17181 = (inp[7]) ? node17185 : node17182;
																assign node17182 = (inp[14]) ? 4'b0011 : 4'b0010;
																assign node17185 = (inp[14]) ? 4'b0010 : 4'b0011;
														assign node17188 = (inp[8]) ? node17192 : node17189;
															assign node17189 = (inp[7]) ? 4'b0011 : 4'b0010;
															assign node17192 = (inp[7]) ? 4'b0010 : 4'b0011;
											assign node17195 = (inp[10]) ? node17219 : node17196;
												assign node17196 = (inp[8]) ? node17208 : node17197;
													assign node17197 = (inp[7]) ? node17203 : node17198;
														assign node17198 = (inp[2]) ? 4'b0010 : node17199;
															assign node17199 = (inp[14]) ? 4'b0010 : 4'b0011;
														assign node17203 = (inp[14]) ? 4'b0011 : node17204;
															assign node17204 = (inp[2]) ? 4'b0011 : 4'b0010;
													assign node17208 = (inp[7]) ? node17214 : node17209;
														assign node17209 = (inp[12]) ? node17211 : 4'b0011;
															assign node17211 = (inp[2]) ? 4'b0011 : 4'b0010;
														assign node17214 = (inp[14]) ? 4'b0010 : node17215;
															assign node17215 = (inp[2]) ? 4'b0010 : 4'b0011;
												assign node17219 = (inp[12]) ? node17243 : node17220;
													assign node17220 = (inp[14]) ? node17236 : node17221;
														assign node17221 = (inp[2]) ? node17229 : node17222;
															assign node17222 = (inp[8]) ? node17226 : node17223;
																assign node17223 = (inp[7]) ? 4'b0010 : 4'b0011;
																assign node17226 = (inp[7]) ? 4'b0011 : 4'b0010;
															assign node17229 = (inp[8]) ? node17233 : node17230;
																assign node17230 = (inp[7]) ? 4'b0011 : 4'b0010;
																assign node17233 = (inp[7]) ? 4'b0010 : 4'b0011;
														assign node17236 = (inp[8]) ? node17240 : node17237;
															assign node17237 = (inp[7]) ? 4'b0011 : 4'b0010;
															assign node17240 = (inp[7]) ? 4'b0010 : 4'b0011;
													assign node17243 = (inp[7]) ? node17249 : node17244;
														assign node17244 = (inp[8]) ? 4'b0101 : node17245;
															assign node17245 = (inp[2]) ? 4'b0100 : 4'b0101;
														assign node17249 = (inp[8]) ? 4'b0100 : node17250;
															assign node17250 = (inp[2]) ? 4'b0101 : node17251;
																assign node17251 = (inp[14]) ? 4'b0101 : 4'b0100;
										assign node17256 = (inp[9]) ? node17314 : node17257;
											assign node17257 = (inp[10]) ? node17281 : node17258;
												assign node17258 = (inp[8]) ? node17270 : node17259;
													assign node17259 = (inp[7]) ? node17265 : node17260;
														assign node17260 = (inp[2]) ? 4'b0010 : node17261;
															assign node17261 = (inp[14]) ? 4'b0010 : 4'b0011;
														assign node17265 = (inp[14]) ? 4'b0011 : node17266;
															assign node17266 = (inp[2]) ? 4'b0011 : 4'b0010;
													assign node17270 = (inp[7]) ? node17276 : node17271;
														assign node17271 = (inp[2]) ? 4'b0011 : node17272;
															assign node17272 = (inp[14]) ? 4'b0011 : 4'b0010;
														assign node17276 = (inp[2]) ? 4'b0010 : node17277;
															assign node17277 = (inp[14]) ? 4'b0010 : 4'b0011;
												assign node17281 = (inp[12]) ? node17297 : node17282;
													assign node17282 = (inp[8]) ? node17292 : node17283;
														assign node17283 = (inp[2]) ? 4'b0011 : node17284;
															assign node17284 = (inp[14]) ? node17288 : node17285;
																assign node17285 = (inp[7]) ? 4'b0010 : 4'b0011;
																assign node17288 = (inp[7]) ? 4'b0011 : 4'b0010;
														assign node17292 = (inp[7]) ? 4'b0010 : node17293;
															assign node17293 = (inp[2]) ? 4'b0011 : 4'b0010;
													assign node17297 = (inp[7]) ? node17307 : node17298;
														assign node17298 = (inp[8]) ? node17304 : node17299;
															assign node17299 = (inp[14]) ? 4'b0100 : node17300;
																assign node17300 = (inp[2]) ? 4'b0100 : 4'b0101;
															assign node17304 = (inp[2]) ? 4'b0101 : 4'b0100;
														assign node17307 = (inp[8]) ? node17309 : 4'b0101;
															assign node17309 = (inp[2]) ? 4'b0100 : node17310;
																assign node17310 = (inp[14]) ? 4'b0100 : 4'b0101;
											assign node17314 = (inp[10]) ? node17338 : node17315;
												assign node17315 = (inp[7]) ? node17327 : node17316;
													assign node17316 = (inp[8]) ? node17322 : node17317;
														assign node17317 = (inp[2]) ? 4'b0100 : node17318;
															assign node17318 = (inp[14]) ? 4'b0100 : 4'b0101;
														assign node17322 = (inp[2]) ? 4'b0101 : node17323;
															assign node17323 = (inp[14]) ? 4'b0101 : 4'b0100;
													assign node17327 = (inp[8]) ? node17333 : node17328;
														assign node17328 = (inp[14]) ? 4'b0101 : node17329;
															assign node17329 = (inp[2]) ? 4'b0101 : 4'b0100;
														assign node17333 = (inp[2]) ? 4'b0100 : node17334;
															assign node17334 = (inp[14]) ? 4'b0100 : 4'b0101;
												assign node17338 = (inp[12]) ? node17354 : node17339;
													assign node17339 = (inp[8]) ? node17351 : node17340;
														assign node17340 = (inp[7]) ? node17346 : node17341;
															assign node17341 = (inp[14]) ? 4'b0100 : node17342;
																assign node17342 = (inp[2]) ? 4'b0100 : 4'b0101;
															assign node17346 = (inp[2]) ? 4'b0101 : node17347;
																assign node17347 = (inp[14]) ? 4'b0101 : 4'b0100;
														assign node17351 = (inp[7]) ? 4'b0100 : 4'b0101;
													assign node17354 = (inp[14]) ? node17364 : node17355;
														assign node17355 = (inp[8]) ? node17357 : 4'b0001;
															assign node17357 = (inp[2]) ? node17361 : node17358;
																assign node17358 = (inp[7]) ? 4'b0001 : 4'b0000;
																assign node17361 = (inp[7]) ? 4'b0000 : 4'b0001;
														assign node17364 = (inp[8]) ? 4'b0001 : node17365;
															assign node17365 = (inp[7]) ? 4'b0001 : 4'b0000;
									assign node17369 = (inp[2]) ? node17499 : node17370;
										assign node17370 = (inp[4]) ? node17436 : node17371;
											assign node17371 = (inp[9]) ? node17399 : node17372;
												assign node17372 = (inp[12]) ? node17384 : node17373;
													assign node17373 = (inp[14]) ? 4'b0100 : node17374;
														assign node17374 = (inp[10]) ? node17376 : 4'b0101;
															assign node17376 = (inp[8]) ? node17380 : node17377;
																assign node17377 = (inp[7]) ? 4'b0100 : 4'b0101;
																assign node17380 = (inp[7]) ? 4'b0101 : 4'b0100;
													assign node17384 = (inp[10]) ? node17392 : node17385;
														assign node17385 = (inp[7]) ? node17387 : 4'b0100;
															assign node17387 = (inp[14]) ? 4'b0100 : node17388;
																assign node17388 = (inp[8]) ? 4'b0101 : 4'b0100;
														assign node17392 = (inp[8]) ? 4'b0000 : node17393;
															assign node17393 = (inp[7]) ? node17395 : 4'b0001;
																assign node17395 = (inp[14]) ? 4'b0001 : 4'b0000;
												assign node17399 = (inp[12]) ? node17421 : node17400;
													assign node17400 = (inp[7]) ? node17414 : node17401;
														assign node17401 = (inp[10]) ? node17409 : node17402;
															assign node17402 = (inp[14]) ? node17406 : node17403;
																assign node17403 = (inp[8]) ? 4'b0000 : 4'b0001;
																assign node17406 = (inp[8]) ? 4'b0001 : 4'b0000;
															assign node17409 = (inp[14]) ? node17411 : 4'b0001;
																assign node17411 = (inp[8]) ? 4'b0001 : 4'b0000;
														assign node17414 = (inp[14]) ? node17418 : node17415;
															assign node17415 = (inp[8]) ? 4'b0001 : 4'b0000;
															assign node17418 = (inp[8]) ? 4'b0000 : 4'b0001;
													assign node17421 = (inp[10]) ? node17429 : node17422;
														assign node17422 = (inp[7]) ? node17426 : node17423;
															assign node17423 = (inp[8]) ? 4'b0000 : 4'b0001;
															assign node17426 = (inp[8]) ? 4'b0001 : 4'b0000;
														assign node17429 = (inp[7]) ? 4'b0100 : node17430;
															assign node17430 = (inp[14]) ? node17432 : 4'b0101;
																assign node17432 = (inp[8]) ? 4'b0101 : 4'b0100;
											assign node17436 = (inp[9]) ? node17470 : node17437;
												assign node17437 = (inp[10]) ? node17453 : node17438;
													assign node17438 = (inp[12]) ? node17444 : node17439;
														assign node17439 = (inp[7]) ? node17441 : 4'b0000;
															assign node17441 = (inp[8]) ? 4'b0000 : 4'b0001;
														assign node17444 = (inp[8]) ? node17446 : 4'b0001;
															assign node17446 = (inp[14]) ? node17450 : node17447;
																assign node17447 = (inp[7]) ? 4'b0001 : 4'b0000;
																assign node17450 = (inp[7]) ? 4'b0000 : 4'b0001;
													assign node17453 = (inp[12]) ? node17457 : node17454;
														assign node17454 = (inp[14]) ? 4'b0000 : 4'b0001;
														assign node17457 = (inp[8]) ? node17465 : node17458;
															assign node17458 = (inp[7]) ? node17462 : node17459;
																assign node17459 = (inp[14]) ? 4'b0100 : 4'b0101;
																assign node17462 = (inp[14]) ? 4'b0101 : 4'b0100;
															assign node17465 = (inp[7]) ? 4'b0100 : node17466;
																assign node17466 = (inp[14]) ? 4'b0101 : 4'b0100;
												assign node17470 = (inp[12]) ? node17486 : node17471;
													assign node17471 = (inp[8]) ? node17479 : node17472;
														assign node17472 = (inp[7]) ? node17476 : node17473;
															assign node17473 = (inp[14]) ? 4'b0100 : 4'b0101;
															assign node17476 = (inp[14]) ? 4'b0101 : 4'b0100;
														assign node17479 = (inp[7]) ? node17483 : node17480;
															assign node17480 = (inp[14]) ? 4'b0101 : 4'b0100;
															assign node17483 = (inp[14]) ? 4'b0100 : 4'b0101;
													assign node17486 = (inp[10]) ? node17492 : node17487;
														assign node17487 = (inp[8]) ? 4'b0100 : node17488;
															assign node17488 = (inp[7]) ? 4'b0100 : 4'b0101;
														assign node17492 = (inp[14]) ? node17494 : 4'b0000;
															assign node17494 = (inp[8]) ? node17496 : 4'b0001;
																assign node17496 = (inp[7]) ? 4'b0000 : 4'b0001;
										assign node17499 = (inp[4]) ? node17549 : node17500;
											assign node17500 = (inp[9]) ? node17524 : node17501;
												assign node17501 = (inp[10]) ? node17509 : node17502;
													assign node17502 = (inp[8]) ? node17506 : node17503;
														assign node17503 = (inp[7]) ? 4'b0101 : 4'b0100;
														assign node17506 = (inp[7]) ? 4'b0100 : 4'b0101;
													assign node17509 = (inp[12]) ? node17517 : node17510;
														assign node17510 = (inp[7]) ? node17514 : node17511;
															assign node17511 = (inp[8]) ? 4'b0101 : 4'b0100;
															assign node17514 = (inp[8]) ? 4'b0100 : 4'b0101;
														assign node17517 = (inp[8]) ? node17521 : node17518;
															assign node17518 = (inp[7]) ? 4'b0001 : 4'b0000;
															assign node17521 = (inp[7]) ? 4'b0000 : 4'b0001;
												assign node17524 = (inp[10]) ? node17532 : node17525;
													assign node17525 = (inp[8]) ? node17529 : node17526;
														assign node17526 = (inp[7]) ? 4'b0001 : 4'b0000;
														assign node17529 = (inp[7]) ? 4'b0000 : 4'b0001;
													assign node17532 = (inp[12]) ? node17542 : node17533;
														assign node17533 = (inp[14]) ? 4'b0001 : node17534;
															assign node17534 = (inp[8]) ? node17538 : node17535;
																assign node17535 = (inp[7]) ? 4'b0001 : 4'b0000;
																assign node17538 = (inp[7]) ? 4'b0000 : 4'b0001;
														assign node17542 = (inp[8]) ? node17546 : node17543;
															assign node17543 = (inp[7]) ? 4'b0101 : 4'b0100;
															assign node17546 = (inp[7]) ? 4'b0100 : 4'b0101;
											assign node17549 = (inp[9]) ? node17577 : node17550;
												assign node17550 = (inp[10]) ? node17558 : node17551;
													assign node17551 = (inp[7]) ? node17555 : node17552;
														assign node17552 = (inp[8]) ? 4'b0001 : 4'b0000;
														assign node17555 = (inp[8]) ? 4'b0000 : 4'b0001;
													assign node17558 = (inp[12]) ? node17572 : node17559;
														assign node17559 = (inp[14]) ? node17565 : node17560;
															assign node17560 = (inp[8]) ? 4'b0001 : node17561;
																assign node17561 = (inp[7]) ? 4'b0001 : 4'b0000;
															assign node17565 = (inp[8]) ? node17569 : node17566;
																assign node17566 = (inp[7]) ? 4'b0001 : 4'b0000;
																assign node17569 = (inp[7]) ? 4'b0000 : 4'b0001;
														assign node17572 = (inp[8]) ? node17574 : 4'b0100;
															assign node17574 = (inp[7]) ? 4'b0100 : 4'b0101;
												assign node17577 = (inp[12]) ? node17585 : node17578;
													assign node17578 = (inp[8]) ? node17582 : node17579;
														assign node17579 = (inp[7]) ? 4'b0101 : 4'b0100;
														assign node17582 = (inp[7]) ? 4'b0100 : 4'b0101;
													assign node17585 = (inp[10]) ? node17595 : node17586;
														assign node17586 = (inp[14]) ? 4'b0101 : node17587;
															assign node17587 = (inp[7]) ? node17591 : node17588;
																assign node17588 = (inp[8]) ? 4'b0101 : 4'b0100;
																assign node17591 = (inp[8]) ? 4'b0100 : 4'b0101;
														assign node17595 = (inp[14]) ? node17601 : node17596;
															assign node17596 = (inp[8]) ? 4'b0000 : node17597;
																assign node17597 = (inp[7]) ? 4'b0001 : 4'b0000;
															assign node17601 = (inp[7]) ? 4'b0000 : 4'b0001;
							assign node17604 = (inp[5]) ? node18172 : node17605;
								assign node17605 = (inp[3]) ? node17897 : node17606;
									assign node17606 = (inp[10]) ? node17736 : node17607;
										assign node17607 = (inp[7]) ? node17671 : node17608;
											assign node17608 = (inp[8]) ? node17644 : node17609;
												assign node17609 = (inp[2]) ? node17627 : node17610;
													assign node17610 = (inp[14]) ? node17618 : node17611;
														assign node17611 = (inp[4]) ? node17615 : node17612;
															assign node17612 = (inp[9]) ? 4'b0001 : 4'b0101;
															assign node17615 = (inp[9]) ? 4'b0101 : 4'b0001;
														assign node17618 = (inp[12]) ? node17620 : 4'b0000;
															assign node17620 = (inp[4]) ? node17624 : node17621;
																assign node17621 = (inp[9]) ? 4'b0000 : 4'b0100;
																assign node17624 = (inp[9]) ? 4'b0100 : 4'b0000;
													assign node17627 = (inp[14]) ? node17635 : node17628;
														assign node17628 = (inp[9]) ? node17632 : node17629;
															assign node17629 = (inp[4]) ? 4'b0000 : 4'b0100;
															assign node17632 = (inp[4]) ? 4'b0100 : 4'b0000;
														assign node17635 = (inp[12]) ? node17641 : node17636;
															assign node17636 = (inp[9]) ? node17638 : 4'b0000;
																assign node17638 = (inp[4]) ? 4'b0100 : 4'b0000;
															assign node17641 = (inp[4]) ? 4'b0000 : 4'b0100;
												assign node17644 = (inp[2]) ? node17658 : node17645;
													assign node17645 = (inp[14]) ? node17651 : node17646;
														assign node17646 = (inp[4]) ? 4'b0100 : node17647;
															assign node17647 = (inp[9]) ? 4'b0000 : 4'b0100;
														assign node17651 = (inp[12]) ? 4'b0001 : node17652;
															assign node17652 = (inp[4]) ? 4'b0101 : node17653;
																assign node17653 = (inp[9]) ? 4'b0001 : 4'b0101;
													assign node17658 = (inp[14]) ? node17666 : node17659;
														assign node17659 = (inp[4]) ? node17663 : node17660;
															assign node17660 = (inp[9]) ? 4'b0001 : 4'b0101;
															assign node17663 = (inp[9]) ? 4'b0101 : 4'b0001;
														assign node17666 = (inp[4]) ? 4'b0101 : node17667;
															assign node17667 = (inp[9]) ? 4'b0001 : 4'b0101;
											assign node17671 = (inp[8]) ? node17707 : node17672;
												assign node17672 = (inp[2]) ? node17688 : node17673;
													assign node17673 = (inp[14]) ? node17679 : node17674;
														assign node17674 = (inp[4]) ? 4'b0100 : node17675;
															assign node17675 = (inp[9]) ? 4'b0000 : 4'b0100;
														assign node17679 = (inp[12]) ? 4'b0101 : node17680;
															assign node17680 = (inp[4]) ? node17684 : node17681;
																assign node17681 = (inp[9]) ? 4'b0001 : 4'b0101;
																assign node17684 = (inp[9]) ? 4'b0101 : 4'b0001;
													assign node17688 = (inp[14]) ? node17702 : node17689;
														assign node17689 = (inp[12]) ? node17697 : node17690;
															assign node17690 = (inp[4]) ? node17694 : node17691;
																assign node17691 = (inp[9]) ? 4'b0001 : 4'b0101;
																assign node17694 = (inp[9]) ? 4'b0101 : 4'b0001;
															assign node17697 = (inp[4]) ? 4'b0101 : node17698;
																assign node17698 = (inp[9]) ? 4'b0001 : 4'b0101;
														assign node17702 = (inp[9]) ? 4'b0101 : node17703;
															assign node17703 = (inp[4]) ? 4'b0001 : 4'b0101;
												assign node17707 = (inp[14]) ? node17721 : node17708;
													assign node17708 = (inp[2]) ? node17716 : node17709;
														assign node17709 = (inp[4]) ? node17713 : node17710;
															assign node17710 = (inp[9]) ? 4'b0001 : 4'b0101;
															assign node17713 = (inp[9]) ? 4'b0101 : 4'b0001;
														assign node17716 = (inp[4]) ? node17718 : 4'b0100;
															assign node17718 = (inp[9]) ? 4'b0100 : 4'b0000;
													assign node17721 = (inp[2]) ? node17729 : node17722;
														assign node17722 = (inp[9]) ? node17726 : node17723;
															assign node17723 = (inp[4]) ? 4'b0000 : 4'b0100;
															assign node17726 = (inp[4]) ? 4'b0100 : 4'b0000;
														assign node17729 = (inp[4]) ? node17733 : node17730;
															assign node17730 = (inp[9]) ? 4'b0000 : 4'b0100;
															assign node17733 = (inp[9]) ? 4'b0100 : 4'b0000;
										assign node17736 = (inp[12]) ? node17816 : node17737;
											assign node17737 = (inp[9]) ? node17775 : node17738;
												assign node17738 = (inp[4]) ? node17760 : node17739;
													assign node17739 = (inp[14]) ? node17749 : node17740;
														assign node17740 = (inp[7]) ? node17742 : 4'b0100;
															assign node17742 = (inp[2]) ? node17746 : node17743;
																assign node17743 = (inp[8]) ? 4'b0101 : 4'b0100;
																assign node17746 = (inp[8]) ? 4'b0100 : 4'b0101;
														assign node17749 = (inp[2]) ? node17755 : node17750;
															assign node17750 = (inp[7]) ? 4'b0100 : node17751;
																assign node17751 = (inp[8]) ? 4'b0101 : 4'b0100;
															assign node17755 = (inp[7]) ? node17757 : 4'b0101;
																assign node17757 = (inp[8]) ? 4'b0100 : 4'b0101;
													assign node17760 = (inp[7]) ? node17766 : node17761;
														assign node17761 = (inp[8]) ? 4'b0001 : node17762;
															assign node17762 = (inp[2]) ? 4'b0000 : 4'b0001;
														assign node17766 = (inp[8]) ? node17770 : node17767;
															assign node17767 = (inp[2]) ? 4'b0001 : 4'b0000;
															assign node17770 = (inp[2]) ? 4'b0000 : node17771;
																assign node17771 = (inp[14]) ? 4'b0000 : 4'b0001;
												assign node17775 = (inp[4]) ? node17805 : node17776;
													assign node17776 = (inp[14]) ? node17790 : node17777;
														assign node17777 = (inp[2]) ? node17783 : node17778;
															assign node17778 = (inp[7]) ? 4'b0001 : node17779;
																assign node17779 = (inp[8]) ? 4'b0000 : 4'b0001;
															assign node17783 = (inp[8]) ? node17787 : node17784;
																assign node17784 = (inp[7]) ? 4'b0001 : 4'b0000;
																assign node17787 = (inp[7]) ? 4'b0000 : 4'b0001;
														assign node17790 = (inp[2]) ? node17798 : node17791;
															assign node17791 = (inp[8]) ? node17795 : node17792;
																assign node17792 = (inp[7]) ? 4'b0001 : 4'b0000;
																assign node17795 = (inp[7]) ? 4'b0000 : 4'b0001;
															assign node17798 = (inp[7]) ? node17802 : node17799;
																assign node17799 = (inp[8]) ? 4'b0001 : 4'b0000;
																assign node17802 = (inp[8]) ? 4'b0000 : 4'b0001;
													assign node17805 = (inp[14]) ? 4'b0101 : node17806;
														assign node17806 = (inp[7]) ? node17808 : 4'b0100;
															assign node17808 = (inp[8]) ? node17812 : node17809;
																assign node17809 = (inp[2]) ? 4'b0101 : 4'b0100;
																assign node17812 = (inp[2]) ? 4'b0100 : 4'b0101;
											assign node17816 = (inp[8]) ? node17852 : node17817;
												assign node17817 = (inp[7]) ? node17839 : node17818;
													assign node17818 = (inp[2]) ? node17826 : node17819;
														assign node17819 = (inp[14]) ? 4'b0100 : node17820;
															assign node17820 = (inp[9]) ? node17822 : 4'b0001;
																assign node17822 = (inp[4]) ? 4'b0001 : 4'b0101;
														assign node17826 = (inp[14]) ? node17832 : node17827;
															assign node17827 = (inp[4]) ? 4'b0000 : node17828;
																assign node17828 = (inp[9]) ? 4'b0100 : 4'b0000;
															assign node17832 = (inp[4]) ? node17836 : node17833;
																assign node17833 = (inp[9]) ? 4'b0100 : 4'b0000;
																assign node17836 = (inp[9]) ? 4'b0000 : 4'b0100;
													assign node17839 = (inp[2]) ? node17845 : node17840;
														assign node17840 = (inp[14]) ? 4'b0001 : node17841;
															assign node17841 = (inp[9]) ? 4'b0100 : 4'b0000;
														assign node17845 = (inp[4]) ? node17849 : node17846;
															assign node17846 = (inp[9]) ? 4'b0101 : 4'b0001;
															assign node17849 = (inp[9]) ? 4'b0001 : 4'b0101;
												assign node17852 = (inp[7]) ? node17872 : node17853;
													assign node17853 = (inp[2]) ? node17865 : node17854;
														assign node17854 = (inp[14]) ? node17862 : node17855;
															assign node17855 = (inp[4]) ? node17859 : node17856;
																assign node17856 = (inp[9]) ? 4'b0100 : 4'b0000;
																assign node17859 = (inp[9]) ? 4'b0000 : 4'b0100;
															assign node17862 = (inp[4]) ? 4'b0101 : 4'b0001;
														assign node17865 = (inp[4]) ? node17869 : node17866;
															assign node17866 = (inp[9]) ? 4'b0101 : 4'b0001;
															assign node17869 = (inp[9]) ? 4'b0001 : 4'b0101;
													assign node17872 = (inp[14]) ? node17882 : node17873;
														assign node17873 = (inp[2]) ? node17877 : node17874;
															assign node17874 = (inp[9]) ? 4'b0101 : 4'b0001;
															assign node17877 = (inp[4]) ? 4'b0100 : node17878;
																assign node17878 = (inp[9]) ? 4'b0100 : 4'b0000;
														assign node17882 = (inp[2]) ? node17890 : node17883;
															assign node17883 = (inp[4]) ? node17887 : node17884;
																assign node17884 = (inp[9]) ? 4'b0100 : 4'b0000;
																assign node17887 = (inp[9]) ? 4'b0000 : 4'b0100;
															assign node17890 = (inp[9]) ? node17894 : node17891;
																assign node17891 = (inp[4]) ? 4'b0100 : 4'b0000;
																assign node17894 = (inp[4]) ? 4'b0000 : 4'b0100;
									assign node17897 = (inp[4]) ? node18043 : node17898;
										assign node17898 = (inp[9]) ? node17968 : node17899;
											assign node17899 = (inp[10]) ? node17929 : node17900;
												assign node17900 = (inp[14]) ? node17924 : node17901;
													assign node17901 = (inp[12]) ? node17911 : node17902;
														assign node17902 = (inp[2]) ? node17904 : 4'b0100;
															assign node17904 = (inp[7]) ? node17908 : node17905;
																assign node17905 = (inp[8]) ? 4'b0101 : 4'b0100;
																assign node17908 = (inp[8]) ? 4'b0100 : 4'b0101;
														assign node17911 = (inp[2]) ? node17917 : node17912;
															assign node17912 = (inp[7]) ? 4'b0101 : node17913;
																assign node17913 = (inp[8]) ? 4'b0100 : 4'b0101;
															assign node17917 = (inp[7]) ? node17921 : node17918;
																assign node17918 = (inp[8]) ? 4'b0101 : 4'b0100;
																assign node17921 = (inp[8]) ? 4'b0100 : 4'b0101;
													assign node17924 = (inp[8]) ? 4'b0101 : node17925;
														assign node17925 = (inp[7]) ? 4'b0101 : 4'b0100;
												assign node17929 = (inp[12]) ? node17951 : node17930;
													assign node17930 = (inp[14]) ? node17946 : node17931;
														assign node17931 = (inp[8]) ? node17939 : node17932;
															assign node17932 = (inp[2]) ? node17936 : node17933;
																assign node17933 = (inp[7]) ? 4'b0100 : 4'b0101;
																assign node17936 = (inp[7]) ? 4'b0101 : 4'b0100;
															assign node17939 = (inp[7]) ? node17943 : node17940;
																assign node17940 = (inp[2]) ? 4'b0101 : 4'b0100;
																assign node17943 = (inp[2]) ? 4'b0100 : 4'b0101;
														assign node17946 = (inp[7]) ? 4'b0100 : node17947;
															assign node17947 = (inp[8]) ? 4'b0101 : 4'b0100;
													assign node17951 = (inp[8]) ? node17957 : node17952;
														assign node17952 = (inp[7]) ? node17954 : 4'b0000;
															assign node17954 = (inp[14]) ? 4'b0001 : 4'b0000;
														assign node17957 = (inp[7]) ? node17963 : node17958;
															assign node17958 = (inp[14]) ? 4'b0001 : node17959;
																assign node17959 = (inp[2]) ? 4'b0001 : 4'b0000;
															assign node17963 = (inp[14]) ? 4'b0000 : node17964;
																assign node17964 = (inp[2]) ? 4'b0000 : 4'b0001;
											assign node17968 = (inp[12]) ? node17990 : node17969;
												assign node17969 = (inp[14]) ? node17983 : node17970;
													assign node17970 = (inp[7]) ? node17976 : node17971;
														assign node17971 = (inp[8]) ? 4'b0000 : node17972;
															assign node17972 = (inp[2]) ? 4'b0000 : 4'b0001;
														assign node17976 = (inp[8]) ? node17980 : node17977;
															assign node17977 = (inp[2]) ? 4'b0001 : 4'b0000;
															assign node17980 = (inp[2]) ? 4'b0000 : 4'b0001;
													assign node17983 = (inp[8]) ? node17987 : node17984;
														assign node17984 = (inp[7]) ? 4'b0001 : 4'b0000;
														assign node17987 = (inp[7]) ? 4'b0000 : 4'b0001;
												assign node17990 = (inp[10]) ? node18014 : node17991;
													assign node17991 = (inp[2]) ? node18005 : node17992;
														assign node17992 = (inp[7]) ? node17998 : node17993;
															assign node17993 = (inp[14]) ? node17995 : 4'b0000;
																assign node17995 = (inp[8]) ? 4'b0001 : 4'b0000;
															assign node17998 = (inp[14]) ? node18002 : node17999;
																assign node17999 = (inp[8]) ? 4'b0001 : 4'b0000;
																assign node18002 = (inp[8]) ? 4'b0000 : 4'b0001;
														assign node18005 = (inp[14]) ? 4'b0001 : node18006;
															assign node18006 = (inp[7]) ? node18010 : node18007;
																assign node18007 = (inp[8]) ? 4'b0001 : 4'b0000;
																assign node18010 = (inp[8]) ? 4'b0000 : 4'b0001;
													assign node18014 = (inp[2]) ? node18030 : node18015;
														assign node18015 = (inp[14]) ? node18023 : node18016;
															assign node18016 = (inp[8]) ? node18020 : node18017;
																assign node18017 = (inp[7]) ? 4'b0110 : 4'b0111;
																assign node18020 = (inp[7]) ? 4'b0111 : 4'b0110;
															assign node18023 = (inp[7]) ? node18027 : node18024;
																assign node18024 = (inp[8]) ? 4'b0111 : 4'b0110;
																assign node18027 = (inp[8]) ? 4'b0110 : 4'b0111;
														assign node18030 = (inp[14]) ? node18036 : node18031;
															assign node18031 = (inp[8]) ? node18033 : 4'b0110;
																assign node18033 = (inp[7]) ? 4'b0110 : 4'b0111;
															assign node18036 = (inp[7]) ? node18040 : node18037;
																assign node18037 = (inp[8]) ? 4'b0111 : 4'b0110;
																assign node18040 = (inp[8]) ? 4'b0110 : 4'b0111;
										assign node18043 = (inp[9]) ? node18109 : node18044;
											assign node18044 = (inp[12]) ? node18076 : node18045;
												assign node18045 = (inp[14]) ? node18069 : node18046;
													assign node18046 = (inp[8]) ? node18054 : node18047;
														assign node18047 = (inp[2]) ? node18051 : node18048;
															assign node18048 = (inp[7]) ? 4'b0000 : 4'b0001;
															assign node18051 = (inp[7]) ? 4'b0001 : 4'b0000;
														assign node18054 = (inp[10]) ? node18062 : node18055;
															assign node18055 = (inp[2]) ? node18059 : node18056;
																assign node18056 = (inp[7]) ? 4'b0001 : 4'b0000;
																assign node18059 = (inp[7]) ? 4'b0000 : 4'b0001;
															assign node18062 = (inp[2]) ? node18066 : node18063;
																assign node18063 = (inp[7]) ? 4'b0001 : 4'b0000;
																assign node18066 = (inp[7]) ? 4'b0000 : 4'b0001;
													assign node18069 = (inp[7]) ? node18073 : node18070;
														assign node18070 = (inp[8]) ? 4'b0001 : 4'b0000;
														assign node18073 = (inp[8]) ? 4'b0000 : 4'b0001;
												assign node18076 = (inp[10]) ? node18086 : node18077;
													assign node18077 = (inp[2]) ? 4'b0001 : node18078;
														assign node18078 = (inp[8]) ? node18080 : 4'b0001;
															assign node18080 = (inp[14]) ? 4'b0000 : node18081;
																assign node18081 = (inp[7]) ? 4'b0001 : 4'b0000;
													assign node18086 = (inp[2]) ? node18102 : node18087;
														assign node18087 = (inp[14]) ? node18095 : node18088;
															assign node18088 = (inp[7]) ? node18092 : node18089;
																assign node18089 = (inp[8]) ? 4'b0110 : 4'b0111;
																assign node18092 = (inp[8]) ? 4'b0111 : 4'b0110;
															assign node18095 = (inp[7]) ? node18099 : node18096;
																assign node18096 = (inp[8]) ? 4'b0111 : 4'b0110;
																assign node18099 = (inp[8]) ? 4'b0110 : 4'b0111;
														assign node18102 = (inp[8]) ? node18106 : node18103;
															assign node18103 = (inp[7]) ? 4'b0111 : 4'b0110;
															assign node18106 = (inp[7]) ? 4'b0110 : 4'b0111;
											assign node18109 = (inp[10]) ? node18145 : node18110;
												assign node18110 = (inp[14]) ? node18126 : node18111;
													assign node18111 = (inp[8]) ? node18119 : node18112;
														assign node18112 = (inp[7]) ? node18116 : node18113;
															assign node18113 = (inp[2]) ? 4'b0110 : 4'b0111;
															assign node18116 = (inp[2]) ? 4'b0111 : 4'b0110;
														assign node18119 = (inp[7]) ? node18123 : node18120;
															assign node18120 = (inp[2]) ? 4'b0111 : 4'b0110;
															assign node18123 = (inp[2]) ? 4'b0110 : 4'b0111;
													assign node18126 = (inp[12]) ? node18134 : node18127;
														assign node18127 = (inp[8]) ? node18131 : node18128;
															assign node18128 = (inp[7]) ? 4'b0111 : 4'b0110;
															assign node18131 = (inp[7]) ? 4'b0110 : 4'b0111;
														assign node18134 = (inp[2]) ? node18140 : node18135;
															assign node18135 = (inp[8]) ? node18137 : 4'b0111;
																assign node18137 = (inp[7]) ? 4'b0110 : 4'b0111;
															assign node18140 = (inp[7]) ? 4'b0111 : node18141;
																assign node18141 = (inp[8]) ? 4'b0111 : 4'b0110;
												assign node18145 = (inp[12]) ? node18161 : node18146;
													assign node18146 = (inp[7]) ? node18156 : node18147;
														assign node18147 = (inp[14]) ? 4'b0110 : node18148;
															assign node18148 = (inp[2]) ? node18152 : node18149;
																assign node18149 = (inp[8]) ? 4'b0110 : 4'b0111;
																assign node18152 = (inp[8]) ? 4'b0111 : 4'b0110;
														assign node18156 = (inp[8]) ? node18158 : 4'b0111;
															assign node18158 = (inp[2]) ? 4'b0110 : 4'b0111;
													assign node18161 = (inp[8]) ? node18167 : node18162;
														assign node18162 = (inp[7]) ? 4'b0011 : node18163;
															assign node18163 = (inp[2]) ? 4'b0010 : 4'b0011;
														assign node18167 = (inp[7]) ? 4'b0010 : node18168;
															assign node18168 = (inp[14]) ? 4'b0011 : 4'b0010;
								assign node18172 = (inp[3]) ? node18426 : node18173;
									assign node18173 = (inp[9]) ? node18291 : node18174;
										assign node18174 = (inp[4]) ? node18232 : node18175;
											assign node18175 = (inp[10]) ? node18199 : node18176;
												assign node18176 = (inp[8]) ? node18188 : node18177;
													assign node18177 = (inp[7]) ? node18183 : node18178;
														assign node18178 = (inp[14]) ? 4'b0100 : node18179;
															assign node18179 = (inp[2]) ? 4'b0100 : 4'b0101;
														assign node18183 = (inp[2]) ? 4'b0101 : node18184;
															assign node18184 = (inp[14]) ? 4'b0101 : 4'b0100;
													assign node18188 = (inp[7]) ? node18194 : node18189;
														assign node18189 = (inp[2]) ? 4'b0101 : node18190;
															assign node18190 = (inp[14]) ? 4'b0101 : 4'b0100;
														assign node18194 = (inp[14]) ? 4'b0100 : node18195;
															assign node18195 = (inp[2]) ? 4'b0100 : 4'b0101;
												assign node18199 = (inp[12]) ? node18217 : node18200;
													assign node18200 = (inp[8]) ? node18210 : node18201;
														assign node18201 = (inp[14]) ? 4'b0100 : node18202;
															assign node18202 = (inp[7]) ? node18206 : node18203;
																assign node18203 = (inp[2]) ? 4'b0100 : 4'b0101;
																assign node18206 = (inp[2]) ? 4'b0101 : 4'b0100;
														assign node18210 = (inp[14]) ? 4'b0101 : node18211;
															assign node18211 = (inp[7]) ? 4'b0100 : node18212;
																assign node18212 = (inp[2]) ? 4'b0101 : 4'b0100;
													assign node18217 = (inp[7]) ? node18225 : node18218;
														assign node18218 = (inp[8]) ? 4'b0001 : node18219;
															assign node18219 = (inp[14]) ? 4'b0000 : node18220;
																assign node18220 = (inp[2]) ? 4'b0000 : 4'b0001;
														assign node18225 = (inp[8]) ? 4'b0000 : node18226;
															assign node18226 = (inp[14]) ? 4'b0001 : node18227;
																assign node18227 = (inp[2]) ? 4'b0001 : 4'b0000;
											assign node18232 = (inp[12]) ? node18256 : node18233;
												assign node18233 = (inp[7]) ? node18245 : node18234;
													assign node18234 = (inp[8]) ? node18240 : node18235;
														assign node18235 = (inp[14]) ? 4'b0000 : node18236;
															assign node18236 = (inp[2]) ? 4'b0000 : 4'b0001;
														assign node18240 = (inp[2]) ? 4'b0001 : node18241;
															assign node18241 = (inp[14]) ? 4'b0001 : 4'b0000;
													assign node18245 = (inp[8]) ? node18251 : node18246;
														assign node18246 = (inp[14]) ? 4'b0001 : node18247;
															assign node18247 = (inp[2]) ? 4'b0001 : 4'b0000;
														assign node18251 = (inp[2]) ? 4'b0000 : node18252;
															assign node18252 = (inp[14]) ? 4'b0000 : 4'b0001;
												assign node18256 = (inp[10]) ? node18274 : node18257;
													assign node18257 = (inp[2]) ? node18269 : node18258;
														assign node18258 = (inp[8]) ? node18264 : node18259;
															assign node18259 = (inp[7]) ? 4'b0001 : node18260;
																assign node18260 = (inp[14]) ? 4'b0000 : 4'b0001;
															assign node18264 = (inp[7]) ? 4'b0000 : node18265;
																assign node18265 = (inp[14]) ? 4'b0001 : 4'b0000;
														assign node18269 = (inp[8]) ? 4'b0001 : node18270;
															assign node18270 = (inp[7]) ? 4'b0001 : 4'b0000;
													assign node18274 = (inp[2]) ? node18284 : node18275;
														assign node18275 = (inp[7]) ? node18277 : 4'b0111;
															assign node18277 = (inp[8]) ? node18281 : node18278;
																assign node18278 = (inp[14]) ? 4'b0111 : 4'b0110;
																assign node18281 = (inp[14]) ? 4'b0110 : 4'b0111;
														assign node18284 = (inp[8]) ? node18288 : node18285;
															assign node18285 = (inp[7]) ? 4'b0111 : 4'b0110;
															assign node18288 = (inp[7]) ? 4'b0110 : 4'b0111;
										assign node18291 = (inp[4]) ? node18347 : node18292;
											assign node18292 = (inp[10]) ? node18310 : node18293;
												assign node18293 = (inp[8]) ? node18303 : node18294;
													assign node18294 = (inp[7]) ? node18300 : node18295;
														assign node18295 = (inp[2]) ? 4'b0000 : node18296;
															assign node18296 = (inp[14]) ? 4'b0000 : 4'b0001;
														assign node18300 = (inp[2]) ? 4'b0001 : 4'b0000;
													assign node18303 = (inp[7]) ? node18305 : 4'b0001;
														assign node18305 = (inp[14]) ? 4'b0000 : node18306;
															assign node18306 = (inp[2]) ? 4'b0000 : 4'b0001;
												assign node18310 = (inp[12]) ? node18328 : node18311;
													assign node18311 = (inp[2]) ? node18321 : node18312;
														assign node18312 = (inp[7]) ? 4'b0001 : node18313;
															assign node18313 = (inp[8]) ? node18317 : node18314;
																assign node18314 = (inp[14]) ? 4'b0000 : 4'b0001;
																assign node18317 = (inp[14]) ? 4'b0001 : 4'b0000;
														assign node18321 = (inp[7]) ? node18325 : node18322;
															assign node18322 = (inp[8]) ? 4'b0001 : 4'b0000;
															assign node18325 = (inp[8]) ? 4'b0000 : 4'b0001;
													assign node18328 = (inp[14]) ? node18340 : node18329;
														assign node18329 = (inp[2]) ? node18335 : node18330;
															assign node18330 = (inp[8]) ? node18332 : 4'b0111;
																assign node18332 = (inp[7]) ? 4'b0111 : 4'b0110;
															assign node18335 = (inp[7]) ? node18337 : 4'b0110;
																assign node18337 = (inp[8]) ? 4'b0110 : 4'b0111;
														assign node18340 = (inp[7]) ? node18344 : node18341;
															assign node18341 = (inp[8]) ? 4'b0111 : 4'b0110;
															assign node18344 = (inp[8]) ? 4'b0110 : 4'b0111;
											assign node18347 = (inp[10]) ? node18389 : node18348;
												assign node18348 = (inp[2]) ? node18368 : node18349;
													assign node18349 = (inp[7]) ? node18363 : node18350;
														assign node18350 = (inp[12]) ? node18358 : node18351;
															assign node18351 = (inp[8]) ? node18355 : node18352;
																assign node18352 = (inp[14]) ? 4'b0110 : 4'b0111;
																assign node18355 = (inp[14]) ? 4'b0111 : 4'b0110;
															assign node18358 = (inp[14]) ? node18360 : 4'b0111;
																assign node18360 = (inp[8]) ? 4'b0111 : 4'b0110;
														assign node18363 = (inp[8]) ? 4'b0110 : node18364;
															assign node18364 = (inp[14]) ? 4'b0111 : 4'b0110;
													assign node18368 = (inp[12]) ? node18376 : node18369;
														assign node18369 = (inp[14]) ? node18371 : 4'b0111;
															assign node18371 = (inp[8]) ? node18373 : 4'b0111;
																assign node18373 = (inp[7]) ? 4'b0110 : 4'b0111;
														assign node18376 = (inp[14]) ? node18382 : node18377;
															assign node18377 = (inp[8]) ? 4'b0111 : node18378;
																assign node18378 = (inp[7]) ? 4'b0111 : 4'b0110;
															assign node18382 = (inp[8]) ? node18386 : node18383;
																assign node18383 = (inp[7]) ? 4'b0111 : 4'b0110;
																assign node18386 = (inp[7]) ? 4'b0110 : 4'b0111;
												assign node18389 = (inp[12]) ? node18407 : node18390;
													assign node18390 = (inp[14]) ? node18400 : node18391;
														assign node18391 = (inp[2]) ? node18393 : 4'b0110;
															assign node18393 = (inp[7]) ? node18397 : node18394;
																assign node18394 = (inp[8]) ? 4'b0111 : 4'b0110;
																assign node18397 = (inp[8]) ? 4'b0110 : 4'b0111;
														assign node18400 = (inp[2]) ? 4'b0110 : node18401;
															assign node18401 = (inp[7]) ? 4'b0111 : node18402;
																assign node18402 = (inp[8]) ? 4'b0111 : 4'b0110;
													assign node18407 = (inp[8]) ? node18417 : node18408;
														assign node18408 = (inp[14]) ? 4'b0011 : node18409;
															assign node18409 = (inp[7]) ? node18413 : node18410;
																assign node18410 = (inp[2]) ? 4'b0010 : 4'b0011;
																assign node18413 = (inp[2]) ? 4'b0011 : 4'b0010;
														assign node18417 = (inp[7]) ? node18423 : node18418;
															assign node18418 = (inp[14]) ? 4'b0011 : node18419;
																assign node18419 = (inp[2]) ? 4'b0011 : 4'b0010;
															assign node18423 = (inp[14]) ? 4'b0010 : 4'b0011;
									assign node18426 = (inp[14]) ? node18566 : node18427;
										assign node18427 = (inp[9]) ? node18487 : node18428;
											assign node18428 = (inp[4]) ? node18456 : node18429;
												assign node18429 = (inp[12]) ? node18443 : node18430;
													assign node18430 = (inp[8]) ? node18436 : node18431;
														assign node18431 = (inp[2]) ? 4'b0110 : node18432;
															assign node18432 = (inp[7]) ? 4'b0110 : 4'b0111;
														assign node18436 = (inp[7]) ? node18440 : node18437;
															assign node18437 = (inp[2]) ? 4'b0111 : 4'b0110;
															assign node18440 = (inp[2]) ? 4'b0110 : 4'b0111;
													assign node18443 = (inp[10]) ? node18445 : 4'b0111;
														assign node18445 = (inp[7]) ? node18451 : node18446;
															assign node18446 = (inp[8]) ? node18448 : 4'b0010;
																assign node18448 = (inp[2]) ? 4'b0011 : 4'b0010;
															assign node18451 = (inp[8]) ? node18453 : 4'b0011;
																assign node18453 = (inp[2]) ? 4'b0010 : 4'b0011;
												assign node18456 = (inp[12]) ? node18474 : node18457;
													assign node18457 = (inp[7]) ? node18467 : node18458;
														assign node18458 = (inp[10]) ? node18460 : 4'b0011;
															assign node18460 = (inp[8]) ? node18464 : node18461;
																assign node18461 = (inp[2]) ? 4'b0010 : 4'b0011;
																assign node18464 = (inp[2]) ? 4'b0011 : 4'b0010;
														assign node18467 = (inp[2]) ? node18471 : node18468;
															assign node18468 = (inp[8]) ? 4'b0011 : 4'b0010;
															assign node18471 = (inp[8]) ? 4'b0010 : 4'b0011;
													assign node18474 = (inp[10]) ? node18484 : node18475;
														assign node18475 = (inp[8]) ? node18477 : 4'b0011;
															assign node18477 = (inp[2]) ? node18481 : node18478;
																assign node18478 = (inp[7]) ? 4'b0011 : 4'b0010;
																assign node18481 = (inp[7]) ? 4'b0010 : 4'b0011;
														assign node18484 = (inp[7]) ? 4'b0110 : 4'b0111;
											assign node18487 = (inp[4]) ? node18531 : node18488;
												assign node18488 = (inp[10]) ? node18510 : node18489;
													assign node18489 = (inp[8]) ? node18505 : node18490;
														assign node18490 = (inp[12]) ? node18498 : node18491;
															assign node18491 = (inp[2]) ? node18495 : node18492;
																assign node18492 = (inp[7]) ? 4'b0010 : 4'b0011;
																assign node18495 = (inp[7]) ? 4'b0011 : 4'b0010;
															assign node18498 = (inp[2]) ? node18502 : node18499;
																assign node18499 = (inp[7]) ? 4'b0010 : 4'b0011;
																assign node18502 = (inp[7]) ? 4'b0011 : 4'b0010;
														assign node18505 = (inp[2]) ? 4'b0010 : node18506;
															assign node18506 = (inp[7]) ? 4'b0011 : 4'b0010;
													assign node18510 = (inp[12]) ? node18520 : node18511;
														assign node18511 = (inp[8]) ? 4'b0011 : node18512;
															assign node18512 = (inp[7]) ? node18516 : node18513;
																assign node18513 = (inp[2]) ? 4'b0010 : 4'b0011;
																assign node18516 = (inp[2]) ? 4'b0011 : 4'b0010;
														assign node18520 = (inp[2]) ? node18526 : node18521;
															assign node18521 = (inp[7]) ? node18523 : 4'b0111;
																assign node18523 = (inp[8]) ? 4'b0111 : 4'b0110;
															assign node18526 = (inp[7]) ? node18528 : 4'b0110;
																assign node18528 = (inp[8]) ? 4'b0110 : 4'b0111;
												assign node18531 = (inp[10]) ? node18547 : node18532;
													assign node18532 = (inp[2]) ? node18540 : node18533;
														assign node18533 = (inp[8]) ? node18537 : node18534;
															assign node18534 = (inp[7]) ? 4'b0110 : 4'b0111;
															assign node18537 = (inp[7]) ? 4'b0111 : 4'b0110;
														assign node18540 = (inp[7]) ? node18544 : node18541;
															assign node18541 = (inp[8]) ? 4'b0111 : 4'b0110;
															assign node18544 = (inp[8]) ? 4'b0110 : 4'b0111;
													assign node18547 = (inp[12]) ? node18557 : node18548;
														assign node18548 = (inp[2]) ? node18550 : 4'b0111;
															assign node18550 = (inp[7]) ? node18554 : node18551;
																assign node18551 = (inp[8]) ? 4'b0111 : 4'b0110;
																assign node18554 = (inp[8]) ? 4'b0110 : 4'b0111;
														assign node18557 = (inp[7]) ? 4'b0011 : node18558;
															assign node18558 = (inp[2]) ? node18562 : node18559;
																assign node18559 = (inp[8]) ? 4'b0010 : 4'b0011;
																assign node18562 = (inp[8]) ? 4'b0011 : 4'b0010;
										assign node18566 = (inp[4]) ? node18618 : node18567;
											assign node18567 = (inp[9]) ? node18587 : node18568;
												assign node18568 = (inp[10]) ? node18576 : node18569;
													assign node18569 = (inp[7]) ? node18573 : node18570;
														assign node18570 = (inp[8]) ? 4'b0111 : 4'b0110;
														assign node18573 = (inp[8]) ? 4'b0110 : 4'b0111;
													assign node18576 = (inp[12]) ? node18582 : node18577;
														assign node18577 = (inp[7]) ? node18579 : 4'b0111;
															assign node18579 = (inp[8]) ? 4'b0110 : 4'b0111;
														assign node18582 = (inp[7]) ? node18584 : 4'b0011;
															assign node18584 = (inp[8]) ? 4'b0010 : 4'b0011;
												assign node18587 = (inp[10]) ? node18603 : node18588;
													assign node18588 = (inp[12]) ? node18598 : node18589;
														assign node18589 = (inp[2]) ? node18591 : 4'b0011;
															assign node18591 = (inp[7]) ? node18595 : node18592;
																assign node18592 = (inp[8]) ? 4'b0011 : 4'b0010;
																assign node18595 = (inp[8]) ? 4'b0010 : 4'b0011;
														assign node18598 = (inp[8]) ? 4'b0010 : node18599;
															assign node18599 = (inp[7]) ? 4'b0011 : 4'b0010;
													assign node18603 = (inp[12]) ? node18611 : node18604;
														assign node18604 = (inp[2]) ? 4'b0010 : node18605;
															assign node18605 = (inp[8]) ? node18607 : 4'b0011;
																assign node18607 = (inp[7]) ? 4'b0010 : 4'b0011;
														assign node18611 = (inp[7]) ? node18615 : node18612;
															assign node18612 = (inp[8]) ? 4'b0111 : 4'b0110;
															assign node18615 = (inp[8]) ? 4'b0110 : 4'b0111;
											assign node18618 = (inp[9]) ? node18652 : node18619;
												assign node18619 = (inp[10]) ? node18637 : node18620;
													assign node18620 = (inp[12]) ? node18630 : node18621;
														assign node18621 = (inp[2]) ? node18623 : 4'b0010;
															assign node18623 = (inp[8]) ? node18627 : node18624;
																assign node18624 = (inp[7]) ? 4'b0011 : 4'b0010;
																assign node18627 = (inp[7]) ? 4'b0010 : 4'b0011;
														assign node18630 = (inp[7]) ? node18634 : node18631;
															assign node18631 = (inp[8]) ? 4'b0011 : 4'b0010;
															assign node18634 = (inp[8]) ? 4'b0010 : 4'b0011;
													assign node18637 = (inp[12]) ? node18645 : node18638;
														assign node18638 = (inp[8]) ? node18642 : node18639;
															assign node18639 = (inp[7]) ? 4'b0011 : 4'b0010;
															assign node18642 = (inp[7]) ? 4'b0010 : 4'b0011;
														assign node18645 = (inp[2]) ? 4'b0110 : node18646;
															assign node18646 = (inp[7]) ? node18648 : 4'b0110;
																assign node18648 = (inp[8]) ? 4'b0110 : 4'b0111;
												assign node18652 = (inp[10]) ? node18666 : node18653;
													assign node18653 = (inp[2]) ? node18659 : node18654;
														assign node18654 = (inp[7]) ? 4'b0110 : node18655;
															assign node18655 = (inp[8]) ? 4'b0111 : 4'b0110;
														assign node18659 = (inp[7]) ? node18663 : node18660;
															assign node18660 = (inp[8]) ? 4'b0111 : 4'b0110;
															assign node18663 = (inp[8]) ? 4'b0110 : 4'b0111;
													assign node18666 = (inp[12]) ? node18670 : node18667;
														assign node18667 = (inp[2]) ? 4'b0111 : 4'b0110;
														assign node18670 = (inp[8]) ? node18674 : node18671;
															assign node18671 = (inp[7]) ? 4'b0011 : 4'b0010;
															assign node18674 = (inp[7]) ? 4'b0010 : 4'b0011;
						assign node18677 = (inp[15]) ? node19751 : node18678;
							assign node18678 = (inp[3]) ? node19194 : node18679;
								assign node18679 = (inp[5]) ? node18933 : node18680;
									assign node18680 = (inp[4]) ? node18796 : node18681;
										assign node18681 = (inp[9]) ? node18735 : node18682;
											assign node18682 = (inp[12]) ? node18704 : node18683;
												assign node18683 = (inp[7]) ? node18695 : node18684;
													assign node18684 = (inp[8]) ? node18690 : node18685;
														assign node18685 = (inp[2]) ? 4'b0100 : node18686;
															assign node18686 = (inp[14]) ? 4'b0100 : 4'b0101;
														assign node18690 = (inp[14]) ? 4'b0101 : node18691;
															assign node18691 = (inp[2]) ? 4'b0101 : 4'b0100;
													assign node18695 = (inp[8]) ? node18699 : node18696;
														assign node18696 = (inp[14]) ? 4'b0101 : 4'b0100;
														assign node18699 = (inp[2]) ? 4'b0100 : node18700;
															assign node18700 = (inp[14]) ? 4'b0100 : 4'b0101;
												assign node18704 = (inp[10]) ? node18718 : node18705;
													assign node18705 = (inp[8]) ? node18715 : node18706;
														assign node18706 = (inp[7]) ? node18710 : node18707;
															assign node18707 = (inp[2]) ? 4'b0100 : 4'b0101;
															assign node18710 = (inp[14]) ? 4'b0101 : node18711;
																assign node18711 = (inp[2]) ? 4'b0101 : 4'b0100;
														assign node18715 = (inp[7]) ? 4'b0100 : 4'b0101;
													assign node18718 = (inp[2]) ? node18720 : 4'b0001;
														assign node18720 = (inp[14]) ? node18728 : node18721;
															assign node18721 = (inp[7]) ? node18725 : node18722;
																assign node18722 = (inp[8]) ? 4'b0001 : 4'b0000;
																assign node18725 = (inp[8]) ? 4'b0000 : 4'b0001;
															assign node18728 = (inp[7]) ? node18732 : node18729;
																assign node18729 = (inp[8]) ? 4'b0001 : 4'b0000;
																assign node18732 = (inp[8]) ? 4'b0000 : 4'b0001;
											assign node18735 = (inp[10]) ? node18767 : node18736;
												assign node18736 = (inp[2]) ? node18754 : node18737;
													assign node18737 = (inp[14]) ? node18745 : node18738;
														assign node18738 = (inp[7]) ? node18742 : node18739;
															assign node18739 = (inp[8]) ? 4'b0000 : 4'b0001;
															assign node18742 = (inp[8]) ? 4'b0001 : 4'b0000;
														assign node18745 = (inp[12]) ? node18747 : 4'b0001;
															assign node18747 = (inp[8]) ? node18751 : node18748;
																assign node18748 = (inp[7]) ? 4'b0001 : 4'b0000;
																assign node18751 = (inp[7]) ? 4'b0000 : 4'b0001;
													assign node18754 = (inp[12]) ? node18762 : node18755;
														assign node18755 = (inp[8]) ? node18759 : node18756;
															assign node18756 = (inp[7]) ? 4'b0001 : 4'b0000;
															assign node18759 = (inp[7]) ? 4'b0000 : 4'b0001;
														assign node18762 = (inp[7]) ? node18764 : 4'b0000;
															assign node18764 = (inp[8]) ? 4'b0000 : 4'b0001;
												assign node18767 = (inp[12]) ? node18777 : node18768;
													assign node18768 = (inp[7]) ? node18774 : node18769;
														assign node18769 = (inp[8]) ? node18771 : 4'b0000;
															assign node18771 = (inp[2]) ? 4'b0001 : 4'b0000;
														assign node18774 = (inp[8]) ? 4'b0000 : 4'b0001;
													assign node18777 = (inp[14]) ? node18787 : node18778;
														assign node18778 = (inp[7]) ? 4'b0101 : node18779;
															assign node18779 = (inp[2]) ? node18783 : node18780;
																assign node18780 = (inp[8]) ? 4'b0100 : 4'b0101;
																assign node18783 = (inp[8]) ? 4'b0101 : 4'b0100;
														assign node18787 = (inp[2]) ? 4'b0100 : node18788;
															assign node18788 = (inp[7]) ? node18792 : node18789;
																assign node18789 = (inp[8]) ? 4'b0101 : 4'b0100;
																assign node18792 = (inp[8]) ? 4'b0100 : 4'b0101;
										assign node18796 = (inp[9]) ? node18866 : node18797;
											assign node18797 = (inp[12]) ? node18831 : node18798;
												assign node18798 = (inp[14]) ? node18816 : node18799;
													assign node18799 = (inp[10]) ? node18801 : 4'b0000;
														assign node18801 = (inp[2]) ? node18809 : node18802;
															assign node18802 = (inp[8]) ? node18806 : node18803;
																assign node18803 = (inp[7]) ? 4'b0000 : 4'b0001;
																assign node18806 = (inp[7]) ? 4'b0001 : 4'b0000;
															assign node18809 = (inp[8]) ? node18813 : node18810;
																assign node18810 = (inp[7]) ? 4'b0001 : 4'b0000;
																assign node18813 = (inp[7]) ? 4'b0000 : 4'b0001;
													assign node18816 = (inp[10]) ? node18824 : node18817;
														assign node18817 = (inp[8]) ? node18821 : node18818;
															assign node18818 = (inp[7]) ? 4'b0001 : 4'b0000;
															assign node18821 = (inp[7]) ? 4'b0000 : 4'b0001;
														assign node18824 = (inp[7]) ? node18828 : node18825;
															assign node18825 = (inp[8]) ? 4'b0001 : 4'b0000;
															assign node18828 = (inp[8]) ? 4'b0000 : 4'b0001;
												assign node18831 = (inp[10]) ? node18847 : node18832;
													assign node18832 = (inp[7]) ? node18844 : node18833;
														assign node18833 = (inp[8]) ? node18839 : node18834;
															assign node18834 = (inp[2]) ? 4'b0000 : node18835;
																assign node18835 = (inp[14]) ? 4'b0000 : 4'b0001;
															assign node18839 = (inp[2]) ? 4'b0001 : node18840;
																assign node18840 = (inp[14]) ? 4'b0001 : 4'b0000;
														assign node18844 = (inp[8]) ? 4'b0000 : 4'b0001;
													assign node18847 = (inp[2]) ? node18857 : node18848;
														assign node18848 = (inp[14]) ? 4'b0100 : node18849;
															assign node18849 = (inp[7]) ? node18853 : node18850;
																assign node18850 = (inp[8]) ? 4'b0100 : 4'b0101;
																assign node18853 = (inp[8]) ? 4'b0101 : 4'b0100;
														assign node18857 = (inp[14]) ? 4'b0101 : node18858;
															assign node18858 = (inp[8]) ? node18862 : node18859;
																assign node18859 = (inp[7]) ? 4'b0101 : 4'b0100;
																assign node18862 = (inp[7]) ? 4'b0100 : 4'b0101;
											assign node18866 = (inp[12]) ? node18900 : node18867;
												assign node18867 = (inp[14]) ? node18883 : node18868;
													assign node18868 = (inp[7]) ? 4'b0100 : node18869;
														assign node18869 = (inp[10]) ? node18877 : node18870;
															assign node18870 = (inp[2]) ? node18874 : node18871;
																assign node18871 = (inp[8]) ? 4'b0100 : 4'b0101;
																assign node18874 = (inp[8]) ? 4'b0101 : 4'b0100;
															assign node18877 = (inp[2]) ? node18879 : 4'b0100;
																assign node18879 = (inp[8]) ? 4'b0101 : 4'b0100;
													assign node18883 = (inp[10]) ? node18893 : node18884;
														assign node18884 = (inp[2]) ? 4'b0101 : node18885;
															assign node18885 = (inp[7]) ? node18889 : node18886;
																assign node18886 = (inp[8]) ? 4'b0101 : 4'b0100;
																assign node18889 = (inp[8]) ? 4'b0100 : 4'b0101;
														assign node18893 = (inp[7]) ? node18897 : node18894;
															assign node18894 = (inp[8]) ? 4'b0101 : 4'b0100;
															assign node18897 = (inp[8]) ? 4'b0100 : 4'b0101;
												assign node18900 = (inp[10]) ? node18914 : node18901;
													assign node18901 = (inp[14]) ? node18909 : node18902;
														assign node18902 = (inp[7]) ? 4'b0101 : node18903;
															assign node18903 = (inp[8]) ? 4'b0100 : node18904;
																assign node18904 = (inp[2]) ? 4'b0100 : 4'b0101;
														assign node18909 = (inp[2]) ? node18911 : 4'b0100;
															assign node18911 = (inp[8]) ? 4'b0101 : 4'b0100;
													assign node18914 = (inp[14]) ? node18926 : node18915;
														assign node18915 = (inp[2]) ? node18921 : node18916;
															assign node18916 = (inp[7]) ? node18918 : 4'b0000;
																assign node18918 = (inp[8]) ? 4'b0001 : 4'b0000;
															assign node18921 = (inp[7]) ? node18923 : 4'b0001;
																assign node18923 = (inp[8]) ? 4'b0000 : 4'b0001;
														assign node18926 = (inp[7]) ? node18930 : node18927;
															assign node18927 = (inp[8]) ? 4'b0001 : 4'b0000;
															assign node18930 = (inp[8]) ? 4'b0000 : 4'b0001;
									assign node18933 = (inp[9]) ? node19069 : node18934;
										assign node18934 = (inp[4]) ? node18994 : node18935;
											assign node18935 = (inp[12]) ? node18959 : node18936;
												assign node18936 = (inp[8]) ? node18948 : node18937;
													assign node18937 = (inp[7]) ? node18943 : node18938;
														assign node18938 = (inp[2]) ? 4'b0100 : node18939;
															assign node18939 = (inp[14]) ? 4'b0100 : 4'b0101;
														assign node18943 = (inp[2]) ? 4'b0101 : node18944;
															assign node18944 = (inp[14]) ? 4'b0101 : 4'b0100;
													assign node18948 = (inp[7]) ? node18954 : node18949;
														assign node18949 = (inp[14]) ? 4'b0101 : node18950;
															assign node18950 = (inp[2]) ? 4'b0101 : 4'b0100;
														assign node18954 = (inp[14]) ? 4'b0100 : node18955;
															assign node18955 = (inp[2]) ? 4'b0100 : 4'b0101;
												assign node18959 = (inp[10]) ? node18981 : node18960;
													assign node18960 = (inp[2]) ? node18970 : node18961;
														assign node18961 = (inp[8]) ? 4'b0101 : node18962;
															assign node18962 = (inp[7]) ? node18966 : node18963;
																assign node18963 = (inp[14]) ? 4'b0100 : 4'b0101;
																assign node18966 = (inp[14]) ? 4'b0101 : 4'b0100;
														assign node18970 = (inp[14]) ? node18976 : node18971;
															assign node18971 = (inp[8]) ? 4'b0100 : node18972;
																assign node18972 = (inp[7]) ? 4'b0101 : 4'b0100;
															assign node18976 = (inp[8]) ? node18978 : 4'b0100;
																assign node18978 = (inp[7]) ? 4'b0100 : 4'b0101;
													assign node18981 = (inp[8]) ? node18991 : node18982;
														assign node18982 = (inp[7]) ? node18986 : node18983;
															assign node18983 = (inp[14]) ? 4'b0000 : 4'b0001;
															assign node18986 = (inp[14]) ? 4'b0001 : node18987;
																assign node18987 = (inp[2]) ? 4'b0001 : 4'b0000;
														assign node18991 = (inp[7]) ? 4'b0000 : 4'b0001;
											assign node18994 = (inp[10]) ? node19038 : node18995;
												assign node18995 = (inp[2]) ? node19015 : node18996;
													assign node18996 = (inp[12]) ? node19008 : node18997;
														assign node18997 = (inp[7]) ? node19003 : node18998;
															assign node18998 = (inp[14]) ? 4'b0001 : node18999;
																assign node18999 = (inp[8]) ? 4'b0000 : 4'b0001;
															assign node19003 = (inp[8]) ? node19005 : 4'b0000;
																assign node19005 = (inp[14]) ? 4'b0000 : 4'b0001;
														assign node19008 = (inp[8]) ? node19010 : 4'b0001;
															assign node19010 = (inp[7]) ? node19012 : 4'b0001;
																assign node19012 = (inp[14]) ? 4'b0000 : 4'b0001;
													assign node19015 = (inp[14]) ? node19023 : node19016;
														assign node19016 = (inp[7]) ? node19020 : node19017;
															assign node19017 = (inp[8]) ? 4'b0001 : 4'b0000;
															assign node19020 = (inp[8]) ? 4'b0000 : 4'b0001;
														assign node19023 = (inp[12]) ? node19031 : node19024;
															assign node19024 = (inp[7]) ? node19028 : node19025;
																assign node19025 = (inp[8]) ? 4'b0001 : 4'b0000;
																assign node19028 = (inp[8]) ? 4'b0000 : 4'b0001;
															assign node19031 = (inp[8]) ? node19035 : node19032;
																assign node19032 = (inp[7]) ? 4'b0001 : 4'b0000;
																assign node19035 = (inp[7]) ? 4'b0000 : 4'b0001;
												assign node19038 = (inp[12]) ? node19058 : node19039;
													assign node19039 = (inp[2]) ? node19051 : node19040;
														assign node19040 = (inp[7]) ? node19046 : node19041;
															assign node19041 = (inp[8]) ? 4'b0001 : node19042;
																assign node19042 = (inp[14]) ? 4'b0000 : 4'b0001;
															assign node19046 = (inp[14]) ? node19048 : 4'b0000;
																assign node19048 = (inp[8]) ? 4'b0000 : 4'b0001;
														assign node19051 = (inp[8]) ? node19055 : node19052;
															assign node19052 = (inp[7]) ? 4'b0001 : 4'b0000;
															assign node19055 = (inp[7]) ? 4'b0000 : 4'b0001;
													assign node19058 = (inp[7]) ? node19062 : node19059;
														assign node19059 = (inp[8]) ? 4'b0111 : 4'b0110;
														assign node19062 = (inp[8]) ? 4'b0110 : node19063;
															assign node19063 = (inp[14]) ? 4'b0111 : node19064;
																assign node19064 = (inp[2]) ? 4'b0111 : 4'b0110;
										assign node19069 = (inp[4]) ? node19129 : node19070;
											assign node19070 = (inp[10]) ? node19094 : node19071;
												assign node19071 = (inp[8]) ? node19083 : node19072;
													assign node19072 = (inp[7]) ? node19078 : node19073;
														assign node19073 = (inp[14]) ? 4'b0000 : node19074;
															assign node19074 = (inp[2]) ? 4'b0000 : 4'b0001;
														assign node19078 = (inp[14]) ? 4'b0001 : node19079;
															assign node19079 = (inp[2]) ? 4'b0001 : 4'b0000;
													assign node19083 = (inp[7]) ? node19089 : node19084;
														assign node19084 = (inp[14]) ? 4'b0001 : node19085;
															assign node19085 = (inp[2]) ? 4'b0001 : 4'b0000;
														assign node19089 = (inp[14]) ? 4'b0000 : node19090;
															assign node19090 = (inp[2]) ? 4'b0000 : 4'b0001;
												assign node19094 = (inp[12]) ? node19106 : node19095;
													assign node19095 = (inp[8]) ? node19101 : node19096;
														assign node19096 = (inp[7]) ? 4'b0001 : node19097;
															assign node19097 = (inp[14]) ? 4'b0000 : 4'b0001;
														assign node19101 = (inp[7]) ? node19103 : 4'b0001;
															assign node19103 = (inp[2]) ? 4'b0000 : 4'b0001;
													assign node19106 = (inp[14]) ? node19120 : node19107;
														assign node19107 = (inp[7]) ? node19113 : node19108;
															assign node19108 = (inp[2]) ? 4'b0110 : node19109;
																assign node19109 = (inp[8]) ? 4'b0110 : 4'b0111;
															assign node19113 = (inp[2]) ? node19117 : node19114;
																assign node19114 = (inp[8]) ? 4'b0111 : 4'b0110;
																assign node19117 = (inp[8]) ? 4'b0110 : 4'b0111;
														assign node19120 = (inp[2]) ? node19122 : 4'b0111;
															assign node19122 = (inp[8]) ? node19126 : node19123;
																assign node19123 = (inp[7]) ? 4'b0111 : 4'b0110;
																assign node19126 = (inp[7]) ? 4'b0110 : 4'b0111;
											assign node19129 = (inp[10]) ? node19157 : node19130;
												assign node19130 = (inp[2]) ? node19150 : node19131;
													assign node19131 = (inp[14]) ? node19143 : node19132;
														assign node19132 = (inp[12]) ? node19138 : node19133;
															assign node19133 = (inp[7]) ? 4'b0111 : node19134;
																assign node19134 = (inp[8]) ? 4'b0110 : 4'b0111;
															assign node19138 = (inp[8]) ? 4'b0111 : node19139;
																assign node19139 = (inp[7]) ? 4'b0110 : 4'b0111;
														assign node19143 = (inp[8]) ? node19147 : node19144;
															assign node19144 = (inp[7]) ? 4'b0111 : 4'b0110;
															assign node19147 = (inp[7]) ? 4'b0110 : 4'b0111;
													assign node19150 = (inp[8]) ? node19154 : node19151;
														assign node19151 = (inp[7]) ? 4'b0111 : 4'b0110;
														assign node19154 = (inp[7]) ? 4'b0110 : 4'b0111;
												assign node19157 = (inp[12]) ? node19171 : node19158;
													assign node19158 = (inp[14]) ? node19166 : node19159;
														assign node19159 = (inp[2]) ? node19161 : 4'b0110;
															assign node19161 = (inp[7]) ? 4'b0110 : node19162;
																assign node19162 = (inp[8]) ? 4'b0111 : 4'b0110;
														assign node19166 = (inp[8]) ? 4'b0111 : node19167;
															assign node19167 = (inp[7]) ? 4'b0111 : 4'b0110;
													assign node19171 = (inp[2]) ? node19185 : node19172;
														assign node19172 = (inp[8]) ? node19180 : node19173;
															assign node19173 = (inp[14]) ? node19177 : node19174;
																assign node19174 = (inp[7]) ? 4'b0010 : 4'b0011;
																assign node19177 = (inp[7]) ? 4'b0011 : 4'b0010;
															assign node19180 = (inp[7]) ? 4'b0010 : node19181;
																assign node19181 = (inp[14]) ? 4'b0011 : 4'b0010;
														assign node19185 = (inp[14]) ? 4'b0010 : node19186;
															assign node19186 = (inp[7]) ? node19190 : node19187;
																assign node19187 = (inp[8]) ? 4'b0011 : 4'b0010;
																assign node19190 = (inp[8]) ? 4'b0010 : 4'b0011;
								assign node19194 = (inp[5]) ? node19470 : node19195;
									assign node19195 = (inp[9]) ? node19341 : node19196;
										assign node19196 = (inp[4]) ? node19274 : node19197;
											assign node19197 = (inp[10]) ? node19235 : node19198;
												assign node19198 = (inp[14]) ? node19214 : node19199;
													assign node19199 = (inp[8]) ? node19207 : node19200;
														assign node19200 = (inp[2]) ? node19204 : node19201;
															assign node19201 = (inp[7]) ? 4'b0100 : 4'b0101;
															assign node19204 = (inp[7]) ? 4'b0101 : 4'b0100;
														assign node19207 = (inp[2]) ? node19211 : node19208;
															assign node19208 = (inp[7]) ? 4'b0101 : 4'b0100;
															assign node19211 = (inp[7]) ? 4'b0100 : 4'b0101;
													assign node19214 = (inp[2]) ? node19230 : node19215;
														assign node19215 = (inp[12]) ? node19223 : node19216;
															assign node19216 = (inp[8]) ? node19220 : node19217;
																assign node19217 = (inp[7]) ? 4'b0101 : 4'b0100;
																assign node19220 = (inp[7]) ? 4'b0100 : 4'b0101;
															assign node19223 = (inp[8]) ? node19227 : node19224;
																assign node19224 = (inp[7]) ? 4'b0101 : 4'b0100;
																assign node19227 = (inp[7]) ? 4'b0100 : 4'b0101;
														assign node19230 = (inp[7]) ? node19232 : 4'b0100;
															assign node19232 = (inp[8]) ? 4'b0100 : 4'b0101;
												assign node19235 = (inp[12]) ? node19255 : node19236;
													assign node19236 = (inp[2]) ? node19250 : node19237;
														assign node19237 = (inp[8]) ? node19243 : node19238;
															assign node19238 = (inp[14]) ? node19240 : 4'b0100;
																assign node19240 = (inp[7]) ? 4'b0101 : 4'b0100;
															assign node19243 = (inp[14]) ? node19247 : node19244;
																assign node19244 = (inp[7]) ? 4'b0101 : 4'b0100;
																assign node19247 = (inp[7]) ? 4'b0100 : 4'b0101;
														assign node19250 = (inp[7]) ? node19252 : 4'b0101;
															assign node19252 = (inp[8]) ? 4'b0100 : 4'b0101;
													assign node19255 = (inp[14]) ? node19265 : node19256;
														assign node19256 = (inp[7]) ? node19258 : 4'b0001;
															assign node19258 = (inp[8]) ? node19262 : node19259;
																assign node19259 = (inp[2]) ? 4'b0001 : 4'b0000;
																assign node19262 = (inp[2]) ? 4'b0000 : 4'b0001;
														assign node19265 = (inp[2]) ? node19267 : 4'b0000;
															assign node19267 = (inp[7]) ? node19271 : node19268;
																assign node19268 = (inp[8]) ? 4'b0001 : 4'b0000;
																assign node19271 = (inp[8]) ? 4'b0000 : 4'b0001;
											assign node19274 = (inp[10]) ? node19312 : node19275;
												assign node19275 = (inp[12]) ? node19297 : node19276;
													assign node19276 = (inp[2]) ? node19290 : node19277;
														assign node19277 = (inp[14]) ? node19285 : node19278;
															assign node19278 = (inp[7]) ? node19282 : node19279;
																assign node19279 = (inp[8]) ? 4'b0000 : 4'b0001;
																assign node19282 = (inp[8]) ? 4'b0001 : 4'b0000;
															assign node19285 = (inp[7]) ? node19287 : 4'b0001;
																assign node19287 = (inp[8]) ? 4'b0000 : 4'b0001;
														assign node19290 = (inp[8]) ? node19294 : node19291;
															assign node19291 = (inp[7]) ? 4'b0001 : 4'b0000;
															assign node19294 = (inp[7]) ? 4'b0000 : 4'b0001;
													assign node19297 = (inp[2]) ? 4'b0001 : node19298;
														assign node19298 = (inp[7]) ? node19306 : node19299;
															assign node19299 = (inp[8]) ? node19303 : node19300;
																assign node19300 = (inp[14]) ? 4'b0000 : 4'b0001;
																assign node19303 = (inp[14]) ? 4'b0001 : 4'b0000;
															assign node19306 = (inp[14]) ? node19308 : 4'b0001;
																assign node19308 = (inp[8]) ? 4'b0000 : 4'b0001;
												assign node19312 = (inp[12]) ? node19326 : node19313;
													assign node19313 = (inp[7]) ? node19317 : node19314;
														assign node19314 = (inp[2]) ? 4'b0000 : 4'b0001;
														assign node19317 = (inp[8]) ? node19321 : node19318;
															assign node19318 = (inp[2]) ? 4'b0001 : 4'b0000;
															assign node19321 = (inp[2]) ? 4'b0000 : node19322;
																assign node19322 = (inp[14]) ? 4'b0000 : 4'b0001;
													assign node19326 = (inp[14]) ? node19334 : node19327;
														assign node19327 = (inp[7]) ? node19329 : 4'b0111;
															assign node19329 = (inp[2]) ? node19331 : 4'b0110;
																assign node19331 = (inp[8]) ? 4'b0110 : 4'b0111;
														assign node19334 = (inp[2]) ? 4'b0110 : node19335;
															assign node19335 = (inp[8]) ? node19337 : 4'b0110;
																assign node19337 = (inp[7]) ? 4'b0110 : 4'b0111;
										assign node19341 = (inp[4]) ? node19397 : node19342;
											assign node19342 = (inp[12]) ? node19366 : node19343;
												assign node19343 = (inp[14]) ? node19359 : node19344;
													assign node19344 = (inp[2]) ? node19352 : node19345;
														assign node19345 = (inp[8]) ? node19349 : node19346;
															assign node19346 = (inp[7]) ? 4'b0000 : 4'b0001;
															assign node19349 = (inp[7]) ? 4'b0001 : 4'b0000;
														assign node19352 = (inp[7]) ? node19356 : node19353;
															assign node19353 = (inp[8]) ? 4'b0001 : 4'b0000;
															assign node19356 = (inp[8]) ? 4'b0000 : 4'b0001;
													assign node19359 = (inp[8]) ? node19363 : node19360;
														assign node19360 = (inp[7]) ? 4'b0001 : 4'b0000;
														assign node19363 = (inp[7]) ? 4'b0000 : 4'b0001;
												assign node19366 = (inp[10]) ? node19378 : node19367;
													assign node19367 = (inp[8]) ? node19373 : node19368;
														assign node19368 = (inp[7]) ? 4'b0001 : node19369;
															assign node19369 = (inp[2]) ? 4'b0000 : 4'b0001;
														assign node19373 = (inp[7]) ? 4'b0000 : node19374;
															assign node19374 = (inp[2]) ? 4'b0001 : 4'b0000;
													assign node19378 = (inp[14]) ? node19390 : node19379;
														assign node19379 = (inp[2]) ? node19385 : node19380;
															assign node19380 = (inp[8]) ? 4'b0110 : node19381;
																assign node19381 = (inp[7]) ? 4'b0110 : 4'b0111;
															assign node19385 = (inp[8]) ? 4'b0111 : node19386;
																assign node19386 = (inp[7]) ? 4'b0111 : 4'b0110;
														assign node19390 = (inp[8]) ? node19394 : node19391;
															assign node19391 = (inp[7]) ? 4'b0111 : 4'b0110;
															assign node19394 = (inp[7]) ? 4'b0110 : 4'b0111;
											assign node19397 = (inp[12]) ? node19433 : node19398;
												assign node19398 = (inp[10]) ? node19410 : node19399;
													assign node19399 = (inp[7]) ? node19405 : node19400;
														assign node19400 = (inp[8]) ? 4'b0111 : node19401;
															assign node19401 = (inp[14]) ? 4'b0110 : 4'b0111;
														assign node19405 = (inp[8]) ? 4'b0110 : node19406;
															assign node19406 = (inp[2]) ? 4'b0111 : 4'b0110;
													assign node19410 = (inp[14]) ? node19426 : node19411;
														assign node19411 = (inp[2]) ? node19419 : node19412;
															assign node19412 = (inp[7]) ? node19416 : node19413;
																assign node19413 = (inp[8]) ? 4'b0110 : 4'b0111;
																assign node19416 = (inp[8]) ? 4'b0111 : 4'b0110;
															assign node19419 = (inp[7]) ? node19423 : node19420;
																assign node19420 = (inp[8]) ? 4'b0111 : 4'b0110;
																assign node19423 = (inp[8]) ? 4'b0110 : 4'b0111;
														assign node19426 = (inp[8]) ? node19430 : node19427;
															assign node19427 = (inp[7]) ? 4'b0111 : 4'b0110;
															assign node19430 = (inp[7]) ? 4'b0110 : 4'b0111;
												assign node19433 = (inp[10]) ? node19453 : node19434;
													assign node19434 = (inp[8]) ? node19444 : node19435;
														assign node19435 = (inp[7]) ? node19441 : node19436;
															assign node19436 = (inp[14]) ? 4'b0110 : node19437;
																assign node19437 = (inp[2]) ? 4'b0110 : 4'b0111;
															assign node19441 = (inp[2]) ? 4'b0111 : 4'b0110;
														assign node19444 = (inp[7]) ? node19450 : node19445;
															assign node19445 = (inp[14]) ? 4'b0111 : node19446;
																assign node19446 = (inp[2]) ? 4'b0111 : 4'b0110;
															assign node19450 = (inp[2]) ? 4'b0110 : 4'b0111;
													assign node19453 = (inp[7]) ? node19459 : node19454;
														assign node19454 = (inp[8]) ? 4'b0011 : node19455;
															assign node19455 = (inp[2]) ? 4'b0010 : 4'b0011;
														assign node19459 = (inp[8]) ? node19465 : node19460;
															assign node19460 = (inp[2]) ? 4'b0011 : node19461;
																assign node19461 = (inp[14]) ? 4'b0011 : 4'b0010;
															assign node19465 = (inp[14]) ? 4'b0010 : node19466;
																assign node19466 = (inp[2]) ? 4'b0010 : 4'b0011;
									assign node19470 = (inp[8]) ? node19588 : node19471;
										assign node19471 = (inp[7]) ? node19529 : node19472;
											assign node19472 = (inp[14]) ? node19508 : node19473;
												assign node19473 = (inp[2]) ? node19491 : node19474;
													assign node19474 = (inp[4]) ? node19484 : node19475;
														assign node19475 = (inp[9]) ? node19481 : node19476;
															assign node19476 = (inp[10]) ? node19478 : 4'b0111;
																assign node19478 = (inp[12]) ? 4'b0011 : 4'b0111;
															assign node19481 = (inp[12]) ? 4'b0111 : 4'b0011;
														assign node19484 = (inp[9]) ? node19486 : 4'b0011;
															assign node19486 = (inp[10]) ? node19488 : 4'b0111;
																assign node19488 = (inp[12]) ? 4'b0011 : 4'b0111;
													assign node19491 = (inp[12]) ? node19499 : node19492;
														assign node19492 = (inp[4]) ? node19496 : node19493;
															assign node19493 = (inp[9]) ? 4'b0010 : 4'b0110;
															assign node19496 = (inp[9]) ? 4'b0110 : 4'b0010;
														assign node19499 = (inp[4]) ? node19501 : 4'b0110;
															assign node19501 = (inp[10]) ? node19505 : node19502;
																assign node19502 = (inp[9]) ? 4'b0110 : 4'b0010;
																assign node19505 = (inp[9]) ? 4'b0010 : 4'b0110;
												assign node19508 = (inp[4]) ? node19518 : node19509;
													assign node19509 = (inp[9]) ? node19513 : node19510;
														assign node19510 = (inp[12]) ? 4'b0010 : 4'b0110;
														assign node19513 = (inp[12]) ? node19515 : 4'b0010;
															assign node19515 = (inp[10]) ? 4'b0110 : 4'b0010;
													assign node19518 = (inp[9]) ? node19524 : node19519;
														assign node19519 = (inp[10]) ? node19521 : 4'b0010;
															assign node19521 = (inp[12]) ? 4'b0110 : 4'b0010;
														assign node19524 = (inp[12]) ? node19526 : 4'b0110;
															assign node19526 = (inp[10]) ? 4'b0010 : 4'b0110;
											assign node19529 = (inp[2]) ? node19569 : node19530;
												assign node19530 = (inp[14]) ? node19552 : node19531;
													assign node19531 = (inp[12]) ? node19539 : node19532;
														assign node19532 = (inp[9]) ? node19536 : node19533;
															assign node19533 = (inp[4]) ? 4'b0010 : 4'b0110;
															assign node19536 = (inp[4]) ? 4'b0110 : 4'b0010;
														assign node19539 = (inp[9]) ? node19545 : node19540;
															assign node19540 = (inp[4]) ? node19542 : 4'b0110;
																assign node19542 = (inp[10]) ? 4'b0110 : 4'b0010;
															assign node19545 = (inp[4]) ? node19549 : node19546;
																assign node19546 = (inp[10]) ? 4'b0110 : 4'b0010;
																assign node19549 = (inp[10]) ? 4'b0010 : 4'b0110;
													assign node19552 = (inp[4]) ? node19562 : node19553;
														assign node19553 = (inp[9]) ? node19559 : node19554;
															assign node19554 = (inp[10]) ? node19556 : 4'b0111;
																assign node19556 = (inp[12]) ? 4'b0011 : 4'b0111;
															assign node19559 = (inp[10]) ? 4'b0111 : 4'b0011;
														assign node19562 = (inp[9]) ? node19564 : 4'b0011;
															assign node19564 = (inp[12]) ? node19566 : 4'b0111;
																assign node19566 = (inp[10]) ? 4'b0011 : 4'b0111;
												assign node19569 = (inp[4]) ? node19581 : node19570;
													assign node19570 = (inp[9]) ? node19576 : node19571;
														assign node19571 = (inp[12]) ? node19573 : 4'b0111;
															assign node19573 = (inp[10]) ? 4'b0011 : 4'b0111;
														assign node19576 = (inp[10]) ? node19578 : 4'b0011;
															assign node19578 = (inp[12]) ? 4'b0111 : 4'b0011;
													assign node19581 = (inp[9]) ? node19583 : 4'b0011;
														assign node19583 = (inp[10]) ? node19585 : 4'b0111;
															assign node19585 = (inp[12]) ? 4'b0011 : 4'b0111;
										assign node19588 = (inp[7]) ? node19662 : node19589;
											assign node19589 = (inp[14]) ? node19627 : node19590;
												assign node19590 = (inp[2]) ? node19608 : node19591;
													assign node19591 = (inp[12]) ? node19599 : node19592;
														assign node19592 = (inp[4]) ? node19596 : node19593;
															assign node19593 = (inp[9]) ? 4'b0010 : 4'b0110;
															assign node19596 = (inp[9]) ? 4'b0110 : 4'b0010;
														assign node19599 = (inp[4]) ? 4'b0110 : node19600;
															assign node19600 = (inp[9]) ? node19604 : node19601;
																assign node19601 = (inp[10]) ? 4'b0010 : 4'b0110;
																assign node19604 = (inp[10]) ? 4'b0110 : 4'b0010;
													assign node19608 = (inp[4]) ? node19616 : node19609;
														assign node19609 = (inp[9]) ? node19611 : 4'b0111;
															assign node19611 = (inp[10]) ? node19613 : 4'b0011;
																assign node19613 = (inp[12]) ? 4'b0111 : 4'b0011;
														assign node19616 = (inp[9]) ? node19622 : node19617;
															assign node19617 = (inp[12]) ? node19619 : 4'b0011;
																assign node19619 = (inp[10]) ? 4'b0111 : 4'b0011;
															assign node19622 = (inp[12]) ? node19624 : 4'b0111;
																assign node19624 = (inp[10]) ? 4'b0011 : 4'b0111;
												assign node19627 = (inp[12]) ? node19647 : node19628;
													assign node19628 = (inp[2]) ? node19636 : node19629;
														assign node19629 = (inp[4]) ? node19633 : node19630;
															assign node19630 = (inp[9]) ? 4'b0011 : 4'b0111;
															assign node19633 = (inp[9]) ? 4'b0111 : 4'b0011;
														assign node19636 = (inp[10]) ? node19642 : node19637;
															assign node19637 = (inp[9]) ? node19639 : 4'b0111;
																assign node19639 = (inp[4]) ? 4'b0111 : 4'b0011;
															assign node19642 = (inp[4]) ? node19644 : 4'b0111;
																assign node19644 = (inp[9]) ? 4'b0111 : 4'b0011;
													assign node19647 = (inp[10]) ? node19655 : node19648;
														assign node19648 = (inp[9]) ? node19652 : node19649;
															assign node19649 = (inp[4]) ? 4'b0011 : 4'b0111;
															assign node19652 = (inp[4]) ? 4'b0111 : 4'b0011;
														assign node19655 = (inp[9]) ? node19659 : node19656;
															assign node19656 = (inp[4]) ? 4'b0111 : 4'b0011;
															assign node19659 = (inp[4]) ? 4'b0011 : 4'b0111;
											assign node19662 = (inp[2]) ? node19708 : node19663;
												assign node19663 = (inp[14]) ? node19683 : node19664;
													assign node19664 = (inp[4]) ? node19674 : node19665;
														assign node19665 = (inp[12]) ? node19667 : 4'b0111;
															assign node19667 = (inp[9]) ? node19671 : node19668;
																assign node19668 = (inp[10]) ? 4'b0011 : 4'b0111;
																assign node19671 = (inp[10]) ? 4'b0111 : 4'b0011;
														assign node19674 = (inp[9]) ? node19678 : node19675;
															assign node19675 = (inp[12]) ? 4'b0111 : 4'b0011;
															assign node19678 = (inp[10]) ? node19680 : 4'b0111;
																assign node19680 = (inp[12]) ? 4'b0011 : 4'b0111;
													assign node19683 = (inp[10]) ? node19693 : node19684;
														assign node19684 = (inp[12]) ? 4'b0110 : node19685;
															assign node19685 = (inp[4]) ? node19689 : node19686;
																assign node19686 = (inp[9]) ? 4'b0010 : 4'b0110;
																assign node19689 = (inp[9]) ? 4'b0110 : 4'b0010;
														assign node19693 = (inp[12]) ? node19701 : node19694;
															assign node19694 = (inp[9]) ? node19698 : node19695;
																assign node19695 = (inp[4]) ? 4'b0010 : 4'b0110;
																assign node19698 = (inp[4]) ? 4'b0110 : 4'b0010;
															assign node19701 = (inp[9]) ? node19705 : node19702;
																assign node19702 = (inp[4]) ? 4'b0110 : 4'b0010;
																assign node19705 = (inp[4]) ? 4'b0010 : 4'b0110;
												assign node19708 = (inp[10]) ? node19736 : node19709;
													assign node19709 = (inp[14]) ? node19723 : node19710;
														assign node19710 = (inp[12]) ? node19718 : node19711;
															assign node19711 = (inp[4]) ? node19715 : node19712;
																assign node19712 = (inp[9]) ? 4'b0010 : 4'b0110;
																assign node19715 = (inp[9]) ? 4'b0110 : 4'b0010;
															assign node19718 = (inp[4]) ? 4'b0110 : node19719;
																assign node19719 = (inp[9]) ? 4'b0010 : 4'b0110;
														assign node19723 = (inp[12]) ? node19729 : node19724;
															assign node19724 = (inp[4]) ? node19726 : 4'b0110;
																assign node19726 = (inp[9]) ? 4'b0110 : 4'b0010;
															assign node19729 = (inp[4]) ? node19733 : node19730;
																assign node19730 = (inp[9]) ? 4'b0010 : 4'b0110;
																assign node19733 = (inp[9]) ? 4'b0110 : 4'b0010;
													assign node19736 = (inp[12]) ? node19744 : node19737;
														assign node19737 = (inp[4]) ? node19741 : node19738;
															assign node19738 = (inp[9]) ? 4'b0010 : 4'b0110;
															assign node19741 = (inp[9]) ? 4'b0110 : 4'b0010;
														assign node19744 = (inp[4]) ? node19748 : node19745;
															assign node19745 = (inp[9]) ? 4'b0110 : 4'b0010;
															assign node19748 = (inp[9]) ? 4'b0010 : 4'b0110;
							assign node19751 = (inp[5]) ? node20321 : node19752;
								assign node19752 = (inp[3]) ? node20046 : node19753;
									assign node19753 = (inp[10]) ? node19891 : node19754;
										assign node19754 = (inp[8]) ? node19818 : node19755;
											assign node19755 = (inp[7]) ? node19797 : node19756;
												assign node19756 = (inp[14]) ? node19782 : node19757;
													assign node19757 = (inp[2]) ? node19767 : node19758;
														assign node19758 = (inp[12]) ? 4'b0111 : node19759;
															assign node19759 = (inp[4]) ? node19763 : node19760;
																assign node19760 = (inp[9]) ? 4'b0011 : 4'b0111;
																assign node19763 = (inp[9]) ? 4'b0111 : 4'b0011;
														assign node19767 = (inp[12]) ? node19775 : node19768;
															assign node19768 = (inp[4]) ? node19772 : node19769;
																assign node19769 = (inp[9]) ? 4'b0010 : 4'b0110;
																assign node19772 = (inp[9]) ? 4'b0110 : 4'b0010;
															assign node19775 = (inp[4]) ? node19779 : node19776;
																assign node19776 = (inp[9]) ? 4'b0010 : 4'b0110;
																assign node19779 = (inp[9]) ? 4'b0110 : 4'b0010;
													assign node19782 = (inp[2]) ? node19790 : node19783;
														assign node19783 = (inp[4]) ? node19787 : node19784;
															assign node19784 = (inp[9]) ? 4'b0010 : 4'b0110;
															assign node19787 = (inp[9]) ? 4'b0110 : 4'b0010;
														assign node19790 = (inp[9]) ? node19794 : node19791;
															assign node19791 = (inp[4]) ? 4'b0010 : 4'b0110;
															assign node19794 = (inp[4]) ? 4'b0110 : 4'b0010;
												assign node19797 = (inp[2]) ? node19811 : node19798;
													assign node19798 = (inp[14]) ? node19804 : node19799;
														assign node19799 = (inp[4]) ? 4'b0010 : node19800;
															assign node19800 = (inp[9]) ? 4'b0010 : 4'b0110;
														assign node19804 = (inp[9]) ? node19808 : node19805;
															assign node19805 = (inp[4]) ? 4'b0011 : 4'b0111;
															assign node19808 = (inp[4]) ? 4'b0111 : 4'b0011;
													assign node19811 = (inp[9]) ? node19815 : node19812;
														assign node19812 = (inp[4]) ? 4'b0011 : 4'b0111;
														assign node19815 = (inp[4]) ? 4'b0111 : 4'b0011;
											assign node19818 = (inp[7]) ? node19856 : node19819;
												assign node19819 = (inp[14]) ? node19835 : node19820;
													assign node19820 = (inp[2]) ? node19828 : node19821;
														assign node19821 = (inp[9]) ? node19825 : node19822;
															assign node19822 = (inp[4]) ? 4'b0010 : 4'b0110;
															assign node19825 = (inp[4]) ? 4'b0110 : 4'b0010;
														assign node19828 = (inp[9]) ? node19832 : node19829;
															assign node19829 = (inp[4]) ? 4'b0011 : 4'b0111;
															assign node19832 = (inp[4]) ? 4'b0111 : 4'b0011;
													assign node19835 = (inp[12]) ? node19843 : node19836;
														assign node19836 = (inp[4]) ? node19840 : node19837;
															assign node19837 = (inp[9]) ? 4'b0011 : 4'b0111;
															assign node19840 = (inp[9]) ? 4'b0111 : 4'b0011;
														assign node19843 = (inp[2]) ? node19851 : node19844;
															assign node19844 = (inp[9]) ? node19848 : node19845;
																assign node19845 = (inp[4]) ? 4'b0011 : 4'b0111;
																assign node19848 = (inp[4]) ? 4'b0111 : 4'b0011;
															assign node19851 = (inp[9]) ? node19853 : 4'b0111;
																assign node19853 = (inp[4]) ? 4'b0111 : 4'b0011;
												assign node19856 = (inp[14]) ? node19878 : node19857;
													assign node19857 = (inp[2]) ? node19867 : node19858;
														assign node19858 = (inp[12]) ? node19860 : 4'b0111;
															assign node19860 = (inp[4]) ? node19864 : node19861;
																assign node19861 = (inp[9]) ? 4'b0011 : 4'b0111;
																assign node19864 = (inp[9]) ? 4'b0111 : 4'b0011;
														assign node19867 = (inp[12]) ? node19873 : node19868;
															assign node19868 = (inp[9]) ? 4'b0110 : node19869;
																assign node19869 = (inp[4]) ? 4'b0010 : 4'b0110;
															assign node19873 = (inp[9]) ? node19875 : 4'b0110;
																assign node19875 = (inp[4]) ? 4'b0110 : 4'b0010;
													assign node19878 = (inp[2]) ? node19886 : node19879;
														assign node19879 = (inp[4]) ? node19883 : node19880;
															assign node19880 = (inp[9]) ? 4'b0010 : 4'b0110;
															assign node19883 = (inp[9]) ? 4'b0110 : 4'b0010;
														assign node19886 = (inp[9]) ? node19888 : 4'b0010;
															assign node19888 = (inp[4]) ? 4'b0110 : 4'b0010;
										assign node19891 = (inp[2]) ? node19977 : node19892;
											assign node19892 = (inp[12]) ? node19930 : node19893;
												assign node19893 = (inp[7]) ? node19913 : node19894;
													assign node19894 = (inp[14]) ? node19904 : node19895;
														assign node19895 = (inp[8]) ? 4'b0110 : node19896;
															assign node19896 = (inp[4]) ? node19900 : node19897;
																assign node19897 = (inp[9]) ? 4'b0011 : 4'b0111;
																assign node19900 = (inp[9]) ? 4'b0111 : 4'b0011;
														assign node19904 = (inp[8]) ? node19906 : 4'b0110;
															assign node19906 = (inp[4]) ? node19910 : node19907;
																assign node19907 = (inp[9]) ? 4'b0011 : 4'b0111;
																assign node19910 = (inp[9]) ? 4'b0111 : 4'b0011;
													assign node19913 = (inp[9]) ? node19921 : node19914;
														assign node19914 = (inp[4]) ? node19916 : 4'b0111;
															assign node19916 = (inp[14]) ? node19918 : 4'b0011;
																assign node19918 = (inp[8]) ? 4'b0010 : 4'b0011;
														assign node19921 = (inp[4]) ? node19927 : node19922;
															assign node19922 = (inp[8]) ? 4'b0010 : node19923;
																assign node19923 = (inp[14]) ? 4'b0011 : 4'b0010;
															assign node19927 = (inp[14]) ? 4'b0111 : 4'b0110;
												assign node19930 = (inp[7]) ? node19954 : node19931;
													assign node19931 = (inp[14]) ? node19945 : node19932;
														assign node19932 = (inp[8]) ? node19940 : node19933;
															assign node19933 = (inp[9]) ? node19937 : node19934;
																assign node19934 = (inp[4]) ? 4'b0111 : 4'b0011;
																assign node19937 = (inp[4]) ? 4'b0011 : 4'b0111;
															assign node19940 = (inp[4]) ? 4'b0110 : node19941;
																assign node19941 = (inp[9]) ? 4'b0110 : 4'b0010;
														assign node19945 = (inp[8]) ? 4'b0011 : node19946;
															assign node19946 = (inp[4]) ? node19950 : node19947;
																assign node19947 = (inp[9]) ? 4'b0110 : 4'b0010;
																assign node19950 = (inp[9]) ? 4'b0010 : 4'b0110;
													assign node19954 = (inp[14]) ? node19970 : node19955;
														assign node19955 = (inp[8]) ? node19963 : node19956;
															assign node19956 = (inp[4]) ? node19960 : node19957;
																assign node19957 = (inp[9]) ? 4'b0110 : 4'b0010;
																assign node19960 = (inp[9]) ? 4'b0010 : 4'b0110;
															assign node19963 = (inp[4]) ? node19967 : node19964;
																assign node19964 = (inp[9]) ? 4'b0111 : 4'b0011;
																assign node19967 = (inp[9]) ? 4'b0011 : 4'b0111;
														assign node19970 = (inp[8]) ? 4'b0110 : node19971;
															assign node19971 = (inp[9]) ? node19973 : 4'b0111;
																assign node19973 = (inp[4]) ? 4'b0011 : 4'b0111;
											assign node19977 = (inp[12]) ? node20011 : node19978;
												assign node19978 = (inp[4]) ? node19994 : node19979;
													assign node19979 = (inp[9]) ? node19987 : node19980;
														assign node19980 = (inp[14]) ? 4'b0111 : node19981;
															assign node19981 = (inp[8]) ? 4'b0110 : node19982;
																assign node19982 = (inp[7]) ? 4'b0111 : 4'b0110;
														assign node19987 = (inp[8]) ? node19991 : node19988;
															assign node19988 = (inp[7]) ? 4'b0011 : 4'b0010;
															assign node19991 = (inp[7]) ? 4'b0010 : 4'b0011;
													assign node19994 = (inp[9]) ? node20004 : node19995;
														assign node19995 = (inp[14]) ? 4'b0010 : node19996;
															assign node19996 = (inp[8]) ? node20000 : node19997;
																assign node19997 = (inp[7]) ? 4'b0011 : 4'b0010;
																assign node20000 = (inp[7]) ? 4'b0010 : 4'b0011;
														assign node20004 = (inp[8]) ? node20008 : node20005;
															assign node20005 = (inp[7]) ? 4'b0111 : 4'b0110;
															assign node20008 = (inp[7]) ? 4'b0110 : 4'b0111;
												assign node20011 = (inp[9]) ? node20033 : node20012;
													assign node20012 = (inp[4]) ? node20020 : node20013;
														assign node20013 = (inp[7]) ? node20017 : node20014;
															assign node20014 = (inp[8]) ? 4'b0011 : 4'b0010;
															assign node20017 = (inp[14]) ? 4'b0010 : 4'b0011;
														assign node20020 = (inp[14]) ? node20028 : node20021;
															assign node20021 = (inp[8]) ? node20025 : node20022;
																assign node20022 = (inp[7]) ? 4'b0111 : 4'b0110;
																assign node20025 = (inp[7]) ? 4'b0110 : 4'b0111;
															assign node20028 = (inp[8]) ? node20030 : 4'b0111;
																assign node20030 = (inp[7]) ? 4'b0110 : 4'b0111;
													assign node20033 = (inp[4]) ? node20041 : node20034;
														assign node20034 = (inp[8]) ? node20038 : node20035;
															assign node20035 = (inp[7]) ? 4'b0111 : 4'b0110;
															assign node20038 = (inp[7]) ? 4'b0110 : 4'b0111;
														assign node20041 = (inp[7]) ? node20043 : 4'b0010;
															assign node20043 = (inp[8]) ? 4'b0010 : 4'b0011;
									assign node20046 = (inp[4]) ? node20180 : node20047;
										assign node20047 = (inp[9]) ? node20117 : node20048;
											assign node20048 = (inp[10]) ? node20084 : node20049;
												assign node20049 = (inp[14]) ? node20071 : node20050;
													assign node20050 = (inp[12]) ? node20056 : node20051;
														assign node20051 = (inp[8]) ? node20053 : 4'b0110;
															assign node20053 = (inp[2]) ? 4'b0111 : 4'b0110;
														assign node20056 = (inp[2]) ? node20064 : node20057;
															assign node20057 = (inp[8]) ? node20061 : node20058;
																assign node20058 = (inp[7]) ? 4'b0110 : 4'b0111;
																assign node20061 = (inp[7]) ? 4'b0111 : 4'b0110;
															assign node20064 = (inp[8]) ? node20068 : node20065;
																assign node20065 = (inp[7]) ? 4'b0111 : 4'b0110;
																assign node20068 = (inp[7]) ? 4'b0110 : 4'b0111;
													assign node20071 = (inp[2]) ? node20077 : node20072;
														assign node20072 = (inp[8]) ? 4'b0111 : node20073;
															assign node20073 = (inp[7]) ? 4'b0111 : 4'b0110;
														assign node20077 = (inp[8]) ? node20081 : node20078;
															assign node20078 = (inp[7]) ? 4'b0111 : 4'b0110;
															assign node20081 = (inp[7]) ? 4'b0110 : 4'b0111;
												assign node20084 = (inp[12]) ? node20098 : node20085;
													assign node20085 = (inp[7]) ? node20093 : node20086;
														assign node20086 = (inp[8]) ? 4'b0111 : node20087;
															assign node20087 = (inp[2]) ? 4'b0110 : node20088;
																assign node20088 = (inp[14]) ? 4'b0110 : 4'b0111;
														assign node20093 = (inp[8]) ? 4'b0110 : node20094;
															assign node20094 = (inp[2]) ? 4'b0111 : 4'b0110;
													assign node20098 = (inp[2]) ? node20108 : node20099;
														assign node20099 = (inp[14]) ? node20101 : 4'b0010;
															assign node20101 = (inp[7]) ? node20105 : node20102;
																assign node20102 = (inp[8]) ? 4'b0011 : 4'b0010;
																assign node20105 = (inp[8]) ? 4'b0010 : 4'b0011;
														assign node20108 = (inp[14]) ? 4'b0010 : node20109;
															assign node20109 = (inp[7]) ? node20113 : node20110;
																assign node20110 = (inp[8]) ? 4'b0011 : 4'b0010;
																assign node20113 = (inp[8]) ? 4'b0010 : 4'b0011;
											assign node20117 = (inp[12]) ? node20141 : node20118;
												assign node20118 = (inp[7]) ? node20130 : node20119;
													assign node20119 = (inp[8]) ? node20125 : node20120;
														assign node20120 = (inp[14]) ? 4'b0010 : node20121;
															assign node20121 = (inp[2]) ? 4'b0010 : 4'b0011;
														assign node20125 = (inp[14]) ? 4'b0011 : node20126;
															assign node20126 = (inp[2]) ? 4'b0011 : 4'b0010;
													assign node20130 = (inp[8]) ? node20136 : node20131;
														assign node20131 = (inp[14]) ? 4'b0011 : node20132;
															assign node20132 = (inp[2]) ? 4'b0011 : 4'b0010;
														assign node20136 = (inp[14]) ? 4'b0010 : node20137;
															assign node20137 = (inp[2]) ? 4'b0010 : 4'b0011;
												assign node20141 = (inp[10]) ? node20163 : node20142;
													assign node20142 = (inp[14]) ? node20156 : node20143;
														assign node20143 = (inp[7]) ? node20149 : node20144;
															assign node20144 = (inp[8]) ? 4'b0010 : node20145;
																assign node20145 = (inp[2]) ? 4'b0010 : 4'b0011;
															assign node20149 = (inp[2]) ? node20153 : node20150;
																assign node20150 = (inp[8]) ? 4'b0011 : 4'b0010;
																assign node20153 = (inp[8]) ? 4'b0010 : 4'b0011;
														assign node20156 = (inp[8]) ? node20160 : node20157;
															assign node20157 = (inp[7]) ? 4'b0011 : 4'b0010;
															assign node20160 = (inp[7]) ? 4'b0010 : 4'b0011;
													assign node20163 = (inp[14]) ? node20173 : node20164;
														assign node20164 = (inp[8]) ? 4'b0101 : node20165;
															assign node20165 = (inp[7]) ? node20169 : node20166;
																assign node20166 = (inp[2]) ? 4'b0100 : 4'b0101;
																assign node20169 = (inp[2]) ? 4'b0101 : 4'b0100;
														assign node20173 = (inp[8]) ? node20177 : node20174;
															assign node20174 = (inp[7]) ? 4'b0101 : 4'b0100;
															assign node20177 = (inp[7]) ? 4'b0100 : 4'b0101;
										assign node20180 = (inp[9]) ? node20246 : node20181;
											assign node20181 = (inp[12]) ? node20211 : node20182;
												assign node20182 = (inp[2]) ? node20198 : node20183;
													assign node20183 = (inp[7]) ? node20191 : node20184;
														assign node20184 = (inp[8]) ? node20188 : node20185;
															assign node20185 = (inp[14]) ? 4'b0010 : 4'b0011;
															assign node20188 = (inp[14]) ? 4'b0011 : 4'b0010;
														assign node20191 = (inp[14]) ? node20195 : node20192;
															assign node20192 = (inp[8]) ? 4'b0011 : 4'b0010;
															assign node20195 = (inp[8]) ? 4'b0010 : 4'b0011;
													assign node20198 = (inp[10]) ? node20204 : node20199;
														assign node20199 = (inp[8]) ? node20201 : 4'b0010;
															assign node20201 = (inp[7]) ? 4'b0010 : 4'b0011;
														assign node20204 = (inp[7]) ? node20208 : node20205;
															assign node20205 = (inp[8]) ? 4'b0011 : 4'b0010;
															assign node20208 = (inp[8]) ? 4'b0010 : 4'b0011;
												assign node20211 = (inp[10]) ? node20229 : node20212;
													assign node20212 = (inp[2]) ? node20222 : node20213;
														assign node20213 = (inp[14]) ? 4'b0010 : node20214;
															assign node20214 = (inp[7]) ? node20218 : node20215;
																assign node20215 = (inp[8]) ? 4'b0010 : 4'b0011;
																assign node20218 = (inp[8]) ? 4'b0011 : 4'b0010;
														assign node20222 = (inp[8]) ? node20226 : node20223;
															assign node20223 = (inp[7]) ? 4'b0011 : 4'b0010;
															assign node20226 = (inp[7]) ? 4'b0010 : 4'b0011;
													assign node20229 = (inp[7]) ? node20241 : node20230;
														assign node20230 = (inp[8]) ? node20236 : node20231;
															assign node20231 = (inp[14]) ? 4'b0100 : node20232;
																assign node20232 = (inp[2]) ? 4'b0100 : 4'b0101;
															assign node20236 = (inp[14]) ? 4'b0101 : node20237;
																assign node20237 = (inp[2]) ? 4'b0101 : 4'b0100;
														assign node20241 = (inp[14]) ? node20243 : 4'b0100;
															assign node20243 = (inp[8]) ? 4'b0100 : 4'b0101;
											assign node20246 = (inp[12]) ? node20282 : node20247;
												assign node20247 = (inp[10]) ? node20261 : node20248;
													assign node20248 = (inp[8]) ? node20254 : node20249;
														assign node20249 = (inp[7]) ? node20251 : 4'b0100;
															assign node20251 = (inp[14]) ? 4'b0101 : 4'b0100;
														assign node20254 = (inp[7]) ? node20256 : 4'b0101;
															assign node20256 = (inp[2]) ? 4'b0100 : node20257;
																assign node20257 = (inp[14]) ? 4'b0100 : 4'b0101;
													assign node20261 = (inp[8]) ? node20273 : node20262;
														assign node20262 = (inp[7]) ? node20268 : node20263;
															assign node20263 = (inp[14]) ? 4'b0100 : node20264;
																assign node20264 = (inp[2]) ? 4'b0100 : 4'b0101;
															assign node20268 = (inp[14]) ? 4'b0101 : node20269;
																assign node20269 = (inp[2]) ? 4'b0101 : 4'b0100;
														assign node20273 = (inp[7]) ? node20279 : node20274;
															assign node20274 = (inp[14]) ? 4'b0101 : node20275;
																assign node20275 = (inp[2]) ? 4'b0101 : 4'b0100;
															assign node20279 = (inp[14]) ? 4'b0100 : 4'b0101;
												assign node20282 = (inp[10]) ? node20298 : node20283;
													assign node20283 = (inp[8]) ? node20291 : node20284;
														assign node20284 = (inp[7]) ? node20286 : 4'b0100;
															assign node20286 = (inp[2]) ? 4'b0101 : node20287;
																assign node20287 = (inp[14]) ? 4'b0101 : 4'b0100;
														assign node20291 = (inp[7]) ? node20293 : 4'b0101;
															assign node20293 = (inp[2]) ? 4'b0100 : node20294;
																assign node20294 = (inp[14]) ? 4'b0100 : 4'b0101;
													assign node20298 = (inp[14]) ? node20314 : node20299;
														assign node20299 = (inp[7]) ? node20307 : node20300;
															assign node20300 = (inp[2]) ? node20304 : node20301;
																assign node20301 = (inp[8]) ? 4'b0000 : 4'b0001;
																assign node20304 = (inp[8]) ? 4'b0001 : 4'b0000;
															assign node20307 = (inp[2]) ? node20311 : node20308;
																assign node20308 = (inp[8]) ? 4'b0001 : 4'b0000;
																assign node20311 = (inp[8]) ? 4'b0000 : 4'b0001;
														assign node20314 = (inp[8]) ? node20318 : node20315;
															assign node20315 = (inp[7]) ? 4'b0001 : 4'b0000;
															assign node20318 = (inp[7]) ? 4'b0000 : 4'b0001;
								assign node20321 = (inp[3]) ? node20559 : node20322;
									assign node20322 = (inp[9]) ? node20440 : node20323;
										assign node20323 = (inp[4]) ? node20385 : node20324;
											assign node20324 = (inp[12]) ? node20348 : node20325;
												assign node20325 = (inp[8]) ? node20337 : node20326;
													assign node20326 = (inp[7]) ? node20332 : node20327;
														assign node20327 = (inp[2]) ? 4'b0110 : node20328;
															assign node20328 = (inp[14]) ? 4'b0110 : 4'b0111;
														assign node20332 = (inp[14]) ? 4'b0111 : node20333;
															assign node20333 = (inp[2]) ? 4'b0111 : 4'b0110;
													assign node20337 = (inp[7]) ? node20343 : node20338;
														assign node20338 = (inp[14]) ? 4'b0111 : node20339;
															assign node20339 = (inp[2]) ? 4'b0111 : 4'b0110;
														assign node20343 = (inp[2]) ? 4'b0110 : node20344;
															assign node20344 = (inp[14]) ? 4'b0110 : 4'b0111;
												assign node20348 = (inp[10]) ? node20370 : node20349;
													assign node20349 = (inp[2]) ? node20359 : node20350;
														assign node20350 = (inp[14]) ? 4'b0111 : node20351;
															assign node20351 = (inp[7]) ? node20355 : node20352;
																assign node20352 = (inp[8]) ? 4'b0110 : 4'b0111;
																assign node20355 = (inp[8]) ? 4'b0111 : 4'b0110;
														assign node20359 = (inp[14]) ? node20365 : node20360;
															assign node20360 = (inp[7]) ? node20362 : 4'b0111;
																assign node20362 = (inp[8]) ? 4'b0110 : 4'b0111;
															assign node20365 = (inp[8]) ? node20367 : 4'b0110;
																assign node20367 = (inp[7]) ? 4'b0110 : 4'b0111;
													assign node20370 = (inp[8]) ? node20380 : node20371;
														assign node20371 = (inp[7]) ? node20375 : node20372;
															assign node20372 = (inp[14]) ? 4'b0010 : 4'b0011;
															assign node20375 = (inp[14]) ? 4'b0011 : node20376;
																assign node20376 = (inp[2]) ? 4'b0011 : 4'b0010;
														assign node20380 = (inp[7]) ? node20382 : 4'b0011;
															assign node20382 = (inp[14]) ? 4'b0010 : 4'b0011;
											assign node20385 = (inp[12]) ? node20405 : node20386;
												assign node20386 = (inp[8]) ? node20394 : node20387;
													assign node20387 = (inp[7]) ? node20389 : 4'b0010;
														assign node20389 = (inp[2]) ? 4'b0011 : node20390;
															assign node20390 = (inp[14]) ? 4'b0011 : 4'b0010;
													assign node20394 = (inp[7]) ? node20400 : node20395;
														assign node20395 = (inp[2]) ? 4'b0011 : node20396;
															assign node20396 = (inp[14]) ? 4'b0011 : 4'b0010;
														assign node20400 = (inp[14]) ? 4'b0010 : node20401;
															assign node20401 = (inp[2]) ? 4'b0010 : 4'b0011;
												assign node20405 = (inp[10]) ? node20425 : node20406;
													assign node20406 = (inp[14]) ? node20418 : node20407;
														assign node20407 = (inp[8]) ? node20413 : node20408;
															assign node20408 = (inp[7]) ? node20410 : 4'b0011;
																assign node20410 = (inp[2]) ? 4'b0011 : 4'b0010;
															assign node20413 = (inp[2]) ? 4'b0010 : node20414;
																assign node20414 = (inp[7]) ? 4'b0011 : 4'b0010;
														assign node20418 = (inp[8]) ? node20422 : node20419;
															assign node20419 = (inp[7]) ? 4'b0011 : 4'b0010;
															assign node20422 = (inp[7]) ? 4'b0010 : 4'b0011;
													assign node20425 = (inp[8]) ? node20433 : node20426;
														assign node20426 = (inp[7]) ? 4'b0101 : node20427;
															assign node20427 = (inp[2]) ? 4'b0100 : node20428;
																assign node20428 = (inp[14]) ? 4'b0100 : 4'b0101;
														assign node20433 = (inp[7]) ? node20435 : 4'b0101;
															assign node20435 = (inp[2]) ? 4'b0100 : node20436;
																assign node20436 = (inp[14]) ? 4'b0100 : 4'b0101;
										assign node20440 = (inp[4]) ? node20494 : node20441;
											assign node20441 = (inp[12]) ? node20465 : node20442;
												assign node20442 = (inp[8]) ? node20454 : node20443;
													assign node20443 = (inp[7]) ? node20449 : node20444;
														assign node20444 = (inp[14]) ? 4'b0010 : node20445;
															assign node20445 = (inp[2]) ? 4'b0010 : 4'b0011;
														assign node20449 = (inp[14]) ? 4'b0011 : node20450;
															assign node20450 = (inp[2]) ? 4'b0011 : 4'b0010;
													assign node20454 = (inp[7]) ? node20460 : node20455;
														assign node20455 = (inp[14]) ? 4'b0011 : node20456;
															assign node20456 = (inp[2]) ? 4'b0011 : 4'b0010;
														assign node20460 = (inp[14]) ? 4'b0010 : node20461;
															assign node20461 = (inp[10]) ? 4'b0011 : 4'b0010;
												assign node20465 = (inp[10]) ? node20483 : node20466;
													assign node20466 = (inp[8]) ? node20474 : node20467;
														assign node20467 = (inp[7]) ? node20469 : 4'b0010;
															assign node20469 = (inp[2]) ? 4'b0011 : node20470;
																assign node20470 = (inp[14]) ? 4'b0011 : 4'b0010;
														assign node20474 = (inp[14]) ? 4'b0011 : node20475;
															assign node20475 = (inp[7]) ? node20479 : node20476;
																assign node20476 = (inp[2]) ? 4'b0011 : 4'b0010;
																assign node20479 = (inp[2]) ? 4'b0010 : 4'b0011;
													assign node20483 = (inp[8]) ? node20491 : node20484;
														assign node20484 = (inp[7]) ? 4'b0101 : node20485;
															assign node20485 = (inp[14]) ? 4'b0100 : node20486;
																assign node20486 = (inp[2]) ? 4'b0100 : 4'b0101;
														assign node20491 = (inp[7]) ? 4'b0100 : 4'b0101;
											assign node20494 = (inp[10]) ? node20526 : node20495;
												assign node20495 = (inp[2]) ? node20519 : node20496;
													assign node20496 = (inp[7]) ? node20504 : node20497;
														assign node20497 = (inp[8]) ? node20501 : node20498;
															assign node20498 = (inp[14]) ? 4'b0100 : 4'b0101;
															assign node20501 = (inp[14]) ? 4'b0101 : 4'b0100;
														assign node20504 = (inp[12]) ? node20512 : node20505;
															assign node20505 = (inp[14]) ? node20509 : node20506;
																assign node20506 = (inp[8]) ? 4'b0101 : 4'b0100;
																assign node20509 = (inp[8]) ? 4'b0100 : 4'b0101;
															assign node20512 = (inp[8]) ? node20516 : node20513;
																assign node20513 = (inp[14]) ? 4'b0101 : 4'b0100;
																assign node20516 = (inp[14]) ? 4'b0100 : 4'b0101;
													assign node20519 = (inp[8]) ? node20523 : node20520;
														assign node20520 = (inp[7]) ? 4'b0101 : 4'b0100;
														assign node20523 = (inp[7]) ? 4'b0100 : 4'b0101;
												assign node20526 = (inp[12]) ? node20544 : node20527;
													assign node20527 = (inp[14]) ? node20537 : node20528;
														assign node20528 = (inp[2]) ? 4'b0101 : node20529;
															assign node20529 = (inp[8]) ? node20533 : node20530;
																assign node20530 = (inp[7]) ? 4'b0100 : 4'b0101;
																assign node20533 = (inp[7]) ? 4'b0101 : 4'b0100;
														assign node20537 = (inp[8]) ? node20541 : node20538;
															assign node20538 = (inp[7]) ? 4'b0101 : 4'b0100;
															assign node20541 = (inp[7]) ? 4'b0100 : 4'b0101;
													assign node20544 = (inp[14]) ? node20554 : node20545;
														assign node20545 = (inp[2]) ? 4'b0001 : node20546;
															assign node20546 = (inp[7]) ? node20550 : node20547;
																assign node20547 = (inp[8]) ? 4'b0000 : 4'b0001;
																assign node20550 = (inp[8]) ? 4'b0001 : 4'b0000;
														assign node20554 = (inp[7]) ? node20556 : 4'b0000;
															assign node20556 = (inp[8]) ? 4'b0000 : 4'b0001;
									assign node20559 = (inp[9]) ? node20723 : node20560;
										assign node20560 = (inp[4]) ? node20632 : node20561;
											assign node20561 = (inp[10]) ? node20597 : node20562;
												assign node20562 = (inp[14]) ? node20576 : node20563;
													assign node20563 = (inp[7]) ? node20571 : node20564;
														assign node20564 = (inp[2]) ? node20568 : node20565;
															assign node20565 = (inp[8]) ? 4'b0100 : 4'b0101;
															assign node20568 = (inp[8]) ? 4'b0101 : 4'b0100;
														assign node20571 = (inp[12]) ? 4'b0100 : node20572;
															assign node20572 = (inp[2]) ? 4'b0101 : 4'b0100;
													assign node20576 = (inp[12]) ? node20590 : node20577;
														assign node20577 = (inp[2]) ? node20585 : node20578;
															assign node20578 = (inp[8]) ? node20582 : node20579;
																assign node20579 = (inp[7]) ? 4'b0101 : 4'b0100;
																assign node20582 = (inp[7]) ? 4'b0100 : 4'b0101;
															assign node20585 = (inp[8]) ? 4'b0101 : node20586;
																assign node20586 = (inp[7]) ? 4'b0101 : 4'b0100;
														assign node20590 = (inp[8]) ? node20594 : node20591;
															assign node20591 = (inp[7]) ? 4'b0101 : 4'b0100;
															assign node20594 = (inp[7]) ? 4'b0100 : 4'b0101;
												assign node20597 = (inp[12]) ? node20615 : node20598;
													assign node20598 = (inp[2]) ? node20608 : node20599;
														assign node20599 = (inp[7]) ? node20601 : 4'b0100;
															assign node20601 = (inp[14]) ? node20605 : node20602;
																assign node20602 = (inp[8]) ? 4'b0101 : 4'b0100;
																assign node20605 = (inp[8]) ? 4'b0100 : 4'b0101;
														assign node20608 = (inp[7]) ? node20612 : node20609;
															assign node20609 = (inp[8]) ? 4'b0101 : 4'b0100;
															assign node20612 = (inp[8]) ? 4'b0100 : 4'b0101;
													assign node20615 = (inp[7]) ? node20627 : node20616;
														assign node20616 = (inp[8]) ? node20622 : node20617;
															assign node20617 = (inp[2]) ? 4'b0000 : node20618;
																assign node20618 = (inp[14]) ? 4'b0000 : 4'b0001;
															assign node20622 = (inp[14]) ? 4'b0001 : node20623;
																assign node20623 = (inp[2]) ? 4'b0001 : 4'b0000;
														assign node20627 = (inp[8]) ? 4'b0000 : node20628;
															assign node20628 = (inp[14]) ? 4'b0001 : 4'b0000;
											assign node20632 = (inp[12]) ? node20682 : node20633;
												assign node20633 = (inp[10]) ? node20665 : node20634;
													assign node20634 = (inp[2]) ? node20650 : node20635;
														assign node20635 = (inp[8]) ? node20643 : node20636;
															assign node20636 = (inp[14]) ? node20640 : node20637;
																assign node20637 = (inp[7]) ? 4'b0000 : 4'b0001;
																assign node20640 = (inp[7]) ? 4'b0001 : 4'b0000;
															assign node20643 = (inp[14]) ? node20647 : node20644;
																assign node20644 = (inp[7]) ? 4'b0001 : 4'b0000;
																assign node20647 = (inp[7]) ? 4'b0000 : 4'b0001;
														assign node20650 = (inp[14]) ? node20658 : node20651;
															assign node20651 = (inp[7]) ? node20655 : node20652;
																assign node20652 = (inp[8]) ? 4'b0001 : 4'b0000;
																assign node20655 = (inp[8]) ? 4'b0000 : 4'b0001;
															assign node20658 = (inp[7]) ? node20662 : node20659;
																assign node20659 = (inp[8]) ? 4'b0001 : 4'b0000;
																assign node20662 = (inp[8]) ? 4'b0000 : 4'b0001;
													assign node20665 = (inp[8]) ? node20675 : node20666;
														assign node20666 = (inp[2]) ? node20672 : node20667;
															assign node20667 = (inp[14]) ? 4'b0001 : node20668;
																assign node20668 = (inp[7]) ? 4'b0000 : 4'b0001;
															assign node20672 = (inp[7]) ? 4'b0001 : 4'b0000;
														assign node20675 = (inp[2]) ? 4'b0000 : node20676;
															assign node20676 = (inp[7]) ? node20678 : 4'b0000;
																assign node20678 = (inp[14]) ? 4'b0000 : 4'b0001;
												assign node20682 = (inp[10]) ? node20694 : node20683;
													assign node20683 = (inp[7]) ? node20689 : node20684;
														assign node20684 = (inp[2]) ? 4'b0000 : node20685;
															assign node20685 = (inp[8]) ? 4'b0000 : 4'b0001;
														assign node20689 = (inp[8]) ? node20691 : 4'b0001;
															assign node20691 = (inp[14]) ? 4'b0000 : 4'b0001;
													assign node20694 = (inp[2]) ? node20710 : node20695;
														assign node20695 = (inp[7]) ? node20703 : node20696;
															assign node20696 = (inp[14]) ? node20700 : node20697;
																assign node20697 = (inp[8]) ? 4'b0100 : 4'b0101;
																assign node20700 = (inp[8]) ? 4'b0101 : 4'b0100;
															assign node20703 = (inp[8]) ? node20707 : node20704;
																assign node20704 = (inp[14]) ? 4'b0101 : 4'b0100;
																assign node20707 = (inp[14]) ? 4'b0100 : 4'b0101;
														assign node20710 = (inp[14]) ? node20716 : node20711;
															assign node20711 = (inp[8]) ? 4'b0101 : node20712;
																assign node20712 = (inp[7]) ? 4'b0101 : 4'b0100;
															assign node20716 = (inp[8]) ? node20720 : node20717;
																assign node20717 = (inp[7]) ? 4'b0101 : 4'b0100;
																assign node20720 = (inp[7]) ? 4'b0100 : 4'b0101;
										assign node20723 = (inp[4]) ? node20789 : node20724;
											assign node20724 = (inp[10]) ? node20758 : node20725;
												assign node20725 = (inp[2]) ? node20745 : node20726;
													assign node20726 = (inp[8]) ? node20738 : node20727;
														assign node20727 = (inp[12]) ? node20733 : node20728;
															assign node20728 = (inp[14]) ? 4'b0001 : node20729;
																assign node20729 = (inp[7]) ? 4'b0000 : 4'b0001;
															assign node20733 = (inp[7]) ? 4'b0001 : node20734;
																assign node20734 = (inp[14]) ? 4'b0000 : 4'b0001;
														assign node20738 = (inp[7]) ? node20742 : node20739;
															assign node20739 = (inp[14]) ? 4'b0001 : 4'b0000;
															assign node20742 = (inp[14]) ? 4'b0000 : 4'b0001;
													assign node20745 = (inp[14]) ? node20753 : node20746;
														assign node20746 = (inp[7]) ? node20750 : node20747;
															assign node20747 = (inp[8]) ? 4'b0001 : 4'b0000;
															assign node20750 = (inp[8]) ? 4'b0000 : 4'b0001;
														assign node20753 = (inp[7]) ? 4'b0000 : node20754;
															assign node20754 = (inp[8]) ? 4'b0001 : 4'b0000;
												assign node20758 = (inp[12]) ? node20778 : node20759;
													assign node20759 = (inp[2]) ? node20769 : node20760;
														assign node20760 = (inp[7]) ? 4'b0001 : node20761;
															assign node20761 = (inp[14]) ? node20765 : node20762;
																assign node20762 = (inp[8]) ? 4'b0000 : 4'b0001;
																assign node20765 = (inp[8]) ? 4'b0001 : 4'b0000;
														assign node20769 = (inp[14]) ? node20773 : node20770;
															assign node20770 = (inp[8]) ? 4'b0000 : 4'b0001;
															assign node20773 = (inp[7]) ? 4'b0000 : node20774;
																assign node20774 = (inp[8]) ? 4'b0001 : 4'b0000;
													assign node20778 = (inp[7]) ? node20784 : node20779;
														assign node20779 = (inp[8]) ? 4'b0101 : node20780;
															assign node20780 = (inp[2]) ? 4'b0100 : 4'b0101;
														assign node20784 = (inp[2]) ? node20786 : 4'b0100;
															assign node20786 = (inp[8]) ? 4'b0100 : 4'b0101;
											assign node20789 = (inp[12]) ? node20819 : node20790;
												assign node20790 = (inp[2]) ? node20806 : node20791;
													assign node20791 = (inp[7]) ? node20799 : node20792;
														assign node20792 = (inp[8]) ? node20796 : node20793;
															assign node20793 = (inp[14]) ? 4'b0100 : 4'b0101;
															assign node20796 = (inp[14]) ? 4'b0101 : 4'b0100;
														assign node20799 = (inp[14]) ? node20803 : node20800;
															assign node20800 = (inp[8]) ? 4'b0101 : 4'b0100;
															assign node20803 = (inp[8]) ? 4'b0100 : 4'b0101;
													assign node20806 = (inp[10]) ? node20814 : node20807;
														assign node20807 = (inp[8]) ? node20811 : node20808;
															assign node20808 = (inp[7]) ? 4'b0101 : 4'b0100;
															assign node20811 = (inp[7]) ? 4'b0100 : 4'b0101;
														assign node20814 = (inp[7]) ? 4'b0101 : node20815;
															assign node20815 = (inp[8]) ? 4'b0101 : 4'b0100;
												assign node20819 = (inp[10]) ? node20839 : node20820;
													assign node20820 = (inp[8]) ? node20832 : node20821;
														assign node20821 = (inp[7]) ? node20827 : node20822;
															assign node20822 = (inp[14]) ? 4'b0100 : node20823;
																assign node20823 = (inp[2]) ? 4'b0100 : 4'b0101;
															assign node20827 = (inp[2]) ? 4'b0101 : node20828;
																assign node20828 = (inp[14]) ? 4'b0101 : 4'b0100;
														assign node20832 = (inp[7]) ? 4'b0100 : node20833;
															assign node20833 = (inp[14]) ? 4'b0101 : node20834;
																assign node20834 = (inp[2]) ? 4'b0101 : 4'b0100;
													assign node20839 = (inp[2]) ? node20847 : node20840;
														assign node20840 = (inp[14]) ? node20842 : 4'b0001;
															assign node20842 = (inp[7]) ? 4'b0000 : node20843;
																assign node20843 = (inp[8]) ? 4'b0001 : 4'b0000;
														assign node20847 = (inp[8]) ? node20851 : node20848;
															assign node20848 = (inp[7]) ? 4'b0001 : 4'b0000;
															assign node20851 = (inp[7]) ? 4'b0000 : 4'b0001;
					assign node20854 = (inp[7]) ? node22788 : node20855;
						assign node20855 = (inp[8]) ? node21869 : node20856;
							assign node20856 = (inp[2]) ? node21404 : node20857;
								assign node20857 = (inp[14]) ? node21147 : node20858;
									assign node20858 = (inp[4]) ? node20994 : node20859;
										assign node20859 = (inp[9]) ? node20917 : node20860;
											assign node20860 = (inp[10]) ? node20892 : node20861;
												assign node20861 = (inp[5]) ? node20879 : node20862;
													assign node20862 = (inp[12]) ? node20872 : node20863;
														assign node20863 = (inp[3]) ? node20865 : 4'b0101;
															assign node20865 = (inp[0]) ? node20869 : node20866;
																assign node20866 = (inp[15]) ? 4'b0101 : 4'b0111;
																assign node20869 = (inp[15]) ? 4'b0111 : 4'b0101;
														assign node20872 = (inp[3]) ? node20874 : 4'b0111;
															assign node20874 = (inp[0]) ? 4'b0111 : node20875;
																assign node20875 = (inp[15]) ? 4'b0101 : 4'b0111;
													assign node20879 = (inp[0]) ? node20887 : node20880;
														assign node20880 = (inp[15]) ? node20884 : node20881;
															assign node20881 = (inp[3]) ? 4'b0101 : 4'b0111;
															assign node20884 = (inp[3]) ? 4'b0111 : 4'b0101;
														assign node20887 = (inp[15]) ? 4'b0101 : node20888;
															assign node20888 = (inp[3]) ? 4'b0111 : 4'b0101;
												assign node20892 = (inp[12]) ? node20904 : node20893;
													assign node20893 = (inp[5]) ? node20895 : 4'b0101;
														assign node20895 = (inp[3]) ? node20897 : 4'b0111;
															assign node20897 = (inp[15]) ? node20901 : node20898;
																assign node20898 = (inp[0]) ? 4'b0111 : 4'b0101;
																assign node20901 = (inp[0]) ? 4'b0101 : 4'b0111;
													assign node20904 = (inp[15]) ? node20914 : node20905;
														assign node20905 = (inp[3]) ? node20907 : 4'b0011;
															assign node20907 = (inp[0]) ? node20911 : node20908;
																assign node20908 = (inp[5]) ? 4'b0001 : 4'b0011;
																assign node20911 = (inp[5]) ? 4'b0011 : 4'b0001;
														assign node20914 = (inp[0]) ? 4'b0011 : 4'b0001;
											assign node20917 = (inp[12]) ? node20953 : node20918;
												assign node20918 = (inp[10]) ? node20938 : node20919;
													assign node20919 = (inp[0]) ? node20931 : node20920;
														assign node20920 = (inp[15]) ? node20926 : node20921;
															assign node20921 = (inp[5]) ? node20923 : 4'b0011;
																assign node20923 = (inp[3]) ? 4'b0001 : 4'b0011;
															assign node20926 = (inp[3]) ? node20928 : 4'b0001;
																assign node20928 = (inp[5]) ? 4'b0011 : 4'b0001;
														assign node20931 = (inp[15]) ? 4'b0011 : node20932;
															assign node20932 = (inp[3]) ? node20934 : 4'b0001;
																assign node20934 = (inp[5]) ? 4'b0011 : 4'b0001;
													assign node20938 = (inp[5]) ? node20946 : node20939;
														assign node20939 = (inp[0]) ? node20943 : node20940;
															assign node20940 = (inp[15]) ? 4'b0001 : 4'b0011;
															assign node20943 = (inp[15]) ? 4'b0011 : 4'b0001;
														assign node20946 = (inp[15]) ? 4'b0001 : node20947;
															assign node20947 = (inp[0]) ? node20949 : 4'b0001;
																assign node20949 = (inp[3]) ? 4'b0011 : 4'b0001;
												assign node20953 = (inp[10]) ? node20971 : node20954;
													assign node20954 = (inp[0]) ? node20960 : node20955;
														assign node20955 = (inp[15]) ? 4'b0001 : node20956;
															assign node20956 = (inp[3]) ? 4'b0001 : 4'b0011;
														assign node20960 = (inp[15]) ? node20966 : node20961;
															assign node20961 = (inp[3]) ? node20963 : 4'b0001;
																assign node20963 = (inp[5]) ? 4'b0011 : 4'b0001;
															assign node20966 = (inp[5]) ? node20968 : 4'b0011;
																assign node20968 = (inp[3]) ? 4'b0001 : 4'b0011;
													assign node20971 = (inp[5]) ? node20985 : node20972;
														assign node20972 = (inp[3]) ? node20980 : node20973;
															assign node20973 = (inp[15]) ? node20977 : node20974;
																assign node20974 = (inp[0]) ? 4'b0101 : 4'b0111;
																assign node20977 = (inp[0]) ? 4'b0111 : 4'b0101;
															assign node20980 = (inp[15]) ? node20982 : 4'b0111;
																assign node20982 = (inp[0]) ? 4'b0101 : 4'b0111;
														assign node20985 = (inp[3]) ? 4'b0101 : node20986;
															assign node20986 = (inp[15]) ? node20990 : node20987;
																assign node20987 = (inp[0]) ? 4'b0111 : 4'b0101;
																assign node20990 = (inp[0]) ? 4'b0101 : 4'b0111;
										assign node20994 = (inp[9]) ? node21066 : node20995;
											assign node20995 = (inp[10]) ? node21029 : node20996;
												assign node20996 = (inp[3]) ? node21010 : node20997;
													assign node20997 = (inp[12]) ? node21003 : node20998;
														assign node20998 = (inp[5]) ? 4'b0011 : node20999;
															assign node20999 = (inp[0]) ? 4'b0011 : 4'b0001;
														assign node21003 = (inp[15]) ? node21007 : node21004;
															assign node21004 = (inp[0]) ? 4'b0001 : 4'b0011;
															assign node21007 = (inp[0]) ? 4'b0011 : 4'b0001;
													assign node21010 = (inp[15]) ? node21018 : node21011;
														assign node21011 = (inp[5]) ? node21015 : node21012;
															assign node21012 = (inp[0]) ? 4'b0001 : 4'b0011;
															assign node21015 = (inp[0]) ? 4'b0011 : 4'b0001;
														assign node21018 = (inp[12]) ? node21024 : node21019;
															assign node21019 = (inp[5]) ? 4'b0001 : node21020;
																assign node21020 = (inp[0]) ? 4'b0011 : 4'b0001;
															assign node21024 = (inp[0]) ? 4'b0001 : node21025;
																assign node21025 = (inp[5]) ? 4'b0011 : 4'b0001;
												assign node21029 = (inp[12]) ? node21045 : node21030;
													assign node21030 = (inp[15]) ? node21036 : node21031;
														assign node21031 = (inp[3]) ? node21033 : 4'b0001;
															assign node21033 = (inp[0]) ? 4'b0011 : 4'b0001;
														assign node21036 = (inp[0]) ? node21042 : node21037;
															assign node21037 = (inp[3]) ? node21039 : 4'b0001;
																assign node21039 = (inp[5]) ? 4'b0011 : 4'b0001;
															assign node21042 = (inp[3]) ? 4'b0001 : 4'b0011;
													assign node21045 = (inp[5]) ? node21059 : node21046;
														assign node21046 = (inp[15]) ? node21052 : node21047;
															assign node21047 = (inp[0]) ? node21049 : 4'b0111;
																assign node21049 = (inp[3]) ? 4'b0111 : 4'b0101;
															assign node21052 = (inp[0]) ? node21056 : node21053;
																assign node21053 = (inp[3]) ? 4'b0111 : 4'b0101;
																assign node21056 = (inp[3]) ? 4'b0101 : 4'b0111;
														assign node21059 = (inp[15]) ? node21063 : node21060;
															assign node21060 = (inp[0]) ? 4'b0111 : 4'b0101;
															assign node21063 = (inp[0]) ? 4'b0101 : 4'b0111;
											assign node21066 = (inp[12]) ? node21108 : node21067;
												assign node21067 = (inp[5]) ? node21091 : node21068;
													assign node21068 = (inp[0]) ? node21078 : node21069;
														assign node21069 = (inp[10]) ? node21071 : 4'b0111;
															assign node21071 = (inp[3]) ? node21075 : node21072;
																assign node21072 = (inp[15]) ? 4'b0101 : 4'b0111;
																assign node21075 = (inp[15]) ? 4'b0111 : 4'b0101;
														assign node21078 = (inp[10]) ? node21086 : node21079;
															assign node21079 = (inp[3]) ? node21083 : node21080;
																assign node21080 = (inp[15]) ? 4'b0111 : 4'b0101;
																assign node21083 = (inp[15]) ? 4'b0101 : 4'b0111;
															assign node21086 = (inp[15]) ? 4'b0111 : node21087;
																assign node21087 = (inp[3]) ? 4'b0111 : 4'b0101;
													assign node21091 = (inp[10]) ? node21099 : node21092;
														assign node21092 = (inp[0]) ? node21096 : node21093;
															assign node21093 = (inp[15]) ? 4'b0111 : 4'b0101;
															assign node21096 = (inp[15]) ? 4'b0101 : 4'b0111;
														assign node21099 = (inp[3]) ? node21103 : node21100;
															assign node21100 = (inp[0]) ? 4'b0101 : 4'b0111;
															assign node21103 = (inp[0]) ? 4'b0111 : node21104;
																assign node21104 = (inp[15]) ? 4'b0111 : 4'b0101;
												assign node21108 = (inp[10]) ? node21128 : node21109;
													assign node21109 = (inp[3]) ? node21121 : node21110;
														assign node21110 = (inp[5]) ? node21116 : node21111;
															assign node21111 = (inp[15]) ? 4'b0101 : node21112;
																assign node21112 = (inp[0]) ? 4'b0101 : 4'b0111;
															assign node21116 = (inp[15]) ? 4'b0111 : node21117;
																assign node21117 = (inp[0]) ? 4'b0111 : 4'b0101;
														assign node21121 = (inp[5]) ? node21123 : 4'b0111;
															assign node21123 = (inp[15]) ? 4'b0111 : node21124;
																assign node21124 = (inp[0]) ? 4'b0111 : 4'b0101;
													assign node21128 = (inp[3]) ? node21140 : node21129;
														assign node21129 = (inp[0]) ? node21135 : node21130;
															assign node21130 = (inp[5]) ? node21132 : 4'b0011;
																assign node21132 = (inp[15]) ? 4'b0011 : 4'b0001;
															assign node21135 = (inp[5]) ? node21137 : 4'b0001;
																assign node21137 = (inp[15]) ? 4'b0001 : 4'b0011;
														assign node21140 = (inp[0]) ? node21144 : node21141;
															assign node21141 = (inp[15]) ? 4'b0011 : 4'b0001;
															assign node21144 = (inp[15]) ? 4'b0001 : 4'b0011;
									assign node21147 = (inp[5]) ? node21271 : node21148;
										assign node21148 = (inp[0]) ? node21220 : node21149;
											assign node21149 = (inp[15]) ? node21179 : node21150;
												assign node21150 = (inp[3]) ? node21162 : node21151;
													assign node21151 = (inp[9]) ? node21153 : 4'b0110;
														assign node21153 = (inp[4]) ? node21157 : node21154;
															assign node21154 = (inp[10]) ? 4'b0110 : 4'b0010;
															assign node21157 = (inp[12]) ? node21159 : 4'b0110;
																assign node21159 = (inp[10]) ? 4'b0010 : 4'b0110;
													assign node21162 = (inp[9]) ? node21170 : node21163;
														assign node21163 = (inp[4]) ? 4'b0010 : node21164;
															assign node21164 = (inp[12]) ? node21166 : 4'b0110;
																assign node21166 = (inp[10]) ? 4'b0010 : 4'b0110;
														assign node21170 = (inp[4]) ? node21174 : node21171;
															assign node21171 = (inp[12]) ? 4'b0100 : 4'b0010;
															assign node21174 = (inp[12]) ? node21176 : 4'b0100;
																assign node21176 = (inp[10]) ? 4'b0000 : 4'b0100;
												assign node21179 = (inp[3]) ? node21199 : node21180;
													assign node21180 = (inp[10]) ? node21188 : node21181;
														assign node21181 = (inp[9]) ? node21185 : node21182;
															assign node21182 = (inp[4]) ? 4'b0000 : 4'b0100;
															assign node21185 = (inp[4]) ? 4'b0100 : 4'b0000;
														assign node21188 = (inp[4]) ? node21194 : node21189;
															assign node21189 = (inp[9]) ? node21191 : 4'b0000;
																assign node21191 = (inp[12]) ? 4'b0100 : 4'b0000;
															assign node21194 = (inp[12]) ? node21196 : 4'b0100;
																assign node21196 = (inp[9]) ? 4'b0000 : 4'b0100;
													assign node21199 = (inp[4]) ? node21211 : node21200;
														assign node21200 = (inp[9]) ? node21206 : node21201;
															assign node21201 = (inp[12]) ? node21203 : 4'b0100;
																assign node21203 = (inp[10]) ? 4'b0000 : 4'b0100;
															assign node21206 = (inp[10]) ? node21208 : 4'b0000;
																assign node21208 = (inp[12]) ? 4'b0110 : 4'b0000;
														assign node21211 = (inp[9]) ? node21215 : node21212;
															assign node21212 = (inp[10]) ? 4'b0110 : 4'b0000;
															assign node21215 = (inp[12]) ? node21217 : 4'b0110;
																assign node21217 = (inp[10]) ? 4'b0010 : 4'b0110;
											assign node21220 = (inp[15]) ? node21248 : node21221;
												assign node21221 = (inp[12]) ? node21235 : node21222;
													assign node21222 = (inp[3]) ? node21230 : node21223;
														assign node21223 = (inp[9]) ? node21227 : node21224;
															assign node21224 = (inp[4]) ? 4'b0000 : 4'b0100;
															assign node21227 = (inp[4]) ? 4'b0100 : 4'b0000;
														assign node21230 = (inp[4]) ? 4'b0110 : node21231;
															assign node21231 = (inp[9]) ? 4'b0000 : 4'b0100;
													assign node21235 = (inp[3]) ? node21237 : 4'b0000;
														assign node21237 = (inp[4]) ? node21243 : node21238;
															assign node21238 = (inp[9]) ? 4'b0000 : node21239;
																assign node21239 = (inp[10]) ? 4'b0000 : 4'b0100;
															assign node21243 = (inp[9]) ? node21245 : 4'b0000;
																assign node21245 = (inp[10]) ? 4'b0010 : 4'b0110;
												assign node21248 = (inp[4]) ? node21260 : node21249;
													assign node21249 = (inp[9]) ? node21255 : node21250;
														assign node21250 = (inp[10]) ? node21252 : 4'b0110;
															assign node21252 = (inp[12]) ? 4'b0010 : 4'b0110;
														assign node21255 = (inp[12]) ? node21257 : 4'b0010;
															assign node21257 = (inp[10]) ? 4'b0110 : 4'b0010;
													assign node21260 = (inp[9]) ? node21268 : node21261;
														assign node21261 = (inp[12]) ? node21263 : 4'b0010;
															assign node21263 = (inp[10]) ? node21265 : 4'b0010;
																assign node21265 = (inp[3]) ? 4'b0100 : 4'b0110;
														assign node21268 = (inp[3]) ? 4'b0100 : 4'b0110;
										assign node21271 = (inp[15]) ? node21337 : node21272;
											assign node21272 = (inp[0]) ? node21306 : node21273;
												assign node21273 = (inp[3]) ? node21293 : node21274;
													assign node21274 = (inp[9]) ? node21282 : node21275;
														assign node21275 = (inp[4]) ? 4'b0010 : node21276;
															assign node21276 = (inp[10]) ? node21278 : 4'b0110;
																assign node21278 = (inp[12]) ? 4'b0010 : 4'b0110;
														assign node21282 = (inp[4]) ? node21288 : node21283;
															assign node21283 = (inp[12]) ? node21285 : 4'b0010;
																assign node21285 = (inp[10]) ? 4'b0100 : 4'b0010;
															assign node21288 = (inp[12]) ? node21290 : 4'b0100;
																assign node21290 = (inp[10]) ? 4'b0000 : 4'b0100;
													assign node21293 = (inp[4]) ? node21301 : node21294;
														assign node21294 = (inp[9]) ? 4'b0000 : node21295;
															assign node21295 = (inp[10]) ? node21297 : 4'b0100;
																assign node21297 = (inp[12]) ? 4'b0000 : 4'b0100;
														assign node21301 = (inp[9]) ? 4'b0100 : node21302;
															assign node21302 = (inp[12]) ? 4'b0100 : 4'b0000;
												assign node21306 = (inp[3]) ? node21328 : node21307;
													assign node21307 = (inp[9]) ? node21319 : node21308;
														assign node21308 = (inp[4]) ? node21314 : node21309;
															assign node21309 = (inp[12]) ? node21311 : 4'b0100;
																assign node21311 = (inp[10]) ? 4'b0000 : 4'b0100;
															assign node21314 = (inp[12]) ? node21316 : 4'b0000;
																assign node21316 = (inp[10]) ? 4'b0110 : 4'b0000;
														assign node21319 = (inp[4]) ? node21323 : node21320;
															assign node21320 = (inp[10]) ? 4'b0110 : 4'b0000;
															assign node21323 = (inp[12]) ? node21325 : 4'b0110;
																assign node21325 = (inp[10]) ? 4'b0010 : 4'b0110;
													assign node21328 = (inp[9]) ? 4'b0010 : node21329;
														assign node21329 = (inp[4]) ? node21331 : 4'b0110;
															assign node21331 = (inp[12]) ? node21333 : 4'b0010;
																assign node21333 = (inp[10]) ? 4'b0110 : 4'b0010;
											assign node21337 = (inp[0]) ? node21367 : node21338;
												assign node21338 = (inp[3]) ? node21356 : node21339;
													assign node21339 = (inp[4]) ? node21351 : node21340;
														assign node21340 = (inp[9]) ? node21346 : node21341;
															assign node21341 = (inp[10]) ? node21343 : 4'b0100;
																assign node21343 = (inp[12]) ? 4'b0000 : 4'b0100;
															assign node21346 = (inp[10]) ? node21348 : 4'b0000;
																assign node21348 = (inp[12]) ? 4'b0110 : 4'b0000;
														assign node21351 = (inp[9]) ? 4'b0110 : node21352;
															assign node21352 = (inp[12]) ? 4'b0110 : 4'b0000;
													assign node21356 = (inp[9]) ? node21362 : node21357;
														assign node21357 = (inp[4]) ? 4'b0010 : node21358;
															assign node21358 = (inp[10]) ? 4'b0010 : 4'b0110;
														assign node21362 = (inp[4]) ? 4'b0110 : node21363;
															assign node21363 = (inp[12]) ? 4'b0110 : 4'b0010;
												assign node21367 = (inp[3]) ? node21383 : node21368;
													assign node21368 = (inp[9]) ? node21378 : node21369;
														assign node21369 = (inp[12]) ? node21373 : node21370;
															assign node21370 = (inp[4]) ? 4'b0010 : 4'b0110;
															assign node21373 = (inp[4]) ? node21375 : 4'b0010;
																assign node21375 = (inp[10]) ? 4'b0100 : 4'b0010;
														assign node21378 = (inp[4]) ? 4'b0100 : node21379;
															assign node21379 = (inp[12]) ? 4'b0100 : 4'b0010;
													assign node21383 = (inp[12]) ? node21391 : node21384;
														assign node21384 = (inp[9]) ? node21388 : node21385;
															assign node21385 = (inp[4]) ? 4'b0000 : 4'b0100;
															assign node21388 = (inp[4]) ? 4'b0100 : 4'b0000;
														assign node21391 = (inp[10]) ? node21399 : node21392;
															assign node21392 = (inp[9]) ? node21396 : node21393;
																assign node21393 = (inp[4]) ? 4'b0000 : 4'b0100;
																assign node21396 = (inp[4]) ? 4'b0100 : 4'b0000;
															assign node21399 = (inp[4]) ? node21401 : 4'b0000;
																assign node21401 = (inp[9]) ? 4'b0000 : 4'b0100;
								assign node21404 = (inp[12]) ? node21666 : node21405;
									assign node21405 = (inp[14]) ? node21555 : node21406;
										assign node21406 = (inp[5]) ? node21488 : node21407;
											assign node21407 = (inp[9]) ? node21447 : node21408;
												assign node21408 = (inp[4]) ? node21424 : node21409;
													assign node21409 = (inp[10]) ? node21417 : node21410;
														assign node21410 = (inp[0]) ? node21414 : node21411;
															assign node21411 = (inp[15]) ? 4'b0100 : 4'b0110;
															assign node21414 = (inp[15]) ? 4'b0110 : 4'b0100;
														assign node21417 = (inp[0]) ? node21421 : node21418;
															assign node21418 = (inp[15]) ? 4'b0100 : 4'b0110;
															assign node21421 = (inp[15]) ? 4'b0110 : 4'b0100;
													assign node21424 = (inp[3]) ? node21438 : node21425;
														assign node21425 = (inp[10]) ? node21433 : node21426;
															assign node21426 = (inp[0]) ? node21430 : node21427;
																assign node21427 = (inp[15]) ? 4'b0000 : 4'b0010;
																assign node21430 = (inp[15]) ? 4'b0010 : 4'b0000;
															assign node21433 = (inp[15]) ? node21435 : 4'b0000;
																assign node21435 = (inp[0]) ? 4'b0010 : 4'b0000;
														assign node21438 = (inp[10]) ? node21440 : 4'b0010;
															assign node21440 = (inp[15]) ? node21444 : node21441;
																assign node21441 = (inp[0]) ? 4'b0000 : 4'b0010;
																assign node21444 = (inp[0]) ? 4'b0010 : 4'b0000;
												assign node21447 = (inp[4]) ? node21471 : node21448;
													assign node21448 = (inp[10]) ? node21464 : node21449;
														assign node21449 = (inp[3]) ? node21457 : node21450;
															assign node21450 = (inp[0]) ? node21454 : node21451;
																assign node21451 = (inp[15]) ? 4'b0000 : 4'b0010;
																assign node21454 = (inp[15]) ? 4'b0010 : 4'b0000;
															assign node21457 = (inp[15]) ? node21461 : node21458;
																assign node21458 = (inp[0]) ? 4'b0000 : 4'b0010;
																assign node21461 = (inp[0]) ? 4'b0010 : 4'b0000;
														assign node21464 = (inp[0]) ? node21468 : node21465;
															assign node21465 = (inp[15]) ? 4'b0000 : 4'b0010;
															assign node21468 = (inp[15]) ? 4'b0010 : 4'b0000;
													assign node21471 = (inp[10]) ? node21481 : node21472;
														assign node21472 = (inp[15]) ? node21474 : 4'b0100;
															assign node21474 = (inp[3]) ? node21478 : node21475;
																assign node21475 = (inp[0]) ? 4'b0110 : 4'b0100;
																assign node21478 = (inp[0]) ? 4'b0100 : 4'b0110;
														assign node21481 = (inp[3]) ? node21483 : 4'b0110;
															assign node21483 = (inp[0]) ? node21485 : 4'b0110;
																assign node21485 = (inp[15]) ? 4'b0100 : 4'b0110;
											assign node21488 = (inp[0]) ? node21526 : node21489;
												assign node21489 = (inp[15]) ? node21507 : node21490;
													assign node21490 = (inp[3]) ? node21498 : node21491;
														assign node21491 = (inp[9]) ? node21495 : node21492;
															assign node21492 = (inp[4]) ? 4'b0010 : 4'b0110;
															assign node21495 = (inp[4]) ? 4'b0100 : 4'b0010;
														assign node21498 = (inp[10]) ? node21500 : 4'b0000;
															assign node21500 = (inp[4]) ? node21504 : node21501;
																assign node21501 = (inp[9]) ? 4'b0000 : 4'b0100;
																assign node21504 = (inp[9]) ? 4'b0100 : 4'b0000;
													assign node21507 = (inp[3]) ? node21515 : node21508;
														assign node21508 = (inp[9]) ? node21512 : node21509;
															assign node21509 = (inp[4]) ? 4'b0000 : 4'b0100;
															assign node21512 = (inp[4]) ? 4'b0110 : 4'b0000;
														assign node21515 = (inp[10]) ? node21521 : node21516;
															assign node21516 = (inp[4]) ? 4'b0010 : node21517;
																assign node21517 = (inp[9]) ? 4'b0010 : 4'b0110;
															assign node21521 = (inp[9]) ? node21523 : 4'b0110;
																assign node21523 = (inp[4]) ? 4'b0110 : 4'b0010;
												assign node21526 = (inp[15]) ? node21542 : node21527;
													assign node21527 = (inp[3]) ? node21535 : node21528;
														assign node21528 = (inp[4]) ? node21532 : node21529;
															assign node21529 = (inp[9]) ? 4'b0000 : 4'b0100;
															assign node21532 = (inp[9]) ? 4'b0110 : 4'b0000;
														assign node21535 = (inp[9]) ? node21539 : node21536;
															assign node21536 = (inp[4]) ? 4'b0010 : 4'b0110;
															assign node21539 = (inp[4]) ? 4'b0110 : 4'b0010;
													assign node21542 = (inp[3]) ? node21548 : node21543;
														assign node21543 = (inp[4]) ? node21545 : 4'b0010;
															assign node21545 = (inp[9]) ? 4'b0100 : 4'b0010;
														assign node21548 = (inp[4]) ? node21552 : node21549;
															assign node21549 = (inp[9]) ? 4'b0000 : 4'b0100;
															assign node21552 = (inp[9]) ? 4'b0100 : 4'b0000;
										assign node21555 = (inp[0]) ? node21607 : node21556;
											assign node21556 = (inp[15]) ? node21582 : node21557;
												assign node21557 = (inp[3]) ? node21567 : node21558;
													assign node21558 = (inp[9]) ? node21562 : node21559;
														assign node21559 = (inp[4]) ? 4'b0010 : 4'b0110;
														assign node21562 = (inp[4]) ? node21564 : 4'b0010;
															assign node21564 = (inp[5]) ? 4'b0100 : 4'b0110;
													assign node21567 = (inp[5]) ? node21575 : node21568;
														assign node21568 = (inp[4]) ? node21572 : node21569;
															assign node21569 = (inp[9]) ? 4'b0010 : 4'b0110;
															assign node21572 = (inp[9]) ? 4'b0100 : 4'b0010;
														assign node21575 = (inp[9]) ? node21579 : node21576;
															assign node21576 = (inp[4]) ? 4'b0000 : 4'b0100;
															assign node21579 = (inp[4]) ? 4'b0100 : 4'b0000;
												assign node21582 = (inp[3]) ? node21592 : node21583;
													assign node21583 = (inp[9]) ? node21587 : node21584;
														assign node21584 = (inp[4]) ? 4'b0000 : 4'b0100;
														assign node21587 = (inp[4]) ? node21589 : 4'b0000;
															assign node21589 = (inp[10]) ? 4'b0100 : 4'b0110;
													assign node21592 = (inp[5]) ? node21600 : node21593;
														assign node21593 = (inp[4]) ? node21597 : node21594;
															assign node21594 = (inp[9]) ? 4'b0000 : 4'b0100;
															assign node21597 = (inp[9]) ? 4'b0110 : 4'b0000;
														assign node21600 = (inp[4]) ? node21604 : node21601;
															assign node21601 = (inp[9]) ? 4'b0010 : 4'b0110;
															assign node21604 = (inp[9]) ? 4'b0110 : 4'b0010;
											assign node21607 = (inp[15]) ? node21637 : node21608;
												assign node21608 = (inp[3]) ? node21616 : node21609;
													assign node21609 = (inp[4]) ? node21613 : node21610;
														assign node21610 = (inp[9]) ? 4'b0000 : 4'b0100;
														assign node21613 = (inp[9]) ? 4'b0110 : 4'b0000;
													assign node21616 = (inp[5]) ? node21624 : node21617;
														assign node21617 = (inp[4]) ? node21621 : node21618;
															assign node21618 = (inp[9]) ? 4'b0000 : 4'b0100;
															assign node21621 = (inp[9]) ? 4'b0110 : 4'b0000;
														assign node21624 = (inp[10]) ? node21632 : node21625;
															assign node21625 = (inp[4]) ? node21629 : node21626;
																assign node21626 = (inp[9]) ? 4'b0010 : 4'b0110;
																assign node21629 = (inp[9]) ? 4'b0110 : 4'b0010;
															assign node21632 = (inp[4]) ? node21634 : 4'b0110;
																assign node21634 = (inp[9]) ? 4'b0110 : 4'b0010;
												assign node21637 = (inp[3]) ? node21647 : node21638;
													assign node21638 = (inp[4]) ? node21642 : node21639;
														assign node21639 = (inp[9]) ? 4'b0010 : 4'b0110;
														assign node21642 = (inp[9]) ? node21644 : 4'b0010;
															assign node21644 = (inp[5]) ? 4'b0100 : 4'b0110;
													assign node21647 = (inp[5]) ? node21653 : node21648;
														assign node21648 = (inp[4]) ? 4'b0100 : node21649;
															assign node21649 = (inp[9]) ? 4'b0010 : 4'b0110;
														assign node21653 = (inp[10]) ? node21661 : node21654;
															assign node21654 = (inp[9]) ? node21658 : node21655;
																assign node21655 = (inp[4]) ? 4'b0000 : 4'b0100;
																assign node21658 = (inp[4]) ? 4'b0100 : 4'b0000;
															assign node21661 = (inp[9]) ? node21663 : 4'b0100;
																assign node21663 = (inp[4]) ? 4'b0100 : 4'b0000;
									assign node21666 = (inp[4]) ? node21752 : node21667;
										assign node21667 = (inp[9]) ? node21709 : node21668;
											assign node21668 = (inp[10]) ? node21688 : node21669;
												assign node21669 = (inp[15]) ? node21677 : node21670;
													assign node21670 = (inp[0]) ? 4'b0100 : node21671;
														assign node21671 = (inp[14]) ? 4'b0110 : node21672;
															assign node21672 = (inp[3]) ? 4'b0100 : 4'b0110;
													assign node21677 = (inp[0]) ? node21683 : node21678;
														assign node21678 = (inp[3]) ? node21680 : 4'b0100;
															assign node21680 = (inp[5]) ? 4'b0110 : 4'b0100;
														assign node21683 = (inp[3]) ? node21685 : 4'b0110;
															assign node21685 = (inp[5]) ? 4'b0100 : 4'b0110;
												assign node21688 = (inp[0]) ? node21700 : node21689;
													assign node21689 = (inp[15]) ? node21695 : node21690;
														assign node21690 = (inp[3]) ? node21692 : 4'b0010;
															assign node21692 = (inp[5]) ? 4'b0000 : 4'b0010;
														assign node21695 = (inp[5]) ? node21697 : 4'b0000;
															assign node21697 = (inp[3]) ? 4'b0010 : 4'b0000;
													assign node21700 = (inp[15]) ? node21706 : node21701;
														assign node21701 = (inp[3]) ? node21703 : 4'b0000;
															assign node21703 = (inp[5]) ? 4'b0010 : 4'b0000;
														assign node21706 = (inp[3]) ? 4'b0000 : 4'b0010;
											assign node21709 = (inp[10]) ? node21729 : node21710;
												assign node21710 = (inp[15]) ? node21718 : node21711;
													assign node21711 = (inp[0]) ? node21713 : 4'b0010;
														assign node21713 = (inp[3]) ? node21715 : 4'b0000;
															assign node21715 = (inp[5]) ? 4'b0010 : 4'b0000;
													assign node21718 = (inp[0]) ? node21724 : node21719;
														assign node21719 = (inp[5]) ? node21721 : 4'b0000;
															assign node21721 = (inp[3]) ? 4'b0010 : 4'b0000;
														assign node21724 = (inp[3]) ? node21726 : 4'b0010;
															assign node21726 = (inp[5]) ? 4'b0000 : 4'b0010;
												assign node21729 = (inp[5]) ? node21745 : node21730;
													assign node21730 = (inp[3]) ? node21738 : node21731;
														assign node21731 = (inp[0]) ? node21735 : node21732;
															assign node21732 = (inp[15]) ? 4'b0100 : 4'b0110;
															assign node21735 = (inp[15]) ? 4'b0110 : 4'b0100;
														assign node21738 = (inp[0]) ? node21742 : node21739;
															assign node21739 = (inp[15]) ? 4'b0110 : 4'b0100;
															assign node21742 = (inp[15]) ? 4'b0100 : 4'b0110;
													assign node21745 = (inp[14]) ? node21747 : 4'b0110;
														assign node21747 = (inp[15]) ? 4'b0110 : node21748;
															assign node21748 = (inp[0]) ? 4'b0110 : 4'b0100;
										assign node21752 = (inp[15]) ? node21820 : node21753;
											assign node21753 = (inp[0]) ? node21781 : node21754;
												assign node21754 = (inp[5]) ? node21766 : node21755;
													assign node21755 = (inp[3]) ? node21763 : node21756;
														assign node21756 = (inp[9]) ? node21760 : node21757;
															assign node21757 = (inp[10]) ? 4'b0110 : 4'b0010;
															assign node21760 = (inp[10]) ? 4'b0010 : 4'b0110;
														assign node21763 = (inp[9]) ? 4'b0100 : 4'b0010;
													assign node21766 = (inp[3]) ? node21774 : node21767;
														assign node21767 = (inp[9]) ? node21771 : node21768;
															assign node21768 = (inp[10]) ? 4'b0100 : 4'b0010;
															assign node21771 = (inp[10]) ? 4'b0000 : 4'b0100;
														assign node21774 = (inp[9]) ? node21778 : node21775;
															assign node21775 = (inp[10]) ? 4'b0100 : 4'b0000;
															assign node21778 = (inp[10]) ? 4'b0000 : 4'b0100;
												assign node21781 = (inp[3]) ? node21801 : node21782;
													assign node21782 = (inp[5]) ? node21794 : node21783;
														assign node21783 = (inp[14]) ? node21789 : node21784;
															assign node21784 = (inp[9]) ? 4'b0100 : node21785;
																assign node21785 = (inp[10]) ? 4'b0100 : 4'b0000;
															assign node21789 = (inp[9]) ? node21791 : 4'b0100;
																assign node21791 = (inp[10]) ? 4'b0000 : 4'b0100;
														assign node21794 = (inp[9]) ? node21798 : node21795;
															assign node21795 = (inp[10]) ? 4'b0110 : 4'b0000;
															assign node21798 = (inp[10]) ? 4'b0010 : 4'b0110;
													assign node21801 = (inp[5]) ? node21807 : node21802;
														assign node21802 = (inp[9]) ? node21804 : 4'b0110;
															assign node21804 = (inp[10]) ? 4'b0010 : 4'b0110;
														assign node21807 = (inp[14]) ? node21815 : node21808;
															assign node21808 = (inp[10]) ? node21812 : node21809;
																assign node21809 = (inp[9]) ? 4'b0110 : 4'b0010;
																assign node21812 = (inp[9]) ? 4'b0010 : 4'b0110;
															assign node21815 = (inp[9]) ? 4'b0010 : node21816;
																assign node21816 = (inp[10]) ? 4'b0110 : 4'b0010;
											assign node21820 = (inp[0]) ? node21844 : node21821;
												assign node21821 = (inp[5]) ? node21835 : node21822;
													assign node21822 = (inp[3]) ? node21828 : node21823;
														assign node21823 = (inp[10]) ? 4'b0000 : node21824;
															assign node21824 = (inp[9]) ? 4'b0100 : 4'b0000;
														assign node21828 = (inp[9]) ? node21832 : node21829;
															assign node21829 = (inp[10]) ? 4'b0110 : 4'b0000;
															assign node21832 = (inp[10]) ? 4'b0010 : 4'b0110;
													assign node21835 = (inp[10]) ? node21841 : node21836;
														assign node21836 = (inp[9]) ? 4'b0110 : node21837;
															assign node21837 = (inp[14]) ? 4'b0000 : 4'b0010;
														assign node21841 = (inp[9]) ? 4'b0010 : 4'b0110;
												assign node21844 = (inp[5]) ? node21860 : node21845;
													assign node21845 = (inp[3]) ? node21853 : node21846;
														assign node21846 = (inp[9]) ? node21850 : node21847;
															assign node21847 = (inp[10]) ? 4'b0110 : 4'b0010;
															assign node21850 = (inp[10]) ? 4'b0010 : 4'b0110;
														assign node21853 = (inp[9]) ? node21857 : node21854;
															assign node21854 = (inp[10]) ? 4'b0100 : 4'b0010;
															assign node21857 = (inp[10]) ? 4'b0000 : 4'b0100;
													assign node21860 = (inp[9]) ? node21866 : node21861;
														assign node21861 = (inp[10]) ? 4'b0100 : node21862;
															assign node21862 = (inp[3]) ? 4'b0000 : 4'b0010;
														assign node21866 = (inp[10]) ? 4'b0000 : 4'b0100;
							assign node21869 = (inp[2]) ? node22459 : node21870;
								assign node21870 = (inp[14]) ? node22152 : node21871;
									assign node21871 = (inp[10]) ? node21983 : node21872;
										assign node21872 = (inp[5]) ? node21908 : node21873;
											assign node21873 = (inp[9]) ? node21889 : node21874;
												assign node21874 = (inp[4]) ? node21882 : node21875;
													assign node21875 = (inp[15]) ? node21879 : node21876;
														assign node21876 = (inp[0]) ? 4'b0100 : 4'b0110;
														assign node21879 = (inp[0]) ? 4'b0110 : 4'b0100;
													assign node21882 = (inp[0]) ? node21886 : node21883;
														assign node21883 = (inp[15]) ? 4'b0000 : 4'b0010;
														assign node21886 = (inp[15]) ? 4'b0010 : 4'b0000;
												assign node21889 = (inp[4]) ? node21897 : node21890;
													assign node21890 = (inp[0]) ? node21894 : node21891;
														assign node21891 = (inp[15]) ? 4'b0000 : 4'b0010;
														assign node21894 = (inp[15]) ? 4'b0010 : 4'b0000;
													assign node21897 = (inp[0]) ? 4'b0110 : node21898;
														assign node21898 = (inp[12]) ? node21900 : 4'b0110;
															assign node21900 = (inp[3]) ? node21904 : node21901;
																assign node21901 = (inp[15]) ? 4'b0100 : 4'b0110;
																assign node21904 = (inp[15]) ? 4'b0110 : 4'b0100;
											assign node21908 = (inp[9]) ? node21948 : node21909;
												assign node21909 = (inp[4]) ? node21929 : node21910;
													assign node21910 = (inp[3]) ? node21916 : node21911;
														assign node21911 = (inp[15]) ? 4'b0110 : node21912;
															assign node21912 = (inp[0]) ? 4'b0100 : 4'b0110;
														assign node21916 = (inp[12]) ? node21924 : node21917;
															assign node21917 = (inp[0]) ? node21921 : node21918;
																assign node21918 = (inp[15]) ? 4'b0110 : 4'b0100;
																assign node21921 = (inp[15]) ? 4'b0100 : 4'b0110;
															assign node21924 = (inp[15]) ? 4'b0110 : node21925;
																assign node21925 = (inp[0]) ? 4'b0110 : 4'b0100;
													assign node21929 = (inp[0]) ? node21941 : node21930;
														assign node21930 = (inp[12]) ? node21936 : node21931;
															assign node21931 = (inp[15]) ? node21933 : 4'b0010;
																assign node21933 = (inp[3]) ? 4'b0010 : 4'b0000;
															assign node21936 = (inp[3]) ? node21938 : 4'b0010;
																assign node21938 = (inp[15]) ? 4'b0010 : 4'b0000;
														assign node21941 = (inp[15]) ? node21945 : node21942;
															assign node21942 = (inp[3]) ? 4'b0010 : 4'b0000;
															assign node21945 = (inp[3]) ? 4'b0000 : 4'b0010;
												assign node21948 = (inp[4]) ? node21976 : node21949;
													assign node21949 = (inp[15]) ? node21965 : node21950;
														assign node21950 = (inp[12]) ? node21958 : node21951;
															assign node21951 = (inp[0]) ? node21955 : node21952;
																assign node21952 = (inp[3]) ? 4'b0000 : 4'b0010;
																assign node21955 = (inp[3]) ? 4'b0010 : 4'b0000;
															assign node21958 = (inp[3]) ? node21962 : node21959;
																assign node21959 = (inp[0]) ? 4'b0000 : 4'b0010;
																assign node21962 = (inp[0]) ? 4'b0010 : 4'b0000;
														assign node21965 = (inp[12]) ? node21971 : node21966;
															assign node21966 = (inp[0]) ? node21968 : 4'b0000;
																assign node21968 = (inp[3]) ? 4'b0000 : 4'b0010;
															assign node21971 = (inp[3]) ? node21973 : 4'b0000;
																assign node21973 = (inp[0]) ? 4'b0000 : 4'b0010;
													assign node21976 = (inp[15]) ? node21980 : node21977;
														assign node21977 = (inp[0]) ? 4'b0110 : 4'b0100;
														assign node21980 = (inp[0]) ? 4'b0100 : 4'b0110;
										assign node21983 = (inp[3]) ? node22069 : node21984;
											assign node21984 = (inp[9]) ? node22018 : node21985;
												assign node21985 = (inp[0]) ? node22005 : node21986;
													assign node21986 = (inp[15]) ? node21996 : node21987;
														assign node21987 = (inp[12]) ? node21991 : node21988;
															assign node21988 = (inp[4]) ? 4'b0010 : 4'b0110;
															assign node21991 = (inp[4]) ? node21993 : 4'b0010;
																assign node21993 = (inp[5]) ? 4'b0100 : 4'b0110;
														assign node21996 = (inp[12]) ? node22000 : node21997;
															assign node21997 = (inp[4]) ? 4'b0000 : 4'b0100;
															assign node22000 = (inp[4]) ? node22002 : 4'b0000;
																assign node22002 = (inp[5]) ? 4'b0110 : 4'b0100;
													assign node22005 = (inp[15]) ? node22015 : node22006;
														assign node22006 = (inp[12]) ? node22010 : node22007;
															assign node22007 = (inp[4]) ? 4'b0000 : 4'b0100;
															assign node22010 = (inp[4]) ? node22012 : 4'b0000;
																assign node22012 = (inp[5]) ? 4'b0110 : 4'b0100;
														assign node22015 = (inp[12]) ? 4'b0100 : 4'b0110;
												assign node22018 = (inp[12]) ? node22046 : node22019;
													assign node22019 = (inp[4]) ? node22033 : node22020;
														assign node22020 = (inp[5]) ? node22028 : node22021;
															assign node22021 = (inp[0]) ? node22025 : node22022;
																assign node22022 = (inp[15]) ? 4'b0000 : 4'b0010;
																assign node22025 = (inp[15]) ? 4'b0010 : 4'b0000;
															assign node22028 = (inp[15]) ? 4'b0010 : node22029;
																assign node22029 = (inp[0]) ? 4'b0000 : 4'b0010;
														assign node22033 = (inp[15]) ? node22041 : node22034;
															assign node22034 = (inp[5]) ? node22038 : node22035;
																assign node22035 = (inp[0]) ? 4'b0100 : 4'b0110;
																assign node22038 = (inp[0]) ? 4'b0110 : 4'b0100;
															assign node22041 = (inp[5]) ? node22043 : 4'b0100;
																assign node22043 = (inp[0]) ? 4'b0100 : 4'b0110;
													assign node22046 = (inp[4]) ? node22062 : node22047;
														assign node22047 = (inp[5]) ? node22055 : node22048;
															assign node22048 = (inp[15]) ? node22052 : node22049;
																assign node22049 = (inp[0]) ? 4'b0100 : 4'b0110;
																assign node22052 = (inp[0]) ? 4'b0110 : 4'b0100;
															assign node22055 = (inp[15]) ? node22059 : node22056;
																assign node22056 = (inp[0]) ? 4'b0110 : 4'b0100;
																assign node22059 = (inp[0]) ? 4'b0100 : 4'b0110;
														assign node22062 = (inp[5]) ? node22064 : 4'b0010;
															assign node22064 = (inp[15]) ? node22066 : 4'b0010;
																assign node22066 = (inp[0]) ? 4'b0000 : 4'b0010;
											assign node22069 = (inp[12]) ? node22111 : node22070;
												assign node22070 = (inp[15]) ? node22088 : node22071;
													assign node22071 = (inp[5]) ? node22081 : node22072;
														assign node22072 = (inp[0]) ? node22076 : node22073;
															assign node22073 = (inp[4]) ? 4'b0010 : 4'b0110;
															assign node22076 = (inp[9]) ? node22078 : 4'b0000;
																assign node22078 = (inp[4]) ? 4'b0110 : 4'b0000;
														assign node22081 = (inp[9]) ? node22085 : node22082;
															assign node22082 = (inp[4]) ? 4'b0010 : 4'b0110;
															assign node22085 = (inp[4]) ? 4'b0110 : 4'b0010;
													assign node22088 = (inp[4]) ? node22104 : node22089;
														assign node22089 = (inp[9]) ? node22097 : node22090;
															assign node22090 = (inp[5]) ? node22094 : node22091;
																assign node22091 = (inp[0]) ? 4'b0110 : 4'b0100;
																assign node22094 = (inp[0]) ? 4'b0100 : 4'b0110;
															assign node22097 = (inp[0]) ? node22101 : node22098;
																assign node22098 = (inp[5]) ? 4'b0010 : 4'b0000;
																assign node22101 = (inp[5]) ? 4'b0000 : 4'b0010;
														assign node22104 = (inp[9]) ? node22108 : node22105;
															assign node22105 = (inp[0]) ? 4'b0010 : 4'b0000;
															assign node22108 = (inp[0]) ? 4'b0100 : 4'b0110;
												assign node22111 = (inp[4]) ? node22133 : node22112;
													assign node22112 = (inp[9]) ? node22126 : node22113;
														assign node22113 = (inp[5]) ? node22119 : node22114;
															assign node22114 = (inp[0]) ? node22116 : 4'b0010;
																assign node22116 = (inp[15]) ? 4'b0010 : 4'b0000;
															assign node22119 = (inp[15]) ? node22123 : node22120;
																assign node22120 = (inp[0]) ? 4'b0010 : 4'b0000;
																assign node22123 = (inp[0]) ? 4'b0000 : 4'b0010;
														assign node22126 = (inp[15]) ? node22130 : node22127;
															assign node22127 = (inp[0]) ? 4'b0110 : 4'b0100;
															assign node22130 = (inp[0]) ? 4'b0100 : 4'b0110;
													assign node22133 = (inp[9]) ? node22145 : node22134;
														assign node22134 = (inp[5]) ? node22140 : node22135;
															assign node22135 = (inp[15]) ? node22137 : 4'b0100;
																assign node22137 = (inp[0]) ? 4'b0100 : 4'b0110;
															assign node22140 = (inp[0]) ? node22142 : 4'b0100;
																assign node22142 = (inp[15]) ? 4'b0100 : 4'b0110;
														assign node22145 = (inp[0]) ? node22149 : node22146;
															assign node22146 = (inp[15]) ? 4'b0010 : 4'b0000;
															assign node22149 = (inp[15]) ? 4'b0000 : 4'b0010;
									assign node22152 = (inp[12]) ? node22308 : node22153;
										assign node22153 = (inp[5]) ? node22223 : node22154;
											assign node22154 = (inp[9]) ? node22190 : node22155;
												assign node22155 = (inp[0]) ? node22173 : node22156;
													assign node22156 = (inp[15]) ? node22166 : node22157;
														assign node22157 = (inp[10]) ? node22161 : node22158;
															assign node22158 = (inp[4]) ? 4'b1011 : 4'b1111;
															assign node22161 = (inp[4]) ? node22163 : 4'b1011;
																assign node22163 = (inp[3]) ? 4'b1101 : 4'b1111;
														assign node22166 = (inp[10]) ? node22168 : 4'b1001;
															assign node22168 = (inp[4]) ? node22170 : 4'b1001;
																assign node22170 = (inp[3]) ? 4'b1111 : 4'b1101;
													assign node22173 = (inp[15]) ? node22183 : node22174;
														assign node22174 = (inp[4]) ? node22178 : node22175;
															assign node22175 = (inp[10]) ? 4'b1001 : 4'b1101;
															assign node22178 = (inp[3]) ? 4'b1111 : node22179;
																assign node22179 = (inp[10]) ? 4'b1101 : 4'b1001;
														assign node22183 = (inp[3]) ? node22185 : 4'b1111;
															assign node22185 = (inp[4]) ? 4'b1011 : node22186;
																assign node22186 = (inp[10]) ? 4'b1011 : 4'b1111;
												assign node22190 = (inp[10]) ? node22214 : node22191;
													assign node22191 = (inp[4]) ? node22201 : node22192;
														assign node22192 = (inp[3]) ? node22198 : node22193;
															assign node22193 = (inp[15]) ? node22195 : 4'b1011;
																assign node22195 = (inp[0]) ? 4'b1011 : 4'b1001;
															assign node22198 = (inp[15]) ? 4'b1011 : 4'b1001;
														assign node22201 = (inp[3]) ? node22207 : node22202;
															assign node22202 = (inp[0]) ? 4'b1111 : node22203;
																assign node22203 = (inp[15]) ? 4'b1101 : 4'b1111;
															assign node22207 = (inp[0]) ? node22211 : node22208;
																assign node22208 = (inp[15]) ? 4'b1111 : 4'b1101;
																assign node22211 = (inp[15]) ? 4'b1101 : 4'b1111;
													assign node22214 = (inp[4]) ? 4'b1011 : node22215;
														assign node22215 = (inp[0]) ? node22217 : 4'b1111;
															assign node22217 = (inp[3]) ? node22219 : 4'b1101;
																assign node22219 = (inp[15]) ? 4'b1101 : 4'b1111;
											assign node22223 = (inp[10]) ? node22261 : node22224;
												assign node22224 = (inp[15]) ? node22246 : node22225;
													assign node22225 = (inp[0]) ? node22235 : node22226;
														assign node22226 = (inp[3]) ? node22230 : node22227;
															assign node22227 = (inp[4]) ? 4'b1101 : 4'b1111;
															assign node22230 = (inp[4]) ? node22232 : 4'b1001;
																assign node22232 = (inp[9]) ? 4'b1101 : 4'b1001;
														assign node22235 = (inp[3]) ? node22241 : node22236;
															assign node22236 = (inp[4]) ? node22238 : 4'b1001;
																assign node22238 = (inp[9]) ? 4'b1111 : 4'b1001;
															assign node22241 = (inp[4]) ? 4'b1011 : node22242;
																assign node22242 = (inp[9]) ? 4'b1011 : 4'b1111;
													assign node22246 = (inp[0]) ? node22258 : node22247;
														assign node22247 = (inp[3]) ? node22253 : node22248;
															assign node22248 = (inp[4]) ? 4'b1111 : node22249;
																assign node22249 = (inp[9]) ? 4'b1001 : 4'b1101;
															assign node22253 = (inp[4]) ? 4'b1111 : node22254;
																assign node22254 = (inp[9]) ? 4'b1011 : 4'b1111;
														assign node22258 = (inp[9]) ? 4'b1101 : 4'b1111;
												assign node22261 = (inp[4]) ? node22287 : node22262;
													assign node22262 = (inp[9]) ? node22276 : node22263;
														assign node22263 = (inp[15]) ? node22269 : node22264;
															assign node22264 = (inp[3]) ? node22266 : 4'b1001;
																assign node22266 = (inp[0]) ? 4'b1011 : 4'b1001;
															assign node22269 = (inp[3]) ? node22273 : node22270;
																assign node22270 = (inp[0]) ? 4'b1011 : 4'b1001;
																assign node22273 = (inp[0]) ? 4'b1001 : 4'b1011;
														assign node22276 = (inp[3]) ? node22282 : node22277;
															assign node22277 = (inp[15]) ? node22279 : 4'b1111;
																assign node22279 = (inp[0]) ? 4'b1101 : 4'b1111;
															assign node22282 = (inp[15]) ? node22284 : 4'b1101;
																assign node22284 = (inp[0]) ? 4'b1101 : 4'b1111;
													assign node22287 = (inp[9]) ? node22293 : node22288;
														assign node22288 = (inp[15]) ? node22290 : 4'b1111;
															assign node22290 = (inp[0]) ? 4'b1101 : 4'b1111;
														assign node22293 = (inp[3]) ? node22301 : node22294;
															assign node22294 = (inp[0]) ? node22298 : node22295;
																assign node22295 = (inp[15]) ? 4'b1011 : 4'b1001;
																assign node22298 = (inp[15]) ? 4'b1001 : 4'b1011;
															assign node22301 = (inp[15]) ? node22305 : node22302;
																assign node22302 = (inp[0]) ? 4'b1011 : 4'b1001;
																assign node22305 = (inp[0]) ? 4'b1001 : 4'b1011;
										assign node22308 = (inp[10]) ? node22376 : node22309;
											assign node22309 = (inp[4]) ? node22345 : node22310;
												assign node22310 = (inp[9]) ? node22330 : node22311;
													assign node22311 = (inp[3]) ? node22319 : node22312;
														assign node22312 = (inp[15]) ? node22316 : node22313;
															assign node22313 = (inp[0]) ? 4'b1001 : 4'b1011;
															assign node22316 = (inp[0]) ? 4'b1011 : 4'b1001;
														assign node22319 = (inp[5]) ? node22325 : node22320;
															assign node22320 = (inp[0]) ? 4'b1001 : node22321;
																assign node22321 = (inp[15]) ? 4'b1001 : 4'b1011;
															assign node22325 = (inp[0]) ? 4'b1011 : node22326;
																assign node22326 = (inp[15]) ? 4'b1011 : 4'b1001;
													assign node22330 = (inp[3]) ? node22338 : node22331;
														assign node22331 = (inp[0]) ? 4'b1101 : node22332;
															assign node22332 = (inp[5]) ? 4'b1101 : node22333;
																assign node22333 = (inp[15]) ? 4'b1101 : 4'b1111;
														assign node22338 = (inp[15]) ? node22342 : node22339;
															assign node22339 = (inp[0]) ? 4'b1111 : 4'b1101;
															assign node22342 = (inp[0]) ? 4'b1101 : 4'b1111;
												assign node22345 = (inp[9]) ? node22359 : node22346;
													assign node22346 = (inp[15]) ? node22354 : node22347;
														assign node22347 = (inp[0]) ? node22351 : node22348;
															assign node22348 = (inp[3]) ? 4'b1101 : 4'b1111;
															assign node22351 = (inp[5]) ? 4'b1111 : 4'b1101;
														assign node22354 = (inp[3]) ? 4'b1111 : node22355;
															assign node22355 = (inp[0]) ? 4'b1111 : 4'b1101;
													assign node22359 = (inp[0]) ? node22369 : node22360;
														assign node22360 = (inp[15]) ? node22366 : node22361;
															assign node22361 = (inp[3]) ? 4'b1001 : node22362;
																assign node22362 = (inp[5]) ? 4'b1001 : 4'b1011;
															assign node22366 = (inp[3]) ? 4'b1011 : 4'b1001;
														assign node22369 = (inp[15]) ? node22371 : 4'b1011;
															assign node22371 = (inp[5]) ? 4'b1001 : node22372;
																assign node22372 = (inp[3]) ? 4'b1001 : 4'b1011;
											assign node22376 = (inp[3]) ? node22426 : node22377;
												assign node22377 = (inp[5]) ? node22403 : node22378;
													assign node22378 = (inp[4]) ? node22390 : node22379;
														assign node22379 = (inp[9]) ? node22383 : node22380;
															assign node22380 = (inp[0]) ? 4'b1001 : 4'b1011;
															assign node22383 = (inp[0]) ? node22387 : node22384;
																assign node22384 = (inp[15]) ? 4'b1101 : 4'b1111;
																assign node22387 = (inp[15]) ? 4'b1111 : 4'b1101;
														assign node22390 = (inp[9]) ? node22396 : node22391;
															assign node22391 = (inp[0]) ? 4'b1101 : node22392;
																assign node22392 = (inp[15]) ? 4'b1101 : 4'b1111;
															assign node22396 = (inp[15]) ? node22400 : node22397;
																assign node22397 = (inp[0]) ? 4'b1001 : 4'b1011;
																assign node22400 = (inp[0]) ? 4'b1011 : 4'b1001;
													assign node22403 = (inp[0]) ? node22417 : node22404;
														assign node22404 = (inp[15]) ? node22410 : node22405;
															assign node22405 = (inp[4]) ? node22407 : 4'b1011;
																assign node22407 = (inp[9]) ? 4'b1001 : 4'b1101;
															assign node22410 = (inp[4]) ? node22414 : node22411;
																assign node22411 = (inp[9]) ? 4'b1111 : 4'b1001;
																assign node22414 = (inp[9]) ? 4'b1011 : 4'b1111;
														assign node22417 = (inp[15]) ? 4'b1011 : node22418;
															assign node22418 = (inp[9]) ? node22422 : node22419;
																assign node22419 = (inp[4]) ? 4'b1111 : 4'b1001;
																assign node22422 = (inp[4]) ? 4'b1011 : 4'b1111;
												assign node22426 = (inp[0]) ? node22444 : node22427;
													assign node22427 = (inp[15]) ? node22439 : node22428;
														assign node22428 = (inp[5]) ? node22434 : node22429;
															assign node22429 = (inp[4]) ? 4'b1101 : node22430;
																assign node22430 = (inp[9]) ? 4'b1101 : 4'b1011;
															assign node22434 = (inp[4]) ? node22436 : 4'b1101;
																assign node22436 = (inp[9]) ? 4'b1001 : 4'b1101;
														assign node22439 = (inp[4]) ? node22441 : 4'b1111;
															assign node22441 = (inp[9]) ? 4'b1011 : 4'b1111;
													assign node22444 = (inp[15]) ? node22452 : node22445;
														assign node22445 = (inp[5]) ? 4'b1111 : node22446;
															assign node22446 = (inp[9]) ? node22448 : 4'b1001;
																assign node22448 = (inp[4]) ? 4'b1011 : 4'b1111;
														assign node22452 = (inp[9]) ? node22456 : node22453;
															assign node22453 = (inp[4]) ? 4'b1101 : 4'b1001;
															assign node22456 = (inp[4]) ? 4'b1001 : 4'b1101;
								assign node22459 = (inp[9]) ? node22639 : node22460;
									assign node22460 = (inp[4]) ? node22546 : node22461;
										assign node22461 = (inp[12]) ? node22523 : node22462;
											assign node22462 = (inp[10]) ? node22482 : node22463;
												assign node22463 = (inp[15]) ? node22473 : node22464;
													assign node22464 = (inp[0]) ? node22468 : node22465;
														assign node22465 = (inp[3]) ? 4'b1101 : 4'b1111;
														assign node22468 = (inp[5]) ? node22470 : 4'b1101;
															assign node22470 = (inp[3]) ? 4'b1111 : 4'b1101;
													assign node22473 = (inp[0]) ? node22477 : node22474;
														assign node22474 = (inp[3]) ? 4'b1111 : 4'b1101;
														assign node22477 = (inp[5]) ? node22479 : 4'b1111;
															assign node22479 = (inp[3]) ? 4'b1101 : 4'b1111;
												assign node22482 = (inp[3]) ? node22502 : node22483;
													assign node22483 = (inp[14]) ? node22489 : node22484;
														assign node22484 = (inp[0]) ? 4'b1001 : node22485;
															assign node22485 = (inp[5]) ? 4'b1011 : 4'b1001;
														assign node22489 = (inp[5]) ? node22495 : node22490;
															assign node22490 = (inp[15]) ? node22492 : 4'b1011;
																assign node22492 = (inp[0]) ? 4'b1011 : 4'b1001;
															assign node22495 = (inp[15]) ? node22499 : node22496;
																assign node22496 = (inp[0]) ? 4'b1001 : 4'b1011;
																assign node22499 = (inp[0]) ? 4'b1011 : 4'b1001;
													assign node22502 = (inp[14]) ? node22516 : node22503;
														assign node22503 = (inp[5]) ? node22509 : node22504;
															assign node22504 = (inp[15]) ? 4'b1011 : node22505;
																assign node22505 = (inp[0]) ? 4'b1001 : 4'b1011;
															assign node22509 = (inp[0]) ? node22513 : node22510;
																assign node22510 = (inp[15]) ? 4'b1011 : 4'b1001;
																assign node22513 = (inp[15]) ? 4'b1001 : 4'b1011;
														assign node22516 = (inp[0]) ? 4'b1011 : node22517;
															assign node22517 = (inp[15]) ? node22519 : 4'b1011;
																assign node22519 = (inp[5]) ? 4'b1011 : 4'b1001;
											assign node22523 = (inp[0]) ? node22535 : node22524;
												assign node22524 = (inp[15]) ? node22530 : node22525;
													assign node22525 = (inp[5]) ? node22527 : 4'b1011;
														assign node22527 = (inp[3]) ? 4'b1001 : 4'b1011;
													assign node22530 = (inp[5]) ? node22532 : 4'b1001;
														assign node22532 = (inp[3]) ? 4'b1011 : 4'b1001;
												assign node22535 = (inp[15]) ? node22541 : node22536;
													assign node22536 = (inp[3]) ? node22538 : 4'b1001;
														assign node22538 = (inp[5]) ? 4'b1011 : 4'b1001;
													assign node22541 = (inp[3]) ? node22543 : 4'b1011;
														assign node22543 = (inp[5]) ? 4'b1001 : 4'b1011;
										assign node22546 = (inp[10]) ? node22618 : node22547;
											assign node22547 = (inp[12]) ? node22585 : node22548;
												assign node22548 = (inp[5]) ? node22558 : node22549;
													assign node22549 = (inp[3]) ? node22551 : 4'b1001;
														assign node22551 = (inp[15]) ? node22555 : node22552;
															assign node22552 = (inp[0]) ? 4'b1001 : 4'b1011;
															assign node22555 = (inp[0]) ? 4'b1011 : 4'b1001;
													assign node22558 = (inp[14]) ? node22572 : node22559;
														assign node22559 = (inp[15]) ? node22567 : node22560;
															assign node22560 = (inp[0]) ? node22564 : node22561;
																assign node22561 = (inp[3]) ? 4'b1001 : 4'b1011;
																assign node22564 = (inp[3]) ? 4'b1011 : 4'b1001;
															assign node22567 = (inp[3]) ? node22569 : 4'b1001;
																assign node22569 = (inp[0]) ? 4'b1001 : 4'b1011;
														assign node22572 = (inp[3]) ? node22578 : node22573;
															assign node22573 = (inp[0]) ? node22575 : 4'b1011;
																assign node22575 = (inp[15]) ? 4'b1011 : 4'b1001;
															assign node22578 = (inp[15]) ? node22582 : node22579;
																assign node22579 = (inp[0]) ? 4'b1011 : 4'b1001;
																assign node22582 = (inp[0]) ? 4'b1001 : 4'b1011;
												assign node22585 = (inp[14]) ? node22601 : node22586;
													assign node22586 = (inp[3]) ? node22594 : node22587;
														assign node22587 = (inp[0]) ? node22589 : 4'b1111;
															assign node22589 = (inp[5]) ? 4'b1111 : node22590;
																assign node22590 = (inp[15]) ? 4'b1111 : 4'b1101;
														assign node22594 = (inp[0]) ? node22598 : node22595;
															assign node22595 = (inp[15]) ? 4'b1111 : 4'b1101;
															assign node22598 = (inp[15]) ? 4'b1101 : 4'b1111;
													assign node22601 = (inp[15]) ? node22607 : node22602;
														assign node22602 = (inp[0]) ? node22604 : 4'b1101;
															assign node22604 = (inp[5]) ? 4'b1111 : 4'b1101;
														assign node22607 = (inp[0]) ? node22613 : node22608;
															assign node22608 = (inp[5]) ? 4'b1111 : node22609;
																assign node22609 = (inp[3]) ? 4'b1111 : 4'b1101;
															assign node22613 = (inp[5]) ? 4'b1101 : node22614;
																assign node22614 = (inp[3]) ? 4'b1101 : 4'b1111;
											assign node22618 = (inp[0]) ? node22628 : node22619;
												assign node22619 = (inp[15]) ? node22625 : node22620;
													assign node22620 = (inp[5]) ? 4'b1101 : node22621;
														assign node22621 = (inp[3]) ? 4'b1101 : 4'b1111;
													assign node22625 = (inp[3]) ? 4'b1111 : 4'b1101;
												assign node22628 = (inp[15]) ? node22634 : node22629;
													assign node22629 = (inp[5]) ? 4'b1111 : node22630;
														assign node22630 = (inp[3]) ? 4'b1111 : 4'b1101;
													assign node22634 = (inp[3]) ? 4'b1101 : node22635;
														assign node22635 = (inp[5]) ? 4'b1101 : 4'b1111;
									assign node22639 = (inp[4]) ? node22703 : node22640;
										assign node22640 = (inp[12]) ? node22680 : node22641;
											assign node22641 = (inp[10]) ? node22659 : node22642;
												assign node22642 = (inp[0]) ? node22654 : node22643;
													assign node22643 = (inp[15]) ? node22649 : node22644;
														assign node22644 = (inp[3]) ? node22646 : 4'b1011;
															assign node22646 = (inp[14]) ? 4'b1001 : 4'b1011;
														assign node22649 = (inp[5]) ? node22651 : 4'b1001;
															assign node22651 = (inp[3]) ? 4'b1011 : 4'b1001;
													assign node22654 = (inp[15]) ? 4'b1011 : node22655;
														assign node22655 = (inp[5]) ? 4'b1011 : 4'b1001;
												assign node22659 = (inp[0]) ? node22669 : node22660;
													assign node22660 = (inp[5]) ? 4'b1101 : node22661;
														assign node22661 = (inp[3]) ? node22665 : node22662;
															assign node22662 = (inp[15]) ? 4'b1101 : 4'b1111;
															assign node22665 = (inp[15]) ? 4'b1111 : 4'b1101;
													assign node22669 = (inp[15]) ? node22675 : node22670;
														assign node22670 = (inp[5]) ? 4'b1111 : node22671;
															assign node22671 = (inp[3]) ? 4'b1111 : 4'b1101;
														assign node22675 = (inp[5]) ? 4'b1101 : node22676;
															assign node22676 = (inp[3]) ? 4'b1101 : 4'b1111;
											assign node22680 = (inp[0]) ? node22692 : node22681;
												assign node22681 = (inp[15]) ? node22687 : node22682;
													assign node22682 = (inp[5]) ? 4'b1101 : node22683;
														assign node22683 = (inp[3]) ? 4'b1101 : 4'b1111;
													assign node22687 = (inp[3]) ? 4'b1111 : node22688;
														assign node22688 = (inp[5]) ? 4'b1111 : 4'b1101;
												assign node22692 = (inp[15]) ? node22698 : node22693;
													assign node22693 = (inp[5]) ? 4'b1111 : node22694;
														assign node22694 = (inp[3]) ? 4'b1111 : 4'b1101;
													assign node22698 = (inp[5]) ? 4'b1101 : node22699;
														assign node22699 = (inp[3]) ? 4'b1101 : 4'b1111;
										assign node22703 = (inp[12]) ? node22765 : node22704;
											assign node22704 = (inp[10]) ? node22738 : node22705;
												assign node22705 = (inp[3]) ? node22731 : node22706;
													assign node22706 = (inp[14]) ? node22722 : node22707;
														assign node22707 = (inp[15]) ? node22715 : node22708;
															assign node22708 = (inp[5]) ? node22712 : node22709;
																assign node22709 = (inp[0]) ? 4'b1101 : 4'b1111;
																assign node22712 = (inp[0]) ? 4'b1111 : 4'b1101;
															assign node22715 = (inp[0]) ? node22719 : node22716;
																assign node22716 = (inp[5]) ? 4'b1111 : 4'b1101;
																assign node22719 = (inp[5]) ? 4'b1101 : 4'b1111;
														assign node22722 = (inp[5]) ? node22724 : 4'b1101;
															assign node22724 = (inp[15]) ? node22728 : node22725;
																assign node22725 = (inp[0]) ? 4'b1111 : 4'b1101;
																assign node22728 = (inp[0]) ? 4'b1101 : 4'b1111;
													assign node22731 = (inp[0]) ? node22735 : node22732;
														assign node22732 = (inp[15]) ? 4'b1111 : 4'b1101;
														assign node22735 = (inp[15]) ? 4'b1101 : 4'b1111;
												assign node22738 = (inp[3]) ? node22750 : node22739;
													assign node22739 = (inp[0]) ? node22745 : node22740;
														assign node22740 = (inp[15]) ? 4'b1011 : node22741;
															assign node22741 = (inp[5]) ? 4'b1001 : 4'b1011;
														assign node22745 = (inp[5]) ? node22747 : 4'b1001;
															assign node22747 = (inp[15]) ? 4'b1001 : 4'b1011;
													assign node22750 = (inp[14]) ? node22758 : node22751;
														assign node22751 = (inp[15]) ? node22755 : node22752;
															assign node22752 = (inp[0]) ? 4'b1011 : 4'b1001;
															assign node22755 = (inp[0]) ? 4'b1001 : 4'b1011;
														assign node22758 = (inp[15]) ? node22762 : node22759;
															assign node22759 = (inp[0]) ? 4'b1011 : 4'b1001;
															assign node22762 = (inp[0]) ? 4'b1001 : 4'b1011;
											assign node22765 = (inp[3]) ? node22781 : node22766;
												assign node22766 = (inp[5]) ? node22774 : node22767;
													assign node22767 = (inp[0]) ? node22771 : node22768;
														assign node22768 = (inp[15]) ? 4'b1001 : 4'b1011;
														assign node22771 = (inp[15]) ? 4'b1011 : 4'b1001;
													assign node22774 = (inp[0]) ? node22778 : node22775;
														assign node22775 = (inp[15]) ? 4'b1011 : 4'b1001;
														assign node22778 = (inp[15]) ? 4'b1001 : 4'b1011;
												assign node22781 = (inp[0]) ? node22785 : node22782;
													assign node22782 = (inp[15]) ? 4'b1011 : 4'b1001;
													assign node22785 = (inp[15]) ? 4'b1001 : 4'b1011;
						assign node22788 = (inp[8]) ? node23832 : node22789;
							assign node22789 = (inp[2]) ? node23409 : node22790;
								assign node22790 = (inp[14]) ? node23084 : node22791;
									assign node22791 = (inp[3]) ? node22929 : node22792;
										assign node22792 = (inp[5]) ? node22850 : node22793;
											assign node22793 = (inp[15]) ? node22821 : node22794;
												assign node22794 = (inp[0]) ? node22812 : node22795;
													assign node22795 = (inp[12]) ? node22801 : node22796;
														assign node22796 = (inp[9]) ? 4'b0110 : node22797;
															assign node22797 = (inp[4]) ? 4'b0010 : 4'b0110;
														assign node22801 = (inp[9]) ? node22807 : node22802;
															assign node22802 = (inp[10]) ? 4'b0010 : node22803;
																assign node22803 = (inp[4]) ? 4'b0010 : 4'b0110;
															assign node22807 = (inp[10]) ? 4'b0110 : node22808;
																assign node22808 = (inp[4]) ? 4'b0110 : 4'b0010;
													assign node22812 = (inp[9]) ? node22814 : 4'b0100;
														assign node22814 = (inp[4]) ? node22818 : node22815;
															assign node22815 = (inp[12]) ? 4'b0100 : 4'b0000;
															assign node22818 = (inp[12]) ? 4'b0000 : 4'b0100;
												assign node22821 = (inp[0]) ? node22833 : node22822;
													assign node22822 = (inp[4]) ? node22828 : node22823;
														assign node22823 = (inp[9]) ? node22825 : 4'b0100;
															assign node22825 = (inp[10]) ? 4'b0100 : 4'b0000;
														assign node22828 = (inp[9]) ? node22830 : 4'b0000;
															assign node22830 = (inp[10]) ? 4'b0000 : 4'b0100;
													assign node22833 = (inp[9]) ? node22841 : node22834;
														assign node22834 = (inp[4]) ? node22838 : node22835;
															assign node22835 = (inp[10]) ? 4'b0010 : 4'b0110;
															assign node22838 = (inp[10]) ? 4'b0110 : 4'b0010;
														assign node22841 = (inp[4]) ? node22845 : node22842;
															assign node22842 = (inp[12]) ? 4'b0110 : 4'b0010;
															assign node22845 = (inp[12]) ? node22847 : 4'b0110;
																assign node22847 = (inp[10]) ? 4'b0010 : 4'b0110;
											assign node22850 = (inp[4]) ? node22888 : node22851;
												assign node22851 = (inp[9]) ? node22873 : node22852;
													assign node22852 = (inp[10]) ? node22866 : node22853;
														assign node22853 = (inp[12]) ? node22859 : node22854;
															assign node22854 = (inp[15]) ? 4'b0110 : node22855;
																assign node22855 = (inp[0]) ? 4'b0100 : 4'b0110;
															assign node22859 = (inp[0]) ? node22863 : node22860;
																assign node22860 = (inp[15]) ? 4'b0100 : 4'b0110;
																assign node22863 = (inp[15]) ? 4'b0110 : 4'b0100;
														assign node22866 = (inp[12]) ? node22868 : 4'b0110;
															assign node22868 = (inp[0]) ? node22870 : 4'b0010;
																assign node22870 = (inp[15]) ? 4'b0010 : 4'b0000;
													assign node22873 = (inp[10]) ? node22881 : node22874;
														assign node22874 = (inp[15]) ? node22878 : node22875;
															assign node22875 = (inp[0]) ? 4'b0000 : 4'b0010;
															assign node22878 = (inp[0]) ? 4'b0010 : 4'b0000;
														assign node22881 = (inp[12]) ? 4'b0110 : node22882;
															assign node22882 = (inp[15]) ? 4'b0010 : node22883;
																assign node22883 = (inp[0]) ? 4'b0000 : 4'b0010;
												assign node22888 = (inp[9]) ? node22912 : node22889;
													assign node22889 = (inp[12]) ? node22897 : node22890;
														assign node22890 = (inp[15]) ? node22894 : node22891;
															assign node22891 = (inp[0]) ? 4'b0000 : 4'b0010;
															assign node22894 = (inp[0]) ? 4'b0010 : 4'b0000;
														assign node22897 = (inp[10]) ? node22905 : node22898;
															assign node22898 = (inp[15]) ? node22902 : node22899;
																assign node22899 = (inp[0]) ? 4'b0000 : 4'b0010;
																assign node22902 = (inp[0]) ? 4'b0010 : 4'b0000;
															assign node22905 = (inp[15]) ? node22909 : node22906;
																assign node22906 = (inp[0]) ? 4'b0110 : 4'b0100;
																assign node22909 = (inp[0]) ? 4'b0100 : 4'b0110;
													assign node22912 = (inp[10]) ? node22920 : node22913;
														assign node22913 = (inp[15]) ? node22917 : node22914;
															assign node22914 = (inp[0]) ? 4'b0110 : 4'b0100;
															assign node22917 = (inp[0]) ? 4'b0100 : 4'b0110;
														assign node22920 = (inp[12]) ? node22926 : node22921;
															assign node22921 = (inp[0]) ? 4'b0100 : node22922;
																assign node22922 = (inp[15]) ? 4'b0110 : 4'b0100;
															assign node22926 = (inp[0]) ? 4'b0000 : 4'b0010;
										assign node22929 = (inp[4]) ? node23015 : node22930;
											assign node22930 = (inp[9]) ? node22976 : node22931;
												assign node22931 = (inp[10]) ? node22953 : node22932;
													assign node22932 = (inp[12]) ? node22940 : node22933;
														assign node22933 = (inp[5]) ? 4'b0100 : node22934;
															assign node22934 = (inp[15]) ? 4'b0100 : node22935;
																assign node22935 = (inp[0]) ? 4'b0100 : 4'b0110;
														assign node22940 = (inp[5]) ? node22946 : node22941;
															assign node22941 = (inp[0]) ? 4'b0110 : node22942;
																assign node22942 = (inp[15]) ? 4'b0100 : 4'b0110;
															assign node22946 = (inp[0]) ? node22950 : node22947;
																assign node22947 = (inp[15]) ? 4'b0110 : 4'b0100;
																assign node22950 = (inp[15]) ? 4'b0100 : 4'b0110;
													assign node22953 = (inp[12]) ? node22965 : node22954;
														assign node22954 = (inp[5]) ? node22960 : node22955;
															assign node22955 = (inp[15]) ? node22957 : 4'b0100;
																assign node22957 = (inp[0]) ? 4'b0110 : 4'b0100;
															assign node22960 = (inp[15]) ? 4'b0110 : node22961;
																assign node22961 = (inp[0]) ? 4'b0110 : 4'b0100;
														assign node22965 = (inp[0]) ? node22971 : node22966;
															assign node22966 = (inp[5]) ? node22968 : 4'b0000;
																assign node22968 = (inp[15]) ? 4'b0010 : 4'b0000;
															assign node22971 = (inp[5]) ? 4'b0010 : node22972;
																assign node22972 = (inp[15]) ? 4'b0010 : 4'b0000;
												assign node22976 = (inp[10]) ? node22994 : node22977;
													assign node22977 = (inp[0]) ? node22987 : node22978;
														assign node22978 = (inp[12]) ? node22980 : 4'b0010;
															assign node22980 = (inp[15]) ? node22984 : node22981;
																assign node22981 = (inp[5]) ? 4'b0000 : 4'b0010;
																assign node22984 = (inp[5]) ? 4'b0010 : 4'b0000;
														assign node22987 = (inp[5]) ? node22991 : node22988;
															assign node22988 = (inp[15]) ? 4'b0010 : 4'b0000;
															assign node22991 = (inp[15]) ? 4'b0000 : 4'b0010;
													assign node22994 = (inp[12]) ? node23008 : node22995;
														assign node22995 = (inp[15]) ? node23003 : node22996;
															assign node22996 = (inp[5]) ? node23000 : node22997;
																assign node22997 = (inp[0]) ? 4'b0000 : 4'b0010;
																assign node23000 = (inp[0]) ? 4'b0010 : 4'b0000;
															assign node23003 = (inp[5]) ? 4'b0010 : node23004;
																assign node23004 = (inp[0]) ? 4'b0010 : 4'b0000;
														assign node23008 = (inp[15]) ? node23012 : node23009;
															assign node23009 = (inp[0]) ? 4'b0110 : 4'b0100;
															assign node23012 = (inp[0]) ? 4'b0100 : 4'b0110;
											assign node23015 = (inp[9]) ? node23061 : node23016;
												assign node23016 = (inp[10]) ? node23038 : node23017;
													assign node23017 = (inp[0]) ? node23031 : node23018;
														assign node23018 = (inp[12]) ? node23024 : node23019;
															assign node23019 = (inp[5]) ? 4'b0000 : node23020;
																assign node23020 = (inp[15]) ? 4'b0000 : 4'b0010;
															assign node23024 = (inp[5]) ? node23028 : node23025;
																assign node23025 = (inp[15]) ? 4'b0000 : 4'b0010;
																assign node23028 = (inp[15]) ? 4'b0010 : 4'b0000;
														assign node23031 = (inp[5]) ? node23035 : node23032;
															assign node23032 = (inp[15]) ? 4'b0010 : 4'b0000;
															assign node23035 = (inp[15]) ? 4'b0000 : 4'b0010;
													assign node23038 = (inp[12]) ? node23054 : node23039;
														assign node23039 = (inp[5]) ? node23047 : node23040;
															assign node23040 = (inp[15]) ? node23044 : node23041;
																assign node23041 = (inp[0]) ? 4'b0000 : 4'b0010;
																assign node23044 = (inp[0]) ? 4'b0010 : 4'b0000;
															assign node23047 = (inp[0]) ? node23051 : node23048;
																assign node23048 = (inp[15]) ? 4'b0010 : 4'b0000;
																assign node23051 = (inp[15]) ? 4'b0000 : 4'b0010;
														assign node23054 = (inp[0]) ? node23058 : node23055;
															assign node23055 = (inp[15]) ? 4'b0110 : 4'b0100;
															assign node23058 = (inp[15]) ? 4'b0100 : 4'b0110;
												assign node23061 = (inp[10]) ? node23069 : node23062;
													assign node23062 = (inp[15]) ? node23066 : node23063;
														assign node23063 = (inp[0]) ? 4'b0110 : 4'b0100;
														assign node23066 = (inp[0]) ? 4'b0100 : 4'b0110;
													assign node23069 = (inp[12]) ? node23077 : node23070;
														assign node23070 = (inp[0]) ? node23074 : node23071;
															assign node23071 = (inp[15]) ? 4'b0110 : 4'b0100;
															assign node23074 = (inp[15]) ? 4'b0100 : 4'b0110;
														assign node23077 = (inp[0]) ? node23081 : node23078;
															assign node23078 = (inp[15]) ? 4'b0010 : 4'b0000;
															assign node23081 = (inp[15]) ? 4'b0000 : 4'b0010;
									assign node23084 = (inp[10]) ? node23272 : node23085;
										assign node23085 = (inp[3]) ? node23183 : node23086;
											assign node23086 = (inp[9]) ? node23128 : node23087;
												assign node23087 = (inp[15]) ? node23109 : node23088;
													assign node23088 = (inp[0]) ? node23096 : node23089;
														assign node23089 = (inp[5]) ? node23093 : node23090;
															assign node23090 = (inp[4]) ? 4'b1011 : 4'b1111;
															assign node23093 = (inp[4]) ? 4'b1101 : 4'b1011;
														assign node23096 = (inp[5]) ? node23104 : node23097;
															assign node23097 = (inp[4]) ? node23101 : node23098;
																assign node23098 = (inp[12]) ? 4'b1001 : 4'b1101;
																assign node23101 = (inp[12]) ? 4'b1101 : 4'b1001;
															assign node23104 = (inp[4]) ? 4'b1001 : node23105;
																assign node23105 = (inp[12]) ? 4'b1001 : 4'b1101;
													assign node23109 = (inp[0]) ? node23123 : node23110;
														assign node23110 = (inp[5]) ? node23118 : node23111;
															assign node23111 = (inp[12]) ? node23115 : node23112;
																assign node23112 = (inp[4]) ? 4'b1001 : 4'b1101;
																assign node23115 = (inp[4]) ? 4'b1101 : 4'b1001;
															assign node23118 = (inp[4]) ? node23120 : 4'b1001;
																assign node23120 = (inp[12]) ? 4'b1111 : 4'b1001;
														assign node23123 = (inp[4]) ? node23125 : 4'b1011;
															assign node23125 = (inp[12]) ? 4'b1101 : 4'b1011;
												assign node23128 = (inp[4]) ? node23154 : node23129;
													assign node23129 = (inp[12]) ? node23141 : node23130;
														assign node23130 = (inp[5]) ? node23136 : node23131;
															assign node23131 = (inp[15]) ? 4'b1001 : node23132;
																assign node23132 = (inp[0]) ? 4'b1001 : 4'b1011;
															assign node23136 = (inp[15]) ? node23138 : 4'b1001;
																assign node23138 = (inp[0]) ? 4'b1011 : 4'b1001;
														assign node23141 = (inp[15]) ? node23149 : node23142;
															assign node23142 = (inp[0]) ? node23146 : node23143;
																assign node23143 = (inp[5]) ? 4'b1101 : 4'b1111;
																assign node23146 = (inp[5]) ? 4'b1111 : 4'b1101;
															assign node23149 = (inp[5]) ? node23151 : 4'b1101;
																assign node23151 = (inp[0]) ? 4'b1101 : 4'b1111;
													assign node23154 = (inp[12]) ? node23170 : node23155;
														assign node23155 = (inp[0]) ? node23163 : node23156;
															assign node23156 = (inp[15]) ? node23160 : node23157;
																assign node23157 = (inp[5]) ? 4'b1101 : 4'b1111;
																assign node23160 = (inp[5]) ? 4'b1111 : 4'b1101;
															assign node23163 = (inp[5]) ? node23167 : node23164;
																assign node23164 = (inp[15]) ? 4'b1111 : 4'b1101;
																assign node23167 = (inp[15]) ? 4'b1101 : 4'b1111;
														assign node23170 = (inp[0]) ? node23176 : node23171;
															assign node23171 = (inp[5]) ? 4'b1001 : node23172;
																assign node23172 = (inp[15]) ? 4'b1001 : 4'b1011;
															assign node23176 = (inp[15]) ? node23180 : node23177;
																assign node23177 = (inp[5]) ? 4'b1011 : 4'b1001;
																assign node23180 = (inp[5]) ? 4'b1001 : 4'b1011;
											assign node23183 = (inp[4]) ? node23229 : node23184;
												assign node23184 = (inp[15]) ? node23208 : node23185;
													assign node23185 = (inp[5]) ? node23199 : node23186;
														assign node23186 = (inp[0]) ? node23194 : node23187;
															assign node23187 = (inp[9]) ? node23191 : node23188;
																assign node23188 = (inp[12]) ? 4'b1011 : 4'b1111;
																assign node23191 = (inp[12]) ? 4'b1101 : 4'b1011;
															assign node23194 = (inp[9]) ? node23196 : 4'b1001;
																assign node23196 = (inp[12]) ? 4'b1111 : 4'b1001;
														assign node23199 = (inp[0]) ? node23201 : 4'b1001;
															assign node23201 = (inp[9]) ? node23205 : node23202;
																assign node23202 = (inp[12]) ? 4'b1011 : 4'b1111;
																assign node23205 = (inp[12]) ? 4'b1111 : 4'b1011;
													assign node23208 = (inp[5]) ? node23220 : node23209;
														assign node23209 = (inp[0]) ? node23213 : node23210;
															assign node23210 = (inp[9]) ? 4'b1001 : 4'b1101;
															assign node23213 = (inp[12]) ? node23217 : node23214;
																assign node23214 = (inp[9]) ? 4'b1011 : 4'b1111;
																assign node23217 = (inp[9]) ? 4'b1101 : 4'b1011;
														assign node23220 = (inp[0]) ? node23222 : 4'b1011;
															assign node23222 = (inp[9]) ? node23226 : node23223;
																assign node23223 = (inp[12]) ? 4'b1001 : 4'b1101;
																assign node23226 = (inp[12]) ? 4'b1101 : 4'b1001;
												assign node23229 = (inp[5]) ? node23255 : node23230;
													assign node23230 = (inp[15]) ? node23246 : node23231;
														assign node23231 = (inp[0]) ? node23239 : node23232;
															assign node23232 = (inp[12]) ? node23236 : node23233;
																assign node23233 = (inp[9]) ? 4'b1101 : 4'b1011;
																assign node23236 = (inp[9]) ? 4'b1001 : 4'b1101;
															assign node23239 = (inp[9]) ? node23243 : node23240;
																assign node23240 = (inp[12]) ? 4'b1111 : 4'b1001;
																assign node23243 = (inp[12]) ? 4'b1011 : 4'b1111;
														assign node23246 = (inp[0]) ? node23252 : node23247;
															assign node23247 = (inp[9]) ? 4'b1111 : node23248;
																assign node23248 = (inp[12]) ? 4'b1111 : 4'b1001;
															assign node23252 = (inp[9]) ? 4'b1001 : 4'b1101;
													assign node23255 = (inp[15]) ? node23261 : node23256;
														assign node23256 = (inp[0]) ? 4'b1111 : node23257;
															assign node23257 = (inp[12]) ? 4'b1001 : 4'b1101;
														assign node23261 = (inp[0]) ? node23269 : node23262;
															assign node23262 = (inp[12]) ? node23266 : node23263;
																assign node23263 = (inp[9]) ? 4'b1111 : 4'b1011;
																assign node23266 = (inp[9]) ? 4'b1011 : 4'b1111;
															assign node23269 = (inp[9]) ? 4'b1101 : 4'b1001;
										assign node23272 = (inp[9]) ? node23348 : node23273;
											assign node23273 = (inp[4]) ? node23321 : node23274;
												assign node23274 = (inp[12]) ? node23296 : node23275;
													assign node23275 = (inp[15]) ? node23285 : node23276;
														assign node23276 = (inp[0]) ? node23282 : node23277;
															assign node23277 = (inp[3]) ? node23279 : 4'b1011;
																assign node23279 = (inp[5]) ? 4'b1001 : 4'b1011;
															assign node23282 = (inp[3]) ? 4'b1011 : 4'b1001;
														assign node23285 = (inp[0]) ? node23291 : node23286;
															assign node23286 = (inp[3]) ? node23288 : 4'b1001;
																assign node23288 = (inp[5]) ? 4'b1011 : 4'b1001;
															assign node23291 = (inp[5]) ? node23293 : 4'b1011;
																assign node23293 = (inp[3]) ? 4'b1001 : 4'b1011;
													assign node23296 = (inp[5]) ? node23306 : node23297;
														assign node23297 = (inp[3]) ? node23299 : 4'b1001;
															assign node23299 = (inp[15]) ? node23303 : node23300;
																assign node23300 = (inp[0]) ? 4'b1001 : 4'b1011;
																assign node23303 = (inp[0]) ? 4'b1011 : 4'b1001;
														assign node23306 = (inp[15]) ? node23314 : node23307;
															assign node23307 = (inp[3]) ? node23311 : node23308;
																assign node23308 = (inp[0]) ? 4'b1001 : 4'b1011;
																assign node23311 = (inp[0]) ? 4'b1011 : 4'b1001;
															assign node23314 = (inp[3]) ? node23318 : node23315;
																assign node23315 = (inp[0]) ? 4'b1011 : 4'b1001;
																assign node23318 = (inp[0]) ? 4'b1001 : 4'b1011;
												assign node23321 = (inp[3]) ? node23335 : node23322;
													assign node23322 = (inp[15]) ? node23328 : node23323;
														assign node23323 = (inp[5]) ? 4'b1111 : node23324;
															assign node23324 = (inp[0]) ? 4'b1101 : 4'b1111;
														assign node23328 = (inp[5]) ? node23332 : node23329;
															assign node23329 = (inp[0]) ? 4'b1111 : 4'b1101;
															assign node23332 = (inp[0]) ? 4'b1101 : 4'b1111;
													assign node23335 = (inp[5]) ? node23343 : node23336;
														assign node23336 = (inp[0]) ? node23340 : node23337;
															assign node23337 = (inp[15]) ? 4'b1111 : 4'b1101;
															assign node23340 = (inp[15]) ? 4'b1101 : 4'b1111;
														assign node23343 = (inp[0]) ? node23345 : 4'b1101;
															assign node23345 = (inp[15]) ? 4'b1101 : 4'b1111;
											assign node23348 = (inp[4]) ? node23388 : node23349;
												assign node23349 = (inp[12]) ? node23371 : node23350;
													assign node23350 = (inp[15]) ? node23360 : node23351;
														assign node23351 = (inp[0]) ? node23357 : node23352;
															assign node23352 = (inp[3]) ? 4'b1101 : node23353;
																assign node23353 = (inp[5]) ? 4'b1101 : 4'b1111;
															assign node23357 = (inp[3]) ? 4'b1111 : 4'b1101;
														assign node23360 = (inp[0]) ? node23366 : node23361;
															assign node23361 = (inp[5]) ? 4'b1111 : node23362;
																assign node23362 = (inp[3]) ? 4'b1111 : 4'b1101;
															assign node23366 = (inp[5]) ? 4'b1101 : node23367;
																assign node23367 = (inp[3]) ? 4'b1101 : 4'b1111;
													assign node23371 = (inp[0]) ? node23383 : node23372;
														assign node23372 = (inp[15]) ? node23378 : node23373;
															assign node23373 = (inp[3]) ? 4'b1101 : node23374;
																assign node23374 = (inp[5]) ? 4'b1101 : 4'b1111;
															assign node23378 = (inp[3]) ? 4'b1111 : node23379;
																assign node23379 = (inp[5]) ? 4'b1111 : 4'b1101;
														assign node23383 = (inp[3]) ? node23385 : 4'b1111;
															assign node23385 = (inp[15]) ? 4'b1101 : 4'b1111;
												assign node23388 = (inp[0]) ? node23398 : node23389;
													assign node23389 = (inp[5]) ? 4'b1011 : node23390;
														assign node23390 = (inp[15]) ? node23394 : node23391;
															assign node23391 = (inp[3]) ? 4'b1001 : 4'b1011;
															assign node23394 = (inp[3]) ? 4'b1011 : 4'b1001;
													assign node23398 = (inp[15]) ? node23404 : node23399;
														assign node23399 = (inp[5]) ? 4'b1011 : node23400;
															assign node23400 = (inp[3]) ? 4'b1011 : 4'b1001;
														assign node23404 = (inp[5]) ? 4'b1001 : node23405;
															assign node23405 = (inp[3]) ? 4'b1001 : 4'b1011;
								assign node23409 = (inp[4]) ? node23591 : node23410;
									assign node23410 = (inp[9]) ? node23484 : node23411;
										assign node23411 = (inp[12]) ? node23461 : node23412;
											assign node23412 = (inp[10]) ? node23436 : node23413;
												assign node23413 = (inp[15]) ? node23427 : node23414;
													assign node23414 = (inp[5]) ? node23416 : 4'b1111;
														assign node23416 = (inp[14]) ? node23422 : node23417;
															assign node23417 = (inp[0]) ? 4'b1111 : node23418;
																assign node23418 = (inp[3]) ? 4'b1101 : 4'b1111;
															assign node23422 = (inp[3]) ? 4'b1101 : node23423;
																assign node23423 = (inp[0]) ? 4'b1101 : 4'b1111;
													assign node23427 = (inp[5]) ? node23431 : node23428;
														assign node23428 = (inp[0]) ? 4'b1111 : 4'b1101;
														assign node23431 = (inp[0]) ? node23433 : 4'b1111;
															assign node23433 = (inp[3]) ? 4'b1101 : 4'b1111;
												assign node23436 = (inp[5]) ? node23444 : node23437;
													assign node23437 = (inp[15]) ? node23441 : node23438;
														assign node23438 = (inp[0]) ? 4'b1001 : 4'b1011;
														assign node23441 = (inp[0]) ? 4'b1011 : 4'b1001;
													assign node23444 = (inp[15]) ? node23454 : node23445;
														assign node23445 = (inp[14]) ? 4'b1011 : node23446;
															assign node23446 = (inp[3]) ? node23450 : node23447;
																assign node23447 = (inp[0]) ? 4'b1001 : 4'b1011;
																assign node23450 = (inp[0]) ? 4'b1011 : 4'b1001;
														assign node23454 = (inp[3]) ? node23458 : node23455;
															assign node23455 = (inp[0]) ? 4'b1011 : 4'b1001;
															assign node23458 = (inp[0]) ? 4'b1001 : 4'b1011;
											assign node23461 = (inp[3]) ? node23469 : node23462;
												assign node23462 = (inp[15]) ? node23466 : node23463;
													assign node23463 = (inp[0]) ? 4'b1001 : 4'b1011;
													assign node23466 = (inp[0]) ? 4'b1011 : 4'b1001;
												assign node23469 = (inp[5]) ? node23477 : node23470;
													assign node23470 = (inp[0]) ? node23474 : node23471;
														assign node23471 = (inp[15]) ? 4'b1001 : 4'b1011;
														assign node23474 = (inp[15]) ? 4'b1011 : 4'b1001;
													assign node23477 = (inp[0]) ? node23481 : node23478;
														assign node23478 = (inp[15]) ? 4'b1011 : 4'b1001;
														assign node23481 = (inp[15]) ? 4'b1001 : 4'b1011;
										assign node23484 = (inp[10]) ? node23532 : node23485;
											assign node23485 = (inp[12]) ? node23509 : node23486;
												assign node23486 = (inp[15]) ? node23498 : node23487;
													assign node23487 = (inp[0]) ? node23493 : node23488;
														assign node23488 = (inp[3]) ? node23490 : 4'b1011;
															assign node23490 = (inp[5]) ? 4'b1001 : 4'b1011;
														assign node23493 = (inp[3]) ? node23495 : 4'b1001;
															assign node23495 = (inp[5]) ? 4'b1011 : 4'b1001;
													assign node23498 = (inp[0]) ? node23504 : node23499;
														assign node23499 = (inp[3]) ? node23501 : 4'b1001;
															assign node23501 = (inp[5]) ? 4'b1011 : 4'b1001;
														assign node23504 = (inp[5]) ? node23506 : 4'b1011;
															assign node23506 = (inp[3]) ? 4'b1001 : 4'b1011;
												assign node23509 = (inp[5]) ? node23525 : node23510;
													assign node23510 = (inp[0]) ? node23518 : node23511;
														assign node23511 = (inp[3]) ? node23515 : node23512;
															assign node23512 = (inp[15]) ? 4'b1101 : 4'b1111;
															assign node23515 = (inp[15]) ? 4'b1111 : 4'b1101;
														assign node23518 = (inp[15]) ? node23522 : node23519;
															assign node23519 = (inp[3]) ? 4'b1111 : 4'b1101;
															assign node23522 = (inp[3]) ? 4'b1101 : 4'b1111;
													assign node23525 = (inp[15]) ? node23529 : node23526;
														assign node23526 = (inp[0]) ? 4'b1111 : 4'b1101;
														assign node23529 = (inp[0]) ? 4'b1101 : 4'b1111;
											assign node23532 = (inp[14]) ? node23556 : node23533;
												assign node23533 = (inp[3]) ? node23549 : node23534;
													assign node23534 = (inp[15]) ? node23542 : node23535;
														assign node23535 = (inp[5]) ? node23539 : node23536;
															assign node23536 = (inp[0]) ? 4'b1101 : 4'b1111;
															assign node23539 = (inp[0]) ? 4'b1111 : 4'b1101;
														assign node23542 = (inp[5]) ? node23546 : node23543;
															assign node23543 = (inp[12]) ? 4'b1101 : 4'b1111;
															assign node23546 = (inp[12]) ? 4'b1111 : 4'b1101;
													assign node23549 = (inp[0]) ? node23553 : node23550;
														assign node23550 = (inp[15]) ? 4'b1111 : 4'b1101;
														assign node23553 = (inp[15]) ? 4'b1101 : 4'b1111;
												assign node23556 = (inp[12]) ? node23574 : node23557;
													assign node23557 = (inp[5]) ? node23567 : node23558;
														assign node23558 = (inp[15]) ? 4'b1111 : node23559;
															assign node23559 = (inp[3]) ? node23563 : node23560;
																assign node23560 = (inp[0]) ? 4'b1101 : 4'b1111;
																assign node23563 = (inp[0]) ? 4'b1111 : 4'b1101;
														assign node23567 = (inp[15]) ? node23571 : node23568;
															assign node23568 = (inp[0]) ? 4'b1111 : 4'b1101;
															assign node23571 = (inp[0]) ? 4'b1101 : 4'b1111;
													assign node23574 = (inp[5]) ? node23584 : node23575;
														assign node23575 = (inp[15]) ? 4'b1101 : node23576;
															assign node23576 = (inp[0]) ? node23580 : node23577;
																assign node23577 = (inp[3]) ? 4'b1101 : 4'b1111;
																assign node23580 = (inp[3]) ? 4'b1111 : 4'b1101;
														assign node23584 = (inp[15]) ? node23588 : node23585;
															assign node23585 = (inp[0]) ? 4'b1111 : 4'b1101;
															assign node23588 = (inp[0]) ? 4'b1101 : 4'b1111;
									assign node23591 = (inp[9]) ? node23727 : node23592;
										assign node23592 = (inp[12]) ? node23658 : node23593;
											assign node23593 = (inp[10]) ? node23621 : node23594;
												assign node23594 = (inp[14]) ? node23612 : node23595;
													assign node23595 = (inp[3]) ? node23601 : node23596;
														assign node23596 = (inp[0]) ? node23598 : 4'b1001;
															assign node23598 = (inp[15]) ? 4'b1011 : 4'b1001;
														assign node23601 = (inp[15]) ? node23607 : node23602;
															assign node23602 = (inp[0]) ? 4'b1011 : node23603;
																assign node23603 = (inp[5]) ? 4'b1001 : 4'b1011;
															assign node23607 = (inp[5]) ? node23609 : 4'b1001;
																assign node23609 = (inp[0]) ? 4'b1001 : 4'b1011;
													assign node23612 = (inp[5]) ? node23618 : node23613;
														assign node23613 = (inp[0]) ? 4'b1011 : node23614;
															assign node23614 = (inp[3]) ? 4'b1011 : 4'b1001;
														assign node23618 = (inp[3]) ? 4'b1001 : 4'b1011;
												assign node23621 = (inp[5]) ? node23645 : node23622;
													assign node23622 = (inp[14]) ? node23630 : node23623;
														assign node23623 = (inp[15]) ? node23625 : 4'b1101;
															assign node23625 = (inp[3]) ? node23627 : 4'b1101;
																assign node23627 = (inp[0]) ? 4'b1101 : 4'b1111;
														assign node23630 = (inp[15]) ? node23638 : node23631;
															assign node23631 = (inp[3]) ? node23635 : node23632;
																assign node23632 = (inp[0]) ? 4'b1101 : 4'b1111;
																assign node23635 = (inp[0]) ? 4'b1111 : 4'b1101;
															assign node23638 = (inp[3]) ? node23642 : node23639;
																assign node23639 = (inp[0]) ? 4'b1111 : 4'b1101;
																assign node23642 = (inp[0]) ? 4'b1101 : 4'b1111;
													assign node23645 = (inp[14]) ? node23653 : node23646;
														assign node23646 = (inp[3]) ? 4'b1111 : node23647;
															assign node23647 = (inp[0]) ? 4'b1111 : node23648;
																assign node23648 = (inp[15]) ? 4'b1111 : 4'b1101;
														assign node23653 = (inp[15]) ? node23655 : 4'b1111;
															assign node23655 = (inp[0]) ? 4'b1101 : 4'b1111;
											assign node23658 = (inp[14]) ? node23704 : node23659;
												assign node23659 = (inp[10]) ? node23681 : node23660;
													assign node23660 = (inp[0]) ? node23672 : node23661;
														assign node23661 = (inp[15]) ? node23667 : node23662;
															assign node23662 = (inp[3]) ? 4'b1101 : node23663;
																assign node23663 = (inp[5]) ? 4'b1101 : 4'b1111;
															assign node23667 = (inp[3]) ? 4'b1111 : node23668;
																assign node23668 = (inp[5]) ? 4'b1111 : 4'b1101;
														assign node23672 = (inp[15]) ? node23676 : node23673;
															assign node23673 = (inp[5]) ? 4'b1111 : 4'b1101;
															assign node23676 = (inp[5]) ? 4'b1101 : node23677;
																assign node23677 = (inp[3]) ? 4'b1101 : 4'b1111;
													assign node23681 = (inp[3]) ? node23697 : node23682;
														assign node23682 = (inp[15]) ? node23690 : node23683;
															assign node23683 = (inp[5]) ? node23687 : node23684;
																assign node23684 = (inp[0]) ? 4'b1101 : 4'b1111;
																assign node23687 = (inp[0]) ? 4'b1111 : 4'b1101;
															assign node23690 = (inp[5]) ? node23694 : node23691;
																assign node23691 = (inp[0]) ? 4'b1111 : 4'b1101;
																assign node23694 = (inp[0]) ? 4'b1101 : 4'b1111;
														assign node23697 = (inp[0]) ? node23701 : node23698;
															assign node23698 = (inp[15]) ? 4'b1111 : 4'b1101;
															assign node23701 = (inp[15]) ? 4'b1101 : 4'b1111;
												assign node23704 = (inp[3]) ? node23720 : node23705;
													assign node23705 = (inp[15]) ? node23711 : node23706;
														assign node23706 = (inp[5]) ? 4'b1101 : node23707;
															assign node23707 = (inp[0]) ? 4'b1101 : 4'b1111;
														assign node23711 = (inp[10]) ? 4'b1111 : node23712;
															assign node23712 = (inp[5]) ? node23716 : node23713;
																assign node23713 = (inp[0]) ? 4'b1111 : 4'b1101;
																assign node23716 = (inp[0]) ? 4'b1101 : 4'b1111;
													assign node23720 = (inp[15]) ? node23724 : node23721;
														assign node23721 = (inp[0]) ? 4'b1111 : 4'b1101;
														assign node23724 = (inp[0]) ? 4'b1101 : 4'b1111;
										assign node23727 = (inp[10]) ? node23797 : node23728;
											assign node23728 = (inp[12]) ? node23768 : node23729;
												assign node23729 = (inp[5]) ? node23761 : node23730;
													assign node23730 = (inp[14]) ? node23746 : node23731;
														assign node23731 = (inp[0]) ? node23739 : node23732;
															assign node23732 = (inp[3]) ? node23736 : node23733;
																assign node23733 = (inp[15]) ? 4'b1101 : 4'b1111;
																assign node23736 = (inp[15]) ? 4'b1111 : 4'b1101;
															assign node23739 = (inp[15]) ? node23743 : node23740;
																assign node23740 = (inp[3]) ? 4'b1111 : 4'b1101;
																assign node23743 = (inp[3]) ? 4'b1101 : 4'b1111;
														assign node23746 = (inp[0]) ? node23754 : node23747;
															assign node23747 = (inp[3]) ? node23751 : node23748;
																assign node23748 = (inp[15]) ? 4'b1101 : 4'b1111;
																assign node23751 = (inp[15]) ? 4'b1111 : 4'b1101;
															assign node23754 = (inp[3]) ? node23758 : node23755;
																assign node23755 = (inp[15]) ? 4'b1111 : 4'b1101;
																assign node23758 = (inp[15]) ? 4'b1101 : 4'b1111;
													assign node23761 = (inp[15]) ? node23765 : node23762;
														assign node23762 = (inp[0]) ? 4'b1111 : 4'b1101;
														assign node23765 = (inp[0]) ? 4'b1101 : 4'b1111;
												assign node23768 = (inp[3]) ? node23784 : node23769;
													assign node23769 = (inp[5]) ? node23777 : node23770;
														assign node23770 = (inp[15]) ? node23774 : node23771;
															assign node23771 = (inp[0]) ? 4'b1001 : 4'b1011;
															assign node23774 = (inp[0]) ? 4'b1011 : 4'b1001;
														assign node23777 = (inp[15]) ? node23781 : node23778;
															assign node23778 = (inp[0]) ? 4'b1011 : 4'b1001;
															assign node23781 = (inp[0]) ? 4'b1001 : 4'b1011;
													assign node23784 = (inp[14]) ? node23790 : node23785;
														assign node23785 = (inp[15]) ? node23787 : 4'b1011;
															assign node23787 = (inp[0]) ? 4'b1001 : 4'b1011;
														assign node23790 = (inp[0]) ? node23794 : node23791;
															assign node23791 = (inp[15]) ? 4'b1011 : 4'b1001;
															assign node23794 = (inp[15]) ? 4'b1001 : 4'b1011;
											assign node23797 = (inp[5]) ? node23825 : node23798;
												assign node23798 = (inp[15]) ? node23820 : node23799;
													assign node23799 = (inp[12]) ? node23813 : node23800;
														assign node23800 = (inp[14]) ? node23806 : node23801;
															assign node23801 = (inp[0]) ? node23803 : 4'b1001;
																assign node23803 = (inp[3]) ? 4'b1011 : 4'b1001;
															assign node23806 = (inp[0]) ? node23810 : node23807;
																assign node23807 = (inp[3]) ? 4'b1001 : 4'b1011;
																assign node23810 = (inp[3]) ? 4'b1011 : 4'b1001;
														assign node23813 = (inp[0]) ? node23817 : node23814;
															assign node23814 = (inp[3]) ? 4'b1001 : 4'b1011;
															assign node23817 = (inp[3]) ? 4'b1011 : 4'b1001;
													assign node23820 = (inp[3]) ? node23822 : 4'b1001;
														assign node23822 = (inp[0]) ? 4'b1001 : 4'b1011;
												assign node23825 = (inp[15]) ? node23829 : node23826;
													assign node23826 = (inp[0]) ? 4'b1011 : 4'b1001;
													assign node23829 = (inp[0]) ? 4'b1001 : 4'b1011;
							assign node23832 = (inp[14]) ? node24382 : node23833;
								assign node23833 = (inp[2]) ? node24085 : node23834;
									assign node23834 = (inp[4]) ? node23952 : node23835;
										assign node23835 = (inp[9]) ? node23899 : node23836;
											assign node23836 = (inp[10]) ? node23880 : node23837;
												assign node23837 = (inp[12]) ? node23859 : node23838;
													assign node23838 = (inp[3]) ? node23846 : node23839;
														assign node23839 = (inp[0]) ? node23843 : node23840;
															assign node23840 = (inp[15]) ? 4'b1101 : 4'b1111;
															assign node23843 = (inp[15]) ? 4'b1111 : 4'b1101;
														assign node23846 = (inp[0]) ? node23854 : node23847;
															assign node23847 = (inp[15]) ? node23851 : node23848;
																assign node23848 = (inp[5]) ? 4'b1101 : 4'b1111;
																assign node23851 = (inp[5]) ? 4'b1111 : 4'b1101;
															assign node23854 = (inp[15]) ? node23856 : 4'b1101;
																assign node23856 = (inp[5]) ? 4'b1101 : 4'b1111;
													assign node23859 = (inp[3]) ? node23871 : node23860;
														assign node23860 = (inp[5]) ? node23866 : node23861;
															assign node23861 = (inp[15]) ? 4'b1011 : node23862;
																assign node23862 = (inp[0]) ? 4'b1001 : 4'b1011;
															assign node23866 = (inp[15]) ? node23868 : 4'b1011;
																assign node23868 = (inp[0]) ? 4'b1011 : 4'b1001;
														assign node23871 = (inp[0]) ? node23873 : 4'b1001;
															assign node23873 = (inp[5]) ? node23877 : node23874;
																assign node23874 = (inp[15]) ? 4'b1011 : 4'b1001;
																assign node23877 = (inp[15]) ? 4'b1001 : 4'b1011;
												assign node23880 = (inp[15]) ? node23892 : node23881;
													assign node23881 = (inp[0]) ? node23887 : node23882;
														assign node23882 = (inp[3]) ? node23884 : 4'b1011;
															assign node23884 = (inp[5]) ? 4'b1001 : 4'b1011;
														assign node23887 = (inp[5]) ? node23889 : 4'b1001;
															assign node23889 = (inp[3]) ? 4'b1011 : 4'b1001;
													assign node23892 = (inp[0]) ? 4'b1011 : node23893;
														assign node23893 = (inp[3]) ? node23895 : 4'b1001;
															assign node23895 = (inp[5]) ? 4'b1011 : 4'b1001;
											assign node23899 = (inp[10]) ? node23935 : node23900;
												assign node23900 = (inp[12]) ? node23920 : node23901;
													assign node23901 = (inp[0]) ? node23913 : node23902;
														assign node23902 = (inp[15]) ? node23908 : node23903;
															assign node23903 = (inp[3]) ? node23905 : 4'b1011;
																assign node23905 = (inp[5]) ? 4'b1001 : 4'b1011;
															assign node23908 = (inp[3]) ? node23910 : 4'b1001;
																assign node23910 = (inp[5]) ? 4'b1011 : 4'b1001;
														assign node23913 = (inp[3]) ? node23915 : 4'b1011;
															assign node23915 = (inp[15]) ? node23917 : 4'b1011;
																assign node23917 = (inp[5]) ? 4'b1001 : 4'b1011;
													assign node23920 = (inp[0]) ? node23926 : node23921;
														assign node23921 = (inp[15]) ? 4'b1111 : node23922;
															assign node23922 = (inp[3]) ? 4'b1101 : 4'b1111;
														assign node23926 = (inp[3]) ? node23932 : node23927;
															assign node23927 = (inp[15]) ? node23929 : 4'b1101;
																assign node23929 = (inp[5]) ? 4'b1101 : 4'b1111;
															assign node23932 = (inp[15]) ? 4'b1101 : 4'b1111;
												assign node23935 = (inp[5]) ? node23945 : node23936;
													assign node23936 = (inp[3]) ? node23938 : 4'b1101;
														assign node23938 = (inp[15]) ? node23942 : node23939;
															assign node23939 = (inp[0]) ? 4'b1111 : 4'b1101;
															assign node23942 = (inp[0]) ? 4'b1101 : 4'b1111;
													assign node23945 = (inp[15]) ? node23949 : node23946;
														assign node23946 = (inp[0]) ? 4'b1111 : 4'b1101;
														assign node23949 = (inp[0]) ? 4'b1101 : 4'b1111;
										assign node23952 = (inp[9]) ? node24028 : node23953;
											assign node23953 = (inp[10]) ? node23993 : node23954;
												assign node23954 = (inp[12]) ? node23972 : node23955;
													assign node23955 = (inp[3]) ? node23963 : node23956;
														assign node23956 = (inp[0]) ? node23960 : node23957;
															assign node23957 = (inp[15]) ? 4'b1001 : 4'b1011;
															assign node23960 = (inp[15]) ? 4'b1011 : 4'b1001;
														assign node23963 = (inp[0]) ? 4'b1011 : node23964;
															assign node23964 = (inp[5]) ? node23968 : node23965;
																assign node23965 = (inp[15]) ? 4'b1001 : 4'b1011;
																assign node23968 = (inp[15]) ? 4'b1011 : 4'b1001;
													assign node23972 = (inp[0]) ? node23982 : node23973;
														assign node23973 = (inp[15]) ? node23979 : node23974;
															assign node23974 = (inp[5]) ? 4'b1101 : node23975;
																assign node23975 = (inp[3]) ? 4'b1101 : 4'b1111;
															assign node23979 = (inp[3]) ? 4'b1111 : 4'b1101;
														assign node23982 = (inp[15]) ? node23988 : node23983;
															assign node23983 = (inp[5]) ? 4'b1111 : node23984;
																assign node23984 = (inp[3]) ? 4'b1111 : 4'b1101;
															assign node23988 = (inp[5]) ? 4'b1101 : node23989;
																assign node23989 = (inp[3]) ? 4'b1101 : 4'b1111;
												assign node23993 = (inp[5]) ? node24009 : node23994;
													assign node23994 = (inp[15]) ? node24002 : node23995;
														assign node23995 = (inp[0]) ? node23999 : node23996;
															assign node23996 = (inp[3]) ? 4'b1101 : 4'b1111;
															assign node23999 = (inp[3]) ? 4'b1111 : 4'b1101;
														assign node24002 = (inp[0]) ? node24006 : node24003;
															assign node24003 = (inp[3]) ? 4'b1111 : 4'b1101;
															assign node24006 = (inp[3]) ? 4'b1101 : 4'b1111;
													assign node24009 = (inp[12]) ? node24021 : node24010;
														assign node24010 = (inp[3]) ? node24016 : node24011;
															assign node24011 = (inp[0]) ? node24013 : 4'b1101;
																assign node24013 = (inp[15]) ? 4'b1101 : 4'b1111;
															assign node24016 = (inp[0]) ? 4'b1101 : node24017;
																assign node24017 = (inp[15]) ? 4'b1111 : 4'b1101;
														assign node24021 = (inp[15]) ? node24025 : node24022;
															assign node24022 = (inp[0]) ? 4'b1111 : 4'b1101;
															assign node24025 = (inp[0]) ? 4'b1101 : 4'b1111;
											assign node24028 = (inp[10]) ? node24060 : node24029;
												assign node24029 = (inp[12]) ? node24045 : node24030;
													assign node24030 = (inp[3]) ? node24038 : node24031;
														assign node24031 = (inp[5]) ? 4'b1101 : node24032;
															assign node24032 = (inp[0]) ? node24034 : 4'b1101;
																assign node24034 = (inp[15]) ? 4'b1111 : 4'b1101;
														assign node24038 = (inp[0]) ? node24042 : node24039;
															assign node24039 = (inp[15]) ? 4'b1111 : 4'b1101;
															assign node24042 = (inp[15]) ? 4'b1101 : 4'b1111;
													assign node24045 = (inp[3]) ? node24055 : node24046;
														assign node24046 = (inp[0]) ? 4'b1011 : node24047;
															assign node24047 = (inp[5]) ? node24051 : node24048;
																assign node24048 = (inp[15]) ? 4'b1001 : 4'b1011;
																assign node24051 = (inp[15]) ? 4'b1011 : 4'b1001;
														assign node24055 = (inp[15]) ? node24057 : 4'b1001;
															assign node24057 = (inp[0]) ? 4'b1001 : 4'b1011;
												assign node24060 = (inp[5]) ? node24078 : node24061;
													assign node24061 = (inp[0]) ? node24071 : node24062;
														assign node24062 = (inp[12]) ? node24064 : 4'b1011;
															assign node24064 = (inp[15]) ? node24068 : node24065;
																assign node24065 = (inp[3]) ? 4'b1001 : 4'b1011;
																assign node24068 = (inp[3]) ? 4'b1011 : 4'b1001;
														assign node24071 = (inp[15]) ? node24075 : node24072;
															assign node24072 = (inp[3]) ? 4'b1011 : 4'b1001;
															assign node24075 = (inp[3]) ? 4'b1001 : 4'b1011;
													assign node24078 = (inp[0]) ? node24082 : node24079;
														assign node24079 = (inp[15]) ? 4'b1011 : 4'b1001;
														assign node24082 = (inp[15]) ? 4'b1001 : 4'b1011;
									assign node24085 = (inp[3]) ? node24231 : node24086;
										assign node24086 = (inp[5]) ? node24156 : node24087;
											assign node24087 = (inp[9]) ? node24121 : node24088;
												assign node24088 = (inp[4]) ? node24102 : node24089;
													assign node24089 = (inp[12]) ? node24097 : node24090;
														assign node24090 = (inp[10]) ? 4'b1010 : node24091;
															assign node24091 = (inp[0]) ? node24093 : 4'b1100;
																assign node24093 = (inp[15]) ? 4'b1110 : 4'b1100;
														assign node24097 = (inp[15]) ? node24099 : 4'b1010;
															assign node24099 = (inp[0]) ? 4'b1010 : 4'b1000;
													assign node24102 = (inp[12]) ? node24110 : node24103;
														assign node24103 = (inp[10]) ? 4'b1110 : node24104;
															assign node24104 = (inp[15]) ? 4'b1000 : node24105;
																assign node24105 = (inp[0]) ? 4'b1000 : 4'b1010;
														assign node24110 = (inp[10]) ? node24116 : node24111;
															assign node24111 = (inp[0]) ? node24113 : 4'b1110;
																assign node24113 = (inp[15]) ? 4'b1110 : 4'b1100;
															assign node24116 = (inp[0]) ? node24118 : 4'b1100;
																assign node24118 = (inp[15]) ? 4'b1110 : 4'b1100;
												assign node24121 = (inp[4]) ? node24141 : node24122;
													assign node24122 = (inp[12]) ? node24134 : node24123;
														assign node24123 = (inp[10]) ? node24129 : node24124;
															assign node24124 = (inp[0]) ? node24126 : 4'b1010;
																assign node24126 = (inp[15]) ? 4'b1010 : 4'b1000;
															assign node24129 = (inp[0]) ? 4'b1100 : node24130;
																assign node24130 = (inp[15]) ? 4'b1100 : 4'b1110;
														assign node24134 = (inp[0]) ? node24138 : node24135;
															assign node24135 = (inp[15]) ? 4'b1100 : 4'b1110;
															assign node24138 = (inp[15]) ? 4'b1110 : 4'b1100;
													assign node24141 = (inp[10]) ? node24149 : node24142;
														assign node24142 = (inp[12]) ? 4'b1010 : node24143;
															assign node24143 = (inp[0]) ? 4'b1100 : node24144;
																assign node24144 = (inp[15]) ? 4'b1100 : 4'b1110;
														assign node24149 = (inp[12]) ? 4'b1000 : node24150;
															assign node24150 = (inp[15]) ? 4'b1010 : node24151;
																assign node24151 = (inp[0]) ? 4'b1000 : 4'b1010;
											assign node24156 = (inp[12]) ? node24204 : node24157;
												assign node24157 = (inp[15]) ? node24179 : node24158;
													assign node24158 = (inp[4]) ? node24170 : node24159;
														assign node24159 = (inp[10]) ? node24163 : node24160;
															assign node24160 = (inp[9]) ? 4'b1010 : 4'b1110;
															assign node24163 = (inp[9]) ? node24167 : node24164;
																assign node24164 = (inp[0]) ? 4'b1000 : 4'b1010;
																assign node24167 = (inp[0]) ? 4'b1110 : 4'b1100;
														assign node24170 = (inp[0]) ? node24174 : node24171;
															assign node24171 = (inp[10]) ? 4'b1000 : 4'b1100;
															assign node24174 = (inp[10]) ? node24176 : 4'b1000;
																assign node24176 = (inp[9]) ? 4'b1010 : 4'b1110;
													assign node24179 = (inp[10]) ? node24195 : node24180;
														assign node24180 = (inp[0]) ? node24188 : node24181;
															assign node24181 = (inp[9]) ? node24185 : node24182;
																assign node24182 = (inp[4]) ? 4'b1000 : 4'b1100;
																assign node24185 = (inp[4]) ? 4'b1110 : 4'b1000;
															assign node24188 = (inp[4]) ? node24192 : node24189;
																assign node24189 = (inp[9]) ? 4'b1010 : 4'b1110;
																assign node24192 = (inp[9]) ? 4'b1100 : 4'b1010;
														assign node24195 = (inp[0]) ? 4'b1100 : node24196;
															assign node24196 = (inp[4]) ? node24200 : node24197;
																assign node24197 = (inp[9]) ? 4'b1110 : 4'b1000;
																assign node24200 = (inp[9]) ? 4'b1010 : 4'b1110;
												assign node24204 = (inp[0]) ? node24214 : node24205;
													assign node24205 = (inp[15]) ? node24211 : node24206;
														assign node24206 = (inp[9]) ? node24208 : 4'b1100;
															assign node24208 = (inp[4]) ? 4'b1000 : 4'b1100;
														assign node24211 = (inp[9]) ? 4'b1110 : 4'b1000;
													assign node24214 = (inp[15]) ? node24222 : node24215;
														assign node24215 = (inp[4]) ? node24219 : node24216;
															assign node24216 = (inp[9]) ? 4'b1110 : 4'b1000;
															assign node24219 = (inp[9]) ? 4'b1010 : 4'b1110;
														assign node24222 = (inp[10]) ? node24224 : 4'b1100;
															assign node24224 = (inp[4]) ? node24228 : node24225;
																assign node24225 = (inp[9]) ? 4'b1100 : 4'b1010;
																assign node24228 = (inp[9]) ? 4'b1000 : 4'b1100;
										assign node24231 = (inp[10]) ? node24311 : node24232;
											assign node24232 = (inp[15]) ? node24270 : node24233;
												assign node24233 = (inp[0]) ? node24251 : node24234;
													assign node24234 = (inp[9]) ? node24244 : node24235;
														assign node24235 = (inp[4]) ? node24241 : node24236;
															assign node24236 = (inp[5]) ? 4'b1100 : node24237;
																assign node24237 = (inp[12]) ? 4'b1010 : 4'b1110;
															assign node24241 = (inp[12]) ? 4'b1100 : 4'b1000;
														assign node24244 = (inp[4]) ? node24248 : node24245;
															assign node24245 = (inp[12]) ? 4'b1100 : 4'b1000;
															assign node24248 = (inp[12]) ? 4'b1000 : 4'b1100;
													assign node24251 = (inp[9]) ? node24261 : node24252;
														assign node24252 = (inp[5]) ? 4'b1010 : node24253;
															assign node24253 = (inp[12]) ? node24257 : node24254;
																assign node24254 = (inp[4]) ? 4'b1000 : 4'b1100;
																assign node24257 = (inp[4]) ? 4'b1110 : 4'b1000;
														assign node24261 = (inp[5]) ? node24265 : node24262;
															assign node24262 = (inp[4]) ? 4'b1010 : 4'b1110;
															assign node24265 = (inp[12]) ? 4'b1010 : node24266;
																assign node24266 = (inp[4]) ? 4'b1110 : 4'b1010;
												assign node24270 = (inp[0]) ? node24290 : node24271;
													assign node24271 = (inp[5]) ? node24281 : node24272;
														assign node24272 = (inp[4]) ? node24274 : 4'b1000;
															assign node24274 = (inp[9]) ? node24278 : node24275;
																assign node24275 = (inp[12]) ? 4'b1110 : 4'b1000;
																assign node24278 = (inp[12]) ? 4'b1010 : 4'b1110;
														assign node24281 = (inp[12]) ? 4'b1010 : node24282;
															assign node24282 = (inp[9]) ? node24286 : node24283;
																assign node24283 = (inp[4]) ? 4'b1010 : 4'b1110;
																assign node24286 = (inp[4]) ? 4'b1110 : 4'b1010;
													assign node24290 = (inp[5]) ? node24304 : node24291;
														assign node24291 = (inp[4]) ? node24297 : node24292;
															assign node24292 = (inp[9]) ? node24294 : 4'b1010;
																assign node24294 = (inp[12]) ? 4'b1100 : 4'b1010;
															assign node24297 = (inp[12]) ? node24301 : node24298;
																assign node24298 = (inp[9]) ? 4'b1100 : 4'b1010;
																assign node24301 = (inp[9]) ? 4'b1000 : 4'b1100;
														assign node24304 = (inp[4]) ? 4'b1000 : node24305;
															assign node24305 = (inp[12]) ? 4'b1000 : node24306;
																assign node24306 = (inp[9]) ? 4'b1000 : 4'b1100;
											assign node24311 = (inp[9]) ? node24353 : node24312;
												assign node24312 = (inp[4]) ? node24334 : node24313;
													assign node24313 = (inp[12]) ? node24321 : node24314;
														assign node24314 = (inp[0]) ? node24316 : 4'b1000;
															assign node24316 = (inp[15]) ? 4'b1000 : node24317;
																assign node24317 = (inp[5]) ? 4'b1010 : 4'b1000;
														assign node24321 = (inp[15]) ? node24329 : node24322;
															assign node24322 = (inp[0]) ? node24326 : node24323;
																assign node24323 = (inp[5]) ? 4'b1000 : 4'b1010;
																assign node24326 = (inp[5]) ? 4'b1010 : 4'b1000;
															assign node24329 = (inp[0]) ? 4'b1000 : node24330;
																assign node24330 = (inp[5]) ? 4'b1010 : 4'b1000;
													assign node24334 = (inp[5]) ? node24340 : node24335;
														assign node24335 = (inp[0]) ? node24337 : 4'b1100;
															assign node24337 = (inp[15]) ? 4'b1100 : 4'b1110;
														assign node24340 = (inp[12]) ? node24346 : node24341;
															assign node24341 = (inp[15]) ? node24343 : 4'b1110;
																assign node24343 = (inp[0]) ? 4'b1100 : 4'b1110;
															assign node24346 = (inp[15]) ? node24350 : node24347;
																assign node24347 = (inp[0]) ? 4'b1110 : 4'b1100;
																assign node24350 = (inp[0]) ? 4'b1100 : 4'b1110;
												assign node24353 = (inp[4]) ? node24375 : node24354;
													assign node24354 = (inp[5]) ? node24362 : node24355;
														assign node24355 = (inp[0]) ? node24359 : node24356;
															assign node24356 = (inp[15]) ? 4'b1110 : 4'b1100;
															assign node24359 = (inp[15]) ? 4'b1100 : 4'b1110;
														assign node24362 = (inp[12]) ? node24370 : node24363;
															assign node24363 = (inp[15]) ? node24367 : node24364;
																assign node24364 = (inp[0]) ? 4'b1110 : 4'b1100;
																assign node24367 = (inp[0]) ? 4'b1100 : 4'b1110;
															assign node24370 = (inp[0]) ? node24372 : 4'b1110;
																assign node24372 = (inp[15]) ? 4'b1100 : 4'b1110;
													assign node24375 = (inp[0]) ? node24379 : node24376;
														assign node24376 = (inp[15]) ? 4'b1010 : 4'b1000;
														assign node24379 = (inp[15]) ? 4'b1000 : 4'b1010;
								assign node24382 = (inp[12]) ? node24644 : node24383;
									assign node24383 = (inp[15]) ? node24521 : node24384;
										assign node24384 = (inp[4]) ? node24450 : node24385;
											assign node24385 = (inp[0]) ? node24421 : node24386;
												assign node24386 = (inp[3]) ? node24400 : node24387;
													assign node24387 = (inp[2]) ? node24393 : node24388;
														assign node24388 = (inp[9]) ? 4'b1010 : node24389;
															assign node24389 = (inp[10]) ? 4'b1010 : 4'b1110;
														assign node24393 = (inp[10]) ? node24397 : node24394;
															assign node24394 = (inp[5]) ? 4'b1110 : 4'b1010;
															assign node24397 = (inp[9]) ? 4'b1110 : 4'b1010;
													assign node24400 = (inp[5]) ? node24408 : node24401;
														assign node24401 = (inp[9]) ? node24405 : node24402;
															assign node24402 = (inp[10]) ? 4'b1010 : 4'b1110;
															assign node24405 = (inp[10]) ? 4'b1100 : 4'b1010;
														assign node24408 = (inp[2]) ? node24416 : node24409;
															assign node24409 = (inp[9]) ? node24413 : node24410;
																assign node24410 = (inp[10]) ? 4'b1000 : 4'b1100;
																assign node24413 = (inp[10]) ? 4'b1100 : 4'b1000;
															assign node24416 = (inp[10]) ? node24418 : 4'b1000;
																assign node24418 = (inp[9]) ? 4'b1100 : 4'b1000;
												assign node24421 = (inp[3]) ? node24431 : node24422;
													assign node24422 = (inp[10]) ? node24426 : node24423;
														assign node24423 = (inp[9]) ? 4'b1000 : 4'b1100;
														assign node24426 = (inp[9]) ? node24428 : 4'b1000;
															assign node24428 = (inp[5]) ? 4'b1110 : 4'b1100;
													assign node24431 = (inp[5]) ? node24439 : node24432;
														assign node24432 = (inp[2]) ? 4'b1000 : node24433;
															assign node24433 = (inp[10]) ? 4'b1110 : node24434;
																assign node24434 = (inp[9]) ? 4'b1000 : 4'b1100;
														assign node24439 = (inp[2]) ? node24445 : node24440;
															assign node24440 = (inp[10]) ? 4'b1110 : node24441;
																assign node24441 = (inp[9]) ? 4'b1010 : 4'b1110;
															assign node24445 = (inp[10]) ? 4'b1010 : node24446;
																assign node24446 = (inp[9]) ? 4'b1010 : 4'b1110;
											assign node24450 = (inp[0]) ? node24490 : node24451;
												assign node24451 = (inp[5]) ? node24467 : node24452;
													assign node24452 = (inp[3]) ? node24460 : node24453;
														assign node24453 = (inp[9]) ? node24457 : node24454;
															assign node24454 = (inp[10]) ? 4'b1110 : 4'b1010;
															assign node24457 = (inp[10]) ? 4'b1010 : 4'b1110;
														assign node24460 = (inp[9]) ? node24464 : node24461;
															assign node24461 = (inp[10]) ? 4'b1100 : 4'b1010;
															assign node24464 = (inp[10]) ? 4'b1000 : 4'b1100;
													assign node24467 = (inp[3]) ? node24475 : node24468;
														assign node24468 = (inp[9]) ? node24472 : node24469;
															assign node24469 = (inp[10]) ? 4'b1100 : 4'b1010;
															assign node24472 = (inp[10]) ? 4'b1000 : 4'b1100;
														assign node24475 = (inp[2]) ? node24483 : node24476;
															assign node24476 = (inp[10]) ? node24480 : node24477;
																assign node24477 = (inp[9]) ? 4'b1100 : 4'b1000;
																assign node24480 = (inp[9]) ? 4'b1000 : 4'b1100;
															assign node24483 = (inp[10]) ? node24487 : node24484;
																assign node24484 = (inp[9]) ? 4'b1100 : 4'b1000;
																assign node24487 = (inp[9]) ? 4'b1000 : 4'b1100;
												assign node24490 = (inp[3]) ? node24512 : node24491;
													assign node24491 = (inp[5]) ? node24501 : node24492;
														assign node24492 = (inp[2]) ? node24494 : 4'b1100;
															assign node24494 = (inp[9]) ? node24498 : node24495;
																assign node24495 = (inp[10]) ? 4'b1100 : 4'b1000;
																assign node24498 = (inp[10]) ? 4'b1000 : 4'b1100;
														assign node24501 = (inp[2]) ? node24507 : node24502;
															assign node24502 = (inp[10]) ? 4'b1110 : node24503;
																assign node24503 = (inp[9]) ? 4'b1110 : 4'b1000;
															assign node24507 = (inp[10]) ? node24509 : 4'b1110;
																assign node24509 = (inp[9]) ? 4'b1010 : 4'b1110;
													assign node24512 = (inp[9]) ? node24518 : node24513;
														assign node24513 = (inp[10]) ? 4'b1110 : node24514;
															assign node24514 = (inp[5]) ? 4'b1010 : 4'b1000;
														assign node24518 = (inp[10]) ? 4'b1010 : 4'b1110;
										assign node24521 = (inp[3]) ? node24575 : node24522;
											assign node24522 = (inp[0]) ? node24552 : node24523;
												assign node24523 = (inp[9]) ? node24531 : node24524;
													assign node24524 = (inp[4]) ? node24528 : node24525;
														assign node24525 = (inp[10]) ? 4'b1000 : 4'b1100;
														assign node24528 = (inp[10]) ? 4'b1100 : 4'b1000;
													assign node24531 = (inp[5]) ? node24545 : node24532;
														assign node24532 = (inp[2]) ? node24538 : node24533;
															assign node24533 = (inp[10]) ? node24535 : 4'b1100;
																assign node24535 = (inp[4]) ? 4'b1000 : 4'b1100;
															assign node24538 = (inp[4]) ? node24542 : node24539;
																assign node24539 = (inp[10]) ? 4'b1100 : 4'b1000;
																assign node24542 = (inp[10]) ? 4'b1000 : 4'b1100;
														assign node24545 = (inp[4]) ? node24549 : node24546;
															assign node24546 = (inp[10]) ? 4'b1110 : 4'b1000;
															assign node24549 = (inp[10]) ? 4'b1010 : 4'b1110;
												assign node24552 = (inp[5]) ? node24562 : node24553;
													assign node24553 = (inp[4]) ? 4'b1010 : node24554;
														assign node24554 = (inp[9]) ? node24558 : node24555;
															assign node24555 = (inp[10]) ? 4'b1010 : 4'b1110;
															assign node24558 = (inp[10]) ? 4'b1110 : 4'b1010;
													assign node24562 = (inp[10]) ? node24568 : node24563;
														assign node24563 = (inp[4]) ? 4'b1010 : node24564;
															assign node24564 = (inp[9]) ? 4'b1010 : 4'b1110;
														assign node24568 = (inp[4]) ? node24572 : node24569;
															assign node24569 = (inp[9]) ? 4'b1100 : 4'b1010;
															assign node24572 = (inp[9]) ? 4'b1000 : 4'b1100;
											assign node24575 = (inp[0]) ? node24605 : node24576;
												assign node24576 = (inp[5]) ? node24590 : node24577;
													assign node24577 = (inp[4]) ? node24583 : node24578;
														assign node24578 = (inp[9]) ? 4'b1000 : node24579;
															assign node24579 = (inp[10]) ? 4'b1000 : 4'b1100;
														assign node24583 = (inp[9]) ? node24587 : node24584;
															assign node24584 = (inp[10]) ? 4'b1110 : 4'b1000;
															assign node24587 = (inp[10]) ? 4'b1010 : 4'b1110;
													assign node24590 = (inp[4]) ? node24598 : node24591;
														assign node24591 = (inp[9]) ? node24595 : node24592;
															assign node24592 = (inp[10]) ? 4'b1010 : 4'b1110;
															assign node24595 = (inp[10]) ? 4'b1110 : 4'b1010;
														assign node24598 = (inp[10]) ? node24602 : node24599;
															assign node24599 = (inp[9]) ? 4'b1110 : 4'b1010;
															assign node24602 = (inp[9]) ? 4'b1010 : 4'b1110;
												assign node24605 = (inp[5]) ? node24623 : node24606;
													assign node24606 = (inp[10]) ? node24616 : node24607;
														assign node24607 = (inp[2]) ? node24609 : 4'b1010;
															assign node24609 = (inp[4]) ? node24613 : node24610;
																assign node24610 = (inp[9]) ? 4'b1010 : 4'b1110;
																assign node24613 = (inp[9]) ? 4'b1100 : 4'b1010;
														assign node24616 = (inp[4]) ? node24620 : node24617;
															assign node24617 = (inp[9]) ? 4'b1100 : 4'b1010;
															assign node24620 = (inp[9]) ? 4'b1000 : 4'b1100;
													assign node24623 = (inp[2]) ? node24639 : node24624;
														assign node24624 = (inp[10]) ? node24632 : node24625;
															assign node24625 = (inp[4]) ? node24629 : node24626;
																assign node24626 = (inp[9]) ? 4'b1000 : 4'b1100;
																assign node24629 = (inp[9]) ? 4'b1100 : 4'b1000;
															assign node24632 = (inp[9]) ? node24636 : node24633;
																assign node24633 = (inp[4]) ? 4'b1100 : 4'b1000;
																assign node24636 = (inp[4]) ? 4'b1000 : 4'b1100;
														assign node24639 = (inp[10]) ? node24641 : 4'b1100;
															assign node24641 = (inp[4]) ? 4'b1000 : 4'b1100;
									assign node24644 = (inp[4]) ? node24704 : node24645;
										assign node24645 = (inp[9]) ? node24681 : node24646;
											assign node24646 = (inp[10]) ? node24666 : node24647;
												assign node24647 = (inp[15]) ? node24659 : node24648;
													assign node24648 = (inp[0]) ? node24654 : node24649;
														assign node24649 = (inp[5]) ? node24651 : 4'b1010;
															assign node24651 = (inp[3]) ? 4'b1000 : 4'b1010;
														assign node24654 = (inp[5]) ? node24656 : 4'b1000;
															assign node24656 = (inp[3]) ? 4'b1010 : 4'b1000;
													assign node24659 = (inp[0]) ? node24661 : 4'b1000;
														assign node24661 = (inp[5]) ? node24663 : 4'b1010;
															assign node24663 = (inp[3]) ? 4'b1000 : 4'b1010;
												assign node24666 = (inp[15]) ? node24676 : node24667;
													assign node24667 = (inp[0]) ? node24671 : node24668;
														assign node24668 = (inp[5]) ? 4'b1000 : 4'b1010;
														assign node24671 = (inp[3]) ? node24673 : 4'b1000;
															assign node24673 = (inp[5]) ? 4'b1010 : 4'b1000;
													assign node24676 = (inp[0]) ? 4'b1010 : node24677;
														assign node24677 = (inp[5]) ? 4'b1010 : 4'b1000;
											assign node24681 = (inp[0]) ? node24693 : node24682;
												assign node24682 = (inp[15]) ? node24688 : node24683;
													assign node24683 = (inp[5]) ? 4'b1100 : node24684;
														assign node24684 = (inp[3]) ? 4'b1100 : 4'b1110;
													assign node24688 = (inp[3]) ? 4'b1110 : node24689;
														assign node24689 = (inp[5]) ? 4'b1110 : 4'b1100;
												assign node24693 = (inp[15]) ? node24699 : node24694;
													assign node24694 = (inp[3]) ? 4'b1110 : node24695;
														assign node24695 = (inp[5]) ? 4'b1110 : 4'b1100;
													assign node24699 = (inp[3]) ? 4'b1100 : node24700;
														assign node24700 = (inp[5]) ? 4'b1100 : 4'b1110;
										assign node24704 = (inp[9]) ? node24728 : node24705;
											assign node24705 = (inp[0]) ? node24717 : node24706;
												assign node24706 = (inp[15]) ? node24712 : node24707;
													assign node24707 = (inp[3]) ? 4'b1100 : node24708;
														assign node24708 = (inp[5]) ? 4'b1100 : 4'b1110;
													assign node24712 = (inp[5]) ? 4'b1110 : node24713;
														assign node24713 = (inp[3]) ? 4'b1110 : 4'b1100;
												assign node24717 = (inp[15]) ? node24723 : node24718;
													assign node24718 = (inp[3]) ? 4'b1110 : node24719;
														assign node24719 = (inp[5]) ? 4'b1110 : 4'b1100;
													assign node24723 = (inp[3]) ? 4'b1100 : node24724;
														assign node24724 = (inp[5]) ? 4'b1100 : 4'b1110;
											assign node24728 = (inp[2]) ? node24748 : node24729;
												assign node24729 = (inp[0]) ? node24741 : node24730;
													assign node24730 = (inp[15]) ? node24736 : node24731;
														assign node24731 = (inp[3]) ? 4'b1000 : node24732;
															assign node24732 = (inp[5]) ? 4'b1000 : 4'b1010;
														assign node24736 = (inp[5]) ? 4'b1010 : node24737;
															assign node24737 = (inp[3]) ? 4'b1010 : 4'b1000;
													assign node24741 = (inp[15]) ? 4'b1000 : node24742;
														assign node24742 = (inp[5]) ? 4'b1010 : node24743;
															assign node24743 = (inp[3]) ? 4'b1010 : 4'b1000;
												assign node24748 = (inp[10]) ? node24766 : node24749;
													assign node24749 = (inp[3]) ? node24759 : node24750;
														assign node24750 = (inp[15]) ? 4'b1010 : node24751;
															assign node24751 = (inp[0]) ? node24755 : node24752;
																assign node24752 = (inp[5]) ? 4'b1000 : 4'b1010;
																assign node24755 = (inp[5]) ? 4'b1010 : 4'b1000;
														assign node24759 = (inp[0]) ? node24763 : node24760;
															assign node24760 = (inp[15]) ? 4'b1010 : 4'b1000;
															assign node24763 = (inp[15]) ? 4'b1000 : 4'b1010;
													assign node24766 = (inp[5]) ? node24780 : node24767;
														assign node24767 = (inp[3]) ? node24775 : node24768;
															assign node24768 = (inp[0]) ? node24772 : node24769;
																assign node24769 = (inp[15]) ? 4'b1000 : 4'b1010;
																assign node24772 = (inp[15]) ? 4'b1010 : 4'b1000;
															assign node24775 = (inp[0]) ? node24777 : 4'b1010;
																assign node24777 = (inp[15]) ? 4'b1000 : 4'b1010;
														assign node24780 = (inp[0]) ? 4'b1010 : node24781;
															assign node24781 = (inp[15]) ? 4'b1010 : 4'b1000;
				assign node24785 = (inp[1]) ? node28811 : node24786;
					assign node24786 = (inp[8]) ? node26648 : node24787;
						assign node24787 = (inp[7]) ? node25755 : node24788;
							assign node24788 = (inp[2]) ? node25336 : node24789;
								assign node24789 = (inp[14]) ? node25061 : node24790;
									assign node24790 = (inp[0]) ? node24918 : node24791;
										assign node24791 = (inp[15]) ? node24845 : node24792;
											assign node24792 = (inp[3]) ? node24814 : node24793;
												assign node24793 = (inp[9]) ? node24803 : node24794;
													assign node24794 = (inp[4]) ? node24800 : node24795;
														assign node24795 = (inp[10]) ? node24797 : 4'b0111;
															assign node24797 = (inp[12]) ? 4'b0011 : 4'b0111;
														assign node24800 = (inp[12]) ? 4'b0111 : 4'b0011;
													assign node24803 = (inp[4]) ? node24809 : node24804;
														assign node24804 = (inp[12]) ? node24806 : 4'b0011;
															assign node24806 = (inp[10]) ? 4'b0101 : 4'b0011;
														assign node24809 = (inp[12]) ? 4'b0001 : node24810;
															assign node24810 = (inp[5]) ? 4'b0101 : 4'b0111;
												assign node24814 = (inp[5]) ? node24830 : node24815;
													assign node24815 = (inp[9]) ? node24821 : node24816;
														assign node24816 = (inp[4]) ? 4'b0011 : node24817;
															assign node24817 = (inp[12]) ? 4'b0011 : 4'b0111;
														assign node24821 = (inp[4]) ? node24825 : node24822;
															assign node24822 = (inp[10]) ? 4'b0101 : 4'b0011;
															assign node24825 = (inp[10]) ? node24827 : 4'b0101;
																assign node24827 = (inp[12]) ? 4'b0001 : 4'b0101;
													assign node24830 = (inp[9]) ? node24840 : node24831;
														assign node24831 = (inp[4]) ? node24837 : node24832;
															assign node24832 = (inp[10]) ? node24834 : 4'b0101;
																assign node24834 = (inp[12]) ? 4'b0001 : 4'b0101;
															assign node24837 = (inp[12]) ? 4'b0101 : 4'b0001;
														assign node24840 = (inp[4]) ? node24842 : 4'b0001;
															assign node24842 = (inp[10]) ? 4'b0001 : 4'b0101;
											assign node24845 = (inp[3]) ? node24881 : node24846;
												assign node24846 = (inp[5]) ? node24864 : node24847;
													assign node24847 = (inp[12]) ? node24853 : node24848;
														assign node24848 = (inp[4]) ? 4'b0101 : node24849;
															assign node24849 = (inp[9]) ? 4'b0001 : 4'b0101;
														assign node24853 = (inp[10]) ? node24859 : node24854;
															assign node24854 = (inp[9]) ? 4'b0101 : node24855;
																assign node24855 = (inp[4]) ? 4'b0001 : 4'b0101;
															assign node24859 = (inp[4]) ? node24861 : 4'b0001;
																assign node24861 = (inp[9]) ? 4'b0001 : 4'b0101;
													assign node24864 = (inp[4]) ? node24876 : node24865;
														assign node24865 = (inp[9]) ? node24871 : node24866;
															assign node24866 = (inp[10]) ? node24868 : 4'b0101;
																assign node24868 = (inp[12]) ? 4'b0001 : 4'b0101;
															assign node24871 = (inp[10]) ? node24873 : 4'b0001;
																assign node24873 = (inp[12]) ? 4'b0111 : 4'b0001;
														assign node24876 = (inp[9]) ? 4'b0111 : node24877;
															assign node24877 = (inp[10]) ? 4'b0111 : 4'b0001;
												assign node24881 = (inp[5]) ? node24897 : node24882;
													assign node24882 = (inp[9]) ? node24890 : node24883;
														assign node24883 = (inp[4]) ? node24885 : 4'b0101;
															assign node24885 = (inp[10]) ? node24887 : 4'b0001;
																assign node24887 = (inp[12]) ? 4'b0111 : 4'b0001;
														assign node24890 = (inp[4]) ? node24894 : node24891;
															assign node24891 = (inp[12]) ? 4'b0111 : 4'b0001;
															assign node24894 = (inp[12]) ? 4'b0011 : 4'b0111;
													assign node24897 = (inp[12]) ? node24905 : node24898;
														assign node24898 = (inp[4]) ? node24902 : node24899;
															assign node24899 = (inp[9]) ? 4'b0011 : 4'b0111;
															assign node24902 = (inp[9]) ? 4'b0111 : 4'b0011;
														assign node24905 = (inp[9]) ? node24911 : node24906;
															assign node24906 = (inp[10]) ? node24908 : 4'b0111;
																assign node24908 = (inp[4]) ? 4'b0111 : 4'b0011;
															assign node24911 = (inp[10]) ? node24915 : node24912;
																assign node24912 = (inp[4]) ? 4'b0111 : 4'b0011;
																assign node24915 = (inp[4]) ? 4'b0011 : 4'b0111;
										assign node24918 = (inp[15]) ? node24982 : node24919;
											assign node24919 = (inp[5]) ? node24947 : node24920;
												assign node24920 = (inp[3]) ? node24934 : node24921;
													assign node24921 = (inp[9]) ? node24929 : node24922;
														assign node24922 = (inp[4]) ? 4'b0001 : node24923;
															assign node24923 = (inp[10]) ? node24925 : 4'b0101;
																assign node24925 = (inp[12]) ? 4'b0001 : 4'b0101;
														assign node24929 = (inp[4]) ? 4'b0101 : node24930;
															assign node24930 = (inp[10]) ? 4'b0101 : 4'b0001;
													assign node24934 = (inp[4]) ? node24942 : node24935;
														assign node24935 = (inp[9]) ? node24937 : 4'b0101;
															assign node24937 = (inp[12]) ? node24939 : 4'b0001;
																assign node24939 = (inp[10]) ? 4'b0111 : 4'b0001;
														assign node24942 = (inp[9]) ? 4'b0111 : node24943;
															assign node24943 = (inp[10]) ? 4'b0111 : 4'b0001;
												assign node24947 = (inp[3]) ? node24969 : node24948;
													assign node24948 = (inp[4]) ? node24960 : node24949;
														assign node24949 = (inp[9]) ? node24955 : node24950;
															assign node24950 = (inp[10]) ? node24952 : 4'b0101;
																assign node24952 = (inp[12]) ? 4'b0001 : 4'b0101;
															assign node24955 = (inp[10]) ? node24957 : 4'b0001;
																assign node24957 = (inp[12]) ? 4'b0111 : 4'b0001;
														assign node24960 = (inp[10]) ? node24962 : 4'b0111;
															assign node24962 = (inp[9]) ? node24966 : node24963;
																assign node24963 = (inp[12]) ? 4'b0111 : 4'b0001;
																assign node24966 = (inp[12]) ? 4'b0011 : 4'b0111;
													assign node24969 = (inp[9]) ? node24977 : node24970;
														assign node24970 = (inp[4]) ? 4'b0011 : node24971;
															assign node24971 = (inp[10]) ? node24973 : 4'b0111;
																assign node24973 = (inp[12]) ? 4'b0011 : 4'b0111;
														assign node24977 = (inp[4]) ? 4'b0111 : node24978;
															assign node24978 = (inp[10]) ? 4'b0111 : 4'b0011;
											assign node24982 = (inp[5]) ? node25026 : node24983;
												assign node24983 = (inp[3]) ? node25009 : node24984;
													assign node24984 = (inp[10]) ? node24994 : node24985;
														assign node24985 = (inp[12]) ? node24987 : 4'b0011;
															assign node24987 = (inp[9]) ? node24991 : node24988;
																assign node24988 = (inp[4]) ? 4'b0011 : 4'b0111;
																assign node24991 = (inp[4]) ? 4'b0111 : 4'b0011;
														assign node24994 = (inp[9]) ? node25002 : node24995;
															assign node24995 = (inp[12]) ? node24999 : node24996;
																assign node24996 = (inp[4]) ? 4'b0011 : 4'b0111;
																assign node24999 = (inp[4]) ? 4'b0111 : 4'b0011;
															assign node25002 = (inp[4]) ? node25006 : node25003;
																assign node25003 = (inp[12]) ? 4'b0111 : 4'b0011;
																assign node25006 = (inp[12]) ? 4'b0011 : 4'b0111;
													assign node25009 = (inp[4]) ? node25021 : node25010;
														assign node25010 = (inp[9]) ? node25016 : node25011;
															assign node25011 = (inp[12]) ? node25013 : 4'b0111;
																assign node25013 = (inp[10]) ? 4'b0011 : 4'b0111;
															assign node25016 = (inp[12]) ? node25018 : 4'b0011;
																assign node25018 = (inp[10]) ? 4'b0101 : 4'b0011;
														assign node25021 = (inp[9]) ? 4'b0101 : node25022;
															assign node25022 = (inp[12]) ? 4'b0101 : 4'b0011;
												assign node25026 = (inp[3]) ? node25042 : node25027;
													assign node25027 = (inp[9]) ? node25035 : node25028;
														assign node25028 = (inp[4]) ? 4'b0011 : node25029;
															assign node25029 = (inp[10]) ? node25031 : 4'b0111;
																assign node25031 = (inp[12]) ? 4'b0011 : 4'b0111;
														assign node25035 = (inp[4]) ? node25037 : 4'b0011;
															assign node25037 = (inp[12]) ? node25039 : 4'b0101;
																assign node25039 = (inp[10]) ? 4'b0001 : 4'b0101;
													assign node25042 = (inp[9]) ? node25052 : node25043;
														assign node25043 = (inp[4]) ? node25049 : node25044;
															assign node25044 = (inp[12]) ? node25046 : 4'b0101;
																assign node25046 = (inp[10]) ? 4'b0001 : 4'b0101;
															assign node25049 = (inp[10]) ? 4'b0101 : 4'b0001;
														assign node25052 = (inp[4]) ? node25056 : node25053;
															assign node25053 = (inp[12]) ? 4'b0101 : 4'b0001;
															assign node25056 = (inp[12]) ? node25058 : 4'b0101;
																assign node25058 = (inp[10]) ? 4'b0001 : 4'b0101;
									assign node25061 = (inp[12]) ? node25167 : node25062;
										assign node25062 = (inp[0]) ? node25110 : node25063;
											assign node25063 = (inp[15]) ? node25087 : node25064;
												assign node25064 = (inp[5]) ? node25070 : node25065;
													assign node25065 = (inp[4]) ? node25067 : 4'b0110;
														assign node25067 = (inp[9]) ? 4'b0110 : 4'b0010;
													assign node25070 = (inp[3]) ? node25080 : node25071;
														assign node25071 = (inp[10]) ? 4'b0010 : node25072;
															assign node25072 = (inp[4]) ? node25076 : node25073;
																assign node25073 = (inp[9]) ? 4'b0010 : 4'b0110;
																assign node25076 = (inp[9]) ? 4'b0100 : 4'b0010;
														assign node25080 = (inp[4]) ? node25084 : node25081;
															assign node25081 = (inp[9]) ? 4'b0000 : 4'b0100;
															assign node25084 = (inp[9]) ? 4'b0100 : 4'b0000;
												assign node25087 = (inp[5]) ? node25097 : node25088;
													assign node25088 = (inp[10]) ? 4'b0000 : node25089;
														assign node25089 = (inp[4]) ? node25093 : node25090;
															assign node25090 = (inp[9]) ? 4'b0000 : 4'b0100;
															assign node25093 = (inp[3]) ? 4'b0000 : 4'b0100;
													assign node25097 = (inp[3]) ? node25103 : node25098;
														assign node25098 = (inp[9]) ? node25100 : 4'b0000;
															assign node25100 = (inp[4]) ? 4'b0110 : 4'b0000;
														assign node25103 = (inp[4]) ? node25107 : node25104;
															assign node25104 = (inp[9]) ? 4'b0010 : 4'b0110;
															assign node25107 = (inp[9]) ? 4'b0110 : 4'b0010;
											assign node25110 = (inp[15]) ? node25142 : node25111;
												assign node25111 = (inp[3]) ? node25121 : node25112;
													assign node25112 = (inp[4]) ? node25116 : node25113;
														assign node25113 = (inp[9]) ? 4'b0000 : 4'b0100;
														assign node25116 = (inp[9]) ? node25118 : 4'b0000;
															assign node25118 = (inp[5]) ? 4'b0110 : 4'b0100;
													assign node25121 = (inp[5]) ? node25127 : node25122;
														assign node25122 = (inp[10]) ? 4'b0000 : node25123;
															assign node25123 = (inp[4]) ? 4'b0110 : 4'b0100;
														assign node25127 = (inp[10]) ? node25135 : node25128;
															assign node25128 = (inp[4]) ? node25132 : node25129;
																assign node25129 = (inp[9]) ? 4'b0010 : 4'b0110;
																assign node25132 = (inp[9]) ? 4'b0110 : 4'b0010;
															assign node25135 = (inp[4]) ? node25139 : node25136;
																assign node25136 = (inp[9]) ? 4'b0010 : 4'b0110;
																assign node25139 = (inp[9]) ? 4'b0110 : 4'b0010;
												assign node25142 = (inp[3]) ? node25152 : node25143;
													assign node25143 = (inp[9]) ? node25147 : node25144;
														assign node25144 = (inp[4]) ? 4'b0010 : 4'b0110;
														assign node25147 = (inp[4]) ? node25149 : 4'b0010;
															assign node25149 = (inp[5]) ? 4'b0100 : 4'b0110;
													assign node25152 = (inp[5]) ? node25160 : node25153;
														assign node25153 = (inp[9]) ? node25157 : node25154;
															assign node25154 = (inp[4]) ? 4'b0010 : 4'b0110;
															assign node25157 = (inp[4]) ? 4'b0100 : 4'b0010;
														assign node25160 = (inp[4]) ? node25164 : node25161;
															assign node25161 = (inp[9]) ? 4'b0000 : 4'b0100;
															assign node25164 = (inp[9]) ? 4'b0100 : 4'b0000;
										assign node25167 = (inp[15]) ? node25255 : node25168;
											assign node25168 = (inp[9]) ? node25218 : node25169;
												assign node25169 = (inp[5]) ? node25193 : node25170;
													assign node25170 = (inp[0]) ? node25178 : node25171;
														assign node25171 = (inp[10]) ? node25175 : node25172;
															assign node25172 = (inp[4]) ? 4'b0010 : 4'b0110;
															assign node25175 = (inp[3]) ? 4'b0100 : 4'b0110;
														assign node25178 = (inp[3]) ? node25186 : node25179;
															assign node25179 = (inp[4]) ? node25183 : node25180;
																assign node25180 = (inp[10]) ? 4'b0000 : 4'b0100;
																assign node25183 = (inp[10]) ? 4'b0100 : 4'b0000;
															assign node25186 = (inp[10]) ? node25190 : node25187;
																assign node25187 = (inp[4]) ? 4'b0000 : 4'b0100;
																assign node25190 = (inp[4]) ? 4'b0110 : 4'b0000;
													assign node25193 = (inp[0]) ? node25207 : node25194;
														assign node25194 = (inp[3]) ? node25202 : node25195;
															assign node25195 = (inp[10]) ? node25199 : node25196;
																assign node25196 = (inp[4]) ? 4'b0010 : 4'b0110;
																assign node25199 = (inp[4]) ? 4'b0100 : 4'b0010;
															assign node25202 = (inp[10]) ? node25204 : 4'b0000;
																assign node25204 = (inp[4]) ? 4'b0100 : 4'b0000;
														assign node25207 = (inp[3]) ? node25211 : node25208;
															assign node25208 = (inp[10]) ? 4'b0110 : 4'b0100;
															assign node25211 = (inp[4]) ? node25215 : node25212;
																assign node25212 = (inp[10]) ? 4'b0010 : 4'b0110;
																assign node25215 = (inp[10]) ? 4'b0110 : 4'b0010;
												assign node25218 = (inp[4]) ? node25234 : node25219;
													assign node25219 = (inp[10]) ? node25231 : node25220;
														assign node25220 = (inp[0]) ? node25226 : node25221;
															assign node25221 = (inp[3]) ? node25223 : 4'b0010;
																assign node25223 = (inp[5]) ? 4'b0000 : 4'b0010;
															assign node25226 = (inp[5]) ? node25228 : 4'b0000;
																assign node25228 = (inp[3]) ? 4'b0010 : 4'b0000;
														assign node25231 = (inp[0]) ? 4'b0110 : 4'b0100;
													assign node25234 = (inp[10]) ? node25244 : node25235;
														assign node25235 = (inp[0]) ? node25241 : node25236;
															assign node25236 = (inp[5]) ? 4'b0100 : node25237;
																assign node25237 = (inp[3]) ? 4'b0100 : 4'b0110;
															assign node25241 = (inp[3]) ? 4'b0110 : 4'b0100;
														assign node25244 = (inp[0]) ? node25250 : node25245;
															assign node25245 = (inp[5]) ? 4'b0000 : node25246;
																assign node25246 = (inp[3]) ? 4'b0000 : 4'b0010;
															assign node25250 = (inp[3]) ? 4'b0010 : node25251;
																assign node25251 = (inp[5]) ? 4'b0010 : 4'b0000;
											assign node25255 = (inp[5]) ? node25299 : node25256;
												assign node25256 = (inp[0]) ? node25284 : node25257;
													assign node25257 = (inp[3]) ? node25271 : node25258;
														assign node25258 = (inp[10]) ? node25264 : node25259;
															assign node25259 = (inp[4]) ? 4'b0100 : node25260;
																assign node25260 = (inp[9]) ? 4'b0000 : 4'b0100;
															assign node25264 = (inp[4]) ? node25268 : node25265;
																assign node25265 = (inp[9]) ? 4'b0100 : 4'b0000;
																assign node25268 = (inp[9]) ? 4'b0000 : 4'b0100;
														assign node25271 = (inp[4]) ? node25279 : node25272;
															assign node25272 = (inp[9]) ? node25276 : node25273;
																assign node25273 = (inp[10]) ? 4'b0000 : 4'b0100;
																assign node25276 = (inp[10]) ? 4'b0110 : 4'b0000;
															assign node25279 = (inp[9]) ? node25281 : 4'b0110;
																assign node25281 = (inp[10]) ? 4'b0010 : 4'b0110;
													assign node25284 = (inp[3]) ? node25292 : node25285;
														assign node25285 = (inp[10]) ? 4'b0110 : node25286;
															assign node25286 = (inp[4]) ? node25288 : 4'b0010;
																assign node25288 = (inp[9]) ? 4'b0110 : 4'b0010;
														assign node25292 = (inp[9]) ? 4'b0100 : node25293;
															assign node25293 = (inp[10]) ? 4'b0100 : node25294;
																assign node25294 = (inp[4]) ? 4'b0010 : 4'b0110;
												assign node25299 = (inp[0]) ? node25315 : node25300;
													assign node25300 = (inp[9]) ? node25308 : node25301;
														assign node25301 = (inp[3]) ? 4'b0110 : node25302;
															assign node25302 = (inp[4]) ? node25304 : 4'b0000;
																assign node25304 = (inp[10]) ? 4'b0110 : 4'b0000;
														assign node25308 = (inp[4]) ? node25312 : node25309;
															assign node25309 = (inp[10]) ? 4'b0110 : 4'b0010;
															assign node25312 = (inp[10]) ? 4'b0010 : 4'b0110;
													assign node25315 = (inp[3]) ? node25327 : node25316;
														assign node25316 = (inp[4]) ? node25322 : node25317;
															assign node25317 = (inp[10]) ? 4'b0010 : node25318;
																assign node25318 = (inp[9]) ? 4'b0010 : 4'b0110;
															assign node25322 = (inp[9]) ? 4'b0100 : node25323;
																assign node25323 = (inp[10]) ? 4'b0100 : 4'b0010;
														assign node25327 = (inp[9]) ? 4'b0100 : node25328;
															assign node25328 = (inp[4]) ? node25332 : node25329;
																assign node25329 = (inp[10]) ? 4'b0000 : 4'b0100;
																assign node25332 = (inp[10]) ? 4'b0100 : 4'b0000;
								assign node25336 = (inp[15]) ? node25556 : node25337;
									assign node25337 = (inp[0]) ? node25443 : node25338;
										assign node25338 = (inp[5]) ? node25396 : node25339;
											assign node25339 = (inp[3]) ? node25373 : node25340;
												assign node25340 = (inp[12]) ? node25348 : node25341;
													assign node25341 = (inp[9]) ? node25345 : node25342;
														assign node25342 = (inp[4]) ? 4'b0010 : 4'b0110;
														assign node25345 = (inp[4]) ? 4'b0110 : 4'b0010;
													assign node25348 = (inp[14]) ? node25358 : node25349;
														assign node25349 = (inp[9]) ? node25351 : 4'b0010;
															assign node25351 = (inp[10]) ? node25355 : node25352;
																assign node25352 = (inp[4]) ? 4'b0110 : 4'b0010;
																assign node25355 = (inp[4]) ? 4'b0010 : 4'b0110;
														assign node25358 = (inp[9]) ? node25366 : node25359;
															assign node25359 = (inp[10]) ? node25363 : node25360;
																assign node25360 = (inp[4]) ? 4'b0010 : 4'b0110;
																assign node25363 = (inp[4]) ? 4'b0110 : 4'b0010;
															assign node25366 = (inp[10]) ? node25370 : node25367;
																assign node25367 = (inp[4]) ? 4'b0110 : 4'b0010;
																assign node25370 = (inp[4]) ? 4'b0010 : 4'b0110;
												assign node25373 = (inp[9]) ? node25385 : node25374;
													assign node25374 = (inp[4]) ? node25380 : node25375;
														assign node25375 = (inp[10]) ? node25377 : 4'b0110;
															assign node25377 = (inp[12]) ? 4'b0010 : 4'b0110;
														assign node25380 = (inp[12]) ? node25382 : 4'b0010;
															assign node25382 = (inp[14]) ? 4'b0100 : 4'b0010;
													assign node25385 = (inp[4]) ? node25391 : node25386;
														assign node25386 = (inp[12]) ? node25388 : 4'b0010;
															assign node25388 = (inp[10]) ? 4'b0100 : 4'b0010;
														assign node25391 = (inp[12]) ? node25393 : 4'b0100;
															assign node25393 = (inp[10]) ? 4'b0000 : 4'b0100;
											assign node25396 = (inp[3]) ? node25420 : node25397;
												assign node25397 = (inp[9]) ? node25409 : node25398;
													assign node25398 = (inp[4]) ? node25404 : node25399;
														assign node25399 = (inp[10]) ? node25401 : 4'b0110;
															assign node25401 = (inp[12]) ? 4'b0010 : 4'b0110;
														assign node25404 = (inp[12]) ? node25406 : 4'b0010;
															assign node25406 = (inp[10]) ? 4'b0100 : 4'b0010;
													assign node25409 = (inp[4]) ? node25415 : node25410;
														assign node25410 = (inp[12]) ? node25412 : 4'b0010;
															assign node25412 = (inp[10]) ? 4'b0100 : 4'b0010;
														assign node25415 = (inp[12]) ? node25417 : 4'b0100;
															assign node25417 = (inp[10]) ? 4'b0000 : 4'b0100;
												assign node25420 = (inp[9]) ? node25432 : node25421;
													assign node25421 = (inp[4]) ? node25427 : node25422;
														assign node25422 = (inp[12]) ? node25424 : 4'b0100;
															assign node25424 = (inp[10]) ? 4'b0000 : 4'b0100;
														assign node25427 = (inp[12]) ? node25429 : 4'b0000;
															assign node25429 = (inp[10]) ? 4'b0100 : 4'b0000;
													assign node25432 = (inp[4]) ? node25438 : node25433;
														assign node25433 = (inp[12]) ? node25435 : 4'b0000;
															assign node25435 = (inp[10]) ? 4'b0100 : 4'b0000;
														assign node25438 = (inp[12]) ? node25440 : 4'b0100;
															assign node25440 = (inp[14]) ? 4'b0000 : 4'b0100;
										assign node25443 = (inp[5]) ? node25497 : node25444;
											assign node25444 = (inp[3]) ? node25476 : node25445;
												assign node25445 = (inp[12]) ? node25461 : node25446;
													assign node25446 = (inp[10]) ? node25454 : node25447;
														assign node25447 = (inp[9]) ? node25451 : node25448;
															assign node25448 = (inp[4]) ? 4'b0000 : 4'b0100;
															assign node25451 = (inp[4]) ? 4'b0100 : 4'b0000;
														assign node25454 = (inp[9]) ? node25458 : node25455;
															assign node25455 = (inp[4]) ? 4'b0000 : 4'b0100;
															assign node25458 = (inp[4]) ? 4'b0100 : 4'b0000;
													assign node25461 = (inp[4]) ? node25469 : node25462;
														assign node25462 = (inp[9]) ? node25466 : node25463;
															assign node25463 = (inp[10]) ? 4'b0000 : 4'b0100;
															assign node25466 = (inp[10]) ? 4'b0100 : 4'b0000;
														assign node25469 = (inp[10]) ? node25473 : node25470;
															assign node25470 = (inp[9]) ? 4'b0100 : 4'b0000;
															assign node25473 = (inp[9]) ? 4'b0000 : 4'b0100;
												assign node25476 = (inp[10]) ? node25482 : node25477;
													assign node25477 = (inp[4]) ? 4'b0000 : node25478;
														assign node25478 = (inp[9]) ? 4'b0000 : 4'b0100;
													assign node25482 = (inp[12]) ? node25490 : node25483;
														assign node25483 = (inp[9]) ? node25487 : node25484;
															assign node25484 = (inp[4]) ? 4'b0000 : 4'b0100;
															assign node25487 = (inp[4]) ? 4'b0110 : 4'b0000;
														assign node25490 = (inp[4]) ? node25494 : node25491;
															assign node25491 = (inp[9]) ? 4'b0110 : 4'b0000;
															assign node25494 = (inp[9]) ? 4'b0010 : 4'b0110;
											assign node25497 = (inp[3]) ? node25519 : node25498;
												assign node25498 = (inp[4]) ? node25510 : node25499;
													assign node25499 = (inp[9]) ? node25505 : node25500;
														assign node25500 = (inp[12]) ? node25502 : 4'b0100;
															assign node25502 = (inp[10]) ? 4'b0000 : 4'b0100;
														assign node25505 = (inp[10]) ? node25507 : 4'b0000;
															assign node25507 = (inp[12]) ? 4'b0110 : 4'b0000;
													assign node25510 = (inp[9]) ? node25516 : node25511;
														assign node25511 = (inp[12]) ? node25513 : 4'b0000;
															assign node25513 = (inp[10]) ? 4'b0110 : 4'b0000;
														assign node25516 = (inp[10]) ? 4'b0010 : 4'b0110;
												assign node25519 = (inp[14]) ? node25537 : node25520;
													assign node25520 = (inp[12]) ? node25528 : node25521;
														assign node25521 = (inp[4]) ? node25525 : node25522;
															assign node25522 = (inp[9]) ? 4'b0010 : 4'b0110;
															assign node25525 = (inp[9]) ? 4'b0110 : 4'b0010;
														assign node25528 = (inp[10]) ? node25530 : 4'b0110;
															assign node25530 = (inp[9]) ? node25534 : node25531;
																assign node25531 = (inp[4]) ? 4'b0110 : 4'b0010;
																assign node25534 = (inp[4]) ? 4'b0010 : 4'b0110;
													assign node25537 = (inp[9]) ? node25547 : node25538;
														assign node25538 = (inp[4]) ? node25544 : node25539;
															assign node25539 = (inp[12]) ? node25541 : 4'b0110;
																assign node25541 = (inp[10]) ? 4'b0010 : 4'b0110;
															assign node25544 = (inp[10]) ? 4'b0110 : 4'b0010;
														assign node25547 = (inp[4]) ? node25553 : node25548;
															assign node25548 = (inp[12]) ? node25550 : 4'b0010;
																assign node25550 = (inp[10]) ? 4'b0110 : 4'b0010;
															assign node25553 = (inp[10]) ? 4'b0010 : 4'b0110;
									assign node25556 = (inp[0]) ? node25652 : node25557;
										assign node25557 = (inp[3]) ? node25607 : node25558;
											assign node25558 = (inp[5]) ? node25584 : node25559;
												assign node25559 = (inp[4]) ? node25571 : node25560;
													assign node25560 = (inp[9]) ? node25566 : node25561;
														assign node25561 = (inp[10]) ? node25563 : 4'b0100;
															assign node25563 = (inp[12]) ? 4'b0000 : 4'b0100;
														assign node25566 = (inp[10]) ? node25568 : 4'b0000;
															assign node25568 = (inp[14]) ? 4'b0000 : 4'b0100;
													assign node25571 = (inp[12]) ? node25573 : 4'b0000;
														assign node25573 = (inp[14]) ? node25579 : node25574;
															assign node25574 = (inp[9]) ? node25576 : 4'b0000;
																assign node25576 = (inp[10]) ? 4'b0000 : 4'b0100;
															assign node25579 = (inp[9]) ? 4'b0100 : node25580;
																assign node25580 = (inp[10]) ? 4'b0100 : 4'b0000;
												assign node25584 = (inp[4]) ? node25596 : node25585;
													assign node25585 = (inp[9]) ? node25591 : node25586;
														assign node25586 = (inp[12]) ? node25588 : 4'b0100;
															assign node25588 = (inp[10]) ? 4'b0000 : 4'b0100;
														assign node25591 = (inp[10]) ? node25593 : 4'b0000;
															assign node25593 = (inp[12]) ? 4'b0110 : 4'b0000;
													assign node25596 = (inp[9]) ? node25602 : node25597;
														assign node25597 = (inp[10]) ? node25599 : 4'b0000;
															assign node25599 = (inp[12]) ? 4'b0110 : 4'b0000;
														assign node25602 = (inp[12]) ? node25604 : 4'b0110;
															assign node25604 = (inp[10]) ? 4'b0010 : 4'b0110;
											assign node25607 = (inp[5]) ? node25629 : node25608;
												assign node25608 = (inp[4]) ? node25620 : node25609;
													assign node25609 = (inp[9]) ? node25615 : node25610;
														assign node25610 = (inp[12]) ? node25612 : 4'b0100;
															assign node25612 = (inp[10]) ? 4'b0000 : 4'b0100;
														assign node25615 = (inp[10]) ? node25617 : 4'b0000;
															assign node25617 = (inp[12]) ? 4'b0110 : 4'b0000;
													assign node25620 = (inp[9]) ? node25624 : node25621;
														assign node25621 = (inp[12]) ? 4'b0110 : 4'b0000;
														assign node25624 = (inp[10]) ? node25626 : 4'b0110;
															assign node25626 = (inp[12]) ? 4'b0010 : 4'b0110;
												assign node25629 = (inp[4]) ? node25641 : node25630;
													assign node25630 = (inp[9]) ? node25636 : node25631;
														assign node25631 = (inp[10]) ? node25633 : 4'b0110;
															assign node25633 = (inp[12]) ? 4'b0010 : 4'b0110;
														assign node25636 = (inp[12]) ? node25638 : 4'b0010;
															assign node25638 = (inp[10]) ? 4'b0110 : 4'b0010;
													assign node25641 = (inp[9]) ? node25647 : node25642;
														assign node25642 = (inp[10]) ? node25644 : 4'b0010;
															assign node25644 = (inp[12]) ? 4'b0110 : 4'b0010;
														assign node25647 = (inp[10]) ? node25649 : 4'b0110;
															assign node25649 = (inp[12]) ? 4'b0010 : 4'b0110;
										assign node25652 = (inp[3]) ? node25696 : node25653;
											assign node25653 = (inp[5]) ? node25673 : node25654;
												assign node25654 = (inp[4]) ? node25666 : node25655;
													assign node25655 = (inp[9]) ? node25661 : node25656;
														assign node25656 = (inp[12]) ? node25658 : 4'b0110;
															assign node25658 = (inp[10]) ? 4'b0010 : 4'b0110;
														assign node25661 = (inp[12]) ? node25663 : 4'b0010;
															assign node25663 = (inp[10]) ? 4'b0110 : 4'b0010;
													assign node25666 = (inp[9]) ? 4'b0110 : node25667;
														assign node25667 = (inp[10]) ? node25669 : 4'b0010;
															assign node25669 = (inp[12]) ? 4'b0110 : 4'b0010;
												assign node25673 = (inp[4]) ? node25685 : node25674;
													assign node25674 = (inp[9]) ? node25680 : node25675;
														assign node25675 = (inp[12]) ? node25677 : 4'b0110;
															assign node25677 = (inp[10]) ? 4'b0010 : 4'b0110;
														assign node25680 = (inp[12]) ? node25682 : 4'b0010;
															assign node25682 = (inp[10]) ? 4'b0100 : 4'b0010;
													assign node25685 = (inp[9]) ? node25691 : node25686;
														assign node25686 = (inp[10]) ? node25688 : 4'b0010;
															assign node25688 = (inp[12]) ? 4'b0100 : 4'b0010;
														assign node25691 = (inp[12]) ? node25693 : 4'b0100;
															assign node25693 = (inp[14]) ? 4'b0000 : 4'b0100;
											assign node25696 = (inp[5]) ? node25720 : node25697;
												assign node25697 = (inp[9]) ? node25709 : node25698;
													assign node25698 = (inp[4]) ? node25704 : node25699;
														assign node25699 = (inp[10]) ? node25701 : 4'b0110;
															assign node25701 = (inp[12]) ? 4'b0010 : 4'b0110;
														assign node25704 = (inp[10]) ? node25706 : 4'b0010;
															assign node25706 = (inp[12]) ? 4'b0100 : 4'b0010;
													assign node25709 = (inp[4]) ? node25715 : node25710;
														assign node25710 = (inp[10]) ? node25712 : 4'b0010;
															assign node25712 = (inp[12]) ? 4'b0100 : 4'b0010;
														assign node25715 = (inp[12]) ? node25717 : 4'b0100;
															assign node25717 = (inp[10]) ? 4'b0000 : 4'b0100;
												assign node25720 = (inp[10]) ? node25740 : node25721;
													assign node25721 = (inp[12]) ? node25729 : node25722;
														assign node25722 = (inp[9]) ? node25726 : node25723;
															assign node25723 = (inp[4]) ? 4'b0000 : 4'b0100;
															assign node25726 = (inp[4]) ? 4'b0100 : 4'b0000;
														assign node25729 = (inp[14]) ? node25735 : node25730;
															assign node25730 = (inp[9]) ? node25732 : 4'b0100;
																assign node25732 = (inp[4]) ? 4'b0100 : 4'b0000;
															assign node25735 = (inp[4]) ? node25737 : 4'b0000;
																assign node25737 = (inp[9]) ? 4'b0100 : 4'b0000;
													assign node25740 = (inp[12]) ? node25748 : node25741;
														assign node25741 = (inp[4]) ? node25745 : node25742;
															assign node25742 = (inp[9]) ? 4'b0000 : 4'b0100;
															assign node25745 = (inp[14]) ? 4'b0100 : 4'b0000;
														assign node25748 = (inp[4]) ? node25752 : node25749;
															assign node25749 = (inp[9]) ? 4'b0100 : 4'b0000;
															assign node25752 = (inp[9]) ? 4'b0000 : 4'b0100;
							assign node25755 = (inp[14]) ? node26287 : node25756;
								assign node25756 = (inp[2]) ? node26036 : node25757;
									assign node25757 = (inp[0]) ? node25911 : node25758;
										assign node25758 = (inp[15]) ? node25834 : node25759;
											assign node25759 = (inp[5]) ? node25799 : node25760;
												assign node25760 = (inp[3]) ? node25784 : node25761;
													assign node25761 = (inp[10]) ? node25775 : node25762;
														assign node25762 = (inp[12]) ? node25768 : node25763;
															assign node25763 = (inp[9]) ? 4'b0110 : node25764;
																assign node25764 = (inp[4]) ? 4'b0010 : 4'b0110;
															assign node25768 = (inp[9]) ? node25772 : node25769;
																assign node25769 = (inp[4]) ? 4'b0010 : 4'b0110;
																assign node25772 = (inp[4]) ? 4'b0110 : 4'b0010;
														assign node25775 = (inp[4]) ? node25777 : 4'b0010;
															assign node25777 = (inp[9]) ? node25781 : node25778;
																assign node25778 = (inp[12]) ? 4'b0110 : 4'b0010;
																assign node25781 = (inp[12]) ? 4'b0010 : 4'b0110;
													assign node25784 = (inp[9]) ? node25794 : node25785;
														assign node25785 = (inp[4]) ? node25789 : node25786;
															assign node25786 = (inp[10]) ? 4'b0010 : 4'b0110;
															assign node25789 = (inp[10]) ? node25791 : 4'b0010;
																assign node25791 = (inp[12]) ? 4'b0100 : 4'b0010;
														assign node25794 = (inp[4]) ? 4'b0100 : node25795;
															assign node25795 = (inp[12]) ? 4'b0100 : 4'b0010;
												assign node25799 = (inp[3]) ? node25817 : node25800;
													assign node25800 = (inp[4]) ? node25808 : node25801;
														assign node25801 = (inp[9]) ? 4'b0010 : node25802;
															assign node25802 = (inp[12]) ? node25804 : 4'b0110;
																assign node25804 = (inp[10]) ? 4'b0010 : 4'b0110;
														assign node25808 = (inp[9]) ? node25812 : node25809;
															assign node25809 = (inp[12]) ? 4'b0100 : 4'b0010;
															assign node25812 = (inp[10]) ? node25814 : 4'b0100;
																assign node25814 = (inp[12]) ? 4'b0000 : 4'b0100;
													assign node25817 = (inp[9]) ? node25829 : node25818;
														assign node25818 = (inp[4]) ? node25824 : node25819;
															assign node25819 = (inp[12]) ? node25821 : 4'b0100;
																assign node25821 = (inp[10]) ? 4'b0000 : 4'b0100;
															assign node25824 = (inp[12]) ? node25826 : 4'b0000;
																assign node25826 = (inp[10]) ? 4'b0100 : 4'b0000;
														assign node25829 = (inp[4]) ? node25831 : 4'b0000;
															assign node25831 = (inp[12]) ? 4'b0000 : 4'b0100;
											assign node25834 = (inp[5]) ? node25866 : node25835;
												assign node25835 = (inp[9]) ? node25847 : node25836;
													assign node25836 = (inp[4]) ? node25842 : node25837;
														assign node25837 = (inp[12]) ? node25839 : 4'b0100;
															assign node25839 = (inp[10]) ? 4'b0000 : 4'b0100;
														assign node25842 = (inp[10]) ? node25844 : 4'b0000;
															assign node25844 = (inp[12]) ? 4'b0100 : 4'b0000;
													assign node25847 = (inp[3]) ? node25855 : node25848;
														assign node25848 = (inp[12]) ? node25850 : 4'b0100;
															assign node25850 = (inp[4]) ? 4'b0000 : node25851;
																assign node25851 = (inp[10]) ? 4'b0100 : 4'b0000;
														assign node25855 = (inp[4]) ? node25861 : node25856;
															assign node25856 = (inp[10]) ? node25858 : 4'b0000;
																assign node25858 = (inp[12]) ? 4'b0110 : 4'b0000;
															assign node25861 = (inp[12]) ? node25863 : 4'b0110;
																assign node25863 = (inp[10]) ? 4'b0010 : 4'b0110;
												assign node25866 = (inp[3]) ? node25888 : node25867;
													assign node25867 = (inp[4]) ? node25879 : node25868;
														assign node25868 = (inp[9]) ? node25874 : node25869;
															assign node25869 = (inp[12]) ? node25871 : 4'b0100;
																assign node25871 = (inp[10]) ? 4'b0000 : 4'b0100;
															assign node25874 = (inp[10]) ? node25876 : 4'b0000;
																assign node25876 = (inp[12]) ? 4'b0110 : 4'b0000;
														assign node25879 = (inp[9]) ? node25883 : node25880;
															assign node25880 = (inp[12]) ? 4'b0110 : 4'b0000;
															assign node25883 = (inp[10]) ? node25885 : 4'b0110;
																assign node25885 = (inp[12]) ? 4'b0010 : 4'b0110;
													assign node25888 = (inp[12]) ? node25898 : node25889;
														assign node25889 = (inp[10]) ? 4'b0110 : node25890;
															assign node25890 = (inp[4]) ? node25894 : node25891;
																assign node25891 = (inp[9]) ? 4'b0010 : 4'b0110;
																assign node25894 = (inp[9]) ? 4'b0110 : 4'b0010;
														assign node25898 = (inp[4]) ? node25906 : node25899;
															assign node25899 = (inp[9]) ? node25903 : node25900;
																assign node25900 = (inp[10]) ? 4'b0010 : 4'b0110;
																assign node25903 = (inp[10]) ? 4'b0110 : 4'b0010;
															assign node25906 = (inp[10]) ? node25908 : 4'b0010;
																assign node25908 = (inp[9]) ? 4'b0010 : 4'b0110;
										assign node25911 = (inp[5]) ? node25967 : node25912;
											assign node25912 = (inp[15]) ? node25944 : node25913;
												assign node25913 = (inp[10]) ? node25921 : node25914;
													assign node25914 = (inp[4]) ? node25918 : node25915;
														assign node25915 = (inp[9]) ? 4'b0000 : 4'b0100;
														assign node25918 = (inp[9]) ? 4'b0100 : 4'b0000;
													assign node25921 = (inp[3]) ? node25935 : node25922;
														assign node25922 = (inp[12]) ? node25928 : node25923;
															assign node25923 = (inp[4]) ? node25925 : 4'b0000;
																assign node25925 = (inp[9]) ? 4'b0100 : 4'b0000;
															assign node25928 = (inp[9]) ? node25932 : node25929;
																assign node25929 = (inp[4]) ? 4'b0100 : 4'b0000;
																assign node25932 = (inp[4]) ? 4'b0000 : 4'b0100;
														assign node25935 = (inp[4]) ? 4'b0110 : node25936;
															assign node25936 = (inp[12]) ? node25940 : node25937;
																assign node25937 = (inp[9]) ? 4'b0000 : 4'b0100;
																assign node25940 = (inp[9]) ? 4'b0110 : 4'b0000;
												assign node25944 = (inp[4]) ? node25952 : node25945;
													assign node25945 = (inp[9]) ? node25949 : node25946;
														assign node25946 = (inp[10]) ? 4'b0010 : 4'b0110;
														assign node25949 = (inp[10]) ? 4'b0110 : 4'b0010;
													assign node25952 = (inp[3]) ? node25960 : node25953;
														assign node25953 = (inp[10]) ? node25955 : 4'b0010;
															assign node25955 = (inp[9]) ? 4'b0010 : node25956;
																assign node25956 = (inp[12]) ? 4'b0110 : 4'b0010;
														assign node25960 = (inp[9]) ? node25964 : node25961;
															assign node25961 = (inp[12]) ? 4'b0100 : 4'b0010;
															assign node25964 = (inp[12]) ? 4'b0000 : 4'b0100;
											assign node25967 = (inp[15]) ? node26005 : node25968;
												assign node25968 = (inp[3]) ? node25988 : node25969;
													assign node25969 = (inp[9]) ? node25977 : node25970;
														assign node25970 = (inp[4]) ? node25972 : 4'b0100;
															assign node25972 = (inp[12]) ? node25974 : 4'b0000;
																assign node25974 = (inp[10]) ? 4'b0110 : 4'b0000;
														assign node25977 = (inp[4]) ? node25983 : node25978;
															assign node25978 = (inp[12]) ? node25980 : 4'b0000;
																assign node25980 = (inp[10]) ? 4'b0110 : 4'b0000;
															assign node25983 = (inp[12]) ? node25985 : 4'b0110;
																assign node25985 = (inp[10]) ? 4'b0010 : 4'b0110;
													assign node25988 = (inp[9]) ? node26000 : node25989;
														assign node25989 = (inp[4]) ? node25995 : node25990;
															assign node25990 = (inp[12]) ? node25992 : 4'b0110;
																assign node25992 = (inp[10]) ? 4'b0010 : 4'b0110;
															assign node25995 = (inp[12]) ? node25997 : 4'b0010;
																assign node25997 = (inp[10]) ? 4'b0110 : 4'b0010;
														assign node26000 = (inp[4]) ? 4'b0110 : node26001;
															assign node26001 = (inp[12]) ? 4'b0110 : 4'b0010;
												assign node26005 = (inp[3]) ? node26019 : node26006;
													assign node26006 = (inp[4]) ? 4'b0100 : node26007;
														assign node26007 = (inp[9]) ? node26013 : node26008;
															assign node26008 = (inp[12]) ? node26010 : 4'b0110;
																assign node26010 = (inp[10]) ? 4'b0010 : 4'b0110;
															assign node26013 = (inp[12]) ? node26015 : 4'b0010;
																assign node26015 = (inp[10]) ? 4'b0100 : 4'b0010;
													assign node26019 = (inp[10]) ? node26027 : node26020;
														assign node26020 = (inp[4]) ? node26024 : node26021;
															assign node26021 = (inp[9]) ? 4'b0000 : 4'b0100;
															assign node26024 = (inp[9]) ? 4'b0100 : 4'b0000;
														assign node26027 = (inp[12]) ? node26029 : 4'b0000;
															assign node26029 = (inp[4]) ? node26033 : node26030;
																assign node26030 = (inp[9]) ? 4'b0100 : 4'b0000;
																assign node26033 = (inp[9]) ? 4'b0000 : 4'b0100;
									assign node26036 = (inp[3]) ? node26178 : node26037;
										assign node26037 = (inp[4]) ? node26103 : node26038;
											assign node26038 = (inp[9]) ? node26070 : node26039;
												assign node26039 = (inp[10]) ? node26055 : node26040;
													assign node26040 = (inp[12]) ? node26048 : node26041;
														assign node26041 = (inp[0]) ? node26045 : node26042;
															assign node26042 = (inp[15]) ? 4'b1101 : 4'b1111;
															assign node26045 = (inp[15]) ? 4'b1111 : 4'b1101;
														assign node26048 = (inp[15]) ? node26052 : node26049;
															assign node26049 = (inp[0]) ? 4'b1001 : 4'b1011;
															assign node26052 = (inp[0]) ? 4'b1011 : 4'b1001;
													assign node26055 = (inp[5]) ? node26063 : node26056;
														assign node26056 = (inp[15]) ? node26060 : node26057;
															assign node26057 = (inp[0]) ? 4'b1001 : 4'b1011;
															assign node26060 = (inp[0]) ? 4'b1011 : 4'b1001;
														assign node26063 = (inp[15]) ? node26067 : node26064;
															assign node26064 = (inp[0]) ? 4'b1001 : 4'b1011;
															assign node26067 = (inp[0]) ? 4'b1011 : 4'b1001;
												assign node26070 = (inp[12]) ? node26082 : node26071;
													assign node26071 = (inp[10]) ? node26077 : node26072;
														assign node26072 = (inp[0]) ? 4'b1001 : node26073;
															assign node26073 = (inp[15]) ? 4'b1001 : 4'b1011;
														assign node26077 = (inp[15]) ? 4'b1101 : node26078;
															assign node26078 = (inp[5]) ? 4'b1101 : 4'b1111;
													assign node26082 = (inp[15]) ? node26096 : node26083;
														assign node26083 = (inp[10]) ? node26089 : node26084;
															assign node26084 = (inp[0]) ? 4'b1101 : node26085;
																assign node26085 = (inp[5]) ? 4'b1101 : 4'b1111;
															assign node26089 = (inp[0]) ? node26093 : node26090;
																assign node26090 = (inp[5]) ? 4'b1101 : 4'b1111;
																assign node26093 = (inp[5]) ? 4'b1111 : 4'b1101;
														assign node26096 = (inp[5]) ? node26100 : node26097;
															assign node26097 = (inp[0]) ? 4'b1111 : 4'b1101;
															assign node26100 = (inp[0]) ? 4'b1101 : 4'b1111;
											assign node26103 = (inp[9]) ? node26141 : node26104;
												assign node26104 = (inp[10]) ? node26118 : node26105;
													assign node26105 = (inp[12]) ? node26113 : node26106;
														assign node26106 = (inp[0]) ? node26110 : node26107;
															assign node26107 = (inp[15]) ? 4'b1001 : 4'b1011;
															assign node26110 = (inp[15]) ? 4'b1011 : 4'b1001;
														assign node26113 = (inp[0]) ? 4'b1101 : node26114;
															assign node26114 = (inp[5]) ? 4'b1101 : 4'b1111;
													assign node26118 = (inp[12]) ? node26128 : node26119;
														assign node26119 = (inp[0]) ? node26121 : 4'b1111;
															assign node26121 = (inp[15]) ? node26125 : node26122;
																assign node26122 = (inp[5]) ? 4'b1111 : 4'b1101;
																assign node26125 = (inp[5]) ? 4'b1101 : 4'b1111;
														assign node26128 = (inp[0]) ? node26134 : node26129;
															assign node26129 = (inp[5]) ? node26131 : 4'b1101;
																assign node26131 = (inp[15]) ? 4'b1111 : 4'b1101;
															assign node26134 = (inp[5]) ? node26138 : node26135;
																assign node26135 = (inp[15]) ? 4'b1111 : 4'b1101;
																assign node26138 = (inp[15]) ? 4'b1101 : 4'b1111;
												assign node26141 = (inp[10]) ? node26163 : node26142;
													assign node26142 = (inp[12]) ? node26150 : node26143;
														assign node26143 = (inp[5]) ? 4'b1111 : node26144;
															assign node26144 = (inp[15]) ? 4'b1101 : node26145;
																assign node26145 = (inp[0]) ? 4'b1101 : 4'b1111;
														assign node26150 = (inp[0]) ? node26158 : node26151;
															assign node26151 = (inp[15]) ? node26155 : node26152;
																assign node26152 = (inp[5]) ? 4'b1001 : 4'b1011;
																assign node26155 = (inp[5]) ? 4'b1011 : 4'b1001;
															assign node26158 = (inp[5]) ? node26160 : 4'b1011;
																assign node26160 = (inp[15]) ? 4'b1001 : 4'b1011;
													assign node26163 = (inp[5]) ? node26171 : node26164;
														assign node26164 = (inp[15]) ? node26168 : node26165;
															assign node26165 = (inp[0]) ? 4'b1001 : 4'b1011;
															assign node26168 = (inp[0]) ? 4'b1011 : 4'b1001;
														assign node26171 = (inp[0]) ? node26175 : node26172;
															assign node26172 = (inp[15]) ? 4'b1011 : 4'b1001;
															assign node26175 = (inp[15]) ? 4'b1001 : 4'b1011;
										assign node26178 = (inp[9]) ? node26234 : node26179;
											assign node26179 = (inp[4]) ? node26211 : node26180;
												assign node26180 = (inp[12]) ? node26198 : node26181;
													assign node26181 = (inp[10]) ? node26193 : node26182;
														assign node26182 = (inp[0]) ? node26188 : node26183;
															assign node26183 = (inp[15]) ? node26185 : 4'b1111;
																assign node26185 = (inp[5]) ? 4'b1111 : 4'b1101;
															assign node26188 = (inp[5]) ? 4'b1101 : node26189;
																assign node26189 = (inp[15]) ? 4'b1111 : 4'b1101;
														assign node26193 = (inp[15]) ? node26195 : 4'b1011;
															assign node26195 = (inp[0]) ? 4'b1011 : 4'b1001;
													assign node26198 = (inp[0]) ? node26204 : node26199;
														assign node26199 = (inp[5]) ? 4'b1011 : node26200;
															assign node26200 = (inp[15]) ? 4'b1001 : 4'b1011;
														assign node26204 = (inp[5]) ? node26208 : node26205;
															assign node26205 = (inp[15]) ? 4'b1011 : 4'b1001;
															assign node26208 = (inp[15]) ? 4'b1001 : 4'b1011;
												assign node26211 = (inp[10]) ? node26227 : node26212;
													assign node26212 = (inp[12]) ? node26222 : node26213;
														assign node26213 = (inp[5]) ? node26215 : 4'b1011;
															assign node26215 = (inp[15]) ? node26219 : node26216;
																assign node26216 = (inp[0]) ? 4'b1011 : 4'b1001;
																assign node26219 = (inp[0]) ? 4'b1001 : 4'b1011;
														assign node26222 = (inp[0]) ? node26224 : 4'b1111;
															assign node26224 = (inp[15]) ? 4'b1101 : 4'b1111;
													assign node26227 = (inp[0]) ? node26231 : node26228;
														assign node26228 = (inp[15]) ? 4'b1111 : 4'b1101;
														assign node26231 = (inp[15]) ? 4'b1101 : 4'b1111;
											assign node26234 = (inp[4]) ? node26266 : node26235;
												assign node26235 = (inp[10]) ? node26251 : node26236;
													assign node26236 = (inp[12]) ? node26244 : node26237;
														assign node26237 = (inp[0]) ? 4'b1001 : node26238;
															assign node26238 = (inp[15]) ? node26240 : 4'b1011;
																assign node26240 = (inp[5]) ? 4'b1011 : 4'b1001;
														assign node26244 = (inp[15]) ? node26248 : node26245;
															assign node26245 = (inp[0]) ? 4'b1111 : 4'b1101;
															assign node26248 = (inp[0]) ? 4'b1101 : 4'b1111;
													assign node26251 = (inp[12]) ? node26259 : node26252;
														assign node26252 = (inp[0]) ? node26256 : node26253;
															assign node26253 = (inp[15]) ? 4'b1111 : 4'b1101;
															assign node26256 = (inp[15]) ? 4'b1101 : 4'b1111;
														assign node26259 = (inp[0]) ? node26263 : node26260;
															assign node26260 = (inp[15]) ? 4'b1111 : 4'b1101;
															assign node26263 = (inp[15]) ? 4'b1101 : 4'b1111;
												assign node26266 = (inp[12]) ? node26280 : node26267;
													assign node26267 = (inp[10]) ? node26273 : node26268;
														assign node26268 = (inp[0]) ? 4'b1111 : node26269;
															assign node26269 = (inp[15]) ? 4'b1111 : 4'b1101;
														assign node26273 = (inp[5]) ? node26275 : 4'b1001;
															assign node26275 = (inp[0]) ? 4'b1011 : node26276;
																assign node26276 = (inp[15]) ? 4'b1011 : 4'b1001;
													assign node26280 = (inp[15]) ? node26284 : node26281;
														assign node26281 = (inp[0]) ? 4'b1011 : 4'b1001;
														assign node26284 = (inp[0]) ? 4'b1001 : 4'b1011;
								assign node26287 = (inp[9]) ? node26485 : node26288;
									assign node26288 = (inp[4]) ? node26398 : node26289;
										assign node26289 = (inp[10]) ? node26353 : node26290;
											assign node26290 = (inp[12]) ? node26310 : node26291;
												assign node26291 = (inp[15]) ? node26299 : node26292;
													assign node26292 = (inp[0]) ? 4'b1101 : node26293;
														assign node26293 = (inp[3]) ? node26295 : 4'b1111;
															assign node26295 = (inp[5]) ? 4'b1101 : 4'b1111;
													assign node26299 = (inp[0]) ? node26305 : node26300;
														assign node26300 = (inp[5]) ? node26302 : 4'b1101;
															assign node26302 = (inp[3]) ? 4'b1111 : 4'b1101;
														assign node26305 = (inp[5]) ? node26307 : 4'b1111;
															assign node26307 = (inp[3]) ? 4'b1101 : 4'b1111;
												assign node26310 = (inp[3]) ? node26328 : node26311;
													assign node26311 = (inp[2]) ? node26321 : node26312;
														assign node26312 = (inp[5]) ? 4'b1011 : node26313;
															assign node26313 = (inp[0]) ? node26317 : node26314;
																assign node26314 = (inp[15]) ? 4'b1001 : 4'b1011;
																assign node26317 = (inp[15]) ? 4'b1011 : 4'b1001;
														assign node26321 = (inp[5]) ? node26323 : 4'b1011;
															assign node26323 = (inp[0]) ? 4'b1011 : node26324;
																assign node26324 = (inp[15]) ? 4'b1001 : 4'b1011;
													assign node26328 = (inp[15]) ? node26338 : node26329;
														assign node26329 = (inp[2]) ? node26333 : node26330;
															assign node26330 = (inp[5]) ? 4'b1011 : 4'b1001;
															assign node26333 = (inp[5]) ? node26335 : 4'b1011;
																assign node26335 = (inp[0]) ? 4'b1011 : 4'b1001;
														assign node26338 = (inp[2]) ? node26346 : node26339;
															assign node26339 = (inp[5]) ? node26343 : node26340;
																assign node26340 = (inp[0]) ? 4'b1011 : 4'b1001;
																assign node26343 = (inp[0]) ? 4'b1001 : 4'b1011;
															assign node26346 = (inp[5]) ? node26350 : node26347;
																assign node26347 = (inp[0]) ? 4'b1011 : 4'b1001;
																assign node26350 = (inp[0]) ? 4'b1001 : 4'b1011;
											assign node26353 = (inp[12]) ? node26369 : node26354;
												assign node26354 = (inp[5]) ? node26362 : node26355;
													assign node26355 = (inp[15]) ? node26359 : node26356;
														assign node26356 = (inp[0]) ? 4'b1001 : 4'b1011;
														assign node26359 = (inp[0]) ? 4'b1011 : 4'b1001;
													assign node26362 = (inp[3]) ? 4'b1011 : node26363;
														assign node26363 = (inp[0]) ? node26365 : 4'b1011;
															assign node26365 = (inp[15]) ? 4'b1011 : 4'b1001;
												assign node26369 = (inp[2]) ? node26383 : node26370;
													assign node26370 = (inp[15]) ? node26376 : node26371;
														assign node26371 = (inp[0]) ? node26373 : 4'b1011;
															assign node26373 = (inp[3]) ? 4'b1011 : 4'b1001;
														assign node26376 = (inp[0]) ? node26378 : 4'b1001;
															assign node26378 = (inp[3]) ? node26380 : 4'b1011;
																assign node26380 = (inp[5]) ? 4'b1001 : 4'b1011;
													assign node26383 = (inp[3]) ? node26391 : node26384;
														assign node26384 = (inp[15]) ? node26388 : node26385;
															assign node26385 = (inp[0]) ? 4'b1001 : 4'b1011;
															assign node26388 = (inp[0]) ? 4'b1011 : 4'b1001;
														assign node26391 = (inp[15]) ? node26393 : 4'b1001;
															assign node26393 = (inp[5]) ? node26395 : 4'b1001;
																assign node26395 = (inp[0]) ? 4'b1001 : 4'b1011;
										assign node26398 = (inp[10]) ? node26462 : node26399;
											assign node26399 = (inp[12]) ? node26417 : node26400;
												assign node26400 = (inp[5]) ? node26406 : node26401;
													assign node26401 = (inp[0]) ? node26403 : 4'b1001;
														assign node26403 = (inp[15]) ? 4'b1011 : 4'b1001;
													assign node26406 = (inp[2]) ? node26408 : 4'b1011;
														assign node26408 = (inp[15]) ? node26410 : 4'b1011;
															assign node26410 = (inp[0]) ? node26414 : node26411;
																assign node26411 = (inp[3]) ? 4'b1011 : 4'b1001;
																assign node26414 = (inp[3]) ? 4'b1001 : 4'b1011;
												assign node26417 = (inp[5]) ? node26439 : node26418;
													assign node26418 = (inp[15]) ? node26426 : node26419;
														assign node26419 = (inp[2]) ? 4'b1101 : node26420;
															assign node26420 = (inp[3]) ? node26422 : 4'b1101;
																assign node26422 = (inp[0]) ? 4'b1111 : 4'b1101;
														assign node26426 = (inp[2]) ? node26434 : node26427;
															assign node26427 = (inp[0]) ? node26431 : node26428;
																assign node26428 = (inp[3]) ? 4'b1111 : 4'b1101;
																assign node26431 = (inp[3]) ? 4'b1101 : 4'b1111;
															assign node26434 = (inp[3]) ? 4'b1111 : node26435;
																assign node26435 = (inp[0]) ? 4'b1111 : 4'b1101;
													assign node26439 = (inp[3]) ? node26447 : node26440;
														assign node26440 = (inp[15]) ? node26444 : node26441;
															assign node26441 = (inp[0]) ? 4'b1111 : 4'b1101;
															assign node26444 = (inp[0]) ? 4'b1101 : 4'b1111;
														assign node26447 = (inp[2]) ? node26455 : node26448;
															assign node26448 = (inp[15]) ? node26452 : node26449;
																assign node26449 = (inp[0]) ? 4'b1111 : 4'b1101;
																assign node26452 = (inp[0]) ? 4'b1101 : 4'b1111;
															assign node26455 = (inp[0]) ? node26459 : node26456;
																assign node26456 = (inp[15]) ? 4'b1111 : 4'b1101;
																assign node26459 = (inp[15]) ? 4'b1101 : 4'b1111;
											assign node26462 = (inp[0]) ? node26474 : node26463;
												assign node26463 = (inp[15]) ? node26469 : node26464;
													assign node26464 = (inp[5]) ? 4'b1101 : node26465;
														assign node26465 = (inp[3]) ? 4'b1101 : 4'b1111;
													assign node26469 = (inp[3]) ? 4'b1111 : node26470;
														assign node26470 = (inp[5]) ? 4'b1111 : 4'b1101;
												assign node26474 = (inp[15]) ? node26480 : node26475;
													assign node26475 = (inp[5]) ? 4'b1111 : node26476;
														assign node26476 = (inp[3]) ? 4'b1111 : 4'b1101;
													assign node26480 = (inp[3]) ? 4'b1101 : node26481;
														assign node26481 = (inp[5]) ? 4'b1101 : 4'b1111;
									assign node26485 = (inp[4]) ? node26565 : node26486;
										assign node26486 = (inp[12]) ? node26532 : node26487;
											assign node26487 = (inp[10]) ? node26511 : node26488;
												assign node26488 = (inp[15]) ? node26500 : node26489;
													assign node26489 = (inp[0]) ? node26495 : node26490;
														assign node26490 = (inp[5]) ? node26492 : 4'b1011;
															assign node26492 = (inp[3]) ? 4'b1001 : 4'b1011;
														assign node26495 = (inp[5]) ? node26497 : 4'b1001;
															assign node26497 = (inp[3]) ? 4'b1011 : 4'b1001;
													assign node26500 = (inp[0]) ? node26506 : node26501;
														assign node26501 = (inp[5]) ? node26503 : 4'b1001;
															assign node26503 = (inp[3]) ? 4'b1011 : 4'b1001;
														assign node26506 = (inp[5]) ? node26508 : 4'b1011;
															assign node26508 = (inp[3]) ? 4'b1001 : 4'b1011;
												assign node26511 = (inp[0]) ? node26523 : node26512;
													assign node26512 = (inp[15]) ? node26518 : node26513;
														assign node26513 = (inp[5]) ? 4'b1101 : node26514;
															assign node26514 = (inp[3]) ? 4'b1101 : 4'b1111;
														assign node26518 = (inp[3]) ? 4'b1111 : node26519;
															assign node26519 = (inp[5]) ? 4'b1111 : 4'b1101;
													assign node26523 = (inp[3]) ? 4'b1111 : node26524;
														assign node26524 = (inp[5]) ? node26528 : node26525;
															assign node26525 = (inp[15]) ? 4'b1111 : 4'b1101;
															assign node26528 = (inp[15]) ? 4'b1101 : 4'b1111;
											assign node26532 = (inp[3]) ? node26558 : node26533;
												assign node26533 = (inp[5]) ? node26543 : node26534;
													assign node26534 = (inp[10]) ? node26536 : 4'b1111;
														assign node26536 = (inp[2]) ? 4'b1111 : node26537;
															assign node26537 = (inp[0]) ? 4'b1101 : node26538;
																assign node26538 = (inp[15]) ? 4'b1101 : 4'b1111;
													assign node26543 = (inp[10]) ? node26551 : node26544;
														assign node26544 = (inp[15]) ? node26548 : node26545;
															assign node26545 = (inp[0]) ? 4'b1111 : 4'b1101;
															assign node26548 = (inp[0]) ? 4'b1101 : 4'b1111;
														assign node26551 = (inp[15]) ? node26555 : node26552;
															assign node26552 = (inp[0]) ? 4'b1111 : 4'b1101;
															assign node26555 = (inp[0]) ? 4'b1101 : 4'b1111;
												assign node26558 = (inp[15]) ? node26562 : node26559;
													assign node26559 = (inp[0]) ? 4'b1111 : 4'b1101;
													assign node26562 = (inp[0]) ? 4'b1101 : 4'b1111;
										assign node26565 = (inp[10]) ? node26629 : node26566;
											assign node26566 = (inp[12]) ? node26608 : node26567;
												assign node26567 = (inp[2]) ? node26587 : node26568;
													assign node26568 = (inp[5]) ? node26582 : node26569;
														assign node26569 = (inp[0]) ? node26575 : node26570;
															assign node26570 = (inp[3]) ? node26572 : 4'b1111;
																assign node26572 = (inp[15]) ? 4'b1111 : 4'b1101;
															assign node26575 = (inp[15]) ? node26579 : node26576;
																assign node26576 = (inp[3]) ? 4'b1111 : 4'b1101;
																assign node26579 = (inp[3]) ? 4'b1101 : 4'b1111;
														assign node26582 = (inp[0]) ? 4'b1111 : node26583;
															assign node26583 = (inp[15]) ? 4'b1111 : 4'b1101;
													assign node26587 = (inp[5]) ? node26601 : node26588;
														assign node26588 = (inp[15]) ? node26594 : node26589;
															assign node26589 = (inp[3]) ? 4'b1111 : node26590;
																assign node26590 = (inp[0]) ? 4'b1101 : 4'b1111;
															assign node26594 = (inp[0]) ? node26598 : node26595;
																assign node26595 = (inp[3]) ? 4'b1111 : 4'b1101;
																assign node26598 = (inp[3]) ? 4'b1101 : 4'b1111;
														assign node26601 = (inp[15]) ? node26605 : node26602;
															assign node26602 = (inp[0]) ? 4'b1111 : 4'b1101;
															assign node26605 = (inp[0]) ? 4'b1101 : 4'b1111;
												assign node26608 = (inp[0]) ? node26620 : node26609;
													assign node26609 = (inp[15]) ? node26615 : node26610;
														assign node26610 = (inp[5]) ? 4'b1001 : node26611;
															assign node26611 = (inp[3]) ? 4'b1001 : 4'b1011;
														assign node26615 = (inp[3]) ? 4'b1011 : node26616;
															assign node26616 = (inp[5]) ? 4'b1011 : 4'b1001;
													assign node26620 = (inp[15]) ? node26626 : node26621;
														assign node26621 = (inp[5]) ? 4'b1011 : node26622;
															assign node26622 = (inp[2]) ? 4'b1001 : 4'b1011;
														assign node26626 = (inp[5]) ? 4'b1001 : 4'b1011;
											assign node26629 = (inp[15]) ? node26637 : node26630;
												assign node26630 = (inp[0]) ? 4'b1011 : node26631;
													assign node26631 = (inp[3]) ? 4'b1001 : node26632;
														assign node26632 = (inp[5]) ? 4'b1001 : 4'b1011;
												assign node26637 = (inp[0]) ? node26643 : node26638;
													assign node26638 = (inp[5]) ? 4'b1011 : node26639;
														assign node26639 = (inp[3]) ? 4'b1011 : 4'b1001;
													assign node26643 = (inp[5]) ? 4'b1001 : node26644;
														assign node26644 = (inp[3]) ? 4'b1001 : 4'b1011;
						assign node26648 = (inp[7]) ? node27750 : node26649;
							assign node26649 = (inp[14]) ? node27157 : node26650;
								assign node26650 = (inp[2]) ? node26908 : node26651;
									assign node26651 = (inp[4]) ? node26785 : node26652;
										assign node26652 = (inp[9]) ? node26712 : node26653;
											assign node26653 = (inp[12]) ? node26683 : node26654;
												assign node26654 = (inp[3]) ? node26670 : node26655;
													assign node26655 = (inp[10]) ? node26663 : node26656;
														assign node26656 = (inp[5]) ? 4'b0100 : node26657;
															assign node26657 = (inp[15]) ? 4'b0100 : node26658;
																assign node26658 = (inp[0]) ? 4'b0100 : 4'b0110;
														assign node26663 = (inp[15]) ? node26667 : node26664;
															assign node26664 = (inp[0]) ? 4'b0100 : 4'b0110;
															assign node26667 = (inp[0]) ? 4'b0110 : 4'b0100;
													assign node26670 = (inp[5]) ? node26672 : 4'b0110;
														assign node26672 = (inp[10]) ? node26678 : node26673;
															assign node26673 = (inp[15]) ? node26675 : 4'b0110;
																assign node26675 = (inp[0]) ? 4'b0100 : 4'b0110;
															assign node26678 = (inp[0]) ? 4'b0100 : node26679;
																assign node26679 = (inp[15]) ? 4'b0110 : 4'b0100;
												assign node26683 = (inp[10]) ? node26693 : node26684;
													assign node26684 = (inp[5]) ? 4'b0100 : node26685;
														assign node26685 = (inp[15]) ? node26689 : node26686;
															assign node26686 = (inp[0]) ? 4'b0100 : 4'b0110;
															assign node26689 = (inp[0]) ? 4'b0110 : 4'b0100;
													assign node26693 = (inp[15]) ? node26703 : node26694;
														assign node26694 = (inp[0]) ? node26698 : node26695;
															assign node26695 = (inp[5]) ? 4'b0000 : 4'b0010;
															assign node26698 = (inp[3]) ? node26700 : 4'b0000;
																assign node26700 = (inp[5]) ? 4'b0010 : 4'b0000;
														assign node26703 = (inp[0]) ? node26709 : node26704;
															assign node26704 = (inp[3]) ? node26706 : 4'b0000;
																assign node26706 = (inp[5]) ? 4'b0010 : 4'b0000;
															assign node26709 = (inp[3]) ? 4'b0000 : 4'b0010;
											assign node26712 = (inp[10]) ? node26752 : node26713;
												assign node26713 = (inp[12]) ? node26735 : node26714;
													assign node26714 = (inp[3]) ? node26728 : node26715;
														assign node26715 = (inp[5]) ? node26721 : node26716;
															assign node26716 = (inp[0]) ? 4'b0010 : node26717;
																assign node26717 = (inp[15]) ? 4'b0000 : 4'b0010;
															assign node26721 = (inp[15]) ? node26725 : node26722;
																assign node26722 = (inp[0]) ? 4'b0000 : 4'b0010;
																assign node26725 = (inp[0]) ? 4'b0010 : 4'b0000;
														assign node26728 = (inp[0]) ? 4'b0010 : node26729;
															assign node26729 = (inp[5]) ? node26731 : 4'b0010;
																assign node26731 = (inp[15]) ? 4'b0010 : 4'b0000;
													assign node26735 = (inp[0]) ? node26743 : node26736;
														assign node26736 = (inp[15]) ? node26738 : 4'b0010;
															assign node26738 = (inp[5]) ? node26740 : 4'b0000;
																assign node26740 = (inp[3]) ? 4'b0010 : 4'b0000;
														assign node26743 = (inp[15]) ? node26749 : node26744;
															assign node26744 = (inp[3]) ? node26746 : 4'b0000;
																assign node26746 = (inp[5]) ? 4'b0010 : 4'b0000;
															assign node26749 = (inp[5]) ? 4'b0000 : 4'b0010;
												assign node26752 = (inp[12]) ? node26762 : node26753;
													assign node26753 = (inp[5]) ? 4'b0010 : node26754;
														assign node26754 = (inp[0]) ? node26758 : node26755;
															assign node26755 = (inp[15]) ? 4'b0000 : 4'b0010;
															assign node26758 = (inp[15]) ? 4'b0010 : 4'b0000;
													assign node26762 = (inp[3]) ? node26776 : node26763;
														assign node26763 = (inp[5]) ? node26769 : node26764;
															assign node26764 = (inp[0]) ? node26766 : 4'b0110;
																assign node26766 = (inp[15]) ? 4'b0110 : 4'b0100;
															assign node26769 = (inp[15]) ? node26773 : node26770;
																assign node26770 = (inp[0]) ? 4'b0110 : 4'b0100;
																assign node26773 = (inp[0]) ? 4'b0100 : 4'b0110;
														assign node26776 = (inp[5]) ? node26778 : 4'b0100;
															assign node26778 = (inp[15]) ? node26782 : node26779;
																assign node26779 = (inp[0]) ? 4'b0110 : 4'b0100;
																assign node26782 = (inp[0]) ? 4'b0100 : 4'b0110;
										assign node26785 = (inp[9]) ? node26839 : node26786;
											assign node26786 = (inp[12]) ? node26808 : node26787;
												assign node26787 = (inp[0]) ? node26797 : node26788;
													assign node26788 = (inp[15]) ? node26792 : node26789;
														assign node26789 = (inp[3]) ? 4'b0000 : 4'b0010;
														assign node26792 = (inp[5]) ? node26794 : 4'b0000;
															assign node26794 = (inp[3]) ? 4'b0010 : 4'b0000;
													assign node26797 = (inp[15]) ? node26803 : node26798;
														assign node26798 = (inp[5]) ? node26800 : 4'b0000;
															assign node26800 = (inp[3]) ? 4'b0010 : 4'b0000;
														assign node26803 = (inp[5]) ? node26805 : 4'b0010;
															assign node26805 = (inp[3]) ? 4'b0000 : 4'b0010;
												assign node26808 = (inp[10]) ? node26818 : node26809;
													assign node26809 = (inp[15]) ? node26813 : node26810;
														assign node26810 = (inp[0]) ? 4'b0000 : 4'b0010;
														assign node26813 = (inp[0]) ? 4'b0010 : node26814;
															assign node26814 = (inp[5]) ? 4'b0010 : 4'b0000;
													assign node26818 = (inp[15]) ? node26828 : node26819;
														assign node26819 = (inp[0]) ? node26823 : node26820;
															assign node26820 = (inp[5]) ? 4'b0100 : 4'b0110;
															assign node26823 = (inp[3]) ? 4'b0110 : node26824;
																assign node26824 = (inp[5]) ? 4'b0110 : 4'b0100;
														assign node26828 = (inp[0]) ? node26834 : node26829;
															assign node26829 = (inp[3]) ? 4'b0110 : node26830;
																assign node26830 = (inp[5]) ? 4'b0110 : 4'b0100;
															assign node26834 = (inp[5]) ? 4'b0100 : node26835;
																assign node26835 = (inp[3]) ? 4'b0100 : 4'b0110;
											assign node26839 = (inp[12]) ? node26875 : node26840;
												assign node26840 = (inp[3]) ? node26860 : node26841;
													assign node26841 = (inp[15]) ? node26849 : node26842;
														assign node26842 = (inp[0]) ? node26846 : node26843;
															assign node26843 = (inp[5]) ? 4'b0100 : 4'b0110;
															assign node26846 = (inp[5]) ? 4'b0110 : 4'b0100;
														assign node26849 = (inp[10]) ? node26855 : node26850;
															assign node26850 = (inp[0]) ? node26852 : 4'b0100;
																assign node26852 = (inp[5]) ? 4'b0100 : 4'b0110;
															assign node26855 = (inp[5]) ? node26857 : 4'b0110;
																assign node26857 = (inp[0]) ? 4'b0100 : 4'b0110;
													assign node26860 = (inp[5]) ? node26868 : node26861;
														assign node26861 = (inp[0]) ? node26865 : node26862;
															assign node26862 = (inp[15]) ? 4'b0110 : 4'b0100;
															assign node26865 = (inp[15]) ? 4'b0100 : 4'b0110;
														assign node26868 = (inp[0]) ? node26872 : node26869;
															assign node26869 = (inp[15]) ? 4'b0110 : 4'b0100;
															assign node26872 = (inp[15]) ? 4'b0100 : 4'b0110;
												assign node26875 = (inp[10]) ? node26885 : node26876;
													assign node26876 = (inp[15]) ? node26878 : 4'b0110;
														assign node26878 = (inp[0]) ? 4'b0100 : node26879;
															assign node26879 = (inp[3]) ? 4'b0110 : node26880;
																assign node26880 = (inp[5]) ? 4'b0110 : 4'b0100;
													assign node26885 = (inp[3]) ? node26901 : node26886;
														assign node26886 = (inp[5]) ? node26894 : node26887;
															assign node26887 = (inp[0]) ? node26891 : node26888;
																assign node26888 = (inp[15]) ? 4'b0000 : 4'b0010;
																assign node26891 = (inp[15]) ? 4'b0010 : 4'b0000;
															assign node26894 = (inp[15]) ? node26898 : node26895;
																assign node26895 = (inp[0]) ? 4'b0010 : 4'b0000;
																assign node26898 = (inp[0]) ? 4'b0000 : 4'b0010;
														assign node26901 = (inp[5]) ? node26903 : 4'b0000;
															assign node26903 = (inp[0]) ? 4'b0000 : node26904;
																assign node26904 = (inp[15]) ? 4'b0010 : 4'b0000;
									assign node26908 = (inp[9]) ? node27026 : node26909;
										assign node26909 = (inp[4]) ? node26975 : node26910;
											assign node26910 = (inp[10]) ? node26952 : node26911;
												assign node26911 = (inp[12]) ? node26931 : node26912;
													assign node26912 = (inp[3]) ? node26920 : node26913;
														assign node26913 = (inp[15]) ? node26917 : node26914;
															assign node26914 = (inp[0]) ? 4'b1101 : 4'b1111;
															assign node26917 = (inp[0]) ? 4'b1111 : 4'b1101;
														assign node26920 = (inp[0]) ? node26926 : node26921;
															assign node26921 = (inp[5]) ? node26923 : 4'b1111;
																assign node26923 = (inp[15]) ? 4'b1111 : 4'b1101;
															assign node26926 = (inp[5]) ? node26928 : 4'b1101;
																assign node26928 = (inp[15]) ? 4'b1101 : 4'b1111;
													assign node26931 = (inp[5]) ? node26939 : node26932;
														assign node26932 = (inp[0]) ? node26936 : node26933;
															assign node26933 = (inp[15]) ? 4'b1001 : 4'b1011;
															assign node26936 = (inp[15]) ? 4'b1011 : 4'b1001;
														assign node26939 = (inp[0]) ? node26947 : node26940;
															assign node26940 = (inp[15]) ? node26944 : node26941;
																assign node26941 = (inp[3]) ? 4'b1001 : 4'b1011;
																assign node26944 = (inp[3]) ? 4'b1011 : 4'b1001;
															assign node26947 = (inp[3]) ? node26949 : 4'b1001;
																assign node26949 = (inp[15]) ? 4'b1001 : 4'b1011;
												assign node26952 = (inp[15]) ? node26964 : node26953;
													assign node26953 = (inp[0]) ? node26959 : node26954;
														assign node26954 = (inp[3]) ? node26956 : 4'b1011;
															assign node26956 = (inp[5]) ? 4'b1001 : 4'b1011;
														assign node26959 = (inp[3]) ? node26961 : 4'b1001;
															assign node26961 = (inp[5]) ? 4'b1011 : 4'b1001;
													assign node26964 = (inp[0]) ? node26970 : node26965;
														assign node26965 = (inp[5]) ? node26967 : 4'b1001;
															assign node26967 = (inp[3]) ? 4'b1011 : 4'b1001;
														assign node26970 = (inp[5]) ? node26972 : 4'b1011;
															assign node26972 = (inp[3]) ? 4'b1001 : 4'b1011;
											assign node26975 = (inp[10]) ? node27005 : node26976;
												assign node26976 = (inp[12]) ? node26990 : node26977;
													assign node26977 = (inp[3]) ? node26985 : node26978;
														assign node26978 = (inp[0]) ? node26982 : node26979;
															assign node26979 = (inp[15]) ? 4'b1001 : 4'b1011;
															assign node26982 = (inp[15]) ? 4'b1011 : 4'b1001;
														assign node26985 = (inp[5]) ? node26987 : 4'b1001;
															assign node26987 = (inp[15]) ? 4'b1001 : 4'b1011;
													assign node26990 = (inp[15]) ? node26998 : node26991;
														assign node26991 = (inp[5]) ? node26995 : node26992;
															assign node26992 = (inp[0]) ? 4'b1101 : 4'b1111;
															assign node26995 = (inp[0]) ? 4'b1111 : 4'b1101;
														assign node26998 = (inp[0]) ? node27002 : node26999;
															assign node26999 = (inp[3]) ? 4'b1111 : 4'b1101;
															assign node27002 = (inp[3]) ? 4'b1101 : 4'b1111;
												assign node27005 = (inp[15]) ? node27017 : node27006;
													assign node27006 = (inp[0]) ? node27012 : node27007;
														assign node27007 = (inp[5]) ? 4'b1101 : node27008;
															assign node27008 = (inp[3]) ? 4'b1101 : 4'b1111;
														assign node27012 = (inp[3]) ? 4'b1111 : node27013;
															assign node27013 = (inp[5]) ? 4'b1111 : 4'b1101;
													assign node27017 = (inp[0]) ? node27023 : node27018;
														assign node27018 = (inp[5]) ? 4'b1111 : node27019;
															assign node27019 = (inp[3]) ? 4'b1111 : 4'b1101;
														assign node27023 = (inp[3]) ? 4'b1101 : 4'b1111;
										assign node27026 = (inp[4]) ? node27086 : node27027;
											assign node27027 = (inp[12]) ? node27063 : node27028;
												assign node27028 = (inp[10]) ? node27048 : node27029;
													assign node27029 = (inp[15]) ? node27039 : node27030;
														assign node27030 = (inp[0]) ? node27034 : node27031;
															assign node27031 = (inp[5]) ? 4'b1001 : 4'b1011;
															assign node27034 = (inp[5]) ? node27036 : 4'b1001;
																assign node27036 = (inp[3]) ? 4'b1011 : 4'b1001;
														assign node27039 = (inp[5]) ? node27041 : 4'b1011;
															assign node27041 = (inp[3]) ? node27045 : node27042;
																assign node27042 = (inp[0]) ? 4'b1011 : 4'b1001;
																assign node27045 = (inp[0]) ? 4'b1001 : 4'b1011;
													assign node27048 = (inp[3]) ? node27058 : node27049;
														assign node27049 = (inp[15]) ? node27051 : 4'b1111;
															assign node27051 = (inp[0]) ? node27055 : node27052;
																assign node27052 = (inp[5]) ? 4'b1111 : 4'b1101;
																assign node27055 = (inp[5]) ? 4'b1101 : 4'b1111;
														assign node27058 = (inp[5]) ? 4'b1101 : node27059;
															assign node27059 = (inp[15]) ? 4'b1111 : 4'b1101;
												assign node27063 = (inp[3]) ? node27079 : node27064;
													assign node27064 = (inp[10]) ? 4'b1101 : node27065;
														assign node27065 = (inp[0]) ? node27073 : node27066;
															assign node27066 = (inp[15]) ? node27070 : node27067;
																assign node27067 = (inp[5]) ? 4'b1101 : 4'b1111;
																assign node27070 = (inp[5]) ? 4'b1111 : 4'b1101;
															assign node27073 = (inp[5]) ? node27075 : 4'b1101;
																assign node27075 = (inp[15]) ? 4'b1101 : 4'b1111;
													assign node27079 = (inp[0]) ? node27083 : node27080;
														assign node27080 = (inp[15]) ? 4'b1111 : 4'b1101;
														assign node27083 = (inp[15]) ? 4'b1101 : 4'b1111;
											assign node27086 = (inp[12]) ? node27128 : node27087;
												assign node27087 = (inp[10]) ? node27107 : node27088;
													assign node27088 = (inp[3]) ? node27100 : node27089;
														assign node27089 = (inp[0]) ? node27095 : node27090;
															assign node27090 = (inp[15]) ? 4'b1111 : node27091;
																assign node27091 = (inp[5]) ? 4'b1101 : 4'b1111;
															assign node27095 = (inp[5]) ? 4'b1101 : node27096;
																assign node27096 = (inp[15]) ? 4'b1111 : 4'b1101;
														assign node27100 = (inp[15]) ? node27104 : node27101;
															assign node27101 = (inp[0]) ? 4'b1111 : 4'b1101;
															assign node27104 = (inp[0]) ? 4'b1101 : 4'b1111;
													assign node27107 = (inp[5]) ? node27123 : node27108;
														assign node27108 = (inp[3]) ? node27116 : node27109;
															assign node27109 = (inp[15]) ? node27113 : node27110;
																assign node27110 = (inp[0]) ? 4'b1001 : 4'b1011;
																assign node27113 = (inp[0]) ? 4'b1011 : 4'b1001;
															assign node27116 = (inp[15]) ? node27120 : node27117;
																assign node27117 = (inp[0]) ? 4'b1011 : 4'b1001;
																assign node27120 = (inp[0]) ? 4'b1001 : 4'b1011;
														assign node27123 = (inp[0]) ? 4'b1001 : node27124;
															assign node27124 = (inp[15]) ? 4'b1011 : 4'b1001;
												assign node27128 = (inp[5]) ? node27150 : node27129;
													assign node27129 = (inp[0]) ? node27143 : node27130;
														assign node27130 = (inp[10]) ? node27138 : node27131;
															assign node27131 = (inp[15]) ? node27135 : node27132;
																assign node27132 = (inp[3]) ? 4'b1001 : 4'b1011;
																assign node27135 = (inp[3]) ? 4'b1011 : 4'b1001;
															assign node27138 = (inp[15]) ? node27140 : 4'b1001;
																assign node27140 = (inp[3]) ? 4'b1011 : 4'b1001;
														assign node27143 = (inp[3]) ? node27147 : node27144;
															assign node27144 = (inp[15]) ? 4'b1011 : 4'b1001;
															assign node27147 = (inp[15]) ? 4'b1001 : 4'b1011;
													assign node27150 = (inp[15]) ? node27154 : node27151;
														assign node27151 = (inp[0]) ? 4'b1011 : 4'b1001;
														assign node27154 = (inp[0]) ? 4'b1001 : 4'b1011;
								assign node27157 = (inp[2]) ? node27427 : node27158;
									assign node27158 = (inp[9]) ? node27290 : node27159;
										assign node27159 = (inp[4]) ? node27225 : node27160;
											assign node27160 = (inp[10]) ? node27194 : node27161;
												assign node27161 = (inp[12]) ? node27183 : node27162;
													assign node27162 = (inp[5]) ? node27176 : node27163;
														assign node27163 = (inp[3]) ? node27171 : node27164;
															assign node27164 = (inp[15]) ? node27168 : node27165;
																assign node27165 = (inp[0]) ? 4'b1101 : 4'b1111;
																assign node27168 = (inp[0]) ? 4'b1111 : 4'b1101;
															assign node27171 = (inp[15]) ? 4'b1101 : node27172;
																assign node27172 = (inp[0]) ? 4'b1101 : 4'b1111;
														assign node27176 = (inp[15]) ? 4'b1111 : node27177;
															assign node27177 = (inp[3]) ? 4'b1111 : node27178;
																assign node27178 = (inp[0]) ? 4'b1101 : 4'b1111;
													assign node27183 = (inp[0]) ? node27191 : node27184;
														assign node27184 = (inp[3]) ? node27186 : 4'b1001;
															assign node27186 = (inp[15]) ? node27188 : 4'b1011;
																assign node27188 = (inp[5]) ? 4'b1011 : 4'b1001;
														assign node27191 = (inp[15]) ? 4'b1011 : 4'b1001;
												assign node27194 = (inp[3]) ? node27210 : node27195;
													assign node27195 = (inp[12]) ? node27203 : node27196;
														assign node27196 = (inp[15]) ? node27200 : node27197;
															assign node27197 = (inp[0]) ? 4'b1001 : 4'b1011;
															assign node27200 = (inp[0]) ? 4'b1011 : 4'b1001;
														assign node27203 = (inp[0]) ? node27207 : node27204;
															assign node27204 = (inp[15]) ? 4'b1001 : 4'b1011;
															assign node27207 = (inp[15]) ? 4'b1011 : 4'b1001;
													assign node27210 = (inp[5]) ? node27220 : node27211;
														assign node27211 = (inp[12]) ? node27217 : node27212;
															assign node27212 = (inp[0]) ? 4'b1011 : node27213;
																assign node27213 = (inp[15]) ? 4'b1001 : 4'b1011;
															assign node27217 = (inp[0]) ? 4'b1001 : 4'b1011;
														assign node27220 = (inp[15]) ? 4'b1011 : node27221;
															assign node27221 = (inp[0]) ? 4'b1011 : 4'b1001;
											assign node27225 = (inp[12]) ? node27263 : node27226;
												assign node27226 = (inp[10]) ? node27246 : node27227;
													assign node27227 = (inp[5]) ? node27233 : node27228;
														assign node27228 = (inp[15]) ? 4'b1011 : node27229;
															assign node27229 = (inp[0]) ? 4'b1001 : 4'b1011;
														assign node27233 = (inp[3]) ? node27239 : node27234;
															assign node27234 = (inp[0]) ? 4'b1001 : node27235;
																assign node27235 = (inp[15]) ? 4'b1001 : 4'b1011;
															assign node27239 = (inp[0]) ? node27243 : node27240;
																assign node27240 = (inp[15]) ? 4'b1011 : 4'b1001;
																assign node27243 = (inp[15]) ? 4'b1001 : 4'b1011;
													assign node27246 = (inp[15]) ? node27256 : node27247;
														assign node27247 = (inp[0]) ? node27251 : node27248;
															assign node27248 = (inp[5]) ? 4'b1101 : 4'b1111;
															assign node27251 = (inp[5]) ? 4'b1111 : node27252;
																assign node27252 = (inp[3]) ? 4'b1111 : 4'b1101;
														assign node27256 = (inp[3]) ? node27260 : node27257;
															assign node27257 = (inp[0]) ? 4'b1111 : 4'b1101;
															assign node27260 = (inp[0]) ? 4'b1101 : 4'b1111;
												assign node27263 = (inp[10]) ? node27281 : node27264;
													assign node27264 = (inp[15]) ? node27276 : node27265;
														assign node27265 = (inp[0]) ? node27271 : node27266;
															assign node27266 = (inp[3]) ? 4'b1101 : node27267;
																assign node27267 = (inp[5]) ? 4'b1101 : 4'b1111;
															assign node27271 = (inp[3]) ? 4'b1111 : node27272;
																assign node27272 = (inp[5]) ? 4'b1111 : 4'b1101;
														assign node27276 = (inp[0]) ? 4'b1101 : node27277;
															assign node27277 = (inp[3]) ? 4'b1111 : 4'b1101;
													assign node27281 = (inp[15]) ? node27285 : node27282;
														assign node27282 = (inp[5]) ? 4'b1111 : 4'b1101;
														assign node27285 = (inp[0]) ? node27287 : 4'b1111;
															assign node27287 = (inp[3]) ? 4'b1101 : 4'b1111;
										assign node27290 = (inp[4]) ? node27370 : node27291;
											assign node27291 = (inp[12]) ? node27331 : node27292;
												assign node27292 = (inp[10]) ? node27314 : node27293;
													assign node27293 = (inp[5]) ? node27301 : node27294;
														assign node27294 = (inp[0]) ? node27298 : node27295;
															assign node27295 = (inp[15]) ? 4'b1001 : 4'b1011;
															assign node27298 = (inp[15]) ? 4'b1011 : 4'b1001;
														assign node27301 = (inp[15]) ? node27309 : node27302;
															assign node27302 = (inp[0]) ? node27306 : node27303;
																assign node27303 = (inp[3]) ? 4'b1001 : 4'b1011;
																assign node27306 = (inp[3]) ? 4'b1011 : 4'b1001;
															assign node27309 = (inp[0]) ? node27311 : 4'b1001;
																assign node27311 = (inp[3]) ? 4'b1001 : 4'b1011;
													assign node27314 = (inp[5]) ? node27326 : node27315;
														assign node27315 = (inp[15]) ? node27321 : node27316;
															assign node27316 = (inp[3]) ? node27318 : 4'b1111;
																assign node27318 = (inp[0]) ? 4'b1111 : 4'b1101;
															assign node27321 = (inp[0]) ? 4'b1101 : node27322;
																assign node27322 = (inp[3]) ? 4'b1111 : 4'b1101;
														assign node27326 = (inp[0]) ? 4'b1101 : node27327;
															assign node27327 = (inp[15]) ? 4'b1111 : 4'b1101;
												assign node27331 = (inp[3]) ? node27357 : node27332;
													assign node27332 = (inp[10]) ? node27342 : node27333;
														assign node27333 = (inp[15]) ? node27335 : 4'b1111;
															assign node27335 = (inp[0]) ? node27339 : node27336;
																assign node27336 = (inp[5]) ? 4'b1111 : 4'b1101;
																assign node27339 = (inp[5]) ? 4'b1101 : 4'b1111;
														assign node27342 = (inp[5]) ? node27350 : node27343;
															assign node27343 = (inp[15]) ? node27347 : node27344;
																assign node27344 = (inp[0]) ? 4'b1101 : 4'b1111;
																assign node27347 = (inp[0]) ? 4'b1111 : 4'b1101;
															assign node27350 = (inp[15]) ? node27354 : node27351;
																assign node27351 = (inp[0]) ? 4'b1111 : 4'b1101;
																assign node27354 = (inp[0]) ? 4'b1101 : 4'b1111;
													assign node27357 = (inp[5]) ? node27365 : node27358;
														assign node27358 = (inp[15]) ? node27362 : node27359;
															assign node27359 = (inp[0]) ? 4'b1111 : 4'b1101;
															assign node27362 = (inp[0]) ? 4'b1101 : 4'b1111;
														assign node27365 = (inp[0]) ? 4'b1101 : node27366;
															assign node27366 = (inp[15]) ? 4'b1111 : 4'b1101;
											assign node27370 = (inp[12]) ? node27406 : node27371;
												assign node27371 = (inp[10]) ? node27385 : node27372;
													assign node27372 = (inp[0]) ? node27376 : node27373;
														assign node27373 = (inp[15]) ? 4'b1111 : 4'b1101;
														assign node27376 = (inp[15]) ? node27380 : node27377;
															assign node27377 = (inp[5]) ? 4'b1111 : 4'b1101;
															assign node27380 = (inp[5]) ? 4'b1101 : node27381;
																assign node27381 = (inp[3]) ? 4'b1101 : 4'b1111;
													assign node27385 = (inp[3]) ? node27399 : node27386;
														assign node27386 = (inp[0]) ? node27392 : node27387;
															assign node27387 = (inp[5]) ? node27389 : 4'b1011;
																assign node27389 = (inp[15]) ? 4'b1011 : 4'b1001;
															assign node27392 = (inp[5]) ? node27396 : node27393;
																assign node27393 = (inp[15]) ? 4'b1011 : 4'b1001;
																assign node27396 = (inp[15]) ? 4'b1001 : 4'b1011;
														assign node27399 = (inp[0]) ? node27403 : node27400;
															assign node27400 = (inp[15]) ? 4'b1011 : 4'b1001;
															assign node27403 = (inp[15]) ? 4'b1001 : 4'b1011;
												assign node27406 = (inp[15]) ? node27418 : node27407;
													assign node27407 = (inp[0]) ? node27413 : node27408;
														assign node27408 = (inp[5]) ? 4'b1001 : node27409;
															assign node27409 = (inp[3]) ? 4'b1001 : 4'b1011;
														assign node27413 = (inp[5]) ? 4'b1011 : node27414;
															assign node27414 = (inp[3]) ? 4'b1011 : 4'b1001;
													assign node27418 = (inp[0]) ? node27422 : node27419;
														assign node27419 = (inp[3]) ? 4'b1011 : 4'b1001;
														assign node27422 = (inp[5]) ? 4'b1001 : node27423;
															assign node27423 = (inp[3]) ? 4'b1001 : 4'b1011;
									assign node27427 = (inp[5]) ? node27581 : node27428;
										assign node27428 = (inp[12]) ? node27516 : node27429;
											assign node27429 = (inp[0]) ? node27479 : node27430;
												assign node27430 = (inp[15]) ? node27456 : node27431;
													assign node27431 = (inp[3]) ? node27441 : node27432;
														assign node27432 = (inp[4]) ? node27434 : 4'b1011;
															assign node27434 = (inp[9]) ? node27438 : node27435;
																assign node27435 = (inp[10]) ? 4'b1111 : 4'b1011;
																assign node27438 = (inp[10]) ? 4'b1011 : 4'b1111;
														assign node27441 = (inp[4]) ? node27449 : node27442;
															assign node27442 = (inp[10]) ? node27446 : node27443;
																assign node27443 = (inp[9]) ? 4'b1011 : 4'b1111;
																assign node27446 = (inp[9]) ? 4'b1101 : 4'b1011;
															assign node27449 = (inp[10]) ? node27453 : node27450;
																assign node27450 = (inp[9]) ? 4'b1101 : 4'b1011;
																assign node27453 = (inp[9]) ? 4'b1001 : 4'b1101;
													assign node27456 = (inp[3]) ? node27466 : node27457;
														assign node27457 = (inp[10]) ? 4'b1001 : node27458;
															assign node27458 = (inp[9]) ? node27462 : node27459;
																assign node27459 = (inp[4]) ? 4'b1001 : 4'b1101;
																assign node27462 = (inp[4]) ? 4'b1101 : 4'b1001;
														assign node27466 = (inp[9]) ? node27472 : node27467;
															assign node27467 = (inp[10]) ? node27469 : 4'b1001;
																assign node27469 = (inp[4]) ? 4'b1111 : 4'b1001;
															assign node27472 = (inp[10]) ? node27476 : node27473;
																assign node27473 = (inp[4]) ? 4'b1111 : 4'b1001;
																assign node27476 = (inp[4]) ? 4'b1011 : 4'b1111;
												assign node27479 = (inp[15]) ? node27503 : node27480;
													assign node27480 = (inp[3]) ? node27494 : node27481;
														assign node27481 = (inp[10]) ? node27489 : node27482;
															assign node27482 = (inp[4]) ? node27486 : node27483;
																assign node27483 = (inp[9]) ? 4'b1001 : 4'b1101;
																assign node27486 = (inp[9]) ? 4'b1101 : 4'b1001;
															assign node27489 = (inp[4]) ? 4'b1101 : node27490;
																assign node27490 = (inp[9]) ? 4'b1101 : 4'b1001;
														assign node27494 = (inp[9]) ? node27498 : node27495;
															assign node27495 = (inp[4]) ? 4'b1001 : 4'b1101;
															assign node27498 = (inp[10]) ? node27500 : 4'b1111;
																assign node27500 = (inp[4]) ? 4'b1011 : 4'b1111;
													assign node27503 = (inp[10]) ? node27509 : node27504;
														assign node27504 = (inp[9]) ? 4'b1011 : node27505;
															assign node27505 = (inp[4]) ? 4'b1011 : 4'b1111;
														assign node27509 = (inp[3]) ? 4'b1101 : node27510;
															assign node27510 = (inp[4]) ? node27512 : 4'b1111;
																assign node27512 = (inp[9]) ? 4'b1011 : 4'b1111;
											assign node27516 = (inp[15]) ? node27548 : node27517;
												assign node27517 = (inp[0]) ? node27533 : node27518;
													assign node27518 = (inp[3]) ? node27526 : node27519;
														assign node27519 = (inp[9]) ? node27523 : node27520;
															assign node27520 = (inp[4]) ? 4'b1111 : 4'b1011;
															assign node27523 = (inp[4]) ? 4'b1011 : 4'b1111;
														assign node27526 = (inp[4]) ? node27530 : node27527;
															assign node27527 = (inp[9]) ? 4'b1101 : 4'b1011;
															assign node27530 = (inp[9]) ? 4'b1001 : 4'b1101;
													assign node27533 = (inp[3]) ? node27541 : node27534;
														assign node27534 = (inp[10]) ? node27536 : 4'b1001;
															assign node27536 = (inp[9]) ? 4'b1001 : node27537;
																assign node27537 = (inp[4]) ? 4'b1101 : 4'b1001;
														assign node27541 = (inp[4]) ? node27545 : node27542;
															assign node27542 = (inp[9]) ? 4'b1111 : 4'b1001;
															assign node27545 = (inp[9]) ? 4'b1011 : 4'b1111;
												assign node27548 = (inp[0]) ? node27562 : node27549;
													assign node27549 = (inp[3]) ? node27557 : node27550;
														assign node27550 = (inp[4]) ? node27554 : node27551;
															assign node27551 = (inp[9]) ? 4'b1101 : 4'b1001;
															assign node27554 = (inp[9]) ? 4'b1001 : 4'b1101;
														assign node27557 = (inp[9]) ? node27559 : 4'b1001;
															assign node27559 = (inp[4]) ? 4'b1011 : 4'b1111;
													assign node27562 = (inp[3]) ? node27570 : node27563;
														assign node27563 = (inp[9]) ? node27567 : node27564;
															assign node27564 = (inp[4]) ? 4'b1111 : 4'b1011;
															assign node27567 = (inp[4]) ? 4'b1011 : 4'b1111;
														assign node27570 = (inp[10]) ? node27576 : node27571;
															assign node27571 = (inp[9]) ? node27573 : 4'b1101;
																assign node27573 = (inp[4]) ? 4'b1001 : 4'b1101;
															assign node27576 = (inp[4]) ? node27578 : 4'b1011;
																assign node27578 = (inp[9]) ? 4'b1001 : 4'b1101;
										assign node27581 = (inp[10]) ? node27675 : node27582;
											assign node27582 = (inp[9]) ? node27632 : node27583;
												assign node27583 = (inp[3]) ? node27613 : node27584;
													assign node27584 = (inp[12]) ? node27600 : node27585;
														assign node27585 = (inp[4]) ? node27593 : node27586;
															assign node27586 = (inp[0]) ? node27590 : node27587;
																assign node27587 = (inp[15]) ? 4'b1101 : 4'b1111;
																assign node27590 = (inp[15]) ? 4'b1111 : 4'b1101;
															assign node27593 = (inp[15]) ? node27597 : node27594;
																assign node27594 = (inp[0]) ? 4'b1001 : 4'b1011;
																assign node27597 = (inp[0]) ? 4'b1011 : 4'b1001;
														assign node27600 = (inp[4]) ? node27606 : node27601;
															assign node27601 = (inp[15]) ? node27603 : 4'b1001;
																assign node27603 = (inp[0]) ? 4'b1011 : 4'b1001;
															assign node27606 = (inp[0]) ? node27610 : node27607;
																assign node27607 = (inp[15]) ? 4'b1111 : 4'b1101;
																assign node27610 = (inp[15]) ? 4'b1101 : 4'b1111;
													assign node27613 = (inp[4]) ? node27625 : node27614;
														assign node27614 = (inp[12]) ? node27620 : node27615;
															assign node27615 = (inp[15]) ? node27617 : 4'b1101;
																assign node27617 = (inp[0]) ? 4'b1101 : 4'b1111;
															assign node27620 = (inp[0]) ? node27622 : 4'b1011;
																assign node27622 = (inp[15]) ? 4'b1001 : 4'b1011;
														assign node27625 = (inp[12]) ? 4'b1111 : node27626;
															assign node27626 = (inp[15]) ? 4'b1011 : node27627;
																assign node27627 = (inp[0]) ? 4'b1011 : 4'b1001;
												assign node27632 = (inp[15]) ? node27656 : node27633;
													assign node27633 = (inp[0]) ? node27649 : node27634;
														assign node27634 = (inp[3]) ? node27642 : node27635;
															assign node27635 = (inp[12]) ? node27639 : node27636;
																assign node27636 = (inp[4]) ? 4'b1101 : 4'b1011;
																assign node27639 = (inp[4]) ? 4'b1001 : 4'b1101;
															assign node27642 = (inp[12]) ? node27646 : node27643;
																assign node27643 = (inp[4]) ? 4'b1101 : 4'b1001;
																assign node27646 = (inp[4]) ? 4'b1001 : 4'b1101;
														assign node27649 = (inp[12]) ? node27653 : node27650;
															assign node27650 = (inp[4]) ? 4'b1111 : 4'b1001;
															assign node27653 = (inp[4]) ? 4'b1011 : 4'b1111;
													assign node27656 = (inp[0]) ? node27666 : node27657;
														assign node27657 = (inp[3]) ? node27663 : node27658;
															assign node27658 = (inp[4]) ? node27660 : 4'b1001;
																assign node27660 = (inp[12]) ? 4'b1011 : 4'b1111;
															assign node27663 = (inp[12]) ? 4'b1111 : 4'b1011;
														assign node27666 = (inp[12]) ? node27672 : node27667;
															assign node27667 = (inp[4]) ? 4'b1101 : node27668;
																assign node27668 = (inp[3]) ? 4'b1001 : 4'b1011;
															assign node27672 = (inp[4]) ? 4'b1001 : 4'b1101;
											assign node27675 = (inp[4]) ? node27713 : node27676;
												assign node27676 = (inp[9]) ? node27694 : node27677;
													assign node27677 = (inp[0]) ? node27687 : node27678;
														assign node27678 = (inp[12]) ? 4'b1001 : node27679;
															assign node27679 = (inp[15]) ? node27683 : node27680;
																assign node27680 = (inp[3]) ? 4'b1001 : 4'b1011;
																assign node27683 = (inp[3]) ? 4'b1011 : 4'b1001;
														assign node27687 = (inp[15]) ? node27691 : node27688;
															assign node27688 = (inp[3]) ? 4'b1011 : 4'b1001;
															assign node27691 = (inp[3]) ? 4'b1001 : 4'b1011;
													assign node27694 = (inp[12]) ? node27702 : node27695;
														assign node27695 = (inp[0]) ? node27699 : node27696;
															assign node27696 = (inp[15]) ? 4'b1111 : 4'b1101;
															assign node27699 = (inp[15]) ? 4'b1101 : 4'b1111;
														assign node27702 = (inp[3]) ? node27708 : node27703;
															assign node27703 = (inp[0]) ? 4'b1111 : node27704;
																assign node27704 = (inp[15]) ? 4'b1111 : 4'b1101;
															assign node27708 = (inp[15]) ? node27710 : 4'b1111;
																assign node27710 = (inp[0]) ? 4'b1101 : 4'b1111;
												assign node27713 = (inp[9]) ? node27733 : node27714;
													assign node27714 = (inp[3]) ? node27722 : node27715;
														assign node27715 = (inp[15]) ? node27719 : node27716;
															assign node27716 = (inp[0]) ? 4'b1111 : 4'b1101;
															assign node27719 = (inp[0]) ? 4'b1101 : 4'b1111;
														assign node27722 = (inp[12]) ? node27728 : node27723;
															assign node27723 = (inp[15]) ? node27725 : 4'b1101;
																assign node27725 = (inp[0]) ? 4'b1101 : 4'b1111;
															assign node27728 = (inp[15]) ? 4'b1101 : node27729;
																assign node27729 = (inp[0]) ? 4'b1111 : 4'b1101;
													assign node27733 = (inp[12]) ? node27739 : node27734;
														assign node27734 = (inp[15]) ? node27736 : 4'b1011;
															assign node27736 = (inp[0]) ? 4'b1001 : 4'b1011;
														assign node27739 = (inp[3]) ? node27745 : node27740;
															assign node27740 = (inp[15]) ? node27742 : 4'b1001;
																assign node27742 = (inp[0]) ? 4'b1001 : 4'b1011;
															assign node27745 = (inp[0]) ? node27747 : 4'b1001;
																assign node27747 = (inp[15]) ? 4'b1001 : 4'b1011;
							assign node27750 = (inp[14]) ? node28364 : node27751;
								assign node27751 = (inp[2]) ? node28037 : node27752;
									assign node27752 = (inp[5]) ? node27904 : node27753;
										assign node27753 = (inp[4]) ? node27821 : node27754;
											assign node27754 = (inp[9]) ? node27786 : node27755;
												assign node27755 = (inp[10]) ? node27771 : node27756;
													assign node27756 = (inp[12]) ? node27764 : node27757;
														assign node27757 = (inp[15]) ? node27761 : node27758;
															assign node27758 = (inp[0]) ? 4'b1101 : 4'b1111;
															assign node27761 = (inp[0]) ? 4'b1111 : 4'b1101;
														assign node27764 = (inp[0]) ? node27768 : node27765;
															assign node27765 = (inp[15]) ? 4'b1001 : 4'b1011;
															assign node27768 = (inp[15]) ? 4'b1011 : 4'b1001;
													assign node27771 = (inp[3]) ? node27773 : 4'b1001;
														assign node27773 = (inp[12]) ? node27781 : node27774;
															assign node27774 = (inp[15]) ? node27778 : node27775;
																assign node27775 = (inp[0]) ? 4'b1001 : 4'b1011;
																assign node27778 = (inp[0]) ? 4'b1011 : 4'b1001;
															assign node27781 = (inp[0]) ? 4'b1001 : node27782;
																assign node27782 = (inp[15]) ? 4'b1001 : 4'b1011;
												assign node27786 = (inp[10]) ? node27800 : node27787;
													assign node27787 = (inp[12]) ? node27791 : node27788;
														assign node27788 = (inp[15]) ? 4'b1011 : 4'b1001;
														assign node27791 = (inp[0]) ? 4'b1111 : node27792;
															assign node27792 = (inp[3]) ? node27796 : node27793;
																assign node27793 = (inp[15]) ? 4'b1101 : 4'b1111;
																assign node27796 = (inp[15]) ? 4'b1111 : 4'b1101;
													assign node27800 = (inp[12]) ? node27814 : node27801;
														assign node27801 = (inp[0]) ? node27807 : node27802;
															assign node27802 = (inp[3]) ? 4'b1111 : node27803;
																assign node27803 = (inp[15]) ? 4'b1101 : 4'b1111;
															assign node27807 = (inp[15]) ? node27811 : node27808;
																assign node27808 = (inp[3]) ? 4'b1111 : 4'b1101;
																assign node27811 = (inp[3]) ? 4'b1101 : 4'b1111;
														assign node27814 = (inp[15]) ? node27816 : 4'b1101;
															assign node27816 = (inp[3]) ? node27818 : 4'b1101;
																assign node27818 = (inp[0]) ? 4'b1101 : 4'b1111;
											assign node27821 = (inp[9]) ? node27863 : node27822;
												assign node27822 = (inp[10]) ? node27850 : node27823;
													assign node27823 = (inp[12]) ? node27839 : node27824;
														assign node27824 = (inp[3]) ? node27832 : node27825;
															assign node27825 = (inp[0]) ? node27829 : node27826;
																assign node27826 = (inp[15]) ? 4'b1001 : 4'b1011;
																assign node27829 = (inp[15]) ? 4'b1011 : 4'b1001;
															assign node27832 = (inp[15]) ? node27836 : node27833;
																assign node27833 = (inp[0]) ? 4'b1001 : 4'b1011;
																assign node27836 = (inp[0]) ? 4'b1011 : 4'b1001;
														assign node27839 = (inp[15]) ? node27845 : node27840;
															assign node27840 = (inp[3]) ? 4'b1111 : node27841;
																assign node27841 = (inp[0]) ? 4'b1101 : 4'b1111;
															assign node27845 = (inp[0]) ? 4'b1101 : node27846;
																assign node27846 = (inp[3]) ? 4'b1111 : 4'b1101;
													assign node27850 = (inp[0]) ? node27858 : node27851;
														assign node27851 = (inp[3]) ? node27855 : node27852;
															assign node27852 = (inp[15]) ? 4'b1101 : 4'b1111;
															assign node27855 = (inp[15]) ? 4'b1111 : 4'b1101;
														assign node27858 = (inp[15]) ? 4'b1111 : node27859;
															assign node27859 = (inp[3]) ? 4'b1111 : 4'b1101;
												assign node27863 = (inp[10]) ? node27881 : node27864;
													assign node27864 = (inp[12]) ? node27878 : node27865;
														assign node27865 = (inp[3]) ? node27873 : node27866;
															assign node27866 = (inp[15]) ? node27870 : node27867;
																assign node27867 = (inp[0]) ? 4'b1101 : 4'b1111;
																assign node27870 = (inp[0]) ? 4'b1111 : 4'b1101;
															assign node27873 = (inp[0]) ? 4'b1101 : node27874;
																assign node27874 = (inp[15]) ? 4'b1111 : 4'b1101;
														assign node27878 = (inp[3]) ? 4'b1001 : 4'b1011;
													assign node27881 = (inp[12]) ? node27895 : node27882;
														assign node27882 = (inp[0]) ? node27890 : node27883;
															assign node27883 = (inp[3]) ? node27887 : node27884;
																assign node27884 = (inp[15]) ? 4'b1001 : 4'b1011;
																assign node27887 = (inp[15]) ? 4'b1011 : 4'b1001;
															assign node27890 = (inp[15]) ? node27892 : 4'b1011;
																assign node27892 = (inp[3]) ? 4'b1001 : 4'b1011;
														assign node27895 = (inp[15]) ? node27897 : 4'b1001;
															assign node27897 = (inp[3]) ? node27901 : node27898;
																assign node27898 = (inp[0]) ? 4'b1011 : 4'b1001;
																assign node27901 = (inp[0]) ? 4'b1001 : 4'b1011;
										assign node27904 = (inp[12]) ? node27986 : node27905;
											assign node27905 = (inp[4]) ? node27945 : node27906;
												assign node27906 = (inp[10]) ? node27928 : node27907;
													assign node27907 = (inp[9]) ? node27915 : node27908;
														assign node27908 = (inp[15]) ? 4'b1111 : node27909;
															assign node27909 = (inp[0]) ? 4'b1101 : node27910;
																assign node27910 = (inp[3]) ? 4'b1101 : 4'b1111;
														assign node27915 = (inp[0]) ? node27923 : node27916;
															assign node27916 = (inp[15]) ? node27920 : node27917;
																assign node27917 = (inp[3]) ? 4'b1001 : 4'b1011;
																assign node27920 = (inp[3]) ? 4'b1011 : 4'b1001;
															assign node27923 = (inp[3]) ? node27925 : 4'b1001;
																assign node27925 = (inp[15]) ? 4'b1001 : 4'b1011;
													assign node27928 = (inp[9]) ? node27938 : node27929;
														assign node27929 = (inp[3]) ? 4'b1011 : node27930;
															assign node27930 = (inp[15]) ? node27934 : node27931;
																assign node27931 = (inp[0]) ? 4'b1001 : 4'b1011;
																assign node27934 = (inp[0]) ? 4'b1011 : 4'b1001;
														assign node27938 = (inp[0]) ? node27942 : node27939;
															assign node27939 = (inp[15]) ? 4'b1111 : 4'b1101;
															assign node27942 = (inp[15]) ? 4'b1101 : 4'b1111;
												assign node27945 = (inp[15]) ? node27963 : node27946;
													assign node27946 = (inp[0]) ? node27956 : node27947;
														assign node27947 = (inp[10]) ? node27953 : node27948;
															assign node27948 = (inp[9]) ? 4'b1101 : node27949;
																assign node27949 = (inp[3]) ? 4'b1001 : 4'b1011;
															assign node27953 = (inp[9]) ? 4'b1001 : 4'b1101;
														assign node27956 = (inp[10]) ? node27960 : node27957;
															assign node27957 = (inp[9]) ? 4'b1111 : 4'b1001;
															assign node27960 = (inp[9]) ? 4'b1011 : 4'b1111;
													assign node27963 = (inp[0]) ? node27973 : node27964;
														assign node27964 = (inp[9]) ? node27970 : node27965;
															assign node27965 = (inp[10]) ? 4'b1111 : node27966;
																assign node27966 = (inp[3]) ? 4'b1011 : 4'b1001;
															assign node27970 = (inp[10]) ? 4'b1011 : 4'b1111;
														assign node27973 = (inp[3]) ? node27979 : node27974;
															assign node27974 = (inp[10]) ? node27976 : 4'b1011;
																assign node27976 = (inp[9]) ? 4'b1001 : 4'b1101;
															assign node27979 = (inp[9]) ? node27983 : node27980;
																assign node27980 = (inp[10]) ? 4'b1101 : 4'b1001;
																assign node27983 = (inp[10]) ? 4'b1001 : 4'b1101;
											assign node27986 = (inp[0]) ? node28006 : node27987;
												assign node27987 = (inp[15]) ? node27997 : node27988;
													assign node27988 = (inp[4]) ? node27994 : node27989;
														assign node27989 = (inp[9]) ? 4'b1101 : node27990;
															assign node27990 = (inp[3]) ? 4'b1001 : 4'b1011;
														assign node27994 = (inp[9]) ? 4'b1001 : 4'b1101;
													assign node27997 = (inp[9]) ? node28003 : node27998;
														assign node27998 = (inp[4]) ? 4'b1111 : node27999;
															assign node27999 = (inp[3]) ? 4'b1011 : 4'b1001;
														assign node28003 = (inp[4]) ? 4'b1011 : 4'b1111;
												assign node28006 = (inp[15]) ? node28028 : node28007;
													assign node28007 = (inp[3]) ? node28013 : node28008;
														assign node28008 = (inp[4]) ? node28010 : 4'b1001;
															assign node28010 = (inp[9]) ? 4'b1011 : 4'b1111;
														assign node28013 = (inp[10]) ? node28021 : node28014;
															assign node28014 = (inp[4]) ? node28018 : node28015;
																assign node28015 = (inp[9]) ? 4'b1111 : 4'b1011;
																assign node28018 = (inp[9]) ? 4'b1011 : 4'b1111;
															assign node28021 = (inp[9]) ? node28025 : node28022;
																assign node28022 = (inp[4]) ? 4'b1111 : 4'b1011;
																assign node28025 = (inp[4]) ? 4'b1011 : 4'b1111;
													assign node28028 = (inp[4]) ? node28034 : node28029;
														assign node28029 = (inp[9]) ? 4'b1101 : node28030;
															assign node28030 = (inp[3]) ? 4'b1001 : 4'b1011;
														assign node28034 = (inp[9]) ? 4'b1001 : 4'b1101;
									assign node28037 = (inp[3]) ? node28179 : node28038;
										assign node28038 = (inp[4]) ? node28098 : node28039;
											assign node28039 = (inp[9]) ? node28065 : node28040;
												assign node28040 = (inp[12]) ? node28050 : node28041;
													assign node28041 = (inp[10]) ? 4'b1000 : node28042;
														assign node28042 = (inp[15]) ? node28046 : node28043;
															assign node28043 = (inp[0]) ? 4'b1100 : 4'b1110;
															assign node28046 = (inp[0]) ? 4'b1110 : 4'b1100;
													assign node28050 = (inp[10]) ? node28058 : node28051;
														assign node28051 = (inp[5]) ? 4'b1000 : node28052;
															assign node28052 = (inp[0]) ? node28054 : 4'b1000;
																assign node28054 = (inp[15]) ? 4'b1010 : 4'b1000;
														assign node28058 = (inp[15]) ? node28062 : node28059;
															assign node28059 = (inp[0]) ? 4'b1000 : 4'b1010;
															assign node28062 = (inp[0]) ? 4'b1010 : 4'b1000;
												assign node28065 = (inp[12]) ? node28085 : node28066;
													assign node28066 = (inp[10]) ? node28076 : node28067;
														assign node28067 = (inp[5]) ? 4'b1000 : node28068;
															assign node28068 = (inp[15]) ? node28072 : node28069;
																assign node28069 = (inp[0]) ? 4'b1000 : 4'b1010;
																assign node28072 = (inp[0]) ? 4'b1010 : 4'b1000;
														assign node28076 = (inp[0]) ? 4'b1100 : node28077;
															assign node28077 = (inp[15]) ? node28081 : node28078;
																assign node28078 = (inp[5]) ? 4'b1100 : 4'b1110;
																assign node28081 = (inp[5]) ? 4'b1110 : 4'b1100;
													assign node28085 = (inp[15]) ? node28093 : node28086;
														assign node28086 = (inp[5]) ? node28090 : node28087;
															assign node28087 = (inp[0]) ? 4'b1100 : 4'b1110;
															assign node28090 = (inp[0]) ? 4'b1110 : 4'b1100;
														assign node28093 = (inp[0]) ? node28095 : 4'b1100;
															assign node28095 = (inp[5]) ? 4'b1100 : 4'b1110;
											assign node28098 = (inp[9]) ? node28136 : node28099;
												assign node28099 = (inp[10]) ? node28121 : node28100;
													assign node28100 = (inp[12]) ? node28108 : node28101;
														assign node28101 = (inp[15]) ? node28105 : node28102;
															assign node28102 = (inp[0]) ? 4'b1000 : 4'b1010;
															assign node28105 = (inp[0]) ? 4'b1010 : 4'b1000;
														assign node28108 = (inp[0]) ? node28116 : node28109;
															assign node28109 = (inp[15]) ? node28113 : node28110;
																assign node28110 = (inp[5]) ? 4'b1100 : 4'b1110;
																assign node28113 = (inp[5]) ? 4'b1110 : 4'b1100;
															assign node28116 = (inp[15]) ? node28118 : 4'b1100;
																assign node28118 = (inp[5]) ? 4'b1100 : 4'b1110;
													assign node28121 = (inp[5]) ? node28129 : node28122;
														assign node28122 = (inp[0]) ? node28126 : node28123;
															assign node28123 = (inp[15]) ? 4'b1100 : 4'b1110;
															assign node28126 = (inp[15]) ? 4'b1110 : 4'b1100;
														assign node28129 = (inp[15]) ? node28133 : node28130;
															assign node28130 = (inp[0]) ? 4'b1110 : 4'b1100;
															assign node28133 = (inp[0]) ? 4'b1100 : 4'b1110;
												assign node28136 = (inp[12]) ? node28164 : node28137;
													assign node28137 = (inp[10]) ? node28151 : node28138;
														assign node28138 = (inp[15]) ? node28146 : node28139;
															assign node28139 = (inp[5]) ? node28143 : node28140;
																assign node28140 = (inp[0]) ? 4'b1100 : 4'b1110;
																assign node28143 = (inp[0]) ? 4'b1110 : 4'b1100;
															assign node28146 = (inp[5]) ? 4'b1100 : node28147;
																assign node28147 = (inp[0]) ? 4'b1110 : 4'b1100;
														assign node28151 = (inp[0]) ? node28159 : node28152;
															assign node28152 = (inp[5]) ? node28156 : node28153;
																assign node28153 = (inp[15]) ? 4'b1000 : 4'b1010;
																assign node28156 = (inp[15]) ? 4'b1010 : 4'b1000;
															assign node28159 = (inp[15]) ? 4'b1000 : node28160;
																assign node28160 = (inp[5]) ? 4'b1010 : 4'b1000;
													assign node28164 = (inp[5]) ? node28172 : node28165;
														assign node28165 = (inp[0]) ? node28169 : node28166;
															assign node28166 = (inp[15]) ? 4'b1000 : 4'b1010;
															assign node28169 = (inp[15]) ? 4'b1010 : 4'b1000;
														assign node28172 = (inp[15]) ? node28176 : node28173;
															assign node28173 = (inp[0]) ? 4'b1010 : 4'b1000;
															assign node28176 = (inp[0]) ? 4'b1000 : 4'b1010;
										assign node28179 = (inp[10]) ? node28283 : node28180;
											assign node28180 = (inp[12]) ? node28242 : node28181;
												assign node28181 = (inp[0]) ? node28211 : node28182;
													assign node28182 = (inp[15]) ? node28198 : node28183;
														assign node28183 = (inp[5]) ? node28191 : node28184;
															assign node28184 = (inp[4]) ? node28188 : node28185;
																assign node28185 = (inp[9]) ? 4'b1010 : 4'b1110;
																assign node28188 = (inp[9]) ? 4'b1100 : 4'b1010;
															assign node28191 = (inp[9]) ? node28195 : node28192;
																assign node28192 = (inp[4]) ? 4'b1000 : 4'b1100;
																assign node28195 = (inp[4]) ? 4'b1100 : 4'b1000;
														assign node28198 = (inp[5]) ? node28204 : node28199;
															assign node28199 = (inp[9]) ? node28201 : 4'b1000;
																assign node28201 = (inp[4]) ? 4'b1110 : 4'b1000;
															assign node28204 = (inp[9]) ? node28208 : node28205;
																assign node28205 = (inp[4]) ? 4'b1010 : 4'b1110;
																assign node28208 = (inp[4]) ? 4'b1110 : 4'b1010;
													assign node28211 = (inp[15]) ? node28227 : node28212;
														assign node28212 = (inp[5]) ? node28220 : node28213;
															assign node28213 = (inp[4]) ? node28217 : node28214;
																assign node28214 = (inp[9]) ? 4'b1000 : 4'b1100;
																assign node28217 = (inp[9]) ? 4'b1110 : 4'b1000;
															assign node28220 = (inp[9]) ? node28224 : node28221;
																assign node28221 = (inp[4]) ? 4'b1010 : 4'b1110;
																assign node28224 = (inp[4]) ? 4'b1110 : 4'b1010;
														assign node28227 = (inp[5]) ? node28235 : node28228;
															assign node28228 = (inp[4]) ? node28232 : node28229;
																assign node28229 = (inp[9]) ? 4'b1010 : 4'b1110;
																assign node28232 = (inp[9]) ? 4'b1100 : 4'b1010;
															assign node28235 = (inp[9]) ? node28239 : node28236;
																assign node28236 = (inp[4]) ? 4'b1000 : 4'b1100;
																assign node28239 = (inp[4]) ? 4'b1100 : 4'b1000;
												assign node28242 = (inp[0]) ? node28260 : node28243;
													assign node28243 = (inp[15]) ? node28251 : node28244;
														assign node28244 = (inp[9]) ? node28248 : node28245;
															assign node28245 = (inp[5]) ? 4'b1000 : 4'b1010;
															assign node28248 = (inp[4]) ? 4'b1000 : 4'b1100;
														assign node28251 = (inp[9]) ? node28257 : node28252;
															assign node28252 = (inp[4]) ? 4'b1110 : node28253;
																assign node28253 = (inp[5]) ? 4'b1010 : 4'b1000;
															assign node28257 = (inp[4]) ? 4'b1010 : 4'b1110;
													assign node28260 = (inp[15]) ? node28274 : node28261;
														assign node28261 = (inp[5]) ? node28267 : node28262;
															assign node28262 = (inp[9]) ? 4'b1110 : node28263;
																assign node28263 = (inp[4]) ? 4'b1110 : 4'b1000;
															assign node28267 = (inp[9]) ? node28271 : node28268;
																assign node28268 = (inp[4]) ? 4'b1110 : 4'b1010;
																assign node28271 = (inp[4]) ? 4'b1010 : 4'b1110;
														assign node28274 = (inp[9]) ? node28280 : node28275;
															assign node28275 = (inp[4]) ? 4'b1100 : node28276;
																assign node28276 = (inp[5]) ? 4'b1000 : 4'b1010;
															assign node28280 = (inp[4]) ? 4'b1000 : 4'b1100;
											assign node28283 = (inp[4]) ? node28327 : node28284;
												assign node28284 = (inp[9]) ? node28304 : node28285;
													assign node28285 = (inp[12]) ? node28291 : node28286;
														assign node28286 = (inp[0]) ? 4'b1010 : node28287;
															assign node28287 = (inp[15]) ? 4'b1010 : 4'b1000;
														assign node28291 = (inp[5]) ? node28297 : node28292;
															assign node28292 = (inp[0]) ? node28294 : 4'b1000;
																assign node28294 = (inp[15]) ? 4'b1010 : 4'b1000;
															assign node28297 = (inp[0]) ? node28301 : node28298;
																assign node28298 = (inp[15]) ? 4'b1010 : 4'b1000;
																assign node28301 = (inp[15]) ? 4'b1000 : 4'b1010;
													assign node28304 = (inp[12]) ? node28320 : node28305;
														assign node28305 = (inp[5]) ? node28313 : node28306;
															assign node28306 = (inp[0]) ? node28310 : node28307;
																assign node28307 = (inp[15]) ? 4'b1110 : 4'b1100;
																assign node28310 = (inp[15]) ? 4'b1100 : 4'b1110;
															assign node28313 = (inp[0]) ? node28317 : node28314;
																assign node28314 = (inp[15]) ? 4'b1110 : 4'b1100;
																assign node28317 = (inp[15]) ? 4'b1100 : 4'b1110;
														assign node28320 = (inp[0]) ? node28324 : node28321;
															assign node28321 = (inp[15]) ? 4'b1110 : 4'b1100;
															assign node28324 = (inp[15]) ? 4'b1100 : 4'b1110;
												assign node28327 = (inp[9]) ? node28345 : node28328;
													assign node28328 = (inp[12]) ? node28336 : node28329;
														assign node28329 = (inp[5]) ? 4'b1100 : node28330;
															assign node28330 = (inp[0]) ? node28332 : 4'b1100;
																assign node28332 = (inp[15]) ? 4'b1100 : 4'b1110;
														assign node28336 = (inp[5]) ? node28342 : node28337;
															assign node28337 = (inp[15]) ? 4'b1110 : node28338;
																assign node28338 = (inp[0]) ? 4'b1110 : 4'b1100;
															assign node28342 = (inp[0]) ? 4'b1100 : 4'b1110;
													assign node28345 = (inp[5]) ? node28357 : node28346;
														assign node28346 = (inp[12]) ? node28352 : node28347;
															assign node28347 = (inp[15]) ? 4'b1000 : node28348;
																assign node28348 = (inp[0]) ? 4'b1010 : 4'b1000;
															assign node28352 = (inp[0]) ? 4'b1000 : node28353;
																assign node28353 = (inp[15]) ? 4'b1010 : 4'b1000;
														assign node28357 = (inp[0]) ? node28361 : node28358;
															assign node28358 = (inp[15]) ? 4'b1010 : 4'b1000;
															assign node28361 = (inp[15]) ? 4'b1000 : 4'b1010;
								assign node28364 = (inp[15]) ? node28586 : node28365;
									assign node28365 = (inp[0]) ? node28479 : node28366;
										assign node28366 = (inp[3]) ? node28436 : node28367;
											assign node28367 = (inp[5]) ? node28415 : node28368;
												assign node28368 = (inp[12]) ? node28394 : node28369;
													assign node28369 = (inp[10]) ? node28379 : node28370;
														assign node28370 = (inp[2]) ? node28374 : node28371;
															assign node28371 = (inp[9]) ? 4'b1010 : 4'b1110;
															assign node28374 = (inp[4]) ? node28376 : 4'b1010;
																assign node28376 = (inp[9]) ? 4'b1110 : 4'b1010;
														assign node28379 = (inp[2]) ? node28387 : node28380;
															assign node28380 = (inp[9]) ? node28384 : node28381;
																assign node28381 = (inp[4]) ? 4'b1110 : 4'b1010;
																assign node28384 = (inp[4]) ? 4'b1010 : 4'b1110;
															assign node28387 = (inp[9]) ? node28391 : node28388;
																assign node28388 = (inp[4]) ? 4'b1110 : 4'b1010;
																assign node28391 = (inp[4]) ? 4'b1010 : 4'b1110;
													assign node28394 = (inp[2]) ? node28410 : node28395;
														assign node28395 = (inp[10]) ? node28403 : node28396;
															assign node28396 = (inp[4]) ? node28400 : node28397;
																assign node28397 = (inp[9]) ? 4'b1110 : 4'b1010;
																assign node28400 = (inp[9]) ? 4'b1010 : 4'b1110;
															assign node28403 = (inp[9]) ? node28407 : node28404;
																assign node28404 = (inp[4]) ? 4'b1110 : 4'b1010;
																assign node28407 = (inp[4]) ? 4'b1010 : 4'b1110;
														assign node28410 = (inp[9]) ? 4'b1110 : node28411;
															assign node28411 = (inp[4]) ? 4'b1110 : 4'b1010;
												assign node28415 = (inp[4]) ? node28427 : node28416;
													assign node28416 = (inp[9]) ? node28422 : node28417;
														assign node28417 = (inp[10]) ? 4'b1010 : node28418;
															assign node28418 = (inp[12]) ? 4'b1010 : 4'b1110;
														assign node28422 = (inp[12]) ? 4'b1100 : node28423;
															assign node28423 = (inp[10]) ? 4'b1100 : 4'b1010;
													assign node28427 = (inp[9]) ? node28433 : node28428;
														assign node28428 = (inp[12]) ? 4'b1100 : node28429;
															assign node28429 = (inp[10]) ? 4'b1100 : 4'b1010;
														assign node28433 = (inp[12]) ? 4'b1000 : 4'b1100;
											assign node28436 = (inp[5]) ? node28458 : node28437;
												assign node28437 = (inp[4]) ? node28447 : node28438;
													assign node28438 = (inp[9]) ? node28444 : node28439;
														assign node28439 = (inp[12]) ? 4'b1010 : node28440;
															assign node28440 = (inp[10]) ? 4'b1010 : 4'b1110;
														assign node28444 = (inp[12]) ? 4'b1100 : 4'b1010;
													assign node28447 = (inp[9]) ? node28453 : node28448;
														assign node28448 = (inp[12]) ? 4'b1100 : node28449;
															assign node28449 = (inp[10]) ? 4'b1100 : 4'b1010;
														assign node28453 = (inp[12]) ? 4'b1000 : node28454;
															assign node28454 = (inp[10]) ? 4'b1000 : 4'b1100;
												assign node28458 = (inp[12]) ? node28474 : node28459;
													assign node28459 = (inp[10]) ? node28467 : node28460;
														assign node28460 = (inp[9]) ? node28464 : node28461;
															assign node28461 = (inp[4]) ? 4'b1000 : 4'b1100;
															assign node28464 = (inp[4]) ? 4'b1100 : 4'b1000;
														assign node28467 = (inp[4]) ? node28471 : node28468;
															assign node28468 = (inp[9]) ? 4'b1100 : 4'b1000;
															assign node28471 = (inp[9]) ? 4'b1000 : 4'b1100;
													assign node28474 = (inp[9]) ? 4'b1100 : node28475;
														assign node28475 = (inp[4]) ? 4'b1100 : 4'b1000;
										assign node28479 = (inp[3]) ? node28545 : node28480;
											assign node28480 = (inp[5]) ? node28520 : node28481;
												assign node28481 = (inp[2]) ? node28503 : node28482;
													assign node28482 = (inp[12]) ? node28496 : node28483;
														assign node28483 = (inp[4]) ? node28491 : node28484;
															assign node28484 = (inp[10]) ? node28488 : node28485;
																assign node28485 = (inp[9]) ? 4'b1000 : 4'b1100;
																assign node28488 = (inp[9]) ? 4'b1100 : 4'b1000;
															assign node28491 = (inp[9]) ? 4'b1000 : node28492;
																assign node28492 = (inp[10]) ? 4'b1100 : 4'b1000;
														assign node28496 = (inp[4]) ? node28500 : node28497;
															assign node28497 = (inp[9]) ? 4'b1100 : 4'b1000;
															assign node28500 = (inp[9]) ? 4'b1000 : 4'b1100;
													assign node28503 = (inp[10]) ? node28515 : node28504;
														assign node28504 = (inp[9]) ? node28510 : node28505;
															assign node28505 = (inp[12]) ? node28507 : 4'b1000;
																assign node28507 = (inp[4]) ? 4'b1100 : 4'b1000;
															assign node28510 = (inp[4]) ? 4'b1100 : node28511;
																assign node28511 = (inp[12]) ? 4'b1100 : 4'b1000;
														assign node28515 = (inp[4]) ? node28517 : 4'b1100;
															assign node28517 = (inp[9]) ? 4'b1000 : 4'b1100;
												assign node28520 = (inp[9]) ? node28534 : node28521;
													assign node28521 = (inp[4]) ? node28527 : node28522;
														assign node28522 = (inp[12]) ? 4'b1000 : node28523;
															assign node28523 = (inp[10]) ? 4'b1000 : 4'b1100;
														assign node28527 = (inp[2]) ? node28529 : 4'b1110;
															assign node28529 = (inp[10]) ? 4'b1110 : node28530;
																assign node28530 = (inp[12]) ? 4'b1110 : 4'b1000;
													assign node28534 = (inp[4]) ? node28540 : node28535;
														assign node28535 = (inp[12]) ? 4'b1110 : node28536;
															assign node28536 = (inp[10]) ? 4'b1110 : 4'b1000;
														assign node28540 = (inp[12]) ? 4'b1010 : node28541;
															assign node28541 = (inp[10]) ? 4'b1010 : 4'b1110;
											assign node28545 = (inp[5]) ? node28563 : node28546;
												assign node28546 = (inp[9]) ? node28558 : node28547;
													assign node28547 = (inp[4]) ? node28553 : node28548;
														assign node28548 = (inp[12]) ? 4'b1000 : node28549;
															assign node28549 = (inp[10]) ? 4'b1000 : 4'b1100;
														assign node28553 = (inp[10]) ? 4'b1110 : node28554;
															assign node28554 = (inp[12]) ? 4'b1110 : 4'b1000;
													assign node28558 = (inp[4]) ? node28560 : 4'b1110;
														assign node28560 = (inp[10]) ? 4'b1010 : 4'b1110;
												assign node28563 = (inp[4]) ? node28575 : node28564;
													assign node28564 = (inp[9]) ? node28570 : node28565;
														assign node28565 = (inp[10]) ? 4'b1010 : node28566;
															assign node28566 = (inp[12]) ? 4'b1010 : 4'b1110;
														assign node28570 = (inp[10]) ? 4'b1110 : node28571;
															assign node28571 = (inp[12]) ? 4'b1110 : 4'b1010;
													assign node28575 = (inp[9]) ? node28581 : node28576;
														assign node28576 = (inp[12]) ? 4'b1110 : node28577;
															assign node28577 = (inp[10]) ? 4'b1110 : 4'b1010;
														assign node28581 = (inp[10]) ? 4'b1010 : node28582;
															assign node28582 = (inp[12]) ? 4'b1010 : 4'b1110;
									assign node28586 = (inp[0]) ? node28702 : node28587;
										assign node28587 = (inp[3]) ? node28655 : node28588;
											assign node28588 = (inp[5]) ? node28634 : node28589;
												assign node28589 = (inp[2]) ? node28615 : node28590;
													assign node28590 = (inp[10]) ? node28600 : node28591;
														assign node28591 = (inp[12]) ? node28593 : 4'b1000;
															assign node28593 = (inp[4]) ? node28597 : node28594;
																assign node28594 = (inp[9]) ? 4'b1100 : 4'b1000;
																assign node28597 = (inp[9]) ? 4'b1000 : 4'b1100;
														assign node28600 = (inp[12]) ? node28608 : node28601;
															assign node28601 = (inp[9]) ? node28605 : node28602;
																assign node28602 = (inp[4]) ? 4'b1100 : 4'b1000;
																assign node28605 = (inp[4]) ? 4'b1000 : 4'b1100;
															assign node28608 = (inp[9]) ? node28612 : node28609;
																assign node28609 = (inp[4]) ? 4'b1100 : 4'b1000;
																assign node28612 = (inp[4]) ? 4'b1000 : 4'b1100;
													assign node28615 = (inp[4]) ? node28623 : node28616;
														assign node28616 = (inp[9]) ? 4'b1100 : node28617;
															assign node28617 = (inp[12]) ? 4'b1000 : node28618;
																assign node28618 = (inp[10]) ? 4'b1000 : 4'b1100;
														assign node28623 = (inp[9]) ? node28629 : node28624;
															assign node28624 = (inp[12]) ? 4'b1100 : node28625;
																assign node28625 = (inp[10]) ? 4'b1100 : 4'b1000;
															assign node28629 = (inp[12]) ? 4'b1000 : node28630;
																assign node28630 = (inp[10]) ? 4'b1000 : 4'b1100;
												assign node28634 = (inp[9]) ? node28644 : node28635;
													assign node28635 = (inp[4]) ? node28641 : node28636;
														assign node28636 = (inp[12]) ? 4'b1000 : node28637;
															assign node28637 = (inp[10]) ? 4'b1000 : 4'b1100;
														assign node28641 = (inp[12]) ? 4'b1110 : 4'b1000;
													assign node28644 = (inp[4]) ? node28650 : node28645;
														assign node28645 = (inp[10]) ? 4'b1110 : node28646;
															assign node28646 = (inp[12]) ? 4'b1110 : 4'b1000;
														assign node28650 = (inp[10]) ? 4'b1010 : node28651;
															assign node28651 = (inp[2]) ? 4'b1110 : 4'b1010;
											assign node28655 = (inp[5]) ? node28679 : node28656;
												assign node28656 = (inp[9]) ? node28668 : node28657;
													assign node28657 = (inp[4]) ? node28663 : node28658;
														assign node28658 = (inp[12]) ? 4'b1000 : node28659;
															assign node28659 = (inp[10]) ? 4'b1000 : 4'b1100;
														assign node28663 = (inp[10]) ? 4'b1110 : node28664;
															assign node28664 = (inp[12]) ? 4'b1110 : 4'b1000;
													assign node28668 = (inp[4]) ? node28674 : node28669;
														assign node28669 = (inp[10]) ? 4'b1110 : node28670;
															assign node28670 = (inp[12]) ? 4'b1110 : 4'b1000;
														assign node28674 = (inp[10]) ? 4'b1010 : node28675;
															assign node28675 = (inp[12]) ? 4'b1010 : 4'b1110;
												assign node28679 = (inp[9]) ? node28691 : node28680;
													assign node28680 = (inp[4]) ? node28686 : node28681;
														assign node28681 = (inp[10]) ? 4'b1010 : node28682;
															assign node28682 = (inp[12]) ? 4'b1010 : 4'b1110;
														assign node28686 = (inp[10]) ? 4'b1110 : node28687;
															assign node28687 = (inp[12]) ? 4'b1110 : 4'b1010;
													assign node28691 = (inp[4]) ? node28697 : node28692;
														assign node28692 = (inp[12]) ? 4'b1110 : node28693;
															assign node28693 = (inp[10]) ? 4'b1110 : 4'b1010;
														assign node28697 = (inp[10]) ? 4'b1010 : node28698;
															assign node28698 = (inp[12]) ? 4'b1010 : 4'b1110;
										assign node28702 = (inp[5]) ? node28748 : node28703;
											assign node28703 = (inp[3]) ? node28725 : node28704;
												assign node28704 = (inp[4]) ? node28716 : node28705;
													assign node28705 = (inp[9]) ? node28711 : node28706;
														assign node28706 = (inp[12]) ? 4'b1010 : node28707;
															assign node28707 = (inp[10]) ? 4'b1010 : 4'b1110;
														assign node28711 = (inp[12]) ? 4'b1110 : node28712;
															assign node28712 = (inp[10]) ? 4'b1110 : 4'b1010;
													assign node28716 = (inp[9]) ? node28720 : node28717;
														assign node28717 = (inp[10]) ? 4'b1110 : 4'b1010;
														assign node28720 = (inp[12]) ? 4'b1010 : node28721;
															assign node28721 = (inp[10]) ? 4'b1010 : 4'b1110;
												assign node28725 = (inp[4]) ? node28737 : node28726;
													assign node28726 = (inp[9]) ? node28732 : node28727;
														assign node28727 = (inp[12]) ? 4'b1010 : node28728;
															assign node28728 = (inp[10]) ? 4'b1010 : 4'b1110;
														assign node28732 = (inp[12]) ? 4'b1100 : node28733;
															assign node28733 = (inp[10]) ? 4'b1100 : 4'b1010;
													assign node28737 = (inp[9]) ? node28743 : node28738;
														assign node28738 = (inp[12]) ? 4'b1100 : node28739;
															assign node28739 = (inp[10]) ? 4'b1100 : 4'b1010;
														assign node28743 = (inp[10]) ? 4'b1000 : node28744;
															assign node28744 = (inp[12]) ? 4'b1000 : 4'b1100;
											assign node28748 = (inp[3]) ? node28770 : node28749;
												assign node28749 = (inp[4]) ? node28761 : node28750;
													assign node28750 = (inp[9]) ? node28756 : node28751;
														assign node28751 = (inp[10]) ? 4'b1010 : node28752;
															assign node28752 = (inp[12]) ? 4'b1010 : 4'b1110;
														assign node28756 = (inp[10]) ? 4'b1100 : node28757;
															assign node28757 = (inp[12]) ? 4'b1100 : 4'b1010;
													assign node28761 = (inp[9]) ? node28767 : node28762;
														assign node28762 = (inp[10]) ? 4'b1100 : node28763;
															assign node28763 = (inp[2]) ? 4'b1010 : 4'b1100;
														assign node28767 = (inp[10]) ? 4'b1000 : 4'b1100;
												assign node28770 = (inp[12]) ? node28798 : node28771;
													assign node28771 = (inp[2]) ? node28785 : node28772;
														assign node28772 = (inp[10]) ? node28780 : node28773;
															assign node28773 = (inp[9]) ? node28777 : node28774;
																assign node28774 = (inp[4]) ? 4'b1000 : 4'b1100;
																assign node28777 = (inp[4]) ? 4'b1100 : 4'b1000;
															assign node28780 = (inp[4]) ? node28782 : 4'b1100;
																assign node28782 = (inp[9]) ? 4'b1000 : 4'b1100;
														assign node28785 = (inp[10]) ? node28791 : node28786;
															assign node28786 = (inp[4]) ? node28788 : 4'b1000;
																assign node28788 = (inp[9]) ? 4'b1100 : 4'b1000;
															assign node28791 = (inp[4]) ? node28795 : node28792;
																assign node28792 = (inp[9]) ? 4'b1100 : 4'b1000;
																assign node28795 = (inp[9]) ? 4'b1000 : 4'b1100;
													assign node28798 = (inp[10]) ? node28806 : node28799;
														assign node28799 = (inp[9]) ? node28803 : node28800;
															assign node28800 = (inp[4]) ? 4'b1100 : 4'b1000;
															assign node28803 = (inp[4]) ? 4'b1000 : 4'b1100;
														assign node28806 = (inp[9]) ? node28808 : 4'b1000;
															assign node28808 = (inp[4]) ? 4'b1000 : 4'b1100;
					assign node28811 = (inp[10]) ? node31063 : node28812;
						assign node28812 = (inp[8]) ? node29978 : node28813;
							assign node28813 = (inp[7]) ? node29319 : node28814;
								assign node28814 = (inp[2]) ? node29136 : node28815;
									assign node28815 = (inp[14]) ? node28991 : node28816;
										assign node28816 = (inp[3]) ? node28916 : node28817;
											assign node28817 = (inp[0]) ? node28863 : node28818;
												assign node28818 = (inp[15]) ? node28846 : node28819;
													assign node28819 = (inp[5]) ? node28835 : node28820;
														assign node28820 = (inp[12]) ? node28828 : node28821;
															assign node28821 = (inp[9]) ? node28825 : node28822;
																assign node28822 = (inp[4]) ? 4'b1011 : 4'b1111;
																assign node28825 = (inp[4]) ? 4'b1111 : 4'b1011;
															assign node28828 = (inp[9]) ? node28832 : node28829;
																assign node28829 = (inp[4]) ? 4'b1111 : 4'b1011;
																assign node28832 = (inp[4]) ? 4'b1011 : 4'b1111;
														assign node28835 = (inp[12]) ? node28841 : node28836;
															assign node28836 = (inp[9]) ? 4'b1011 : node28837;
																assign node28837 = (inp[4]) ? 4'b1011 : 4'b1111;
															assign node28841 = (inp[9]) ? node28843 : 4'b1011;
																assign node28843 = (inp[4]) ? 4'b1001 : 4'b1101;
													assign node28846 = (inp[5]) ? node28852 : node28847;
														assign node28847 = (inp[12]) ? node28849 : 4'b1001;
															assign node28849 = (inp[4]) ? 4'b1101 : 4'b1001;
														assign node28852 = (inp[12]) ? node28856 : node28853;
															assign node28853 = (inp[4]) ? 4'b1001 : 4'b1101;
															assign node28856 = (inp[9]) ? node28860 : node28857;
																assign node28857 = (inp[4]) ? 4'b1111 : 4'b1001;
																assign node28860 = (inp[4]) ? 4'b1011 : 4'b1111;
												assign node28863 = (inp[15]) ? node28893 : node28864;
													assign node28864 = (inp[5]) ? node28880 : node28865;
														assign node28865 = (inp[4]) ? node28873 : node28866;
															assign node28866 = (inp[12]) ? node28870 : node28867;
																assign node28867 = (inp[9]) ? 4'b1001 : 4'b1101;
																assign node28870 = (inp[9]) ? 4'b1101 : 4'b1001;
															assign node28873 = (inp[9]) ? node28877 : node28874;
																assign node28874 = (inp[12]) ? 4'b1101 : 4'b1001;
																assign node28877 = (inp[12]) ? 4'b1001 : 4'b1101;
														assign node28880 = (inp[12]) ? node28888 : node28881;
															assign node28881 = (inp[9]) ? node28885 : node28882;
																assign node28882 = (inp[4]) ? 4'b1001 : 4'b1101;
																assign node28885 = (inp[4]) ? 4'b1111 : 4'b1001;
															assign node28888 = (inp[4]) ? 4'b1111 : node28889;
																assign node28889 = (inp[9]) ? 4'b1111 : 4'b1001;
													assign node28893 = (inp[5]) ? node28907 : node28894;
														assign node28894 = (inp[4]) ? node28900 : node28895;
															assign node28895 = (inp[12]) ? 4'b1011 : node28896;
																assign node28896 = (inp[9]) ? 4'b1011 : 4'b1111;
															assign node28900 = (inp[9]) ? node28904 : node28901;
																assign node28901 = (inp[12]) ? 4'b1111 : 4'b1011;
																assign node28904 = (inp[12]) ? 4'b1011 : 4'b1111;
														assign node28907 = (inp[9]) ? 4'b1101 : node28908;
															assign node28908 = (inp[12]) ? node28912 : node28909;
																assign node28909 = (inp[4]) ? 4'b1011 : 4'b1111;
																assign node28912 = (inp[4]) ? 4'b1101 : 4'b1011;
											assign node28916 = (inp[5]) ? node28960 : node28917;
												assign node28917 = (inp[4]) ? node28939 : node28918;
													assign node28918 = (inp[15]) ? node28928 : node28919;
														assign node28919 = (inp[0]) ? node28921 : 4'b1101;
															assign node28921 = (inp[12]) ? node28925 : node28922;
																assign node28922 = (inp[9]) ? 4'b1001 : 4'b1101;
																assign node28925 = (inp[9]) ? 4'b1111 : 4'b1001;
														assign node28928 = (inp[9]) ? node28936 : node28929;
															assign node28929 = (inp[0]) ? node28933 : node28930;
																assign node28930 = (inp[12]) ? 4'b1001 : 4'b1101;
																assign node28933 = (inp[12]) ? 4'b1011 : 4'b1111;
															assign node28936 = (inp[0]) ? 4'b1101 : 4'b1111;
													assign node28939 = (inp[0]) ? node28949 : node28940;
														assign node28940 = (inp[15]) ? node28946 : node28941;
															assign node28941 = (inp[9]) ? 4'b1101 : node28942;
																assign node28942 = (inp[12]) ? 4'b1101 : 4'b1011;
															assign node28946 = (inp[9]) ? 4'b1011 : 4'b1111;
														assign node28949 = (inp[9]) ? node28953 : node28950;
															assign node28950 = (inp[15]) ? 4'b1011 : 4'b1001;
															assign node28953 = (inp[12]) ? node28957 : node28954;
																assign node28954 = (inp[15]) ? 4'b1101 : 4'b1111;
																assign node28957 = (inp[15]) ? 4'b1001 : 4'b1011;
												assign node28960 = (inp[0]) ? node28980 : node28961;
													assign node28961 = (inp[15]) ? node28973 : node28962;
														assign node28962 = (inp[4]) ? node28968 : node28963;
															assign node28963 = (inp[9]) ? 4'b1101 : node28964;
																assign node28964 = (inp[12]) ? 4'b1001 : 4'b1101;
															assign node28968 = (inp[12]) ? node28970 : 4'b1001;
																assign node28970 = (inp[9]) ? 4'b1001 : 4'b1101;
														assign node28973 = (inp[4]) ? node28975 : 4'b1011;
															assign node28975 = (inp[12]) ? 4'b1111 : node28976;
																assign node28976 = (inp[9]) ? 4'b1111 : 4'b1011;
													assign node28980 = (inp[15]) ? node28982 : 4'b1011;
														assign node28982 = (inp[12]) ? 4'b1001 : node28983;
															assign node28983 = (inp[4]) ? node28987 : node28984;
																assign node28984 = (inp[9]) ? 4'b1001 : 4'b1101;
																assign node28987 = (inp[9]) ? 4'b1101 : 4'b1001;
										assign node28991 = (inp[4]) ? node29057 : node28992;
											assign node28992 = (inp[15]) ? node29028 : node28993;
												assign node28993 = (inp[12]) ? node29013 : node28994;
													assign node28994 = (inp[9]) ? node29002 : node28995;
														assign node28995 = (inp[5]) ? node28999 : node28996;
															assign node28996 = (inp[0]) ? 4'b1100 : 4'b1110;
															assign node28999 = (inp[0]) ? 4'b1110 : 4'b1100;
														assign node29002 = (inp[0]) ? node29008 : node29003;
															assign node29003 = (inp[5]) ? node29005 : 4'b1010;
																assign node29005 = (inp[3]) ? 4'b1000 : 4'b1010;
															assign node29008 = (inp[3]) ? node29010 : 4'b1000;
																assign node29010 = (inp[5]) ? 4'b1010 : 4'b1000;
													assign node29013 = (inp[9]) ? node29021 : node29014;
														assign node29014 = (inp[0]) ? node29016 : 4'b1010;
															assign node29016 = (inp[3]) ? node29018 : 4'b1000;
																assign node29018 = (inp[5]) ? 4'b1010 : 4'b1000;
														assign node29021 = (inp[0]) ? node29023 : 4'b1100;
															assign node29023 = (inp[5]) ? 4'b1110 : node29024;
																assign node29024 = (inp[3]) ? 4'b1110 : 4'b1100;
												assign node29028 = (inp[5]) ? node29036 : node29029;
													assign node29029 = (inp[0]) ? node29031 : 4'b1000;
														assign node29031 = (inp[12]) ? node29033 : 4'b1010;
															assign node29033 = (inp[9]) ? 4'b1110 : 4'b1010;
													assign node29036 = (inp[0]) ? node29048 : node29037;
														assign node29037 = (inp[3]) ? node29041 : node29038;
															assign node29038 = (inp[9]) ? 4'b1110 : 4'b1100;
															assign node29041 = (inp[9]) ? node29045 : node29042;
																assign node29042 = (inp[12]) ? 4'b1010 : 4'b1110;
																assign node29045 = (inp[12]) ? 4'b1110 : 4'b1010;
														assign node29048 = (inp[3]) ? node29054 : node29049;
															assign node29049 = (inp[9]) ? node29051 : 4'b1010;
																assign node29051 = (inp[12]) ? 4'b1100 : 4'b1010;
															assign node29054 = (inp[12]) ? 4'b1000 : 4'b1100;
											assign node29057 = (inp[3]) ? node29103 : node29058;
												assign node29058 = (inp[9]) ? node29074 : node29059;
													assign node29059 = (inp[12]) ? node29067 : node29060;
														assign node29060 = (inp[15]) ? node29064 : node29061;
															assign node29061 = (inp[0]) ? 4'b1000 : 4'b1010;
															assign node29064 = (inp[0]) ? 4'b1010 : 4'b1000;
														assign node29067 = (inp[0]) ? 4'b1110 : node29068;
															assign node29068 = (inp[5]) ? 4'b1100 : node29069;
																assign node29069 = (inp[15]) ? 4'b1100 : 4'b1110;
													assign node29074 = (inp[12]) ? node29090 : node29075;
														assign node29075 = (inp[5]) ? node29083 : node29076;
															assign node29076 = (inp[15]) ? node29080 : node29077;
																assign node29077 = (inp[0]) ? 4'b1100 : 4'b1110;
																assign node29080 = (inp[0]) ? 4'b1110 : 4'b1100;
															assign node29083 = (inp[0]) ? node29087 : node29084;
																assign node29084 = (inp[15]) ? 4'b1110 : 4'b1100;
																assign node29087 = (inp[15]) ? 4'b1100 : 4'b1110;
														assign node29090 = (inp[15]) ? node29098 : node29091;
															assign node29091 = (inp[5]) ? node29095 : node29092;
																assign node29092 = (inp[0]) ? 4'b1000 : 4'b1010;
																assign node29095 = (inp[0]) ? 4'b1010 : 4'b1000;
															assign node29098 = (inp[0]) ? 4'b1000 : node29099;
																assign node29099 = (inp[5]) ? 4'b1010 : 4'b1000;
												assign node29103 = (inp[5]) ? node29119 : node29104;
													assign node29104 = (inp[9]) ? node29114 : node29105;
														assign node29105 = (inp[12]) ? node29111 : node29106;
															assign node29106 = (inp[15]) ? node29108 : 4'b1010;
																assign node29108 = (inp[0]) ? 4'b1010 : 4'b1000;
															assign node29111 = (inp[15]) ? 4'b1110 : 4'b1100;
														assign node29114 = (inp[12]) ? 4'b1000 : node29115;
															assign node29115 = (inp[0]) ? 4'b1100 : 4'b1110;
													assign node29119 = (inp[9]) ? node29129 : node29120;
														assign node29120 = (inp[12]) ? node29122 : 4'b1000;
															assign node29122 = (inp[0]) ? node29126 : node29123;
																assign node29123 = (inp[15]) ? 4'b1110 : 4'b1100;
																assign node29126 = (inp[15]) ? 4'b1100 : 4'b1110;
														assign node29129 = (inp[12]) ? 4'b1000 : node29130;
															assign node29130 = (inp[15]) ? node29132 : 4'b1110;
																assign node29132 = (inp[0]) ? 4'b1100 : 4'b1110;
									assign node29136 = (inp[12]) ? node29228 : node29137;
										assign node29137 = (inp[9]) ? node29183 : node29138;
											assign node29138 = (inp[4]) ? node29162 : node29139;
												assign node29139 = (inp[0]) ? node29151 : node29140;
													assign node29140 = (inp[15]) ? node29146 : node29141;
														assign node29141 = (inp[5]) ? node29143 : 4'b1110;
															assign node29143 = (inp[3]) ? 4'b1100 : 4'b1110;
														assign node29146 = (inp[5]) ? node29148 : 4'b1100;
															assign node29148 = (inp[3]) ? 4'b1110 : 4'b1100;
													assign node29151 = (inp[15]) ? node29157 : node29152;
														assign node29152 = (inp[5]) ? node29154 : 4'b1100;
															assign node29154 = (inp[3]) ? 4'b1110 : 4'b1100;
														assign node29157 = (inp[5]) ? node29159 : 4'b1110;
															assign node29159 = (inp[3]) ? 4'b1100 : 4'b1110;
												assign node29162 = (inp[15]) ? node29172 : node29163;
													assign node29163 = (inp[5]) ? node29165 : 4'b1010;
														assign node29165 = (inp[0]) ? node29169 : node29166;
															assign node29166 = (inp[3]) ? 4'b1000 : 4'b1010;
															assign node29169 = (inp[3]) ? 4'b1010 : 4'b1000;
													assign node29172 = (inp[0]) ? node29178 : node29173;
														assign node29173 = (inp[3]) ? node29175 : 4'b1000;
															assign node29175 = (inp[5]) ? 4'b1010 : 4'b1000;
														assign node29178 = (inp[5]) ? node29180 : 4'b1010;
															assign node29180 = (inp[3]) ? 4'b1000 : 4'b1010;
											assign node29183 = (inp[4]) ? node29205 : node29184;
												assign node29184 = (inp[15]) ? node29196 : node29185;
													assign node29185 = (inp[0]) ? node29191 : node29186;
														assign node29186 = (inp[3]) ? node29188 : 4'b1010;
															assign node29188 = (inp[5]) ? 4'b1000 : 4'b1010;
														assign node29191 = (inp[5]) ? node29193 : 4'b1000;
															assign node29193 = (inp[3]) ? 4'b1010 : 4'b1000;
													assign node29196 = (inp[0]) ? node29202 : node29197;
														assign node29197 = (inp[5]) ? node29199 : 4'b1000;
															assign node29199 = (inp[3]) ? 4'b1010 : 4'b1000;
														assign node29202 = (inp[5]) ? 4'b1000 : 4'b1010;
												assign node29205 = (inp[0]) ? node29217 : node29206;
													assign node29206 = (inp[15]) ? node29212 : node29207;
														assign node29207 = (inp[5]) ? 4'b1100 : node29208;
															assign node29208 = (inp[3]) ? 4'b1100 : 4'b1110;
														assign node29212 = (inp[3]) ? 4'b1110 : node29213;
															assign node29213 = (inp[14]) ? 4'b1110 : 4'b1100;
													assign node29217 = (inp[14]) ? 4'b1100 : node29218;
														assign node29218 = (inp[15]) ? node29222 : node29219;
															assign node29219 = (inp[3]) ? 4'b1110 : 4'b1100;
															assign node29222 = (inp[5]) ? 4'b1100 : node29223;
																assign node29223 = (inp[3]) ? 4'b1100 : 4'b1110;
										assign node29228 = (inp[9]) ? node29274 : node29229;
											assign node29229 = (inp[4]) ? node29251 : node29230;
												assign node29230 = (inp[15]) ? node29242 : node29231;
													assign node29231 = (inp[0]) ? node29237 : node29232;
														assign node29232 = (inp[5]) ? node29234 : 4'b1010;
															assign node29234 = (inp[3]) ? 4'b1000 : 4'b1010;
														assign node29237 = (inp[5]) ? node29239 : 4'b1000;
															assign node29239 = (inp[3]) ? 4'b1010 : 4'b1000;
													assign node29242 = (inp[0]) ? node29246 : node29243;
														assign node29243 = (inp[3]) ? 4'b1010 : 4'b1000;
														assign node29246 = (inp[3]) ? node29248 : 4'b1010;
															assign node29248 = (inp[5]) ? 4'b1000 : 4'b1010;
												assign node29251 = (inp[0]) ? node29259 : node29252;
													assign node29252 = (inp[15]) ? node29256 : node29253;
														assign node29253 = (inp[3]) ? 4'b1100 : 4'b1110;
														assign node29256 = (inp[3]) ? 4'b1110 : 4'b1100;
													assign node29259 = (inp[3]) ? 4'b1100 : node29260;
														assign node29260 = (inp[14]) ? node29266 : node29261;
															assign node29261 = (inp[15]) ? node29263 : 4'b1100;
																assign node29263 = (inp[5]) ? 4'b1100 : 4'b1110;
															assign node29266 = (inp[5]) ? node29270 : node29267;
																assign node29267 = (inp[15]) ? 4'b1110 : 4'b1100;
																assign node29270 = (inp[15]) ? 4'b1100 : 4'b1110;
											assign node29274 = (inp[4]) ? node29294 : node29275;
												assign node29275 = (inp[0]) ? node29289 : node29276;
													assign node29276 = (inp[15]) ? node29284 : node29277;
														assign node29277 = (inp[14]) ? 4'b1100 : node29278;
															assign node29278 = (inp[3]) ? 4'b1100 : node29279;
																assign node29279 = (inp[5]) ? 4'b1100 : 4'b1110;
														assign node29284 = (inp[5]) ? 4'b1110 : node29285;
															assign node29285 = (inp[3]) ? 4'b1110 : 4'b1100;
													assign node29289 = (inp[15]) ? node29291 : 4'b1110;
														assign node29291 = (inp[3]) ? 4'b1100 : 4'b1110;
												assign node29294 = (inp[3]) ? node29312 : node29295;
													assign node29295 = (inp[0]) ? node29303 : node29296;
														assign node29296 = (inp[15]) ? node29300 : node29297;
															assign node29297 = (inp[5]) ? 4'b1000 : 4'b1010;
															assign node29300 = (inp[5]) ? 4'b1010 : 4'b1000;
														assign node29303 = (inp[14]) ? node29305 : 4'b1010;
															assign node29305 = (inp[15]) ? node29309 : node29306;
																assign node29306 = (inp[5]) ? 4'b1010 : 4'b1000;
																assign node29309 = (inp[5]) ? 4'b1000 : 4'b1010;
													assign node29312 = (inp[0]) ? node29316 : node29313;
														assign node29313 = (inp[15]) ? 4'b1010 : 4'b1000;
														assign node29316 = (inp[15]) ? 4'b1000 : 4'b1010;
								assign node29319 = (inp[14]) ? node29657 : node29320;
									assign node29320 = (inp[2]) ? node29480 : node29321;
										assign node29321 = (inp[12]) ? node29397 : node29322;
											assign node29322 = (inp[4]) ? node29360 : node29323;
												assign node29323 = (inp[9]) ? node29347 : node29324;
													assign node29324 = (inp[0]) ? node29336 : node29325;
														assign node29325 = (inp[15]) ? node29331 : node29326;
															assign node29326 = (inp[3]) ? node29328 : 4'b1110;
																assign node29328 = (inp[5]) ? 4'b1100 : 4'b1110;
															assign node29331 = (inp[3]) ? node29333 : 4'b1100;
																assign node29333 = (inp[5]) ? 4'b1110 : 4'b1100;
														assign node29336 = (inp[15]) ? node29342 : node29337;
															assign node29337 = (inp[5]) ? node29339 : 4'b1100;
																assign node29339 = (inp[3]) ? 4'b1110 : 4'b1100;
															assign node29342 = (inp[3]) ? node29344 : 4'b1110;
																assign node29344 = (inp[5]) ? 4'b1100 : 4'b1110;
													assign node29347 = (inp[3]) ? node29349 : 4'b1000;
														assign node29349 = (inp[0]) ? node29355 : node29350;
															assign node29350 = (inp[15]) ? node29352 : 4'b1000;
																assign node29352 = (inp[5]) ? 4'b1010 : 4'b1000;
															assign node29355 = (inp[15]) ? node29357 : 4'b1010;
																assign node29357 = (inp[5]) ? 4'b1000 : 4'b1010;
												assign node29360 = (inp[9]) ? node29380 : node29361;
													assign node29361 = (inp[3]) ? node29367 : node29362;
														assign node29362 = (inp[5]) ? 4'b1010 : node29363;
															assign node29363 = (inp[0]) ? 4'b1010 : 4'b1000;
														assign node29367 = (inp[5]) ? node29373 : node29368;
															assign node29368 = (inp[15]) ? node29370 : 4'b1000;
																assign node29370 = (inp[0]) ? 4'b1010 : 4'b1000;
															assign node29373 = (inp[0]) ? node29377 : node29374;
																assign node29374 = (inp[15]) ? 4'b1010 : 4'b1000;
																assign node29377 = (inp[15]) ? 4'b1000 : 4'b1010;
													assign node29380 = (inp[5]) ? node29390 : node29381;
														assign node29381 = (inp[3]) ? node29383 : 4'b1110;
															assign node29383 = (inp[0]) ? node29387 : node29384;
																assign node29384 = (inp[15]) ? 4'b1110 : 4'b1100;
																assign node29387 = (inp[15]) ? 4'b1100 : 4'b1110;
														assign node29390 = (inp[15]) ? node29394 : node29391;
															assign node29391 = (inp[0]) ? 4'b1110 : 4'b1100;
															assign node29394 = (inp[0]) ? 4'b1100 : 4'b1110;
											assign node29397 = (inp[0]) ? node29435 : node29398;
												assign node29398 = (inp[4]) ? node29416 : node29399;
													assign node29399 = (inp[9]) ? node29407 : node29400;
														assign node29400 = (inp[15]) ? 4'b1000 : node29401;
															assign node29401 = (inp[3]) ? node29403 : 4'b1010;
																assign node29403 = (inp[5]) ? 4'b1000 : 4'b1010;
														assign node29407 = (inp[3]) ? node29413 : node29408;
															assign node29408 = (inp[5]) ? 4'b1110 : node29409;
																assign node29409 = (inp[15]) ? 4'b1100 : 4'b1110;
															assign node29413 = (inp[15]) ? 4'b1110 : 4'b1100;
													assign node29416 = (inp[9]) ? node29426 : node29417;
														assign node29417 = (inp[15]) ? node29421 : node29418;
															assign node29418 = (inp[5]) ? 4'b1100 : 4'b1110;
															assign node29421 = (inp[5]) ? 4'b1110 : node29422;
																assign node29422 = (inp[3]) ? 4'b1110 : 4'b1100;
														assign node29426 = (inp[15]) ? node29430 : node29427;
															assign node29427 = (inp[3]) ? 4'b1000 : 4'b1010;
															assign node29430 = (inp[3]) ? 4'b1010 : node29431;
																assign node29431 = (inp[5]) ? 4'b1010 : 4'b1000;
												assign node29435 = (inp[3]) ? node29461 : node29436;
													assign node29436 = (inp[15]) ? node29448 : node29437;
														assign node29437 = (inp[5]) ? node29443 : node29438;
															assign node29438 = (inp[4]) ? 4'b1100 : node29439;
																assign node29439 = (inp[9]) ? 4'b1100 : 4'b1000;
															assign node29443 = (inp[9]) ? node29445 : 4'b1000;
																assign node29445 = (inp[4]) ? 4'b1010 : 4'b1110;
														assign node29448 = (inp[5]) ? node29456 : node29449;
															assign node29449 = (inp[4]) ? node29453 : node29450;
																assign node29450 = (inp[9]) ? 4'b1110 : 4'b1010;
																assign node29453 = (inp[9]) ? 4'b1010 : 4'b1110;
															assign node29456 = (inp[4]) ? node29458 : 4'b1010;
																assign node29458 = (inp[9]) ? 4'b1000 : 4'b1100;
													assign node29461 = (inp[15]) ? node29471 : node29462;
														assign node29462 = (inp[5]) ? node29466 : node29463;
															assign node29463 = (inp[9]) ? 4'b1010 : 4'b1000;
															assign node29466 = (inp[9]) ? 4'b1110 : node29467;
																assign node29467 = (inp[4]) ? 4'b1110 : 4'b1010;
														assign node29471 = (inp[4]) ? node29477 : node29472;
															assign node29472 = (inp[9]) ? 4'b1100 : node29473;
																assign node29473 = (inp[5]) ? 4'b1000 : 4'b1010;
															assign node29477 = (inp[9]) ? 4'b1000 : 4'b1100;
										assign node29480 = (inp[3]) ? node29570 : node29481;
											assign node29481 = (inp[4]) ? node29519 : node29482;
												assign node29482 = (inp[9]) ? node29494 : node29483;
													assign node29483 = (inp[12]) ? node29491 : node29484;
														assign node29484 = (inp[15]) ? node29488 : node29485;
															assign node29485 = (inp[0]) ? 4'b1101 : 4'b1111;
															assign node29488 = (inp[0]) ? 4'b1111 : 4'b1101;
														assign node29491 = (inp[5]) ? 4'b1001 : 4'b1011;
													assign node29494 = (inp[12]) ? node29508 : node29495;
														assign node29495 = (inp[5]) ? node29503 : node29496;
															assign node29496 = (inp[0]) ? node29500 : node29497;
																assign node29497 = (inp[15]) ? 4'b1001 : 4'b1011;
																assign node29500 = (inp[15]) ? 4'b1011 : 4'b1001;
															assign node29503 = (inp[0]) ? node29505 : 4'b1011;
																assign node29505 = (inp[15]) ? 4'b1011 : 4'b1001;
														assign node29508 = (inp[5]) ? node29514 : node29509;
															assign node29509 = (inp[0]) ? 4'b1111 : node29510;
																assign node29510 = (inp[15]) ? 4'b1101 : 4'b1111;
															assign node29514 = (inp[0]) ? node29516 : 4'b1101;
																assign node29516 = (inp[15]) ? 4'b1101 : 4'b1111;
												assign node29519 = (inp[5]) ? node29545 : node29520;
													assign node29520 = (inp[12]) ? node29534 : node29521;
														assign node29521 = (inp[9]) ? node29529 : node29522;
															assign node29522 = (inp[0]) ? node29526 : node29523;
																assign node29523 = (inp[15]) ? 4'b1001 : 4'b1011;
																assign node29526 = (inp[15]) ? 4'b1011 : 4'b1001;
															assign node29529 = (inp[15]) ? 4'b1101 : node29530;
																assign node29530 = (inp[0]) ? 4'b1101 : 4'b1111;
														assign node29534 = (inp[9]) ? node29540 : node29535;
															assign node29535 = (inp[15]) ? node29537 : 4'b1101;
																assign node29537 = (inp[0]) ? 4'b1111 : 4'b1101;
															assign node29540 = (inp[0]) ? node29542 : 4'b1001;
																assign node29542 = (inp[15]) ? 4'b1011 : 4'b1001;
													assign node29545 = (inp[9]) ? node29559 : node29546;
														assign node29546 = (inp[12]) ? node29554 : node29547;
															assign node29547 = (inp[0]) ? node29551 : node29548;
																assign node29548 = (inp[15]) ? 4'b1001 : 4'b1011;
																assign node29551 = (inp[15]) ? 4'b1011 : 4'b1001;
															assign node29554 = (inp[0]) ? node29556 : 4'b1101;
																assign node29556 = (inp[15]) ? 4'b1101 : 4'b1111;
														assign node29559 = (inp[12]) ? node29565 : node29560;
															assign node29560 = (inp[15]) ? 4'b1111 : node29561;
																assign node29561 = (inp[0]) ? 4'b1111 : 4'b1101;
															assign node29565 = (inp[0]) ? node29567 : 4'b1011;
																assign node29567 = (inp[15]) ? 4'b1001 : 4'b1011;
											assign node29570 = (inp[15]) ? node29618 : node29571;
												assign node29571 = (inp[0]) ? node29597 : node29572;
													assign node29572 = (inp[5]) ? node29584 : node29573;
														assign node29573 = (inp[4]) ? node29579 : node29574;
															assign node29574 = (inp[9]) ? 4'b1011 : node29575;
																assign node29575 = (inp[12]) ? 4'b1011 : 4'b1111;
															assign node29579 = (inp[12]) ? node29581 : 4'b1011;
																assign node29581 = (inp[9]) ? 4'b1001 : 4'b1101;
														assign node29584 = (inp[12]) ? node29590 : node29585;
															assign node29585 = (inp[9]) ? 4'b1001 : node29586;
																assign node29586 = (inp[4]) ? 4'b1001 : 4'b1101;
															assign node29590 = (inp[9]) ? node29594 : node29591;
																assign node29591 = (inp[4]) ? 4'b1101 : 4'b1001;
																assign node29594 = (inp[4]) ? 4'b1001 : 4'b1101;
													assign node29597 = (inp[4]) ? node29607 : node29598;
														assign node29598 = (inp[5]) ? node29604 : node29599;
															assign node29599 = (inp[9]) ? node29601 : 4'b1001;
																assign node29601 = (inp[12]) ? 4'b1111 : 4'b1001;
															assign node29604 = (inp[12]) ? 4'b1011 : 4'b1111;
														assign node29607 = (inp[5]) ? node29613 : node29608;
															assign node29608 = (inp[12]) ? node29610 : 4'b1111;
																assign node29610 = (inp[9]) ? 4'b1011 : 4'b1111;
															assign node29613 = (inp[9]) ? node29615 : 4'b1011;
																assign node29615 = (inp[12]) ? 4'b1011 : 4'b1111;
												assign node29618 = (inp[0]) ? node29636 : node29619;
													assign node29619 = (inp[5]) ? node29627 : node29620;
														assign node29620 = (inp[4]) ? node29622 : 4'b1001;
															assign node29622 = (inp[12]) ? node29624 : 4'b1001;
																assign node29624 = (inp[9]) ? 4'b1011 : 4'b1111;
														assign node29627 = (inp[9]) ? 4'b1111 : node29628;
															assign node29628 = (inp[12]) ? node29632 : node29629;
																assign node29629 = (inp[4]) ? 4'b1011 : 4'b1111;
																assign node29632 = (inp[4]) ? 4'b1111 : 4'b1011;
													assign node29636 = (inp[5]) ? node29648 : node29637;
														assign node29637 = (inp[9]) ? node29643 : node29638;
															assign node29638 = (inp[4]) ? 4'b1101 : node29639;
																assign node29639 = (inp[12]) ? 4'b1011 : 4'b1111;
															assign node29643 = (inp[4]) ? node29645 : 4'b1101;
																assign node29645 = (inp[12]) ? 4'b1001 : 4'b1101;
														assign node29648 = (inp[4]) ? 4'b1001 : node29649;
															assign node29649 = (inp[12]) ? node29653 : node29650;
																assign node29650 = (inp[9]) ? 4'b1001 : 4'b1101;
																assign node29653 = (inp[9]) ? 4'b1101 : 4'b1001;
									assign node29657 = (inp[3]) ? node29841 : node29658;
										assign node29658 = (inp[12]) ? node29744 : node29659;
											assign node29659 = (inp[5]) ? node29691 : node29660;
												assign node29660 = (inp[9]) ? node29674 : node29661;
													assign node29661 = (inp[4]) ? node29669 : node29662;
														assign node29662 = (inp[15]) ? node29666 : node29663;
															assign node29663 = (inp[0]) ? 4'b1101 : 4'b1111;
															assign node29666 = (inp[0]) ? 4'b1111 : 4'b1101;
														assign node29669 = (inp[15]) ? node29671 : 4'b1011;
															assign node29671 = (inp[0]) ? 4'b1011 : 4'b1001;
													assign node29674 = (inp[4]) ? node29682 : node29675;
														assign node29675 = (inp[15]) ? node29679 : node29676;
															assign node29676 = (inp[0]) ? 4'b1001 : 4'b1011;
															assign node29679 = (inp[0]) ? 4'b1011 : 4'b1001;
														assign node29682 = (inp[2]) ? 4'b1101 : node29683;
															assign node29683 = (inp[15]) ? node29687 : node29684;
																assign node29684 = (inp[0]) ? 4'b1101 : 4'b1111;
																assign node29687 = (inp[0]) ? 4'b1111 : 4'b1101;
												assign node29691 = (inp[2]) ? node29717 : node29692;
													assign node29692 = (inp[9]) ? node29706 : node29693;
														assign node29693 = (inp[4]) ? node29699 : node29694;
															assign node29694 = (inp[15]) ? node29696 : 4'b1111;
																assign node29696 = (inp[0]) ? 4'b1111 : 4'b1101;
															assign node29699 = (inp[15]) ? node29703 : node29700;
																assign node29700 = (inp[0]) ? 4'b1001 : 4'b1011;
																assign node29703 = (inp[0]) ? 4'b1011 : 4'b1001;
														assign node29706 = (inp[4]) ? node29710 : node29707;
															assign node29707 = (inp[0]) ? 4'b1001 : 4'b1011;
															assign node29710 = (inp[0]) ? node29714 : node29711;
																assign node29711 = (inp[15]) ? 4'b1111 : 4'b1101;
																assign node29714 = (inp[15]) ? 4'b1101 : 4'b1111;
													assign node29717 = (inp[9]) ? node29729 : node29718;
														assign node29718 = (inp[4]) ? node29724 : node29719;
															assign node29719 = (inp[15]) ? node29721 : 4'b1101;
																assign node29721 = (inp[0]) ? 4'b1111 : 4'b1101;
															assign node29724 = (inp[0]) ? node29726 : 4'b1001;
																assign node29726 = (inp[15]) ? 4'b1011 : 4'b1001;
														assign node29729 = (inp[4]) ? node29737 : node29730;
															assign node29730 = (inp[15]) ? node29734 : node29731;
																assign node29731 = (inp[0]) ? 4'b1001 : 4'b1011;
																assign node29734 = (inp[0]) ? 4'b1011 : 4'b1001;
															assign node29737 = (inp[15]) ? node29741 : node29738;
																assign node29738 = (inp[0]) ? 4'b1111 : 4'b1101;
																assign node29741 = (inp[0]) ? 4'b1101 : 4'b1111;
											assign node29744 = (inp[2]) ? node29802 : node29745;
												assign node29745 = (inp[15]) ? node29773 : node29746;
													assign node29746 = (inp[0]) ? node29760 : node29747;
														assign node29747 = (inp[5]) ? node29753 : node29748;
															assign node29748 = (inp[9]) ? node29750 : 4'b1111;
																assign node29750 = (inp[4]) ? 4'b1011 : 4'b1111;
															assign node29753 = (inp[4]) ? node29757 : node29754;
																assign node29754 = (inp[9]) ? 4'b1101 : 4'b1011;
																assign node29757 = (inp[9]) ? 4'b1001 : 4'b1101;
														assign node29760 = (inp[5]) ? node29768 : node29761;
															assign node29761 = (inp[4]) ? node29765 : node29762;
																assign node29762 = (inp[9]) ? 4'b1101 : 4'b1001;
																assign node29765 = (inp[9]) ? 4'b1001 : 4'b1101;
															assign node29768 = (inp[4]) ? node29770 : 4'b1001;
																assign node29770 = (inp[9]) ? 4'b1011 : 4'b1111;
													assign node29773 = (inp[0]) ? node29787 : node29774;
														assign node29774 = (inp[5]) ? node29780 : node29775;
															assign node29775 = (inp[4]) ? 4'b1001 : node29776;
																assign node29776 = (inp[9]) ? 4'b1101 : 4'b1001;
															assign node29780 = (inp[4]) ? node29784 : node29781;
																assign node29781 = (inp[9]) ? 4'b1111 : 4'b1001;
																assign node29784 = (inp[9]) ? 4'b1011 : 4'b1111;
														assign node29787 = (inp[5]) ? node29795 : node29788;
															assign node29788 = (inp[4]) ? node29792 : node29789;
																assign node29789 = (inp[9]) ? 4'b1111 : 4'b1011;
																assign node29792 = (inp[9]) ? 4'b1011 : 4'b1111;
															assign node29795 = (inp[9]) ? node29799 : node29796;
																assign node29796 = (inp[4]) ? 4'b1101 : 4'b1011;
																assign node29799 = (inp[4]) ? 4'b1001 : 4'b1101;
												assign node29802 = (inp[4]) ? node29820 : node29803;
													assign node29803 = (inp[9]) ? node29811 : node29804;
														assign node29804 = (inp[15]) ? node29808 : node29805;
															assign node29805 = (inp[0]) ? 4'b1001 : 4'b1011;
															assign node29808 = (inp[0]) ? 4'b1011 : 4'b1001;
														assign node29811 = (inp[5]) ? 4'b1101 : node29812;
															assign node29812 = (inp[0]) ? node29816 : node29813;
																assign node29813 = (inp[15]) ? 4'b1101 : 4'b1111;
																assign node29816 = (inp[15]) ? 4'b1111 : 4'b1101;
													assign node29820 = (inp[9]) ? node29834 : node29821;
														assign node29821 = (inp[15]) ? node29829 : node29822;
															assign node29822 = (inp[0]) ? node29826 : node29823;
																assign node29823 = (inp[5]) ? 4'b1101 : 4'b1111;
																assign node29826 = (inp[5]) ? 4'b1111 : 4'b1101;
															assign node29829 = (inp[5]) ? node29831 : 4'b1101;
																assign node29831 = (inp[0]) ? 4'b1101 : 4'b1111;
														assign node29834 = (inp[5]) ? node29836 : 4'b1001;
															assign node29836 = (inp[0]) ? 4'b1011 : node29837;
																assign node29837 = (inp[15]) ? 4'b1011 : 4'b1001;
										assign node29841 = (inp[4]) ? node29919 : node29842;
											assign node29842 = (inp[9]) ? node29884 : node29843;
												assign node29843 = (inp[12]) ? node29855 : node29844;
													assign node29844 = (inp[15]) ? 4'b1111 : node29845;
														assign node29845 = (inp[2]) ? 4'b1101 : node29846;
															assign node29846 = (inp[5]) ? node29850 : node29847;
																assign node29847 = (inp[0]) ? 4'b1101 : 4'b1111;
																assign node29850 = (inp[0]) ? 4'b1111 : 4'b1101;
													assign node29855 = (inp[2]) ? node29869 : node29856;
														assign node29856 = (inp[5]) ? node29864 : node29857;
															assign node29857 = (inp[15]) ? node29861 : node29858;
																assign node29858 = (inp[0]) ? 4'b1001 : 4'b1011;
																assign node29861 = (inp[0]) ? 4'b1011 : 4'b1001;
															assign node29864 = (inp[0]) ? node29866 : 4'b1011;
																assign node29866 = (inp[15]) ? 4'b1001 : 4'b1011;
														assign node29869 = (inp[0]) ? node29877 : node29870;
															assign node29870 = (inp[15]) ? node29874 : node29871;
																assign node29871 = (inp[5]) ? 4'b1001 : 4'b1011;
																assign node29874 = (inp[5]) ? 4'b1011 : 4'b1001;
															assign node29877 = (inp[15]) ? node29881 : node29878;
																assign node29878 = (inp[5]) ? 4'b1011 : 4'b1001;
																assign node29881 = (inp[5]) ? 4'b1001 : 4'b1011;
												assign node29884 = (inp[12]) ? node29908 : node29885;
													assign node29885 = (inp[2]) ? node29899 : node29886;
														assign node29886 = (inp[15]) ? node29892 : node29887;
															assign node29887 = (inp[0]) ? 4'b1001 : node29888;
																assign node29888 = (inp[5]) ? 4'b1001 : 4'b1011;
															assign node29892 = (inp[0]) ? node29896 : node29893;
																assign node29893 = (inp[5]) ? 4'b1011 : 4'b1001;
																assign node29896 = (inp[5]) ? 4'b1001 : 4'b1011;
														assign node29899 = (inp[15]) ? 4'b1001 : node29900;
															assign node29900 = (inp[5]) ? node29904 : node29901;
																assign node29901 = (inp[0]) ? 4'b1001 : 4'b1011;
																assign node29904 = (inp[0]) ? 4'b1011 : 4'b1001;
													assign node29908 = (inp[5]) ? node29914 : node29909;
														assign node29909 = (inp[0]) ? node29911 : 4'b1111;
															assign node29911 = (inp[15]) ? 4'b1101 : 4'b1111;
														assign node29914 = (inp[0]) ? node29916 : 4'b1101;
															assign node29916 = (inp[15]) ? 4'b1101 : 4'b1111;
											assign node29919 = (inp[9]) ? node29955 : node29920;
												assign node29920 = (inp[12]) ? node29942 : node29921;
													assign node29921 = (inp[2]) ? node29933 : node29922;
														assign node29922 = (inp[0]) ? node29928 : node29923;
															assign node29923 = (inp[15]) ? node29925 : 4'b1011;
																assign node29925 = (inp[5]) ? 4'b1011 : 4'b1001;
															assign node29928 = (inp[5]) ? node29930 : 4'b1001;
																assign node29930 = (inp[15]) ? 4'b1001 : 4'b1011;
														assign node29933 = (inp[0]) ? node29935 : 4'b1001;
															assign node29935 = (inp[5]) ? node29939 : node29936;
																assign node29936 = (inp[15]) ? 4'b1011 : 4'b1001;
																assign node29939 = (inp[15]) ? 4'b1001 : 4'b1011;
													assign node29942 = (inp[5]) ? node29950 : node29943;
														assign node29943 = (inp[0]) ? node29947 : node29944;
															assign node29944 = (inp[15]) ? 4'b1111 : 4'b1101;
															assign node29947 = (inp[15]) ? 4'b1101 : 4'b1111;
														assign node29950 = (inp[0]) ? node29952 : 4'b1101;
															assign node29952 = (inp[15]) ? 4'b1101 : 4'b1111;
												assign node29955 = (inp[12]) ? node29963 : node29956;
													assign node29956 = (inp[0]) ? node29960 : node29957;
														assign node29957 = (inp[15]) ? 4'b1111 : 4'b1101;
														assign node29960 = (inp[15]) ? 4'b1101 : 4'b1111;
													assign node29963 = (inp[2]) ? node29971 : node29964;
														assign node29964 = (inp[0]) ? node29968 : node29965;
															assign node29965 = (inp[15]) ? 4'b1011 : 4'b1001;
															assign node29968 = (inp[15]) ? 4'b1001 : 4'b1011;
														assign node29971 = (inp[15]) ? node29975 : node29972;
															assign node29972 = (inp[0]) ? 4'b1011 : 4'b1001;
															assign node29975 = (inp[0]) ? 4'b1001 : 4'b1011;
							assign node29978 = (inp[7]) ? node30510 : node29979;
								assign node29979 = (inp[14]) ? node30303 : node29980;
									assign node29980 = (inp[2]) ? node30148 : node29981;
										assign node29981 = (inp[15]) ? node30065 : node29982;
											assign node29982 = (inp[12]) ? node30022 : node29983;
												assign node29983 = (inp[9]) ? node30005 : node29984;
													assign node29984 = (inp[4]) ? node29996 : node29985;
														assign node29985 = (inp[0]) ? node29991 : node29986;
															assign node29986 = (inp[5]) ? node29988 : 4'b1110;
																assign node29988 = (inp[3]) ? 4'b1100 : 4'b1110;
															assign node29991 = (inp[5]) ? node29993 : 4'b1100;
																assign node29993 = (inp[3]) ? 4'b1110 : 4'b1100;
														assign node29996 = (inp[5]) ? node30000 : node29997;
															assign node29997 = (inp[0]) ? 4'b1000 : 4'b1010;
															assign node30000 = (inp[3]) ? node30002 : 4'b1010;
																assign node30002 = (inp[0]) ? 4'b1010 : 4'b1000;
													assign node30005 = (inp[4]) ? node30011 : node30006;
														assign node30006 = (inp[5]) ? node30008 : 4'b1010;
															assign node30008 = (inp[0]) ? 4'b1010 : 4'b1000;
														assign node30011 = (inp[0]) ? node30017 : node30012;
															assign node30012 = (inp[3]) ? 4'b1100 : node30013;
																assign node30013 = (inp[5]) ? 4'b1100 : 4'b1110;
															assign node30017 = (inp[5]) ? 4'b1110 : node30018;
																assign node30018 = (inp[3]) ? 4'b1110 : 4'b1100;
												assign node30022 = (inp[0]) ? node30046 : node30023;
													assign node30023 = (inp[5]) ? node30037 : node30024;
														assign node30024 = (inp[3]) ? node30032 : node30025;
															assign node30025 = (inp[4]) ? node30029 : node30026;
																assign node30026 = (inp[9]) ? 4'b1110 : 4'b1010;
																assign node30029 = (inp[9]) ? 4'b1010 : 4'b1110;
															assign node30032 = (inp[9]) ? node30034 : 4'b1010;
																assign node30034 = (inp[4]) ? 4'b1000 : 4'b1100;
														assign node30037 = (inp[4]) ? node30043 : node30038;
															assign node30038 = (inp[9]) ? 4'b1100 : node30039;
																assign node30039 = (inp[3]) ? 4'b1000 : 4'b1010;
															assign node30043 = (inp[9]) ? 4'b1000 : 4'b1100;
													assign node30046 = (inp[3]) ? node30060 : node30047;
														assign node30047 = (inp[5]) ? node30055 : node30048;
															assign node30048 = (inp[9]) ? node30052 : node30049;
																assign node30049 = (inp[4]) ? 4'b1100 : 4'b1000;
																assign node30052 = (inp[4]) ? 4'b1000 : 4'b1100;
															assign node30055 = (inp[4]) ? node30057 : 4'b1000;
																assign node30057 = (inp[9]) ? 4'b1010 : 4'b1110;
														assign node30060 = (inp[4]) ? node30062 : 4'b1110;
															assign node30062 = (inp[9]) ? 4'b1010 : 4'b1110;
											assign node30065 = (inp[12]) ? node30111 : node30066;
												assign node30066 = (inp[0]) ? node30090 : node30067;
													assign node30067 = (inp[3]) ? node30075 : node30068;
														assign node30068 = (inp[4]) ? node30072 : node30069;
															assign node30069 = (inp[9]) ? 4'b1000 : 4'b1100;
															assign node30072 = (inp[9]) ? 4'b1110 : 4'b1000;
														assign node30075 = (inp[5]) ? node30083 : node30076;
															assign node30076 = (inp[9]) ? node30080 : node30077;
																assign node30077 = (inp[4]) ? 4'b1000 : 4'b1100;
																assign node30080 = (inp[4]) ? 4'b1110 : 4'b1000;
															assign node30083 = (inp[4]) ? node30087 : node30084;
																assign node30084 = (inp[9]) ? 4'b1010 : 4'b1110;
																assign node30087 = (inp[9]) ? 4'b1110 : 4'b1010;
													assign node30090 = (inp[3]) ? node30100 : node30091;
														assign node30091 = (inp[4]) ? node30095 : node30092;
															assign node30092 = (inp[9]) ? 4'b1010 : 4'b1110;
															assign node30095 = (inp[9]) ? node30097 : 4'b1010;
																assign node30097 = (inp[5]) ? 4'b1100 : 4'b1110;
														assign node30100 = (inp[5]) ? node30106 : node30101;
															assign node30101 = (inp[4]) ? node30103 : 4'b1010;
																assign node30103 = (inp[9]) ? 4'b1100 : 4'b1010;
															assign node30106 = (inp[4]) ? 4'b1000 : node30107;
																assign node30107 = (inp[9]) ? 4'b1000 : 4'b1100;
												assign node30111 = (inp[0]) ? node30129 : node30112;
													assign node30112 = (inp[5]) ? node30122 : node30113;
														assign node30113 = (inp[9]) ? node30117 : node30114;
															assign node30114 = (inp[4]) ? 4'b1100 : 4'b1000;
															assign node30117 = (inp[4]) ? 4'b1000 : node30118;
																assign node30118 = (inp[3]) ? 4'b1110 : 4'b1100;
														assign node30122 = (inp[9]) ? node30126 : node30123;
															assign node30123 = (inp[4]) ? 4'b1110 : 4'b1000;
															assign node30126 = (inp[4]) ? 4'b1010 : 4'b1110;
													assign node30129 = (inp[5]) ? node30141 : node30130;
														assign node30130 = (inp[3]) ? node30138 : node30131;
															assign node30131 = (inp[4]) ? node30135 : node30132;
																assign node30132 = (inp[9]) ? 4'b1110 : 4'b1010;
																assign node30135 = (inp[9]) ? 4'b1010 : 4'b1110;
															assign node30138 = (inp[4]) ? 4'b1000 : 4'b1100;
														assign node30141 = (inp[4]) ? node30145 : node30142;
															assign node30142 = (inp[9]) ? 4'b1100 : 4'b1000;
															assign node30145 = (inp[9]) ? 4'b1000 : 4'b1100;
										assign node30148 = (inp[15]) ? node30220 : node30149;
											assign node30149 = (inp[4]) ? node30181 : node30150;
												assign node30150 = (inp[3]) ? node30166 : node30151;
													assign node30151 = (inp[0]) ? node30157 : node30152;
														assign node30152 = (inp[9]) ? node30154 : 4'b1011;
															assign node30154 = (inp[12]) ? 4'b1101 : 4'b1011;
														assign node30157 = (inp[5]) ? node30163 : node30158;
															assign node30158 = (inp[12]) ? node30160 : 4'b1001;
																assign node30160 = (inp[9]) ? 4'b1101 : 4'b1001;
															assign node30163 = (inp[12]) ? 4'b1001 : 4'b1101;
													assign node30166 = (inp[0]) ? node30176 : node30167;
														assign node30167 = (inp[5]) ? node30171 : node30168;
															assign node30168 = (inp[12]) ? 4'b1101 : 4'b1111;
															assign node30171 = (inp[9]) ? 4'b1101 : node30172;
																assign node30172 = (inp[12]) ? 4'b1001 : 4'b1101;
														assign node30176 = (inp[12]) ? 4'b1111 : node30177;
															assign node30177 = (inp[9]) ? 4'b1001 : 4'b1101;
												assign node30181 = (inp[3]) ? node30205 : node30182;
													assign node30182 = (inp[0]) ? node30192 : node30183;
														assign node30183 = (inp[5]) ? node30185 : 4'b1111;
															assign node30185 = (inp[9]) ? node30189 : node30186;
																assign node30186 = (inp[12]) ? 4'b1101 : 4'b1011;
																assign node30189 = (inp[12]) ? 4'b1001 : 4'b1101;
														assign node30192 = (inp[5]) ? node30200 : node30193;
															assign node30193 = (inp[9]) ? node30197 : node30194;
																assign node30194 = (inp[12]) ? 4'b1101 : 4'b1001;
																assign node30197 = (inp[12]) ? 4'b1001 : 4'b1101;
															assign node30200 = (inp[12]) ? 4'b1111 : node30201;
																assign node30201 = (inp[9]) ? 4'b1111 : 4'b1001;
													assign node30205 = (inp[0]) ? node30211 : node30206;
														assign node30206 = (inp[12]) ? 4'b1001 : node30207;
															assign node30207 = (inp[9]) ? 4'b1101 : 4'b1001;
														assign node30211 = (inp[12]) ? node30217 : node30212;
															assign node30212 = (inp[5]) ? node30214 : 4'b1001;
																assign node30214 = (inp[9]) ? 4'b1111 : 4'b1011;
															assign node30217 = (inp[9]) ? 4'b1011 : 4'b1111;
											assign node30220 = (inp[12]) ? node30264 : node30221;
												assign node30221 = (inp[0]) ? node30243 : node30222;
													assign node30222 = (inp[5]) ? node30230 : node30223;
														assign node30223 = (inp[9]) ? node30227 : node30224;
															assign node30224 = (inp[4]) ? 4'b1001 : 4'b1101;
															assign node30227 = (inp[3]) ? 4'b1111 : 4'b1101;
														assign node30230 = (inp[3]) ? node30236 : node30231;
															assign node30231 = (inp[4]) ? 4'b1111 : node30232;
																assign node30232 = (inp[9]) ? 4'b1001 : 4'b1101;
															assign node30236 = (inp[9]) ? node30240 : node30237;
																assign node30237 = (inp[4]) ? 4'b1011 : 4'b1111;
																assign node30240 = (inp[4]) ? 4'b1111 : 4'b1011;
													assign node30243 = (inp[3]) ? node30257 : node30244;
														assign node30244 = (inp[5]) ? node30252 : node30245;
															assign node30245 = (inp[9]) ? node30249 : node30246;
																assign node30246 = (inp[4]) ? 4'b1011 : 4'b1111;
																assign node30249 = (inp[4]) ? 4'b1111 : 4'b1011;
															assign node30252 = (inp[4]) ? 4'b1101 : node30253;
																assign node30253 = (inp[9]) ? 4'b1011 : 4'b1111;
														assign node30257 = (inp[5]) ? 4'b1001 : node30258;
															assign node30258 = (inp[4]) ? 4'b1101 : node30259;
																assign node30259 = (inp[9]) ? 4'b1011 : 4'b1111;
												assign node30264 = (inp[0]) ? node30284 : node30265;
													assign node30265 = (inp[5]) ? node30271 : node30266;
														assign node30266 = (inp[9]) ? node30268 : 4'b1001;
															assign node30268 = (inp[4]) ? 4'b1001 : 4'b1111;
														assign node30271 = (inp[3]) ? node30277 : node30272;
															assign node30272 = (inp[4]) ? 4'b1111 : node30273;
																assign node30273 = (inp[9]) ? 4'b1111 : 4'b1001;
															assign node30277 = (inp[9]) ? node30281 : node30278;
																assign node30278 = (inp[4]) ? 4'b1111 : 4'b1011;
																assign node30281 = (inp[4]) ? 4'b1011 : 4'b1111;
													assign node30284 = (inp[5]) ? node30292 : node30285;
														assign node30285 = (inp[3]) ? node30287 : 4'b1111;
															assign node30287 = (inp[4]) ? node30289 : 4'b1101;
																assign node30289 = (inp[9]) ? 4'b1001 : 4'b1101;
														assign node30292 = (inp[3]) ? node30298 : node30293;
															assign node30293 = (inp[9]) ? node30295 : 4'b1101;
																assign node30295 = (inp[4]) ? 4'b1001 : 4'b1101;
															assign node30298 = (inp[9]) ? node30300 : 4'b1001;
																assign node30300 = (inp[4]) ? 4'b1001 : 4'b1101;
									assign node30303 = (inp[12]) ? node30415 : node30304;
										assign node30304 = (inp[15]) ? node30344 : node30305;
											assign node30305 = (inp[0]) ? node30329 : node30306;
												assign node30306 = (inp[5]) ? node30320 : node30307;
													assign node30307 = (inp[3]) ? node30315 : node30308;
														assign node30308 = (inp[9]) ? node30312 : node30309;
															assign node30309 = (inp[4]) ? 4'b1011 : 4'b1111;
															assign node30312 = (inp[4]) ? 4'b1111 : 4'b1011;
														assign node30315 = (inp[4]) ? node30317 : 4'b1011;
															assign node30317 = (inp[9]) ? 4'b1101 : 4'b1011;
													assign node30320 = (inp[9]) ? node30326 : node30321;
														assign node30321 = (inp[4]) ? node30323 : 4'b1101;
															assign node30323 = (inp[3]) ? 4'b1001 : 4'b1011;
														assign node30326 = (inp[4]) ? 4'b1101 : 4'b1001;
												assign node30329 = (inp[9]) ? node30333 : node30330;
													assign node30330 = (inp[4]) ? 4'b1001 : 4'b1101;
													assign node30333 = (inp[4]) ? node30339 : node30334;
														assign node30334 = (inp[5]) ? node30336 : 4'b1001;
															assign node30336 = (inp[2]) ? 4'b1001 : 4'b1011;
														assign node30339 = (inp[5]) ? 4'b1111 : node30340;
															assign node30340 = (inp[3]) ? 4'b1111 : 4'b1101;
											assign node30344 = (inp[0]) ? node30392 : node30345;
												assign node30345 = (inp[3]) ? node30371 : node30346;
													assign node30346 = (inp[5]) ? node30362 : node30347;
														assign node30347 = (inp[2]) ? node30355 : node30348;
															assign node30348 = (inp[9]) ? node30352 : node30349;
																assign node30349 = (inp[4]) ? 4'b1001 : 4'b1101;
																assign node30352 = (inp[4]) ? 4'b1101 : 4'b1001;
															assign node30355 = (inp[9]) ? node30359 : node30356;
																assign node30356 = (inp[4]) ? 4'b1001 : 4'b1101;
																assign node30359 = (inp[4]) ? 4'b1101 : 4'b1001;
														assign node30362 = (inp[2]) ? 4'b1001 : node30363;
															assign node30363 = (inp[9]) ? node30367 : node30364;
																assign node30364 = (inp[4]) ? 4'b1001 : 4'b1101;
																assign node30367 = (inp[4]) ? 4'b1111 : 4'b1001;
													assign node30371 = (inp[5]) ? node30379 : node30372;
														assign node30372 = (inp[4]) ? node30376 : node30373;
															assign node30373 = (inp[9]) ? 4'b1001 : 4'b1101;
															assign node30376 = (inp[9]) ? 4'b1111 : 4'b1001;
														assign node30379 = (inp[2]) ? node30387 : node30380;
															assign node30380 = (inp[9]) ? node30384 : node30381;
																assign node30381 = (inp[4]) ? 4'b1011 : 4'b1111;
																assign node30384 = (inp[4]) ? 4'b1111 : 4'b1011;
															assign node30387 = (inp[9]) ? 4'b1111 : node30388;
																assign node30388 = (inp[4]) ? 4'b1011 : 4'b1111;
												assign node30392 = (inp[5]) ? node30402 : node30393;
													assign node30393 = (inp[4]) ? node30397 : node30394;
														assign node30394 = (inp[9]) ? 4'b1011 : 4'b1111;
														assign node30397 = (inp[9]) ? node30399 : 4'b1011;
															assign node30399 = (inp[3]) ? 4'b1101 : 4'b1111;
													assign node30402 = (inp[3]) ? node30408 : node30403;
														assign node30403 = (inp[4]) ? 4'b1101 : node30404;
															assign node30404 = (inp[9]) ? 4'b1011 : 4'b1111;
														assign node30408 = (inp[9]) ? node30412 : node30409;
															assign node30409 = (inp[4]) ? 4'b1001 : 4'b1101;
															assign node30412 = (inp[4]) ? 4'b1101 : 4'b1001;
										assign node30415 = (inp[4]) ? node30461 : node30416;
											assign node30416 = (inp[9]) ? node30438 : node30417;
												assign node30417 = (inp[15]) ? node30427 : node30418;
													assign node30418 = (inp[0]) ? node30424 : node30419;
														assign node30419 = (inp[5]) ? node30421 : 4'b1011;
															assign node30421 = (inp[3]) ? 4'b1001 : 4'b1011;
														assign node30424 = (inp[5]) ? 4'b1011 : 4'b1001;
													assign node30427 = (inp[0]) ? node30433 : node30428;
														assign node30428 = (inp[3]) ? node30430 : 4'b1001;
															assign node30430 = (inp[5]) ? 4'b1011 : 4'b1001;
														assign node30433 = (inp[3]) ? node30435 : 4'b1011;
															assign node30435 = (inp[5]) ? 4'b1001 : 4'b1011;
												assign node30438 = (inp[5]) ? node30454 : node30439;
													assign node30439 = (inp[15]) ? node30447 : node30440;
														assign node30440 = (inp[0]) ? node30444 : node30441;
															assign node30441 = (inp[3]) ? 4'b1101 : 4'b1111;
															assign node30444 = (inp[3]) ? 4'b1111 : 4'b1101;
														assign node30447 = (inp[0]) ? node30451 : node30448;
															assign node30448 = (inp[3]) ? 4'b1111 : 4'b1101;
															assign node30451 = (inp[3]) ? 4'b1101 : 4'b1111;
													assign node30454 = (inp[15]) ? node30458 : node30455;
														assign node30455 = (inp[0]) ? 4'b1111 : 4'b1101;
														assign node30458 = (inp[0]) ? 4'b1101 : 4'b1111;
											assign node30461 = (inp[9]) ? node30483 : node30462;
												assign node30462 = (inp[3]) ? node30476 : node30463;
													assign node30463 = (inp[5]) ? node30471 : node30464;
														assign node30464 = (inp[15]) ? node30468 : node30465;
															assign node30465 = (inp[0]) ? 4'b1101 : 4'b1111;
															assign node30468 = (inp[0]) ? 4'b1111 : 4'b1101;
														assign node30471 = (inp[15]) ? 4'b1101 : node30472;
															assign node30472 = (inp[0]) ? 4'b1111 : 4'b1101;
													assign node30476 = (inp[15]) ? node30480 : node30477;
														assign node30477 = (inp[0]) ? 4'b1111 : 4'b1101;
														assign node30480 = (inp[0]) ? 4'b1101 : 4'b1111;
												assign node30483 = (inp[15]) ? node30501 : node30484;
													assign node30484 = (inp[2]) ? node30494 : node30485;
														assign node30485 = (inp[0]) ? node30491 : node30486;
															assign node30486 = (inp[3]) ? 4'b1001 : node30487;
																assign node30487 = (inp[5]) ? 4'b1001 : 4'b1011;
															assign node30491 = (inp[5]) ? 4'b1011 : 4'b1001;
														assign node30494 = (inp[5]) ? 4'b1001 : node30495;
															assign node30495 = (inp[0]) ? 4'b1001 : node30496;
																assign node30496 = (inp[3]) ? 4'b1001 : 4'b1011;
													assign node30501 = (inp[0]) ? node30507 : node30502;
														assign node30502 = (inp[5]) ? 4'b1011 : node30503;
															assign node30503 = (inp[3]) ? 4'b1011 : 4'b1001;
														assign node30507 = (inp[3]) ? 4'b1001 : 4'b1011;
								assign node30510 = (inp[2]) ? node30810 : node30511;
									assign node30511 = (inp[14]) ? node30659 : node30512;
										assign node30512 = (inp[0]) ? node30584 : node30513;
											assign node30513 = (inp[12]) ? node30545 : node30514;
												assign node30514 = (inp[15]) ? node30530 : node30515;
													assign node30515 = (inp[5]) ? node30521 : node30516;
														assign node30516 = (inp[9]) ? 4'b1011 : node30517;
															assign node30517 = (inp[4]) ? 4'b1011 : 4'b1111;
														assign node30521 = (inp[3]) ? 4'b1101 : node30522;
															assign node30522 = (inp[4]) ? node30526 : node30523;
																assign node30523 = (inp[9]) ? 4'b1011 : 4'b1111;
																assign node30526 = (inp[9]) ? 4'b1101 : 4'b1011;
													assign node30530 = (inp[9]) ? node30538 : node30531;
														assign node30531 = (inp[4]) ? 4'b1001 : node30532;
															assign node30532 = (inp[5]) ? node30534 : 4'b1101;
																assign node30534 = (inp[3]) ? 4'b1111 : 4'b1101;
														assign node30538 = (inp[4]) ? node30540 : 4'b1001;
															assign node30540 = (inp[5]) ? 4'b1111 : node30541;
																assign node30541 = (inp[3]) ? 4'b1111 : 4'b1101;
												assign node30545 = (inp[3]) ? node30565 : node30546;
													assign node30546 = (inp[15]) ? node30554 : node30547;
														assign node30547 = (inp[5]) ? node30549 : 4'b1111;
															assign node30549 = (inp[4]) ? 4'b1101 : node30550;
																assign node30550 = (inp[9]) ? 4'b1101 : 4'b1011;
														assign node30554 = (inp[5]) ? node30560 : node30555;
															assign node30555 = (inp[9]) ? node30557 : 4'b1101;
																assign node30557 = (inp[4]) ? 4'b1001 : 4'b1101;
															assign node30560 = (inp[9]) ? 4'b1111 : node30561;
																assign node30561 = (inp[4]) ? 4'b1111 : 4'b1001;
													assign node30565 = (inp[15]) ? node30575 : node30566;
														assign node30566 = (inp[4]) ? node30572 : node30567;
															assign node30567 = (inp[5]) ? node30569 : 4'b1011;
																assign node30569 = (inp[9]) ? 4'b1101 : 4'b1001;
															assign node30572 = (inp[9]) ? 4'b1001 : 4'b1101;
														assign node30575 = (inp[9]) ? node30581 : node30576;
															assign node30576 = (inp[4]) ? 4'b1111 : node30577;
																assign node30577 = (inp[5]) ? 4'b1011 : 4'b1001;
															assign node30581 = (inp[4]) ? 4'b1011 : 4'b1111;
											assign node30584 = (inp[3]) ? node30624 : node30585;
												assign node30585 = (inp[15]) ? node30605 : node30586;
													assign node30586 = (inp[9]) ? node30592 : node30587;
														assign node30587 = (inp[12]) ? 4'b1001 : node30588;
															assign node30588 = (inp[4]) ? 4'b1001 : 4'b1101;
														assign node30592 = (inp[5]) ? node30598 : node30593;
															assign node30593 = (inp[4]) ? node30595 : 4'b1101;
																assign node30595 = (inp[12]) ? 4'b1001 : 4'b1101;
															assign node30598 = (inp[12]) ? node30602 : node30599;
																assign node30599 = (inp[4]) ? 4'b1111 : 4'b1001;
																assign node30602 = (inp[4]) ? 4'b1011 : 4'b1111;
													assign node30605 = (inp[5]) ? node30615 : node30606;
														assign node30606 = (inp[4]) ? 4'b1011 : node30607;
															assign node30607 = (inp[9]) ? node30611 : node30608;
																assign node30608 = (inp[12]) ? 4'b1011 : 4'b1111;
																assign node30611 = (inp[12]) ? 4'b1111 : 4'b1011;
														assign node30615 = (inp[9]) ? node30617 : 4'b1011;
															assign node30617 = (inp[4]) ? node30621 : node30618;
																assign node30618 = (inp[12]) ? 4'b1101 : 4'b1011;
																assign node30621 = (inp[12]) ? 4'b1001 : 4'b1101;
												assign node30624 = (inp[15]) ? node30642 : node30625;
													assign node30625 = (inp[12]) ? node30635 : node30626;
														assign node30626 = (inp[9]) ? node30630 : node30627;
															assign node30627 = (inp[5]) ? 4'b1111 : 4'b1101;
															assign node30630 = (inp[4]) ? 4'b1111 : node30631;
																assign node30631 = (inp[5]) ? 4'b1011 : 4'b1001;
														assign node30635 = (inp[4]) ? node30639 : node30636;
															assign node30636 = (inp[9]) ? 4'b1111 : 4'b1011;
															assign node30639 = (inp[9]) ? 4'b1011 : 4'b1111;
													assign node30642 = (inp[12]) ? node30652 : node30643;
														assign node30643 = (inp[9]) ? node30647 : node30644;
															assign node30644 = (inp[5]) ? 4'b1101 : 4'b1111;
															assign node30647 = (inp[4]) ? 4'b1101 : node30648;
																assign node30648 = (inp[5]) ? 4'b1001 : 4'b1011;
														assign node30652 = (inp[9]) ? node30656 : node30653;
															assign node30653 = (inp[4]) ? 4'b1101 : 4'b1001;
															assign node30656 = (inp[4]) ? 4'b1001 : 4'b1101;
										assign node30659 = (inp[5]) ? node30733 : node30660;
											assign node30660 = (inp[4]) ? node30690 : node30661;
												assign node30661 = (inp[9]) ? node30679 : node30662;
													assign node30662 = (inp[12]) ? node30672 : node30663;
														assign node30663 = (inp[3]) ? node30665 : 4'b1110;
															assign node30665 = (inp[0]) ? node30669 : node30666;
																assign node30666 = (inp[15]) ? 4'b1100 : 4'b1110;
																assign node30669 = (inp[15]) ? 4'b1110 : 4'b1100;
														assign node30672 = (inp[0]) ? node30676 : node30673;
															assign node30673 = (inp[15]) ? 4'b1000 : 4'b1010;
															assign node30676 = (inp[3]) ? 4'b1010 : 4'b1000;
													assign node30679 = (inp[12]) ? node30687 : node30680;
														assign node30680 = (inp[15]) ? node30684 : node30681;
															assign node30681 = (inp[0]) ? 4'b1000 : 4'b1010;
															assign node30684 = (inp[0]) ? 4'b1010 : 4'b1000;
														assign node30687 = (inp[15]) ? 4'b1100 : 4'b1110;
												assign node30690 = (inp[0]) ? node30710 : node30691;
													assign node30691 = (inp[15]) ? node30699 : node30692;
														assign node30692 = (inp[3]) ? node30694 : 4'b1110;
															assign node30694 = (inp[9]) ? node30696 : 4'b1100;
																assign node30696 = (inp[12]) ? 4'b1000 : 4'b1100;
														assign node30699 = (inp[3]) ? node30707 : node30700;
															assign node30700 = (inp[12]) ? node30704 : node30701;
																assign node30701 = (inp[9]) ? 4'b1100 : 4'b1000;
																assign node30704 = (inp[9]) ? 4'b1000 : 4'b1100;
															assign node30707 = (inp[9]) ? 4'b1010 : 4'b1110;
													assign node30710 = (inp[15]) ? node30724 : node30711;
														assign node30711 = (inp[3]) ? node30717 : node30712;
															assign node30712 = (inp[12]) ? 4'b1000 : node30713;
																assign node30713 = (inp[9]) ? 4'b1100 : 4'b1000;
															assign node30717 = (inp[9]) ? node30721 : node30718;
																assign node30718 = (inp[12]) ? 4'b1110 : 4'b1000;
																assign node30721 = (inp[12]) ? 4'b1010 : 4'b1110;
														assign node30724 = (inp[3]) ? node30726 : 4'b1110;
															assign node30726 = (inp[9]) ? node30730 : node30727;
																assign node30727 = (inp[12]) ? 4'b1100 : 4'b1010;
																assign node30730 = (inp[12]) ? 4'b1000 : 4'b1100;
											assign node30733 = (inp[4]) ? node30773 : node30734;
												assign node30734 = (inp[9]) ? node30756 : node30735;
													assign node30735 = (inp[12]) ? node30749 : node30736;
														assign node30736 = (inp[15]) ? node30744 : node30737;
															assign node30737 = (inp[3]) ? node30741 : node30738;
																assign node30738 = (inp[0]) ? 4'b1100 : 4'b1110;
																assign node30741 = (inp[0]) ? 4'b1110 : 4'b1100;
															assign node30744 = (inp[0]) ? node30746 : 4'b1100;
																assign node30746 = (inp[3]) ? 4'b1100 : 4'b1110;
														assign node30749 = (inp[0]) ? 4'b1010 : node30750;
															assign node30750 = (inp[15]) ? 4'b1000 : node30751;
																assign node30751 = (inp[3]) ? 4'b1000 : 4'b1010;
													assign node30756 = (inp[12]) ? node30766 : node30757;
														assign node30757 = (inp[15]) ? 4'b1010 : node30758;
															assign node30758 = (inp[0]) ? node30762 : node30759;
																assign node30759 = (inp[3]) ? 4'b1000 : 4'b1010;
																assign node30762 = (inp[3]) ? 4'b1010 : 4'b1000;
														assign node30766 = (inp[15]) ? node30770 : node30767;
															assign node30767 = (inp[0]) ? 4'b1110 : 4'b1100;
															assign node30770 = (inp[0]) ? 4'b1100 : 4'b1110;
												assign node30773 = (inp[0]) ? node30793 : node30774;
													assign node30774 = (inp[15]) ? node30778 : node30775;
														assign node30775 = (inp[12]) ? 4'b1000 : 4'b1010;
														assign node30778 = (inp[3]) ? node30786 : node30779;
															assign node30779 = (inp[9]) ? node30783 : node30780;
																assign node30780 = (inp[12]) ? 4'b1110 : 4'b1000;
																assign node30783 = (inp[12]) ? 4'b1010 : 4'b1110;
															assign node30786 = (inp[9]) ? node30790 : node30787;
																assign node30787 = (inp[12]) ? 4'b1110 : 4'b1010;
																assign node30790 = (inp[12]) ? 4'b1010 : 4'b1110;
													assign node30793 = (inp[15]) ? node30803 : node30794;
														assign node30794 = (inp[3]) ? 4'b1010 : node30795;
															assign node30795 = (inp[12]) ? node30799 : node30796;
																assign node30796 = (inp[9]) ? 4'b1110 : 4'b1000;
																assign node30799 = (inp[9]) ? 4'b1010 : 4'b1110;
														assign node30803 = (inp[9]) ? node30807 : node30804;
															assign node30804 = (inp[3]) ? 4'b1000 : 4'b1010;
															assign node30807 = (inp[12]) ? 4'b1000 : 4'b1100;
									assign node30810 = (inp[0]) ? node30928 : node30811;
										assign node30811 = (inp[4]) ? node30873 : node30812;
											assign node30812 = (inp[15]) ? node30836 : node30813;
												assign node30813 = (inp[3]) ? node30823 : node30814;
													assign node30814 = (inp[9]) ? node30818 : node30815;
														assign node30815 = (inp[12]) ? 4'b1010 : 4'b1110;
														assign node30818 = (inp[12]) ? node30820 : 4'b1010;
															assign node30820 = (inp[5]) ? 4'b1100 : 4'b1110;
													assign node30823 = (inp[5]) ? node30829 : node30824;
														assign node30824 = (inp[14]) ? node30826 : 4'b1010;
															assign node30826 = (inp[12]) ? 4'b1100 : 4'b1010;
														assign node30829 = (inp[12]) ? node30833 : node30830;
															assign node30830 = (inp[9]) ? 4'b1000 : 4'b1100;
															assign node30833 = (inp[9]) ? 4'b1100 : 4'b1000;
												assign node30836 = (inp[5]) ? node30850 : node30837;
													assign node30837 = (inp[3]) ? node30845 : node30838;
														assign node30838 = (inp[12]) ? node30842 : node30839;
															assign node30839 = (inp[9]) ? 4'b1000 : 4'b1100;
															assign node30842 = (inp[9]) ? 4'b1100 : 4'b1000;
														assign node30845 = (inp[9]) ? 4'b1000 : node30846;
															assign node30846 = (inp[12]) ? 4'b1000 : 4'b1100;
													assign node30850 = (inp[3]) ? node30860 : node30851;
														assign node30851 = (inp[14]) ? node30853 : 4'b1000;
															assign node30853 = (inp[12]) ? node30857 : node30854;
																assign node30854 = (inp[9]) ? 4'b1000 : 4'b1100;
																assign node30857 = (inp[9]) ? 4'b1110 : 4'b1000;
														assign node30860 = (inp[14]) ? node30866 : node30861;
															assign node30861 = (inp[12]) ? 4'b1010 : node30862;
																assign node30862 = (inp[9]) ? 4'b1010 : 4'b1110;
															assign node30866 = (inp[12]) ? node30870 : node30867;
																assign node30867 = (inp[9]) ? 4'b1010 : 4'b1110;
																assign node30870 = (inp[9]) ? 4'b1110 : 4'b1010;
											assign node30873 = (inp[15]) ? node30905 : node30874;
												assign node30874 = (inp[3]) ? node30890 : node30875;
													assign node30875 = (inp[5]) ? node30883 : node30876;
														assign node30876 = (inp[12]) ? node30880 : node30877;
															assign node30877 = (inp[9]) ? 4'b1110 : 4'b1010;
															assign node30880 = (inp[9]) ? 4'b1010 : 4'b1110;
														assign node30883 = (inp[9]) ? node30887 : node30884;
															assign node30884 = (inp[12]) ? 4'b1100 : 4'b1010;
															assign node30887 = (inp[12]) ? 4'b1000 : 4'b1100;
													assign node30890 = (inp[5]) ? node30898 : node30891;
														assign node30891 = (inp[12]) ? node30895 : node30892;
															assign node30892 = (inp[9]) ? 4'b1100 : 4'b1010;
															assign node30895 = (inp[9]) ? 4'b1000 : 4'b1100;
														assign node30898 = (inp[9]) ? node30902 : node30899;
															assign node30899 = (inp[12]) ? 4'b1100 : 4'b1000;
															assign node30902 = (inp[12]) ? 4'b1000 : 4'b1100;
												assign node30905 = (inp[3]) ? node30921 : node30906;
													assign node30906 = (inp[5]) ? node30916 : node30907;
														assign node30907 = (inp[14]) ? node30909 : 4'b1000;
															assign node30909 = (inp[12]) ? node30913 : node30910;
																assign node30910 = (inp[9]) ? 4'b1100 : 4'b1000;
																assign node30913 = (inp[9]) ? 4'b1000 : 4'b1100;
														assign node30916 = (inp[9]) ? node30918 : 4'b1000;
															assign node30918 = (inp[12]) ? 4'b1010 : 4'b1110;
													assign node30921 = (inp[12]) ? node30925 : node30922;
														assign node30922 = (inp[9]) ? 4'b1110 : 4'b1010;
														assign node30925 = (inp[9]) ? 4'b1010 : 4'b1110;
										assign node30928 = (inp[5]) ? node30994 : node30929;
											assign node30929 = (inp[15]) ? node30967 : node30930;
												assign node30930 = (inp[3]) ? node30950 : node30931;
													assign node30931 = (inp[9]) ? node30939 : node30932;
														assign node30932 = (inp[12]) ? node30936 : node30933;
															assign node30933 = (inp[4]) ? 4'b1000 : 4'b1100;
															assign node30936 = (inp[4]) ? 4'b1100 : 4'b1000;
														assign node30939 = (inp[14]) ? node30945 : node30940;
															assign node30940 = (inp[4]) ? 4'b1100 : node30941;
																assign node30941 = (inp[12]) ? 4'b1100 : 4'b1000;
															assign node30945 = (inp[4]) ? node30947 : 4'b1100;
																assign node30947 = (inp[12]) ? 4'b1000 : 4'b1100;
													assign node30950 = (inp[12]) ? node30956 : node30951;
														assign node30951 = (inp[4]) ? 4'b1000 : node30952;
															assign node30952 = (inp[9]) ? 4'b1000 : 4'b1100;
														assign node30956 = (inp[14]) ? node30962 : node30957;
															assign node30957 = (inp[9]) ? node30959 : 4'b1000;
																assign node30959 = (inp[4]) ? 4'b1010 : 4'b1110;
															assign node30962 = (inp[4]) ? node30964 : 4'b1110;
																assign node30964 = (inp[9]) ? 4'b1010 : 4'b1110;
												assign node30967 = (inp[3]) ? node30979 : node30968;
													assign node30968 = (inp[12]) ? node30974 : node30969;
														assign node30969 = (inp[9]) ? node30971 : 4'b1010;
															assign node30971 = (inp[4]) ? 4'b1110 : 4'b1010;
														assign node30974 = (inp[9]) ? node30976 : 4'b1110;
															assign node30976 = (inp[4]) ? 4'b1010 : 4'b1110;
													assign node30979 = (inp[4]) ? node30987 : node30980;
														assign node30980 = (inp[9]) ? node30984 : node30981;
															assign node30981 = (inp[12]) ? 4'b1010 : 4'b1110;
															assign node30984 = (inp[12]) ? 4'b1100 : 4'b1010;
														assign node30987 = (inp[12]) ? node30991 : node30988;
															assign node30988 = (inp[9]) ? 4'b1100 : 4'b1010;
															assign node30991 = (inp[9]) ? 4'b1000 : 4'b1100;
											assign node30994 = (inp[15]) ? node31030 : node30995;
												assign node30995 = (inp[3]) ? node31009 : node30996;
													assign node30996 = (inp[4]) ? node31004 : node30997;
														assign node30997 = (inp[9]) ? node31001 : node30998;
															assign node30998 = (inp[12]) ? 4'b1000 : 4'b1100;
															assign node31001 = (inp[12]) ? 4'b1110 : 4'b1000;
														assign node31004 = (inp[9]) ? node31006 : 4'b1110;
															assign node31006 = (inp[12]) ? 4'b1010 : 4'b1110;
													assign node31009 = (inp[14]) ? node31015 : node31010;
														assign node31010 = (inp[9]) ? 4'b1110 : node31011;
															assign node31011 = (inp[12]) ? 4'b1010 : 4'b1110;
														assign node31015 = (inp[4]) ? node31023 : node31016;
															assign node31016 = (inp[12]) ? node31020 : node31017;
																assign node31017 = (inp[9]) ? 4'b1010 : 4'b1110;
																assign node31020 = (inp[9]) ? 4'b1110 : 4'b1010;
															assign node31023 = (inp[9]) ? node31027 : node31024;
																assign node31024 = (inp[12]) ? 4'b1110 : 4'b1010;
																assign node31027 = (inp[12]) ? 4'b1010 : 4'b1110;
												assign node31030 = (inp[3]) ? node31044 : node31031;
													assign node31031 = (inp[4]) ? node31039 : node31032;
														assign node31032 = (inp[12]) ? node31036 : node31033;
															assign node31033 = (inp[9]) ? 4'b1010 : 4'b1110;
															assign node31036 = (inp[9]) ? 4'b1100 : 4'b1010;
														assign node31039 = (inp[9]) ? node31041 : 4'b1100;
															assign node31041 = (inp[12]) ? 4'b1000 : 4'b1100;
													assign node31044 = (inp[14]) ? node31058 : node31045;
														assign node31045 = (inp[9]) ? node31053 : node31046;
															assign node31046 = (inp[4]) ? node31050 : node31047;
																assign node31047 = (inp[12]) ? 4'b1000 : 4'b1100;
																assign node31050 = (inp[12]) ? 4'b1100 : 4'b1000;
															assign node31053 = (inp[12]) ? node31055 : 4'b1000;
																assign node31055 = (inp[4]) ? 4'b1000 : 4'b1100;
														assign node31058 = (inp[9]) ? node31060 : 4'b1000;
															assign node31060 = (inp[4]) ? 4'b1100 : 4'b1000;
						assign node31063 = (inp[12]) ? node32263 : node31064;
							assign node31064 = (inp[9]) ? node31662 : node31065;
								assign node31065 = (inp[4]) ? node31411 : node31066;
									assign node31066 = (inp[14]) ? node31232 : node31067;
										assign node31067 = (inp[5]) ? node31157 : node31068;
											assign node31068 = (inp[8]) ? node31110 : node31069;
												assign node31069 = (inp[0]) ? node31091 : node31070;
													assign node31070 = (inp[15]) ? node31086 : node31071;
														assign node31071 = (inp[3]) ? node31079 : node31072;
															assign node31072 = (inp[2]) ? node31076 : node31073;
																assign node31073 = (inp[7]) ? 4'b1010 : 4'b1011;
																assign node31076 = (inp[7]) ? 4'b1011 : 4'b1010;
															assign node31079 = (inp[7]) ? node31083 : node31080;
																assign node31080 = (inp[2]) ? 4'b1010 : 4'b1011;
																assign node31083 = (inp[2]) ? 4'b1011 : 4'b1010;
														assign node31086 = (inp[7]) ? node31088 : 4'b1000;
															assign node31088 = (inp[2]) ? 4'b1001 : 4'b1000;
													assign node31091 = (inp[15]) ? node31103 : node31092;
														assign node31092 = (inp[3]) ? node31098 : node31093;
															assign node31093 = (inp[7]) ? 4'b1000 : node31094;
																assign node31094 = (inp[2]) ? 4'b1000 : 4'b1001;
															assign node31098 = (inp[2]) ? node31100 : 4'b1001;
																assign node31100 = (inp[7]) ? 4'b1001 : 4'b1000;
														assign node31103 = (inp[3]) ? 4'b1010 : node31104;
															assign node31104 = (inp[7]) ? 4'b1011 : node31105;
																assign node31105 = (inp[2]) ? 4'b1010 : 4'b1011;
												assign node31110 = (inp[3]) ? node31132 : node31111;
													assign node31111 = (inp[15]) ? node31119 : node31112;
														assign node31112 = (inp[0]) ? node31114 : 4'b1011;
															assign node31114 = (inp[2]) ? node31116 : 4'b1001;
																assign node31116 = (inp[7]) ? 4'b1000 : 4'b1001;
														assign node31119 = (inp[0]) ? node31127 : node31120;
															assign node31120 = (inp[2]) ? node31124 : node31121;
																assign node31121 = (inp[7]) ? 4'b1001 : 4'b1000;
																assign node31124 = (inp[7]) ? 4'b1000 : 4'b1001;
															assign node31127 = (inp[7]) ? 4'b1010 : node31128;
																assign node31128 = (inp[2]) ? 4'b1011 : 4'b1010;
													assign node31132 = (inp[0]) ? node31144 : node31133;
														assign node31133 = (inp[15]) ? node31139 : node31134;
															assign node31134 = (inp[7]) ? node31136 : 4'b1010;
																assign node31136 = (inp[2]) ? 4'b1010 : 4'b1011;
															assign node31139 = (inp[2]) ? node31141 : 4'b1001;
																assign node31141 = (inp[7]) ? 4'b1000 : 4'b1001;
														assign node31144 = (inp[15]) ? node31150 : node31145;
															assign node31145 = (inp[7]) ? 4'b1001 : node31146;
																assign node31146 = (inp[2]) ? 4'b1001 : 4'b1000;
															assign node31150 = (inp[7]) ? node31154 : node31151;
																assign node31151 = (inp[2]) ? 4'b1011 : 4'b1010;
																assign node31154 = (inp[2]) ? 4'b1010 : 4'b1011;
											assign node31157 = (inp[2]) ? node31195 : node31158;
												assign node31158 = (inp[3]) ? node31176 : node31159;
													assign node31159 = (inp[0]) ? node31167 : node31160;
														assign node31160 = (inp[15]) ? 4'b1000 : node31161;
															assign node31161 = (inp[8]) ? node31163 : 4'b1010;
																assign node31163 = (inp[7]) ? 4'b1011 : 4'b1010;
														assign node31167 = (inp[15]) ? node31173 : node31168;
															assign node31168 = (inp[8]) ? 4'b1000 : node31169;
																assign node31169 = (inp[7]) ? 4'b1000 : 4'b1001;
															assign node31173 = (inp[8]) ? 4'b1010 : 4'b1011;
													assign node31176 = (inp[15]) ? node31186 : node31177;
														assign node31177 = (inp[0]) ? 4'b1010 : node31178;
															assign node31178 = (inp[8]) ? node31182 : node31179;
																assign node31179 = (inp[7]) ? 4'b1000 : 4'b1001;
																assign node31182 = (inp[7]) ? 4'b1001 : 4'b1000;
														assign node31186 = (inp[0]) ? node31188 : 4'b1010;
															assign node31188 = (inp[7]) ? node31192 : node31189;
																assign node31189 = (inp[8]) ? 4'b1000 : 4'b1001;
																assign node31192 = (inp[8]) ? 4'b1001 : 4'b1000;
												assign node31195 = (inp[8]) ? node31209 : node31196;
													assign node31196 = (inp[7]) ? node31200 : node31197;
														assign node31197 = (inp[15]) ? 4'b1010 : 4'b1000;
														assign node31200 = (inp[15]) ? node31202 : 4'b1001;
															assign node31202 = (inp[0]) ? node31206 : node31203;
																assign node31203 = (inp[3]) ? 4'b1011 : 4'b1001;
																assign node31206 = (inp[3]) ? 4'b1001 : 4'b1011;
													assign node31209 = (inp[7]) ? node31221 : node31210;
														assign node31210 = (inp[15]) ? node31216 : node31211;
															assign node31211 = (inp[3]) ? 4'b1001 : node31212;
																assign node31212 = (inp[0]) ? 4'b1001 : 4'b1011;
															assign node31216 = (inp[3]) ? node31218 : 4'b1011;
																assign node31218 = (inp[0]) ? 4'b1001 : 4'b1011;
														assign node31221 = (inp[15]) ? node31227 : node31222;
															assign node31222 = (inp[3]) ? 4'b1010 : node31223;
																assign node31223 = (inp[0]) ? 4'b1000 : 4'b1010;
															assign node31227 = (inp[0]) ? node31229 : 4'b1000;
																assign node31229 = (inp[3]) ? 4'b1000 : 4'b1010;
										assign node31232 = (inp[2]) ? node31318 : node31233;
											assign node31233 = (inp[3]) ? node31271 : node31234;
												assign node31234 = (inp[0]) ? node31248 : node31235;
													assign node31235 = (inp[15]) ? node31243 : node31236;
														assign node31236 = (inp[7]) ? node31240 : node31237;
															assign node31237 = (inp[8]) ? 4'b1011 : 4'b1010;
															assign node31240 = (inp[8]) ? 4'b1010 : 4'b1011;
														assign node31243 = (inp[7]) ? node31245 : 4'b1000;
															assign node31245 = (inp[8]) ? 4'b1000 : 4'b1001;
													assign node31248 = (inp[15]) ? node31264 : node31249;
														assign node31249 = (inp[5]) ? node31257 : node31250;
															assign node31250 = (inp[7]) ? node31254 : node31251;
																assign node31251 = (inp[8]) ? 4'b1001 : 4'b1000;
																assign node31254 = (inp[8]) ? 4'b1000 : 4'b1001;
															assign node31257 = (inp[8]) ? node31261 : node31258;
																assign node31258 = (inp[7]) ? 4'b1001 : 4'b1000;
																assign node31261 = (inp[7]) ? 4'b1000 : 4'b1001;
														assign node31264 = (inp[8]) ? node31268 : node31265;
															assign node31265 = (inp[7]) ? 4'b1011 : 4'b1010;
															assign node31268 = (inp[7]) ? 4'b1010 : 4'b1011;
												assign node31271 = (inp[5]) ? node31299 : node31272;
													assign node31272 = (inp[7]) ? node31288 : node31273;
														assign node31273 = (inp[8]) ? node31281 : node31274;
															assign node31274 = (inp[0]) ? node31278 : node31275;
																assign node31275 = (inp[15]) ? 4'b1000 : 4'b1010;
																assign node31278 = (inp[15]) ? 4'b1010 : 4'b1000;
															assign node31281 = (inp[0]) ? node31285 : node31282;
																assign node31282 = (inp[15]) ? 4'b1001 : 4'b1011;
																assign node31285 = (inp[15]) ? 4'b1011 : 4'b1001;
														assign node31288 = (inp[8]) ? node31294 : node31289;
															assign node31289 = (inp[15]) ? 4'b1011 : node31290;
																assign node31290 = (inp[0]) ? 4'b1001 : 4'b1011;
															assign node31294 = (inp[0]) ? 4'b1010 : node31295;
																assign node31295 = (inp[15]) ? 4'b1000 : 4'b1010;
													assign node31299 = (inp[7]) ? node31309 : node31300;
														assign node31300 = (inp[8]) ? node31302 : 4'b1010;
															assign node31302 = (inp[0]) ? node31306 : node31303;
																assign node31303 = (inp[15]) ? 4'b1011 : 4'b1001;
																assign node31306 = (inp[15]) ? 4'b1001 : 4'b1011;
														assign node31309 = (inp[8]) ? 4'b1000 : node31310;
															assign node31310 = (inp[15]) ? node31314 : node31311;
																assign node31311 = (inp[0]) ? 4'b1011 : 4'b1001;
																assign node31314 = (inp[0]) ? 4'b1001 : 4'b1011;
											assign node31318 = (inp[5]) ? node31364 : node31319;
												assign node31319 = (inp[15]) ? node31345 : node31320;
													assign node31320 = (inp[0]) ? node31336 : node31321;
														assign node31321 = (inp[3]) ? node31329 : node31322;
															assign node31322 = (inp[7]) ? node31326 : node31323;
																assign node31323 = (inp[8]) ? 4'b1011 : 4'b1010;
																assign node31326 = (inp[8]) ? 4'b1010 : 4'b1011;
															assign node31329 = (inp[7]) ? node31333 : node31330;
																assign node31330 = (inp[8]) ? 4'b1011 : 4'b1010;
																assign node31333 = (inp[8]) ? 4'b1010 : 4'b1011;
														assign node31336 = (inp[3]) ? node31342 : node31337;
															assign node31337 = (inp[8]) ? 4'b1001 : node31338;
																assign node31338 = (inp[7]) ? 4'b1001 : 4'b1000;
															assign node31342 = (inp[7]) ? 4'b1000 : 4'b1001;
													assign node31345 = (inp[0]) ? node31353 : node31346;
														assign node31346 = (inp[8]) ? node31350 : node31347;
															assign node31347 = (inp[7]) ? 4'b1001 : 4'b1000;
															assign node31350 = (inp[7]) ? 4'b1000 : 4'b1001;
														assign node31353 = (inp[3]) ? node31359 : node31354;
															assign node31354 = (inp[8]) ? node31356 : 4'b1011;
																assign node31356 = (inp[7]) ? 4'b1010 : 4'b1011;
															assign node31359 = (inp[7]) ? 4'b1010 : node31360;
																assign node31360 = (inp[8]) ? 4'b1011 : 4'b1010;
												assign node31364 = (inp[3]) ? node31386 : node31365;
													assign node31365 = (inp[8]) ? node31373 : node31366;
														assign node31366 = (inp[7]) ? 4'b1011 : node31367;
															assign node31367 = (inp[15]) ? 4'b1010 : node31368;
																assign node31368 = (inp[0]) ? 4'b1000 : 4'b1010;
														assign node31373 = (inp[7]) ? node31381 : node31374;
															assign node31374 = (inp[15]) ? node31378 : node31375;
																assign node31375 = (inp[0]) ? 4'b1001 : 4'b1011;
																assign node31378 = (inp[0]) ? 4'b1011 : 4'b1001;
															assign node31381 = (inp[15]) ? node31383 : 4'b1010;
																assign node31383 = (inp[0]) ? 4'b1010 : 4'b1000;
													assign node31386 = (inp[7]) ? node31396 : node31387;
														assign node31387 = (inp[8]) ? 4'b1011 : node31388;
															assign node31388 = (inp[15]) ? node31392 : node31389;
																assign node31389 = (inp[0]) ? 4'b1010 : 4'b1000;
																assign node31392 = (inp[0]) ? 4'b1000 : 4'b1010;
														assign node31396 = (inp[8]) ? node31404 : node31397;
															assign node31397 = (inp[0]) ? node31401 : node31398;
																assign node31398 = (inp[15]) ? 4'b1011 : 4'b1001;
																assign node31401 = (inp[15]) ? 4'b1001 : 4'b1011;
															assign node31404 = (inp[0]) ? node31408 : node31405;
																assign node31405 = (inp[15]) ? 4'b1010 : 4'b1000;
																assign node31408 = (inp[15]) ? 4'b1000 : 4'b1010;
									assign node31411 = (inp[0]) ? node31527 : node31412;
										assign node31412 = (inp[15]) ? node31470 : node31413;
											assign node31413 = (inp[5]) ? node31447 : node31414;
												assign node31414 = (inp[3]) ? node31436 : node31415;
													assign node31415 = (inp[14]) ? node31429 : node31416;
														assign node31416 = (inp[7]) ? node31424 : node31417;
															assign node31417 = (inp[8]) ? node31421 : node31418;
																assign node31418 = (inp[2]) ? 4'b1110 : 4'b1111;
																assign node31421 = (inp[2]) ? 4'b1111 : 4'b1110;
															assign node31424 = (inp[2]) ? 4'b1111 : node31425;
																assign node31425 = (inp[8]) ? 4'b1111 : 4'b1110;
														assign node31429 = (inp[2]) ? 4'b1111 : node31430;
															assign node31430 = (inp[7]) ? node31432 : 4'b1111;
																assign node31432 = (inp[8]) ? 4'b1110 : 4'b1111;
													assign node31436 = (inp[8]) ? node31442 : node31437;
														assign node31437 = (inp[14]) ? 4'b1100 : node31438;
															assign node31438 = (inp[7]) ? 4'b1100 : 4'b1101;
														assign node31442 = (inp[14]) ? 4'b1101 : node31443;
															assign node31443 = (inp[7]) ? 4'b1101 : 4'b1100;
												assign node31447 = (inp[8]) ? node31459 : node31448;
													assign node31448 = (inp[7]) ? node31454 : node31449;
														assign node31449 = (inp[14]) ? 4'b1100 : node31450;
															assign node31450 = (inp[2]) ? 4'b1100 : 4'b1101;
														assign node31454 = (inp[2]) ? 4'b1101 : node31455;
															assign node31455 = (inp[14]) ? 4'b1101 : 4'b1100;
													assign node31459 = (inp[7]) ? node31465 : node31460;
														assign node31460 = (inp[2]) ? 4'b1101 : node31461;
															assign node31461 = (inp[14]) ? 4'b1101 : 4'b1100;
														assign node31465 = (inp[14]) ? 4'b1100 : node31466;
															assign node31466 = (inp[2]) ? 4'b1100 : 4'b1101;
											assign node31470 = (inp[5]) ? node31496 : node31471;
												assign node31471 = (inp[3]) ? node31485 : node31472;
													assign node31472 = (inp[8]) ? node31480 : node31473;
														assign node31473 = (inp[7]) ? 4'b1101 : node31474;
															assign node31474 = (inp[2]) ? 4'b1100 : node31475;
																assign node31475 = (inp[14]) ? 4'b1100 : 4'b1101;
														assign node31480 = (inp[7]) ? node31482 : 4'b1101;
															assign node31482 = (inp[2]) ? 4'b1100 : 4'b1101;
													assign node31485 = (inp[2]) ? node31491 : node31486;
														assign node31486 = (inp[14]) ? node31488 : 4'b1111;
															assign node31488 = (inp[8]) ? 4'b1110 : 4'b1111;
														assign node31491 = (inp[8]) ? node31493 : 4'b1110;
															assign node31493 = (inp[7]) ? 4'b1110 : 4'b1111;
												assign node31496 = (inp[14]) ? node31512 : node31497;
													assign node31497 = (inp[2]) ? node31505 : node31498;
														assign node31498 = (inp[7]) ? node31502 : node31499;
															assign node31499 = (inp[8]) ? 4'b1110 : 4'b1111;
															assign node31502 = (inp[8]) ? 4'b1111 : 4'b1110;
														assign node31505 = (inp[8]) ? node31509 : node31506;
															assign node31506 = (inp[7]) ? 4'b1111 : 4'b1110;
															assign node31509 = (inp[7]) ? 4'b1110 : 4'b1111;
													assign node31512 = (inp[2]) ? node31520 : node31513;
														assign node31513 = (inp[3]) ? node31515 : 4'b1110;
															assign node31515 = (inp[7]) ? 4'b1111 : node31516;
																assign node31516 = (inp[8]) ? 4'b1111 : 4'b1110;
														assign node31520 = (inp[3]) ? 4'b1110 : node31521;
															assign node31521 = (inp[7]) ? 4'b1110 : node31522;
																assign node31522 = (inp[8]) ? 4'b1111 : 4'b1110;
										assign node31527 = (inp[15]) ? node31603 : node31528;
											assign node31528 = (inp[3]) ? node31566 : node31529;
												assign node31529 = (inp[5]) ? node31549 : node31530;
													assign node31530 = (inp[8]) ? node31538 : node31531;
														assign node31531 = (inp[2]) ? 4'b1101 : node31532;
															assign node31532 = (inp[14]) ? 4'b1101 : node31533;
																assign node31533 = (inp[7]) ? 4'b1100 : 4'b1101;
														assign node31538 = (inp[7]) ? node31544 : node31539;
															assign node31539 = (inp[14]) ? 4'b1101 : node31540;
																assign node31540 = (inp[2]) ? 4'b1101 : 4'b1100;
															assign node31544 = (inp[14]) ? 4'b1100 : node31545;
																assign node31545 = (inp[2]) ? 4'b1100 : 4'b1101;
													assign node31549 = (inp[2]) ? node31559 : node31550;
														assign node31550 = (inp[8]) ? 4'b1111 : node31551;
															assign node31551 = (inp[14]) ? node31555 : node31552;
																assign node31552 = (inp[7]) ? 4'b1110 : 4'b1111;
																assign node31555 = (inp[7]) ? 4'b1111 : 4'b1110;
														assign node31559 = (inp[7]) ? node31563 : node31560;
															assign node31560 = (inp[8]) ? 4'b1111 : 4'b1110;
															assign node31563 = (inp[8]) ? 4'b1110 : 4'b1111;
												assign node31566 = (inp[2]) ? node31586 : node31567;
													assign node31567 = (inp[7]) ? node31579 : node31568;
														assign node31568 = (inp[5]) ? node31574 : node31569;
															assign node31569 = (inp[8]) ? node31571 : 4'b1111;
																assign node31571 = (inp[14]) ? 4'b1111 : 4'b1110;
															assign node31574 = (inp[14]) ? node31576 : 4'b1111;
																assign node31576 = (inp[8]) ? 4'b1111 : 4'b1110;
														assign node31579 = (inp[14]) ? node31583 : node31580;
															assign node31580 = (inp[8]) ? 4'b1111 : 4'b1110;
															assign node31583 = (inp[8]) ? 4'b1110 : 4'b1111;
													assign node31586 = (inp[14]) ? node31594 : node31587;
														assign node31587 = (inp[7]) ? node31591 : node31588;
															assign node31588 = (inp[8]) ? 4'b1111 : 4'b1110;
															assign node31591 = (inp[8]) ? 4'b1110 : 4'b1111;
														assign node31594 = (inp[5]) ? 4'b1110 : node31595;
															assign node31595 = (inp[8]) ? node31599 : node31596;
																assign node31596 = (inp[7]) ? 4'b1111 : 4'b1110;
																assign node31599 = (inp[7]) ? 4'b1110 : 4'b1111;
											assign node31603 = (inp[3]) ? node31637 : node31604;
												assign node31604 = (inp[5]) ? node31632 : node31605;
													assign node31605 = (inp[14]) ? node31619 : node31606;
														assign node31606 = (inp[8]) ? node31614 : node31607;
															assign node31607 = (inp[7]) ? node31611 : node31608;
																assign node31608 = (inp[2]) ? 4'b1110 : 4'b1111;
																assign node31611 = (inp[2]) ? 4'b1111 : 4'b1110;
															assign node31614 = (inp[7]) ? 4'b1110 : node31615;
																assign node31615 = (inp[2]) ? 4'b1111 : 4'b1110;
														assign node31619 = (inp[2]) ? node31625 : node31620;
															assign node31620 = (inp[7]) ? node31622 : 4'b1111;
																assign node31622 = (inp[8]) ? 4'b1110 : 4'b1111;
															assign node31625 = (inp[7]) ? node31629 : node31626;
																assign node31626 = (inp[8]) ? 4'b1111 : 4'b1110;
																assign node31629 = (inp[8]) ? 4'b1110 : 4'b1111;
													assign node31632 = (inp[7]) ? 4'b1101 : node31633;
														assign node31633 = (inp[8]) ? 4'b1101 : 4'b1100;
												assign node31637 = (inp[14]) ? node31647 : node31638;
													assign node31638 = (inp[5]) ? node31640 : 4'b1101;
														assign node31640 = (inp[7]) ? node31642 : 4'b1101;
															assign node31642 = (inp[2]) ? node31644 : 4'b1100;
																assign node31644 = (inp[8]) ? 4'b1100 : 4'b1101;
													assign node31647 = (inp[2]) ? node31655 : node31648;
														assign node31648 = (inp[8]) ? node31652 : node31649;
															assign node31649 = (inp[7]) ? 4'b1101 : 4'b1100;
															assign node31652 = (inp[7]) ? 4'b1100 : 4'b1101;
														assign node31655 = (inp[8]) ? node31659 : node31656;
															assign node31656 = (inp[7]) ? 4'b1101 : 4'b1100;
															assign node31659 = (inp[7]) ? 4'b1100 : 4'b1101;
								assign node31662 = (inp[4]) ? node31992 : node31663;
									assign node31663 = (inp[5]) ? node31853 : node31664;
										assign node31664 = (inp[2]) ? node31756 : node31665;
											assign node31665 = (inp[8]) ? node31705 : node31666;
												assign node31666 = (inp[3]) ? node31680 : node31667;
													assign node31667 = (inp[15]) ? node31671 : node31668;
														assign node31668 = (inp[0]) ? 4'b1101 : 4'b1111;
														assign node31671 = (inp[0]) ? 4'b1111 : node31672;
															assign node31672 = (inp[7]) ? node31676 : node31673;
																assign node31673 = (inp[14]) ? 4'b1100 : 4'b1101;
																assign node31676 = (inp[14]) ? 4'b1101 : 4'b1100;
													assign node31680 = (inp[0]) ? node31694 : node31681;
														assign node31681 = (inp[15]) ? node31689 : node31682;
															assign node31682 = (inp[14]) ? node31686 : node31683;
																assign node31683 = (inp[7]) ? 4'b1100 : 4'b1101;
																assign node31686 = (inp[7]) ? 4'b1101 : 4'b1100;
															assign node31689 = (inp[14]) ? node31691 : 4'b1110;
																assign node31691 = (inp[7]) ? 4'b1111 : 4'b1110;
														assign node31694 = (inp[15]) ? node31700 : node31695;
															assign node31695 = (inp[7]) ? node31697 : 4'b1111;
																assign node31697 = (inp[14]) ? 4'b1111 : 4'b1110;
															assign node31700 = (inp[7]) ? 4'b1101 : node31701;
																assign node31701 = (inp[14]) ? 4'b1100 : 4'b1101;
												assign node31705 = (inp[15]) ? node31733 : node31706;
													assign node31706 = (inp[14]) ? node31720 : node31707;
														assign node31707 = (inp[7]) ? node31715 : node31708;
															assign node31708 = (inp[0]) ? node31712 : node31709;
																assign node31709 = (inp[3]) ? 4'b1100 : 4'b1110;
																assign node31712 = (inp[3]) ? 4'b1110 : 4'b1100;
															assign node31715 = (inp[0]) ? node31717 : 4'b1101;
																assign node31717 = (inp[3]) ? 4'b1111 : 4'b1101;
														assign node31720 = (inp[7]) ? node31728 : node31721;
															assign node31721 = (inp[0]) ? node31725 : node31722;
																assign node31722 = (inp[3]) ? 4'b1101 : 4'b1111;
																assign node31725 = (inp[3]) ? 4'b1111 : 4'b1101;
															assign node31728 = (inp[0]) ? node31730 : 4'b1110;
																assign node31730 = (inp[3]) ? 4'b1110 : 4'b1100;
													assign node31733 = (inp[3]) ? node31747 : node31734;
														assign node31734 = (inp[0]) ? node31742 : node31735;
															assign node31735 = (inp[7]) ? node31739 : node31736;
																assign node31736 = (inp[14]) ? 4'b1101 : 4'b1100;
																assign node31739 = (inp[14]) ? 4'b1100 : 4'b1101;
															assign node31742 = (inp[14]) ? 4'b1111 : node31743;
																assign node31743 = (inp[7]) ? 4'b1111 : 4'b1110;
														assign node31747 = (inp[0]) ? node31751 : node31748;
															assign node31748 = (inp[14]) ? 4'b1110 : 4'b1111;
															assign node31751 = (inp[14]) ? node31753 : 4'b1100;
																assign node31753 = (inp[7]) ? 4'b1100 : 4'b1101;
											assign node31756 = (inp[14]) ? node31802 : node31757;
												assign node31757 = (inp[0]) ? node31785 : node31758;
													assign node31758 = (inp[7]) ? node31772 : node31759;
														assign node31759 = (inp[8]) ? node31767 : node31760;
															assign node31760 = (inp[15]) ? node31764 : node31761;
																assign node31761 = (inp[3]) ? 4'b1100 : 4'b1110;
																assign node31764 = (inp[3]) ? 4'b1110 : 4'b1100;
															assign node31767 = (inp[3]) ? 4'b1101 : node31768;
																assign node31768 = (inp[15]) ? 4'b1101 : 4'b1111;
														assign node31772 = (inp[8]) ? node31778 : node31773;
															assign node31773 = (inp[3]) ? node31775 : 4'b1101;
																assign node31775 = (inp[15]) ? 4'b1111 : 4'b1101;
															assign node31778 = (inp[15]) ? node31782 : node31779;
																assign node31779 = (inp[3]) ? 4'b1100 : 4'b1110;
																assign node31782 = (inp[3]) ? 4'b1110 : 4'b1100;
													assign node31785 = (inp[15]) ? node31793 : node31786;
														assign node31786 = (inp[3]) ? node31788 : 4'b1100;
															assign node31788 = (inp[8]) ? 4'b1110 : node31789;
																assign node31789 = (inp[7]) ? 4'b1111 : 4'b1110;
														assign node31793 = (inp[3]) ? node31797 : node31794;
															assign node31794 = (inp[8]) ? 4'b1111 : 4'b1110;
															assign node31797 = (inp[8]) ? 4'b1100 : node31798;
																assign node31798 = (inp[7]) ? 4'b1101 : 4'b1100;
												assign node31802 = (inp[7]) ? node31826 : node31803;
													assign node31803 = (inp[8]) ? node31813 : node31804;
														assign node31804 = (inp[0]) ? node31806 : 4'b1100;
															assign node31806 = (inp[3]) ? node31810 : node31807;
																assign node31807 = (inp[15]) ? 4'b1110 : 4'b1100;
																assign node31810 = (inp[15]) ? 4'b1100 : 4'b1110;
														assign node31813 = (inp[15]) ? node31819 : node31814;
															assign node31814 = (inp[0]) ? 4'b1101 : node31815;
																assign node31815 = (inp[3]) ? 4'b1101 : 4'b1111;
															assign node31819 = (inp[3]) ? node31823 : node31820;
																assign node31820 = (inp[0]) ? 4'b1111 : 4'b1101;
																assign node31823 = (inp[0]) ? 4'b1101 : 4'b1111;
													assign node31826 = (inp[8]) ? node31838 : node31827;
														assign node31827 = (inp[3]) ? node31833 : node31828;
															assign node31828 = (inp[0]) ? node31830 : 4'b1111;
																assign node31830 = (inp[15]) ? 4'b1111 : 4'b1101;
															assign node31833 = (inp[15]) ? 4'b1101 : node31834;
																assign node31834 = (inp[0]) ? 4'b1111 : 4'b1101;
														assign node31838 = (inp[0]) ? node31846 : node31839;
															assign node31839 = (inp[15]) ? node31843 : node31840;
																assign node31840 = (inp[3]) ? 4'b1100 : 4'b1110;
																assign node31843 = (inp[3]) ? 4'b1110 : 4'b1100;
															assign node31846 = (inp[15]) ? node31850 : node31847;
																assign node31847 = (inp[3]) ? 4'b1110 : 4'b1100;
																assign node31850 = (inp[3]) ? 4'b1100 : 4'b1110;
										assign node31853 = (inp[14]) ? node31929 : node31854;
											assign node31854 = (inp[0]) ? node31886 : node31855;
												assign node31855 = (inp[15]) ? node31871 : node31856;
													assign node31856 = (inp[2]) ? node31864 : node31857;
														assign node31857 = (inp[8]) ? node31861 : node31858;
															assign node31858 = (inp[7]) ? 4'b1100 : 4'b1101;
															assign node31861 = (inp[7]) ? 4'b1101 : 4'b1100;
														assign node31864 = (inp[8]) ? node31868 : node31865;
															assign node31865 = (inp[7]) ? 4'b1101 : 4'b1100;
															assign node31868 = (inp[7]) ? 4'b1100 : 4'b1101;
													assign node31871 = (inp[8]) ? node31881 : node31872;
														assign node31872 = (inp[3]) ? node31874 : 4'b1111;
															assign node31874 = (inp[7]) ? node31878 : node31875;
																assign node31875 = (inp[2]) ? 4'b1110 : 4'b1111;
																assign node31878 = (inp[2]) ? 4'b1111 : 4'b1110;
														assign node31881 = (inp[2]) ? 4'b1110 : node31882;
															assign node31882 = (inp[7]) ? 4'b1111 : 4'b1110;
												assign node31886 = (inp[15]) ? node31906 : node31887;
													assign node31887 = (inp[7]) ? node31901 : node31888;
														assign node31888 = (inp[3]) ? node31894 : node31889;
															assign node31889 = (inp[8]) ? 4'b1111 : node31890;
																assign node31890 = (inp[2]) ? 4'b1110 : 4'b1111;
															assign node31894 = (inp[2]) ? node31898 : node31895;
																assign node31895 = (inp[8]) ? 4'b1110 : 4'b1111;
																assign node31898 = (inp[8]) ? 4'b1111 : 4'b1110;
														assign node31901 = (inp[2]) ? 4'b1111 : node31902;
															assign node31902 = (inp[8]) ? 4'b1111 : 4'b1110;
													assign node31906 = (inp[3]) ? node31920 : node31907;
														assign node31907 = (inp[7]) ? node31913 : node31908;
															assign node31908 = (inp[8]) ? 4'b1101 : node31909;
																assign node31909 = (inp[2]) ? 4'b1100 : 4'b1101;
															assign node31913 = (inp[2]) ? node31917 : node31914;
																assign node31914 = (inp[8]) ? 4'b1101 : 4'b1100;
																assign node31917 = (inp[8]) ? 4'b1100 : 4'b1101;
														assign node31920 = (inp[8]) ? node31922 : 4'b1101;
															assign node31922 = (inp[2]) ? node31926 : node31923;
																assign node31923 = (inp[7]) ? 4'b1101 : 4'b1100;
																assign node31926 = (inp[7]) ? 4'b1100 : 4'b1101;
											assign node31929 = (inp[3]) ? node31961 : node31930;
												assign node31930 = (inp[0]) ? node31946 : node31931;
													assign node31931 = (inp[15]) ? node31939 : node31932;
														assign node31932 = (inp[7]) ? node31936 : node31933;
															assign node31933 = (inp[8]) ? 4'b1101 : 4'b1100;
															assign node31936 = (inp[8]) ? 4'b1100 : 4'b1101;
														assign node31939 = (inp[8]) ? node31943 : node31940;
															assign node31940 = (inp[7]) ? 4'b1111 : 4'b1110;
															assign node31943 = (inp[7]) ? 4'b1110 : 4'b1111;
													assign node31946 = (inp[15]) ? node31954 : node31947;
														assign node31947 = (inp[8]) ? node31951 : node31948;
															assign node31948 = (inp[7]) ? 4'b1111 : 4'b1110;
															assign node31951 = (inp[7]) ? 4'b1110 : 4'b1111;
														assign node31954 = (inp[7]) ? node31958 : node31955;
															assign node31955 = (inp[8]) ? 4'b1101 : 4'b1100;
															assign node31958 = (inp[8]) ? 4'b1100 : 4'b1101;
												assign node31961 = (inp[7]) ? node31975 : node31962;
													assign node31962 = (inp[8]) ? node31968 : node31963;
														assign node31963 = (inp[0]) ? node31965 : 4'b1110;
															assign node31965 = (inp[15]) ? 4'b1100 : 4'b1110;
														assign node31968 = (inp[0]) ? node31972 : node31969;
															assign node31969 = (inp[15]) ? 4'b1111 : 4'b1101;
															assign node31972 = (inp[15]) ? 4'b1101 : 4'b1111;
													assign node31975 = (inp[8]) ? node31983 : node31976;
														assign node31976 = (inp[15]) ? node31980 : node31977;
															assign node31977 = (inp[0]) ? 4'b1111 : 4'b1101;
															assign node31980 = (inp[0]) ? 4'b1101 : 4'b1111;
														assign node31983 = (inp[2]) ? 4'b1110 : node31984;
															assign node31984 = (inp[0]) ? node31988 : node31985;
																assign node31985 = (inp[15]) ? 4'b1110 : 4'b1100;
																assign node31988 = (inp[15]) ? 4'b1100 : 4'b1110;
									assign node31992 = (inp[7]) ? node32128 : node31993;
										assign node31993 = (inp[8]) ? node32071 : node31994;
											assign node31994 = (inp[14]) ? node32022 : node31995;
												assign node31995 = (inp[2]) ? node32011 : node31996;
													assign node31996 = (inp[15]) ? node32006 : node31997;
														assign node31997 = (inp[0]) ? node32001 : node31998;
															assign node31998 = (inp[5]) ? 4'b1001 : 4'b1011;
															assign node32001 = (inp[5]) ? 4'b1011 : node32002;
																assign node32002 = (inp[3]) ? 4'b1011 : 4'b1001;
														assign node32006 = (inp[5]) ? node32008 : 4'b1001;
															assign node32008 = (inp[0]) ? 4'b1001 : 4'b1011;
													assign node32011 = (inp[5]) ? 4'b1000 : node32012;
														assign node32012 = (inp[15]) ? 4'b1010 : node32013;
															assign node32013 = (inp[0]) ? node32017 : node32014;
																assign node32014 = (inp[3]) ? 4'b1000 : 4'b1010;
																assign node32017 = (inp[3]) ? 4'b1010 : 4'b1000;
												assign node32022 = (inp[2]) ? node32046 : node32023;
													assign node32023 = (inp[0]) ? node32035 : node32024;
														assign node32024 = (inp[15]) ? node32030 : node32025;
															assign node32025 = (inp[3]) ? 4'b1000 : node32026;
																assign node32026 = (inp[5]) ? 4'b1000 : 4'b1010;
															assign node32030 = (inp[3]) ? 4'b1010 : node32031;
																assign node32031 = (inp[5]) ? 4'b1010 : 4'b1000;
														assign node32035 = (inp[15]) ? node32041 : node32036;
															assign node32036 = (inp[5]) ? 4'b1010 : node32037;
																assign node32037 = (inp[3]) ? 4'b1010 : 4'b1000;
															assign node32041 = (inp[5]) ? 4'b1000 : node32042;
																assign node32042 = (inp[3]) ? 4'b1000 : 4'b1010;
													assign node32046 = (inp[3]) ? node32062 : node32047;
														assign node32047 = (inp[5]) ? node32055 : node32048;
															assign node32048 = (inp[0]) ? node32052 : node32049;
																assign node32049 = (inp[15]) ? 4'b1000 : 4'b1010;
																assign node32052 = (inp[15]) ? 4'b1010 : 4'b1000;
															assign node32055 = (inp[15]) ? node32059 : node32056;
																assign node32056 = (inp[0]) ? 4'b1010 : 4'b1000;
																assign node32059 = (inp[0]) ? 4'b1000 : 4'b1010;
														assign node32062 = (inp[5]) ? 4'b1000 : node32063;
															assign node32063 = (inp[0]) ? node32067 : node32064;
																assign node32064 = (inp[15]) ? 4'b1010 : 4'b1000;
																assign node32067 = (inp[15]) ? 4'b1000 : 4'b1010;
											assign node32071 = (inp[2]) ? node32105 : node32072;
												assign node32072 = (inp[14]) ? node32090 : node32073;
													assign node32073 = (inp[15]) ? node32079 : node32074;
														assign node32074 = (inp[0]) ? node32076 : 4'b1000;
															assign node32076 = (inp[5]) ? 4'b1010 : 4'b1000;
														assign node32079 = (inp[0]) ? node32085 : node32080;
															assign node32080 = (inp[3]) ? 4'b1010 : node32081;
																assign node32081 = (inp[5]) ? 4'b1010 : 4'b1000;
															assign node32085 = (inp[5]) ? 4'b1000 : node32086;
																assign node32086 = (inp[3]) ? 4'b1000 : 4'b1010;
													assign node32090 = (inp[3]) ? node32100 : node32091;
														assign node32091 = (inp[15]) ? node32093 : 4'b1001;
															assign node32093 = (inp[5]) ? node32097 : node32094;
																assign node32094 = (inp[0]) ? 4'b1011 : 4'b1001;
																assign node32097 = (inp[0]) ? 4'b1001 : 4'b1011;
														assign node32100 = (inp[5]) ? node32102 : 4'b1011;
															assign node32102 = (inp[15]) ? 4'b1001 : 4'b1011;
												assign node32105 = (inp[15]) ? node32117 : node32106;
													assign node32106 = (inp[0]) ? node32112 : node32107;
														assign node32107 = (inp[3]) ? 4'b1001 : node32108;
															assign node32108 = (inp[5]) ? 4'b1001 : 4'b1011;
														assign node32112 = (inp[5]) ? 4'b1011 : node32113;
															assign node32113 = (inp[3]) ? 4'b1011 : 4'b1001;
													assign node32117 = (inp[0]) ? node32123 : node32118;
														assign node32118 = (inp[3]) ? 4'b1011 : node32119;
															assign node32119 = (inp[5]) ? 4'b1011 : 4'b1001;
														assign node32123 = (inp[3]) ? 4'b1001 : node32124;
															assign node32124 = (inp[5]) ? 4'b1001 : 4'b1011;
										assign node32128 = (inp[8]) ? node32204 : node32129;
											assign node32129 = (inp[14]) ? node32161 : node32130;
												assign node32130 = (inp[2]) ? node32142 : node32131;
													assign node32131 = (inp[0]) ? node32137 : node32132;
														assign node32132 = (inp[5]) ? node32134 : 4'b1000;
															assign node32134 = (inp[15]) ? 4'b1010 : 4'b1000;
														assign node32137 = (inp[15]) ? node32139 : 4'b1010;
															assign node32139 = (inp[3]) ? 4'b1000 : 4'b1010;
													assign node32142 = (inp[0]) ? node32152 : node32143;
														assign node32143 = (inp[15]) ? node32149 : node32144;
															assign node32144 = (inp[3]) ? 4'b1001 : node32145;
																assign node32145 = (inp[5]) ? 4'b1001 : 4'b1011;
															assign node32149 = (inp[5]) ? 4'b1011 : 4'b1001;
														assign node32152 = (inp[15]) ? node32156 : node32153;
															assign node32153 = (inp[3]) ? 4'b1011 : 4'b1001;
															assign node32156 = (inp[3]) ? 4'b1001 : node32157;
																assign node32157 = (inp[5]) ? 4'b1001 : 4'b1011;
												assign node32161 = (inp[3]) ? node32183 : node32162;
													assign node32162 = (inp[0]) ? node32178 : node32163;
														assign node32163 = (inp[2]) ? node32171 : node32164;
															assign node32164 = (inp[15]) ? node32168 : node32165;
																assign node32165 = (inp[5]) ? 4'b1001 : 4'b1011;
																assign node32168 = (inp[5]) ? 4'b1011 : 4'b1001;
															assign node32171 = (inp[15]) ? node32175 : node32172;
																assign node32172 = (inp[5]) ? 4'b1001 : 4'b1011;
																assign node32175 = (inp[5]) ? 4'b1011 : 4'b1001;
														assign node32178 = (inp[5]) ? node32180 : 4'b1011;
															assign node32180 = (inp[2]) ? 4'b1011 : 4'b1001;
													assign node32183 = (inp[2]) ? node32197 : node32184;
														assign node32184 = (inp[5]) ? node32192 : node32185;
															assign node32185 = (inp[0]) ? node32189 : node32186;
																assign node32186 = (inp[15]) ? 4'b1011 : 4'b1001;
																assign node32189 = (inp[15]) ? 4'b1001 : 4'b1011;
															assign node32192 = (inp[15]) ? node32194 : 4'b1001;
																assign node32194 = (inp[0]) ? 4'b1001 : 4'b1011;
														assign node32197 = (inp[15]) ? node32201 : node32198;
															assign node32198 = (inp[0]) ? 4'b1011 : 4'b1001;
															assign node32201 = (inp[0]) ? 4'b1001 : 4'b1011;
											assign node32204 = (inp[2]) ? node32234 : node32205;
												assign node32205 = (inp[14]) ? node32223 : node32206;
													assign node32206 = (inp[3]) ? node32216 : node32207;
														assign node32207 = (inp[15]) ? node32209 : 4'b1001;
															assign node32209 = (inp[0]) ? node32213 : node32210;
																assign node32210 = (inp[5]) ? 4'b1011 : 4'b1001;
																assign node32213 = (inp[5]) ? 4'b1001 : 4'b1011;
														assign node32216 = (inp[0]) ? node32220 : node32217;
															assign node32217 = (inp[15]) ? 4'b1011 : 4'b1001;
															assign node32220 = (inp[15]) ? 4'b1001 : 4'b1011;
													assign node32223 = (inp[15]) ? node32227 : node32224;
														assign node32224 = (inp[0]) ? 4'b1010 : 4'b1000;
														assign node32227 = (inp[0]) ? 4'b1000 : node32228;
															assign node32228 = (inp[3]) ? 4'b1010 : node32229;
																assign node32229 = (inp[5]) ? 4'b1010 : 4'b1000;
												assign node32234 = (inp[3]) ? node32256 : node32235;
													assign node32235 = (inp[14]) ? node32251 : node32236;
														assign node32236 = (inp[5]) ? node32244 : node32237;
															assign node32237 = (inp[15]) ? node32241 : node32238;
																assign node32238 = (inp[0]) ? 4'b1000 : 4'b1010;
																assign node32241 = (inp[0]) ? 4'b1010 : 4'b1000;
															assign node32244 = (inp[0]) ? node32248 : node32245;
																assign node32245 = (inp[15]) ? 4'b1010 : 4'b1000;
																assign node32248 = (inp[15]) ? 4'b1000 : 4'b1010;
														assign node32251 = (inp[15]) ? node32253 : 4'b1010;
															assign node32253 = (inp[5]) ? 4'b1010 : 4'b1000;
													assign node32256 = (inp[0]) ? node32260 : node32257;
														assign node32257 = (inp[15]) ? 4'b1010 : 4'b1000;
														assign node32260 = (inp[15]) ? 4'b1000 : 4'b1010;
							assign node32263 = (inp[3]) ? node32861 : node32264;
								assign node32264 = (inp[0]) ? node32558 : node32265;
									assign node32265 = (inp[15]) ? node32403 : node32266;
										assign node32266 = (inp[5]) ? node32334 : node32267;
											assign node32267 = (inp[4]) ? node32303 : node32268;
												assign node32268 = (inp[9]) ? node32286 : node32269;
													assign node32269 = (inp[8]) ? node32279 : node32270;
														assign node32270 = (inp[14]) ? node32276 : node32271;
															assign node32271 = (inp[2]) ? 4'b1010 : node32272;
																assign node32272 = (inp[7]) ? 4'b1010 : 4'b1011;
															assign node32276 = (inp[7]) ? 4'b1011 : 4'b1010;
														assign node32279 = (inp[14]) ? 4'b1011 : node32280;
															assign node32280 = (inp[2]) ? 4'b1011 : node32281;
																assign node32281 = (inp[7]) ? 4'b1011 : 4'b1010;
													assign node32286 = (inp[8]) ? node32296 : node32287;
														assign node32287 = (inp[7]) ? node32293 : node32288;
															assign node32288 = (inp[2]) ? 4'b1110 : node32289;
																assign node32289 = (inp[14]) ? 4'b1110 : 4'b1111;
															assign node32293 = (inp[14]) ? 4'b1111 : 4'b1110;
														assign node32296 = (inp[7]) ? 4'b1110 : node32297;
															assign node32297 = (inp[2]) ? 4'b1111 : node32298;
																assign node32298 = (inp[14]) ? 4'b1111 : 4'b1110;
												assign node32303 = (inp[9]) ? node32319 : node32304;
													assign node32304 = (inp[2]) ? node32312 : node32305;
														assign node32305 = (inp[8]) ? node32307 : 4'b1110;
															assign node32307 = (inp[7]) ? node32309 : 4'b1110;
																assign node32309 = (inp[14]) ? 4'b1110 : 4'b1111;
														assign node32312 = (inp[7]) ? node32316 : node32313;
															assign node32313 = (inp[8]) ? 4'b1111 : 4'b1110;
															assign node32316 = (inp[8]) ? 4'b1110 : 4'b1111;
													assign node32319 = (inp[7]) ? node32327 : node32320;
														assign node32320 = (inp[14]) ? 4'b1010 : node32321;
															assign node32321 = (inp[2]) ? 4'b1010 : node32322;
																assign node32322 = (inp[8]) ? 4'b1010 : 4'b1011;
														assign node32327 = (inp[8]) ? node32331 : node32328;
															assign node32328 = (inp[14]) ? 4'b1011 : 4'b1010;
															assign node32331 = (inp[14]) ? 4'b1010 : 4'b1011;
											assign node32334 = (inp[9]) ? node32370 : node32335;
												assign node32335 = (inp[4]) ? node32359 : node32336;
													assign node32336 = (inp[14]) ? node32352 : node32337;
														assign node32337 = (inp[2]) ? node32345 : node32338;
															assign node32338 = (inp[7]) ? node32342 : node32339;
																assign node32339 = (inp[8]) ? 4'b1010 : 4'b1011;
																assign node32342 = (inp[8]) ? 4'b1011 : 4'b1010;
															assign node32345 = (inp[8]) ? node32349 : node32346;
																assign node32346 = (inp[7]) ? 4'b1011 : 4'b1010;
																assign node32349 = (inp[7]) ? 4'b1010 : 4'b1011;
														assign node32352 = (inp[8]) ? node32356 : node32353;
															assign node32353 = (inp[7]) ? 4'b1011 : 4'b1010;
															assign node32356 = (inp[7]) ? 4'b1010 : 4'b1011;
													assign node32359 = (inp[8]) ? node32365 : node32360;
														assign node32360 = (inp[14]) ? node32362 : 4'b1101;
															assign node32362 = (inp[7]) ? 4'b1101 : 4'b1100;
														assign node32365 = (inp[7]) ? 4'b1100 : node32366;
															assign node32366 = (inp[2]) ? 4'b1101 : 4'b1100;
												assign node32370 = (inp[4]) ? node32384 : node32371;
													assign node32371 = (inp[2]) ? node32377 : node32372;
														assign node32372 = (inp[14]) ? 4'b1101 : node32373;
															assign node32373 = (inp[8]) ? 4'b1101 : 4'b1100;
														assign node32377 = (inp[8]) ? node32381 : node32378;
															assign node32378 = (inp[7]) ? 4'b1101 : 4'b1100;
															assign node32381 = (inp[7]) ? 4'b1100 : 4'b1101;
													assign node32384 = (inp[8]) ? node32396 : node32385;
														assign node32385 = (inp[7]) ? node32391 : node32386;
															assign node32386 = (inp[2]) ? 4'b1000 : node32387;
																assign node32387 = (inp[14]) ? 4'b1000 : 4'b1001;
															assign node32391 = (inp[2]) ? 4'b1001 : node32392;
																assign node32392 = (inp[14]) ? 4'b1001 : 4'b1000;
														assign node32396 = (inp[7]) ? 4'b1000 : node32397;
															assign node32397 = (inp[14]) ? 4'b1001 : node32398;
																assign node32398 = (inp[2]) ? 4'b1001 : 4'b1000;
										assign node32403 = (inp[5]) ? node32489 : node32404;
											assign node32404 = (inp[14]) ? node32446 : node32405;
												assign node32405 = (inp[7]) ? node32429 : node32406;
													assign node32406 = (inp[8]) ? node32420 : node32407;
														assign node32407 = (inp[2]) ? node32413 : node32408;
															assign node32408 = (inp[4]) ? node32410 : 4'b1001;
																assign node32410 = (inp[9]) ? 4'b1001 : 4'b1101;
															assign node32413 = (inp[4]) ? node32417 : node32414;
																assign node32414 = (inp[9]) ? 4'b1100 : 4'b1000;
																assign node32417 = (inp[9]) ? 4'b1000 : 4'b1100;
														assign node32420 = (inp[2]) ? node32424 : node32421;
															assign node32421 = (inp[9]) ? 4'b1100 : 4'b1000;
															assign node32424 = (inp[9]) ? 4'b1101 : node32425;
																assign node32425 = (inp[4]) ? 4'b1101 : 4'b1001;
													assign node32429 = (inp[2]) ? node32437 : node32430;
														assign node32430 = (inp[8]) ? 4'b1101 : node32431;
															assign node32431 = (inp[4]) ? node32433 : 4'b1100;
																assign node32433 = (inp[9]) ? 4'b1000 : 4'b1100;
														assign node32437 = (inp[8]) ? node32439 : 4'b1001;
															assign node32439 = (inp[9]) ? node32443 : node32440;
																assign node32440 = (inp[4]) ? 4'b1100 : 4'b1000;
																assign node32443 = (inp[4]) ? 4'b1000 : 4'b1100;
												assign node32446 = (inp[2]) ? node32464 : node32447;
													assign node32447 = (inp[4]) ? node32455 : node32448;
														assign node32448 = (inp[9]) ? 4'b1100 : node32449;
															assign node32449 = (inp[7]) ? node32451 : 4'b1000;
																assign node32451 = (inp[8]) ? 4'b1000 : 4'b1001;
														assign node32455 = (inp[9]) ? node32457 : 4'b1101;
															assign node32457 = (inp[7]) ? node32461 : node32458;
																assign node32458 = (inp[8]) ? 4'b1001 : 4'b1000;
																assign node32461 = (inp[8]) ? 4'b1000 : 4'b1001;
													assign node32464 = (inp[7]) ? node32480 : node32465;
														assign node32465 = (inp[8]) ? node32473 : node32466;
															assign node32466 = (inp[9]) ? node32470 : node32467;
																assign node32467 = (inp[4]) ? 4'b1100 : 4'b1000;
																assign node32470 = (inp[4]) ? 4'b1000 : 4'b1100;
															assign node32473 = (inp[4]) ? node32477 : node32474;
																assign node32474 = (inp[9]) ? 4'b1101 : 4'b1001;
																assign node32477 = (inp[9]) ? 4'b1001 : 4'b1101;
														assign node32480 = (inp[8]) ? 4'b1100 : node32481;
															assign node32481 = (inp[9]) ? node32485 : node32482;
																assign node32482 = (inp[4]) ? 4'b1101 : 4'b1001;
																assign node32485 = (inp[4]) ? 4'b1001 : 4'b1101;
											assign node32489 = (inp[4]) ? node32519 : node32490;
												assign node32490 = (inp[9]) ? node32506 : node32491;
													assign node32491 = (inp[14]) ? node32499 : node32492;
														assign node32492 = (inp[7]) ? node32494 : 4'b1000;
															assign node32494 = (inp[8]) ? node32496 : 4'b1000;
																assign node32496 = (inp[2]) ? 4'b1000 : 4'b1001;
														assign node32499 = (inp[7]) ? node32503 : node32500;
															assign node32500 = (inp[8]) ? 4'b1001 : 4'b1000;
															assign node32503 = (inp[8]) ? 4'b1000 : 4'b1001;
													assign node32506 = (inp[7]) ? node32514 : node32507;
														assign node32507 = (inp[8]) ? 4'b1111 : node32508;
															assign node32508 = (inp[14]) ? 4'b1110 : node32509;
																assign node32509 = (inp[2]) ? 4'b1110 : 4'b1111;
														assign node32514 = (inp[14]) ? node32516 : 4'b1110;
															assign node32516 = (inp[2]) ? 4'b1110 : 4'b1111;
												assign node32519 = (inp[9]) ? node32537 : node32520;
													assign node32520 = (inp[7]) ? node32532 : node32521;
														assign node32521 = (inp[8]) ? node32527 : node32522;
															assign node32522 = (inp[14]) ? 4'b1110 : node32523;
																assign node32523 = (inp[2]) ? 4'b1110 : 4'b1111;
															assign node32527 = (inp[14]) ? 4'b1111 : node32528;
																assign node32528 = (inp[2]) ? 4'b1111 : 4'b1110;
														assign node32532 = (inp[8]) ? 4'b1110 : node32533;
															assign node32533 = (inp[14]) ? 4'b1111 : 4'b1110;
													assign node32537 = (inp[14]) ? node32551 : node32538;
														assign node32538 = (inp[2]) ? node32546 : node32539;
															assign node32539 = (inp[8]) ? node32543 : node32540;
																assign node32540 = (inp[7]) ? 4'b1010 : 4'b1011;
																assign node32543 = (inp[7]) ? 4'b1011 : 4'b1010;
															assign node32546 = (inp[8]) ? 4'b1011 : node32547;
																assign node32547 = (inp[7]) ? 4'b1011 : 4'b1010;
														assign node32551 = (inp[8]) ? node32555 : node32552;
															assign node32552 = (inp[7]) ? 4'b1011 : 4'b1010;
															assign node32555 = (inp[7]) ? 4'b1010 : 4'b1011;
									assign node32558 = (inp[15]) ? node32714 : node32559;
										assign node32559 = (inp[5]) ? node32633 : node32560;
											assign node32560 = (inp[7]) ? node32598 : node32561;
												assign node32561 = (inp[8]) ? node32581 : node32562;
													assign node32562 = (inp[14]) ? node32572 : node32563;
														assign node32563 = (inp[2]) ? node32567 : node32564;
															assign node32564 = (inp[9]) ? 4'b1001 : 4'b1101;
															assign node32567 = (inp[4]) ? node32569 : 4'b1000;
																assign node32569 = (inp[9]) ? 4'b1000 : 4'b1100;
														assign node32572 = (inp[2]) ? 4'b1100 : node32573;
															assign node32573 = (inp[4]) ? node32577 : node32574;
																assign node32574 = (inp[9]) ? 4'b1100 : 4'b1000;
																assign node32577 = (inp[9]) ? 4'b1000 : 4'b1100;
													assign node32581 = (inp[2]) ? node32591 : node32582;
														assign node32582 = (inp[14]) ? 4'b1101 : node32583;
															assign node32583 = (inp[4]) ? node32587 : node32584;
																assign node32584 = (inp[9]) ? 4'b1100 : 4'b1000;
																assign node32587 = (inp[9]) ? 4'b1000 : 4'b1100;
														assign node32591 = (inp[9]) ? node32595 : node32592;
															assign node32592 = (inp[4]) ? 4'b1101 : 4'b1001;
															assign node32595 = (inp[4]) ? 4'b1001 : 4'b1101;
												assign node32598 = (inp[8]) ? node32616 : node32599;
													assign node32599 = (inp[14]) ? node32609 : node32600;
														assign node32600 = (inp[2]) ? node32602 : 4'b1100;
															assign node32602 = (inp[9]) ? node32606 : node32603;
																assign node32603 = (inp[4]) ? 4'b1101 : 4'b1001;
																assign node32606 = (inp[4]) ? 4'b1001 : 4'b1101;
														assign node32609 = (inp[9]) ? node32613 : node32610;
															assign node32610 = (inp[4]) ? 4'b1101 : 4'b1001;
															assign node32613 = (inp[4]) ? 4'b1001 : 4'b1101;
													assign node32616 = (inp[2]) ? node32626 : node32617;
														assign node32617 = (inp[14]) ? 4'b1000 : node32618;
															assign node32618 = (inp[4]) ? node32622 : node32619;
																assign node32619 = (inp[9]) ? 4'b1101 : 4'b1001;
																assign node32622 = (inp[9]) ? 4'b1001 : 4'b1101;
														assign node32626 = (inp[9]) ? node32630 : node32627;
															assign node32627 = (inp[4]) ? 4'b1100 : 4'b1000;
															assign node32630 = (inp[4]) ? 4'b1000 : 4'b1100;
											assign node32633 = (inp[4]) ? node32675 : node32634;
												assign node32634 = (inp[9]) ? node32654 : node32635;
													assign node32635 = (inp[2]) ? node32649 : node32636;
														assign node32636 = (inp[14]) ? node32642 : node32637;
															assign node32637 = (inp[8]) ? 4'b1001 : node32638;
																assign node32638 = (inp[7]) ? 4'b1000 : 4'b1001;
															assign node32642 = (inp[8]) ? node32646 : node32643;
																assign node32643 = (inp[7]) ? 4'b1001 : 4'b1000;
																assign node32646 = (inp[7]) ? 4'b1000 : 4'b1001;
														assign node32649 = (inp[7]) ? 4'b1000 : node32650;
															assign node32650 = (inp[8]) ? 4'b1001 : 4'b1000;
													assign node32654 = (inp[2]) ? node32668 : node32655;
														assign node32655 = (inp[7]) ? node32663 : node32656;
															assign node32656 = (inp[8]) ? node32660 : node32657;
																assign node32657 = (inp[14]) ? 4'b1110 : 4'b1111;
																assign node32660 = (inp[14]) ? 4'b1111 : 4'b1110;
															assign node32663 = (inp[8]) ? node32665 : 4'b1110;
																assign node32665 = (inp[14]) ? 4'b1110 : 4'b1111;
														assign node32668 = (inp[8]) ? node32672 : node32669;
															assign node32669 = (inp[7]) ? 4'b1111 : 4'b1110;
															assign node32672 = (inp[7]) ? 4'b1110 : 4'b1111;
												assign node32675 = (inp[9]) ? node32699 : node32676;
													assign node32676 = (inp[2]) ? node32692 : node32677;
														assign node32677 = (inp[8]) ? node32685 : node32678;
															assign node32678 = (inp[14]) ? node32682 : node32679;
																assign node32679 = (inp[7]) ? 4'b1110 : 4'b1111;
																assign node32682 = (inp[7]) ? 4'b1111 : 4'b1110;
															assign node32685 = (inp[14]) ? node32689 : node32686;
																assign node32686 = (inp[7]) ? 4'b1111 : 4'b1110;
																assign node32689 = (inp[7]) ? 4'b1110 : 4'b1111;
														assign node32692 = (inp[8]) ? node32696 : node32693;
															assign node32693 = (inp[7]) ? 4'b1111 : 4'b1110;
															assign node32696 = (inp[7]) ? 4'b1110 : 4'b1111;
													assign node32699 = (inp[8]) ? node32709 : node32700;
														assign node32700 = (inp[7]) ? node32706 : node32701;
															assign node32701 = (inp[14]) ? 4'b1010 : node32702;
																assign node32702 = (inp[2]) ? 4'b1010 : 4'b1011;
															assign node32706 = (inp[2]) ? 4'b1011 : 4'b1010;
														assign node32709 = (inp[7]) ? node32711 : 4'b1011;
															assign node32711 = (inp[2]) ? 4'b1010 : 4'b1011;
										assign node32714 = (inp[5]) ? node32792 : node32715;
											assign node32715 = (inp[2]) ? node32763 : node32716;
												assign node32716 = (inp[9]) ? node32740 : node32717;
													assign node32717 = (inp[4]) ? node32725 : node32718;
														assign node32718 = (inp[7]) ? 4'b1010 : node32719;
															assign node32719 = (inp[8]) ? node32721 : 4'b1010;
																assign node32721 = (inp[14]) ? 4'b1011 : 4'b1010;
														assign node32725 = (inp[7]) ? node32733 : node32726;
															assign node32726 = (inp[8]) ? node32730 : node32727;
																assign node32727 = (inp[14]) ? 4'b1110 : 4'b1111;
																assign node32730 = (inp[14]) ? 4'b1111 : 4'b1110;
															assign node32733 = (inp[14]) ? node32737 : node32734;
																assign node32734 = (inp[8]) ? 4'b1111 : 4'b1110;
																assign node32737 = (inp[8]) ? 4'b1110 : 4'b1111;
													assign node32740 = (inp[4]) ? node32750 : node32741;
														assign node32741 = (inp[14]) ? node32743 : 4'b1111;
															assign node32743 = (inp[7]) ? node32747 : node32744;
																assign node32744 = (inp[8]) ? 4'b1111 : 4'b1110;
																assign node32747 = (inp[8]) ? 4'b1110 : 4'b1111;
														assign node32750 = (inp[7]) ? node32756 : node32751;
															assign node32751 = (inp[8]) ? node32753 : 4'b1010;
																assign node32753 = (inp[14]) ? 4'b1011 : 4'b1010;
															assign node32756 = (inp[8]) ? node32760 : node32757;
																assign node32757 = (inp[14]) ? 4'b1011 : 4'b1010;
																assign node32760 = (inp[14]) ? 4'b1010 : 4'b1011;
												assign node32763 = (inp[4]) ? node32775 : node32764;
													assign node32764 = (inp[9]) ? node32772 : node32765;
														assign node32765 = (inp[7]) ? node32769 : node32766;
															assign node32766 = (inp[8]) ? 4'b1011 : 4'b1010;
															assign node32769 = (inp[8]) ? 4'b1010 : 4'b1011;
														assign node32772 = (inp[14]) ? 4'b1110 : 4'b1111;
													assign node32775 = (inp[9]) ? node32783 : node32776;
														assign node32776 = (inp[7]) ? node32780 : node32777;
															assign node32777 = (inp[8]) ? 4'b1111 : 4'b1110;
															assign node32780 = (inp[8]) ? 4'b1110 : 4'b1111;
														assign node32783 = (inp[14]) ? node32785 : 4'b1011;
															assign node32785 = (inp[7]) ? node32789 : node32786;
																assign node32786 = (inp[8]) ? 4'b1011 : 4'b1010;
																assign node32789 = (inp[8]) ? 4'b1010 : 4'b1011;
											assign node32792 = (inp[4]) ? node32830 : node32793;
												assign node32793 = (inp[9]) ? node32815 : node32794;
													assign node32794 = (inp[2]) ? node32804 : node32795;
														assign node32795 = (inp[8]) ? node32797 : 4'b1011;
															assign node32797 = (inp[7]) ? node32801 : node32798;
																assign node32798 = (inp[14]) ? 4'b1011 : 4'b1010;
																assign node32801 = (inp[14]) ? 4'b1010 : 4'b1011;
														assign node32804 = (inp[14]) ? node32810 : node32805;
															assign node32805 = (inp[7]) ? 4'b1010 : node32806;
																assign node32806 = (inp[8]) ? 4'b1011 : 4'b1010;
															assign node32810 = (inp[8]) ? 4'b1010 : node32811;
																assign node32811 = (inp[7]) ? 4'b1011 : 4'b1010;
													assign node32815 = (inp[2]) ? 4'b1101 : node32816;
														assign node32816 = (inp[14]) ? node32822 : node32817;
															assign node32817 = (inp[7]) ? 4'b1101 : node32818;
																assign node32818 = (inp[8]) ? 4'b1100 : 4'b1101;
															assign node32822 = (inp[7]) ? node32826 : node32823;
																assign node32823 = (inp[8]) ? 4'b1101 : 4'b1100;
																assign node32826 = (inp[8]) ? 4'b1100 : 4'b1101;
												assign node32830 = (inp[9]) ? node32852 : node32831;
													assign node32831 = (inp[2]) ? node32839 : node32832;
														assign node32832 = (inp[7]) ? 4'b1101 : node32833;
															assign node32833 = (inp[8]) ? node32835 : 4'b1101;
																assign node32835 = (inp[14]) ? 4'b1101 : 4'b1100;
														assign node32839 = (inp[14]) ? node32847 : node32840;
															assign node32840 = (inp[8]) ? node32844 : node32841;
																assign node32841 = (inp[7]) ? 4'b1101 : 4'b1100;
																assign node32844 = (inp[7]) ? 4'b1100 : 4'b1101;
															assign node32847 = (inp[8]) ? 4'b1101 : node32848;
																assign node32848 = (inp[7]) ? 4'b1101 : 4'b1100;
													assign node32852 = (inp[14]) ? node32854 : 4'b1000;
														assign node32854 = (inp[8]) ? node32858 : node32855;
															assign node32855 = (inp[7]) ? 4'b1001 : 4'b1000;
															assign node32858 = (inp[7]) ? 4'b1000 : 4'b1001;
								assign node32861 = (inp[0]) ? node33129 : node32862;
									assign node32862 = (inp[15]) ? node33022 : node32863;
										assign node32863 = (inp[5]) ? node32941 : node32864;
											assign node32864 = (inp[9]) ? node32906 : node32865;
												assign node32865 = (inp[4]) ? node32887 : node32866;
													assign node32866 = (inp[14]) ? node32880 : node32867;
														assign node32867 = (inp[2]) ? node32873 : node32868;
															assign node32868 = (inp[7]) ? 4'b1011 : node32869;
																assign node32869 = (inp[8]) ? 4'b1010 : 4'b1011;
															assign node32873 = (inp[7]) ? node32877 : node32874;
																assign node32874 = (inp[8]) ? 4'b1011 : 4'b1010;
																assign node32877 = (inp[8]) ? 4'b1010 : 4'b1011;
														assign node32880 = (inp[7]) ? node32884 : node32881;
															assign node32881 = (inp[8]) ? 4'b1011 : 4'b1010;
															assign node32884 = (inp[8]) ? 4'b1010 : 4'b1011;
													assign node32887 = (inp[2]) ? node32899 : node32888;
														assign node32888 = (inp[14]) ? node32894 : node32889;
															assign node32889 = (inp[7]) ? 4'b1101 : node32890;
																assign node32890 = (inp[8]) ? 4'b1100 : 4'b1101;
															assign node32894 = (inp[8]) ? node32896 : 4'b1100;
																assign node32896 = (inp[7]) ? 4'b1100 : 4'b1101;
														assign node32899 = (inp[8]) ? node32903 : node32900;
															assign node32900 = (inp[7]) ? 4'b1101 : 4'b1100;
															assign node32903 = (inp[7]) ? 4'b1100 : 4'b1101;
												assign node32906 = (inp[4]) ? node32924 : node32907;
													assign node32907 = (inp[2]) ? node32917 : node32908;
														assign node32908 = (inp[8]) ? node32910 : 4'b1100;
															assign node32910 = (inp[7]) ? node32914 : node32911;
																assign node32911 = (inp[14]) ? 4'b1101 : 4'b1100;
																assign node32914 = (inp[14]) ? 4'b1100 : 4'b1101;
														assign node32917 = (inp[8]) ? node32921 : node32918;
															assign node32918 = (inp[7]) ? 4'b1101 : 4'b1100;
															assign node32921 = (inp[7]) ? 4'b1100 : 4'b1101;
													assign node32924 = (inp[7]) ? node32934 : node32925;
														assign node32925 = (inp[14]) ? 4'b1000 : node32926;
															assign node32926 = (inp[2]) ? node32930 : node32927;
																assign node32927 = (inp[8]) ? 4'b1000 : 4'b1001;
																assign node32930 = (inp[8]) ? 4'b1001 : 4'b1000;
														assign node32934 = (inp[8]) ? node32938 : node32935;
															assign node32935 = (inp[14]) ? 4'b1001 : 4'b1000;
															assign node32938 = (inp[14]) ? 4'b1000 : 4'b1001;
											assign node32941 = (inp[14]) ? node32973 : node32942;
												assign node32942 = (inp[8]) ? node32958 : node32943;
													assign node32943 = (inp[4]) ? node32953 : node32944;
														assign node32944 = (inp[9]) ? node32946 : 4'b1000;
															assign node32946 = (inp[7]) ? node32950 : node32947;
																assign node32947 = (inp[2]) ? 4'b1100 : 4'b1101;
																assign node32950 = (inp[2]) ? 4'b1101 : 4'b1100;
														assign node32953 = (inp[9]) ? node32955 : 4'b1100;
															assign node32955 = (inp[7]) ? 4'b1001 : 4'b1000;
													assign node32958 = (inp[9]) ? node32966 : node32959;
														assign node32959 = (inp[4]) ? node32961 : 4'b1001;
															assign node32961 = (inp[7]) ? 4'b1100 : node32962;
																assign node32962 = (inp[2]) ? 4'b1101 : 4'b1100;
														assign node32966 = (inp[4]) ? 4'b1001 : node32967;
															assign node32967 = (inp[2]) ? 4'b1100 : node32968;
																assign node32968 = (inp[7]) ? 4'b1101 : 4'b1100;
												assign node32973 = (inp[4]) ? node32997 : node32974;
													assign node32974 = (inp[9]) ? node32988 : node32975;
														assign node32975 = (inp[2]) ? node32981 : node32976;
															assign node32976 = (inp[8]) ? 4'b1000 : node32977;
																assign node32977 = (inp[7]) ? 4'b1001 : 4'b1000;
															assign node32981 = (inp[7]) ? node32985 : node32982;
																assign node32982 = (inp[8]) ? 4'b1001 : 4'b1000;
																assign node32985 = (inp[8]) ? 4'b1000 : 4'b1001;
														assign node32988 = (inp[2]) ? node32990 : 4'b1100;
															assign node32990 = (inp[8]) ? node32994 : node32991;
																assign node32991 = (inp[7]) ? 4'b1101 : 4'b1100;
																assign node32994 = (inp[7]) ? 4'b1100 : 4'b1101;
													assign node32997 = (inp[9]) ? node33011 : node32998;
														assign node32998 = (inp[2]) ? node33006 : node32999;
															assign node32999 = (inp[7]) ? node33003 : node33000;
																assign node33000 = (inp[8]) ? 4'b1101 : 4'b1100;
																assign node33003 = (inp[8]) ? 4'b1100 : 4'b1101;
															assign node33006 = (inp[8]) ? 4'b1100 : node33007;
																assign node33007 = (inp[7]) ? 4'b1101 : 4'b1100;
														assign node33011 = (inp[2]) ? node33017 : node33012;
															assign node33012 = (inp[7]) ? 4'b1001 : node33013;
																assign node33013 = (inp[8]) ? 4'b1001 : 4'b1000;
															assign node33017 = (inp[8]) ? node33019 : 4'b1000;
																assign node33019 = (inp[7]) ? 4'b1000 : 4'b1001;
										assign node33022 = (inp[4]) ? node33072 : node33023;
											assign node33023 = (inp[9]) ? node33051 : node33024;
												assign node33024 = (inp[5]) ? node33034 : node33025;
													assign node33025 = (inp[8]) ? 4'b1001 : node33026;
														assign node33026 = (inp[7]) ? node33028 : 4'b1000;
															assign node33028 = (inp[14]) ? 4'b1001 : node33029;
																assign node33029 = (inp[2]) ? 4'b1001 : 4'b1000;
													assign node33034 = (inp[14]) ? node33044 : node33035;
														assign node33035 = (inp[7]) ? 4'b1010 : node33036;
															assign node33036 = (inp[2]) ? node33040 : node33037;
																assign node33037 = (inp[8]) ? 4'b1010 : 4'b1011;
																assign node33040 = (inp[8]) ? 4'b1011 : 4'b1010;
														assign node33044 = (inp[7]) ? node33048 : node33045;
															assign node33045 = (inp[8]) ? 4'b1011 : 4'b1010;
															assign node33048 = (inp[8]) ? 4'b1010 : 4'b1011;
												assign node33051 = (inp[8]) ? node33063 : node33052;
													assign node33052 = (inp[7]) ? node33058 : node33053;
														assign node33053 = (inp[14]) ? 4'b1110 : node33054;
															assign node33054 = (inp[2]) ? 4'b1110 : 4'b1111;
														assign node33058 = (inp[2]) ? 4'b1111 : node33059;
															assign node33059 = (inp[14]) ? 4'b1111 : 4'b1110;
													assign node33063 = (inp[7]) ? node33069 : node33064;
														assign node33064 = (inp[2]) ? 4'b1111 : node33065;
															assign node33065 = (inp[14]) ? 4'b1111 : 4'b1110;
														assign node33069 = (inp[2]) ? 4'b1110 : 4'b1111;
											assign node33072 = (inp[9]) ? node33104 : node33073;
												assign node33073 = (inp[2]) ? node33089 : node33074;
													assign node33074 = (inp[5]) ? 4'b1111 : node33075;
														assign node33075 = (inp[8]) ? node33081 : node33076;
															assign node33076 = (inp[14]) ? node33078 : 4'b1111;
																assign node33078 = (inp[7]) ? 4'b1111 : 4'b1110;
															assign node33081 = (inp[14]) ? node33085 : node33082;
																assign node33082 = (inp[7]) ? 4'b1111 : 4'b1110;
																assign node33085 = (inp[7]) ? 4'b1110 : 4'b1111;
													assign node33089 = (inp[14]) ? node33097 : node33090;
														assign node33090 = (inp[7]) ? node33094 : node33091;
															assign node33091 = (inp[8]) ? 4'b1111 : 4'b1110;
															assign node33094 = (inp[8]) ? 4'b1110 : 4'b1111;
														assign node33097 = (inp[7]) ? node33101 : node33098;
															assign node33098 = (inp[8]) ? 4'b1111 : 4'b1110;
															assign node33101 = (inp[8]) ? 4'b1110 : 4'b1111;
												assign node33104 = (inp[14]) ? node33122 : node33105;
													assign node33105 = (inp[7]) ? node33111 : node33106;
														assign node33106 = (inp[8]) ? 4'b1010 : node33107;
															assign node33107 = (inp[2]) ? 4'b1010 : 4'b1011;
														assign node33111 = (inp[5]) ? node33117 : node33112;
															assign node33112 = (inp[8]) ? node33114 : 4'b1010;
																assign node33114 = (inp[2]) ? 4'b1010 : 4'b1011;
															assign node33117 = (inp[8]) ? 4'b1011 : node33118;
																assign node33118 = (inp[2]) ? 4'b1011 : 4'b1010;
													assign node33122 = (inp[7]) ? node33126 : node33123;
														assign node33123 = (inp[8]) ? 4'b1011 : 4'b1010;
														assign node33126 = (inp[8]) ? 4'b1010 : 4'b1011;
									assign node33129 = (inp[15]) ? node33313 : node33130;
										assign node33130 = (inp[5]) ? node33212 : node33131;
											assign node33131 = (inp[4]) ? node33169 : node33132;
												assign node33132 = (inp[9]) ? node33156 : node33133;
													assign node33133 = (inp[2]) ? node33147 : node33134;
														assign node33134 = (inp[8]) ? node33140 : node33135;
															assign node33135 = (inp[14]) ? 4'b1001 : node33136;
																assign node33136 = (inp[7]) ? 4'b1000 : 4'b1001;
															assign node33140 = (inp[14]) ? node33144 : node33141;
																assign node33141 = (inp[7]) ? 4'b1001 : 4'b1000;
																assign node33144 = (inp[7]) ? 4'b1000 : 4'b1001;
														assign node33147 = (inp[14]) ? 4'b1000 : node33148;
															assign node33148 = (inp[8]) ? node33152 : node33149;
																assign node33149 = (inp[7]) ? 4'b1001 : 4'b1000;
																assign node33152 = (inp[7]) ? 4'b1000 : 4'b1001;
													assign node33156 = (inp[8]) ? node33162 : node33157;
														assign node33157 = (inp[7]) ? node33159 : 4'b1110;
															assign node33159 = (inp[14]) ? 4'b1111 : 4'b1110;
														assign node33162 = (inp[7]) ? node33166 : node33163;
															assign node33163 = (inp[14]) ? 4'b1111 : 4'b1110;
															assign node33166 = (inp[14]) ? 4'b1110 : 4'b1111;
												assign node33169 = (inp[9]) ? node33193 : node33170;
													assign node33170 = (inp[8]) ? node33182 : node33171;
														assign node33171 = (inp[7]) ? node33177 : node33172;
															assign node33172 = (inp[14]) ? 4'b1110 : node33173;
																assign node33173 = (inp[2]) ? 4'b1110 : 4'b1111;
															assign node33177 = (inp[2]) ? 4'b1111 : node33178;
																assign node33178 = (inp[14]) ? 4'b1111 : 4'b1110;
														assign node33182 = (inp[7]) ? node33188 : node33183;
															assign node33183 = (inp[2]) ? 4'b1111 : node33184;
																assign node33184 = (inp[14]) ? 4'b1111 : 4'b1110;
															assign node33188 = (inp[14]) ? 4'b1110 : node33189;
																assign node33189 = (inp[2]) ? 4'b1110 : 4'b1111;
													assign node33193 = (inp[14]) ? node33207 : node33194;
														assign node33194 = (inp[2]) ? node33202 : node33195;
															assign node33195 = (inp[8]) ? node33199 : node33196;
																assign node33196 = (inp[7]) ? 4'b1010 : 4'b1011;
																assign node33199 = (inp[7]) ? 4'b1011 : 4'b1010;
															assign node33202 = (inp[8]) ? node33204 : 4'b1011;
																assign node33204 = (inp[7]) ? 4'b1010 : 4'b1011;
														assign node33207 = (inp[8]) ? 4'b1010 : node33208;
															assign node33208 = (inp[7]) ? 4'b1011 : 4'b1010;
											assign node33212 = (inp[2]) ? node33272 : node33213;
												assign node33213 = (inp[7]) ? node33241 : node33214;
													assign node33214 = (inp[8]) ? node33226 : node33215;
														assign node33215 = (inp[14]) ? node33221 : node33216;
															assign node33216 = (inp[9]) ? 4'b1111 : node33217;
																assign node33217 = (inp[4]) ? 4'b1111 : 4'b1011;
															assign node33221 = (inp[9]) ? node33223 : 4'b1110;
																assign node33223 = (inp[4]) ? 4'b1010 : 4'b1110;
														assign node33226 = (inp[14]) ? node33234 : node33227;
															assign node33227 = (inp[4]) ? node33231 : node33228;
																assign node33228 = (inp[9]) ? 4'b1110 : 4'b1010;
																assign node33231 = (inp[9]) ? 4'b1010 : 4'b1110;
															assign node33234 = (inp[9]) ? node33238 : node33235;
																assign node33235 = (inp[4]) ? 4'b1111 : 4'b1011;
																assign node33238 = (inp[4]) ? 4'b1011 : 4'b1111;
													assign node33241 = (inp[4]) ? node33257 : node33242;
														assign node33242 = (inp[9]) ? node33250 : node33243;
															assign node33243 = (inp[14]) ? node33247 : node33244;
																assign node33244 = (inp[8]) ? 4'b1011 : 4'b1010;
																assign node33247 = (inp[8]) ? 4'b1010 : 4'b1011;
															assign node33250 = (inp[8]) ? node33254 : node33251;
																assign node33251 = (inp[14]) ? 4'b1111 : 4'b1110;
																assign node33254 = (inp[14]) ? 4'b1110 : 4'b1111;
														assign node33257 = (inp[9]) ? node33265 : node33258;
															assign node33258 = (inp[14]) ? node33262 : node33259;
																assign node33259 = (inp[8]) ? 4'b1111 : 4'b1110;
																assign node33262 = (inp[8]) ? 4'b1110 : 4'b1111;
															assign node33265 = (inp[14]) ? node33269 : node33266;
																assign node33266 = (inp[8]) ? 4'b1011 : 4'b1010;
																assign node33269 = (inp[8]) ? 4'b1010 : 4'b1011;
												assign node33272 = (inp[14]) ? node33294 : node33273;
													assign node33273 = (inp[9]) ? node33281 : node33274;
														assign node33274 = (inp[4]) ? 4'b1111 : node33275;
															assign node33275 = (inp[7]) ? node33277 : 4'b1011;
																assign node33277 = (inp[8]) ? 4'b1010 : 4'b1011;
														assign node33281 = (inp[4]) ? node33287 : node33282;
															assign node33282 = (inp[7]) ? 4'b1110 : node33283;
																assign node33283 = (inp[8]) ? 4'b1111 : 4'b1110;
															assign node33287 = (inp[7]) ? node33291 : node33288;
																assign node33288 = (inp[8]) ? 4'b1011 : 4'b1010;
																assign node33291 = (inp[8]) ? 4'b1010 : 4'b1011;
													assign node33294 = (inp[7]) ? node33302 : node33295;
														assign node33295 = (inp[8]) ? 4'b1011 : node33296;
															assign node33296 = (inp[9]) ? node33298 : 4'b1010;
																assign node33298 = (inp[4]) ? 4'b1010 : 4'b1110;
														assign node33302 = (inp[8]) ? node33306 : node33303;
															assign node33303 = (inp[4]) ? 4'b1111 : 4'b1011;
															assign node33306 = (inp[9]) ? node33310 : node33307;
																assign node33307 = (inp[4]) ? 4'b1110 : 4'b1010;
																assign node33310 = (inp[4]) ? 4'b1010 : 4'b1110;
										assign node33313 = (inp[4]) ? node33385 : node33314;
											assign node33314 = (inp[9]) ? node33358 : node33315;
												assign node33315 = (inp[5]) ? node33333 : node33316;
													assign node33316 = (inp[2]) ? node33326 : node33317;
														assign node33317 = (inp[8]) ? node33319 : 4'b1010;
															assign node33319 = (inp[14]) ? node33323 : node33320;
																assign node33320 = (inp[7]) ? 4'b1011 : 4'b1010;
																assign node33323 = (inp[7]) ? 4'b1010 : 4'b1011;
														assign node33326 = (inp[7]) ? node33330 : node33327;
															assign node33327 = (inp[8]) ? 4'b1011 : 4'b1010;
															assign node33330 = (inp[8]) ? 4'b1010 : 4'b1011;
													assign node33333 = (inp[2]) ? node33349 : node33334;
														assign node33334 = (inp[8]) ? node33342 : node33335;
															assign node33335 = (inp[7]) ? node33339 : node33336;
																assign node33336 = (inp[14]) ? 4'b1000 : 4'b1001;
																assign node33339 = (inp[14]) ? 4'b1001 : 4'b1000;
															assign node33342 = (inp[7]) ? node33346 : node33343;
																assign node33343 = (inp[14]) ? 4'b1001 : 4'b1000;
																assign node33346 = (inp[14]) ? 4'b1000 : 4'b1001;
														assign node33349 = (inp[14]) ? node33353 : node33350;
															assign node33350 = (inp[7]) ? 4'b1001 : 4'b1000;
															assign node33353 = (inp[7]) ? node33355 : 4'b1001;
																assign node33355 = (inp[8]) ? 4'b1000 : 4'b1001;
												assign node33358 = (inp[5]) ? node33376 : node33359;
													assign node33359 = (inp[14]) ? node33369 : node33360;
														assign node33360 = (inp[7]) ? node33362 : 4'b1101;
															assign node33362 = (inp[2]) ? node33366 : node33363;
																assign node33363 = (inp[8]) ? 4'b1101 : 4'b1100;
																assign node33366 = (inp[8]) ? 4'b1100 : 4'b1101;
														assign node33369 = (inp[8]) ? node33373 : node33370;
															assign node33370 = (inp[7]) ? 4'b1101 : 4'b1100;
															assign node33373 = (inp[7]) ? 4'b1100 : 4'b1101;
													assign node33376 = (inp[14]) ? node33378 : 4'b1100;
														assign node33378 = (inp[8]) ? node33382 : node33379;
															assign node33379 = (inp[7]) ? 4'b1101 : 4'b1100;
															assign node33382 = (inp[7]) ? 4'b1100 : 4'b1101;
											assign node33385 = (inp[9]) ? node33409 : node33386;
												assign node33386 = (inp[14]) ? node33402 : node33387;
													assign node33387 = (inp[7]) ? node33395 : node33388;
														assign node33388 = (inp[2]) ? node33392 : node33389;
															assign node33389 = (inp[8]) ? 4'b1100 : 4'b1101;
															assign node33392 = (inp[8]) ? 4'b1101 : 4'b1100;
														assign node33395 = (inp[2]) ? node33399 : node33396;
															assign node33396 = (inp[8]) ? 4'b1101 : 4'b1100;
															assign node33399 = (inp[8]) ? 4'b1100 : 4'b1101;
													assign node33402 = (inp[7]) ? node33406 : node33403;
														assign node33403 = (inp[8]) ? 4'b1101 : 4'b1100;
														assign node33406 = (inp[8]) ? 4'b1100 : 4'b1101;
												assign node33409 = (inp[2]) ? node33423 : node33410;
													assign node33410 = (inp[14]) ? 4'b1000 : node33411;
														assign node33411 = (inp[5]) ? node33417 : node33412;
															assign node33412 = (inp[8]) ? 4'b1000 : node33413;
																assign node33413 = (inp[7]) ? 4'b1000 : 4'b1001;
															assign node33417 = (inp[8]) ? node33419 : 4'b1000;
																assign node33419 = (inp[7]) ? 4'b1001 : 4'b1000;
													assign node33423 = (inp[8]) ? node33427 : node33424;
														assign node33424 = (inp[7]) ? 4'b1001 : 4'b1000;
														assign node33427 = (inp[7]) ? 4'b1000 : 4'b1001;
		assign node33430 = (inp[11]) ? node49852 : node33431;
			assign node33431 = (inp[13]) ? node41539 : node33432;
				assign node33432 = (inp[1]) ? node37382 : node33433;
					assign node33433 = (inp[12]) ? node35081 : node33434;
						assign node33434 = (inp[8]) ? node34176 : node33435;
							assign node33435 = (inp[7]) ? node33837 : node33436;
								assign node33436 = (inp[14]) ? node33702 : node33437;
									assign node33437 = (inp[2]) ? node33567 : node33438;
										assign node33438 = (inp[0]) ? node33500 : node33439;
											assign node33439 = (inp[15]) ? node33463 : node33440;
												assign node33440 = (inp[5]) ? node33450 : node33441;
													assign node33441 = (inp[9]) ? node33445 : node33442;
														assign node33442 = (inp[4]) ? 4'b0011 : 4'b0111;
														assign node33445 = (inp[4]) ? node33447 : 4'b0011;
															assign node33447 = (inp[3]) ? 4'b0101 : 4'b0111;
													assign node33450 = (inp[3]) ? node33456 : node33451;
														assign node33451 = (inp[9]) ? 4'b0101 : node33452;
															assign node33452 = (inp[4]) ? 4'b0011 : 4'b0111;
														assign node33456 = (inp[10]) ? 4'b0101 : node33457;
															assign node33457 = (inp[9]) ? node33459 : 4'b0101;
																assign node33459 = (inp[4]) ? 4'b0101 : 4'b0001;
												assign node33463 = (inp[5]) ? node33481 : node33464;
													assign node33464 = (inp[3]) ? node33474 : node33465;
														assign node33465 = (inp[10]) ? 4'b0001 : node33466;
															assign node33466 = (inp[9]) ? node33470 : node33467;
																assign node33467 = (inp[4]) ? 4'b0001 : 4'b0101;
																assign node33470 = (inp[4]) ? 4'b0101 : 4'b0001;
														assign node33474 = (inp[9]) ? node33478 : node33475;
															assign node33475 = (inp[4]) ? 4'b0001 : 4'b0101;
															assign node33478 = (inp[4]) ? 4'b0111 : 4'b0001;
													assign node33481 = (inp[3]) ? node33487 : node33482;
														assign node33482 = (inp[4]) ? 4'b0111 : node33483;
															assign node33483 = (inp[9]) ? 4'b0001 : 4'b0101;
														assign node33487 = (inp[10]) ? node33495 : node33488;
															assign node33488 = (inp[4]) ? node33492 : node33489;
																assign node33489 = (inp[9]) ? 4'b0011 : 4'b0111;
																assign node33492 = (inp[9]) ? 4'b0111 : 4'b0011;
															assign node33495 = (inp[9]) ? node33497 : 4'b0011;
																assign node33497 = (inp[4]) ? 4'b0111 : 4'b0011;
											assign node33500 = (inp[15]) ? node33534 : node33501;
												assign node33501 = (inp[3]) ? node33519 : node33502;
													assign node33502 = (inp[5]) ? node33510 : node33503;
														assign node33503 = (inp[9]) ? node33507 : node33504;
															assign node33504 = (inp[4]) ? 4'b0001 : 4'b0101;
															assign node33507 = (inp[4]) ? 4'b0101 : 4'b0001;
														assign node33510 = (inp[10]) ? node33512 : 4'b0001;
															assign node33512 = (inp[9]) ? node33516 : node33513;
																assign node33513 = (inp[4]) ? 4'b0001 : 4'b0101;
																assign node33516 = (inp[4]) ? 4'b0111 : 4'b0001;
													assign node33519 = (inp[5]) ? node33527 : node33520;
														assign node33520 = (inp[9]) ? node33524 : node33521;
															assign node33521 = (inp[4]) ? 4'b0001 : 4'b0101;
															assign node33524 = (inp[4]) ? 4'b0111 : 4'b0001;
														assign node33527 = (inp[9]) ? node33531 : node33528;
															assign node33528 = (inp[4]) ? 4'b0011 : 4'b0111;
															assign node33531 = (inp[4]) ? 4'b0111 : 4'b0011;
												assign node33534 = (inp[3]) ? node33544 : node33535;
													assign node33535 = (inp[9]) ? node33539 : node33536;
														assign node33536 = (inp[4]) ? 4'b0011 : 4'b0111;
														assign node33539 = (inp[4]) ? node33541 : 4'b0011;
															assign node33541 = (inp[5]) ? 4'b0101 : 4'b0111;
													assign node33544 = (inp[5]) ? node33554 : node33545;
														assign node33545 = (inp[10]) ? node33551 : node33546;
															assign node33546 = (inp[9]) ? 4'b0011 : node33547;
																assign node33547 = (inp[4]) ? 4'b0011 : 4'b0111;
															assign node33551 = (inp[4]) ? 4'b0101 : 4'b0111;
														assign node33554 = (inp[10]) ? node33562 : node33555;
															assign node33555 = (inp[9]) ? node33559 : node33556;
																assign node33556 = (inp[4]) ? 4'b0001 : 4'b0101;
																assign node33559 = (inp[4]) ? 4'b0101 : 4'b0001;
															assign node33562 = (inp[9]) ? 4'b0001 : node33563;
																assign node33563 = (inp[4]) ? 4'b0001 : 4'b0101;
										assign node33567 = (inp[5]) ? node33621 : node33568;
											assign node33568 = (inp[0]) ? node33594 : node33569;
												assign node33569 = (inp[15]) ? node33585 : node33570;
													assign node33570 = (inp[3]) ? node33578 : node33571;
														assign node33571 = (inp[4]) ? node33575 : node33572;
															assign node33572 = (inp[9]) ? 4'b0010 : 4'b0110;
															assign node33575 = (inp[9]) ? 4'b0110 : 4'b0010;
														assign node33578 = (inp[4]) ? node33582 : node33579;
															assign node33579 = (inp[9]) ? 4'b0010 : 4'b0110;
															assign node33582 = (inp[10]) ? 4'b0010 : 4'b0100;
													assign node33585 = (inp[4]) ? node33589 : node33586;
														assign node33586 = (inp[9]) ? 4'b0000 : 4'b0100;
														assign node33589 = (inp[9]) ? node33591 : 4'b0000;
															assign node33591 = (inp[3]) ? 4'b0110 : 4'b0100;
												assign node33594 = (inp[15]) ? node33614 : node33595;
													assign node33595 = (inp[3]) ? node33603 : node33596;
														assign node33596 = (inp[4]) ? node33600 : node33597;
															assign node33597 = (inp[9]) ? 4'b0000 : 4'b0100;
															assign node33600 = (inp[9]) ? 4'b0100 : 4'b0000;
														assign node33603 = (inp[10]) ? node33609 : node33604;
															assign node33604 = (inp[4]) ? node33606 : 4'b0000;
																assign node33606 = (inp[9]) ? 4'b0110 : 4'b0000;
															assign node33609 = (inp[9]) ? 4'b0000 : node33610;
																assign node33610 = (inp[4]) ? 4'b0000 : 4'b0100;
													assign node33614 = (inp[9]) ? node33618 : node33615;
														assign node33615 = (inp[4]) ? 4'b0010 : 4'b0110;
														assign node33618 = (inp[4]) ? 4'b0100 : 4'b0010;
											assign node33621 = (inp[10]) ? node33665 : node33622;
												assign node33622 = (inp[0]) ? node33650 : node33623;
													assign node33623 = (inp[15]) ? node33635 : node33624;
														assign node33624 = (inp[3]) ? node33630 : node33625;
															assign node33625 = (inp[9]) ? 4'b0100 : node33626;
																assign node33626 = (inp[4]) ? 4'b0010 : 4'b0110;
															assign node33630 = (inp[9]) ? 4'b0000 : node33631;
																assign node33631 = (inp[4]) ? 4'b0000 : 4'b0100;
														assign node33635 = (inp[3]) ? node33643 : node33636;
															assign node33636 = (inp[4]) ? node33640 : node33637;
																assign node33637 = (inp[9]) ? 4'b0000 : 4'b0100;
																assign node33640 = (inp[9]) ? 4'b0110 : 4'b0000;
															assign node33643 = (inp[9]) ? node33647 : node33644;
																assign node33644 = (inp[4]) ? 4'b0010 : 4'b0110;
																assign node33647 = (inp[4]) ? 4'b0110 : 4'b0010;
													assign node33650 = (inp[15]) ? node33654 : node33651;
														assign node33651 = (inp[9]) ? 4'b0110 : 4'b0010;
														assign node33654 = (inp[3]) ? node33660 : node33655;
															assign node33655 = (inp[4]) ? 4'b0100 : node33656;
																assign node33656 = (inp[9]) ? 4'b0010 : 4'b0110;
															assign node33660 = (inp[4]) ? node33662 : 4'b0100;
																assign node33662 = (inp[9]) ? 4'b0100 : 4'b0000;
												assign node33665 = (inp[3]) ? node33687 : node33666;
													assign node33666 = (inp[0]) ? node33678 : node33667;
														assign node33667 = (inp[9]) ? node33671 : node33668;
															assign node33668 = (inp[4]) ? 4'b0000 : 4'b0100;
															assign node33671 = (inp[4]) ? node33675 : node33672;
																assign node33672 = (inp[15]) ? 4'b0000 : 4'b0010;
																assign node33675 = (inp[15]) ? 4'b0110 : 4'b0100;
														assign node33678 = (inp[15]) ? node33684 : node33679;
															assign node33679 = (inp[9]) ? node33681 : 4'b0000;
																assign node33681 = (inp[4]) ? 4'b0110 : 4'b0000;
															assign node33684 = (inp[4]) ? 4'b0010 : 4'b0110;
													assign node33687 = (inp[15]) ? node33695 : node33688;
														assign node33688 = (inp[0]) ? node33690 : 4'b0000;
															assign node33690 = (inp[4]) ? 4'b0110 : node33691;
																assign node33691 = (inp[9]) ? 4'b0010 : 4'b0110;
														assign node33695 = (inp[0]) ? 4'b0000 : node33696;
															assign node33696 = (inp[9]) ? node33698 : 4'b0010;
																assign node33698 = (inp[4]) ? 4'b0110 : 4'b0010;
									assign node33702 = (inp[0]) ? node33780 : node33703;
										assign node33703 = (inp[15]) ? node33749 : node33704;
											assign node33704 = (inp[5]) ? node33714 : node33705;
												assign node33705 = (inp[4]) ? node33709 : node33706;
													assign node33706 = (inp[9]) ? 4'b0010 : 4'b0110;
													assign node33709 = (inp[9]) ? node33711 : 4'b0010;
														assign node33711 = (inp[3]) ? 4'b0100 : 4'b0110;
												assign node33714 = (inp[3]) ? node33722 : node33715;
													assign node33715 = (inp[9]) ? node33719 : node33716;
														assign node33716 = (inp[4]) ? 4'b0010 : 4'b0110;
														assign node33719 = (inp[4]) ? 4'b0100 : 4'b0010;
													assign node33722 = (inp[10]) ? node33736 : node33723;
														assign node33723 = (inp[2]) ? node33731 : node33724;
															assign node33724 = (inp[9]) ? node33728 : node33725;
																assign node33725 = (inp[4]) ? 4'b0000 : 4'b0100;
																assign node33728 = (inp[4]) ? 4'b0100 : 4'b0000;
															assign node33731 = (inp[4]) ? 4'b0000 : node33732;
																assign node33732 = (inp[9]) ? 4'b0000 : 4'b0100;
														assign node33736 = (inp[2]) ? node33742 : node33737;
															assign node33737 = (inp[9]) ? node33739 : 4'b0100;
																assign node33739 = (inp[4]) ? 4'b0100 : 4'b0000;
															assign node33742 = (inp[4]) ? node33746 : node33743;
																assign node33743 = (inp[9]) ? 4'b0000 : 4'b0100;
																assign node33746 = (inp[9]) ? 4'b0100 : 4'b0000;
											assign node33749 = (inp[5]) ? node33759 : node33750;
												assign node33750 = (inp[4]) ? node33754 : node33751;
													assign node33751 = (inp[9]) ? 4'b0000 : 4'b0100;
													assign node33754 = (inp[9]) ? node33756 : 4'b0000;
														assign node33756 = (inp[3]) ? 4'b0110 : 4'b0100;
												assign node33759 = (inp[3]) ? node33767 : node33760;
													assign node33760 = (inp[9]) ? node33764 : node33761;
														assign node33761 = (inp[4]) ? 4'b0000 : 4'b0100;
														assign node33764 = (inp[4]) ? 4'b0110 : 4'b0000;
													assign node33767 = (inp[2]) ? node33773 : node33768;
														assign node33768 = (inp[9]) ? 4'b0010 : node33769;
															assign node33769 = (inp[4]) ? 4'b0010 : 4'b0110;
														assign node33773 = (inp[9]) ? node33777 : node33774;
															assign node33774 = (inp[4]) ? 4'b0010 : 4'b0110;
															assign node33777 = (inp[4]) ? 4'b0110 : 4'b0010;
										assign node33780 = (inp[15]) ? node33812 : node33781;
											assign node33781 = (inp[3]) ? node33797 : node33782;
												assign node33782 = (inp[5]) ? node33790 : node33783;
													assign node33783 = (inp[9]) ? node33787 : node33784;
														assign node33784 = (inp[4]) ? 4'b0000 : 4'b0100;
														assign node33787 = (inp[4]) ? 4'b0100 : 4'b0000;
													assign node33790 = (inp[4]) ? node33794 : node33791;
														assign node33791 = (inp[9]) ? 4'b0000 : 4'b0100;
														assign node33794 = (inp[9]) ? 4'b0110 : 4'b0000;
												assign node33797 = (inp[5]) ? node33805 : node33798;
													assign node33798 = (inp[4]) ? node33802 : node33799;
														assign node33799 = (inp[9]) ? 4'b0000 : 4'b0100;
														assign node33802 = (inp[9]) ? 4'b0110 : 4'b0000;
													assign node33805 = (inp[2]) ? 4'b0110 : node33806;
														assign node33806 = (inp[9]) ? 4'b0110 : node33807;
															assign node33807 = (inp[4]) ? 4'b0010 : 4'b0110;
											assign node33812 = (inp[3]) ? node33822 : node33813;
												assign node33813 = (inp[4]) ? node33817 : node33814;
													assign node33814 = (inp[9]) ? 4'b0010 : 4'b0110;
													assign node33817 = (inp[9]) ? node33819 : 4'b0010;
														assign node33819 = (inp[5]) ? 4'b0100 : 4'b0110;
												assign node33822 = (inp[5]) ? node33830 : node33823;
													assign node33823 = (inp[9]) ? node33827 : node33824;
														assign node33824 = (inp[4]) ? 4'b0010 : 4'b0110;
														assign node33827 = (inp[4]) ? 4'b0100 : 4'b0010;
													assign node33830 = (inp[4]) ? node33834 : node33831;
														assign node33831 = (inp[9]) ? 4'b0000 : 4'b0100;
														assign node33834 = (inp[9]) ? 4'b0100 : 4'b0000;
								assign node33837 = (inp[2]) ? node34059 : node33838;
									assign node33838 = (inp[14]) ? node33946 : node33839;
										assign node33839 = (inp[0]) ? node33885 : node33840;
											assign node33840 = (inp[15]) ? node33862 : node33841;
												assign node33841 = (inp[5]) ? node33849 : node33842;
													assign node33842 = (inp[9]) ? node33846 : node33843;
														assign node33843 = (inp[4]) ? 4'b0010 : 4'b0110;
														assign node33846 = (inp[4]) ? 4'b0110 : 4'b0010;
													assign node33849 = (inp[3]) ? node33855 : node33850;
														assign node33850 = (inp[4]) ? 4'b0100 : node33851;
															assign node33851 = (inp[9]) ? 4'b0010 : 4'b0110;
														assign node33855 = (inp[9]) ? node33859 : node33856;
															assign node33856 = (inp[4]) ? 4'b0000 : 4'b0100;
															assign node33859 = (inp[4]) ? 4'b0100 : 4'b0000;
												assign node33862 = (inp[3]) ? node33872 : node33863;
													assign node33863 = (inp[9]) ? node33867 : node33864;
														assign node33864 = (inp[4]) ? 4'b0000 : 4'b0100;
														assign node33867 = (inp[4]) ? node33869 : 4'b0000;
															assign node33869 = (inp[5]) ? 4'b0110 : 4'b0100;
													assign node33872 = (inp[5]) ? node33878 : node33873;
														assign node33873 = (inp[9]) ? 4'b0110 : node33874;
															assign node33874 = (inp[4]) ? 4'b0000 : 4'b0100;
														assign node33878 = (inp[4]) ? node33882 : node33879;
															assign node33879 = (inp[9]) ? 4'b0010 : 4'b0110;
															assign node33882 = (inp[9]) ? 4'b0110 : 4'b0010;
											assign node33885 = (inp[15]) ? node33921 : node33886;
												assign node33886 = (inp[3]) ? node33902 : node33887;
													assign node33887 = (inp[5]) ? node33895 : node33888;
														assign node33888 = (inp[9]) ? node33892 : node33889;
															assign node33889 = (inp[4]) ? 4'b0000 : 4'b0100;
															assign node33892 = (inp[4]) ? 4'b0100 : 4'b0000;
														assign node33895 = (inp[4]) ? node33899 : node33896;
															assign node33896 = (inp[9]) ? 4'b0000 : 4'b0100;
															assign node33899 = (inp[9]) ? 4'b0110 : 4'b0000;
													assign node33902 = (inp[5]) ? node33910 : node33903;
														assign node33903 = (inp[9]) ? node33907 : node33904;
															assign node33904 = (inp[4]) ? 4'b0000 : 4'b0100;
															assign node33907 = (inp[4]) ? 4'b0110 : 4'b0000;
														assign node33910 = (inp[10]) ? node33916 : node33911;
															assign node33911 = (inp[9]) ? node33913 : 4'b0010;
																assign node33913 = (inp[4]) ? 4'b0110 : 4'b0010;
															assign node33916 = (inp[9]) ? 4'b0010 : node33917;
																assign node33917 = (inp[4]) ? 4'b0010 : 4'b0110;
												assign node33921 = (inp[5]) ? node33931 : node33922;
													assign node33922 = (inp[4]) ? node33926 : node33923;
														assign node33923 = (inp[9]) ? 4'b0010 : 4'b0110;
														assign node33926 = (inp[9]) ? node33928 : 4'b0010;
															assign node33928 = (inp[10]) ? 4'b0110 : 4'b0100;
													assign node33931 = (inp[3]) ? node33939 : node33932;
														assign node33932 = (inp[9]) ? node33936 : node33933;
															assign node33933 = (inp[4]) ? 4'b0010 : 4'b0110;
															assign node33936 = (inp[4]) ? 4'b0100 : 4'b0010;
														assign node33939 = (inp[9]) ? node33943 : node33940;
															assign node33940 = (inp[4]) ? 4'b0000 : 4'b0100;
															assign node33943 = (inp[4]) ? 4'b0100 : 4'b0000;
										assign node33946 = (inp[5]) ? node33986 : node33947;
											assign node33947 = (inp[0]) ? node33967 : node33948;
												assign node33948 = (inp[15]) ? node33958 : node33949;
													assign node33949 = (inp[4]) ? node33953 : node33950;
														assign node33950 = (inp[9]) ? 4'b0011 : 4'b0111;
														assign node33953 = (inp[9]) ? node33955 : 4'b0011;
															assign node33955 = (inp[3]) ? 4'b0101 : 4'b0111;
													assign node33958 = (inp[9]) ? node33962 : node33959;
														assign node33959 = (inp[4]) ? 4'b0001 : 4'b0101;
														assign node33962 = (inp[4]) ? node33964 : 4'b0001;
															assign node33964 = (inp[3]) ? 4'b0111 : 4'b0101;
												assign node33967 = (inp[15]) ? node33977 : node33968;
													assign node33968 = (inp[4]) ? node33972 : node33969;
														assign node33969 = (inp[9]) ? 4'b0001 : 4'b0101;
														assign node33972 = (inp[3]) ? 4'b0111 : node33973;
															assign node33973 = (inp[10]) ? 4'b0101 : 4'b0001;
													assign node33977 = (inp[9]) ? node33981 : node33978;
														assign node33978 = (inp[4]) ? 4'b0011 : 4'b0111;
														assign node33981 = (inp[4]) ? node33983 : 4'b0011;
															assign node33983 = (inp[3]) ? 4'b0101 : 4'b0111;
											assign node33986 = (inp[4]) ? node34024 : node33987;
												assign node33987 = (inp[9]) ? node34001 : node33988;
													assign node33988 = (inp[10]) ? node33996 : node33989;
														assign node33989 = (inp[15]) ? node33991 : 4'b0111;
															assign node33991 = (inp[3]) ? 4'b0101 : node33992;
																assign node33992 = (inp[0]) ? 4'b0111 : 4'b0101;
														assign node33996 = (inp[3]) ? 4'b0101 : node33997;
															assign node33997 = (inp[0]) ? 4'b0101 : 4'b0111;
													assign node34001 = (inp[3]) ? node34009 : node34002;
														assign node34002 = (inp[15]) ? node34006 : node34003;
															assign node34003 = (inp[0]) ? 4'b0001 : 4'b0011;
															assign node34006 = (inp[0]) ? 4'b0011 : 4'b0001;
														assign node34009 = (inp[10]) ? node34017 : node34010;
															assign node34010 = (inp[15]) ? node34014 : node34011;
																assign node34011 = (inp[0]) ? 4'b0011 : 4'b0001;
																assign node34014 = (inp[0]) ? 4'b0001 : 4'b0011;
															assign node34017 = (inp[0]) ? node34021 : node34018;
																assign node34018 = (inp[15]) ? 4'b0011 : 4'b0001;
																assign node34021 = (inp[15]) ? 4'b0001 : 4'b0011;
												assign node34024 = (inp[9]) ? node34044 : node34025;
													assign node34025 = (inp[3]) ? node34031 : node34026;
														assign node34026 = (inp[15]) ? 4'b0001 : node34027;
															assign node34027 = (inp[0]) ? 4'b0001 : 4'b0011;
														assign node34031 = (inp[10]) ? node34039 : node34032;
															assign node34032 = (inp[15]) ? node34036 : node34033;
																assign node34033 = (inp[0]) ? 4'b0011 : 4'b0001;
																assign node34036 = (inp[0]) ? 4'b0001 : 4'b0011;
															assign node34039 = (inp[15]) ? 4'b0011 : node34040;
																assign node34040 = (inp[0]) ? 4'b0011 : 4'b0001;
													assign node34044 = (inp[3]) ? node34052 : node34045;
														assign node34045 = (inp[15]) ? node34049 : node34046;
															assign node34046 = (inp[0]) ? 4'b0111 : 4'b0101;
															assign node34049 = (inp[0]) ? 4'b0101 : 4'b0111;
														assign node34052 = (inp[0]) ? node34056 : node34053;
															assign node34053 = (inp[15]) ? 4'b0111 : 4'b0101;
															assign node34056 = (inp[15]) ? 4'b0101 : 4'b0111;
									assign node34059 = (inp[15]) ? node34117 : node34060;
										assign node34060 = (inp[0]) ? node34086 : node34061;
											assign node34061 = (inp[3]) ? node34071 : node34062;
												assign node34062 = (inp[4]) ? node34066 : node34063;
													assign node34063 = (inp[9]) ? 4'b0011 : 4'b0111;
													assign node34066 = (inp[9]) ? node34068 : 4'b0011;
														assign node34068 = (inp[5]) ? 4'b0101 : 4'b0111;
												assign node34071 = (inp[5]) ? node34079 : node34072;
													assign node34072 = (inp[4]) ? node34076 : node34073;
														assign node34073 = (inp[9]) ? 4'b0011 : 4'b0111;
														assign node34076 = (inp[9]) ? 4'b0101 : 4'b0011;
													assign node34079 = (inp[9]) ? node34083 : node34080;
														assign node34080 = (inp[4]) ? 4'b0001 : 4'b0101;
														assign node34083 = (inp[4]) ? 4'b0101 : 4'b0001;
											assign node34086 = (inp[5]) ? node34096 : node34087;
												assign node34087 = (inp[4]) ? node34091 : node34088;
													assign node34088 = (inp[9]) ? 4'b0001 : 4'b0101;
													assign node34091 = (inp[9]) ? node34093 : 4'b0001;
														assign node34093 = (inp[3]) ? 4'b0111 : 4'b0101;
												assign node34096 = (inp[3]) ? node34104 : node34097;
													assign node34097 = (inp[9]) ? node34101 : node34098;
														assign node34098 = (inp[4]) ? 4'b0001 : 4'b0101;
														assign node34101 = (inp[4]) ? 4'b0111 : 4'b0001;
													assign node34104 = (inp[10]) ? node34112 : node34105;
														assign node34105 = (inp[9]) ? node34109 : node34106;
															assign node34106 = (inp[4]) ? 4'b0011 : 4'b0111;
															assign node34109 = (inp[4]) ? 4'b0111 : 4'b0011;
														assign node34112 = (inp[9]) ? 4'b0011 : node34113;
															assign node34113 = (inp[4]) ? 4'b0011 : 4'b0111;
										assign node34117 = (inp[0]) ? node34151 : node34118;
											assign node34118 = (inp[3]) ? node34128 : node34119;
												assign node34119 = (inp[4]) ? node34123 : node34120;
													assign node34120 = (inp[9]) ? 4'b0001 : 4'b0101;
													assign node34123 = (inp[9]) ? node34125 : 4'b0001;
														assign node34125 = (inp[5]) ? 4'b0111 : 4'b0101;
												assign node34128 = (inp[5]) ? node34136 : node34129;
													assign node34129 = (inp[9]) ? node34133 : node34130;
														assign node34130 = (inp[4]) ? 4'b0001 : 4'b0101;
														assign node34133 = (inp[4]) ? 4'b0111 : 4'b0001;
													assign node34136 = (inp[10]) ? node34144 : node34137;
														assign node34137 = (inp[9]) ? node34141 : node34138;
															assign node34138 = (inp[4]) ? 4'b0011 : 4'b0111;
															assign node34141 = (inp[4]) ? 4'b0111 : 4'b0011;
														assign node34144 = (inp[14]) ? node34146 : 4'b0011;
															assign node34146 = (inp[9]) ? 4'b0011 : node34147;
																assign node34147 = (inp[4]) ? 4'b0011 : 4'b0111;
											assign node34151 = (inp[5]) ? node34161 : node34152;
												assign node34152 = (inp[9]) ? node34156 : node34153;
													assign node34153 = (inp[4]) ? 4'b0011 : 4'b0111;
													assign node34156 = (inp[4]) ? node34158 : 4'b0011;
														assign node34158 = (inp[3]) ? 4'b0101 : 4'b0111;
												assign node34161 = (inp[3]) ? node34169 : node34162;
													assign node34162 = (inp[4]) ? node34166 : node34163;
														assign node34163 = (inp[9]) ? 4'b0011 : 4'b0111;
														assign node34166 = (inp[9]) ? 4'b0101 : 4'b0011;
													assign node34169 = (inp[4]) ? node34173 : node34170;
														assign node34170 = (inp[9]) ? 4'b0001 : 4'b0101;
														assign node34173 = (inp[9]) ? 4'b0101 : 4'b0001;
							assign node34176 = (inp[7]) ? node34708 : node34177;
								assign node34177 = (inp[2]) ? node34419 : node34178;
									assign node34178 = (inp[14]) ? node34272 : node34179;
										assign node34179 = (inp[15]) ? node34237 : node34180;
											assign node34180 = (inp[0]) ? node34214 : node34181;
												assign node34181 = (inp[3]) ? node34195 : node34182;
													assign node34182 = (inp[5]) ? node34188 : node34183;
														assign node34183 = (inp[4]) ? 4'b0010 : node34184;
															assign node34184 = (inp[9]) ? 4'b0010 : 4'b0110;
														assign node34188 = (inp[4]) ? node34192 : node34189;
															assign node34189 = (inp[9]) ? 4'b0010 : 4'b0110;
															assign node34192 = (inp[9]) ? 4'b0100 : 4'b0010;
													assign node34195 = (inp[5]) ? node34201 : node34196;
														assign node34196 = (inp[9]) ? node34198 : 4'b0010;
															assign node34198 = (inp[4]) ? 4'b0100 : 4'b0010;
														assign node34201 = (inp[10]) ? node34207 : node34202;
															assign node34202 = (inp[9]) ? 4'b0100 : node34203;
																assign node34203 = (inp[4]) ? 4'b0000 : 4'b0100;
															assign node34207 = (inp[9]) ? node34211 : node34208;
																assign node34208 = (inp[4]) ? 4'b0000 : 4'b0100;
																assign node34211 = (inp[4]) ? 4'b0100 : 4'b0000;
												assign node34214 = (inp[3]) ? node34224 : node34215;
													assign node34215 = (inp[4]) ? node34219 : node34216;
														assign node34216 = (inp[9]) ? 4'b0000 : 4'b0100;
														assign node34219 = (inp[9]) ? node34221 : 4'b0000;
															assign node34221 = (inp[5]) ? 4'b0110 : 4'b0100;
													assign node34224 = (inp[5]) ? node34232 : node34225;
														assign node34225 = (inp[9]) ? node34229 : node34226;
															assign node34226 = (inp[4]) ? 4'b0000 : 4'b0100;
															assign node34229 = (inp[4]) ? 4'b0110 : 4'b0000;
														assign node34232 = (inp[4]) ? node34234 : 4'b0010;
															assign node34234 = (inp[9]) ? 4'b0110 : 4'b0010;
											assign node34237 = (inp[0]) ? node34253 : node34238;
												assign node34238 = (inp[4]) ? node34246 : node34239;
													assign node34239 = (inp[9]) ? 4'b0000 : node34240;
														assign node34240 = (inp[3]) ? node34242 : 4'b0100;
															assign node34242 = (inp[10]) ? 4'b0110 : 4'b0100;
													assign node34246 = (inp[9]) ? 4'b0110 : node34247;
														assign node34247 = (inp[3]) ? node34249 : 4'b0000;
															assign node34249 = (inp[5]) ? 4'b0010 : 4'b0000;
												assign node34253 = (inp[5]) ? node34263 : node34254;
													assign node34254 = (inp[4]) ? node34258 : node34255;
														assign node34255 = (inp[9]) ? 4'b0010 : 4'b0110;
														assign node34258 = (inp[9]) ? node34260 : 4'b0010;
															assign node34260 = (inp[10]) ? 4'b0110 : 4'b0100;
													assign node34263 = (inp[3]) ? 4'b0000 : node34264;
														assign node34264 = (inp[9]) ? node34268 : node34265;
															assign node34265 = (inp[4]) ? 4'b0010 : 4'b0110;
															assign node34268 = (inp[4]) ? 4'b0100 : 4'b0010;
										assign node34272 = (inp[3]) ? node34346 : node34273;
											assign node34273 = (inp[9]) ? node34311 : node34274;
												assign node34274 = (inp[4]) ? node34290 : node34275;
													assign node34275 = (inp[5]) ? node34283 : node34276;
														assign node34276 = (inp[0]) ? node34280 : node34277;
															assign node34277 = (inp[15]) ? 4'b0101 : 4'b0111;
															assign node34280 = (inp[15]) ? 4'b0111 : 4'b0101;
														assign node34283 = (inp[0]) ? node34287 : node34284;
															assign node34284 = (inp[15]) ? 4'b0101 : 4'b0111;
															assign node34287 = (inp[15]) ? 4'b0111 : 4'b0101;
													assign node34290 = (inp[10]) ? node34306 : node34291;
														assign node34291 = (inp[5]) ? node34299 : node34292;
															assign node34292 = (inp[15]) ? node34296 : node34293;
																assign node34293 = (inp[0]) ? 4'b0001 : 4'b0011;
																assign node34296 = (inp[0]) ? 4'b0011 : 4'b0001;
															assign node34299 = (inp[0]) ? node34303 : node34300;
																assign node34300 = (inp[15]) ? 4'b0001 : 4'b0011;
																assign node34303 = (inp[15]) ? 4'b0011 : 4'b0001;
														assign node34306 = (inp[0]) ? 4'b0011 : node34307;
															assign node34307 = (inp[15]) ? 4'b0001 : 4'b0011;
												assign node34311 = (inp[4]) ? node34327 : node34312;
													assign node34312 = (inp[5]) ? node34320 : node34313;
														assign node34313 = (inp[0]) ? node34317 : node34314;
															assign node34314 = (inp[15]) ? 4'b0001 : 4'b0011;
															assign node34317 = (inp[15]) ? 4'b0011 : 4'b0001;
														assign node34320 = (inp[10]) ? 4'b0001 : node34321;
															assign node34321 = (inp[0]) ? node34323 : 4'b0001;
																assign node34323 = (inp[15]) ? 4'b0011 : 4'b0001;
													assign node34327 = (inp[10]) ? node34335 : node34328;
														assign node34328 = (inp[15]) ? node34330 : 4'b0101;
															assign node34330 = (inp[0]) ? node34332 : 4'b0101;
																assign node34332 = (inp[5]) ? 4'b0101 : 4'b0111;
														assign node34335 = (inp[0]) ? node34341 : node34336;
															assign node34336 = (inp[5]) ? 4'b0111 : node34337;
																assign node34337 = (inp[15]) ? 4'b0101 : 4'b0111;
															assign node34341 = (inp[5]) ? 4'b0101 : node34342;
																assign node34342 = (inp[15]) ? 4'b0111 : 4'b0101;
											assign node34346 = (inp[10]) ? node34388 : node34347;
												assign node34347 = (inp[5]) ? node34371 : node34348;
													assign node34348 = (inp[15]) ? node34360 : node34349;
														assign node34349 = (inp[4]) ? node34355 : node34350;
															assign node34350 = (inp[9]) ? 4'b0011 : node34351;
																assign node34351 = (inp[0]) ? 4'b0101 : 4'b0111;
															assign node34355 = (inp[9]) ? node34357 : 4'b0001;
																assign node34357 = (inp[0]) ? 4'b0111 : 4'b0101;
														assign node34360 = (inp[0]) ? node34366 : node34361;
															assign node34361 = (inp[4]) ? 4'b0111 : node34362;
																assign node34362 = (inp[9]) ? 4'b0001 : 4'b0101;
															assign node34366 = (inp[9]) ? 4'b0011 : node34367;
																assign node34367 = (inp[4]) ? 4'b0011 : 4'b0111;
													assign node34371 = (inp[9]) ? node34381 : node34372;
														assign node34372 = (inp[4]) ? 4'b0011 : node34373;
															assign node34373 = (inp[15]) ? node34377 : node34374;
																assign node34374 = (inp[0]) ? 4'b0111 : 4'b0101;
																assign node34377 = (inp[0]) ? 4'b0101 : 4'b0111;
														assign node34381 = (inp[0]) ? node34385 : node34382;
															assign node34382 = (inp[15]) ? 4'b0111 : 4'b0101;
															assign node34385 = (inp[15]) ? 4'b0101 : 4'b0111;
												assign node34388 = (inp[9]) ? node34404 : node34389;
													assign node34389 = (inp[4]) ? node34397 : node34390;
														assign node34390 = (inp[5]) ? node34392 : 4'b0101;
															assign node34392 = (inp[0]) ? 4'b0101 : node34393;
																assign node34393 = (inp[15]) ? 4'b0111 : 4'b0101;
														assign node34397 = (inp[5]) ? node34399 : 4'b0001;
															assign node34399 = (inp[0]) ? node34401 : 4'b0001;
																assign node34401 = (inp[15]) ? 4'b0001 : 4'b0011;
													assign node34404 = (inp[4]) ? node34412 : node34405;
														assign node34405 = (inp[0]) ? 4'b0001 : node34406;
															assign node34406 = (inp[5]) ? 4'b0011 : node34407;
																assign node34407 = (inp[15]) ? 4'b0001 : 4'b0011;
														assign node34412 = (inp[15]) ? node34416 : node34413;
															assign node34413 = (inp[0]) ? 4'b0111 : 4'b0101;
															assign node34416 = (inp[0]) ? 4'b0101 : 4'b0111;
									assign node34419 = (inp[5]) ? node34533 : node34420;
										assign node34420 = (inp[4]) ? node34460 : node34421;
											assign node34421 = (inp[9]) ? node34453 : node34422;
												assign node34422 = (inp[3]) ? node34440 : node34423;
													assign node34423 = (inp[10]) ? node34431 : node34424;
														assign node34424 = (inp[0]) ? node34428 : node34425;
															assign node34425 = (inp[15]) ? 4'b0101 : 4'b0111;
															assign node34428 = (inp[15]) ? 4'b0111 : 4'b0101;
														assign node34431 = (inp[14]) ? node34433 : 4'b0101;
															assign node34433 = (inp[15]) ? node34437 : node34434;
																assign node34434 = (inp[0]) ? 4'b0101 : 4'b0111;
																assign node34437 = (inp[0]) ? 4'b0111 : 4'b0101;
													assign node34440 = (inp[14]) ? node34448 : node34441;
														assign node34441 = (inp[0]) ? node34445 : node34442;
															assign node34442 = (inp[15]) ? 4'b0101 : 4'b0111;
															assign node34445 = (inp[15]) ? 4'b0111 : 4'b0101;
														assign node34448 = (inp[0]) ? node34450 : 4'b0101;
															assign node34450 = (inp[15]) ? 4'b0111 : 4'b0101;
												assign node34453 = (inp[15]) ? node34457 : node34454;
													assign node34454 = (inp[0]) ? 4'b0001 : 4'b0011;
													assign node34457 = (inp[0]) ? 4'b0011 : 4'b0001;
											assign node34460 = (inp[9]) ? node34496 : node34461;
												assign node34461 = (inp[3]) ? node34489 : node34462;
													assign node34462 = (inp[10]) ? node34478 : node34463;
														assign node34463 = (inp[14]) ? node34471 : node34464;
															assign node34464 = (inp[15]) ? node34468 : node34465;
																assign node34465 = (inp[0]) ? 4'b0001 : 4'b0011;
																assign node34468 = (inp[0]) ? 4'b0011 : 4'b0001;
															assign node34471 = (inp[0]) ? node34475 : node34472;
																assign node34472 = (inp[15]) ? 4'b0001 : 4'b0011;
																assign node34475 = (inp[15]) ? 4'b0011 : 4'b0001;
														assign node34478 = (inp[14]) ? node34484 : node34479;
															assign node34479 = (inp[0]) ? 4'b0001 : node34480;
																assign node34480 = (inp[15]) ? 4'b0001 : 4'b0011;
															assign node34484 = (inp[0]) ? node34486 : 4'b0001;
																assign node34486 = (inp[15]) ? 4'b0011 : 4'b0001;
													assign node34489 = (inp[0]) ? node34493 : node34490;
														assign node34490 = (inp[15]) ? 4'b0001 : 4'b0011;
														assign node34493 = (inp[15]) ? 4'b0011 : 4'b0001;
												assign node34496 = (inp[15]) ? node34510 : node34497;
													assign node34497 = (inp[10]) ? node34503 : node34498;
														assign node34498 = (inp[0]) ? node34500 : 4'b0111;
															assign node34500 = (inp[3]) ? 4'b0111 : 4'b0101;
														assign node34503 = (inp[0]) ? node34507 : node34504;
															assign node34504 = (inp[3]) ? 4'b0101 : 4'b0111;
															assign node34507 = (inp[3]) ? 4'b0111 : 4'b0101;
													assign node34510 = (inp[10]) ? node34526 : node34511;
														assign node34511 = (inp[14]) ? node34519 : node34512;
															assign node34512 = (inp[0]) ? node34516 : node34513;
																assign node34513 = (inp[3]) ? 4'b0111 : 4'b0101;
																assign node34516 = (inp[3]) ? 4'b0101 : 4'b0111;
															assign node34519 = (inp[0]) ? node34523 : node34520;
																assign node34520 = (inp[3]) ? 4'b0111 : 4'b0101;
																assign node34523 = (inp[3]) ? 4'b0101 : 4'b0111;
														assign node34526 = (inp[3]) ? node34530 : node34527;
															assign node34527 = (inp[0]) ? 4'b0111 : 4'b0101;
															assign node34530 = (inp[0]) ? 4'b0101 : 4'b0111;
										assign node34533 = (inp[10]) ? node34637 : node34534;
											assign node34534 = (inp[14]) ? node34588 : node34535;
												assign node34535 = (inp[3]) ? node34565 : node34536;
													assign node34536 = (inp[9]) ? node34550 : node34537;
														assign node34537 = (inp[4]) ? node34543 : node34538;
															assign node34538 = (inp[15]) ? 4'b0101 : node34539;
																assign node34539 = (inp[0]) ? 4'b0101 : 4'b0111;
															assign node34543 = (inp[15]) ? node34547 : node34544;
																assign node34544 = (inp[0]) ? 4'b0001 : 4'b0011;
																assign node34547 = (inp[0]) ? 4'b0011 : 4'b0001;
														assign node34550 = (inp[4]) ? node34558 : node34551;
															assign node34551 = (inp[15]) ? node34555 : node34552;
																assign node34552 = (inp[0]) ? 4'b0001 : 4'b0011;
																assign node34555 = (inp[0]) ? 4'b0011 : 4'b0001;
															assign node34558 = (inp[15]) ? node34562 : node34559;
																assign node34559 = (inp[0]) ? 4'b0111 : 4'b0101;
																assign node34562 = (inp[0]) ? 4'b0101 : 4'b0111;
													assign node34565 = (inp[0]) ? node34579 : node34566;
														assign node34566 = (inp[15]) ? node34574 : node34567;
															assign node34567 = (inp[4]) ? node34571 : node34568;
																assign node34568 = (inp[9]) ? 4'b0001 : 4'b0101;
																assign node34571 = (inp[9]) ? 4'b0101 : 4'b0001;
															assign node34574 = (inp[4]) ? node34576 : 4'b0011;
																assign node34576 = (inp[9]) ? 4'b0111 : 4'b0011;
														assign node34579 = (inp[15]) ? 4'b0101 : node34580;
															assign node34580 = (inp[9]) ? node34584 : node34581;
																assign node34581 = (inp[4]) ? 4'b0011 : 4'b0111;
																assign node34584 = (inp[4]) ? 4'b0111 : 4'b0011;
												assign node34588 = (inp[15]) ? node34608 : node34589;
													assign node34589 = (inp[9]) ? node34601 : node34590;
														assign node34590 = (inp[4]) ? node34598 : node34591;
															assign node34591 = (inp[0]) ? node34595 : node34592;
																assign node34592 = (inp[3]) ? 4'b0101 : 4'b0111;
																assign node34595 = (inp[3]) ? 4'b0111 : 4'b0101;
															assign node34598 = (inp[3]) ? 4'b0011 : 4'b0001;
														assign node34601 = (inp[4]) ? 4'b0101 : node34602;
															assign node34602 = (inp[3]) ? 4'b0001 : node34603;
																assign node34603 = (inp[0]) ? 4'b0001 : 4'b0011;
													assign node34608 = (inp[0]) ? node34622 : node34609;
														assign node34609 = (inp[3]) ? node34617 : node34610;
															assign node34610 = (inp[9]) ? node34614 : node34611;
																assign node34611 = (inp[4]) ? 4'b0001 : 4'b0101;
																assign node34614 = (inp[4]) ? 4'b0111 : 4'b0001;
															assign node34617 = (inp[9]) ? node34619 : 4'b0011;
																assign node34619 = (inp[4]) ? 4'b0111 : 4'b0011;
														assign node34622 = (inp[3]) ? node34630 : node34623;
															assign node34623 = (inp[9]) ? node34627 : node34624;
																assign node34624 = (inp[4]) ? 4'b0011 : 4'b0111;
																assign node34627 = (inp[4]) ? 4'b0101 : 4'b0011;
															assign node34630 = (inp[4]) ? node34634 : node34631;
																assign node34631 = (inp[9]) ? 4'b0001 : 4'b0101;
																assign node34634 = (inp[9]) ? 4'b0101 : 4'b0001;
											assign node34637 = (inp[9]) ? node34681 : node34638;
												assign node34638 = (inp[4]) ? node34662 : node34639;
													assign node34639 = (inp[3]) ? node34655 : node34640;
														assign node34640 = (inp[14]) ? node34648 : node34641;
															assign node34641 = (inp[0]) ? node34645 : node34642;
																assign node34642 = (inp[15]) ? 4'b0101 : 4'b0111;
																assign node34645 = (inp[15]) ? 4'b0111 : 4'b0101;
															assign node34648 = (inp[0]) ? node34652 : node34649;
																assign node34649 = (inp[15]) ? 4'b0101 : 4'b0111;
																assign node34652 = (inp[15]) ? 4'b0111 : 4'b0101;
														assign node34655 = (inp[0]) ? node34659 : node34656;
															assign node34656 = (inp[15]) ? 4'b0111 : 4'b0101;
															assign node34659 = (inp[15]) ? 4'b0101 : 4'b0111;
													assign node34662 = (inp[0]) ? node34674 : node34663;
														assign node34663 = (inp[14]) ? node34669 : node34664;
															assign node34664 = (inp[3]) ? 4'b0001 : node34665;
																assign node34665 = (inp[15]) ? 4'b0001 : 4'b0011;
															assign node34669 = (inp[3]) ? node34671 : 4'b0001;
																assign node34671 = (inp[15]) ? 4'b0011 : 4'b0001;
														assign node34674 = (inp[3]) ? node34678 : node34675;
															assign node34675 = (inp[15]) ? 4'b0011 : 4'b0001;
															assign node34678 = (inp[15]) ? 4'b0001 : 4'b0011;
												assign node34681 = (inp[4]) ? node34701 : node34682;
													assign node34682 = (inp[0]) ? node34696 : node34683;
														assign node34683 = (inp[14]) ? node34689 : node34684;
															assign node34684 = (inp[3]) ? 4'b0011 : node34685;
																assign node34685 = (inp[15]) ? 4'b0001 : 4'b0011;
															assign node34689 = (inp[15]) ? node34693 : node34690;
																assign node34690 = (inp[3]) ? 4'b0001 : 4'b0011;
																assign node34693 = (inp[3]) ? 4'b0011 : 4'b0001;
														assign node34696 = (inp[14]) ? node34698 : 4'b0001;
															assign node34698 = (inp[15]) ? 4'b0011 : 4'b0001;
													assign node34701 = (inp[15]) ? node34705 : node34702;
														assign node34702 = (inp[0]) ? 4'b0111 : 4'b0101;
														assign node34705 = (inp[0]) ? 4'b0101 : 4'b0111;
								assign node34708 = (inp[14]) ? node34916 : node34709;
									assign node34709 = (inp[2]) ? node34809 : node34710;
										assign node34710 = (inp[9]) ? node34762 : node34711;
											assign node34711 = (inp[4]) ? node34733 : node34712;
												assign node34712 = (inp[0]) ? node34722 : node34713;
													assign node34713 = (inp[15]) ? node34717 : node34714;
														assign node34714 = (inp[3]) ? 4'b0101 : 4'b0111;
														assign node34717 = (inp[3]) ? node34719 : 4'b0101;
															assign node34719 = (inp[5]) ? 4'b0111 : 4'b0101;
													assign node34722 = (inp[15]) ? node34728 : node34723;
														assign node34723 = (inp[3]) ? node34725 : 4'b0101;
															assign node34725 = (inp[5]) ? 4'b0111 : 4'b0101;
														assign node34728 = (inp[3]) ? node34730 : 4'b0111;
															assign node34730 = (inp[5]) ? 4'b0101 : 4'b0111;
												assign node34733 = (inp[3]) ? node34747 : node34734;
													assign node34734 = (inp[5]) ? node34740 : node34735;
														assign node34735 = (inp[15]) ? node34737 : 4'b0011;
															assign node34737 = (inp[0]) ? 4'b0011 : 4'b0001;
														assign node34740 = (inp[0]) ? node34744 : node34741;
															assign node34741 = (inp[15]) ? 4'b0001 : 4'b0011;
															assign node34744 = (inp[15]) ? 4'b0011 : 4'b0001;
													assign node34747 = (inp[5]) ? node34755 : node34748;
														assign node34748 = (inp[0]) ? node34752 : node34749;
															assign node34749 = (inp[15]) ? 4'b0001 : 4'b0011;
															assign node34752 = (inp[10]) ? 4'b0001 : 4'b0011;
														assign node34755 = (inp[0]) ? node34759 : node34756;
															assign node34756 = (inp[15]) ? 4'b0011 : 4'b0001;
															assign node34759 = (inp[15]) ? 4'b0001 : 4'b0011;
											assign node34762 = (inp[4]) ? node34786 : node34763;
												assign node34763 = (inp[15]) ? node34775 : node34764;
													assign node34764 = (inp[0]) ? node34770 : node34765;
														assign node34765 = (inp[5]) ? node34767 : 4'b0011;
															assign node34767 = (inp[3]) ? 4'b0001 : 4'b0011;
														assign node34770 = (inp[3]) ? node34772 : 4'b0001;
															assign node34772 = (inp[5]) ? 4'b0011 : 4'b0001;
													assign node34775 = (inp[0]) ? node34781 : node34776;
														assign node34776 = (inp[5]) ? node34778 : 4'b0001;
															assign node34778 = (inp[3]) ? 4'b0011 : 4'b0001;
														assign node34781 = (inp[3]) ? node34783 : 4'b0011;
															assign node34783 = (inp[5]) ? 4'b0001 : 4'b0011;
												assign node34786 = (inp[0]) ? node34798 : node34787;
													assign node34787 = (inp[15]) ? node34793 : node34788;
														assign node34788 = (inp[3]) ? 4'b0101 : node34789;
															assign node34789 = (inp[5]) ? 4'b0101 : 4'b0111;
														assign node34793 = (inp[5]) ? 4'b0111 : node34794;
															assign node34794 = (inp[3]) ? 4'b0111 : 4'b0101;
													assign node34798 = (inp[15]) ? node34804 : node34799;
														assign node34799 = (inp[3]) ? 4'b0111 : node34800;
															assign node34800 = (inp[5]) ? 4'b0111 : 4'b0101;
														assign node34804 = (inp[5]) ? 4'b0101 : node34805;
															assign node34805 = (inp[3]) ? 4'b0101 : 4'b0111;
										assign node34809 = (inp[15]) ? node34863 : node34810;
											assign node34810 = (inp[0]) ? node34834 : node34811;
												assign node34811 = (inp[5]) ? node34821 : node34812;
													assign node34812 = (inp[9]) ? node34816 : node34813;
														assign node34813 = (inp[4]) ? 4'b0010 : 4'b0110;
														assign node34816 = (inp[4]) ? node34818 : 4'b0010;
															assign node34818 = (inp[3]) ? 4'b0100 : 4'b0110;
													assign node34821 = (inp[3]) ? node34829 : node34822;
														assign node34822 = (inp[4]) ? node34826 : node34823;
															assign node34823 = (inp[9]) ? 4'b0010 : 4'b0110;
															assign node34826 = (inp[9]) ? 4'b0100 : 4'b0010;
														assign node34829 = (inp[4]) ? 4'b0100 : node34830;
															assign node34830 = (inp[9]) ? 4'b0000 : 4'b0100;
												assign node34834 = (inp[5]) ? node34848 : node34835;
													assign node34835 = (inp[3]) ? node34843 : node34836;
														assign node34836 = (inp[9]) ? node34840 : node34837;
															assign node34837 = (inp[4]) ? 4'b0000 : 4'b0100;
															assign node34840 = (inp[4]) ? 4'b0100 : 4'b0000;
														assign node34843 = (inp[4]) ? node34845 : 4'b0000;
															assign node34845 = (inp[9]) ? 4'b0110 : 4'b0000;
													assign node34848 = (inp[3]) ? node34856 : node34849;
														assign node34849 = (inp[4]) ? node34853 : node34850;
															assign node34850 = (inp[9]) ? 4'b0000 : 4'b0100;
															assign node34853 = (inp[9]) ? 4'b0110 : 4'b0000;
														assign node34856 = (inp[10]) ? 4'b0110 : node34857;
															assign node34857 = (inp[9]) ? node34859 : 4'b0110;
																assign node34859 = (inp[4]) ? 4'b0110 : 4'b0010;
											assign node34863 = (inp[0]) ? node34895 : node34864;
												assign node34864 = (inp[3]) ? node34880 : node34865;
													assign node34865 = (inp[5]) ? node34873 : node34866;
														assign node34866 = (inp[10]) ? node34868 : 4'b0100;
															assign node34868 = (inp[9]) ? node34870 : 4'b0000;
																assign node34870 = (inp[4]) ? 4'b0100 : 4'b0000;
														assign node34873 = (inp[9]) ? node34877 : node34874;
															assign node34874 = (inp[4]) ? 4'b0000 : 4'b0100;
															assign node34877 = (inp[4]) ? 4'b0110 : 4'b0000;
													assign node34880 = (inp[5]) ? node34888 : node34881;
														assign node34881 = (inp[9]) ? node34885 : node34882;
															assign node34882 = (inp[4]) ? 4'b0000 : 4'b0100;
															assign node34885 = (inp[4]) ? 4'b0110 : 4'b0000;
														assign node34888 = (inp[9]) ? node34892 : node34889;
															assign node34889 = (inp[4]) ? 4'b0010 : 4'b0110;
															assign node34892 = (inp[4]) ? 4'b0110 : 4'b0010;
												assign node34895 = (inp[3]) ? node34903 : node34896;
													assign node34896 = (inp[4]) ? node34900 : node34897;
														assign node34897 = (inp[9]) ? 4'b0010 : 4'b0110;
														assign node34900 = (inp[9]) ? 4'b0110 : 4'b0010;
													assign node34903 = (inp[5]) ? node34911 : node34904;
														assign node34904 = (inp[9]) ? node34908 : node34905;
															assign node34905 = (inp[4]) ? 4'b0010 : 4'b0110;
															assign node34908 = (inp[4]) ? 4'b0100 : 4'b0010;
														assign node34911 = (inp[4]) ? 4'b0000 : node34912;
															assign node34912 = (inp[9]) ? 4'b0000 : 4'b0100;
									assign node34916 = (inp[3]) ? node34978 : node34917;
										assign node34917 = (inp[9]) ? node34955 : node34918;
											assign node34918 = (inp[4]) ? node34926 : node34919;
												assign node34919 = (inp[0]) ? node34923 : node34920;
													assign node34920 = (inp[15]) ? 4'b0100 : 4'b0110;
													assign node34923 = (inp[15]) ? 4'b0110 : 4'b0100;
												assign node34926 = (inp[5]) ? node34942 : node34927;
													assign node34927 = (inp[2]) ? node34935 : node34928;
														assign node34928 = (inp[15]) ? node34932 : node34929;
															assign node34929 = (inp[0]) ? 4'b0000 : 4'b0010;
															assign node34932 = (inp[0]) ? 4'b0010 : 4'b0000;
														assign node34935 = (inp[0]) ? node34939 : node34936;
															assign node34936 = (inp[15]) ? 4'b0000 : 4'b0010;
															assign node34939 = (inp[15]) ? 4'b0010 : 4'b0000;
													assign node34942 = (inp[10]) ? node34950 : node34943;
														assign node34943 = (inp[0]) ? node34947 : node34944;
															assign node34944 = (inp[15]) ? 4'b0000 : 4'b0010;
															assign node34947 = (inp[15]) ? 4'b0010 : 4'b0000;
														assign node34950 = (inp[0]) ? 4'b0010 : node34951;
															assign node34951 = (inp[2]) ? 4'b0010 : 4'b0000;
											assign node34955 = (inp[4]) ? node34963 : node34956;
												assign node34956 = (inp[0]) ? node34960 : node34957;
													assign node34957 = (inp[15]) ? 4'b0000 : 4'b0010;
													assign node34960 = (inp[15]) ? 4'b0010 : 4'b0000;
												assign node34963 = (inp[15]) ? node34971 : node34964;
													assign node34964 = (inp[0]) ? node34968 : node34965;
														assign node34965 = (inp[5]) ? 4'b0100 : 4'b0110;
														assign node34968 = (inp[5]) ? 4'b0110 : 4'b0100;
													assign node34971 = (inp[2]) ? node34973 : 4'b0110;
														assign node34973 = (inp[0]) ? 4'b0100 : node34974;
															assign node34974 = (inp[5]) ? 4'b0110 : 4'b0100;
										assign node34978 = (inp[0]) ? node35038 : node34979;
											assign node34979 = (inp[2]) ? node35007 : node34980;
												assign node34980 = (inp[9]) ? node34996 : node34981;
													assign node34981 = (inp[4]) ? node34987 : node34982;
														assign node34982 = (inp[15]) ? node34984 : 4'b0110;
															assign node34984 = (inp[5]) ? 4'b0110 : 4'b0100;
														assign node34987 = (inp[10]) ? 4'b0010 : node34988;
															assign node34988 = (inp[5]) ? node34992 : node34989;
																assign node34989 = (inp[15]) ? 4'b0000 : 4'b0010;
																assign node34992 = (inp[15]) ? 4'b0010 : 4'b0000;
													assign node34996 = (inp[4]) ? node35004 : node34997;
														assign node34997 = (inp[15]) ? node35001 : node34998;
															assign node34998 = (inp[5]) ? 4'b0000 : 4'b0010;
															assign node35001 = (inp[5]) ? 4'b0010 : 4'b0000;
														assign node35004 = (inp[15]) ? 4'b0110 : 4'b0100;
												assign node35007 = (inp[15]) ? node35027 : node35008;
													assign node35008 = (inp[5]) ? node35014 : node35009;
														assign node35009 = (inp[10]) ? 4'b0010 : node35010;
															assign node35010 = (inp[9]) ? 4'b0100 : 4'b0110;
														assign node35014 = (inp[10]) ? node35020 : node35015;
															assign node35015 = (inp[4]) ? node35017 : 4'b0100;
																assign node35017 = (inp[9]) ? 4'b0100 : 4'b0000;
															assign node35020 = (inp[4]) ? node35024 : node35021;
																assign node35021 = (inp[9]) ? 4'b0000 : 4'b0100;
																assign node35024 = (inp[9]) ? 4'b0100 : 4'b0000;
													assign node35027 = (inp[5]) ? node35033 : node35028;
														assign node35028 = (inp[4]) ? 4'b0000 : node35029;
															assign node35029 = (inp[9]) ? 4'b0000 : 4'b0100;
														assign node35033 = (inp[4]) ? node35035 : 4'b0010;
															assign node35035 = (inp[9]) ? 4'b0110 : 4'b0010;
											assign node35038 = (inp[15]) ? node35054 : node35039;
												assign node35039 = (inp[5]) ? node35047 : node35040;
													assign node35040 = (inp[4]) ? node35044 : node35041;
														assign node35041 = (inp[9]) ? 4'b0000 : 4'b0100;
														assign node35044 = (inp[9]) ? 4'b0110 : 4'b0000;
													assign node35047 = (inp[4]) ? node35051 : node35048;
														assign node35048 = (inp[9]) ? 4'b0010 : 4'b0110;
														assign node35051 = (inp[9]) ? 4'b0110 : 4'b0010;
												assign node35054 = (inp[5]) ? node35062 : node35055;
													assign node35055 = (inp[4]) ? node35059 : node35056;
														assign node35056 = (inp[9]) ? 4'b0010 : 4'b0110;
														assign node35059 = (inp[9]) ? 4'b0100 : 4'b0010;
													assign node35062 = (inp[2]) ? node35076 : node35063;
														assign node35063 = (inp[10]) ? node35071 : node35064;
															assign node35064 = (inp[9]) ? node35068 : node35065;
																assign node35065 = (inp[4]) ? 4'b0000 : 4'b0100;
																assign node35068 = (inp[4]) ? 4'b0100 : 4'b0000;
															assign node35071 = (inp[9]) ? node35073 : 4'b0100;
																assign node35073 = (inp[4]) ? 4'b0100 : 4'b0000;
														assign node35076 = (inp[4]) ? node35078 : 4'b0100;
															assign node35078 = (inp[9]) ? 4'b0100 : 4'b0000;
						assign node35081 = (inp[10]) ? node36197 : node35082;
							assign node35082 = (inp[15]) ? node35632 : node35083;
								assign node35083 = (inp[0]) ? node35349 : node35084;
									assign node35084 = (inp[5]) ? node35200 : node35085;
										assign node35085 = (inp[4]) ? node35143 : node35086;
											assign node35086 = (inp[9]) ? node35120 : node35087;
												assign node35087 = (inp[2]) ? node35113 : node35088;
													assign node35088 = (inp[3]) ? node35098 : node35089;
														assign node35089 = (inp[7]) ? node35091 : 4'b0111;
															assign node35091 = (inp[14]) ? node35095 : node35092;
																assign node35092 = (inp[8]) ? 4'b0111 : 4'b0110;
																assign node35095 = (inp[8]) ? 4'b0110 : 4'b0111;
														assign node35098 = (inp[7]) ? node35106 : node35099;
															assign node35099 = (inp[14]) ? node35103 : node35100;
																assign node35100 = (inp[8]) ? 4'b0110 : 4'b0111;
																assign node35103 = (inp[8]) ? 4'b0111 : 4'b0110;
															assign node35106 = (inp[14]) ? node35110 : node35107;
																assign node35107 = (inp[8]) ? 4'b0111 : 4'b0110;
																assign node35110 = (inp[8]) ? 4'b0110 : 4'b0111;
													assign node35113 = (inp[7]) ? node35117 : node35114;
														assign node35114 = (inp[8]) ? 4'b0111 : 4'b0110;
														assign node35117 = (inp[8]) ? 4'b0110 : 4'b0111;
												assign node35120 = (inp[7]) ? node35132 : node35121;
													assign node35121 = (inp[8]) ? node35127 : node35122;
														assign node35122 = (inp[14]) ? 4'b0010 : node35123;
															assign node35123 = (inp[2]) ? 4'b0010 : 4'b0011;
														assign node35127 = (inp[14]) ? 4'b0011 : node35128;
															assign node35128 = (inp[2]) ? 4'b0011 : 4'b0010;
													assign node35132 = (inp[8]) ? node35138 : node35133;
														assign node35133 = (inp[14]) ? 4'b0011 : node35134;
															assign node35134 = (inp[2]) ? 4'b0011 : 4'b0010;
														assign node35138 = (inp[14]) ? 4'b0010 : node35139;
															assign node35139 = (inp[2]) ? 4'b0010 : 4'b0011;
											assign node35143 = (inp[9]) ? node35161 : node35144;
												assign node35144 = (inp[8]) ? node35150 : node35145;
													assign node35145 = (inp[7]) ? 4'b0011 : node35146;
														assign node35146 = (inp[2]) ? 4'b0010 : 4'b0011;
													assign node35150 = (inp[7]) ? node35156 : node35151;
														assign node35151 = (inp[14]) ? 4'b0011 : node35152;
															assign node35152 = (inp[2]) ? 4'b0011 : 4'b0010;
														assign node35156 = (inp[14]) ? 4'b0010 : node35157;
															assign node35157 = (inp[2]) ? 4'b0010 : 4'b0011;
												assign node35161 = (inp[3]) ? node35179 : node35162;
													assign node35162 = (inp[8]) ? node35168 : node35163;
														assign node35163 = (inp[7]) ? node35165 : 4'b0110;
															assign node35165 = (inp[14]) ? 4'b0111 : 4'b0110;
														assign node35168 = (inp[7]) ? node35174 : node35169;
															assign node35169 = (inp[2]) ? 4'b0111 : node35170;
																assign node35170 = (inp[14]) ? 4'b0111 : 4'b0110;
															assign node35174 = (inp[14]) ? 4'b0110 : node35175;
																assign node35175 = (inp[2]) ? 4'b0110 : 4'b0111;
													assign node35179 = (inp[2]) ? node35193 : node35180;
														assign node35180 = (inp[8]) ? node35188 : node35181;
															assign node35181 = (inp[7]) ? node35185 : node35182;
																assign node35182 = (inp[14]) ? 4'b0100 : 4'b0101;
																assign node35185 = (inp[14]) ? 4'b0101 : 4'b0100;
															assign node35188 = (inp[7]) ? node35190 : 4'b0101;
																assign node35190 = (inp[14]) ? 4'b0100 : 4'b0101;
														assign node35193 = (inp[7]) ? node35197 : node35194;
															assign node35194 = (inp[8]) ? 4'b0101 : 4'b0100;
															assign node35197 = (inp[8]) ? 4'b0100 : 4'b0101;
										assign node35200 = (inp[3]) ? node35282 : node35201;
											assign node35201 = (inp[4]) ? node35237 : node35202;
												assign node35202 = (inp[9]) ? node35220 : node35203;
													assign node35203 = (inp[2]) ? node35217 : node35204;
														assign node35204 = (inp[7]) ? node35212 : node35205;
															assign node35205 = (inp[8]) ? node35209 : node35206;
																assign node35206 = (inp[14]) ? 4'b0110 : 4'b0111;
																assign node35209 = (inp[14]) ? 4'b0111 : 4'b0110;
															assign node35212 = (inp[14]) ? 4'b0110 : node35213;
																assign node35213 = (inp[8]) ? 4'b0111 : 4'b0110;
														assign node35217 = (inp[8]) ? 4'b0110 : 4'b0111;
													assign node35220 = (inp[8]) ? node35226 : node35221;
														assign node35221 = (inp[7]) ? node35223 : 4'b0010;
															assign node35223 = (inp[14]) ? 4'b0011 : 4'b0010;
														assign node35226 = (inp[7]) ? node35232 : node35227;
															assign node35227 = (inp[14]) ? 4'b0011 : node35228;
																assign node35228 = (inp[2]) ? 4'b0011 : 4'b0010;
															assign node35232 = (inp[14]) ? 4'b0010 : node35233;
																assign node35233 = (inp[2]) ? 4'b0010 : 4'b0011;
												assign node35237 = (inp[9]) ? node35259 : node35238;
													assign node35238 = (inp[14]) ? node35252 : node35239;
														assign node35239 = (inp[2]) ? node35247 : node35240;
															assign node35240 = (inp[8]) ? node35244 : node35241;
																assign node35241 = (inp[7]) ? 4'b0010 : 4'b0011;
																assign node35244 = (inp[7]) ? 4'b0011 : 4'b0010;
															assign node35247 = (inp[7]) ? node35249 : 4'b0011;
																assign node35249 = (inp[8]) ? 4'b0010 : 4'b0011;
														assign node35252 = (inp[7]) ? node35256 : node35253;
															assign node35253 = (inp[8]) ? 4'b0011 : 4'b0010;
															assign node35256 = (inp[8]) ? 4'b0010 : 4'b0011;
													assign node35259 = (inp[2]) ? node35271 : node35260;
														assign node35260 = (inp[7]) ? node35266 : node35261;
															assign node35261 = (inp[8]) ? 4'b0101 : node35262;
																assign node35262 = (inp[14]) ? 4'b0100 : 4'b0101;
															assign node35266 = (inp[8]) ? 4'b0100 : node35267;
																assign node35267 = (inp[14]) ? 4'b0101 : 4'b0100;
														assign node35271 = (inp[14]) ? node35277 : node35272;
															assign node35272 = (inp[7]) ? 4'b0100 : node35273;
																assign node35273 = (inp[8]) ? 4'b0101 : 4'b0100;
															assign node35277 = (inp[7]) ? node35279 : 4'b0100;
																assign node35279 = (inp[8]) ? 4'b0100 : 4'b0101;
											assign node35282 = (inp[4]) ? node35320 : node35283;
												assign node35283 = (inp[9]) ? node35299 : node35284;
													assign node35284 = (inp[8]) ? node35290 : node35285;
														assign node35285 = (inp[7]) ? node35287 : 4'b0100;
															assign node35287 = (inp[14]) ? 4'b0101 : 4'b0100;
														assign node35290 = (inp[14]) ? node35296 : node35291;
															assign node35291 = (inp[2]) ? 4'b0101 : node35292;
																assign node35292 = (inp[7]) ? 4'b0101 : 4'b0100;
															assign node35296 = (inp[7]) ? 4'b0100 : 4'b0101;
													assign node35299 = (inp[14]) ? node35307 : node35300;
														assign node35300 = (inp[2]) ? node35302 : 4'b0000;
															assign node35302 = (inp[8]) ? 4'b0000 : node35303;
																assign node35303 = (inp[7]) ? 4'b0001 : 4'b0000;
														assign node35307 = (inp[2]) ? node35315 : node35308;
															assign node35308 = (inp[7]) ? node35312 : node35309;
																assign node35309 = (inp[8]) ? 4'b0001 : 4'b0000;
																assign node35312 = (inp[8]) ? 4'b0000 : 4'b0001;
															assign node35315 = (inp[8]) ? 4'b0000 : node35316;
																assign node35316 = (inp[7]) ? 4'b0001 : 4'b0000;
												assign node35320 = (inp[9]) ? node35338 : node35321;
													assign node35321 = (inp[2]) ? node35331 : node35322;
														assign node35322 = (inp[8]) ? 4'b0000 : node35323;
															assign node35323 = (inp[7]) ? node35327 : node35324;
																assign node35324 = (inp[14]) ? 4'b0000 : 4'b0001;
																assign node35327 = (inp[14]) ? 4'b0001 : 4'b0000;
														assign node35331 = (inp[8]) ? node35335 : node35332;
															assign node35332 = (inp[7]) ? 4'b0001 : 4'b0000;
															assign node35335 = (inp[7]) ? 4'b0000 : 4'b0001;
													assign node35338 = (inp[7]) ? node35344 : node35339;
														assign node35339 = (inp[14]) ? node35341 : 4'b0100;
															assign node35341 = (inp[8]) ? 4'b0101 : 4'b0100;
														assign node35344 = (inp[8]) ? node35346 : 4'b0101;
															assign node35346 = (inp[2]) ? 4'b0100 : 4'b0101;
									assign node35349 = (inp[3]) ? node35505 : node35350;
										assign node35350 = (inp[5]) ? node35436 : node35351;
											assign node35351 = (inp[7]) ? node35393 : node35352;
												assign node35352 = (inp[8]) ? node35378 : node35353;
													assign node35353 = (inp[14]) ? node35363 : node35354;
														assign node35354 = (inp[2]) ? node35358 : node35355;
															assign node35355 = (inp[9]) ? 4'b0001 : 4'b0101;
															assign node35358 = (inp[9]) ? 4'b0100 : node35359;
																assign node35359 = (inp[4]) ? 4'b0000 : 4'b0100;
														assign node35363 = (inp[2]) ? node35371 : node35364;
															assign node35364 = (inp[4]) ? node35368 : node35365;
																assign node35365 = (inp[9]) ? 4'b0000 : 4'b0100;
																assign node35368 = (inp[9]) ? 4'b0100 : 4'b0000;
															assign node35371 = (inp[4]) ? node35375 : node35372;
																assign node35372 = (inp[9]) ? 4'b0000 : 4'b0100;
																assign node35375 = (inp[9]) ? 4'b0100 : 4'b0000;
													assign node35378 = (inp[14]) ? node35386 : node35379;
														assign node35379 = (inp[2]) ? 4'b0001 : node35380;
															assign node35380 = (inp[9]) ? 4'b0100 : node35381;
																assign node35381 = (inp[4]) ? 4'b0000 : 4'b0100;
														assign node35386 = (inp[9]) ? node35390 : node35387;
															assign node35387 = (inp[4]) ? 4'b0001 : 4'b0101;
															assign node35390 = (inp[4]) ? 4'b0101 : 4'b0001;
												assign node35393 = (inp[8]) ? node35413 : node35394;
													assign node35394 = (inp[2]) ? node35404 : node35395;
														assign node35395 = (inp[14]) ? node35399 : node35396;
															assign node35396 = (inp[4]) ? 4'b0100 : 4'b0000;
															assign node35399 = (inp[9]) ? 4'b0101 : node35400;
																assign node35400 = (inp[4]) ? 4'b0001 : 4'b0101;
														assign node35404 = (inp[14]) ? 4'b0001 : node35405;
															assign node35405 = (inp[9]) ? node35409 : node35406;
																assign node35406 = (inp[4]) ? 4'b0001 : 4'b0101;
																assign node35409 = (inp[4]) ? 4'b0101 : 4'b0001;
													assign node35413 = (inp[14]) ? node35423 : node35414;
														assign node35414 = (inp[2]) ? node35420 : node35415;
															assign node35415 = (inp[4]) ? node35417 : 4'b0001;
																assign node35417 = (inp[9]) ? 4'b0101 : 4'b0001;
															assign node35420 = (inp[9]) ? 4'b0100 : 4'b0000;
														assign node35423 = (inp[2]) ? node35429 : node35424;
															assign node35424 = (inp[9]) ? 4'b0000 : node35425;
																assign node35425 = (inp[4]) ? 4'b0000 : 4'b0100;
															assign node35429 = (inp[9]) ? node35433 : node35430;
																assign node35430 = (inp[4]) ? 4'b0000 : 4'b0100;
																assign node35433 = (inp[4]) ? 4'b0100 : 4'b0000;
											assign node35436 = (inp[9]) ? node35474 : node35437;
												assign node35437 = (inp[4]) ? node35455 : node35438;
													assign node35438 = (inp[14]) ? node35448 : node35439;
														assign node35439 = (inp[8]) ? node35441 : 4'b0101;
															assign node35441 = (inp[2]) ? node35445 : node35442;
																assign node35442 = (inp[7]) ? 4'b0101 : 4'b0100;
																assign node35445 = (inp[7]) ? 4'b0100 : 4'b0101;
														assign node35448 = (inp[8]) ? node35452 : node35449;
															assign node35449 = (inp[7]) ? 4'b0101 : 4'b0100;
															assign node35452 = (inp[7]) ? 4'b0100 : 4'b0101;
													assign node35455 = (inp[14]) ? node35469 : node35456;
														assign node35456 = (inp[8]) ? node35462 : node35457;
															assign node35457 = (inp[2]) ? 4'b0001 : node35458;
																assign node35458 = (inp[7]) ? 4'b0000 : 4'b0001;
															assign node35462 = (inp[7]) ? node35466 : node35463;
																assign node35463 = (inp[2]) ? 4'b0001 : 4'b0000;
																assign node35466 = (inp[2]) ? 4'b0000 : 4'b0001;
														assign node35469 = (inp[7]) ? node35471 : 4'b0000;
															assign node35471 = (inp[8]) ? 4'b0000 : 4'b0001;
												assign node35474 = (inp[4]) ? node35490 : node35475;
													assign node35475 = (inp[2]) ? node35485 : node35476;
														assign node35476 = (inp[14]) ? node35478 : 4'b0000;
															assign node35478 = (inp[8]) ? node35482 : node35479;
																assign node35479 = (inp[7]) ? 4'b0001 : 4'b0000;
																assign node35482 = (inp[7]) ? 4'b0000 : 4'b0001;
														assign node35485 = (inp[7]) ? node35487 : 4'b0001;
															assign node35487 = (inp[14]) ? 4'b0000 : 4'b0001;
													assign node35490 = (inp[2]) ? node35500 : node35491;
														assign node35491 = (inp[14]) ? 4'b0111 : node35492;
															assign node35492 = (inp[7]) ? node35496 : node35493;
																assign node35493 = (inp[8]) ? 4'b0110 : 4'b0111;
																assign node35496 = (inp[8]) ? 4'b0111 : 4'b0110;
														assign node35500 = (inp[7]) ? node35502 : 4'b0110;
															assign node35502 = (inp[8]) ? 4'b0110 : 4'b0111;
										assign node35505 = (inp[5]) ? node35567 : node35506;
											assign node35506 = (inp[4]) ? node35530 : node35507;
												assign node35507 = (inp[9]) ? node35517 : node35508;
													assign node35508 = (inp[7]) ? node35510 : 4'b0100;
														assign node35510 = (inp[8]) ? node35512 : 4'b0101;
															assign node35512 = (inp[14]) ? 4'b0100 : node35513;
																assign node35513 = (inp[2]) ? 4'b0100 : 4'b0101;
													assign node35517 = (inp[8]) ? node35523 : node35518;
														assign node35518 = (inp[7]) ? node35520 : 4'b0000;
															assign node35520 = (inp[2]) ? 4'b0001 : 4'b0000;
														assign node35523 = (inp[7]) ? node35527 : node35524;
															assign node35524 = (inp[14]) ? 4'b0001 : 4'b0000;
															assign node35527 = (inp[2]) ? 4'b0000 : 4'b0001;
												assign node35530 = (inp[9]) ? node35548 : node35531;
													assign node35531 = (inp[14]) ? node35537 : node35532;
														assign node35532 = (inp[7]) ? 4'b0000 : node35533;
															assign node35533 = (inp[8]) ? 4'b0001 : 4'b0000;
														assign node35537 = (inp[2]) ? node35543 : node35538;
															assign node35538 = (inp[7]) ? node35540 : 4'b0000;
																assign node35540 = (inp[8]) ? 4'b0000 : 4'b0001;
															assign node35543 = (inp[7]) ? node35545 : 4'b0001;
																assign node35545 = (inp[8]) ? 4'b0000 : 4'b0001;
													assign node35548 = (inp[7]) ? node35560 : node35549;
														assign node35549 = (inp[8]) ? node35555 : node35550;
															assign node35550 = (inp[2]) ? 4'b0110 : node35551;
																assign node35551 = (inp[14]) ? 4'b0110 : 4'b0111;
															assign node35555 = (inp[14]) ? 4'b0111 : node35556;
																assign node35556 = (inp[2]) ? 4'b0111 : 4'b0110;
														assign node35560 = (inp[8]) ? node35562 : 4'b0111;
															assign node35562 = (inp[14]) ? 4'b0110 : node35563;
																assign node35563 = (inp[2]) ? 4'b0110 : 4'b0111;
											assign node35567 = (inp[9]) ? node35599 : node35568;
												assign node35568 = (inp[4]) ? node35582 : node35569;
													assign node35569 = (inp[7]) ? node35575 : node35570;
														assign node35570 = (inp[8]) ? 4'b0111 : node35571;
															assign node35571 = (inp[2]) ? 4'b0110 : 4'b0111;
														assign node35575 = (inp[8]) ? node35577 : 4'b0111;
															assign node35577 = (inp[14]) ? 4'b0110 : node35578;
																assign node35578 = (inp[2]) ? 4'b0110 : 4'b0111;
													assign node35582 = (inp[2]) ? node35592 : node35583;
														assign node35583 = (inp[7]) ? 4'b0011 : node35584;
															assign node35584 = (inp[14]) ? node35588 : node35585;
																assign node35585 = (inp[8]) ? 4'b0010 : 4'b0011;
																assign node35588 = (inp[8]) ? 4'b0011 : 4'b0010;
														assign node35592 = (inp[8]) ? node35596 : node35593;
															assign node35593 = (inp[7]) ? 4'b0011 : 4'b0010;
															assign node35596 = (inp[7]) ? 4'b0010 : 4'b0011;
												assign node35599 = (inp[4]) ? node35613 : node35600;
													assign node35600 = (inp[14]) ? node35606 : node35601;
														assign node35601 = (inp[2]) ? node35603 : 4'b0010;
															assign node35603 = (inp[8]) ? 4'b0010 : 4'b0011;
														assign node35606 = (inp[8]) ? node35610 : node35607;
															assign node35607 = (inp[7]) ? 4'b0011 : 4'b0010;
															assign node35610 = (inp[7]) ? 4'b0010 : 4'b0011;
													assign node35613 = (inp[2]) ? node35627 : node35614;
														assign node35614 = (inp[8]) ? node35622 : node35615;
															assign node35615 = (inp[7]) ? node35619 : node35616;
																assign node35616 = (inp[14]) ? 4'b0110 : 4'b0111;
																assign node35619 = (inp[14]) ? 4'b0111 : 4'b0110;
															assign node35622 = (inp[7]) ? 4'b0111 : node35623;
																assign node35623 = (inp[14]) ? 4'b0111 : 4'b0110;
														assign node35627 = (inp[8]) ? 4'b0110 : node35628;
															assign node35628 = (inp[7]) ? 4'b0111 : 4'b0110;
								assign node35632 = (inp[0]) ? node35918 : node35633;
									assign node35633 = (inp[5]) ? node35763 : node35634;
										assign node35634 = (inp[4]) ? node35680 : node35635;
											assign node35635 = (inp[9]) ? node35659 : node35636;
												assign node35636 = (inp[8]) ? node35648 : node35637;
													assign node35637 = (inp[7]) ? node35643 : node35638;
														assign node35638 = (inp[14]) ? 4'b0100 : node35639;
															assign node35639 = (inp[2]) ? 4'b0100 : 4'b0101;
														assign node35643 = (inp[2]) ? 4'b0101 : node35644;
															assign node35644 = (inp[14]) ? 4'b0101 : 4'b0100;
													assign node35648 = (inp[7]) ? node35654 : node35649;
														assign node35649 = (inp[2]) ? 4'b0101 : node35650;
															assign node35650 = (inp[3]) ? 4'b0100 : 4'b0101;
														assign node35654 = (inp[2]) ? 4'b0100 : node35655;
															assign node35655 = (inp[14]) ? 4'b0100 : 4'b0101;
												assign node35659 = (inp[8]) ? node35669 : node35660;
													assign node35660 = (inp[7]) ? node35666 : node35661;
														assign node35661 = (inp[14]) ? 4'b0000 : node35662;
															assign node35662 = (inp[2]) ? 4'b0000 : 4'b0001;
														assign node35666 = (inp[2]) ? 4'b0001 : 4'b0000;
													assign node35669 = (inp[7]) ? node35675 : node35670;
														assign node35670 = (inp[2]) ? 4'b0001 : node35671;
															assign node35671 = (inp[14]) ? 4'b0001 : 4'b0000;
														assign node35675 = (inp[2]) ? 4'b0000 : node35676;
															assign node35676 = (inp[14]) ? 4'b0000 : 4'b0001;
											assign node35680 = (inp[9]) ? node35718 : node35681;
												assign node35681 = (inp[2]) ? node35705 : node35682;
													assign node35682 = (inp[8]) ? node35690 : node35683;
														assign node35683 = (inp[14]) ? node35687 : node35684;
															assign node35684 = (inp[7]) ? 4'b0000 : 4'b0001;
															assign node35687 = (inp[7]) ? 4'b0001 : 4'b0000;
														assign node35690 = (inp[3]) ? node35698 : node35691;
															assign node35691 = (inp[7]) ? node35695 : node35692;
																assign node35692 = (inp[14]) ? 4'b0001 : 4'b0000;
																assign node35695 = (inp[14]) ? 4'b0000 : 4'b0001;
															assign node35698 = (inp[7]) ? node35702 : node35699;
																assign node35699 = (inp[14]) ? 4'b0001 : 4'b0000;
																assign node35702 = (inp[14]) ? 4'b0000 : 4'b0001;
													assign node35705 = (inp[14]) ? node35711 : node35706;
														assign node35706 = (inp[8]) ? node35708 : 4'b0000;
															assign node35708 = (inp[7]) ? 4'b0000 : 4'b0001;
														assign node35711 = (inp[7]) ? node35715 : node35712;
															assign node35712 = (inp[8]) ? 4'b0001 : 4'b0000;
															assign node35715 = (inp[8]) ? 4'b0000 : 4'b0001;
												assign node35718 = (inp[3]) ? node35738 : node35719;
													assign node35719 = (inp[14]) ? node35727 : node35720;
														assign node35720 = (inp[7]) ? 4'b0101 : node35721;
															assign node35721 = (inp[8]) ? node35723 : 4'b0101;
																assign node35723 = (inp[2]) ? 4'b0101 : 4'b0100;
														assign node35727 = (inp[2]) ? node35733 : node35728;
															assign node35728 = (inp[7]) ? 4'b0101 : node35729;
																assign node35729 = (inp[8]) ? 4'b0101 : 4'b0100;
															assign node35733 = (inp[8]) ? node35735 : 4'b0100;
																assign node35735 = (inp[7]) ? 4'b0100 : 4'b0101;
													assign node35738 = (inp[2]) ? node35754 : node35739;
														assign node35739 = (inp[7]) ? node35747 : node35740;
															assign node35740 = (inp[14]) ? node35744 : node35741;
																assign node35741 = (inp[8]) ? 4'b0110 : 4'b0111;
																assign node35744 = (inp[8]) ? 4'b0111 : 4'b0110;
															assign node35747 = (inp[14]) ? node35751 : node35748;
																assign node35748 = (inp[8]) ? 4'b0111 : 4'b0110;
																assign node35751 = (inp[8]) ? 4'b0110 : 4'b0111;
														assign node35754 = (inp[14]) ? node35760 : node35755;
															assign node35755 = (inp[8]) ? 4'b0110 : node35756;
																assign node35756 = (inp[7]) ? 4'b0111 : 4'b0110;
															assign node35760 = (inp[8]) ? 4'b0111 : 4'b0110;
										assign node35763 = (inp[3]) ? node35843 : node35764;
											assign node35764 = (inp[9]) ? node35810 : node35765;
												assign node35765 = (inp[4]) ? node35787 : node35766;
													assign node35766 = (inp[2]) ? node35774 : node35767;
														assign node35767 = (inp[14]) ? 4'b0101 : node35768;
															assign node35768 = (inp[8]) ? 4'b0101 : node35769;
																assign node35769 = (inp[7]) ? 4'b0100 : 4'b0101;
														assign node35774 = (inp[14]) ? node35782 : node35775;
															assign node35775 = (inp[7]) ? node35779 : node35776;
																assign node35776 = (inp[8]) ? 4'b0101 : 4'b0100;
																assign node35779 = (inp[8]) ? 4'b0100 : 4'b0101;
															assign node35782 = (inp[7]) ? node35784 : 4'b0100;
																assign node35784 = (inp[8]) ? 4'b0100 : 4'b0101;
													assign node35787 = (inp[8]) ? node35799 : node35788;
														assign node35788 = (inp[7]) ? node35794 : node35789;
															assign node35789 = (inp[2]) ? 4'b0000 : node35790;
																assign node35790 = (inp[14]) ? 4'b0000 : 4'b0001;
															assign node35794 = (inp[2]) ? 4'b0001 : node35795;
																assign node35795 = (inp[14]) ? 4'b0001 : 4'b0000;
														assign node35799 = (inp[7]) ? node35805 : node35800;
															assign node35800 = (inp[2]) ? 4'b0001 : node35801;
																assign node35801 = (inp[14]) ? 4'b0001 : 4'b0000;
															assign node35805 = (inp[2]) ? 4'b0000 : node35806;
																assign node35806 = (inp[14]) ? 4'b0000 : 4'b0001;
												assign node35810 = (inp[4]) ? node35828 : node35811;
													assign node35811 = (inp[14]) ? node35821 : node35812;
														assign node35812 = (inp[2]) ? node35814 : 4'b0000;
															assign node35814 = (inp[7]) ? node35818 : node35815;
																assign node35815 = (inp[8]) ? 4'b0001 : 4'b0000;
																assign node35818 = (inp[8]) ? 4'b0000 : 4'b0001;
														assign node35821 = (inp[7]) ? node35825 : node35822;
															assign node35822 = (inp[8]) ? 4'b0001 : 4'b0000;
															assign node35825 = (inp[8]) ? 4'b0000 : 4'b0001;
													assign node35828 = (inp[8]) ? node35836 : node35829;
														assign node35829 = (inp[7]) ? 4'b0111 : node35830;
															assign node35830 = (inp[14]) ? 4'b0110 : node35831;
																assign node35831 = (inp[2]) ? 4'b0110 : 4'b0111;
														assign node35836 = (inp[7]) ? 4'b0110 : node35837;
															assign node35837 = (inp[2]) ? 4'b0111 : node35838;
																assign node35838 = (inp[14]) ? 4'b0111 : 4'b0110;
											assign node35843 = (inp[4]) ? node35879 : node35844;
												assign node35844 = (inp[9]) ? node35862 : node35845;
													assign node35845 = (inp[2]) ? node35855 : node35846;
														assign node35846 = (inp[7]) ? 4'b0110 : node35847;
															assign node35847 = (inp[14]) ? node35851 : node35848;
																assign node35848 = (inp[8]) ? 4'b0110 : 4'b0111;
																assign node35851 = (inp[8]) ? 4'b0111 : 4'b0110;
														assign node35855 = (inp[7]) ? node35859 : node35856;
															assign node35856 = (inp[8]) ? 4'b0111 : 4'b0110;
															assign node35859 = (inp[8]) ? 4'b0110 : 4'b0111;
													assign node35862 = (inp[7]) ? node35874 : node35863;
														assign node35863 = (inp[8]) ? node35869 : node35864;
															assign node35864 = (inp[2]) ? 4'b0010 : node35865;
																assign node35865 = (inp[14]) ? 4'b0010 : 4'b0011;
															assign node35869 = (inp[2]) ? 4'b0011 : node35870;
																assign node35870 = (inp[14]) ? 4'b0011 : 4'b0010;
														assign node35874 = (inp[8]) ? node35876 : 4'b0011;
															assign node35876 = (inp[14]) ? 4'b0010 : 4'b0011;
												assign node35879 = (inp[9]) ? node35905 : node35880;
													assign node35880 = (inp[2]) ? node35896 : node35881;
														assign node35881 = (inp[14]) ? node35889 : node35882;
															assign node35882 = (inp[7]) ? node35886 : node35883;
																assign node35883 = (inp[8]) ? 4'b0010 : 4'b0011;
																assign node35886 = (inp[8]) ? 4'b0011 : 4'b0010;
															assign node35889 = (inp[7]) ? node35893 : node35890;
																assign node35890 = (inp[8]) ? 4'b0011 : 4'b0010;
																assign node35893 = (inp[8]) ? 4'b0010 : 4'b0011;
														assign node35896 = (inp[14]) ? 4'b0010 : node35897;
															assign node35897 = (inp[7]) ? node35901 : node35898;
																assign node35898 = (inp[8]) ? 4'b0011 : 4'b0010;
																assign node35901 = (inp[8]) ? 4'b0010 : 4'b0011;
													assign node35905 = (inp[8]) ? node35911 : node35906;
														assign node35906 = (inp[7]) ? node35908 : 4'b0110;
															assign node35908 = (inp[2]) ? 4'b0111 : 4'b0110;
														assign node35911 = (inp[7]) ? node35915 : node35912;
															assign node35912 = (inp[14]) ? 4'b0111 : 4'b0110;
															assign node35915 = (inp[14]) ? 4'b0110 : 4'b0111;
									assign node35918 = (inp[5]) ? node36020 : node35919;
										assign node35919 = (inp[9]) ? node35959 : node35920;
											assign node35920 = (inp[4]) ? node35944 : node35921;
												assign node35921 = (inp[8]) ? node35933 : node35922;
													assign node35922 = (inp[7]) ? node35928 : node35923;
														assign node35923 = (inp[14]) ? 4'b0110 : node35924;
															assign node35924 = (inp[2]) ? 4'b0110 : 4'b0111;
														assign node35928 = (inp[2]) ? 4'b0111 : node35929;
															assign node35929 = (inp[14]) ? 4'b0111 : 4'b0110;
													assign node35933 = (inp[7]) ? node35939 : node35934;
														assign node35934 = (inp[14]) ? 4'b0111 : node35935;
															assign node35935 = (inp[2]) ? 4'b0111 : 4'b0110;
														assign node35939 = (inp[14]) ? 4'b0110 : node35940;
															assign node35940 = (inp[2]) ? 4'b0110 : 4'b0111;
												assign node35944 = (inp[7]) ? node35954 : node35945;
													assign node35945 = (inp[8]) ? node35951 : node35946;
														assign node35946 = (inp[14]) ? 4'b0010 : node35947;
															assign node35947 = (inp[2]) ? 4'b0010 : 4'b0011;
														assign node35951 = (inp[14]) ? 4'b0011 : 4'b0010;
													assign node35954 = (inp[8]) ? node35956 : 4'b0011;
														assign node35956 = (inp[14]) ? 4'b0010 : 4'b0011;
											assign node35959 = (inp[4]) ? node35983 : node35960;
												assign node35960 = (inp[2]) ? node35976 : node35961;
													assign node35961 = (inp[8]) ? node35969 : node35962;
														assign node35962 = (inp[7]) ? node35966 : node35963;
															assign node35963 = (inp[14]) ? 4'b0010 : 4'b0011;
															assign node35966 = (inp[14]) ? 4'b0011 : 4'b0010;
														assign node35969 = (inp[7]) ? node35973 : node35970;
															assign node35970 = (inp[14]) ? 4'b0011 : 4'b0010;
															assign node35973 = (inp[14]) ? 4'b0010 : 4'b0011;
													assign node35976 = (inp[7]) ? node35980 : node35977;
														assign node35977 = (inp[8]) ? 4'b0011 : 4'b0010;
														assign node35980 = (inp[8]) ? 4'b0010 : 4'b0011;
												assign node35983 = (inp[3]) ? node35997 : node35984;
													assign node35984 = (inp[8]) ? node35990 : node35985;
														assign node35985 = (inp[7]) ? 4'b0111 : node35986;
															assign node35986 = (inp[2]) ? 4'b0110 : 4'b0111;
														assign node35990 = (inp[7]) ? 4'b0110 : node35991;
															assign node35991 = (inp[14]) ? 4'b0111 : node35992;
																assign node35992 = (inp[2]) ? 4'b0111 : 4'b0110;
													assign node35997 = (inp[2]) ? node36013 : node35998;
														assign node35998 = (inp[7]) ? node36006 : node35999;
															assign node35999 = (inp[8]) ? node36003 : node36000;
																assign node36000 = (inp[14]) ? 4'b0100 : 4'b0101;
																assign node36003 = (inp[14]) ? 4'b0101 : 4'b0100;
															assign node36006 = (inp[8]) ? node36010 : node36007;
																assign node36007 = (inp[14]) ? 4'b0101 : 4'b0100;
																assign node36010 = (inp[14]) ? 4'b0100 : 4'b0101;
														assign node36013 = (inp[8]) ? node36017 : node36014;
															assign node36014 = (inp[7]) ? 4'b0101 : 4'b0100;
															assign node36017 = (inp[7]) ? 4'b0100 : 4'b0101;
										assign node36020 = (inp[3]) ? node36102 : node36021;
											assign node36021 = (inp[9]) ? node36055 : node36022;
												assign node36022 = (inp[4]) ? node36038 : node36023;
													assign node36023 = (inp[8]) ? node36027 : node36024;
														assign node36024 = (inp[7]) ? 4'b0111 : 4'b0110;
														assign node36027 = (inp[7]) ? node36033 : node36028;
															assign node36028 = (inp[14]) ? 4'b0111 : node36029;
																assign node36029 = (inp[2]) ? 4'b0111 : 4'b0110;
															assign node36033 = (inp[2]) ? 4'b0110 : node36034;
																assign node36034 = (inp[14]) ? 4'b0110 : 4'b0111;
													assign node36038 = (inp[2]) ? node36046 : node36039;
														assign node36039 = (inp[8]) ? 4'b0010 : node36040;
															assign node36040 = (inp[14]) ? 4'b0010 : node36041;
																assign node36041 = (inp[7]) ? 4'b0010 : 4'b0011;
														assign node36046 = (inp[14]) ? 4'b0011 : node36047;
															assign node36047 = (inp[8]) ? node36051 : node36048;
																assign node36048 = (inp[7]) ? 4'b0011 : 4'b0010;
																assign node36051 = (inp[7]) ? 4'b0010 : 4'b0011;
												assign node36055 = (inp[4]) ? node36075 : node36056;
													assign node36056 = (inp[14]) ? node36066 : node36057;
														assign node36057 = (inp[7]) ? 4'b0011 : node36058;
															assign node36058 = (inp[8]) ? node36062 : node36059;
																assign node36059 = (inp[2]) ? 4'b0010 : 4'b0011;
																assign node36062 = (inp[2]) ? 4'b0011 : 4'b0010;
														assign node36066 = (inp[2]) ? node36068 : 4'b0010;
															assign node36068 = (inp[8]) ? node36072 : node36069;
																assign node36069 = (inp[7]) ? 4'b0011 : 4'b0010;
																assign node36072 = (inp[7]) ? 4'b0010 : 4'b0011;
													assign node36075 = (inp[14]) ? node36089 : node36076;
														assign node36076 = (inp[8]) ? node36082 : node36077;
															assign node36077 = (inp[2]) ? 4'b0101 : node36078;
																assign node36078 = (inp[7]) ? 4'b0100 : 4'b0101;
															assign node36082 = (inp[7]) ? node36086 : node36083;
																assign node36083 = (inp[2]) ? 4'b0101 : 4'b0100;
																assign node36086 = (inp[2]) ? 4'b0100 : 4'b0101;
														assign node36089 = (inp[2]) ? node36095 : node36090;
															assign node36090 = (inp[8]) ? 4'b0100 : node36091;
																assign node36091 = (inp[7]) ? 4'b0101 : 4'b0100;
															assign node36095 = (inp[8]) ? node36099 : node36096;
																assign node36096 = (inp[7]) ? 4'b0101 : 4'b0100;
																assign node36099 = (inp[7]) ? 4'b0100 : 4'b0101;
											assign node36102 = (inp[14]) ? node36158 : node36103;
												assign node36103 = (inp[9]) ? node36133 : node36104;
													assign node36104 = (inp[4]) ? node36118 : node36105;
														assign node36105 = (inp[2]) ? node36113 : node36106;
															assign node36106 = (inp[8]) ? node36110 : node36107;
																assign node36107 = (inp[7]) ? 4'b0100 : 4'b0101;
																assign node36110 = (inp[7]) ? 4'b0101 : 4'b0100;
															assign node36113 = (inp[8]) ? node36115 : 4'b0100;
																assign node36115 = (inp[7]) ? 4'b0100 : 4'b0101;
														assign node36118 = (inp[2]) ? node36126 : node36119;
															assign node36119 = (inp[7]) ? node36123 : node36120;
																assign node36120 = (inp[8]) ? 4'b0000 : 4'b0001;
																assign node36123 = (inp[8]) ? 4'b0001 : 4'b0000;
															assign node36126 = (inp[7]) ? node36130 : node36127;
																assign node36127 = (inp[8]) ? 4'b0001 : 4'b0000;
																assign node36130 = (inp[8]) ? 4'b0000 : 4'b0001;
													assign node36133 = (inp[4]) ? node36149 : node36134;
														assign node36134 = (inp[7]) ? node36142 : node36135;
															assign node36135 = (inp[2]) ? node36139 : node36136;
																assign node36136 = (inp[8]) ? 4'b0000 : 4'b0001;
																assign node36139 = (inp[8]) ? 4'b0001 : 4'b0000;
															assign node36142 = (inp[8]) ? node36146 : node36143;
																assign node36143 = (inp[2]) ? 4'b0001 : 4'b0000;
																assign node36146 = (inp[2]) ? 4'b0000 : 4'b0001;
														assign node36149 = (inp[2]) ? node36151 : 4'b0101;
															assign node36151 = (inp[7]) ? node36155 : node36152;
																assign node36152 = (inp[8]) ? 4'b0101 : 4'b0100;
																assign node36155 = (inp[8]) ? 4'b0100 : 4'b0101;
												assign node36158 = (inp[7]) ? node36174 : node36159;
													assign node36159 = (inp[8]) ? node36167 : node36160;
														assign node36160 = (inp[9]) ? node36164 : node36161;
															assign node36161 = (inp[4]) ? 4'b0000 : 4'b0100;
															assign node36164 = (inp[4]) ? 4'b0100 : 4'b0000;
														assign node36167 = (inp[9]) ? node36171 : node36168;
															assign node36168 = (inp[4]) ? 4'b0001 : 4'b0101;
															assign node36171 = (inp[4]) ? 4'b0101 : 4'b0001;
													assign node36174 = (inp[8]) ? node36190 : node36175;
														assign node36175 = (inp[2]) ? node36183 : node36176;
															assign node36176 = (inp[4]) ? node36180 : node36177;
																assign node36177 = (inp[9]) ? 4'b0001 : 4'b0101;
																assign node36180 = (inp[9]) ? 4'b0101 : 4'b0001;
															assign node36183 = (inp[9]) ? node36187 : node36184;
																assign node36184 = (inp[4]) ? 4'b0001 : 4'b0101;
																assign node36187 = (inp[4]) ? 4'b0101 : 4'b0001;
														assign node36190 = (inp[2]) ? 4'b0100 : node36191;
															assign node36191 = (inp[9]) ? 4'b0100 : node36192;
																assign node36192 = (inp[4]) ? 4'b0000 : 4'b0100;
							assign node36197 = (inp[15]) ? node36729 : node36198;
								assign node36198 = (inp[0]) ? node36458 : node36199;
									assign node36199 = (inp[3]) ? node36345 : node36200;
										assign node36200 = (inp[5]) ? node36280 : node36201;
											assign node36201 = (inp[14]) ? node36247 : node36202;
												assign node36202 = (inp[8]) ? node36226 : node36203;
													assign node36203 = (inp[2]) ? node36213 : node36204;
														assign node36204 = (inp[7]) ? node36206 : 4'b0011;
															assign node36206 = (inp[9]) ? node36210 : node36207;
																assign node36207 = (inp[4]) ? 4'b0110 : 4'b0010;
																assign node36210 = (inp[4]) ? 4'b0010 : 4'b0110;
														assign node36213 = (inp[7]) ? node36219 : node36214;
															assign node36214 = (inp[4]) ? node36216 : 4'b0110;
																assign node36216 = (inp[9]) ? 4'b0010 : 4'b0110;
															assign node36219 = (inp[9]) ? node36223 : node36220;
																assign node36220 = (inp[4]) ? 4'b0111 : 4'b0011;
																assign node36223 = (inp[4]) ? 4'b0011 : 4'b0111;
													assign node36226 = (inp[9]) ? node36236 : node36227;
														assign node36227 = (inp[4]) ? node36231 : node36228;
															assign node36228 = (inp[2]) ? 4'b0011 : 4'b0010;
															assign node36231 = (inp[2]) ? 4'b0111 : node36232;
																assign node36232 = (inp[7]) ? 4'b0111 : 4'b0110;
														assign node36236 = (inp[4]) ? node36242 : node36237;
															assign node36237 = (inp[2]) ? node36239 : 4'b0111;
																assign node36239 = (inp[7]) ? 4'b0110 : 4'b0111;
															assign node36242 = (inp[7]) ? node36244 : 4'b0011;
																assign node36244 = (inp[2]) ? 4'b0010 : 4'b0011;
												assign node36247 = (inp[4]) ? node36267 : node36248;
													assign node36248 = (inp[9]) ? node36260 : node36249;
														assign node36249 = (inp[2]) ? node36255 : node36250;
															assign node36250 = (inp[7]) ? node36252 : 4'b0010;
																assign node36252 = (inp[8]) ? 4'b0010 : 4'b0011;
															assign node36255 = (inp[8]) ? 4'b0011 : node36256;
																assign node36256 = (inp[7]) ? 4'b0011 : 4'b0010;
														assign node36260 = (inp[7]) ? node36264 : node36261;
															assign node36261 = (inp[8]) ? 4'b0111 : 4'b0110;
															assign node36264 = (inp[8]) ? 4'b0110 : 4'b0111;
													assign node36267 = (inp[9]) ? node36275 : node36268;
														assign node36268 = (inp[8]) ? node36272 : node36269;
															assign node36269 = (inp[7]) ? 4'b0111 : 4'b0110;
															assign node36272 = (inp[7]) ? 4'b0110 : 4'b0111;
														assign node36275 = (inp[7]) ? 4'b0010 : node36276;
															assign node36276 = (inp[8]) ? 4'b0011 : 4'b0010;
											assign node36280 = (inp[9]) ? node36318 : node36281;
												assign node36281 = (inp[4]) ? node36299 : node36282;
													assign node36282 = (inp[7]) ? node36290 : node36283;
														assign node36283 = (inp[8]) ? node36285 : 4'b0010;
															assign node36285 = (inp[14]) ? 4'b0011 : node36286;
																assign node36286 = (inp[2]) ? 4'b0011 : 4'b0010;
														assign node36290 = (inp[2]) ? node36296 : node36291;
															assign node36291 = (inp[14]) ? 4'b0011 : node36292;
																assign node36292 = (inp[8]) ? 4'b0011 : 4'b0010;
															assign node36296 = (inp[8]) ? 4'b0010 : 4'b0011;
													assign node36299 = (inp[2]) ? node36311 : node36300;
														assign node36300 = (inp[14]) ? node36306 : node36301;
															assign node36301 = (inp[8]) ? node36303 : 4'b0101;
																assign node36303 = (inp[7]) ? 4'b0101 : 4'b0100;
															assign node36306 = (inp[8]) ? 4'b0100 : node36307;
																assign node36307 = (inp[7]) ? 4'b0101 : 4'b0100;
														assign node36311 = (inp[8]) ? node36315 : node36312;
															assign node36312 = (inp[14]) ? 4'b0101 : 4'b0100;
															assign node36315 = (inp[7]) ? 4'b0100 : 4'b0101;
												assign node36318 = (inp[4]) ? node36334 : node36319;
													assign node36319 = (inp[8]) ? node36323 : node36320;
														assign node36320 = (inp[7]) ? 4'b0101 : 4'b0100;
														assign node36323 = (inp[7]) ? node36329 : node36324;
															assign node36324 = (inp[2]) ? 4'b0101 : node36325;
																assign node36325 = (inp[14]) ? 4'b0101 : 4'b0100;
															assign node36329 = (inp[2]) ? 4'b0100 : node36330;
																assign node36330 = (inp[14]) ? 4'b0100 : 4'b0101;
													assign node36334 = (inp[8]) ? node36340 : node36335;
														assign node36335 = (inp[2]) ? node36337 : 4'b0000;
															assign node36337 = (inp[7]) ? 4'b0001 : 4'b0000;
														assign node36340 = (inp[7]) ? node36342 : 4'b0001;
															assign node36342 = (inp[2]) ? 4'b0000 : 4'b0001;
										assign node36345 = (inp[4]) ? node36413 : node36346;
											assign node36346 = (inp[9]) ? node36368 : node36347;
												assign node36347 = (inp[5]) ? node36361 : node36348;
													assign node36348 = (inp[2]) ? node36354 : node36349;
														assign node36349 = (inp[14]) ? node36351 : 4'b0011;
															assign node36351 = (inp[7]) ? 4'b0011 : 4'b0010;
														assign node36354 = (inp[8]) ? node36358 : node36355;
															assign node36355 = (inp[7]) ? 4'b0011 : 4'b0010;
															assign node36358 = (inp[7]) ? 4'b0010 : 4'b0011;
													assign node36361 = (inp[7]) ? 4'b0001 : node36362;
														assign node36362 = (inp[14]) ? 4'b0000 : node36363;
															assign node36363 = (inp[2]) ? 4'b0000 : 4'b0001;
												assign node36368 = (inp[2]) ? node36398 : node36369;
													assign node36369 = (inp[5]) ? node36385 : node36370;
														assign node36370 = (inp[7]) ? node36378 : node36371;
															assign node36371 = (inp[8]) ? node36375 : node36372;
																assign node36372 = (inp[14]) ? 4'b0100 : 4'b0101;
																assign node36375 = (inp[14]) ? 4'b0101 : 4'b0100;
															assign node36378 = (inp[8]) ? node36382 : node36379;
																assign node36379 = (inp[14]) ? 4'b0101 : 4'b0100;
																assign node36382 = (inp[14]) ? 4'b0100 : 4'b0101;
														assign node36385 = (inp[14]) ? node36391 : node36386;
															assign node36386 = (inp[7]) ? node36388 : 4'b0100;
																assign node36388 = (inp[8]) ? 4'b0101 : 4'b0100;
															assign node36391 = (inp[7]) ? node36395 : node36392;
																assign node36392 = (inp[8]) ? 4'b0101 : 4'b0100;
																assign node36395 = (inp[8]) ? 4'b0100 : 4'b0101;
													assign node36398 = (inp[5]) ? node36406 : node36399;
														assign node36399 = (inp[8]) ? node36403 : node36400;
															assign node36400 = (inp[7]) ? 4'b0101 : 4'b0100;
															assign node36403 = (inp[7]) ? 4'b0100 : 4'b0101;
														assign node36406 = (inp[14]) ? 4'b0100 : node36407;
															assign node36407 = (inp[8]) ? node36409 : 4'b0100;
																assign node36409 = (inp[7]) ? 4'b0100 : 4'b0101;
											assign node36413 = (inp[9]) ? node36437 : node36414;
												assign node36414 = (inp[7]) ? node36426 : node36415;
													assign node36415 = (inp[8]) ? node36421 : node36416;
														assign node36416 = (inp[14]) ? 4'b0100 : node36417;
															assign node36417 = (inp[2]) ? 4'b0100 : 4'b0101;
														assign node36421 = (inp[14]) ? 4'b0101 : node36422;
															assign node36422 = (inp[2]) ? 4'b0101 : 4'b0100;
													assign node36426 = (inp[8]) ? node36432 : node36427;
														assign node36427 = (inp[14]) ? 4'b0101 : node36428;
															assign node36428 = (inp[2]) ? 4'b0101 : 4'b0100;
														assign node36432 = (inp[14]) ? 4'b0100 : node36433;
															assign node36433 = (inp[2]) ? 4'b0100 : 4'b0101;
												assign node36437 = (inp[2]) ? node36451 : node36438;
													assign node36438 = (inp[14]) ? node36444 : node36439;
														assign node36439 = (inp[8]) ? 4'b0001 : node36440;
															assign node36440 = (inp[7]) ? 4'b0000 : 4'b0001;
														assign node36444 = (inp[7]) ? node36448 : node36445;
															assign node36445 = (inp[8]) ? 4'b0001 : 4'b0000;
															assign node36448 = (inp[8]) ? 4'b0000 : 4'b0001;
													assign node36451 = (inp[8]) ? node36455 : node36452;
														assign node36452 = (inp[7]) ? 4'b0001 : 4'b0000;
														assign node36455 = (inp[7]) ? 4'b0000 : 4'b0001;
									assign node36458 = (inp[5]) ? node36602 : node36459;
										assign node36459 = (inp[3]) ? node36537 : node36460;
											assign node36460 = (inp[4]) ? node36500 : node36461;
												assign node36461 = (inp[9]) ? node36477 : node36462;
													assign node36462 = (inp[8]) ? node36468 : node36463;
														assign node36463 = (inp[14]) ? node36465 : 4'b0001;
															assign node36465 = (inp[7]) ? 4'b0001 : 4'b0000;
														assign node36468 = (inp[14]) ? 4'b0000 : node36469;
															assign node36469 = (inp[2]) ? node36473 : node36470;
																assign node36470 = (inp[7]) ? 4'b0001 : 4'b0000;
																assign node36473 = (inp[7]) ? 4'b0000 : 4'b0001;
													assign node36477 = (inp[2]) ? node36493 : node36478;
														assign node36478 = (inp[7]) ? node36486 : node36479;
															assign node36479 = (inp[8]) ? node36483 : node36480;
																assign node36480 = (inp[14]) ? 4'b0100 : 4'b0101;
																assign node36483 = (inp[14]) ? 4'b0101 : 4'b0100;
															assign node36486 = (inp[8]) ? node36490 : node36487;
																assign node36487 = (inp[14]) ? 4'b0101 : 4'b0100;
																assign node36490 = (inp[14]) ? 4'b0100 : 4'b0101;
														assign node36493 = (inp[8]) ? node36497 : node36494;
															assign node36494 = (inp[7]) ? 4'b0101 : 4'b0100;
															assign node36497 = (inp[7]) ? 4'b0100 : 4'b0101;
												assign node36500 = (inp[9]) ? node36518 : node36501;
													assign node36501 = (inp[14]) ? node36513 : node36502;
														assign node36502 = (inp[7]) ? node36508 : node36503;
															assign node36503 = (inp[8]) ? node36505 : 4'b0101;
																assign node36505 = (inp[2]) ? 4'b0101 : 4'b0100;
															assign node36508 = (inp[2]) ? 4'b0100 : node36509;
																assign node36509 = (inp[8]) ? 4'b0101 : 4'b0100;
														assign node36513 = (inp[8]) ? 4'b0100 : node36514;
															assign node36514 = (inp[7]) ? 4'b0101 : 4'b0100;
													assign node36518 = (inp[14]) ? node36532 : node36519;
														assign node36519 = (inp[7]) ? node36525 : node36520;
															assign node36520 = (inp[8]) ? 4'b0000 : node36521;
																assign node36521 = (inp[2]) ? 4'b0000 : 4'b0001;
															assign node36525 = (inp[2]) ? node36529 : node36526;
																assign node36526 = (inp[8]) ? 4'b0001 : 4'b0000;
																assign node36529 = (inp[8]) ? 4'b0000 : 4'b0001;
														assign node36532 = (inp[8]) ? 4'b0001 : node36533;
															assign node36533 = (inp[2]) ? 4'b0001 : 4'b0000;
											assign node36537 = (inp[9]) ? node36571 : node36538;
												assign node36538 = (inp[4]) ? node36554 : node36539;
													assign node36539 = (inp[7]) ? node36547 : node36540;
														assign node36540 = (inp[8]) ? node36544 : node36541;
															assign node36541 = (inp[14]) ? 4'b0000 : 4'b0001;
															assign node36544 = (inp[14]) ? 4'b0001 : 4'b0000;
														assign node36547 = (inp[8]) ? node36549 : 4'b0001;
															assign node36549 = (inp[14]) ? 4'b0000 : node36550;
																assign node36550 = (inp[2]) ? 4'b0000 : 4'b0001;
													assign node36554 = (inp[7]) ? node36564 : node36555;
														assign node36555 = (inp[14]) ? node36561 : node36556;
															assign node36556 = (inp[2]) ? 4'b0110 : node36557;
																assign node36557 = (inp[8]) ? 4'b0110 : 4'b0111;
															assign node36561 = (inp[8]) ? 4'b0111 : 4'b0110;
														assign node36564 = (inp[2]) ? 4'b0111 : node36565;
															assign node36565 = (inp[14]) ? 4'b0111 : node36566;
																assign node36566 = (inp[8]) ? 4'b0111 : 4'b0110;
												assign node36571 = (inp[4]) ? node36589 : node36572;
													assign node36572 = (inp[8]) ? node36578 : node36573;
														assign node36573 = (inp[7]) ? node36575 : 4'b0110;
															assign node36575 = (inp[2]) ? 4'b0111 : 4'b0110;
														assign node36578 = (inp[7]) ? node36584 : node36579;
															assign node36579 = (inp[2]) ? 4'b0111 : node36580;
																assign node36580 = (inp[14]) ? 4'b0111 : 4'b0110;
															assign node36584 = (inp[14]) ? 4'b0110 : node36585;
																assign node36585 = (inp[2]) ? 4'b0110 : 4'b0111;
													assign node36589 = (inp[14]) ? node36595 : node36590;
														assign node36590 = (inp[7]) ? 4'b0011 : node36591;
															assign node36591 = (inp[2]) ? 4'b0011 : 4'b0010;
														assign node36595 = (inp[7]) ? node36599 : node36596;
															assign node36596 = (inp[8]) ? 4'b0011 : 4'b0010;
															assign node36599 = (inp[8]) ? 4'b0010 : 4'b0011;
										assign node36602 = (inp[4]) ? node36670 : node36603;
											assign node36603 = (inp[9]) ? node36645 : node36604;
												assign node36604 = (inp[3]) ? node36620 : node36605;
													assign node36605 = (inp[2]) ? node36615 : node36606;
														assign node36606 = (inp[8]) ? node36608 : 4'b0001;
															assign node36608 = (inp[7]) ? node36612 : node36609;
																assign node36609 = (inp[14]) ? 4'b0001 : 4'b0000;
																assign node36612 = (inp[14]) ? 4'b0000 : 4'b0001;
														assign node36615 = (inp[7]) ? 4'b0000 : node36616;
															assign node36616 = (inp[8]) ? 4'b0001 : 4'b0000;
													assign node36620 = (inp[2]) ? node36636 : node36621;
														assign node36621 = (inp[7]) ? node36629 : node36622;
															assign node36622 = (inp[14]) ? node36626 : node36623;
																assign node36623 = (inp[8]) ? 4'b0010 : 4'b0011;
																assign node36626 = (inp[8]) ? 4'b0011 : 4'b0010;
															assign node36629 = (inp[14]) ? node36633 : node36630;
																assign node36630 = (inp[8]) ? 4'b0011 : 4'b0010;
																assign node36633 = (inp[8]) ? 4'b0010 : 4'b0011;
														assign node36636 = (inp[14]) ? 4'b0010 : node36637;
															assign node36637 = (inp[8]) ? node36641 : node36638;
																assign node36638 = (inp[7]) ? 4'b0011 : 4'b0010;
																assign node36641 = (inp[7]) ? 4'b0010 : 4'b0011;
												assign node36645 = (inp[8]) ? node36659 : node36646;
													assign node36646 = (inp[3]) ? node36648 : 4'b0110;
														assign node36648 = (inp[7]) ? node36654 : node36649;
															assign node36649 = (inp[14]) ? 4'b0110 : node36650;
																assign node36650 = (inp[2]) ? 4'b0110 : 4'b0111;
															assign node36654 = (inp[14]) ? 4'b0111 : node36655;
																assign node36655 = (inp[2]) ? 4'b0111 : 4'b0110;
													assign node36659 = (inp[7]) ? node36665 : node36660;
														assign node36660 = (inp[2]) ? 4'b0111 : node36661;
															assign node36661 = (inp[14]) ? 4'b0111 : 4'b0110;
														assign node36665 = (inp[3]) ? node36667 : 4'b0110;
															assign node36667 = (inp[2]) ? 4'b0110 : 4'b0111;
											assign node36670 = (inp[9]) ? node36706 : node36671;
												assign node36671 = (inp[3]) ? node36687 : node36672;
													assign node36672 = (inp[8]) ? node36676 : node36673;
														assign node36673 = (inp[7]) ? 4'b0111 : 4'b0110;
														assign node36676 = (inp[7]) ? node36682 : node36677;
															assign node36677 = (inp[2]) ? 4'b0111 : node36678;
																assign node36678 = (inp[14]) ? 4'b0111 : 4'b0110;
															assign node36682 = (inp[14]) ? 4'b0110 : node36683;
																assign node36683 = (inp[2]) ? 4'b0110 : 4'b0111;
													assign node36687 = (inp[8]) ? node36695 : node36688;
														assign node36688 = (inp[2]) ? 4'b0111 : node36689;
															assign node36689 = (inp[7]) ? node36691 : 4'b0111;
																assign node36691 = (inp[14]) ? 4'b0111 : 4'b0110;
														assign node36695 = (inp[7]) ? node36701 : node36696;
															assign node36696 = (inp[14]) ? 4'b0111 : node36697;
																assign node36697 = (inp[2]) ? 4'b0111 : 4'b0110;
															assign node36701 = (inp[14]) ? 4'b0110 : node36702;
																assign node36702 = (inp[2]) ? 4'b0110 : 4'b0111;
												assign node36706 = (inp[8]) ? node36718 : node36707;
													assign node36707 = (inp[7]) ? node36713 : node36708;
														assign node36708 = (inp[14]) ? 4'b0010 : node36709;
															assign node36709 = (inp[2]) ? 4'b0010 : 4'b0011;
														assign node36713 = (inp[14]) ? 4'b0011 : node36714;
															assign node36714 = (inp[2]) ? 4'b0011 : 4'b0010;
													assign node36718 = (inp[7]) ? node36724 : node36719;
														assign node36719 = (inp[14]) ? 4'b0011 : node36720;
															assign node36720 = (inp[2]) ? 4'b0011 : 4'b0010;
														assign node36724 = (inp[14]) ? 4'b0010 : node36725;
															assign node36725 = (inp[2]) ? 4'b0010 : 4'b0011;
								assign node36729 = (inp[0]) ? node37089 : node36730;
									assign node36730 = (inp[5]) ? node36890 : node36731;
										assign node36731 = (inp[3]) ? node36801 : node36732;
											assign node36732 = (inp[4]) ? node36762 : node36733;
												assign node36733 = (inp[9]) ? node36749 : node36734;
													assign node36734 = (inp[7]) ? node36742 : node36735;
														assign node36735 = (inp[8]) ? 4'b0001 : node36736;
															assign node36736 = (inp[2]) ? 4'b0000 : node36737;
																assign node36737 = (inp[14]) ? 4'b0000 : 4'b0001;
														assign node36742 = (inp[2]) ? node36746 : node36743;
															assign node36743 = (inp[8]) ? 4'b0001 : 4'b0000;
															assign node36746 = (inp[8]) ? 4'b0000 : 4'b0001;
													assign node36749 = (inp[7]) ? 4'b0101 : node36750;
														assign node36750 = (inp[8]) ? node36756 : node36751;
															assign node36751 = (inp[14]) ? 4'b0100 : node36752;
																assign node36752 = (inp[2]) ? 4'b0100 : 4'b0101;
															assign node36756 = (inp[2]) ? 4'b0101 : node36757;
																assign node36757 = (inp[14]) ? 4'b0101 : 4'b0100;
												assign node36762 = (inp[9]) ? node36780 : node36763;
													assign node36763 = (inp[2]) ? node36773 : node36764;
														assign node36764 = (inp[8]) ? 4'b0100 : node36765;
															assign node36765 = (inp[7]) ? node36769 : node36766;
																assign node36766 = (inp[14]) ? 4'b0100 : 4'b0101;
																assign node36769 = (inp[14]) ? 4'b0101 : 4'b0100;
														assign node36773 = (inp[14]) ? 4'b0101 : node36774;
															assign node36774 = (inp[7]) ? node36776 : 4'b0101;
																assign node36776 = (inp[8]) ? 4'b0100 : 4'b0101;
													assign node36780 = (inp[2]) ? node36792 : node36781;
														assign node36781 = (inp[14]) ? node36787 : node36782;
															assign node36782 = (inp[8]) ? node36784 : 4'b0001;
																assign node36784 = (inp[7]) ? 4'b0001 : 4'b0000;
															assign node36787 = (inp[8]) ? node36789 : 4'b0000;
																assign node36789 = (inp[7]) ? 4'b0000 : 4'b0001;
														assign node36792 = (inp[14]) ? node36798 : node36793;
															assign node36793 = (inp[7]) ? 4'b0000 : node36794;
																assign node36794 = (inp[8]) ? 4'b0001 : 4'b0000;
															assign node36798 = (inp[8]) ? 4'b0000 : 4'b0001;
											assign node36801 = (inp[9]) ? node36839 : node36802;
												assign node36802 = (inp[4]) ? node36822 : node36803;
													assign node36803 = (inp[7]) ? node36813 : node36804;
														assign node36804 = (inp[8]) ? node36808 : node36805;
															assign node36805 = (inp[14]) ? 4'b0000 : 4'b0001;
															assign node36808 = (inp[14]) ? 4'b0001 : node36809;
																assign node36809 = (inp[2]) ? 4'b0001 : 4'b0000;
														assign node36813 = (inp[8]) ? node36817 : node36814;
															assign node36814 = (inp[14]) ? 4'b0001 : 4'b0000;
															assign node36817 = (inp[2]) ? 4'b0000 : node36818;
																assign node36818 = (inp[14]) ? 4'b0000 : 4'b0001;
													assign node36822 = (inp[8]) ? node36830 : node36823;
														assign node36823 = (inp[7]) ? node36825 : 4'b0110;
															assign node36825 = (inp[2]) ? 4'b0111 : node36826;
																assign node36826 = (inp[14]) ? 4'b0111 : 4'b0110;
														assign node36830 = (inp[7]) ? node36836 : node36831;
															assign node36831 = (inp[14]) ? 4'b0111 : node36832;
																assign node36832 = (inp[2]) ? 4'b0111 : 4'b0110;
															assign node36836 = (inp[14]) ? 4'b0110 : 4'b0111;
												assign node36839 = (inp[4]) ? node36869 : node36840;
													assign node36840 = (inp[14]) ? node36854 : node36841;
														assign node36841 = (inp[7]) ? node36849 : node36842;
															assign node36842 = (inp[8]) ? node36846 : node36843;
																assign node36843 = (inp[2]) ? 4'b0110 : 4'b0111;
																assign node36846 = (inp[2]) ? 4'b0111 : 4'b0110;
															assign node36849 = (inp[2]) ? 4'b0110 : node36850;
																assign node36850 = (inp[8]) ? 4'b0111 : 4'b0110;
														assign node36854 = (inp[2]) ? node36862 : node36855;
															assign node36855 = (inp[7]) ? node36859 : node36856;
																assign node36856 = (inp[8]) ? 4'b0111 : 4'b0110;
																assign node36859 = (inp[8]) ? 4'b0110 : 4'b0111;
															assign node36862 = (inp[8]) ? node36866 : node36863;
																assign node36863 = (inp[7]) ? 4'b0111 : 4'b0110;
																assign node36866 = (inp[7]) ? 4'b0110 : 4'b0111;
													assign node36869 = (inp[14]) ? node36883 : node36870;
														assign node36870 = (inp[7]) ? node36878 : node36871;
															assign node36871 = (inp[8]) ? node36875 : node36872;
																assign node36872 = (inp[2]) ? 4'b0010 : 4'b0011;
																assign node36875 = (inp[2]) ? 4'b0011 : 4'b0010;
															assign node36878 = (inp[8]) ? node36880 : 4'b0010;
																assign node36880 = (inp[2]) ? 4'b0010 : 4'b0011;
														assign node36883 = (inp[7]) ? node36887 : node36884;
															assign node36884 = (inp[8]) ? 4'b0011 : 4'b0010;
															assign node36887 = (inp[8]) ? 4'b0010 : 4'b0011;
										assign node36890 = (inp[3]) ? node36988 : node36891;
											assign node36891 = (inp[4]) ? node36941 : node36892;
												assign node36892 = (inp[9]) ? node36914 : node36893;
													assign node36893 = (inp[2]) ? node36907 : node36894;
														assign node36894 = (inp[14]) ? node36900 : node36895;
															assign node36895 = (inp[8]) ? 4'b0000 : node36896;
																assign node36896 = (inp[7]) ? 4'b0000 : 4'b0001;
															assign node36900 = (inp[8]) ? node36904 : node36901;
																assign node36901 = (inp[7]) ? 4'b0001 : 4'b0000;
																assign node36904 = (inp[7]) ? 4'b0000 : 4'b0001;
														assign node36907 = (inp[7]) ? node36911 : node36908;
															assign node36908 = (inp[8]) ? 4'b0001 : 4'b0000;
															assign node36911 = (inp[8]) ? 4'b0000 : 4'b0001;
													assign node36914 = (inp[2]) ? node36928 : node36915;
														assign node36915 = (inp[7]) ? node36923 : node36916;
															assign node36916 = (inp[8]) ? node36920 : node36917;
																assign node36917 = (inp[14]) ? 4'b0110 : 4'b0111;
																assign node36920 = (inp[14]) ? 4'b0111 : 4'b0110;
															assign node36923 = (inp[8]) ? 4'b0110 : node36924;
																assign node36924 = (inp[14]) ? 4'b0111 : 4'b0110;
														assign node36928 = (inp[14]) ? node36934 : node36929;
															assign node36929 = (inp[7]) ? 4'b0111 : node36930;
																assign node36930 = (inp[8]) ? 4'b0111 : 4'b0110;
															assign node36934 = (inp[8]) ? node36938 : node36935;
																assign node36935 = (inp[7]) ? 4'b0111 : 4'b0110;
																assign node36938 = (inp[7]) ? 4'b0110 : 4'b0111;
												assign node36941 = (inp[9]) ? node36963 : node36942;
													assign node36942 = (inp[7]) ? node36952 : node36943;
														assign node36943 = (inp[14]) ? 4'b0111 : node36944;
															assign node36944 = (inp[8]) ? node36948 : node36945;
																assign node36945 = (inp[2]) ? 4'b0110 : 4'b0111;
																assign node36948 = (inp[2]) ? 4'b0111 : 4'b0110;
														assign node36952 = (inp[8]) ? node36958 : node36953;
															assign node36953 = (inp[2]) ? 4'b0111 : node36954;
																assign node36954 = (inp[14]) ? 4'b0111 : 4'b0110;
															assign node36958 = (inp[14]) ? 4'b0110 : node36959;
																assign node36959 = (inp[2]) ? 4'b0110 : 4'b0111;
													assign node36963 = (inp[2]) ? node36977 : node36964;
														assign node36964 = (inp[14]) ? node36972 : node36965;
															assign node36965 = (inp[7]) ? node36969 : node36966;
																assign node36966 = (inp[8]) ? 4'b0010 : 4'b0011;
																assign node36969 = (inp[8]) ? 4'b0011 : 4'b0010;
															assign node36972 = (inp[7]) ? node36974 : 4'b0010;
																assign node36974 = (inp[8]) ? 4'b0010 : 4'b0011;
														assign node36977 = (inp[14]) ? node36983 : node36978;
															assign node36978 = (inp[7]) ? node36980 : 4'b0011;
																assign node36980 = (inp[8]) ? 4'b0010 : 4'b0011;
															assign node36983 = (inp[8]) ? 4'b0011 : node36984;
																assign node36984 = (inp[7]) ? 4'b0011 : 4'b0010;
											assign node36988 = (inp[2]) ? node37034 : node36989;
												assign node36989 = (inp[8]) ? node37015 : node36990;
													assign node36990 = (inp[7]) ? node37004 : node36991;
														assign node36991 = (inp[14]) ? node36999 : node36992;
															assign node36992 = (inp[9]) ? node36996 : node36993;
																assign node36993 = (inp[4]) ? 4'b0111 : 4'b0011;
																assign node36996 = (inp[4]) ? 4'b0011 : 4'b0111;
															assign node36999 = (inp[4]) ? node37001 : 4'b0110;
																assign node37001 = (inp[9]) ? 4'b0010 : 4'b0110;
														assign node37004 = (inp[14]) ? node37010 : node37005;
															assign node37005 = (inp[9]) ? node37007 : 4'b0010;
																assign node37007 = (inp[4]) ? 4'b0010 : 4'b0110;
															assign node37010 = (inp[4]) ? node37012 : 4'b0011;
																assign node37012 = (inp[9]) ? 4'b0011 : 4'b0111;
													assign node37015 = (inp[4]) ? node37027 : node37016;
														assign node37016 = (inp[9]) ? node37024 : node37017;
															assign node37017 = (inp[7]) ? node37021 : node37018;
																assign node37018 = (inp[14]) ? 4'b0011 : 4'b0010;
																assign node37021 = (inp[14]) ? 4'b0010 : 4'b0011;
															assign node37024 = (inp[7]) ? 4'b0111 : 4'b0110;
														assign node37027 = (inp[9]) ? node37029 : 4'b0110;
															assign node37029 = (inp[14]) ? node37031 : 4'b0010;
																assign node37031 = (inp[7]) ? 4'b0010 : 4'b0011;
												assign node37034 = (inp[14]) ? node37062 : node37035;
													assign node37035 = (inp[7]) ? node37051 : node37036;
														assign node37036 = (inp[8]) ? node37044 : node37037;
															assign node37037 = (inp[4]) ? node37041 : node37038;
																assign node37038 = (inp[9]) ? 4'b0110 : 4'b0010;
																assign node37041 = (inp[9]) ? 4'b0010 : 4'b0110;
															assign node37044 = (inp[9]) ? node37048 : node37045;
																assign node37045 = (inp[4]) ? 4'b0111 : 4'b0011;
																assign node37048 = (inp[4]) ? 4'b0011 : 4'b0111;
														assign node37051 = (inp[8]) ? node37059 : node37052;
															assign node37052 = (inp[9]) ? node37056 : node37053;
																assign node37053 = (inp[4]) ? 4'b0111 : 4'b0011;
																assign node37056 = (inp[4]) ? 4'b0011 : 4'b0111;
															assign node37059 = (inp[9]) ? 4'b0010 : 4'b0110;
													assign node37062 = (inp[9]) ? node37078 : node37063;
														assign node37063 = (inp[4]) ? node37071 : node37064;
															assign node37064 = (inp[8]) ? node37068 : node37065;
																assign node37065 = (inp[7]) ? 4'b0011 : 4'b0010;
																assign node37068 = (inp[7]) ? 4'b0010 : 4'b0011;
															assign node37071 = (inp[7]) ? node37075 : node37072;
																assign node37072 = (inp[8]) ? 4'b0111 : 4'b0110;
																assign node37075 = (inp[8]) ? 4'b0110 : 4'b0111;
														assign node37078 = (inp[4]) ? node37084 : node37079;
															assign node37079 = (inp[8]) ? node37081 : 4'b0110;
																assign node37081 = (inp[7]) ? 4'b0110 : 4'b0111;
															assign node37084 = (inp[8]) ? 4'b0010 : node37085;
																assign node37085 = (inp[7]) ? 4'b0011 : 4'b0010;
									assign node37089 = (inp[5]) ? node37233 : node37090;
										assign node37090 = (inp[3]) ? node37176 : node37091;
											assign node37091 = (inp[7]) ? node37127 : node37092;
												assign node37092 = (inp[8]) ? node37110 : node37093;
													assign node37093 = (inp[14]) ? node37103 : node37094;
														assign node37094 = (inp[2]) ? 4'b0110 : node37095;
															assign node37095 = (inp[9]) ? node37099 : node37096;
																assign node37096 = (inp[4]) ? 4'b0111 : 4'b0011;
																assign node37099 = (inp[4]) ? 4'b0011 : 4'b0111;
														assign node37103 = (inp[4]) ? node37107 : node37104;
															assign node37104 = (inp[9]) ? 4'b0110 : 4'b0010;
															assign node37107 = (inp[9]) ? 4'b0010 : 4'b0110;
													assign node37110 = (inp[2]) ? node37120 : node37111;
														assign node37111 = (inp[14]) ? 4'b0111 : node37112;
															assign node37112 = (inp[9]) ? node37116 : node37113;
																assign node37113 = (inp[4]) ? 4'b0110 : 4'b0010;
																assign node37116 = (inp[4]) ? 4'b0010 : 4'b0110;
														assign node37120 = (inp[4]) ? node37124 : node37121;
															assign node37121 = (inp[9]) ? 4'b0111 : 4'b0011;
															assign node37124 = (inp[9]) ? 4'b0011 : 4'b0111;
												assign node37127 = (inp[8]) ? node37155 : node37128;
													assign node37128 = (inp[14]) ? node37140 : node37129;
														assign node37129 = (inp[2]) ? node37135 : node37130;
															assign node37130 = (inp[4]) ? node37132 : 4'b0010;
																assign node37132 = (inp[9]) ? 4'b0010 : 4'b0110;
															assign node37135 = (inp[4]) ? node37137 : 4'b0111;
																assign node37137 = (inp[9]) ? 4'b0011 : 4'b0111;
														assign node37140 = (inp[2]) ? node37148 : node37141;
															assign node37141 = (inp[9]) ? node37145 : node37142;
																assign node37142 = (inp[4]) ? 4'b0111 : 4'b0011;
																assign node37145 = (inp[4]) ? 4'b0011 : 4'b0111;
															assign node37148 = (inp[4]) ? node37152 : node37149;
																assign node37149 = (inp[9]) ? 4'b0111 : 4'b0011;
																assign node37152 = (inp[9]) ? 4'b0011 : 4'b0111;
													assign node37155 = (inp[14]) ? node37169 : node37156;
														assign node37156 = (inp[2]) ? node37164 : node37157;
															assign node37157 = (inp[9]) ? node37161 : node37158;
																assign node37158 = (inp[4]) ? 4'b0111 : 4'b0011;
																assign node37161 = (inp[4]) ? 4'b0011 : 4'b0111;
															assign node37164 = (inp[9]) ? node37166 : 4'b0110;
																assign node37166 = (inp[4]) ? 4'b0010 : 4'b0110;
														assign node37169 = (inp[2]) ? 4'b0010 : node37170;
															assign node37170 = (inp[9]) ? 4'b0110 : node37171;
																assign node37171 = (inp[4]) ? 4'b0110 : 4'b0010;
											assign node37176 = (inp[4]) ? node37202 : node37177;
												assign node37177 = (inp[9]) ? node37193 : node37178;
													assign node37178 = (inp[8]) ? node37182 : node37179;
														assign node37179 = (inp[7]) ? 4'b0011 : 4'b0010;
														assign node37182 = (inp[7]) ? node37188 : node37183;
															assign node37183 = (inp[14]) ? 4'b0011 : node37184;
																assign node37184 = (inp[2]) ? 4'b0011 : 4'b0010;
															assign node37188 = (inp[14]) ? 4'b0010 : node37189;
																assign node37189 = (inp[2]) ? 4'b0010 : 4'b0011;
													assign node37193 = (inp[2]) ? node37195 : 4'b0100;
														assign node37195 = (inp[14]) ? 4'b0101 : node37196;
															assign node37196 = (inp[7]) ? node37198 : 4'b0100;
																assign node37198 = (inp[8]) ? 4'b0100 : 4'b0101;
												assign node37202 = (inp[9]) ? node37220 : node37203;
													assign node37203 = (inp[7]) ? node37211 : node37204;
														assign node37204 = (inp[8]) ? 4'b0101 : node37205;
															assign node37205 = (inp[14]) ? 4'b0100 : node37206;
																assign node37206 = (inp[2]) ? 4'b0100 : 4'b0101;
														assign node37211 = (inp[8]) ? node37215 : node37212;
															assign node37212 = (inp[2]) ? 4'b0101 : 4'b0100;
															assign node37215 = (inp[2]) ? 4'b0100 : node37216;
																assign node37216 = (inp[14]) ? 4'b0100 : 4'b0101;
													assign node37220 = (inp[7]) ? node37228 : node37221;
														assign node37221 = (inp[8]) ? 4'b0001 : node37222;
															assign node37222 = (inp[2]) ? 4'b0000 : node37223;
																assign node37223 = (inp[14]) ? 4'b0000 : 4'b0001;
														assign node37228 = (inp[2]) ? node37230 : 4'b0000;
															assign node37230 = (inp[8]) ? 4'b0000 : 4'b0001;
										assign node37233 = (inp[9]) ? node37301 : node37234;
											assign node37234 = (inp[4]) ? node37266 : node37235;
												assign node37235 = (inp[3]) ? node37251 : node37236;
													assign node37236 = (inp[7]) ? node37244 : node37237;
														assign node37237 = (inp[8]) ? node37239 : 4'b0010;
															assign node37239 = (inp[2]) ? 4'b0011 : node37240;
																assign node37240 = (inp[14]) ? 4'b0011 : 4'b0010;
														assign node37244 = (inp[8]) ? node37246 : 4'b0011;
															assign node37246 = (inp[14]) ? 4'b0010 : node37247;
																assign node37247 = (inp[2]) ? 4'b0010 : 4'b0011;
													assign node37251 = (inp[14]) ? node37259 : node37252;
														assign node37252 = (inp[2]) ? node37254 : 4'b0001;
															assign node37254 = (inp[8]) ? node37256 : 4'b0001;
																assign node37256 = (inp[7]) ? 4'b0000 : 4'b0001;
														assign node37259 = (inp[8]) ? node37263 : node37260;
															assign node37260 = (inp[7]) ? 4'b0001 : 4'b0000;
															assign node37263 = (inp[7]) ? 4'b0000 : 4'b0001;
												assign node37266 = (inp[3]) ? node37286 : node37267;
													assign node37267 = (inp[7]) ? node37279 : node37268;
														assign node37268 = (inp[8]) ? node37274 : node37269;
															assign node37269 = (inp[14]) ? 4'b0100 : node37270;
																assign node37270 = (inp[2]) ? 4'b0100 : 4'b0101;
															assign node37274 = (inp[2]) ? 4'b0101 : node37275;
																assign node37275 = (inp[14]) ? 4'b0101 : 4'b0100;
														assign node37279 = (inp[8]) ? 4'b0100 : node37280;
															assign node37280 = (inp[2]) ? 4'b0101 : node37281;
																assign node37281 = (inp[14]) ? 4'b0101 : 4'b0100;
													assign node37286 = (inp[8]) ? node37292 : node37287;
														assign node37287 = (inp[7]) ? 4'b0101 : node37288;
															assign node37288 = (inp[2]) ? 4'b0100 : 4'b0101;
														assign node37292 = (inp[7]) ? node37298 : node37293;
															assign node37293 = (inp[14]) ? 4'b0101 : node37294;
																assign node37294 = (inp[2]) ? 4'b0101 : 4'b0100;
															assign node37298 = (inp[14]) ? 4'b0100 : 4'b0101;
											assign node37301 = (inp[4]) ? node37333 : node37302;
												assign node37302 = (inp[2]) ? node37326 : node37303;
													assign node37303 = (inp[14]) ? node37313 : node37304;
														assign node37304 = (inp[3]) ? 4'b0101 : node37305;
															assign node37305 = (inp[7]) ? node37309 : node37306;
																assign node37306 = (inp[8]) ? 4'b0100 : 4'b0101;
																assign node37309 = (inp[8]) ? 4'b0101 : 4'b0100;
														assign node37313 = (inp[3]) ? node37319 : node37314;
															assign node37314 = (inp[7]) ? node37316 : 4'b0101;
																assign node37316 = (inp[8]) ? 4'b0100 : 4'b0101;
															assign node37319 = (inp[8]) ? node37323 : node37320;
																assign node37320 = (inp[7]) ? 4'b0101 : 4'b0100;
																assign node37323 = (inp[7]) ? 4'b0100 : 4'b0101;
													assign node37326 = (inp[8]) ? node37330 : node37327;
														assign node37327 = (inp[7]) ? 4'b0101 : 4'b0100;
														assign node37330 = (inp[7]) ? 4'b0100 : 4'b0101;
												assign node37333 = (inp[3]) ? node37361 : node37334;
													assign node37334 = (inp[14]) ? node37350 : node37335;
														assign node37335 = (inp[8]) ? node37343 : node37336;
															assign node37336 = (inp[7]) ? node37340 : node37337;
																assign node37337 = (inp[2]) ? 4'b0000 : 4'b0001;
																assign node37340 = (inp[2]) ? 4'b0001 : 4'b0000;
															assign node37343 = (inp[7]) ? node37347 : node37344;
																assign node37344 = (inp[2]) ? 4'b0001 : 4'b0000;
																assign node37347 = (inp[2]) ? 4'b0000 : 4'b0001;
														assign node37350 = (inp[2]) ? node37356 : node37351;
															assign node37351 = (inp[7]) ? node37353 : 4'b0000;
																assign node37353 = (inp[8]) ? 4'b0000 : 4'b0001;
															assign node37356 = (inp[8]) ? node37358 : 4'b0000;
																assign node37358 = (inp[7]) ? 4'b0000 : 4'b0001;
													assign node37361 = (inp[2]) ? node37371 : node37362;
														assign node37362 = (inp[7]) ? 4'b0001 : node37363;
															assign node37363 = (inp[8]) ? node37367 : node37364;
																assign node37364 = (inp[14]) ? 4'b0000 : 4'b0001;
																assign node37367 = (inp[14]) ? 4'b0001 : 4'b0000;
														assign node37371 = (inp[14]) ? node37377 : node37372;
															assign node37372 = (inp[7]) ? node37374 : 4'b0000;
																assign node37374 = (inp[8]) ? 4'b0000 : 4'b0001;
															assign node37377 = (inp[8]) ? node37379 : 4'b0001;
																assign node37379 = (inp[7]) ? 4'b0000 : 4'b0001;
					assign node37382 = (inp[7]) ? node39416 : node37383;
						assign node37383 = (inp[8]) ? node38377 : node37384;
							assign node37384 = (inp[14]) ? node37948 : node37385;
								assign node37385 = (inp[2]) ? node37687 : node37386;
									assign node37386 = (inp[5]) ? node37532 : node37387;
										assign node37387 = (inp[12]) ? node37425 : node37388;
											assign node37388 = (inp[4]) ? node37404 : node37389;
												assign node37389 = (inp[9]) ? node37397 : node37390;
													assign node37390 = (inp[15]) ? node37394 : node37391;
														assign node37391 = (inp[0]) ? 4'b0101 : 4'b0111;
														assign node37394 = (inp[0]) ? 4'b0111 : 4'b0101;
													assign node37397 = (inp[0]) ? node37401 : node37398;
														assign node37398 = (inp[15]) ? 4'b0001 : 4'b0011;
														assign node37401 = (inp[15]) ? 4'b0011 : 4'b0001;
												assign node37404 = (inp[9]) ? node37412 : node37405;
													assign node37405 = (inp[15]) ? node37409 : node37406;
														assign node37406 = (inp[0]) ? 4'b0001 : 4'b0011;
														assign node37409 = (inp[0]) ? 4'b0011 : 4'b0001;
													assign node37412 = (inp[3]) ? node37418 : node37413;
														assign node37413 = (inp[0]) ? 4'b0101 : node37414;
															assign node37414 = (inp[15]) ? 4'b0101 : 4'b0111;
														assign node37418 = (inp[10]) ? node37422 : node37419;
															assign node37419 = (inp[0]) ? 4'b0111 : 4'b0101;
															assign node37422 = (inp[0]) ? 4'b0101 : 4'b0111;
											assign node37425 = (inp[15]) ? node37477 : node37426;
												assign node37426 = (inp[0]) ? node37450 : node37427;
													assign node37427 = (inp[3]) ? node37441 : node37428;
														assign node37428 = (inp[9]) ? node37434 : node37429;
															assign node37429 = (inp[10]) ? 4'b0011 : node37430;
																assign node37430 = (inp[4]) ? 4'b0011 : 4'b0111;
															assign node37434 = (inp[4]) ? node37438 : node37435;
																assign node37435 = (inp[10]) ? 4'b0111 : 4'b0011;
																assign node37438 = (inp[10]) ? 4'b0011 : 4'b0111;
														assign node37441 = (inp[10]) ? 4'b0101 : node37442;
															assign node37442 = (inp[4]) ? node37446 : node37443;
																assign node37443 = (inp[9]) ? 4'b0011 : 4'b0111;
																assign node37446 = (inp[9]) ? 4'b0101 : 4'b0011;
													assign node37450 = (inp[3]) ? node37462 : node37451;
														assign node37451 = (inp[9]) ? node37457 : node37452;
															assign node37452 = (inp[10]) ? 4'b0101 : node37453;
																assign node37453 = (inp[4]) ? 4'b0001 : 4'b0101;
															assign node37457 = (inp[10]) ? 4'b0001 : node37458;
																assign node37458 = (inp[4]) ? 4'b0101 : 4'b0001;
														assign node37462 = (inp[9]) ? node37470 : node37463;
															assign node37463 = (inp[10]) ? node37467 : node37464;
																assign node37464 = (inp[4]) ? 4'b0001 : 4'b0101;
																assign node37467 = (inp[4]) ? 4'b0111 : 4'b0001;
															assign node37470 = (inp[4]) ? node37474 : node37471;
																assign node37471 = (inp[10]) ? 4'b0111 : 4'b0001;
																assign node37474 = (inp[10]) ? 4'b0011 : 4'b0111;
												assign node37477 = (inp[0]) ? node37509 : node37478;
													assign node37478 = (inp[3]) ? node37494 : node37479;
														assign node37479 = (inp[10]) ? node37487 : node37480;
															assign node37480 = (inp[4]) ? node37484 : node37481;
																assign node37481 = (inp[9]) ? 4'b0001 : 4'b0101;
																assign node37484 = (inp[9]) ? 4'b0101 : 4'b0001;
															assign node37487 = (inp[9]) ? node37491 : node37488;
																assign node37488 = (inp[4]) ? 4'b0101 : 4'b0001;
																assign node37491 = (inp[4]) ? 4'b0001 : 4'b0101;
														assign node37494 = (inp[9]) ? node37502 : node37495;
															assign node37495 = (inp[4]) ? node37499 : node37496;
																assign node37496 = (inp[10]) ? 4'b0001 : 4'b0101;
																assign node37499 = (inp[10]) ? 4'b0111 : 4'b0001;
															assign node37502 = (inp[10]) ? node37506 : node37503;
																assign node37503 = (inp[4]) ? 4'b0111 : 4'b0001;
																assign node37506 = (inp[4]) ? 4'b0011 : 4'b0111;
													assign node37509 = (inp[3]) ? node37519 : node37510;
														assign node37510 = (inp[9]) ? 4'b0111 : node37511;
															assign node37511 = (inp[10]) ? node37515 : node37512;
																assign node37512 = (inp[4]) ? 4'b0011 : 4'b0111;
																assign node37515 = (inp[4]) ? 4'b0111 : 4'b0011;
														assign node37519 = (inp[9]) ? node37525 : node37520;
															assign node37520 = (inp[10]) ? node37522 : 4'b0011;
																assign node37522 = (inp[4]) ? 4'b0101 : 4'b0011;
															assign node37525 = (inp[10]) ? node37529 : node37526;
																assign node37526 = (inp[4]) ? 4'b0101 : 4'b0011;
																assign node37529 = (inp[4]) ? 4'b0001 : 4'b0101;
										assign node37532 = (inp[0]) ? node37606 : node37533;
											assign node37533 = (inp[15]) ? node37571 : node37534;
												assign node37534 = (inp[3]) ? node37554 : node37535;
													assign node37535 = (inp[4]) ? node37547 : node37536;
														assign node37536 = (inp[9]) ? node37542 : node37537;
															assign node37537 = (inp[12]) ? node37539 : 4'b0111;
																assign node37539 = (inp[10]) ? 4'b0011 : 4'b0111;
															assign node37542 = (inp[10]) ? node37544 : 4'b0011;
																assign node37544 = (inp[12]) ? 4'b0101 : 4'b0011;
														assign node37547 = (inp[9]) ? 4'b0101 : node37548;
															assign node37548 = (inp[10]) ? node37550 : 4'b0011;
																assign node37550 = (inp[12]) ? 4'b0101 : 4'b0011;
													assign node37554 = (inp[10]) ? node37564 : node37555;
														assign node37555 = (inp[12]) ? 4'b0101 : node37556;
															assign node37556 = (inp[4]) ? node37560 : node37557;
																assign node37557 = (inp[9]) ? 4'b0001 : 4'b0101;
																assign node37560 = (inp[9]) ? 4'b0101 : 4'b0001;
														assign node37564 = (inp[9]) ? 4'b0001 : node37565;
															assign node37565 = (inp[4]) ? 4'b0001 : node37566;
																assign node37566 = (inp[12]) ? 4'b0001 : 4'b0101;
												assign node37571 = (inp[3]) ? node37585 : node37572;
													assign node37572 = (inp[4]) ? node37576 : node37573;
														assign node37573 = (inp[9]) ? 4'b0001 : 4'b0101;
														assign node37576 = (inp[10]) ? node37580 : node37577;
															assign node37577 = (inp[9]) ? 4'b0111 : 4'b0001;
															assign node37580 = (inp[9]) ? node37582 : 4'b0111;
																assign node37582 = (inp[12]) ? 4'b0011 : 4'b0111;
													assign node37585 = (inp[10]) ? node37593 : node37586;
														assign node37586 = (inp[9]) ? node37590 : node37587;
															assign node37587 = (inp[4]) ? 4'b0011 : 4'b0111;
															assign node37590 = (inp[4]) ? 4'b0111 : 4'b0011;
														assign node37593 = (inp[12]) ? node37599 : node37594;
															assign node37594 = (inp[9]) ? node37596 : 4'b0011;
																assign node37596 = (inp[4]) ? 4'b0111 : 4'b0011;
															assign node37599 = (inp[9]) ? node37603 : node37600;
																assign node37600 = (inp[4]) ? 4'b0111 : 4'b0011;
																assign node37603 = (inp[4]) ? 4'b0011 : 4'b0111;
											assign node37606 = (inp[15]) ? node37646 : node37607;
												assign node37607 = (inp[3]) ? node37627 : node37608;
													assign node37608 = (inp[4]) ? node37616 : node37609;
														assign node37609 = (inp[9]) ? 4'b0001 : node37610;
															assign node37610 = (inp[10]) ? node37612 : 4'b0101;
																assign node37612 = (inp[12]) ? 4'b0001 : 4'b0101;
														assign node37616 = (inp[9]) ? node37622 : node37617;
															assign node37617 = (inp[12]) ? node37619 : 4'b0001;
																assign node37619 = (inp[10]) ? 4'b0111 : 4'b0001;
															assign node37622 = (inp[12]) ? node37624 : 4'b0111;
																assign node37624 = (inp[10]) ? 4'b0011 : 4'b0111;
													assign node37627 = (inp[12]) ? node37637 : node37628;
														assign node37628 = (inp[10]) ? node37630 : 4'b0111;
															assign node37630 = (inp[4]) ? node37634 : node37631;
																assign node37631 = (inp[9]) ? 4'b0011 : 4'b0111;
																assign node37634 = (inp[9]) ? 4'b0111 : 4'b0011;
														assign node37637 = (inp[10]) ? 4'b0111 : node37638;
															assign node37638 = (inp[9]) ? node37642 : node37639;
																assign node37639 = (inp[4]) ? 4'b0011 : 4'b0111;
																assign node37642 = (inp[4]) ? 4'b0111 : 4'b0011;
												assign node37646 = (inp[3]) ? node37668 : node37647;
													assign node37647 = (inp[9]) ? node37657 : node37648;
														assign node37648 = (inp[4]) ? node37652 : node37649;
															assign node37649 = (inp[10]) ? 4'b0011 : 4'b0111;
															assign node37652 = (inp[12]) ? node37654 : 4'b0011;
																assign node37654 = (inp[10]) ? 4'b0101 : 4'b0011;
														assign node37657 = (inp[4]) ? node37663 : node37658;
															assign node37658 = (inp[12]) ? node37660 : 4'b0011;
																assign node37660 = (inp[10]) ? 4'b0101 : 4'b0011;
															assign node37663 = (inp[10]) ? node37665 : 4'b0101;
																assign node37665 = (inp[12]) ? 4'b0001 : 4'b0101;
													assign node37668 = (inp[12]) ? node37674 : node37669;
														assign node37669 = (inp[9]) ? 4'b0001 : node37670;
															assign node37670 = (inp[4]) ? 4'b0001 : 4'b0101;
														assign node37674 = (inp[4]) ? node37682 : node37675;
															assign node37675 = (inp[10]) ? node37679 : node37676;
																assign node37676 = (inp[9]) ? 4'b0001 : 4'b0101;
																assign node37679 = (inp[9]) ? 4'b0101 : 4'b0001;
															assign node37682 = (inp[9]) ? 4'b0101 : node37683;
																assign node37683 = (inp[10]) ? 4'b0101 : 4'b0001;
									assign node37687 = (inp[3]) ? node37807 : node37688;
										assign node37688 = (inp[15]) ? node37752 : node37689;
											assign node37689 = (inp[0]) ? node37733 : node37690;
												assign node37690 = (inp[5]) ? node37712 : node37691;
													assign node37691 = (inp[10]) ? node37697 : node37692;
														assign node37692 = (inp[4]) ? 4'b0010 : node37693;
															assign node37693 = (inp[9]) ? 4'b0010 : 4'b0110;
														assign node37697 = (inp[4]) ? node37705 : node37698;
															assign node37698 = (inp[9]) ? node37702 : node37699;
																assign node37699 = (inp[12]) ? 4'b0010 : 4'b0110;
																assign node37702 = (inp[12]) ? 4'b0110 : 4'b0010;
															assign node37705 = (inp[12]) ? node37709 : node37706;
																assign node37706 = (inp[9]) ? 4'b0110 : 4'b0010;
																assign node37709 = (inp[9]) ? 4'b0010 : 4'b0110;
													assign node37712 = (inp[9]) ? node37722 : node37713;
														assign node37713 = (inp[10]) ? node37715 : 4'b0010;
															assign node37715 = (inp[12]) ? node37719 : node37716;
																assign node37716 = (inp[4]) ? 4'b0010 : 4'b0110;
																assign node37719 = (inp[4]) ? 4'b0100 : 4'b0010;
														assign node37722 = (inp[4]) ? node37728 : node37723;
															assign node37723 = (inp[10]) ? node37725 : 4'b0010;
																assign node37725 = (inp[12]) ? 4'b0100 : 4'b0010;
															assign node37728 = (inp[12]) ? node37730 : 4'b0100;
																assign node37730 = (inp[10]) ? 4'b0000 : 4'b0100;
												assign node37733 = (inp[5]) ? node37747 : node37734;
													assign node37734 = (inp[4]) ? node37742 : node37735;
														assign node37735 = (inp[9]) ? node37737 : 4'b0100;
															assign node37737 = (inp[12]) ? node37739 : 4'b0000;
																assign node37739 = (inp[10]) ? 4'b0100 : 4'b0000;
														assign node37742 = (inp[9]) ? node37744 : 4'b0000;
															assign node37744 = (inp[10]) ? 4'b0000 : 4'b0100;
													assign node37747 = (inp[9]) ? node37749 : 4'b0000;
														assign node37749 = (inp[10]) ? 4'b0110 : 4'b0000;
											assign node37752 = (inp[0]) ? node37780 : node37753;
												assign node37753 = (inp[10]) ? node37769 : node37754;
													assign node37754 = (inp[5]) ? node37762 : node37755;
														assign node37755 = (inp[9]) ? node37759 : node37756;
															assign node37756 = (inp[4]) ? 4'b0000 : 4'b0100;
															assign node37759 = (inp[4]) ? 4'b0100 : 4'b0000;
														assign node37762 = (inp[9]) ? node37766 : node37763;
															assign node37763 = (inp[4]) ? 4'b0000 : 4'b0100;
															assign node37766 = (inp[4]) ? 4'b0110 : 4'b0000;
													assign node37769 = (inp[4]) ? node37775 : node37770;
														assign node37770 = (inp[12]) ? 4'b0000 : node37771;
															assign node37771 = (inp[9]) ? 4'b0000 : 4'b0100;
														assign node37775 = (inp[5]) ? node37777 : 4'b0000;
															assign node37777 = (inp[12]) ? 4'b0010 : 4'b0000;
												assign node37780 = (inp[5]) ? node37792 : node37781;
													assign node37781 = (inp[4]) ? 4'b0010 : node37782;
														assign node37782 = (inp[10]) ? node37786 : node37783;
															assign node37783 = (inp[9]) ? 4'b0010 : 4'b0110;
															assign node37786 = (inp[9]) ? 4'b0110 : node37787;
																assign node37787 = (inp[12]) ? 4'b0010 : 4'b0110;
													assign node37792 = (inp[12]) ? node37800 : node37793;
														assign node37793 = (inp[4]) ? node37797 : node37794;
															assign node37794 = (inp[9]) ? 4'b0010 : 4'b0110;
															assign node37797 = (inp[9]) ? 4'b0100 : 4'b0010;
														assign node37800 = (inp[9]) ? node37802 : 4'b0100;
															assign node37802 = (inp[4]) ? node37804 : 4'b0100;
																assign node37804 = (inp[10]) ? 4'b0000 : 4'b0100;
										assign node37807 = (inp[9]) ? node37871 : node37808;
											assign node37808 = (inp[4]) ? node37842 : node37809;
												assign node37809 = (inp[12]) ? node37825 : node37810;
													assign node37810 = (inp[15]) ? node37818 : node37811;
														assign node37811 = (inp[5]) ? node37815 : node37812;
															assign node37812 = (inp[0]) ? 4'b0100 : 4'b0110;
															assign node37815 = (inp[0]) ? 4'b0110 : 4'b0100;
														assign node37818 = (inp[5]) ? node37822 : node37819;
															assign node37819 = (inp[0]) ? 4'b0110 : 4'b0100;
															assign node37822 = (inp[0]) ? 4'b0100 : 4'b0110;
													assign node37825 = (inp[10]) ? node37835 : node37826;
														assign node37826 = (inp[5]) ? 4'b0110 : node37827;
															assign node37827 = (inp[0]) ? node37831 : node37828;
																assign node37828 = (inp[15]) ? 4'b0100 : 4'b0110;
																assign node37831 = (inp[15]) ? 4'b0110 : 4'b0100;
														assign node37835 = (inp[15]) ? node37837 : 4'b0010;
															assign node37837 = (inp[0]) ? 4'b0000 : node37838;
																assign node37838 = (inp[5]) ? 4'b0010 : 4'b0000;
												assign node37842 = (inp[12]) ? node37856 : node37843;
													assign node37843 = (inp[0]) ? node37849 : node37844;
														assign node37844 = (inp[10]) ? node37846 : 4'b0000;
															assign node37846 = (inp[5]) ? 4'b0000 : 4'b0010;
														assign node37849 = (inp[15]) ? node37853 : node37850;
															assign node37850 = (inp[5]) ? 4'b0010 : 4'b0000;
															assign node37853 = (inp[5]) ? 4'b0000 : 4'b0010;
													assign node37856 = (inp[10]) ? node37864 : node37857;
														assign node37857 = (inp[15]) ? 4'b0000 : node37858;
															assign node37858 = (inp[5]) ? 4'b0000 : node37859;
																assign node37859 = (inp[0]) ? 4'b0000 : 4'b0010;
														assign node37864 = (inp[15]) ? node37868 : node37865;
															assign node37865 = (inp[0]) ? 4'b0110 : 4'b0100;
															assign node37868 = (inp[0]) ? 4'b0100 : 4'b0110;
											assign node37871 = (inp[4]) ? node37917 : node37872;
												assign node37872 = (inp[12]) ? node37900 : node37873;
													assign node37873 = (inp[10]) ? node37887 : node37874;
														assign node37874 = (inp[15]) ? node37880 : node37875;
															assign node37875 = (inp[5]) ? 4'b0000 : node37876;
																assign node37876 = (inp[0]) ? 4'b0000 : 4'b0010;
															assign node37880 = (inp[0]) ? node37884 : node37881;
																assign node37881 = (inp[5]) ? 4'b0010 : 4'b0000;
																assign node37884 = (inp[5]) ? 4'b0000 : 4'b0010;
														assign node37887 = (inp[15]) ? node37895 : node37888;
															assign node37888 = (inp[5]) ? node37892 : node37889;
																assign node37889 = (inp[0]) ? 4'b0000 : 4'b0010;
																assign node37892 = (inp[0]) ? 4'b0010 : 4'b0000;
															assign node37895 = (inp[0]) ? 4'b0010 : node37896;
																assign node37896 = (inp[5]) ? 4'b0010 : 4'b0000;
													assign node37900 = (inp[10]) ? node37910 : node37901;
														assign node37901 = (inp[15]) ? node37903 : 4'b0000;
															assign node37903 = (inp[0]) ? node37907 : node37904;
																assign node37904 = (inp[5]) ? 4'b0010 : 4'b0000;
																assign node37907 = (inp[5]) ? 4'b0000 : 4'b0010;
														assign node37910 = (inp[0]) ? node37914 : node37911;
															assign node37911 = (inp[15]) ? 4'b0110 : 4'b0100;
															assign node37914 = (inp[15]) ? 4'b0100 : 4'b0110;
												assign node37917 = (inp[12]) ? node37925 : node37918;
													assign node37918 = (inp[15]) ? node37922 : node37919;
														assign node37919 = (inp[0]) ? 4'b0110 : 4'b0100;
														assign node37922 = (inp[0]) ? 4'b0100 : 4'b0110;
													assign node37925 = (inp[10]) ? node37935 : node37926;
														assign node37926 = (inp[5]) ? node37928 : 4'b0110;
															assign node37928 = (inp[15]) ? node37932 : node37929;
																assign node37929 = (inp[0]) ? 4'b0110 : 4'b0100;
																assign node37932 = (inp[0]) ? 4'b0100 : 4'b0110;
														assign node37935 = (inp[5]) ? node37943 : node37936;
															assign node37936 = (inp[15]) ? node37940 : node37937;
																assign node37937 = (inp[0]) ? 4'b0010 : 4'b0000;
																assign node37940 = (inp[0]) ? 4'b0000 : 4'b0010;
															assign node37943 = (inp[0]) ? 4'b0010 : node37944;
																assign node37944 = (inp[15]) ? 4'b0010 : 4'b0000;
								assign node37948 = (inp[5]) ? node38176 : node37949;
									assign node37949 = (inp[9]) ? node38037 : node37950;
										assign node37950 = (inp[4]) ? node37982 : node37951;
											assign node37951 = (inp[12]) ? node37959 : node37952;
												assign node37952 = (inp[0]) ? node37956 : node37953;
													assign node37953 = (inp[15]) ? 4'b0100 : 4'b0110;
													assign node37956 = (inp[15]) ? 4'b0110 : 4'b0100;
												assign node37959 = (inp[10]) ? node37967 : node37960;
													assign node37960 = (inp[0]) ? node37964 : node37961;
														assign node37961 = (inp[15]) ? 4'b0100 : 4'b0110;
														assign node37964 = (inp[15]) ? 4'b0110 : 4'b0100;
													assign node37967 = (inp[3]) ? node37975 : node37968;
														assign node37968 = (inp[2]) ? 4'b0000 : node37969;
															assign node37969 = (inp[15]) ? node37971 : 4'b0000;
																assign node37971 = (inp[0]) ? 4'b0010 : 4'b0000;
														assign node37975 = (inp[15]) ? node37979 : node37976;
															assign node37976 = (inp[0]) ? 4'b0000 : 4'b0010;
															assign node37979 = (inp[0]) ? 4'b0010 : 4'b0000;
											assign node37982 = (inp[12]) ? node38006 : node37983;
												assign node37983 = (inp[10]) ? node37991 : node37984;
													assign node37984 = (inp[0]) ? node37988 : node37985;
														assign node37985 = (inp[15]) ? 4'b0000 : 4'b0010;
														assign node37988 = (inp[15]) ? 4'b0010 : 4'b0000;
													assign node37991 = (inp[3]) ? node37999 : node37992;
														assign node37992 = (inp[0]) ? node37996 : node37993;
															assign node37993 = (inp[15]) ? 4'b0000 : 4'b0010;
															assign node37996 = (inp[15]) ? 4'b0010 : 4'b0000;
														assign node37999 = (inp[15]) ? node38003 : node38000;
															assign node38000 = (inp[0]) ? 4'b0000 : 4'b0010;
															assign node38003 = (inp[0]) ? 4'b0010 : 4'b0000;
												assign node38006 = (inp[10]) ? node38022 : node38007;
													assign node38007 = (inp[3]) ? node38013 : node38008;
														assign node38008 = (inp[15]) ? node38010 : 4'b0000;
															assign node38010 = (inp[0]) ? 4'b0010 : 4'b0000;
														assign node38013 = (inp[2]) ? node38019 : node38014;
															assign node38014 = (inp[15]) ? node38016 : 4'b0000;
																assign node38016 = (inp[0]) ? 4'b0010 : 4'b0000;
															assign node38019 = (inp[15]) ? 4'b0000 : 4'b0010;
													assign node38022 = (inp[15]) ? node38030 : node38023;
														assign node38023 = (inp[0]) ? node38027 : node38024;
															assign node38024 = (inp[3]) ? 4'b0100 : 4'b0110;
															assign node38027 = (inp[3]) ? 4'b0110 : 4'b0100;
														assign node38030 = (inp[0]) ? node38034 : node38031;
															assign node38031 = (inp[2]) ? 4'b0100 : 4'b0110;
															assign node38034 = (inp[3]) ? 4'b0100 : 4'b0110;
										assign node38037 = (inp[4]) ? node38093 : node38038;
											assign node38038 = (inp[10]) ? node38068 : node38039;
												assign node38039 = (inp[3]) ? node38053 : node38040;
													assign node38040 = (inp[12]) ? node38046 : node38041;
														assign node38041 = (inp[15]) ? 4'b0000 : node38042;
															assign node38042 = (inp[0]) ? 4'b0000 : 4'b0010;
														assign node38046 = (inp[15]) ? node38050 : node38047;
															assign node38047 = (inp[0]) ? 4'b0000 : 4'b0010;
															assign node38050 = (inp[0]) ? 4'b0010 : 4'b0000;
													assign node38053 = (inp[2]) ? node38061 : node38054;
														assign node38054 = (inp[0]) ? node38058 : node38055;
															assign node38055 = (inp[12]) ? 4'b0000 : 4'b0010;
															assign node38058 = (inp[15]) ? 4'b0010 : 4'b0000;
														assign node38061 = (inp[0]) ? node38065 : node38062;
															assign node38062 = (inp[15]) ? 4'b0000 : 4'b0010;
															assign node38065 = (inp[15]) ? 4'b0010 : 4'b0000;
												assign node38068 = (inp[12]) ? node38078 : node38069;
													assign node38069 = (inp[2]) ? node38075 : node38070;
														assign node38070 = (inp[15]) ? node38072 : 4'b0000;
															assign node38072 = (inp[0]) ? 4'b0010 : 4'b0000;
														assign node38075 = (inp[3]) ? 4'b0000 : 4'b0010;
													assign node38078 = (inp[15]) ? node38086 : node38079;
														assign node38079 = (inp[3]) ? node38083 : node38080;
															assign node38080 = (inp[0]) ? 4'b0100 : 4'b0110;
															assign node38083 = (inp[0]) ? 4'b0110 : 4'b0100;
														assign node38086 = (inp[0]) ? node38090 : node38087;
															assign node38087 = (inp[3]) ? 4'b0110 : 4'b0100;
															assign node38090 = (inp[3]) ? 4'b0100 : 4'b0110;
											assign node38093 = (inp[10]) ? node38143 : node38094;
												assign node38094 = (inp[15]) ? node38114 : node38095;
													assign node38095 = (inp[12]) ? node38107 : node38096;
														assign node38096 = (inp[2]) ? node38102 : node38097;
															assign node38097 = (inp[3]) ? 4'b0110 : node38098;
																assign node38098 = (inp[0]) ? 4'b0100 : 4'b0110;
															assign node38102 = (inp[0]) ? 4'b0110 : node38103;
																assign node38103 = (inp[3]) ? 4'b0100 : 4'b0110;
														assign node38107 = (inp[3]) ? node38111 : node38108;
															assign node38108 = (inp[0]) ? 4'b0100 : 4'b0110;
															assign node38111 = (inp[0]) ? 4'b0110 : 4'b0100;
													assign node38114 = (inp[12]) ? node38130 : node38115;
														assign node38115 = (inp[2]) ? node38123 : node38116;
															assign node38116 = (inp[0]) ? node38120 : node38117;
																assign node38117 = (inp[3]) ? 4'b0110 : 4'b0100;
																assign node38120 = (inp[3]) ? 4'b0100 : 4'b0110;
															assign node38123 = (inp[3]) ? node38127 : node38124;
																assign node38124 = (inp[0]) ? 4'b0110 : 4'b0100;
																assign node38127 = (inp[0]) ? 4'b0100 : 4'b0110;
														assign node38130 = (inp[2]) ? node38136 : node38131;
															assign node38131 = (inp[0]) ? node38133 : 4'b0100;
																assign node38133 = (inp[3]) ? 4'b0100 : 4'b0110;
															assign node38136 = (inp[3]) ? node38140 : node38137;
																assign node38137 = (inp[0]) ? 4'b0110 : 4'b0100;
																assign node38140 = (inp[0]) ? 4'b0100 : 4'b0110;
												assign node38143 = (inp[12]) ? node38159 : node38144;
													assign node38144 = (inp[3]) ? node38152 : node38145;
														assign node38145 = (inp[0]) ? node38149 : node38146;
															assign node38146 = (inp[15]) ? 4'b0100 : 4'b0110;
															assign node38149 = (inp[15]) ? 4'b0110 : 4'b0100;
														assign node38152 = (inp[0]) ? node38156 : node38153;
															assign node38153 = (inp[15]) ? 4'b0110 : 4'b0100;
															assign node38156 = (inp[15]) ? 4'b0100 : 4'b0110;
													assign node38159 = (inp[2]) ? node38169 : node38160;
														assign node38160 = (inp[0]) ? node38162 : 4'b0010;
															assign node38162 = (inp[15]) ? node38166 : node38163;
																assign node38163 = (inp[3]) ? 4'b0010 : 4'b0000;
																assign node38166 = (inp[3]) ? 4'b0000 : 4'b0010;
														assign node38169 = (inp[3]) ? node38171 : 4'b0000;
															assign node38171 = (inp[0]) ? node38173 : 4'b0000;
																assign node38173 = (inp[15]) ? 4'b0000 : 4'b0010;
									assign node38176 = (inp[3]) ? node38260 : node38177;
										assign node38177 = (inp[15]) ? node38217 : node38178;
											assign node38178 = (inp[0]) ? node38198 : node38179;
												assign node38179 = (inp[4]) ? node38191 : node38180;
													assign node38180 = (inp[9]) ? node38186 : node38181;
														assign node38181 = (inp[10]) ? node38183 : 4'b0110;
															assign node38183 = (inp[12]) ? 4'b0010 : 4'b0110;
														assign node38186 = (inp[10]) ? node38188 : 4'b0010;
															assign node38188 = (inp[12]) ? 4'b0100 : 4'b0010;
													assign node38191 = (inp[9]) ? 4'b0100 : node38192;
														assign node38192 = (inp[10]) ? node38194 : 4'b0010;
															assign node38194 = (inp[12]) ? 4'b0100 : 4'b0010;
												assign node38198 = (inp[4]) ? node38206 : node38199;
													assign node38199 = (inp[9]) ? 4'b0000 : node38200;
														assign node38200 = (inp[12]) ? node38202 : 4'b0100;
															assign node38202 = (inp[10]) ? 4'b0000 : 4'b0100;
													assign node38206 = (inp[9]) ? node38212 : node38207;
														assign node38207 = (inp[10]) ? node38209 : 4'b0000;
															assign node38209 = (inp[12]) ? 4'b0110 : 4'b0000;
														assign node38212 = (inp[10]) ? node38214 : 4'b0110;
															assign node38214 = (inp[2]) ? 4'b0110 : 4'b0010;
											assign node38217 = (inp[0]) ? node38237 : node38218;
												assign node38218 = (inp[9]) ? node38226 : node38219;
													assign node38219 = (inp[4]) ? 4'b0000 : node38220;
														assign node38220 = (inp[10]) ? node38222 : 4'b0100;
															assign node38222 = (inp[12]) ? 4'b0000 : 4'b0100;
													assign node38226 = (inp[4]) ? node38232 : node38227;
														assign node38227 = (inp[12]) ? node38229 : 4'b0000;
															assign node38229 = (inp[10]) ? 4'b0110 : 4'b0000;
														assign node38232 = (inp[12]) ? node38234 : 4'b0110;
															assign node38234 = (inp[10]) ? 4'b0010 : 4'b0110;
												assign node38237 = (inp[10]) ? node38247 : node38238;
													assign node38238 = (inp[12]) ? node38240 : 4'b0010;
														assign node38240 = (inp[4]) ? node38244 : node38241;
															assign node38241 = (inp[9]) ? 4'b0010 : 4'b0110;
															assign node38244 = (inp[9]) ? 4'b0100 : 4'b0010;
													assign node38247 = (inp[9]) ? node38253 : node38248;
														assign node38248 = (inp[12]) ? node38250 : 4'b0010;
															assign node38250 = (inp[4]) ? 4'b0100 : 4'b0010;
														assign node38253 = (inp[12]) ? node38257 : node38254;
															assign node38254 = (inp[4]) ? 4'b0100 : 4'b0010;
															assign node38257 = (inp[4]) ? 4'b0000 : 4'b0100;
										assign node38260 = (inp[0]) ? node38330 : node38261;
											assign node38261 = (inp[15]) ? node38287 : node38262;
												assign node38262 = (inp[12]) ? node38278 : node38263;
													assign node38263 = (inp[2]) ? node38271 : node38264;
														assign node38264 = (inp[9]) ? node38268 : node38265;
															assign node38265 = (inp[4]) ? 4'b0000 : 4'b0100;
															assign node38268 = (inp[10]) ? 4'b0100 : 4'b0000;
														assign node38271 = (inp[9]) ? node38275 : node38272;
															assign node38272 = (inp[4]) ? 4'b0000 : 4'b0100;
															assign node38275 = (inp[4]) ? 4'b0100 : 4'b0000;
													assign node38278 = (inp[10]) ? 4'b0000 : node38279;
														assign node38279 = (inp[4]) ? node38283 : node38280;
															assign node38280 = (inp[9]) ? 4'b0000 : 4'b0100;
															assign node38283 = (inp[9]) ? 4'b0100 : 4'b0000;
												assign node38287 = (inp[2]) ? node38309 : node38288;
													assign node38288 = (inp[9]) ? node38300 : node38289;
														assign node38289 = (inp[4]) ? node38295 : node38290;
															assign node38290 = (inp[10]) ? node38292 : 4'b0110;
																assign node38292 = (inp[12]) ? 4'b0010 : 4'b0110;
															assign node38295 = (inp[10]) ? node38297 : 4'b0010;
																assign node38297 = (inp[12]) ? 4'b0110 : 4'b0010;
														assign node38300 = (inp[10]) ? node38302 : 4'b0010;
															assign node38302 = (inp[12]) ? node38306 : node38303;
																assign node38303 = (inp[4]) ? 4'b0110 : 4'b0010;
																assign node38306 = (inp[4]) ? 4'b0010 : 4'b0110;
													assign node38309 = (inp[4]) ? node38321 : node38310;
														assign node38310 = (inp[9]) ? node38316 : node38311;
															assign node38311 = (inp[12]) ? node38313 : 4'b0110;
																assign node38313 = (inp[10]) ? 4'b0010 : 4'b0110;
															assign node38316 = (inp[10]) ? node38318 : 4'b0010;
																assign node38318 = (inp[12]) ? 4'b0110 : 4'b0010;
														assign node38321 = (inp[9]) ? node38325 : node38322;
															assign node38322 = (inp[10]) ? 4'b0110 : 4'b0010;
															assign node38325 = (inp[10]) ? node38327 : 4'b0110;
																assign node38327 = (inp[12]) ? 4'b0010 : 4'b0110;
											assign node38330 = (inp[15]) ? node38360 : node38331;
												assign node38331 = (inp[2]) ? node38343 : node38332;
													assign node38332 = (inp[4]) ? 4'b0010 : node38333;
														assign node38333 = (inp[9]) ? node38339 : node38334;
															assign node38334 = (inp[12]) ? node38336 : 4'b0110;
																assign node38336 = (inp[10]) ? 4'b0010 : 4'b0110;
															assign node38339 = (inp[10]) ? 4'b0110 : 4'b0010;
													assign node38343 = (inp[12]) ? node38351 : node38344;
														assign node38344 = (inp[4]) ? node38348 : node38345;
															assign node38345 = (inp[9]) ? 4'b0010 : 4'b0110;
															assign node38348 = (inp[9]) ? 4'b0110 : 4'b0010;
														assign node38351 = (inp[9]) ? 4'b0110 : node38352;
															assign node38352 = (inp[4]) ? node38356 : node38353;
																assign node38353 = (inp[10]) ? 4'b0010 : 4'b0110;
																assign node38356 = (inp[10]) ? 4'b0110 : 4'b0010;
												assign node38360 = (inp[4]) ? node38368 : node38361;
													assign node38361 = (inp[9]) ? 4'b0000 : node38362;
														assign node38362 = (inp[12]) ? node38364 : 4'b0100;
															assign node38364 = (inp[10]) ? 4'b0000 : 4'b0100;
													assign node38368 = (inp[9]) ? node38372 : node38369;
														assign node38369 = (inp[12]) ? 4'b0100 : 4'b0000;
														assign node38372 = (inp[10]) ? node38374 : 4'b0100;
															assign node38374 = (inp[12]) ? 4'b0000 : 4'b0100;
							assign node38377 = (inp[2]) ? node38915 : node38378;
								assign node38378 = (inp[14]) ? node38644 : node38379;
									assign node38379 = (inp[12]) ? node38485 : node38380;
										assign node38380 = (inp[4]) ? node38428 : node38381;
											assign node38381 = (inp[9]) ? node38407 : node38382;
												assign node38382 = (inp[3]) ? node38392 : node38383;
													assign node38383 = (inp[10]) ? 4'b0100 : node38384;
														assign node38384 = (inp[15]) ? node38388 : node38385;
															assign node38385 = (inp[0]) ? 4'b0100 : 4'b0110;
															assign node38388 = (inp[0]) ? 4'b0110 : 4'b0100;
													assign node38392 = (inp[0]) ? node38400 : node38393;
														assign node38393 = (inp[5]) ? node38397 : node38394;
															assign node38394 = (inp[15]) ? 4'b0100 : 4'b0110;
															assign node38397 = (inp[15]) ? 4'b0110 : 4'b0100;
														assign node38400 = (inp[5]) ? node38404 : node38401;
															assign node38401 = (inp[15]) ? 4'b0110 : 4'b0100;
															assign node38404 = (inp[15]) ? 4'b0100 : 4'b0110;
												assign node38407 = (inp[0]) ? node38417 : node38408;
													assign node38408 = (inp[15]) ? node38412 : node38409;
														assign node38409 = (inp[5]) ? 4'b0000 : 4'b0010;
														assign node38412 = (inp[5]) ? node38414 : 4'b0000;
															assign node38414 = (inp[3]) ? 4'b0010 : 4'b0000;
													assign node38417 = (inp[15]) ? node38423 : node38418;
														assign node38418 = (inp[5]) ? node38420 : 4'b0000;
															assign node38420 = (inp[3]) ? 4'b0010 : 4'b0000;
														assign node38423 = (inp[3]) ? node38425 : 4'b0010;
															assign node38425 = (inp[5]) ? 4'b0000 : 4'b0010;
											assign node38428 = (inp[9]) ? node38466 : node38429;
												assign node38429 = (inp[5]) ? node38445 : node38430;
													assign node38430 = (inp[10]) ? node38438 : node38431;
														assign node38431 = (inp[15]) ? node38435 : node38432;
															assign node38432 = (inp[0]) ? 4'b0000 : 4'b0010;
															assign node38435 = (inp[0]) ? 4'b0010 : 4'b0000;
														assign node38438 = (inp[15]) ? node38442 : node38439;
															assign node38439 = (inp[0]) ? 4'b0000 : 4'b0010;
															assign node38442 = (inp[0]) ? 4'b0010 : 4'b0000;
													assign node38445 = (inp[3]) ? node38461 : node38446;
														assign node38446 = (inp[10]) ? node38454 : node38447;
															assign node38447 = (inp[15]) ? node38451 : node38448;
																assign node38448 = (inp[0]) ? 4'b0000 : 4'b0010;
																assign node38451 = (inp[0]) ? 4'b0010 : 4'b0000;
															assign node38454 = (inp[15]) ? node38458 : node38455;
																assign node38455 = (inp[0]) ? 4'b0000 : 4'b0010;
																assign node38458 = (inp[0]) ? 4'b0010 : 4'b0000;
														assign node38461 = (inp[15]) ? node38463 : 4'b0000;
															assign node38463 = (inp[0]) ? 4'b0000 : 4'b0010;
												assign node38466 = (inp[0]) ? node38474 : node38467;
													assign node38467 = (inp[15]) ? 4'b0110 : node38468;
														assign node38468 = (inp[5]) ? 4'b0100 : node38469;
															assign node38469 = (inp[3]) ? 4'b0100 : 4'b0110;
													assign node38474 = (inp[15]) ? node38480 : node38475;
														assign node38475 = (inp[3]) ? 4'b0110 : node38476;
															assign node38476 = (inp[5]) ? 4'b0110 : 4'b0100;
														assign node38480 = (inp[3]) ? 4'b0100 : node38481;
															assign node38481 = (inp[5]) ? 4'b0100 : 4'b0110;
										assign node38485 = (inp[10]) ? node38563 : node38486;
											assign node38486 = (inp[3]) ? node38524 : node38487;
												assign node38487 = (inp[15]) ? node38507 : node38488;
													assign node38488 = (inp[0]) ? node38498 : node38489;
														assign node38489 = (inp[4]) ? node38493 : node38490;
															assign node38490 = (inp[9]) ? 4'b0010 : 4'b0110;
															assign node38493 = (inp[9]) ? node38495 : 4'b0010;
																assign node38495 = (inp[5]) ? 4'b0100 : 4'b0110;
														assign node38498 = (inp[9]) ? node38502 : node38499;
															assign node38499 = (inp[4]) ? 4'b0000 : 4'b0100;
															assign node38502 = (inp[4]) ? node38504 : 4'b0000;
																assign node38504 = (inp[5]) ? 4'b0110 : 4'b0100;
													assign node38507 = (inp[0]) ? node38515 : node38508;
														assign node38508 = (inp[9]) ? node38512 : node38509;
															assign node38509 = (inp[4]) ? 4'b0000 : 4'b0100;
															assign node38512 = (inp[4]) ? 4'b0110 : 4'b0000;
														assign node38515 = (inp[9]) ? node38519 : node38516;
															assign node38516 = (inp[4]) ? 4'b0010 : 4'b0110;
															assign node38519 = (inp[4]) ? node38521 : 4'b0010;
																assign node38521 = (inp[5]) ? 4'b0100 : 4'b0110;
												assign node38524 = (inp[15]) ? node38544 : node38525;
													assign node38525 = (inp[9]) ? node38537 : node38526;
														assign node38526 = (inp[4]) ? node38530 : node38527;
															assign node38527 = (inp[0]) ? 4'b0100 : 4'b0110;
															assign node38530 = (inp[0]) ? node38534 : node38531;
																assign node38531 = (inp[5]) ? 4'b0000 : 4'b0010;
																assign node38534 = (inp[5]) ? 4'b0010 : 4'b0000;
														assign node38537 = (inp[4]) ? node38541 : node38538;
															assign node38538 = (inp[5]) ? 4'b0010 : 4'b0000;
															assign node38541 = (inp[0]) ? 4'b0110 : 4'b0100;
													assign node38544 = (inp[0]) ? node38556 : node38545;
														assign node38545 = (inp[5]) ? node38553 : node38546;
															assign node38546 = (inp[9]) ? node38550 : node38547;
																assign node38547 = (inp[4]) ? 4'b0000 : 4'b0100;
																assign node38550 = (inp[4]) ? 4'b0110 : 4'b0000;
															assign node38553 = (inp[4]) ? 4'b0010 : 4'b0110;
														assign node38556 = (inp[4]) ? 4'b0100 : node38557;
															assign node38557 = (inp[5]) ? 4'b0100 : node38558;
																assign node38558 = (inp[9]) ? 4'b0010 : 4'b0110;
											assign node38563 = (inp[4]) ? node38599 : node38564;
												assign node38564 = (inp[9]) ? node38586 : node38565;
													assign node38565 = (inp[5]) ? node38571 : node38566;
														assign node38566 = (inp[15]) ? node38568 : 4'b0010;
															assign node38568 = (inp[0]) ? 4'b0010 : 4'b0000;
														assign node38571 = (inp[15]) ? node38579 : node38572;
															assign node38572 = (inp[0]) ? node38576 : node38573;
																assign node38573 = (inp[3]) ? 4'b0000 : 4'b0010;
																assign node38576 = (inp[3]) ? 4'b0010 : 4'b0000;
															assign node38579 = (inp[0]) ? node38583 : node38580;
																assign node38580 = (inp[3]) ? 4'b0010 : 4'b0000;
																assign node38583 = (inp[3]) ? 4'b0000 : 4'b0010;
													assign node38586 = (inp[5]) ? node38592 : node38587;
														assign node38587 = (inp[3]) ? 4'b0110 : node38588;
															assign node38588 = (inp[15]) ? 4'b0110 : 4'b0100;
														assign node38592 = (inp[15]) ? node38596 : node38593;
															assign node38593 = (inp[0]) ? 4'b0110 : 4'b0100;
															assign node38596 = (inp[0]) ? 4'b0100 : 4'b0110;
												assign node38599 = (inp[9]) ? node38629 : node38600;
													assign node38600 = (inp[3]) ? node38614 : node38601;
														assign node38601 = (inp[15]) ? node38609 : node38602;
															assign node38602 = (inp[0]) ? node38606 : node38603;
																assign node38603 = (inp[5]) ? 4'b0100 : 4'b0110;
																assign node38606 = (inp[5]) ? 4'b0110 : 4'b0100;
															assign node38609 = (inp[5]) ? 4'b0110 : node38610;
																assign node38610 = (inp[0]) ? 4'b0110 : 4'b0100;
														assign node38614 = (inp[5]) ? node38622 : node38615;
															assign node38615 = (inp[0]) ? node38619 : node38616;
																assign node38616 = (inp[15]) ? 4'b0110 : 4'b0100;
																assign node38619 = (inp[15]) ? 4'b0100 : 4'b0110;
															assign node38622 = (inp[0]) ? node38626 : node38623;
																assign node38623 = (inp[15]) ? 4'b0110 : 4'b0100;
																assign node38626 = (inp[15]) ? 4'b0100 : 4'b0110;
													assign node38629 = (inp[15]) ? node38639 : node38630;
														assign node38630 = (inp[5]) ? node38636 : node38631;
															assign node38631 = (inp[3]) ? 4'b0000 : node38632;
																assign node38632 = (inp[0]) ? 4'b0000 : 4'b0010;
															assign node38636 = (inp[0]) ? 4'b0010 : 4'b0000;
														assign node38639 = (inp[0]) ? node38641 : 4'b0010;
															assign node38641 = (inp[5]) ? 4'b0000 : 4'b0010;
									assign node38644 = (inp[10]) ? node38802 : node38645;
										assign node38645 = (inp[3]) ? node38727 : node38646;
											assign node38646 = (inp[0]) ? node38696 : node38647;
												assign node38647 = (inp[15]) ? node38669 : node38648;
													assign node38648 = (inp[5]) ? node38660 : node38649;
														assign node38649 = (inp[4]) ? node38655 : node38650;
															assign node38650 = (inp[9]) ? node38652 : 4'b1011;
																assign node38652 = (inp[12]) ? 4'b1111 : 4'b1011;
															assign node38655 = (inp[12]) ? node38657 : 4'b1111;
																assign node38657 = (inp[9]) ? 4'b1011 : 4'b1111;
														assign node38660 = (inp[12]) ? 4'b1101 : node38661;
															assign node38661 = (inp[9]) ? node38665 : node38662;
																assign node38662 = (inp[4]) ? 4'b1011 : 4'b1111;
																assign node38665 = (inp[4]) ? 4'b1101 : 4'b1011;
													assign node38669 = (inp[5]) ? node38683 : node38670;
														assign node38670 = (inp[9]) ? node38676 : node38671;
															assign node38671 = (inp[4]) ? 4'b1101 : node38672;
																assign node38672 = (inp[12]) ? 4'b1001 : 4'b1101;
															assign node38676 = (inp[12]) ? node38680 : node38677;
																assign node38677 = (inp[4]) ? 4'b1101 : 4'b1001;
																assign node38680 = (inp[4]) ? 4'b1001 : 4'b1101;
														assign node38683 = (inp[4]) ? node38691 : node38684;
															assign node38684 = (inp[12]) ? node38688 : node38685;
																assign node38685 = (inp[9]) ? 4'b1001 : 4'b1101;
																assign node38688 = (inp[9]) ? 4'b1111 : 4'b1001;
															assign node38691 = (inp[9]) ? node38693 : 4'b1111;
																assign node38693 = (inp[12]) ? 4'b1011 : 4'b1111;
												assign node38696 = (inp[15]) ? node38714 : node38697;
													assign node38697 = (inp[12]) ? node38703 : node38698;
														assign node38698 = (inp[5]) ? node38700 : 4'b1001;
															assign node38700 = (inp[4]) ? 4'b1001 : 4'b1101;
														assign node38703 = (inp[5]) ? node38709 : node38704;
															assign node38704 = (inp[9]) ? node38706 : 4'b1101;
																assign node38706 = (inp[4]) ? 4'b1001 : 4'b1101;
															assign node38709 = (inp[9]) ? node38711 : 4'b1111;
																assign node38711 = (inp[4]) ? 4'b1011 : 4'b1111;
													assign node38714 = (inp[4]) ? node38722 : node38715;
														assign node38715 = (inp[12]) ? node38719 : node38716;
															assign node38716 = (inp[9]) ? 4'b1011 : 4'b1111;
															assign node38719 = (inp[9]) ? 4'b1111 : 4'b1011;
														assign node38722 = (inp[5]) ? node38724 : 4'b1011;
															assign node38724 = (inp[12]) ? 4'b1001 : 4'b1101;
											assign node38727 = (inp[9]) ? node38771 : node38728;
												assign node38728 = (inp[15]) ? node38750 : node38729;
													assign node38729 = (inp[12]) ? node38739 : node38730;
														assign node38730 = (inp[4]) ? 4'b1011 : node38731;
															assign node38731 = (inp[0]) ? node38735 : node38732;
																assign node38732 = (inp[5]) ? 4'b1101 : 4'b1111;
																assign node38735 = (inp[5]) ? 4'b1111 : 4'b1101;
														assign node38739 = (inp[4]) ? node38747 : node38740;
															assign node38740 = (inp[5]) ? node38744 : node38741;
																assign node38741 = (inp[0]) ? 4'b1001 : 4'b1011;
																assign node38744 = (inp[0]) ? 4'b1011 : 4'b1001;
															assign node38747 = (inp[0]) ? 4'b1111 : 4'b1101;
													assign node38750 = (inp[0]) ? node38764 : node38751;
														assign node38751 = (inp[5]) ? node38759 : node38752;
															assign node38752 = (inp[4]) ? node38756 : node38753;
																assign node38753 = (inp[12]) ? 4'b1001 : 4'b1101;
																assign node38756 = (inp[12]) ? 4'b1111 : 4'b1001;
															assign node38759 = (inp[4]) ? node38761 : 4'b1011;
																assign node38761 = (inp[12]) ? 4'b1111 : 4'b1011;
														assign node38764 = (inp[12]) ? 4'b1101 : node38765;
															assign node38765 = (inp[5]) ? node38767 : 4'b1011;
																assign node38767 = (inp[4]) ? 4'b1001 : 4'b1101;
												assign node38771 = (inp[12]) ? node38787 : node38772;
													assign node38772 = (inp[4]) ? node38774 : 4'b1011;
														assign node38774 = (inp[5]) ? node38782 : node38775;
															assign node38775 = (inp[15]) ? node38779 : node38776;
																assign node38776 = (inp[0]) ? 4'b1111 : 4'b1101;
																assign node38779 = (inp[0]) ? 4'b1101 : 4'b1111;
															assign node38782 = (inp[15]) ? node38784 : 4'b1111;
																assign node38784 = (inp[0]) ? 4'b1101 : 4'b1111;
													assign node38787 = (inp[4]) ? node38797 : node38788;
														assign node38788 = (inp[5]) ? 4'b1101 : node38789;
															assign node38789 = (inp[15]) ? node38793 : node38790;
																assign node38790 = (inp[0]) ? 4'b1111 : 4'b1101;
																assign node38793 = (inp[0]) ? 4'b1101 : 4'b1111;
														assign node38797 = (inp[15]) ? node38799 : 4'b1001;
															assign node38799 = (inp[0]) ? 4'b1001 : 4'b1011;
										assign node38802 = (inp[0]) ? node38852 : node38803;
											assign node38803 = (inp[15]) ? node38823 : node38804;
												assign node38804 = (inp[3]) ? node38814 : node38805;
													assign node38805 = (inp[4]) ? node38809 : node38806;
														assign node38806 = (inp[9]) ? 4'b1111 : 4'b1011;
														assign node38809 = (inp[5]) ? node38811 : 4'b1011;
															assign node38811 = (inp[9]) ? 4'b1001 : 4'b1101;
													assign node38814 = (inp[4]) ? node38820 : node38815;
														assign node38815 = (inp[5]) ? node38817 : 4'b1011;
															assign node38817 = (inp[9]) ? 4'b1101 : 4'b1001;
														assign node38820 = (inp[9]) ? 4'b1001 : 4'b1101;
												assign node38823 = (inp[3]) ? node38837 : node38824;
													assign node38824 = (inp[5]) ? node38832 : node38825;
														assign node38825 = (inp[9]) ? node38829 : node38826;
															assign node38826 = (inp[4]) ? 4'b1101 : 4'b1001;
															assign node38829 = (inp[4]) ? 4'b1001 : 4'b1101;
														assign node38832 = (inp[12]) ? 4'b1001 : node38833;
															assign node38833 = (inp[9]) ? 4'b1011 : 4'b1111;
													assign node38837 = (inp[5]) ? node38845 : node38838;
														assign node38838 = (inp[9]) ? node38842 : node38839;
															assign node38839 = (inp[4]) ? 4'b1111 : 4'b1001;
															assign node38842 = (inp[4]) ? 4'b1011 : 4'b1111;
														assign node38845 = (inp[4]) ? node38849 : node38846;
															assign node38846 = (inp[9]) ? 4'b1111 : 4'b1011;
															assign node38849 = (inp[9]) ? 4'b1011 : 4'b1111;
											assign node38852 = (inp[15]) ? node38886 : node38853;
												assign node38853 = (inp[5]) ? node38869 : node38854;
													assign node38854 = (inp[3]) ? node38862 : node38855;
														assign node38855 = (inp[9]) ? node38859 : node38856;
															assign node38856 = (inp[4]) ? 4'b1101 : 4'b1001;
															assign node38859 = (inp[4]) ? 4'b1001 : 4'b1101;
														assign node38862 = (inp[9]) ? node38866 : node38863;
															assign node38863 = (inp[4]) ? 4'b1111 : 4'b1001;
															assign node38866 = (inp[4]) ? 4'b1011 : 4'b1111;
													assign node38869 = (inp[3]) ? node38877 : node38870;
														assign node38870 = (inp[4]) ? node38874 : node38871;
															assign node38871 = (inp[9]) ? 4'b1111 : 4'b1001;
															assign node38874 = (inp[9]) ? 4'b1011 : 4'b1111;
														assign node38877 = (inp[12]) ? 4'b1011 : node38878;
															assign node38878 = (inp[4]) ? node38882 : node38879;
																assign node38879 = (inp[9]) ? 4'b1111 : 4'b1011;
																assign node38882 = (inp[9]) ? 4'b1011 : 4'b1111;
												assign node38886 = (inp[3]) ? node38908 : node38887;
													assign node38887 = (inp[5]) ? node38901 : node38888;
														assign node38888 = (inp[12]) ? node38894 : node38889;
															assign node38889 = (inp[9]) ? node38891 : 4'b1111;
																assign node38891 = (inp[4]) ? 4'b1011 : 4'b1111;
															assign node38894 = (inp[9]) ? node38898 : node38895;
																assign node38895 = (inp[4]) ? 4'b1111 : 4'b1011;
																assign node38898 = (inp[4]) ? 4'b1011 : 4'b1111;
														assign node38901 = (inp[4]) ? node38905 : node38902;
															assign node38902 = (inp[9]) ? 4'b1101 : 4'b1011;
															assign node38905 = (inp[9]) ? 4'b1001 : 4'b1101;
													assign node38908 = (inp[9]) ? node38912 : node38909;
														assign node38909 = (inp[4]) ? 4'b1101 : 4'b1001;
														assign node38912 = (inp[4]) ? 4'b1001 : 4'b1101;
								assign node38915 = (inp[10]) ? node39191 : node38916;
									assign node38916 = (inp[5]) ? node39054 : node38917;
										assign node38917 = (inp[4]) ? node38975 : node38918;
											assign node38918 = (inp[15]) ? node38946 : node38919;
												assign node38919 = (inp[0]) ? node38931 : node38920;
													assign node38920 = (inp[3]) ? node38926 : node38921;
														assign node38921 = (inp[9]) ? 4'b1111 : node38922;
															assign node38922 = (inp[12]) ? 4'b1011 : 4'b1111;
														assign node38926 = (inp[12]) ? node38928 : 4'b1011;
															assign node38928 = (inp[9]) ? 4'b1101 : 4'b1011;
													assign node38931 = (inp[3]) ? node38939 : node38932;
														assign node38932 = (inp[9]) ? node38936 : node38933;
															assign node38933 = (inp[12]) ? 4'b1001 : 4'b1101;
															assign node38936 = (inp[12]) ? 4'b1101 : 4'b1001;
														assign node38939 = (inp[12]) ? node38943 : node38940;
															assign node38940 = (inp[9]) ? 4'b1001 : 4'b1101;
															assign node38943 = (inp[9]) ? 4'b1111 : 4'b1001;
												assign node38946 = (inp[0]) ? node38962 : node38947;
													assign node38947 = (inp[3]) ? node38955 : node38948;
														assign node38948 = (inp[9]) ? node38952 : node38949;
															assign node38949 = (inp[12]) ? 4'b1001 : 4'b1101;
															assign node38952 = (inp[12]) ? 4'b1101 : 4'b1001;
														assign node38955 = (inp[9]) ? node38959 : node38956;
															assign node38956 = (inp[12]) ? 4'b1001 : 4'b1101;
															assign node38959 = (inp[12]) ? 4'b1111 : 4'b1001;
													assign node38962 = (inp[3]) ? node38968 : node38963;
														assign node38963 = (inp[12]) ? 4'b1011 : node38964;
															assign node38964 = (inp[9]) ? 4'b1011 : 4'b1111;
														assign node38968 = (inp[14]) ? node38970 : 4'b1011;
															assign node38970 = (inp[9]) ? node38972 : 4'b1011;
																assign node38972 = (inp[12]) ? 4'b1101 : 4'b1011;
											assign node38975 = (inp[3]) ? node39025 : node38976;
												assign node38976 = (inp[14]) ? node39004 : node38977;
													assign node38977 = (inp[15]) ? node38991 : node38978;
														assign node38978 = (inp[0]) ? node38984 : node38979;
															assign node38979 = (inp[12]) ? 4'b1011 : node38980;
																assign node38980 = (inp[9]) ? 4'b1111 : 4'b1011;
															assign node38984 = (inp[12]) ? node38988 : node38985;
																assign node38985 = (inp[9]) ? 4'b1101 : 4'b1001;
																assign node38988 = (inp[9]) ? 4'b1001 : 4'b1101;
														assign node38991 = (inp[0]) ? node38997 : node38992;
															assign node38992 = (inp[9]) ? node38994 : 4'b1101;
																assign node38994 = (inp[12]) ? 4'b1001 : 4'b1101;
															assign node38997 = (inp[12]) ? node39001 : node38998;
																assign node38998 = (inp[9]) ? 4'b1111 : 4'b1011;
																assign node39001 = (inp[9]) ? 4'b1011 : 4'b1111;
													assign node39004 = (inp[12]) ? node39014 : node39005;
														assign node39005 = (inp[9]) ? node39011 : node39006;
															assign node39006 = (inp[15]) ? node39008 : 4'b1001;
																assign node39008 = (inp[0]) ? 4'b1011 : 4'b1001;
															assign node39011 = (inp[0]) ? 4'b1101 : 4'b1111;
														assign node39014 = (inp[9]) ? node39020 : node39015;
															assign node39015 = (inp[15]) ? node39017 : 4'b1101;
																assign node39017 = (inp[0]) ? 4'b1111 : 4'b1101;
															assign node39020 = (inp[0]) ? 4'b1001 : node39021;
																assign node39021 = (inp[15]) ? 4'b1001 : 4'b1011;
												assign node39025 = (inp[0]) ? node39041 : node39026;
													assign node39026 = (inp[15]) ? node39034 : node39027;
														assign node39027 = (inp[9]) ? node39031 : node39028;
															assign node39028 = (inp[12]) ? 4'b1101 : 4'b1011;
															assign node39031 = (inp[12]) ? 4'b1001 : 4'b1101;
														assign node39034 = (inp[12]) ? node39038 : node39035;
															assign node39035 = (inp[9]) ? 4'b1111 : 4'b1001;
															assign node39038 = (inp[9]) ? 4'b1011 : 4'b1111;
													assign node39041 = (inp[15]) ? node39047 : node39042;
														assign node39042 = (inp[9]) ? node39044 : 4'b1111;
															assign node39044 = (inp[12]) ? 4'b1011 : 4'b1111;
														assign node39047 = (inp[14]) ? 4'b1101 : node39048;
															assign node39048 = (inp[9]) ? node39050 : 4'b1101;
																assign node39050 = (inp[12]) ? 4'b1001 : 4'b1101;
										assign node39054 = (inp[15]) ? node39118 : node39055;
											assign node39055 = (inp[0]) ? node39085 : node39056;
												assign node39056 = (inp[3]) ? node39070 : node39057;
													assign node39057 = (inp[9]) ? node39065 : node39058;
														assign node39058 = (inp[12]) ? node39062 : node39059;
															assign node39059 = (inp[4]) ? 4'b1011 : 4'b1111;
															assign node39062 = (inp[4]) ? 4'b1101 : 4'b1011;
														assign node39065 = (inp[12]) ? node39067 : 4'b1101;
															assign node39067 = (inp[4]) ? 4'b1001 : 4'b1101;
													assign node39070 = (inp[9]) ? node39078 : node39071;
														assign node39071 = (inp[4]) ? node39075 : node39072;
															assign node39072 = (inp[12]) ? 4'b1001 : 4'b1101;
															assign node39075 = (inp[12]) ? 4'b1101 : 4'b1001;
														assign node39078 = (inp[4]) ? node39082 : node39079;
															assign node39079 = (inp[12]) ? 4'b1101 : 4'b1001;
															assign node39082 = (inp[12]) ? 4'b1001 : 4'b1101;
												assign node39085 = (inp[3]) ? node39103 : node39086;
													assign node39086 = (inp[9]) ? node39094 : node39087;
														assign node39087 = (inp[4]) ? node39091 : node39088;
															assign node39088 = (inp[12]) ? 4'b1001 : 4'b1101;
															assign node39091 = (inp[12]) ? 4'b1111 : 4'b1001;
														assign node39094 = (inp[14]) ? node39096 : 4'b1111;
															assign node39096 = (inp[12]) ? node39100 : node39097;
																assign node39097 = (inp[4]) ? 4'b1111 : 4'b1001;
																assign node39100 = (inp[4]) ? 4'b1011 : 4'b1111;
													assign node39103 = (inp[12]) ? 4'b1111 : node39104;
														assign node39104 = (inp[14]) ? node39110 : node39105;
															assign node39105 = (inp[4]) ? node39107 : 4'b1111;
																assign node39107 = (inp[9]) ? 4'b1111 : 4'b1011;
															assign node39110 = (inp[9]) ? node39114 : node39111;
																assign node39111 = (inp[4]) ? 4'b1011 : 4'b1111;
																assign node39114 = (inp[4]) ? 4'b1111 : 4'b1011;
											assign node39118 = (inp[0]) ? node39162 : node39119;
												assign node39119 = (inp[3]) ? node39139 : node39120;
													assign node39120 = (inp[12]) ? node39128 : node39121;
														assign node39121 = (inp[4]) ? node39125 : node39122;
															assign node39122 = (inp[9]) ? 4'b1001 : 4'b1101;
															assign node39125 = (inp[9]) ? 4'b1111 : 4'b1001;
														assign node39128 = (inp[14]) ? node39134 : node39129;
															assign node39129 = (inp[4]) ? node39131 : 4'b1111;
																assign node39131 = (inp[9]) ? 4'b1011 : 4'b1111;
															assign node39134 = (inp[9]) ? 4'b1111 : node39135;
																assign node39135 = (inp[4]) ? 4'b1111 : 4'b1001;
													assign node39139 = (inp[9]) ? node39147 : node39140;
														assign node39140 = (inp[4]) ? node39144 : node39141;
															assign node39141 = (inp[12]) ? 4'b1011 : 4'b1111;
															assign node39144 = (inp[12]) ? 4'b1111 : 4'b1011;
														assign node39147 = (inp[14]) ? node39155 : node39148;
															assign node39148 = (inp[12]) ? node39152 : node39149;
																assign node39149 = (inp[4]) ? 4'b1111 : 4'b1011;
																assign node39152 = (inp[4]) ? 4'b1011 : 4'b1111;
															assign node39155 = (inp[12]) ? node39159 : node39156;
																assign node39156 = (inp[4]) ? 4'b1111 : 4'b1011;
																assign node39159 = (inp[4]) ? 4'b1011 : 4'b1111;
												assign node39162 = (inp[3]) ? node39178 : node39163;
													assign node39163 = (inp[4]) ? node39171 : node39164;
														assign node39164 = (inp[9]) ? node39168 : node39165;
															assign node39165 = (inp[12]) ? 4'b1011 : 4'b1111;
															assign node39168 = (inp[14]) ? 4'b1101 : 4'b1011;
														assign node39171 = (inp[12]) ? node39175 : node39172;
															assign node39172 = (inp[9]) ? 4'b1101 : 4'b1011;
															assign node39175 = (inp[9]) ? 4'b1001 : 4'b1101;
													assign node39178 = (inp[12]) ? node39184 : node39179;
														assign node39179 = (inp[4]) ? node39181 : 4'b1101;
															assign node39181 = (inp[9]) ? 4'b1101 : 4'b1001;
														assign node39184 = (inp[4]) ? node39188 : node39185;
															assign node39185 = (inp[9]) ? 4'b1101 : 4'b1001;
															assign node39188 = (inp[9]) ? 4'b1001 : 4'b1101;
									assign node39191 = (inp[4]) ? node39307 : node39192;
										assign node39192 = (inp[9]) ? node39240 : node39193;
											assign node39193 = (inp[3]) ? node39201 : node39194;
												assign node39194 = (inp[0]) ? node39198 : node39195;
													assign node39195 = (inp[15]) ? 4'b1001 : 4'b1011;
													assign node39198 = (inp[15]) ? 4'b1011 : 4'b1001;
												assign node39201 = (inp[14]) ? node39219 : node39202;
													assign node39202 = (inp[15]) ? node39212 : node39203;
														assign node39203 = (inp[12]) ? 4'b1001 : node39204;
															assign node39204 = (inp[0]) ? node39208 : node39205;
																assign node39205 = (inp[5]) ? 4'b1001 : 4'b1011;
																assign node39208 = (inp[5]) ? 4'b1011 : 4'b1001;
														assign node39212 = (inp[0]) ? node39216 : node39213;
															assign node39213 = (inp[5]) ? 4'b1011 : 4'b1001;
															assign node39216 = (inp[5]) ? 4'b1001 : 4'b1011;
													assign node39219 = (inp[5]) ? node39227 : node39220;
														assign node39220 = (inp[12]) ? node39222 : 4'b1011;
															assign node39222 = (inp[15]) ? node39224 : 4'b1011;
																assign node39224 = (inp[0]) ? 4'b1011 : 4'b1001;
														assign node39227 = (inp[12]) ? node39235 : node39228;
															assign node39228 = (inp[0]) ? node39232 : node39229;
																assign node39229 = (inp[15]) ? 4'b1011 : 4'b1001;
																assign node39232 = (inp[15]) ? 4'b1001 : 4'b1011;
															assign node39235 = (inp[15]) ? node39237 : 4'b1011;
																assign node39237 = (inp[0]) ? 4'b1001 : 4'b1011;
											assign node39240 = (inp[14]) ? node39282 : node39241;
												assign node39241 = (inp[12]) ? node39259 : node39242;
													assign node39242 = (inp[15]) ? node39248 : node39243;
														assign node39243 = (inp[0]) ? node39245 : 4'b1101;
															assign node39245 = (inp[5]) ? 4'b1111 : 4'b1101;
														assign node39248 = (inp[0]) ? node39254 : node39249;
															assign node39249 = (inp[5]) ? 4'b1111 : node39250;
																assign node39250 = (inp[3]) ? 4'b1111 : 4'b1101;
															assign node39254 = (inp[3]) ? 4'b1101 : node39255;
																assign node39255 = (inp[5]) ? 4'b1101 : 4'b1111;
													assign node39259 = (inp[3]) ? node39273 : node39260;
														assign node39260 = (inp[0]) ? node39268 : node39261;
															assign node39261 = (inp[5]) ? node39265 : node39262;
																assign node39262 = (inp[15]) ? 4'b1101 : 4'b1111;
																assign node39265 = (inp[15]) ? 4'b1111 : 4'b1101;
															assign node39268 = (inp[5]) ? 4'b1111 : node39269;
																assign node39269 = (inp[15]) ? 4'b1111 : 4'b1101;
														assign node39273 = (inp[5]) ? node39275 : 4'b1111;
															assign node39275 = (inp[15]) ? node39279 : node39276;
																assign node39276 = (inp[0]) ? 4'b1111 : 4'b1101;
																assign node39279 = (inp[0]) ? 4'b1101 : 4'b1111;
												assign node39282 = (inp[12]) ? node39294 : node39283;
													assign node39283 = (inp[5]) ? node39285 : 4'b1111;
														assign node39285 = (inp[3]) ? 4'b1111 : node39286;
															assign node39286 = (inp[15]) ? node39290 : node39287;
																assign node39287 = (inp[0]) ? 4'b1111 : 4'b1101;
																assign node39290 = (inp[0]) ? 4'b1101 : 4'b1111;
													assign node39294 = (inp[3]) ? node39300 : node39295;
														assign node39295 = (inp[0]) ? 4'b1111 : node39296;
															assign node39296 = (inp[5]) ? 4'b1111 : 4'b1101;
														assign node39300 = (inp[0]) ? node39304 : node39301;
															assign node39301 = (inp[15]) ? 4'b1111 : 4'b1101;
															assign node39304 = (inp[15]) ? 4'b1101 : 4'b1111;
										assign node39307 = (inp[9]) ? node39357 : node39308;
											assign node39308 = (inp[12]) ? node39336 : node39309;
												assign node39309 = (inp[0]) ? node39321 : node39310;
													assign node39310 = (inp[15]) ? node39316 : node39311;
														assign node39311 = (inp[3]) ? 4'b1101 : node39312;
															assign node39312 = (inp[5]) ? 4'b1101 : 4'b1111;
														assign node39316 = (inp[5]) ? 4'b1111 : node39317;
															assign node39317 = (inp[3]) ? 4'b1111 : 4'b1101;
													assign node39321 = (inp[5]) ? 4'b1101 : node39322;
														assign node39322 = (inp[14]) ? node39330 : node39323;
															assign node39323 = (inp[3]) ? node39327 : node39324;
																assign node39324 = (inp[15]) ? 4'b1111 : 4'b1101;
																assign node39327 = (inp[15]) ? 4'b1101 : 4'b1111;
															assign node39330 = (inp[15]) ? 4'b1101 : node39331;
																assign node39331 = (inp[3]) ? 4'b1111 : 4'b1101;
												assign node39336 = (inp[3]) ? node39350 : node39337;
													assign node39337 = (inp[15]) ? node39345 : node39338;
														assign node39338 = (inp[5]) ? node39342 : node39339;
															assign node39339 = (inp[0]) ? 4'b1101 : 4'b1111;
															assign node39342 = (inp[0]) ? 4'b1111 : 4'b1101;
														assign node39345 = (inp[0]) ? node39347 : 4'b1111;
															assign node39347 = (inp[5]) ? 4'b1101 : 4'b1111;
													assign node39350 = (inp[0]) ? node39354 : node39351;
														assign node39351 = (inp[15]) ? 4'b1111 : 4'b1101;
														assign node39354 = (inp[15]) ? 4'b1101 : 4'b1111;
											assign node39357 = (inp[14]) ? node39395 : node39358;
												assign node39358 = (inp[5]) ? node39374 : node39359;
													assign node39359 = (inp[12]) ? node39361 : 4'b1011;
														assign node39361 = (inp[15]) ? node39369 : node39362;
															assign node39362 = (inp[0]) ? node39366 : node39363;
																assign node39363 = (inp[3]) ? 4'b1001 : 4'b1011;
																assign node39366 = (inp[3]) ? 4'b1011 : 4'b1001;
															assign node39369 = (inp[3]) ? node39371 : 4'b1011;
																assign node39371 = (inp[0]) ? 4'b1001 : 4'b1011;
													assign node39374 = (inp[3]) ? node39382 : node39375;
														assign node39375 = (inp[0]) ? node39379 : node39376;
															assign node39376 = (inp[15]) ? 4'b1011 : 4'b1001;
															assign node39379 = (inp[15]) ? 4'b1001 : 4'b1011;
														assign node39382 = (inp[12]) ? node39388 : node39383;
															assign node39383 = (inp[0]) ? node39385 : 4'b1001;
																assign node39385 = (inp[15]) ? 4'b1001 : 4'b1011;
															assign node39388 = (inp[15]) ? node39392 : node39389;
																assign node39389 = (inp[0]) ? 4'b1011 : 4'b1001;
																assign node39392 = (inp[0]) ? 4'b1001 : 4'b1011;
												assign node39395 = (inp[15]) ? node39407 : node39396;
													assign node39396 = (inp[0]) ? node39402 : node39397;
														assign node39397 = (inp[5]) ? 4'b1001 : node39398;
															assign node39398 = (inp[3]) ? 4'b1001 : 4'b1011;
														assign node39402 = (inp[5]) ? 4'b1011 : node39403;
															assign node39403 = (inp[3]) ? 4'b1011 : 4'b1001;
													assign node39407 = (inp[0]) ? node39411 : node39408;
														assign node39408 = (inp[3]) ? 4'b1011 : 4'b1001;
														assign node39411 = (inp[3]) ? 4'b1001 : node39412;
															assign node39412 = (inp[5]) ? 4'b1001 : 4'b1011;
						assign node39416 = (inp[8]) ? node40584 : node39417;
							assign node39417 = (inp[14]) ? node40023 : node39418;
								assign node39418 = (inp[2]) ? node39754 : node39419;
									assign node39419 = (inp[12]) ? node39585 : node39420;
										assign node39420 = (inp[3]) ? node39496 : node39421;
											assign node39421 = (inp[5]) ? node39449 : node39422;
												assign node39422 = (inp[4]) ? node39434 : node39423;
													assign node39423 = (inp[9]) ? node39431 : node39424;
														assign node39424 = (inp[15]) ? node39428 : node39425;
															assign node39425 = (inp[0]) ? 4'b0100 : 4'b0110;
															assign node39428 = (inp[0]) ? 4'b0110 : 4'b0100;
														assign node39431 = (inp[15]) ? 4'b0000 : 4'b0010;
													assign node39434 = (inp[9]) ? node39442 : node39435;
														assign node39435 = (inp[0]) ? node39439 : node39436;
															assign node39436 = (inp[15]) ? 4'b0000 : 4'b0010;
															assign node39439 = (inp[15]) ? 4'b0010 : 4'b0000;
														assign node39442 = (inp[15]) ? node39446 : node39443;
															assign node39443 = (inp[0]) ? 4'b0100 : 4'b0110;
															assign node39446 = (inp[0]) ? 4'b0110 : 4'b0100;
												assign node39449 = (inp[9]) ? node39473 : node39450;
													assign node39450 = (inp[4]) ? node39458 : node39451;
														assign node39451 = (inp[15]) ? node39455 : node39452;
															assign node39452 = (inp[0]) ? 4'b0100 : 4'b0110;
															assign node39455 = (inp[0]) ? 4'b0110 : 4'b0100;
														assign node39458 = (inp[10]) ? node39466 : node39459;
															assign node39459 = (inp[15]) ? node39463 : node39460;
																assign node39460 = (inp[0]) ? 4'b0000 : 4'b0010;
																assign node39463 = (inp[0]) ? 4'b0010 : 4'b0000;
															assign node39466 = (inp[15]) ? node39470 : node39467;
																assign node39467 = (inp[0]) ? 4'b0000 : 4'b0010;
																assign node39470 = (inp[0]) ? 4'b0010 : 4'b0000;
													assign node39473 = (inp[4]) ? node39489 : node39474;
														assign node39474 = (inp[10]) ? node39482 : node39475;
															assign node39475 = (inp[0]) ? node39479 : node39476;
																assign node39476 = (inp[15]) ? 4'b0000 : 4'b0010;
																assign node39479 = (inp[15]) ? 4'b0010 : 4'b0000;
															assign node39482 = (inp[15]) ? node39486 : node39483;
																assign node39483 = (inp[0]) ? 4'b0000 : 4'b0010;
																assign node39486 = (inp[0]) ? 4'b0010 : 4'b0000;
														assign node39489 = (inp[0]) ? node39493 : node39490;
															assign node39490 = (inp[15]) ? 4'b0110 : 4'b0100;
															assign node39493 = (inp[15]) ? 4'b0100 : 4'b0110;
											assign node39496 = (inp[10]) ? node39540 : node39497;
												assign node39497 = (inp[0]) ? node39521 : node39498;
													assign node39498 = (inp[15]) ? node39512 : node39499;
														assign node39499 = (inp[5]) ? node39507 : node39500;
															assign node39500 = (inp[4]) ? node39504 : node39501;
																assign node39501 = (inp[9]) ? 4'b0010 : 4'b0110;
																assign node39504 = (inp[9]) ? 4'b0100 : 4'b0010;
															assign node39507 = (inp[4]) ? 4'b0100 : node39508;
																assign node39508 = (inp[9]) ? 4'b0000 : 4'b0100;
														assign node39512 = (inp[5]) ? node39516 : node39513;
															assign node39513 = (inp[4]) ? 4'b0110 : 4'b0100;
															assign node39516 = (inp[9]) ? node39518 : 4'b0110;
																assign node39518 = (inp[4]) ? 4'b0110 : 4'b0010;
													assign node39521 = (inp[5]) ? node39529 : node39522;
														assign node39522 = (inp[15]) ? 4'b0010 : node39523;
															assign node39523 = (inp[4]) ? 4'b0000 : node39524;
																assign node39524 = (inp[9]) ? 4'b0000 : 4'b0100;
														assign node39529 = (inp[15]) ? node39535 : node39530;
															assign node39530 = (inp[4]) ? 4'b0110 : node39531;
																assign node39531 = (inp[9]) ? 4'b0010 : 4'b0110;
															assign node39535 = (inp[4]) ? 4'b0100 : node39536;
																assign node39536 = (inp[9]) ? 4'b0000 : 4'b0100;
												assign node39540 = (inp[4]) ? node39562 : node39541;
													assign node39541 = (inp[9]) ? node39555 : node39542;
														assign node39542 = (inp[5]) ? node39550 : node39543;
															assign node39543 = (inp[15]) ? node39547 : node39544;
																assign node39544 = (inp[0]) ? 4'b0100 : 4'b0110;
																assign node39547 = (inp[0]) ? 4'b0110 : 4'b0100;
															assign node39550 = (inp[15]) ? 4'b0100 : node39551;
																assign node39551 = (inp[0]) ? 4'b0110 : 4'b0100;
														assign node39555 = (inp[5]) ? 4'b0000 : node39556;
															assign node39556 = (inp[15]) ? node39558 : 4'b0000;
																assign node39558 = (inp[0]) ? 4'b0010 : 4'b0000;
													assign node39562 = (inp[9]) ? node39578 : node39563;
														assign node39563 = (inp[15]) ? node39571 : node39564;
															assign node39564 = (inp[5]) ? node39568 : node39565;
																assign node39565 = (inp[0]) ? 4'b0000 : 4'b0010;
																assign node39568 = (inp[0]) ? 4'b0010 : 4'b0000;
															assign node39571 = (inp[5]) ? node39575 : node39572;
																assign node39572 = (inp[0]) ? 4'b0010 : 4'b0000;
																assign node39575 = (inp[0]) ? 4'b0000 : 4'b0010;
														assign node39578 = (inp[0]) ? node39582 : node39579;
															assign node39579 = (inp[15]) ? 4'b0110 : 4'b0100;
															assign node39582 = (inp[15]) ? 4'b0100 : 4'b0110;
										assign node39585 = (inp[0]) ? node39671 : node39586;
											assign node39586 = (inp[4]) ? node39630 : node39587;
												assign node39587 = (inp[15]) ? node39609 : node39588;
													assign node39588 = (inp[5]) ? node39594 : node39589;
														assign node39589 = (inp[10]) ? node39591 : 4'b0010;
															assign node39591 = (inp[9]) ? 4'b0110 : 4'b0010;
														assign node39594 = (inp[3]) ? node39602 : node39595;
															assign node39595 = (inp[10]) ? node39599 : node39596;
																assign node39596 = (inp[9]) ? 4'b0010 : 4'b0110;
																assign node39599 = (inp[9]) ? 4'b0100 : 4'b0010;
															assign node39602 = (inp[10]) ? node39606 : node39603;
																assign node39603 = (inp[9]) ? 4'b0000 : 4'b0100;
																assign node39606 = (inp[9]) ? 4'b0100 : 4'b0000;
													assign node39609 = (inp[3]) ? node39617 : node39610;
														assign node39610 = (inp[10]) ? node39614 : node39611;
															assign node39611 = (inp[9]) ? 4'b0000 : 4'b0100;
															assign node39614 = (inp[9]) ? 4'b0100 : 4'b0000;
														assign node39617 = (inp[5]) ? node39625 : node39618;
															assign node39618 = (inp[9]) ? node39622 : node39619;
																assign node39619 = (inp[10]) ? 4'b0000 : 4'b0100;
																assign node39622 = (inp[10]) ? 4'b0110 : 4'b0000;
															assign node39625 = (inp[9]) ? 4'b0010 : node39626;
																assign node39626 = (inp[10]) ? 4'b0010 : 4'b0110;
												assign node39630 = (inp[15]) ? node39648 : node39631;
													assign node39631 = (inp[3]) ? node39641 : node39632;
														assign node39632 = (inp[5]) ? node39636 : node39633;
															assign node39633 = (inp[9]) ? 4'b0010 : 4'b0110;
															assign node39636 = (inp[10]) ? 4'b0100 : node39637;
																assign node39637 = (inp[9]) ? 4'b0100 : 4'b0010;
														assign node39641 = (inp[10]) ? node39645 : node39642;
															assign node39642 = (inp[9]) ? 4'b0100 : 4'b0010;
															assign node39645 = (inp[9]) ? 4'b0000 : 4'b0100;
													assign node39648 = (inp[5]) ? node39662 : node39649;
														assign node39649 = (inp[3]) ? node39655 : node39650;
															assign node39650 = (inp[10]) ? 4'b0000 : node39651;
																assign node39651 = (inp[9]) ? 4'b0100 : 4'b0000;
															assign node39655 = (inp[10]) ? node39659 : node39656;
																assign node39656 = (inp[9]) ? 4'b0110 : 4'b0000;
																assign node39659 = (inp[9]) ? 4'b0010 : 4'b0110;
														assign node39662 = (inp[9]) ? node39668 : node39663;
															assign node39663 = (inp[10]) ? 4'b0110 : node39664;
																assign node39664 = (inp[3]) ? 4'b0010 : 4'b0000;
															assign node39668 = (inp[10]) ? 4'b0010 : 4'b0110;
											assign node39671 = (inp[15]) ? node39707 : node39672;
												assign node39672 = (inp[5]) ? node39684 : node39673;
													assign node39673 = (inp[9]) ? 4'b0100 : node39674;
														assign node39674 = (inp[4]) ? node39678 : node39675;
															assign node39675 = (inp[10]) ? 4'b0000 : 4'b0100;
															assign node39678 = (inp[10]) ? node39680 : 4'b0000;
																assign node39680 = (inp[3]) ? 4'b0110 : 4'b0100;
													assign node39684 = (inp[3]) ? node39694 : node39685;
														assign node39685 = (inp[10]) ? 4'b0010 : node39686;
															assign node39686 = (inp[4]) ? node39690 : node39687;
																assign node39687 = (inp[9]) ? 4'b0000 : 4'b0100;
																assign node39690 = (inp[9]) ? 4'b0110 : 4'b0000;
														assign node39694 = (inp[10]) ? node39700 : node39695;
															assign node39695 = (inp[9]) ? node39697 : 4'b0010;
																assign node39697 = (inp[4]) ? 4'b0110 : 4'b0010;
															assign node39700 = (inp[9]) ? node39704 : node39701;
																assign node39701 = (inp[4]) ? 4'b0110 : 4'b0010;
																assign node39704 = (inp[4]) ? 4'b0010 : 4'b0110;
												assign node39707 = (inp[5]) ? node39735 : node39708;
													assign node39708 = (inp[3]) ? node39724 : node39709;
														assign node39709 = (inp[10]) ? node39717 : node39710;
															assign node39710 = (inp[9]) ? node39714 : node39711;
																assign node39711 = (inp[4]) ? 4'b0010 : 4'b0110;
																assign node39714 = (inp[4]) ? 4'b0110 : 4'b0010;
															assign node39717 = (inp[4]) ? node39721 : node39718;
																assign node39718 = (inp[9]) ? 4'b0110 : 4'b0010;
																assign node39721 = (inp[9]) ? 4'b0010 : 4'b0110;
														assign node39724 = (inp[4]) ? node39730 : node39725;
															assign node39725 = (inp[10]) ? 4'b0010 : node39726;
																assign node39726 = (inp[9]) ? 4'b0010 : 4'b0110;
															assign node39730 = (inp[10]) ? node39732 : 4'b0010;
																assign node39732 = (inp[9]) ? 4'b0000 : 4'b0100;
													assign node39735 = (inp[3]) ? node39749 : node39736;
														assign node39736 = (inp[4]) ? node39742 : node39737;
															assign node39737 = (inp[9]) ? 4'b0010 : node39738;
																assign node39738 = (inp[10]) ? 4'b0010 : 4'b0110;
															assign node39742 = (inp[10]) ? node39746 : node39743;
																assign node39743 = (inp[9]) ? 4'b0100 : 4'b0010;
																assign node39746 = (inp[9]) ? 4'b0000 : 4'b0100;
														assign node39749 = (inp[9]) ? node39751 : 4'b0100;
															assign node39751 = (inp[4]) ? 4'b0000 : 4'b0100;
									assign node39754 = (inp[0]) ? node39876 : node39755;
										assign node39755 = (inp[15]) ? node39817 : node39756;
											assign node39756 = (inp[3]) ? node39792 : node39757;
												assign node39757 = (inp[5]) ? node39773 : node39758;
													assign node39758 = (inp[12]) ? 4'b1111 : node39759;
														assign node39759 = (inp[4]) ? node39767 : node39760;
															assign node39760 = (inp[9]) ? node39764 : node39761;
																assign node39761 = (inp[10]) ? 4'b1011 : 4'b1111;
																assign node39764 = (inp[10]) ? 4'b1111 : 4'b1011;
															assign node39767 = (inp[9]) ? 4'b1111 : node39768;
																assign node39768 = (inp[10]) ? 4'b1111 : 4'b1011;
													assign node39773 = (inp[10]) ? node39785 : node39774;
														assign node39774 = (inp[4]) ? node39780 : node39775;
															assign node39775 = (inp[9]) ? 4'b1011 : node39776;
																assign node39776 = (inp[12]) ? 4'b1011 : 4'b1111;
															assign node39780 = (inp[9]) ? 4'b1101 : node39781;
																assign node39781 = (inp[12]) ? 4'b1101 : 4'b1011;
														assign node39785 = (inp[4]) ? node39789 : node39786;
															assign node39786 = (inp[9]) ? 4'b1101 : 4'b1011;
															assign node39789 = (inp[9]) ? 4'b1001 : 4'b1101;
												assign node39792 = (inp[9]) ? node39806 : node39793;
													assign node39793 = (inp[4]) ? node39801 : node39794;
														assign node39794 = (inp[5]) ? node39798 : node39795;
															assign node39795 = (inp[12]) ? 4'b1011 : 4'b1111;
															assign node39798 = (inp[12]) ? 4'b1001 : 4'b1101;
														assign node39801 = (inp[10]) ? 4'b1101 : node39802;
															assign node39802 = (inp[12]) ? 4'b1101 : 4'b1011;
													assign node39806 = (inp[4]) ? node39812 : node39807;
														assign node39807 = (inp[12]) ? 4'b1101 : node39808;
															assign node39808 = (inp[10]) ? 4'b1101 : 4'b1001;
														assign node39812 = (inp[10]) ? 4'b1001 : node39813;
															assign node39813 = (inp[12]) ? 4'b1001 : 4'b1101;
											assign node39817 = (inp[5]) ? node39853 : node39818;
												assign node39818 = (inp[3]) ? node39840 : node39819;
													assign node39819 = (inp[12]) ? node39831 : node39820;
														assign node39820 = (inp[10]) ? node39826 : node39821;
															assign node39821 = (inp[9]) ? node39823 : 4'b1101;
																assign node39823 = (inp[4]) ? 4'b1101 : 4'b1001;
															assign node39826 = (inp[4]) ? 4'b1001 : node39827;
																assign node39827 = (inp[9]) ? 4'b1101 : 4'b1001;
														assign node39831 = (inp[10]) ? node39837 : node39832;
															assign node39832 = (inp[4]) ? node39834 : 4'b1001;
																assign node39834 = (inp[9]) ? 4'b1001 : 4'b1101;
															assign node39837 = (inp[4]) ? 4'b1001 : 4'b1101;
													assign node39840 = (inp[9]) ? node39846 : node39841;
														assign node39841 = (inp[4]) ? node39843 : 4'b1001;
															assign node39843 = (inp[12]) ? 4'b1111 : 4'b1001;
														assign node39846 = (inp[4]) ? 4'b1011 : node39847;
															assign node39847 = (inp[12]) ? 4'b1111 : node39848;
																assign node39848 = (inp[10]) ? 4'b1111 : 4'b1001;
												assign node39853 = (inp[9]) ? node39865 : node39854;
													assign node39854 = (inp[3]) ? node39862 : node39855;
														assign node39855 = (inp[4]) ? node39859 : node39856;
															assign node39856 = (inp[12]) ? 4'b1001 : 4'b1101;
															assign node39859 = (inp[10]) ? 4'b1111 : 4'b1001;
														assign node39862 = (inp[4]) ? 4'b1111 : 4'b1011;
													assign node39865 = (inp[4]) ? node39871 : node39866;
														assign node39866 = (inp[10]) ? 4'b1111 : node39867;
															assign node39867 = (inp[12]) ? 4'b1111 : 4'b1011;
														assign node39871 = (inp[12]) ? 4'b1011 : node39872;
															assign node39872 = (inp[10]) ? 4'b1011 : 4'b1111;
										assign node39876 = (inp[15]) ? node39954 : node39877;
											assign node39877 = (inp[3]) ? node39907 : node39878;
												assign node39878 = (inp[5]) ? node39892 : node39879;
													assign node39879 = (inp[10]) ? node39885 : node39880;
														assign node39880 = (inp[12]) ? 4'b1001 : node39881;
															assign node39881 = (inp[9]) ? 4'b1001 : 4'b1101;
														assign node39885 = (inp[4]) ? node39889 : node39886;
															assign node39886 = (inp[9]) ? 4'b1101 : 4'b1001;
															assign node39889 = (inp[9]) ? 4'b1001 : 4'b1101;
													assign node39892 = (inp[4]) ? node39900 : node39893;
														assign node39893 = (inp[9]) ? node39897 : node39894;
															assign node39894 = (inp[10]) ? 4'b1001 : 4'b1101;
															assign node39897 = (inp[10]) ? 4'b1111 : 4'b1001;
														assign node39900 = (inp[12]) ? node39904 : node39901;
															assign node39901 = (inp[9]) ? 4'b1111 : 4'b1001;
															assign node39904 = (inp[9]) ? 4'b1011 : 4'b1111;
												assign node39907 = (inp[5]) ? node39929 : node39908;
													assign node39908 = (inp[9]) ? node39918 : node39909;
														assign node39909 = (inp[4]) ? node39913 : node39910;
															assign node39910 = (inp[10]) ? 4'b1001 : 4'b1101;
															assign node39913 = (inp[10]) ? 4'b1111 : node39914;
																assign node39914 = (inp[12]) ? 4'b1111 : 4'b1001;
														assign node39918 = (inp[4]) ? node39924 : node39919;
															assign node39919 = (inp[12]) ? 4'b1111 : node39920;
																assign node39920 = (inp[10]) ? 4'b1111 : 4'b1001;
															assign node39924 = (inp[10]) ? 4'b1011 : node39925;
																assign node39925 = (inp[12]) ? 4'b1011 : 4'b1111;
													assign node39929 = (inp[10]) ? node39939 : node39930;
														assign node39930 = (inp[4]) ? 4'b1111 : node39931;
															assign node39931 = (inp[9]) ? node39935 : node39932;
																assign node39932 = (inp[12]) ? 4'b1011 : 4'b1111;
																assign node39935 = (inp[12]) ? 4'b1111 : 4'b1011;
														assign node39939 = (inp[12]) ? node39947 : node39940;
															assign node39940 = (inp[4]) ? node39944 : node39941;
																assign node39941 = (inp[9]) ? 4'b1111 : 4'b1011;
																assign node39944 = (inp[9]) ? 4'b1011 : 4'b1111;
															assign node39947 = (inp[9]) ? node39951 : node39948;
																assign node39948 = (inp[4]) ? 4'b1111 : 4'b1011;
																assign node39951 = (inp[4]) ? 4'b1011 : 4'b1111;
											assign node39954 = (inp[5]) ? node39994 : node39955;
												assign node39955 = (inp[3]) ? node39971 : node39956;
													assign node39956 = (inp[9]) ? node39964 : node39957;
														assign node39957 = (inp[4]) ? 4'b1111 : node39958;
															assign node39958 = (inp[10]) ? 4'b1011 : node39959;
																assign node39959 = (inp[12]) ? 4'b1011 : 4'b1111;
														assign node39964 = (inp[4]) ? 4'b1011 : node39965;
															assign node39965 = (inp[12]) ? 4'b1111 : node39966;
																assign node39966 = (inp[10]) ? 4'b1111 : 4'b1011;
													assign node39971 = (inp[12]) ? node39983 : node39972;
														assign node39972 = (inp[4]) ? node39978 : node39973;
															assign node39973 = (inp[9]) ? 4'b1011 : node39974;
																assign node39974 = (inp[10]) ? 4'b1011 : 4'b1111;
															assign node39978 = (inp[10]) ? 4'b1101 : node39979;
																assign node39979 = (inp[9]) ? 4'b1101 : 4'b1011;
														assign node39983 = (inp[10]) ? node39989 : node39984;
															assign node39984 = (inp[9]) ? node39986 : 4'b1011;
																assign node39986 = (inp[4]) ? 4'b1001 : 4'b1101;
															assign node39989 = (inp[9]) ? node39991 : 4'b1101;
																assign node39991 = (inp[4]) ? 4'b1001 : 4'b1101;
												assign node39994 = (inp[3]) ? node40008 : node39995;
													assign node39995 = (inp[12]) ? node40001 : node39996;
														assign node39996 = (inp[4]) ? node39998 : 4'b1011;
															assign node39998 = (inp[9]) ? 4'b1101 : 4'b1011;
														assign node40001 = (inp[4]) ? node40005 : node40002;
															assign node40002 = (inp[9]) ? 4'b1101 : 4'b1011;
															assign node40005 = (inp[9]) ? 4'b1001 : 4'b1101;
													assign node40008 = (inp[12]) ? node40018 : node40009;
														assign node40009 = (inp[10]) ? 4'b1001 : node40010;
															assign node40010 = (inp[4]) ? node40014 : node40011;
																assign node40011 = (inp[9]) ? 4'b1001 : 4'b1101;
																assign node40014 = (inp[9]) ? 4'b1101 : 4'b1001;
														assign node40018 = (inp[9]) ? 4'b1101 : node40019;
															assign node40019 = (inp[4]) ? 4'b1101 : 4'b1001;
								assign node40023 = (inp[10]) ? node40301 : node40024;
									assign node40024 = (inp[3]) ? node40160 : node40025;
										assign node40025 = (inp[15]) ? node40087 : node40026;
											assign node40026 = (inp[0]) ? node40058 : node40027;
												assign node40027 = (inp[5]) ? node40043 : node40028;
													assign node40028 = (inp[9]) ? node40038 : node40029;
														assign node40029 = (inp[2]) ? node40031 : 4'b1111;
															assign node40031 = (inp[4]) ? node40035 : node40032;
																assign node40032 = (inp[12]) ? 4'b1011 : 4'b1111;
																assign node40035 = (inp[12]) ? 4'b1111 : 4'b1011;
														assign node40038 = (inp[4]) ? node40040 : 4'b1011;
															assign node40040 = (inp[12]) ? 4'b1011 : 4'b1111;
													assign node40043 = (inp[9]) ? node40051 : node40044;
														assign node40044 = (inp[4]) ? node40048 : node40045;
															assign node40045 = (inp[12]) ? 4'b1011 : 4'b1111;
															assign node40048 = (inp[12]) ? 4'b1101 : 4'b1011;
														assign node40051 = (inp[4]) ? node40055 : node40052;
															assign node40052 = (inp[12]) ? 4'b1101 : 4'b1011;
															assign node40055 = (inp[12]) ? 4'b1001 : 4'b1101;
												assign node40058 = (inp[5]) ? node40074 : node40059;
													assign node40059 = (inp[4]) ? node40065 : node40060;
														assign node40060 = (inp[2]) ? node40062 : 4'b1001;
															assign node40062 = (inp[9]) ? 4'b1101 : 4'b1001;
														assign node40065 = (inp[2]) ? 4'b1101 : node40066;
															assign node40066 = (inp[12]) ? node40070 : node40067;
																assign node40067 = (inp[9]) ? 4'b1101 : 4'b1001;
																assign node40070 = (inp[9]) ? 4'b1001 : 4'b1101;
													assign node40074 = (inp[9]) ? node40080 : node40075;
														assign node40075 = (inp[12]) ? node40077 : 4'b1001;
															assign node40077 = (inp[4]) ? 4'b1111 : 4'b1001;
														assign node40080 = (inp[12]) ? node40084 : node40081;
															assign node40081 = (inp[4]) ? 4'b1111 : 4'b1001;
															assign node40084 = (inp[4]) ? 4'b1011 : 4'b1111;
											assign node40087 = (inp[0]) ? node40133 : node40088;
												assign node40088 = (inp[5]) ? node40114 : node40089;
													assign node40089 = (inp[4]) ? node40103 : node40090;
														assign node40090 = (inp[2]) ? node40098 : node40091;
															assign node40091 = (inp[9]) ? node40095 : node40092;
																assign node40092 = (inp[12]) ? 4'b1001 : 4'b1101;
																assign node40095 = (inp[12]) ? 4'b1101 : 4'b1001;
															assign node40098 = (inp[9]) ? 4'b1101 : node40099;
																assign node40099 = (inp[12]) ? 4'b1001 : 4'b1101;
														assign node40103 = (inp[2]) ? node40109 : node40104;
															assign node40104 = (inp[12]) ? node40106 : 4'b1001;
																assign node40106 = (inp[9]) ? 4'b1001 : 4'b1101;
															assign node40109 = (inp[12]) ? 4'b1001 : node40110;
																assign node40110 = (inp[9]) ? 4'b1101 : 4'b1001;
													assign node40114 = (inp[12]) ? node40122 : node40115;
														assign node40115 = (inp[4]) ? node40119 : node40116;
															assign node40116 = (inp[9]) ? 4'b1001 : 4'b1101;
															assign node40119 = (inp[9]) ? 4'b1111 : 4'b1001;
														assign node40122 = (inp[2]) ? node40128 : node40123;
															assign node40123 = (inp[9]) ? node40125 : 4'b1111;
																assign node40125 = (inp[4]) ? 4'b1011 : 4'b1111;
															assign node40128 = (inp[4]) ? node40130 : 4'b1001;
																assign node40130 = (inp[9]) ? 4'b1011 : 4'b1111;
												assign node40133 = (inp[5]) ? node40147 : node40134;
													assign node40134 = (inp[9]) ? node40142 : node40135;
														assign node40135 = (inp[12]) ? node40139 : node40136;
															assign node40136 = (inp[4]) ? 4'b1011 : 4'b1111;
															assign node40139 = (inp[4]) ? 4'b1111 : 4'b1011;
														assign node40142 = (inp[4]) ? 4'b1011 : node40143;
															assign node40143 = (inp[12]) ? 4'b1111 : 4'b1011;
													assign node40147 = (inp[12]) ? node40155 : node40148;
														assign node40148 = (inp[2]) ? node40150 : 4'b1011;
															assign node40150 = (inp[9]) ? 4'b1101 : node40151;
																assign node40151 = (inp[4]) ? 4'b1011 : 4'b1111;
														assign node40155 = (inp[4]) ? node40157 : 4'b1101;
															assign node40157 = (inp[9]) ? 4'b1001 : 4'b1101;
										assign node40160 = (inp[12]) ? node40222 : node40161;
											assign node40161 = (inp[9]) ? node40193 : node40162;
												assign node40162 = (inp[4]) ? node40178 : node40163;
													assign node40163 = (inp[5]) ? node40171 : node40164;
														assign node40164 = (inp[0]) ? node40168 : node40165;
															assign node40165 = (inp[15]) ? 4'b1101 : 4'b1111;
															assign node40168 = (inp[15]) ? 4'b1111 : 4'b1101;
														assign node40171 = (inp[0]) ? node40175 : node40172;
															assign node40172 = (inp[15]) ? 4'b1111 : 4'b1101;
															assign node40175 = (inp[15]) ? 4'b1101 : 4'b1111;
													assign node40178 = (inp[2]) ? node40184 : node40179;
														assign node40179 = (inp[5]) ? 4'b1001 : node40180;
															assign node40180 = (inp[0]) ? 4'b1011 : 4'b1001;
														assign node40184 = (inp[0]) ? node40186 : 4'b1011;
															assign node40186 = (inp[15]) ? node40190 : node40187;
																assign node40187 = (inp[5]) ? 4'b1011 : 4'b1001;
																assign node40190 = (inp[5]) ? 4'b1001 : 4'b1011;
												assign node40193 = (inp[4]) ? node40215 : node40194;
													assign node40194 = (inp[5]) ? node40208 : node40195;
														assign node40195 = (inp[2]) ? node40203 : node40196;
															assign node40196 = (inp[0]) ? node40200 : node40197;
																assign node40197 = (inp[15]) ? 4'b1001 : 4'b1011;
																assign node40200 = (inp[15]) ? 4'b1011 : 4'b1001;
															assign node40203 = (inp[15]) ? node40205 : 4'b1001;
																assign node40205 = (inp[0]) ? 4'b1011 : 4'b1001;
														assign node40208 = (inp[0]) ? node40212 : node40209;
															assign node40209 = (inp[15]) ? 4'b1011 : 4'b1001;
															assign node40212 = (inp[15]) ? 4'b1001 : 4'b1011;
													assign node40215 = (inp[0]) ? node40219 : node40216;
														assign node40216 = (inp[15]) ? 4'b1111 : 4'b1101;
														assign node40219 = (inp[15]) ? 4'b1101 : 4'b1111;
											assign node40222 = (inp[4]) ? node40268 : node40223;
												assign node40223 = (inp[9]) ? node40243 : node40224;
													assign node40224 = (inp[15]) ? node40236 : node40225;
														assign node40225 = (inp[2]) ? node40231 : node40226;
															assign node40226 = (inp[5]) ? node40228 : 4'b1001;
																assign node40228 = (inp[0]) ? 4'b1011 : 4'b1001;
															assign node40231 = (inp[0]) ? node40233 : 4'b1011;
																assign node40233 = (inp[5]) ? 4'b1011 : 4'b1001;
														assign node40236 = (inp[2]) ? 4'b1001 : node40237;
															assign node40237 = (inp[5]) ? 4'b1001 : node40238;
																assign node40238 = (inp[0]) ? 4'b1011 : 4'b1001;
													assign node40243 = (inp[5]) ? node40255 : node40244;
														assign node40244 = (inp[2]) ? node40250 : node40245;
															assign node40245 = (inp[0]) ? 4'b1101 : node40246;
																assign node40246 = (inp[15]) ? 4'b1111 : 4'b1101;
															assign node40250 = (inp[15]) ? 4'b1101 : node40251;
																assign node40251 = (inp[0]) ? 4'b1111 : 4'b1101;
														assign node40255 = (inp[2]) ? node40263 : node40256;
															assign node40256 = (inp[15]) ? node40260 : node40257;
																assign node40257 = (inp[0]) ? 4'b1111 : 4'b1101;
																assign node40260 = (inp[0]) ? 4'b1101 : 4'b1111;
															assign node40263 = (inp[0]) ? 4'b1111 : node40264;
																assign node40264 = (inp[15]) ? 4'b1111 : 4'b1101;
												assign node40268 = (inp[9]) ? node40280 : node40269;
													assign node40269 = (inp[2]) ? node40277 : node40270;
														assign node40270 = (inp[5]) ? node40272 : 4'b1101;
															assign node40272 = (inp[0]) ? 4'b1101 : node40273;
																assign node40273 = (inp[15]) ? 4'b1111 : 4'b1101;
														assign node40277 = (inp[15]) ? 4'b1101 : 4'b1111;
													assign node40280 = (inp[5]) ? node40288 : node40281;
														assign node40281 = (inp[15]) ? node40285 : node40282;
															assign node40282 = (inp[0]) ? 4'b1011 : 4'b1001;
															assign node40285 = (inp[0]) ? 4'b1001 : 4'b1011;
														assign node40288 = (inp[2]) ? node40296 : node40289;
															assign node40289 = (inp[0]) ? node40293 : node40290;
																assign node40290 = (inp[15]) ? 4'b1011 : 4'b1001;
																assign node40293 = (inp[15]) ? 4'b1001 : 4'b1011;
															assign node40296 = (inp[0]) ? 4'b1001 : node40297;
																assign node40297 = (inp[15]) ? 4'b1011 : 4'b1001;
									assign node40301 = (inp[12]) ? node40477 : node40302;
										assign node40302 = (inp[2]) ? node40396 : node40303;
											assign node40303 = (inp[3]) ? node40341 : node40304;
												assign node40304 = (inp[9]) ? node40322 : node40305;
													assign node40305 = (inp[4]) ? node40309 : node40306;
														assign node40306 = (inp[5]) ? 4'b1001 : 4'b1011;
														assign node40309 = (inp[0]) ? node40317 : node40310;
															assign node40310 = (inp[5]) ? node40314 : node40311;
																assign node40311 = (inp[15]) ? 4'b1101 : 4'b1111;
																assign node40314 = (inp[15]) ? 4'b1111 : 4'b1101;
															assign node40317 = (inp[5]) ? 4'b1101 : node40318;
																assign node40318 = (inp[15]) ? 4'b1111 : 4'b1101;
													assign node40322 = (inp[4]) ? node40328 : node40323;
														assign node40323 = (inp[5]) ? node40325 : 4'b1101;
															assign node40325 = (inp[15]) ? 4'b1101 : 4'b1111;
														assign node40328 = (inp[15]) ? node40336 : node40329;
															assign node40329 = (inp[0]) ? node40333 : node40330;
																assign node40330 = (inp[5]) ? 4'b1001 : 4'b1011;
																assign node40333 = (inp[5]) ? 4'b1011 : 4'b1001;
															assign node40336 = (inp[0]) ? node40338 : 4'b1001;
																assign node40338 = (inp[5]) ? 4'b1001 : 4'b1011;
												assign node40341 = (inp[5]) ? node40371 : node40342;
													assign node40342 = (inp[0]) ? node40358 : node40343;
														assign node40343 = (inp[15]) ? node40351 : node40344;
															assign node40344 = (inp[9]) ? node40348 : node40345;
																assign node40345 = (inp[4]) ? 4'b1101 : 4'b1011;
																assign node40348 = (inp[4]) ? 4'b1001 : 4'b1101;
															assign node40351 = (inp[9]) ? node40355 : node40352;
																assign node40352 = (inp[4]) ? 4'b1111 : 4'b1001;
																assign node40355 = (inp[4]) ? 4'b1011 : 4'b1111;
														assign node40358 = (inp[15]) ? node40364 : node40359;
															assign node40359 = (inp[4]) ? 4'b1111 : node40360;
																assign node40360 = (inp[9]) ? 4'b1111 : 4'b1001;
															assign node40364 = (inp[4]) ? node40368 : node40365;
																assign node40365 = (inp[9]) ? 4'b1101 : 4'b1011;
																assign node40368 = (inp[9]) ? 4'b1001 : 4'b1101;
													assign node40371 = (inp[15]) ? node40385 : node40372;
														assign node40372 = (inp[0]) ? node40378 : node40373;
															assign node40373 = (inp[9]) ? node40375 : 4'b1001;
																assign node40375 = (inp[4]) ? 4'b1001 : 4'b1101;
															assign node40378 = (inp[9]) ? node40382 : node40379;
																assign node40379 = (inp[4]) ? 4'b1111 : 4'b1011;
																assign node40382 = (inp[4]) ? 4'b1011 : 4'b1111;
														assign node40385 = (inp[0]) ? node40393 : node40386;
															assign node40386 = (inp[4]) ? node40390 : node40387;
																assign node40387 = (inp[9]) ? 4'b1111 : 4'b1011;
																assign node40390 = (inp[9]) ? 4'b1011 : 4'b1111;
															assign node40393 = (inp[4]) ? 4'b1101 : 4'b1001;
											assign node40396 = (inp[9]) ? node40440 : node40397;
												assign node40397 = (inp[4]) ? node40415 : node40398;
													assign node40398 = (inp[15]) ? node40408 : node40399;
														assign node40399 = (inp[0]) ? node40403 : node40400;
															assign node40400 = (inp[5]) ? 4'b1001 : 4'b1011;
															assign node40403 = (inp[3]) ? node40405 : 4'b1001;
																assign node40405 = (inp[5]) ? 4'b1011 : 4'b1001;
														assign node40408 = (inp[0]) ? 4'b1011 : node40409;
															assign node40409 = (inp[3]) ? node40411 : 4'b1001;
																assign node40411 = (inp[5]) ? 4'b1011 : 4'b1001;
													assign node40415 = (inp[5]) ? node40425 : node40416;
														assign node40416 = (inp[3]) ? 4'b1101 : node40417;
															assign node40417 = (inp[15]) ? node40421 : node40418;
																assign node40418 = (inp[0]) ? 4'b1101 : 4'b1111;
																assign node40421 = (inp[0]) ? 4'b1111 : 4'b1101;
														assign node40425 = (inp[3]) ? node40433 : node40426;
															assign node40426 = (inp[15]) ? node40430 : node40427;
																assign node40427 = (inp[0]) ? 4'b1111 : 4'b1101;
																assign node40430 = (inp[0]) ? 4'b1101 : 4'b1111;
															assign node40433 = (inp[15]) ? node40437 : node40434;
																assign node40434 = (inp[0]) ? 4'b1111 : 4'b1101;
																assign node40437 = (inp[0]) ? 4'b1101 : 4'b1111;
												assign node40440 = (inp[4]) ? node40462 : node40441;
													assign node40441 = (inp[15]) ? node40453 : node40442;
														assign node40442 = (inp[0]) ? node40448 : node40443;
															assign node40443 = (inp[3]) ? 4'b1101 : node40444;
																assign node40444 = (inp[5]) ? 4'b1101 : 4'b1111;
															assign node40448 = (inp[5]) ? 4'b1111 : node40449;
																assign node40449 = (inp[3]) ? 4'b1111 : 4'b1101;
														assign node40453 = (inp[0]) ? node40457 : node40454;
															assign node40454 = (inp[3]) ? 4'b1111 : 4'b1101;
															assign node40457 = (inp[5]) ? 4'b1101 : node40458;
																assign node40458 = (inp[3]) ? 4'b1101 : 4'b1111;
													assign node40462 = (inp[0]) ? node40472 : node40463;
														assign node40463 = (inp[5]) ? 4'b1011 : node40464;
															assign node40464 = (inp[3]) ? node40468 : node40465;
																assign node40465 = (inp[15]) ? 4'b1001 : 4'b1011;
																assign node40468 = (inp[15]) ? 4'b1011 : 4'b1001;
														assign node40472 = (inp[15]) ? node40474 : 4'b1011;
															assign node40474 = (inp[5]) ? 4'b1001 : 4'b1011;
										assign node40477 = (inp[15]) ? node40533 : node40478;
											assign node40478 = (inp[0]) ? node40510 : node40479;
												assign node40479 = (inp[5]) ? node40495 : node40480;
													assign node40480 = (inp[3]) ? node40488 : node40481;
														assign node40481 = (inp[4]) ? node40485 : node40482;
															assign node40482 = (inp[9]) ? 4'b1111 : 4'b1011;
															assign node40485 = (inp[9]) ? 4'b1011 : 4'b1111;
														assign node40488 = (inp[9]) ? node40492 : node40489;
															assign node40489 = (inp[4]) ? 4'b1101 : 4'b1011;
															assign node40492 = (inp[4]) ? 4'b1001 : 4'b1101;
													assign node40495 = (inp[3]) ? node40503 : node40496;
														assign node40496 = (inp[4]) ? node40500 : node40497;
															assign node40497 = (inp[9]) ? 4'b1101 : 4'b1011;
															assign node40500 = (inp[9]) ? 4'b1001 : 4'b1101;
														assign node40503 = (inp[4]) ? node40507 : node40504;
															assign node40504 = (inp[9]) ? 4'b1101 : 4'b1001;
															assign node40507 = (inp[9]) ? 4'b1001 : 4'b1101;
												assign node40510 = (inp[3]) ? node40524 : node40511;
													assign node40511 = (inp[5]) ? node40517 : node40512;
														assign node40512 = (inp[9]) ? 4'b1101 : node40513;
															assign node40513 = (inp[4]) ? 4'b1101 : 4'b1001;
														assign node40517 = (inp[4]) ? node40521 : node40518;
															assign node40518 = (inp[9]) ? 4'b1111 : 4'b1001;
															assign node40521 = (inp[9]) ? 4'b1011 : 4'b1111;
													assign node40524 = (inp[4]) ? node40530 : node40525;
														assign node40525 = (inp[9]) ? 4'b1111 : node40526;
															assign node40526 = (inp[5]) ? 4'b1011 : 4'b1001;
														assign node40530 = (inp[9]) ? 4'b1011 : 4'b1111;
											assign node40533 = (inp[0]) ? node40561 : node40534;
												assign node40534 = (inp[3]) ? node40552 : node40535;
													assign node40535 = (inp[5]) ? node40545 : node40536;
														assign node40536 = (inp[2]) ? node40538 : 4'b1101;
															assign node40538 = (inp[9]) ? node40542 : node40539;
																assign node40539 = (inp[4]) ? 4'b1101 : 4'b1001;
																assign node40542 = (inp[4]) ? 4'b1001 : 4'b1101;
														assign node40545 = (inp[4]) ? node40549 : node40546;
															assign node40546 = (inp[9]) ? 4'b1111 : 4'b1001;
															assign node40549 = (inp[9]) ? 4'b1011 : 4'b1111;
													assign node40552 = (inp[9]) ? node40558 : node40553;
														assign node40553 = (inp[4]) ? 4'b1111 : node40554;
															assign node40554 = (inp[5]) ? 4'b1011 : 4'b1001;
														assign node40558 = (inp[4]) ? 4'b1011 : 4'b1111;
												assign node40561 = (inp[3]) ? node40575 : node40562;
													assign node40562 = (inp[5]) ? node40568 : node40563;
														assign node40563 = (inp[9]) ? node40565 : 4'b1111;
															assign node40565 = (inp[4]) ? 4'b1011 : 4'b1111;
														assign node40568 = (inp[4]) ? node40572 : node40569;
															assign node40569 = (inp[9]) ? 4'b1101 : 4'b1011;
															assign node40572 = (inp[9]) ? 4'b1001 : 4'b1101;
													assign node40575 = (inp[4]) ? node40581 : node40576;
														assign node40576 = (inp[9]) ? 4'b1101 : node40577;
															assign node40577 = (inp[5]) ? 4'b1001 : 4'b1011;
														assign node40581 = (inp[9]) ? 4'b1001 : 4'b1101;
							assign node40584 = (inp[2]) ? node41150 : node40585;
								assign node40585 = (inp[14]) ? node40873 : node40586;
									assign node40586 = (inp[3]) ? node40758 : node40587;
										assign node40587 = (inp[10]) ? node40673 : node40588;
											assign node40588 = (inp[12]) ? node40634 : node40589;
												assign node40589 = (inp[9]) ? node40613 : node40590;
													assign node40590 = (inp[4]) ? node40600 : node40591;
														assign node40591 = (inp[5]) ? node40593 : 4'b1101;
															assign node40593 = (inp[15]) ? node40597 : node40594;
																assign node40594 = (inp[0]) ? 4'b1101 : 4'b1111;
																assign node40597 = (inp[0]) ? 4'b1111 : 4'b1101;
														assign node40600 = (inp[5]) ? node40608 : node40601;
															assign node40601 = (inp[0]) ? node40605 : node40602;
																assign node40602 = (inp[15]) ? 4'b1001 : 4'b1011;
																assign node40605 = (inp[15]) ? 4'b1011 : 4'b1001;
															assign node40608 = (inp[0]) ? node40610 : 4'b1001;
																assign node40610 = (inp[15]) ? 4'b1011 : 4'b1001;
													assign node40613 = (inp[4]) ? node40621 : node40614;
														assign node40614 = (inp[15]) ? node40618 : node40615;
															assign node40615 = (inp[0]) ? 4'b1001 : 4'b1011;
															assign node40618 = (inp[0]) ? 4'b1011 : 4'b1001;
														assign node40621 = (inp[5]) ? node40627 : node40622;
															assign node40622 = (inp[15]) ? 4'b1111 : node40623;
																assign node40623 = (inp[0]) ? 4'b1101 : 4'b1111;
															assign node40627 = (inp[15]) ? node40631 : node40628;
																assign node40628 = (inp[0]) ? 4'b1111 : 4'b1101;
																assign node40631 = (inp[0]) ? 4'b1101 : 4'b1111;
												assign node40634 = (inp[5]) ? node40656 : node40635;
													assign node40635 = (inp[9]) ? node40649 : node40636;
														assign node40636 = (inp[4]) ? node40644 : node40637;
															assign node40637 = (inp[0]) ? node40641 : node40638;
																assign node40638 = (inp[15]) ? 4'b1001 : 4'b1011;
																assign node40641 = (inp[15]) ? 4'b1011 : 4'b1001;
															assign node40644 = (inp[0]) ? 4'b1101 : node40645;
																assign node40645 = (inp[15]) ? 4'b1101 : 4'b1111;
														assign node40649 = (inp[4]) ? node40651 : 4'b1101;
															assign node40651 = (inp[15]) ? node40653 : 4'b1001;
																assign node40653 = (inp[0]) ? 4'b1011 : 4'b1001;
													assign node40656 = (inp[9]) ? node40664 : node40657;
														assign node40657 = (inp[15]) ? node40661 : node40658;
															assign node40658 = (inp[0]) ? 4'b1001 : 4'b1011;
															assign node40661 = (inp[0]) ? 4'b1011 : 4'b1001;
														assign node40664 = (inp[4]) ? node40668 : node40665;
															assign node40665 = (inp[0]) ? 4'b1101 : 4'b1111;
															assign node40668 = (inp[15]) ? node40670 : 4'b1001;
																assign node40670 = (inp[0]) ? 4'b1001 : 4'b1011;
											assign node40673 = (inp[5]) ? node40709 : node40674;
												assign node40674 = (inp[4]) ? node40688 : node40675;
													assign node40675 = (inp[9]) ? node40683 : node40676;
														assign node40676 = (inp[15]) ? node40680 : node40677;
															assign node40677 = (inp[0]) ? 4'b1001 : 4'b1011;
															assign node40680 = (inp[0]) ? 4'b1011 : 4'b1001;
														assign node40683 = (inp[0]) ? node40685 : 4'b1101;
															assign node40685 = (inp[15]) ? 4'b1111 : 4'b1101;
													assign node40688 = (inp[9]) ? node40694 : node40689;
														assign node40689 = (inp[15]) ? 4'b1101 : node40690;
															assign node40690 = (inp[0]) ? 4'b1101 : 4'b1111;
														assign node40694 = (inp[12]) ? node40702 : node40695;
															assign node40695 = (inp[0]) ? node40699 : node40696;
																assign node40696 = (inp[15]) ? 4'b1001 : 4'b1011;
																assign node40699 = (inp[15]) ? 4'b1011 : 4'b1001;
															assign node40702 = (inp[15]) ? node40706 : node40703;
																assign node40703 = (inp[0]) ? 4'b1001 : 4'b1011;
																assign node40706 = (inp[0]) ? 4'b1011 : 4'b1001;
												assign node40709 = (inp[12]) ? node40729 : node40710;
													assign node40710 = (inp[0]) ? node40722 : node40711;
														assign node40711 = (inp[15]) ? node40717 : node40712;
															assign node40712 = (inp[4]) ? node40714 : 4'b1101;
																assign node40714 = (inp[9]) ? 4'b1001 : 4'b1101;
															assign node40717 = (inp[9]) ? 4'b1111 : node40718;
																assign node40718 = (inp[4]) ? 4'b1111 : 4'b1001;
														assign node40722 = (inp[4]) ? node40726 : node40723;
															assign node40723 = (inp[15]) ? 4'b1011 : 4'b1111;
															assign node40726 = (inp[15]) ? 4'b1101 : 4'b1111;
													assign node40729 = (inp[9]) ? node40745 : node40730;
														assign node40730 = (inp[4]) ? node40738 : node40731;
															assign node40731 = (inp[15]) ? node40735 : node40732;
																assign node40732 = (inp[0]) ? 4'b1001 : 4'b1011;
																assign node40735 = (inp[0]) ? 4'b1011 : 4'b1001;
															assign node40738 = (inp[15]) ? node40742 : node40739;
																assign node40739 = (inp[0]) ? 4'b1111 : 4'b1101;
																assign node40742 = (inp[0]) ? 4'b1101 : 4'b1111;
														assign node40745 = (inp[4]) ? node40751 : node40746;
															assign node40746 = (inp[15]) ? node40748 : 4'b1111;
																assign node40748 = (inp[0]) ? 4'b1101 : 4'b1111;
															assign node40751 = (inp[15]) ? node40755 : node40752;
																assign node40752 = (inp[0]) ? 4'b1011 : 4'b1001;
																assign node40755 = (inp[0]) ? 4'b1001 : 4'b1011;
										assign node40758 = (inp[10]) ? node40834 : node40759;
											assign node40759 = (inp[0]) ? node40793 : node40760;
												assign node40760 = (inp[15]) ? node40780 : node40761;
													assign node40761 = (inp[4]) ? node40773 : node40762;
														assign node40762 = (inp[5]) ? node40768 : node40763;
															assign node40763 = (inp[9]) ? 4'b1011 : node40764;
																assign node40764 = (inp[12]) ? 4'b1011 : 4'b1111;
															assign node40768 = (inp[9]) ? node40770 : 4'b1101;
																assign node40770 = (inp[12]) ? 4'b1101 : 4'b1001;
														assign node40773 = (inp[9]) ? node40777 : node40774;
															assign node40774 = (inp[12]) ? 4'b1101 : 4'b1001;
															assign node40777 = (inp[12]) ? 4'b1001 : 4'b1101;
													assign node40780 = (inp[9]) ? node40786 : node40781;
														assign node40781 = (inp[4]) ? node40783 : 4'b1001;
															assign node40783 = (inp[12]) ? 4'b1111 : 4'b1001;
														assign node40786 = (inp[4]) ? node40790 : node40787;
															assign node40787 = (inp[12]) ? 4'b1111 : 4'b1011;
															assign node40790 = (inp[12]) ? 4'b1011 : 4'b1111;
												assign node40793 = (inp[15]) ? node40817 : node40794;
													assign node40794 = (inp[5]) ? node40804 : node40795;
														assign node40795 = (inp[9]) ? 4'b1111 : node40796;
															assign node40796 = (inp[12]) ? node40800 : node40797;
																assign node40797 = (inp[4]) ? 4'b1001 : 4'b1101;
																assign node40800 = (inp[4]) ? 4'b1111 : 4'b1001;
														assign node40804 = (inp[4]) ? node40810 : node40805;
															assign node40805 = (inp[12]) ? node40807 : 4'b1111;
																assign node40807 = (inp[9]) ? 4'b1111 : 4'b1011;
															assign node40810 = (inp[9]) ? node40814 : node40811;
																assign node40811 = (inp[12]) ? 4'b1111 : 4'b1011;
																assign node40814 = (inp[12]) ? 4'b1011 : 4'b1111;
													assign node40817 = (inp[9]) ? node40827 : node40818;
														assign node40818 = (inp[5]) ? node40822 : node40819;
															assign node40819 = (inp[12]) ? 4'b1011 : 4'b1111;
															assign node40822 = (inp[12]) ? node40824 : 4'b1101;
																assign node40824 = (inp[4]) ? 4'b1101 : 4'b1001;
														assign node40827 = (inp[4]) ? node40831 : node40828;
															assign node40828 = (inp[12]) ? 4'b1101 : 4'b1001;
															assign node40831 = (inp[12]) ? 4'b1001 : 4'b1101;
											assign node40834 = (inp[0]) ? node40854 : node40835;
												assign node40835 = (inp[15]) ? node40845 : node40836;
													assign node40836 = (inp[9]) ? node40842 : node40837;
														assign node40837 = (inp[4]) ? 4'b1101 : node40838;
															assign node40838 = (inp[5]) ? 4'b1001 : 4'b1011;
														assign node40842 = (inp[4]) ? 4'b1001 : 4'b1101;
													assign node40845 = (inp[9]) ? node40851 : node40846;
														assign node40846 = (inp[4]) ? 4'b1111 : node40847;
															assign node40847 = (inp[5]) ? 4'b1011 : 4'b1001;
														assign node40851 = (inp[4]) ? 4'b1011 : 4'b1111;
												assign node40854 = (inp[15]) ? node40864 : node40855;
													assign node40855 = (inp[4]) ? node40861 : node40856;
														assign node40856 = (inp[9]) ? 4'b1111 : node40857;
															assign node40857 = (inp[5]) ? 4'b1011 : 4'b1001;
														assign node40861 = (inp[9]) ? 4'b1011 : 4'b1111;
													assign node40864 = (inp[4]) ? node40870 : node40865;
														assign node40865 = (inp[9]) ? 4'b1101 : node40866;
															assign node40866 = (inp[5]) ? 4'b1001 : 4'b1011;
														assign node40870 = (inp[9]) ? 4'b1001 : 4'b1101;
									assign node40873 = (inp[5]) ? node41007 : node40874;
										assign node40874 = (inp[4]) ? node40932 : node40875;
											assign node40875 = (inp[9]) ? node40897 : node40876;
												assign node40876 = (inp[12]) ? node40890 : node40877;
													assign node40877 = (inp[10]) ? node40883 : node40878;
														assign node40878 = (inp[0]) ? 4'b1100 : node40879;
															assign node40879 = (inp[15]) ? 4'b1100 : 4'b1110;
														assign node40883 = (inp[15]) ? node40887 : node40884;
															assign node40884 = (inp[3]) ? 4'b1000 : 4'b1010;
															assign node40887 = (inp[0]) ? 4'b1010 : 4'b1000;
													assign node40890 = (inp[15]) ? node40894 : node40891;
														assign node40891 = (inp[0]) ? 4'b1000 : 4'b1010;
														assign node40894 = (inp[0]) ? 4'b1010 : 4'b1000;
												assign node40897 = (inp[10]) ? node40913 : node40898;
													assign node40898 = (inp[12]) ? node40906 : node40899;
														assign node40899 = (inp[15]) ? node40903 : node40900;
															assign node40900 = (inp[0]) ? 4'b1000 : 4'b1010;
															assign node40903 = (inp[0]) ? 4'b1010 : 4'b1000;
														assign node40906 = (inp[15]) ? node40908 : 4'b1100;
															assign node40908 = (inp[0]) ? 4'b1100 : node40909;
																assign node40909 = (inp[3]) ? 4'b1110 : 4'b1100;
													assign node40913 = (inp[0]) ? node40923 : node40914;
														assign node40914 = (inp[12]) ? node40916 : 4'b1100;
															assign node40916 = (inp[15]) ? node40920 : node40917;
																assign node40917 = (inp[3]) ? 4'b1100 : 4'b1110;
																assign node40920 = (inp[3]) ? 4'b1110 : 4'b1100;
														assign node40923 = (inp[12]) ? 4'b1100 : node40924;
															assign node40924 = (inp[3]) ? node40928 : node40925;
																assign node40925 = (inp[15]) ? 4'b1110 : 4'b1100;
																assign node40928 = (inp[15]) ? 4'b1100 : 4'b1110;
											assign node40932 = (inp[9]) ? node40978 : node40933;
												assign node40933 = (inp[12]) ? node40955 : node40934;
													assign node40934 = (inp[10]) ? node40944 : node40935;
														assign node40935 = (inp[3]) ? 4'b1000 : node40936;
															assign node40936 = (inp[15]) ? node40940 : node40937;
																assign node40937 = (inp[0]) ? 4'b1000 : 4'b1010;
																assign node40940 = (inp[0]) ? 4'b1010 : 4'b1000;
														assign node40944 = (inp[15]) ? node40950 : node40945;
															assign node40945 = (inp[3]) ? node40947 : 4'b1110;
																assign node40947 = (inp[0]) ? 4'b1110 : 4'b1100;
															assign node40950 = (inp[3]) ? node40952 : 4'b1100;
																assign node40952 = (inp[0]) ? 4'b1100 : 4'b1110;
													assign node40955 = (inp[10]) ? node40969 : node40956;
														assign node40956 = (inp[15]) ? node40962 : node40957;
															assign node40957 = (inp[3]) ? node40959 : 4'b1110;
																assign node40959 = (inp[0]) ? 4'b1110 : 4'b1100;
															assign node40962 = (inp[0]) ? node40966 : node40963;
																assign node40963 = (inp[3]) ? 4'b1110 : 4'b1100;
																assign node40966 = (inp[3]) ? 4'b1100 : 4'b1110;
														assign node40969 = (inp[3]) ? 4'b1100 : node40970;
															assign node40970 = (inp[15]) ? node40974 : node40971;
																assign node40971 = (inp[0]) ? 4'b1100 : 4'b1110;
																assign node40974 = (inp[0]) ? 4'b1110 : 4'b1100;
												assign node40978 = (inp[12]) ? node40998 : node40979;
													assign node40979 = (inp[10]) ? node40991 : node40980;
														assign node40980 = (inp[0]) ? node40986 : node40981;
															assign node40981 = (inp[15]) ? node40983 : 4'b1100;
																assign node40983 = (inp[3]) ? 4'b1110 : 4'b1100;
															assign node40986 = (inp[3]) ? 4'b1110 : node40987;
																assign node40987 = (inp[15]) ? 4'b1110 : 4'b1100;
														assign node40991 = (inp[15]) ? 4'b1000 : node40992;
															assign node40992 = (inp[3]) ? node40994 : 4'b1000;
																assign node40994 = (inp[0]) ? 4'b1010 : 4'b1000;
													assign node40998 = (inp[3]) ? 4'b1010 : node40999;
														assign node40999 = (inp[15]) ? node41003 : node41000;
															assign node41000 = (inp[0]) ? 4'b1000 : 4'b1010;
															assign node41003 = (inp[0]) ? 4'b1010 : 4'b1000;
										assign node41007 = (inp[3]) ? node41089 : node41008;
											assign node41008 = (inp[4]) ? node41044 : node41009;
												assign node41009 = (inp[9]) ? node41029 : node41010;
													assign node41010 = (inp[10]) ? node41022 : node41011;
														assign node41011 = (inp[12]) ? node41017 : node41012;
															assign node41012 = (inp[0]) ? 4'b1110 : node41013;
																assign node41013 = (inp[15]) ? 4'b1100 : 4'b1110;
															assign node41017 = (inp[0]) ? node41019 : 4'b1010;
																assign node41019 = (inp[15]) ? 4'b1010 : 4'b1000;
														assign node41022 = (inp[15]) ? node41026 : node41023;
															assign node41023 = (inp[0]) ? 4'b1000 : 4'b1010;
															assign node41026 = (inp[0]) ? 4'b1010 : 4'b1000;
													assign node41029 = (inp[10]) ? node41037 : node41030;
														assign node41030 = (inp[12]) ? 4'b1110 : node41031;
															assign node41031 = (inp[0]) ? 4'b1000 : node41032;
																assign node41032 = (inp[15]) ? 4'b1000 : 4'b1010;
														assign node41037 = (inp[0]) ? node41041 : node41038;
															assign node41038 = (inp[15]) ? 4'b1110 : 4'b1100;
															assign node41041 = (inp[15]) ? 4'b1100 : 4'b1110;
												assign node41044 = (inp[9]) ? node41066 : node41045;
													assign node41045 = (inp[10]) ? node41059 : node41046;
														assign node41046 = (inp[12]) ? node41054 : node41047;
															assign node41047 = (inp[0]) ? node41051 : node41048;
																assign node41048 = (inp[15]) ? 4'b1000 : 4'b1010;
																assign node41051 = (inp[15]) ? 4'b1010 : 4'b1000;
															assign node41054 = (inp[0]) ? 4'b1100 : node41055;
																assign node41055 = (inp[15]) ? 4'b1110 : 4'b1100;
														assign node41059 = (inp[0]) ? node41063 : node41060;
															assign node41060 = (inp[15]) ? 4'b1110 : 4'b1100;
															assign node41063 = (inp[15]) ? 4'b1100 : 4'b1110;
													assign node41066 = (inp[10]) ? node41082 : node41067;
														assign node41067 = (inp[12]) ? node41075 : node41068;
															assign node41068 = (inp[15]) ? node41072 : node41069;
																assign node41069 = (inp[0]) ? 4'b1110 : 4'b1100;
																assign node41072 = (inp[0]) ? 4'b1100 : 4'b1110;
															assign node41075 = (inp[15]) ? node41079 : node41076;
																assign node41076 = (inp[0]) ? 4'b1010 : 4'b1000;
																assign node41079 = (inp[0]) ? 4'b1000 : 4'b1010;
														assign node41082 = (inp[15]) ? node41086 : node41083;
															assign node41083 = (inp[0]) ? 4'b1010 : 4'b1000;
															assign node41086 = (inp[0]) ? 4'b1000 : 4'b1010;
											assign node41089 = (inp[10]) ? node41123 : node41090;
												assign node41090 = (inp[15]) ? node41110 : node41091;
													assign node41091 = (inp[0]) ? node41097 : node41092;
														assign node41092 = (inp[12]) ? node41094 : 4'b1000;
															assign node41094 = (inp[9]) ? 4'b1100 : 4'b1000;
														assign node41097 = (inp[9]) ? node41105 : node41098;
															assign node41098 = (inp[12]) ? node41102 : node41099;
																assign node41099 = (inp[4]) ? 4'b1010 : 4'b1110;
																assign node41102 = (inp[4]) ? 4'b1110 : 4'b1010;
															assign node41105 = (inp[12]) ? node41107 : 4'b1010;
																assign node41107 = (inp[4]) ? 4'b1010 : 4'b1110;
													assign node41110 = (inp[0]) ? 4'b1100 : node41111;
														assign node41111 = (inp[9]) ? node41117 : node41112;
															assign node41112 = (inp[12]) ? node41114 : 4'b1110;
																assign node41114 = (inp[4]) ? 4'b1110 : 4'b1010;
															assign node41117 = (inp[12]) ? node41119 : 4'b1010;
																assign node41119 = (inp[4]) ? 4'b1010 : 4'b1110;
												assign node41123 = (inp[15]) ? node41137 : node41124;
													assign node41124 = (inp[0]) ? node41130 : node41125;
														assign node41125 = (inp[9]) ? 4'b1100 : node41126;
															assign node41126 = (inp[4]) ? 4'b1100 : 4'b1000;
														assign node41130 = (inp[9]) ? node41134 : node41131;
															assign node41131 = (inp[4]) ? 4'b1110 : 4'b1010;
															assign node41134 = (inp[4]) ? 4'b1010 : 4'b1110;
													assign node41137 = (inp[0]) ? node41141 : node41138;
														assign node41138 = (inp[4]) ? 4'b1010 : 4'b1110;
														assign node41141 = (inp[12]) ? node41145 : node41142;
															assign node41142 = (inp[4]) ? 4'b1000 : 4'b1100;
															assign node41145 = (inp[9]) ? 4'b1000 : node41146;
																assign node41146 = (inp[4]) ? 4'b1100 : 4'b1000;
								assign node41150 = (inp[9]) ? node41354 : node41151;
									assign node41151 = (inp[4]) ? node41229 : node41152;
										assign node41152 = (inp[10]) ? node41206 : node41153;
											assign node41153 = (inp[12]) ? node41187 : node41154;
												assign node41154 = (inp[14]) ? node41172 : node41155;
													assign node41155 = (inp[15]) ? node41163 : node41156;
														assign node41156 = (inp[0]) ? 4'b1100 : node41157;
															assign node41157 = (inp[3]) ? node41159 : 4'b1110;
																assign node41159 = (inp[5]) ? 4'b1100 : 4'b1110;
														assign node41163 = (inp[0]) ? node41167 : node41164;
															assign node41164 = (inp[5]) ? 4'b1110 : 4'b1100;
															assign node41167 = (inp[3]) ? node41169 : 4'b1110;
																assign node41169 = (inp[5]) ? 4'b1100 : 4'b1110;
													assign node41172 = (inp[5]) ? node41180 : node41173;
														assign node41173 = (inp[15]) ? node41177 : node41174;
															assign node41174 = (inp[0]) ? 4'b1100 : 4'b1110;
															assign node41177 = (inp[0]) ? 4'b1110 : 4'b1100;
														assign node41180 = (inp[15]) ? 4'b1100 : node41181;
															assign node41181 = (inp[0]) ? node41183 : 4'b1100;
																assign node41183 = (inp[3]) ? 4'b1110 : 4'b1100;
												assign node41187 = (inp[0]) ? node41197 : node41188;
													assign node41188 = (inp[3]) ? node41190 : 4'b1010;
														assign node41190 = (inp[15]) ? node41194 : node41191;
															assign node41191 = (inp[5]) ? 4'b1000 : 4'b1010;
															assign node41194 = (inp[5]) ? 4'b1010 : 4'b1000;
													assign node41197 = (inp[15]) ? node41203 : node41198;
														assign node41198 = (inp[5]) ? node41200 : 4'b1000;
															assign node41200 = (inp[3]) ? 4'b1010 : 4'b1000;
														assign node41203 = (inp[5]) ? 4'b1000 : 4'b1010;
											assign node41206 = (inp[5]) ? node41214 : node41207;
												assign node41207 = (inp[15]) ? node41211 : node41208;
													assign node41208 = (inp[0]) ? 4'b1000 : 4'b1010;
													assign node41211 = (inp[0]) ? 4'b1010 : 4'b1000;
												assign node41214 = (inp[3]) ? node41222 : node41215;
													assign node41215 = (inp[15]) ? node41219 : node41216;
														assign node41216 = (inp[0]) ? 4'b1000 : 4'b1010;
														assign node41219 = (inp[0]) ? 4'b1010 : 4'b1000;
													assign node41222 = (inp[0]) ? node41226 : node41223;
														assign node41223 = (inp[15]) ? 4'b1010 : 4'b1000;
														assign node41226 = (inp[15]) ? 4'b1000 : 4'b1010;
										assign node41229 = (inp[10]) ? node41281 : node41230;
											assign node41230 = (inp[12]) ? node41252 : node41231;
												assign node41231 = (inp[0]) ? node41241 : node41232;
													assign node41232 = (inp[15]) ? node41236 : node41233;
														assign node41233 = (inp[5]) ? 4'b1000 : 4'b1010;
														assign node41236 = (inp[3]) ? node41238 : 4'b1000;
															assign node41238 = (inp[5]) ? 4'b1010 : 4'b1000;
													assign node41241 = (inp[15]) ? node41247 : node41242;
														assign node41242 = (inp[3]) ? node41244 : 4'b1000;
															assign node41244 = (inp[5]) ? 4'b1010 : 4'b1000;
														assign node41247 = (inp[3]) ? node41249 : 4'b1010;
															assign node41249 = (inp[5]) ? 4'b1000 : 4'b1010;
												assign node41252 = (inp[3]) ? node41268 : node41253;
													assign node41253 = (inp[14]) ? node41261 : node41254;
														assign node41254 = (inp[5]) ? node41256 : 4'b1110;
															assign node41256 = (inp[15]) ? node41258 : 4'b1100;
																assign node41258 = (inp[0]) ? 4'b1100 : 4'b1110;
														assign node41261 = (inp[5]) ? 4'b1110 : node41262;
															assign node41262 = (inp[0]) ? 4'b1110 : node41263;
																assign node41263 = (inp[15]) ? 4'b1100 : 4'b1110;
													assign node41268 = (inp[5]) ? node41276 : node41269;
														assign node41269 = (inp[15]) ? node41273 : node41270;
															assign node41270 = (inp[0]) ? 4'b1110 : 4'b1100;
															assign node41273 = (inp[0]) ? 4'b1100 : 4'b1110;
														assign node41276 = (inp[0]) ? node41278 : 4'b1110;
															assign node41278 = (inp[15]) ? 4'b1100 : 4'b1110;
											assign node41281 = (inp[3]) ? node41319 : node41282;
												assign node41282 = (inp[14]) ? node41304 : node41283;
													assign node41283 = (inp[15]) ? node41291 : node41284;
														assign node41284 = (inp[5]) ? node41288 : node41285;
															assign node41285 = (inp[0]) ? 4'b1100 : 4'b1110;
															assign node41288 = (inp[0]) ? 4'b1110 : 4'b1100;
														assign node41291 = (inp[12]) ? node41299 : node41292;
															assign node41292 = (inp[0]) ? node41296 : node41293;
																assign node41293 = (inp[5]) ? 4'b1110 : 4'b1100;
																assign node41296 = (inp[5]) ? 4'b1100 : 4'b1110;
															assign node41299 = (inp[0]) ? node41301 : 4'b1100;
																assign node41301 = (inp[5]) ? 4'b1100 : 4'b1110;
													assign node41304 = (inp[0]) ? node41310 : node41305;
														assign node41305 = (inp[15]) ? 4'b1110 : node41306;
															assign node41306 = (inp[5]) ? 4'b1100 : 4'b1110;
														assign node41310 = (inp[12]) ? node41312 : 4'b1110;
															assign node41312 = (inp[5]) ? node41316 : node41313;
																assign node41313 = (inp[15]) ? 4'b1110 : 4'b1100;
																assign node41316 = (inp[15]) ? 4'b1100 : 4'b1110;
												assign node41319 = (inp[5]) ? node41335 : node41320;
													assign node41320 = (inp[14]) ? node41328 : node41321;
														assign node41321 = (inp[15]) ? node41325 : node41322;
															assign node41322 = (inp[0]) ? 4'b1110 : 4'b1100;
															assign node41325 = (inp[0]) ? 4'b1100 : 4'b1110;
														assign node41328 = (inp[0]) ? node41332 : node41329;
															assign node41329 = (inp[15]) ? 4'b1110 : 4'b1100;
															assign node41332 = (inp[15]) ? 4'b1100 : 4'b1110;
													assign node41335 = (inp[14]) ? node41343 : node41336;
														assign node41336 = (inp[0]) ? node41340 : node41337;
															assign node41337 = (inp[15]) ? 4'b1110 : 4'b1100;
															assign node41340 = (inp[15]) ? 4'b1100 : 4'b1110;
														assign node41343 = (inp[12]) ? node41349 : node41344;
															assign node41344 = (inp[15]) ? node41346 : 4'b1100;
																assign node41346 = (inp[0]) ? 4'b1100 : 4'b1110;
															assign node41349 = (inp[0]) ? node41351 : 4'b1100;
																assign node41351 = (inp[15]) ? 4'b1100 : 4'b1110;
									assign node41354 = (inp[4]) ? node41456 : node41355;
										assign node41355 = (inp[10]) ? node41397 : node41356;
											assign node41356 = (inp[12]) ? node41380 : node41357;
												assign node41357 = (inp[0]) ? node41369 : node41358;
													assign node41358 = (inp[15]) ? node41364 : node41359;
														assign node41359 = (inp[5]) ? node41361 : 4'b1010;
															assign node41361 = (inp[3]) ? 4'b1000 : 4'b1010;
														assign node41364 = (inp[5]) ? node41366 : 4'b1000;
															assign node41366 = (inp[3]) ? 4'b1010 : 4'b1000;
													assign node41369 = (inp[15]) ? node41375 : node41370;
														assign node41370 = (inp[3]) ? node41372 : 4'b1000;
															assign node41372 = (inp[5]) ? 4'b1010 : 4'b1000;
														assign node41375 = (inp[3]) ? node41377 : 4'b1010;
															assign node41377 = (inp[5]) ? 4'b1000 : 4'b1010;
												assign node41380 = (inp[15]) ? node41390 : node41381;
													assign node41381 = (inp[0]) ? node41385 : node41382;
														assign node41382 = (inp[3]) ? 4'b1100 : 4'b1110;
														assign node41385 = (inp[3]) ? 4'b1110 : node41386;
															assign node41386 = (inp[5]) ? 4'b1110 : 4'b1100;
													assign node41390 = (inp[0]) ? 4'b1100 : node41391;
														assign node41391 = (inp[5]) ? 4'b1110 : node41392;
															assign node41392 = (inp[3]) ? 4'b1110 : 4'b1100;
											assign node41397 = (inp[3]) ? node41441 : node41398;
												assign node41398 = (inp[14]) ? node41422 : node41399;
													assign node41399 = (inp[12]) ? node41413 : node41400;
														assign node41400 = (inp[15]) ? node41408 : node41401;
															assign node41401 = (inp[5]) ? node41405 : node41402;
																assign node41402 = (inp[0]) ? 4'b1100 : 4'b1110;
																assign node41405 = (inp[0]) ? 4'b1110 : 4'b1100;
															assign node41408 = (inp[0]) ? 4'b1110 : node41409;
																assign node41409 = (inp[5]) ? 4'b1110 : 4'b1100;
														assign node41413 = (inp[5]) ? node41415 : 4'b1110;
															assign node41415 = (inp[15]) ? node41419 : node41416;
																assign node41416 = (inp[0]) ? 4'b1110 : 4'b1100;
																assign node41419 = (inp[0]) ? 4'b1100 : 4'b1110;
													assign node41422 = (inp[12]) ? node41432 : node41423;
														assign node41423 = (inp[5]) ? 4'b1110 : node41424;
															assign node41424 = (inp[0]) ? node41428 : node41425;
																assign node41425 = (inp[15]) ? 4'b1100 : 4'b1110;
																assign node41428 = (inp[15]) ? 4'b1110 : 4'b1100;
														assign node41432 = (inp[5]) ? 4'b1100 : node41433;
															assign node41433 = (inp[15]) ? node41437 : node41434;
																assign node41434 = (inp[0]) ? 4'b1100 : 4'b1110;
																assign node41437 = (inp[0]) ? 4'b1110 : 4'b1100;
												assign node41441 = (inp[12]) ? node41449 : node41442;
													assign node41442 = (inp[0]) ? node41446 : node41443;
														assign node41443 = (inp[15]) ? 4'b1110 : 4'b1100;
														assign node41446 = (inp[15]) ? 4'b1100 : 4'b1110;
													assign node41449 = (inp[0]) ? node41453 : node41450;
														assign node41450 = (inp[15]) ? 4'b1110 : 4'b1100;
														assign node41453 = (inp[15]) ? 4'b1100 : 4'b1110;
										assign node41456 = (inp[10]) ? node41516 : node41457;
											assign node41457 = (inp[12]) ? node41493 : node41458;
												assign node41458 = (inp[14]) ? node41468 : node41459;
													assign node41459 = (inp[3]) ? 4'b1110 : node41460;
														assign node41460 = (inp[5]) ? node41464 : node41461;
															assign node41461 = (inp[0]) ? 4'b1110 : 4'b1100;
															assign node41464 = (inp[0]) ? 4'b1100 : 4'b1110;
													assign node41468 = (inp[5]) ? node41478 : node41469;
														assign node41469 = (inp[3]) ? 4'b1100 : node41470;
															assign node41470 = (inp[15]) ? node41474 : node41471;
																assign node41471 = (inp[0]) ? 4'b1100 : 4'b1110;
																assign node41474 = (inp[0]) ? 4'b1110 : 4'b1100;
														assign node41478 = (inp[3]) ? node41486 : node41479;
															assign node41479 = (inp[0]) ? node41483 : node41480;
																assign node41480 = (inp[15]) ? 4'b1110 : 4'b1100;
																assign node41483 = (inp[15]) ? 4'b1100 : 4'b1110;
															assign node41486 = (inp[0]) ? node41490 : node41487;
																assign node41487 = (inp[15]) ? 4'b1110 : 4'b1100;
																assign node41490 = (inp[15]) ? 4'b1100 : 4'b1110;
												assign node41493 = (inp[0]) ? node41505 : node41494;
													assign node41494 = (inp[15]) ? node41500 : node41495;
														assign node41495 = (inp[5]) ? 4'b1000 : node41496;
															assign node41496 = (inp[3]) ? 4'b1000 : 4'b1010;
														assign node41500 = (inp[5]) ? 4'b1010 : node41501;
															assign node41501 = (inp[3]) ? 4'b1010 : 4'b1000;
													assign node41505 = (inp[15]) ? node41511 : node41506;
														assign node41506 = (inp[14]) ? 4'b1010 : node41507;
															assign node41507 = (inp[5]) ? 4'b1010 : 4'b1000;
														assign node41511 = (inp[3]) ? 4'b1000 : node41512;
															assign node41512 = (inp[5]) ? 4'b1000 : 4'b1010;
											assign node41516 = (inp[0]) ? node41528 : node41517;
												assign node41517 = (inp[15]) ? node41523 : node41518;
													assign node41518 = (inp[3]) ? 4'b1000 : node41519;
														assign node41519 = (inp[5]) ? 4'b1000 : 4'b1010;
													assign node41523 = (inp[3]) ? 4'b1010 : node41524;
														assign node41524 = (inp[5]) ? 4'b1010 : 4'b1000;
												assign node41528 = (inp[15]) ? node41534 : node41529;
													assign node41529 = (inp[5]) ? 4'b1010 : node41530;
														assign node41530 = (inp[3]) ? 4'b1010 : 4'b1000;
													assign node41534 = (inp[5]) ? 4'b1000 : node41535;
														assign node41535 = (inp[3]) ? 4'b1000 : 4'b1010;
				assign node41539 = (inp[1]) ? node45539 : node41540;
					assign node41540 = (inp[8]) ? node43602 : node41541;
						assign node41541 = (inp[7]) ? node42555 : node41542;
							assign node41542 = (inp[2]) ? node42156 : node41543;
								assign node41543 = (inp[14]) ? node41805 : node41544;
									assign node41544 = (inp[3]) ? node41662 : node41545;
										assign node41545 = (inp[0]) ? node41599 : node41546;
											assign node41546 = (inp[15]) ? node41574 : node41547;
												assign node41547 = (inp[5]) ? node41565 : node41548;
													assign node41548 = (inp[10]) ? node41556 : node41549;
														assign node41549 = (inp[4]) ? node41553 : node41550;
															assign node41550 = (inp[9]) ? 4'b0011 : 4'b0111;
															assign node41553 = (inp[9]) ? 4'b0111 : 4'b0011;
														assign node41556 = (inp[12]) ? node41558 : 4'b0111;
															assign node41558 = (inp[4]) ? node41562 : node41559;
																assign node41559 = (inp[9]) ? 4'b0111 : 4'b0011;
																assign node41562 = (inp[9]) ? 4'b0011 : 4'b0111;
													assign node41565 = (inp[9]) ? node41569 : node41566;
														assign node41566 = (inp[4]) ? 4'b0011 : 4'b0111;
														assign node41569 = (inp[4]) ? 4'b0101 : node41570;
															assign node41570 = (inp[12]) ? 4'b0101 : 4'b0011;
												assign node41574 = (inp[5]) ? node41588 : node41575;
													assign node41575 = (inp[9]) ? node41579 : node41576;
														assign node41576 = (inp[4]) ? 4'b0001 : 4'b0101;
														assign node41579 = (inp[4]) ? node41583 : node41580;
															assign node41580 = (inp[10]) ? 4'b0101 : 4'b0001;
															assign node41583 = (inp[10]) ? node41585 : 4'b0101;
																assign node41585 = (inp[12]) ? 4'b0001 : 4'b0101;
													assign node41588 = (inp[4]) ? node41596 : node41589;
														assign node41589 = (inp[9]) ? 4'b0001 : node41590;
															assign node41590 = (inp[10]) ? node41592 : 4'b0101;
																assign node41592 = (inp[12]) ? 4'b0001 : 4'b0101;
														assign node41596 = (inp[9]) ? 4'b0111 : 4'b0001;
											assign node41599 = (inp[15]) ? node41631 : node41600;
												assign node41600 = (inp[9]) ? node41614 : node41601;
													assign node41601 = (inp[4]) ? node41607 : node41602;
														assign node41602 = (inp[12]) ? node41604 : 4'b0101;
															assign node41604 = (inp[10]) ? 4'b0001 : 4'b0101;
														assign node41607 = (inp[5]) ? 4'b0001 : node41608;
															assign node41608 = (inp[12]) ? node41610 : 4'b0001;
																assign node41610 = (inp[10]) ? 4'b0101 : 4'b0001;
													assign node41614 = (inp[5]) ? node41624 : node41615;
														assign node41615 = (inp[4]) ? node41621 : node41616;
															assign node41616 = (inp[12]) ? node41618 : 4'b0001;
																assign node41618 = (inp[10]) ? 4'b0101 : 4'b0001;
															assign node41621 = (inp[10]) ? 4'b0001 : 4'b0101;
														assign node41624 = (inp[12]) ? node41626 : 4'b0001;
															assign node41626 = (inp[10]) ? node41628 : 4'b0111;
																assign node41628 = (inp[4]) ? 4'b0011 : 4'b0111;
												assign node41631 = (inp[5]) ? node41649 : node41632;
													assign node41632 = (inp[9]) ? node41644 : node41633;
														assign node41633 = (inp[4]) ? node41639 : node41634;
															assign node41634 = (inp[10]) ? node41636 : 4'b0111;
																assign node41636 = (inp[12]) ? 4'b0011 : 4'b0111;
															assign node41639 = (inp[12]) ? node41641 : 4'b0011;
																assign node41641 = (inp[10]) ? 4'b0111 : 4'b0011;
														assign node41644 = (inp[4]) ? 4'b0111 : node41645;
															assign node41645 = (inp[10]) ? 4'b0111 : 4'b0011;
													assign node41649 = (inp[9]) ? node41655 : node41650;
														assign node41650 = (inp[4]) ? 4'b0011 : node41651;
															assign node41651 = (inp[10]) ? 4'b0011 : 4'b0111;
														assign node41655 = (inp[4]) ? node41657 : 4'b0011;
															assign node41657 = (inp[10]) ? node41659 : 4'b0101;
																assign node41659 = (inp[12]) ? 4'b0001 : 4'b0101;
										assign node41662 = (inp[12]) ? node41730 : node41663;
											assign node41663 = (inp[4]) ? node41695 : node41664;
												assign node41664 = (inp[9]) ? node41686 : node41665;
													assign node41665 = (inp[10]) ? node41673 : node41666;
														assign node41666 = (inp[15]) ? 4'b0111 : node41667;
															assign node41667 = (inp[5]) ? 4'b0111 : node41668;
																assign node41668 = (inp[0]) ? 4'b0101 : 4'b0111;
														assign node41673 = (inp[15]) ? node41679 : node41674;
															assign node41674 = (inp[5]) ? 4'b0111 : node41675;
																assign node41675 = (inp[0]) ? 4'b0101 : 4'b0111;
															assign node41679 = (inp[5]) ? node41683 : node41680;
																assign node41680 = (inp[0]) ? 4'b0111 : 4'b0101;
																assign node41683 = (inp[0]) ? 4'b0101 : 4'b0111;
													assign node41686 = (inp[5]) ? 4'b0011 : node41687;
														assign node41687 = (inp[15]) ? node41691 : node41688;
															assign node41688 = (inp[0]) ? 4'b0001 : 4'b0011;
															assign node41691 = (inp[0]) ? 4'b0011 : 4'b0001;
												assign node41695 = (inp[9]) ? node41719 : node41696;
													assign node41696 = (inp[0]) ? node41704 : node41697;
														assign node41697 = (inp[15]) ? node41701 : node41698;
															assign node41698 = (inp[5]) ? 4'b0001 : 4'b0011;
															assign node41701 = (inp[5]) ? 4'b0011 : 4'b0001;
														assign node41704 = (inp[10]) ? node41712 : node41705;
															assign node41705 = (inp[5]) ? node41709 : node41706;
																assign node41706 = (inp[15]) ? 4'b0011 : 4'b0001;
																assign node41709 = (inp[15]) ? 4'b0001 : 4'b0011;
															assign node41712 = (inp[5]) ? node41716 : node41713;
																assign node41713 = (inp[15]) ? 4'b0011 : 4'b0001;
																assign node41716 = (inp[15]) ? 4'b0001 : 4'b0011;
													assign node41719 = (inp[10]) ? node41725 : node41720;
														assign node41720 = (inp[0]) ? node41722 : 4'b0101;
															assign node41722 = (inp[15]) ? 4'b0101 : 4'b0111;
														assign node41725 = (inp[15]) ? node41727 : 4'b0111;
															assign node41727 = (inp[0]) ? 4'b0101 : 4'b0111;
											assign node41730 = (inp[9]) ? node41772 : node41731;
												assign node41731 = (inp[5]) ? node41755 : node41732;
													assign node41732 = (inp[0]) ? node41742 : node41733;
														assign node41733 = (inp[15]) ? node41739 : node41734;
															assign node41734 = (inp[4]) ? 4'b0101 : node41735;
																assign node41735 = (inp[10]) ? 4'b0011 : 4'b0111;
															assign node41739 = (inp[4]) ? 4'b0111 : 4'b0101;
														assign node41742 = (inp[15]) ? node41750 : node41743;
															assign node41743 = (inp[4]) ? node41747 : node41744;
																assign node41744 = (inp[10]) ? 4'b0001 : 4'b0101;
																assign node41747 = (inp[10]) ? 4'b0111 : 4'b0001;
															assign node41750 = (inp[10]) ? 4'b0101 : node41751;
																assign node41751 = (inp[4]) ? 4'b0011 : 4'b0111;
													assign node41755 = (inp[10]) ? node41765 : node41756;
														assign node41756 = (inp[4]) ? 4'b0011 : node41757;
															assign node41757 = (inp[15]) ? node41761 : node41758;
																assign node41758 = (inp[0]) ? 4'b0111 : 4'b0101;
																assign node41761 = (inp[0]) ? 4'b0101 : 4'b0111;
														assign node41765 = (inp[4]) ? node41767 : 4'b0011;
															assign node41767 = (inp[15]) ? 4'b0111 : node41768;
																assign node41768 = (inp[0]) ? 4'b0111 : 4'b0101;
												assign node41772 = (inp[4]) ? node41792 : node41773;
													assign node41773 = (inp[10]) ? node41787 : node41774;
														assign node41774 = (inp[5]) ? node41782 : node41775;
															assign node41775 = (inp[15]) ? node41779 : node41776;
																assign node41776 = (inp[0]) ? 4'b0001 : 4'b0011;
																assign node41779 = (inp[0]) ? 4'b0011 : 4'b0001;
															assign node41782 = (inp[15]) ? node41784 : 4'b0001;
																assign node41784 = (inp[0]) ? 4'b0001 : 4'b0011;
														assign node41787 = (inp[5]) ? node41789 : 4'b0101;
															assign node41789 = (inp[15]) ? 4'b0101 : 4'b0111;
													assign node41792 = (inp[10]) ? node41800 : node41793;
														assign node41793 = (inp[15]) ? node41797 : node41794;
															assign node41794 = (inp[0]) ? 4'b0111 : 4'b0101;
															assign node41797 = (inp[0]) ? 4'b0101 : 4'b0111;
														assign node41800 = (inp[0]) ? node41802 : 4'b0001;
															assign node41802 = (inp[15]) ? 4'b0001 : 4'b0011;
									assign node41805 = (inp[5]) ? node41995 : node41806;
										assign node41806 = (inp[3]) ? node41908 : node41807;
											assign node41807 = (inp[12]) ? node41857 : node41808;
												assign node41808 = (inp[10]) ? node41832 : node41809;
													assign node41809 = (inp[9]) ? node41821 : node41810;
														assign node41810 = (inp[4]) ? node41814 : node41811;
															assign node41811 = (inp[15]) ? 4'b0100 : 4'b0110;
															assign node41814 = (inp[15]) ? node41818 : node41815;
																assign node41815 = (inp[0]) ? 4'b0000 : 4'b0010;
																assign node41818 = (inp[0]) ? 4'b0010 : 4'b0000;
														assign node41821 = (inp[4]) ? node41827 : node41822;
															assign node41822 = (inp[0]) ? 4'b0010 : node41823;
																assign node41823 = (inp[15]) ? 4'b0000 : 4'b0010;
															assign node41827 = (inp[0]) ? node41829 : 4'b0110;
																assign node41829 = (inp[15]) ? 4'b0110 : 4'b0100;
													assign node41832 = (inp[9]) ? node41846 : node41833;
														assign node41833 = (inp[4]) ? node41841 : node41834;
															assign node41834 = (inp[15]) ? node41838 : node41835;
																assign node41835 = (inp[0]) ? 4'b0100 : 4'b0110;
																assign node41838 = (inp[0]) ? 4'b0110 : 4'b0100;
															assign node41841 = (inp[15]) ? 4'b0010 : node41842;
																assign node41842 = (inp[0]) ? 4'b0000 : 4'b0010;
														assign node41846 = (inp[4]) ? node41852 : node41847;
															assign node41847 = (inp[0]) ? 4'b0000 : node41848;
																assign node41848 = (inp[15]) ? 4'b0000 : 4'b0010;
															assign node41852 = (inp[0]) ? node41854 : 4'b0100;
																assign node41854 = (inp[15]) ? 4'b0110 : 4'b0100;
												assign node41857 = (inp[9]) ? node41881 : node41858;
													assign node41858 = (inp[4]) ? node41872 : node41859;
														assign node41859 = (inp[10]) ? node41867 : node41860;
															assign node41860 = (inp[15]) ? node41864 : node41861;
																assign node41861 = (inp[0]) ? 4'b0100 : 4'b0110;
																assign node41864 = (inp[0]) ? 4'b0110 : 4'b0100;
															assign node41867 = (inp[0]) ? 4'b0010 : node41868;
																assign node41868 = (inp[15]) ? 4'b0000 : 4'b0010;
														assign node41872 = (inp[10]) ? node41874 : 4'b0000;
															assign node41874 = (inp[0]) ? node41878 : node41875;
																assign node41875 = (inp[15]) ? 4'b0100 : 4'b0110;
																assign node41878 = (inp[15]) ? 4'b0110 : 4'b0100;
													assign node41881 = (inp[0]) ? node41893 : node41882;
														assign node41882 = (inp[15]) ? node41890 : node41883;
															assign node41883 = (inp[4]) ? node41887 : node41884;
																assign node41884 = (inp[10]) ? 4'b0110 : 4'b0010;
																assign node41887 = (inp[10]) ? 4'b0010 : 4'b0110;
															assign node41890 = (inp[4]) ? 4'b0000 : 4'b0100;
														assign node41893 = (inp[15]) ? node41901 : node41894;
															assign node41894 = (inp[10]) ? node41898 : node41895;
																assign node41895 = (inp[4]) ? 4'b0100 : 4'b0000;
																assign node41898 = (inp[4]) ? 4'b0000 : 4'b0100;
															assign node41901 = (inp[10]) ? node41905 : node41902;
																assign node41902 = (inp[4]) ? 4'b0110 : 4'b0010;
																assign node41905 = (inp[4]) ? 4'b0010 : 4'b0110;
											assign node41908 = (inp[12]) ? node41956 : node41909;
												assign node41909 = (inp[10]) ? node41929 : node41910;
													assign node41910 = (inp[9]) ? node41920 : node41911;
														assign node41911 = (inp[4]) ? 4'b0000 : node41912;
															assign node41912 = (inp[0]) ? node41916 : node41913;
																assign node41913 = (inp[15]) ? 4'b0100 : 4'b0110;
																assign node41916 = (inp[15]) ? 4'b0110 : 4'b0100;
														assign node41920 = (inp[4]) ? node41922 : 4'b0000;
															assign node41922 = (inp[0]) ? node41926 : node41923;
																assign node41923 = (inp[15]) ? 4'b0110 : 4'b0100;
																assign node41926 = (inp[15]) ? 4'b0100 : 4'b0110;
													assign node41929 = (inp[15]) ? node41941 : node41930;
														assign node41930 = (inp[4]) ? node41938 : node41931;
															assign node41931 = (inp[9]) ? node41935 : node41932;
																assign node41932 = (inp[0]) ? 4'b0100 : 4'b0110;
																assign node41935 = (inp[0]) ? 4'b0000 : 4'b0010;
															assign node41938 = (inp[0]) ? 4'b0110 : 4'b0100;
														assign node41941 = (inp[0]) ? node41949 : node41942;
															assign node41942 = (inp[9]) ? node41946 : node41943;
																assign node41943 = (inp[4]) ? 4'b0000 : 4'b0100;
																assign node41946 = (inp[4]) ? 4'b0110 : 4'b0000;
															assign node41949 = (inp[9]) ? node41953 : node41950;
																assign node41950 = (inp[4]) ? 4'b0010 : 4'b0110;
																assign node41953 = (inp[4]) ? 4'b0100 : 4'b0010;
												assign node41956 = (inp[4]) ? node41972 : node41957;
													assign node41957 = (inp[9]) ? node41963 : node41958;
														assign node41958 = (inp[10]) ? 4'b0000 : node41959;
															assign node41959 = (inp[0]) ? 4'b0110 : 4'b0100;
														assign node41963 = (inp[10]) ? node41965 : 4'b0000;
															assign node41965 = (inp[0]) ? node41969 : node41966;
																assign node41966 = (inp[15]) ? 4'b0110 : 4'b0100;
																assign node41969 = (inp[15]) ? 4'b0100 : 4'b0110;
													assign node41972 = (inp[15]) ? node41988 : node41973;
														assign node41973 = (inp[0]) ? node41981 : node41974;
															assign node41974 = (inp[10]) ? node41978 : node41975;
																assign node41975 = (inp[9]) ? 4'b0100 : 4'b0010;
																assign node41978 = (inp[9]) ? 4'b0000 : 4'b0100;
															assign node41981 = (inp[9]) ? node41985 : node41982;
																assign node41982 = (inp[10]) ? 4'b0110 : 4'b0000;
																assign node41985 = (inp[10]) ? 4'b0010 : 4'b0110;
														assign node41988 = (inp[0]) ? node41992 : node41989;
															assign node41989 = (inp[9]) ? 4'b0010 : 4'b0000;
															assign node41992 = (inp[9]) ? 4'b0000 : 4'b0010;
										assign node41995 = (inp[10]) ? node42049 : node41996;
											assign node41996 = (inp[0]) ? node42022 : node41997;
												assign node41997 = (inp[4]) ? node42011 : node41998;
													assign node41998 = (inp[9]) ? node42004 : node41999;
														assign node41999 = (inp[3]) ? node42001 : 4'b0110;
															assign node42001 = (inp[15]) ? 4'b0110 : 4'b0100;
														assign node42004 = (inp[15]) ? node42008 : node42005;
															assign node42005 = (inp[3]) ? 4'b0000 : 4'b0010;
															assign node42008 = (inp[3]) ? 4'b0010 : 4'b0000;
													assign node42011 = (inp[9]) ? node42019 : node42012;
														assign node42012 = (inp[15]) ? node42016 : node42013;
															assign node42013 = (inp[3]) ? 4'b0000 : 4'b0010;
															assign node42016 = (inp[3]) ? 4'b0010 : 4'b0000;
														assign node42019 = (inp[15]) ? 4'b0110 : 4'b0100;
												assign node42022 = (inp[15]) ? node42034 : node42023;
													assign node42023 = (inp[3]) ? node42029 : node42024;
														assign node42024 = (inp[9]) ? 4'b0110 : node42025;
															assign node42025 = (inp[4]) ? 4'b0000 : 4'b0100;
														assign node42029 = (inp[4]) ? node42031 : 4'b0110;
															assign node42031 = (inp[9]) ? 4'b0110 : 4'b0010;
													assign node42034 = (inp[3]) ? node42040 : node42035;
														assign node42035 = (inp[4]) ? 4'b0100 : node42036;
															assign node42036 = (inp[9]) ? 4'b0010 : 4'b0110;
														assign node42040 = (inp[12]) ? node42042 : 4'b0000;
															assign node42042 = (inp[4]) ? node42046 : node42043;
																assign node42043 = (inp[9]) ? 4'b0000 : 4'b0100;
																assign node42046 = (inp[9]) ? 4'b0100 : 4'b0000;
											assign node42049 = (inp[3]) ? node42107 : node42050;
												assign node42050 = (inp[15]) ? node42078 : node42051;
													assign node42051 = (inp[12]) ? node42067 : node42052;
														assign node42052 = (inp[0]) ? node42060 : node42053;
															assign node42053 = (inp[9]) ? node42057 : node42054;
																assign node42054 = (inp[4]) ? 4'b0010 : 4'b0110;
																assign node42057 = (inp[4]) ? 4'b0100 : 4'b0010;
															assign node42060 = (inp[4]) ? node42064 : node42061;
																assign node42061 = (inp[9]) ? 4'b0000 : 4'b0100;
																assign node42064 = (inp[9]) ? 4'b0110 : 4'b0000;
														assign node42067 = (inp[0]) ? node42073 : node42068;
															assign node42068 = (inp[4]) ? node42070 : 4'b0100;
																assign node42070 = (inp[9]) ? 4'b0000 : 4'b0100;
															assign node42073 = (inp[4]) ? 4'b0110 : node42074;
																assign node42074 = (inp[9]) ? 4'b0110 : 4'b0000;
													assign node42078 = (inp[12]) ? node42092 : node42079;
														assign node42079 = (inp[0]) ? node42085 : node42080;
															assign node42080 = (inp[4]) ? 4'b0000 : node42081;
																assign node42081 = (inp[9]) ? 4'b0000 : 4'b0100;
															assign node42085 = (inp[9]) ? node42089 : node42086;
																assign node42086 = (inp[4]) ? 4'b0010 : 4'b0110;
																assign node42089 = (inp[4]) ? 4'b0100 : 4'b0010;
														assign node42092 = (inp[0]) ? node42100 : node42093;
															assign node42093 = (inp[9]) ? node42097 : node42094;
																assign node42094 = (inp[4]) ? 4'b0110 : 4'b0000;
																assign node42097 = (inp[4]) ? 4'b0010 : 4'b0110;
															assign node42100 = (inp[4]) ? node42104 : node42101;
																assign node42101 = (inp[9]) ? 4'b0100 : 4'b0010;
																assign node42104 = (inp[9]) ? 4'b0000 : 4'b0100;
												assign node42107 = (inp[15]) ? node42135 : node42108;
													assign node42108 = (inp[0]) ? node42122 : node42109;
														assign node42109 = (inp[9]) ? node42115 : node42110;
															assign node42110 = (inp[12]) ? node42112 : 4'b0000;
																assign node42112 = (inp[4]) ? 4'b0100 : 4'b0000;
															assign node42115 = (inp[4]) ? node42119 : node42116;
																assign node42116 = (inp[12]) ? 4'b0100 : 4'b0000;
																assign node42119 = (inp[12]) ? 4'b0000 : 4'b0100;
														assign node42122 = (inp[4]) ? node42130 : node42123;
															assign node42123 = (inp[12]) ? node42127 : node42124;
																assign node42124 = (inp[9]) ? 4'b0010 : 4'b0110;
																assign node42127 = (inp[9]) ? 4'b0110 : 4'b0010;
															assign node42130 = (inp[9]) ? 4'b0010 : node42131;
																assign node42131 = (inp[12]) ? 4'b0110 : 4'b0010;
													assign node42135 = (inp[0]) ? node42143 : node42136;
														assign node42136 = (inp[9]) ? node42138 : 4'b0010;
															assign node42138 = (inp[12]) ? 4'b0010 : node42139;
																assign node42139 = (inp[4]) ? 4'b0110 : 4'b0010;
														assign node42143 = (inp[12]) ? node42149 : node42144;
															assign node42144 = (inp[4]) ? 4'b0000 : node42145;
																assign node42145 = (inp[9]) ? 4'b0000 : 4'b0100;
															assign node42149 = (inp[9]) ? node42153 : node42150;
																assign node42150 = (inp[4]) ? 4'b0100 : 4'b0000;
																assign node42153 = (inp[4]) ? 4'b0000 : 4'b0100;
								assign node42156 = (inp[9]) ? node42356 : node42157;
									assign node42157 = (inp[4]) ? node42249 : node42158;
										assign node42158 = (inp[12]) ? node42182 : node42159;
											assign node42159 = (inp[0]) ? node42171 : node42160;
												assign node42160 = (inp[15]) ? node42166 : node42161;
													assign node42161 = (inp[3]) ? node42163 : 4'b0110;
														assign node42163 = (inp[5]) ? 4'b0100 : 4'b0110;
													assign node42166 = (inp[3]) ? node42168 : 4'b0100;
														assign node42168 = (inp[5]) ? 4'b0110 : 4'b0100;
												assign node42171 = (inp[15]) ? node42177 : node42172;
													assign node42172 = (inp[3]) ? node42174 : 4'b0100;
														assign node42174 = (inp[5]) ? 4'b0110 : 4'b0100;
													assign node42177 = (inp[5]) ? node42179 : 4'b0110;
														assign node42179 = (inp[3]) ? 4'b0100 : 4'b0110;
											assign node42182 = (inp[10]) ? node42206 : node42183;
												assign node42183 = (inp[15]) ? node42195 : node42184;
													assign node42184 = (inp[0]) ? node42190 : node42185;
														assign node42185 = (inp[5]) ? node42187 : 4'b0110;
															assign node42187 = (inp[3]) ? 4'b0100 : 4'b0110;
														assign node42190 = (inp[5]) ? node42192 : 4'b0100;
															assign node42192 = (inp[3]) ? 4'b0110 : 4'b0100;
													assign node42195 = (inp[0]) ? node42201 : node42196;
														assign node42196 = (inp[5]) ? node42198 : 4'b0100;
															assign node42198 = (inp[3]) ? 4'b0110 : 4'b0100;
														assign node42201 = (inp[5]) ? node42203 : 4'b0110;
															assign node42203 = (inp[3]) ? 4'b0100 : 4'b0110;
												assign node42206 = (inp[5]) ? node42220 : node42207;
													assign node42207 = (inp[3]) ? node42215 : node42208;
														assign node42208 = (inp[0]) ? node42212 : node42209;
															assign node42209 = (inp[15]) ? 4'b0000 : 4'b0010;
															assign node42212 = (inp[15]) ? 4'b0010 : 4'b0000;
														assign node42215 = (inp[0]) ? node42217 : 4'b0000;
															assign node42217 = (inp[15]) ? 4'b0010 : 4'b0000;
													assign node42220 = (inp[14]) ? node42236 : node42221;
														assign node42221 = (inp[3]) ? node42229 : node42222;
															assign node42222 = (inp[15]) ? node42226 : node42223;
																assign node42223 = (inp[0]) ? 4'b0000 : 4'b0010;
																assign node42226 = (inp[0]) ? 4'b0010 : 4'b0000;
															assign node42229 = (inp[0]) ? node42233 : node42230;
																assign node42230 = (inp[15]) ? 4'b0010 : 4'b0000;
																assign node42233 = (inp[15]) ? 4'b0000 : 4'b0010;
														assign node42236 = (inp[3]) ? node42244 : node42237;
															assign node42237 = (inp[0]) ? node42241 : node42238;
																assign node42238 = (inp[15]) ? 4'b0000 : 4'b0010;
																assign node42241 = (inp[15]) ? 4'b0010 : 4'b0000;
															assign node42244 = (inp[15]) ? 4'b0010 : node42245;
																assign node42245 = (inp[0]) ? 4'b0010 : 4'b0000;
										assign node42249 = (inp[10]) ? node42305 : node42250;
											assign node42250 = (inp[12]) ? node42266 : node42251;
												assign node42251 = (inp[15]) ? node42263 : node42252;
													assign node42252 = (inp[0]) ? node42258 : node42253;
														assign node42253 = (inp[5]) ? node42255 : 4'b0010;
															assign node42255 = (inp[3]) ? 4'b0000 : 4'b0010;
														assign node42258 = (inp[3]) ? node42260 : 4'b0000;
															assign node42260 = (inp[5]) ? 4'b0010 : 4'b0000;
													assign node42263 = (inp[0]) ? 4'b0010 : 4'b0000;
												assign node42266 = (inp[3]) ? node42290 : node42267;
													assign node42267 = (inp[5]) ? node42275 : node42268;
														assign node42268 = (inp[0]) ? node42272 : node42269;
															assign node42269 = (inp[14]) ? 4'b0000 : 4'b0010;
															assign node42272 = (inp[15]) ? 4'b0010 : 4'b0000;
														assign node42275 = (inp[14]) ? node42283 : node42276;
															assign node42276 = (inp[15]) ? node42280 : node42277;
																assign node42277 = (inp[0]) ? 4'b0000 : 4'b0010;
																assign node42280 = (inp[0]) ? 4'b0010 : 4'b0000;
															assign node42283 = (inp[0]) ? node42287 : node42284;
																assign node42284 = (inp[15]) ? 4'b0000 : 4'b0010;
																assign node42287 = (inp[15]) ? 4'b0010 : 4'b0000;
													assign node42290 = (inp[5]) ? node42298 : node42291;
														assign node42291 = (inp[15]) ? node42295 : node42292;
															assign node42292 = (inp[0]) ? 4'b0000 : 4'b0010;
															assign node42295 = (inp[0]) ? 4'b0010 : 4'b0000;
														assign node42298 = (inp[15]) ? node42302 : node42299;
															assign node42299 = (inp[0]) ? 4'b0010 : 4'b0000;
															assign node42302 = (inp[0]) ? 4'b0000 : 4'b0010;
											assign node42305 = (inp[12]) ? node42327 : node42306;
												assign node42306 = (inp[15]) ? node42318 : node42307;
													assign node42307 = (inp[0]) ? node42313 : node42308;
														assign node42308 = (inp[5]) ? node42310 : 4'b0010;
															assign node42310 = (inp[3]) ? 4'b0000 : 4'b0010;
														assign node42313 = (inp[3]) ? node42315 : 4'b0000;
															assign node42315 = (inp[5]) ? 4'b0010 : 4'b0000;
													assign node42318 = (inp[0]) ? node42324 : node42319;
														assign node42319 = (inp[3]) ? node42321 : 4'b0000;
															assign node42321 = (inp[5]) ? 4'b0010 : 4'b0000;
														assign node42324 = (inp[3]) ? 4'b0000 : 4'b0010;
												assign node42327 = (inp[0]) ? node42339 : node42328;
													assign node42328 = (inp[15]) ? node42334 : node42329;
														assign node42329 = (inp[3]) ? 4'b0100 : node42330;
															assign node42330 = (inp[5]) ? 4'b0100 : 4'b0110;
														assign node42334 = (inp[3]) ? 4'b0110 : node42335;
															assign node42335 = (inp[5]) ? 4'b0110 : 4'b0100;
													assign node42339 = (inp[3]) ? node42353 : node42340;
														assign node42340 = (inp[14]) ? node42348 : node42341;
															assign node42341 = (inp[5]) ? node42345 : node42342;
																assign node42342 = (inp[15]) ? 4'b0110 : 4'b0100;
																assign node42345 = (inp[15]) ? 4'b0100 : 4'b0110;
															assign node42348 = (inp[15]) ? 4'b0110 : node42349;
																assign node42349 = (inp[5]) ? 4'b0110 : 4'b0100;
														assign node42353 = (inp[15]) ? 4'b0100 : 4'b0110;
									assign node42356 = (inp[4]) ? node42454 : node42357;
										assign node42357 = (inp[10]) ? node42387 : node42358;
											assign node42358 = (inp[5]) ? node42366 : node42359;
												assign node42359 = (inp[15]) ? node42363 : node42360;
													assign node42360 = (inp[0]) ? 4'b0000 : 4'b0010;
													assign node42363 = (inp[0]) ? 4'b0010 : 4'b0000;
												assign node42366 = (inp[15]) ? node42380 : node42367;
													assign node42367 = (inp[12]) ? node42373 : node42368;
														assign node42368 = (inp[3]) ? 4'b0000 : node42369;
															assign node42369 = (inp[0]) ? 4'b0000 : 4'b0010;
														assign node42373 = (inp[3]) ? node42377 : node42374;
															assign node42374 = (inp[0]) ? 4'b0000 : 4'b0010;
															assign node42377 = (inp[0]) ? 4'b0010 : 4'b0000;
													assign node42380 = (inp[0]) ? node42384 : node42381;
														assign node42381 = (inp[3]) ? 4'b0010 : 4'b0000;
														assign node42384 = (inp[3]) ? 4'b0000 : 4'b0010;
											assign node42387 = (inp[12]) ? node42429 : node42388;
												assign node42388 = (inp[3]) ? node42406 : node42389;
													assign node42389 = (inp[14]) ? node42397 : node42390;
														assign node42390 = (inp[15]) ? node42394 : node42391;
															assign node42391 = (inp[0]) ? 4'b0000 : 4'b0010;
															assign node42394 = (inp[0]) ? 4'b0010 : 4'b0000;
														assign node42397 = (inp[5]) ? node42399 : 4'b0010;
															assign node42399 = (inp[0]) ? node42403 : node42400;
																assign node42400 = (inp[15]) ? 4'b0000 : 4'b0010;
																assign node42403 = (inp[15]) ? 4'b0010 : 4'b0000;
													assign node42406 = (inp[0]) ? node42414 : node42407;
														assign node42407 = (inp[15]) ? node42411 : node42408;
															assign node42408 = (inp[5]) ? 4'b0000 : 4'b0010;
															assign node42411 = (inp[5]) ? 4'b0010 : 4'b0000;
														assign node42414 = (inp[14]) ? node42422 : node42415;
															assign node42415 = (inp[5]) ? node42419 : node42416;
																assign node42416 = (inp[15]) ? 4'b0010 : 4'b0000;
																assign node42419 = (inp[15]) ? 4'b0000 : 4'b0010;
															assign node42422 = (inp[5]) ? node42426 : node42423;
																assign node42423 = (inp[15]) ? 4'b0010 : 4'b0000;
																assign node42426 = (inp[15]) ? 4'b0000 : 4'b0010;
												assign node42429 = (inp[5]) ? node42447 : node42430;
													assign node42430 = (inp[3]) ? node42440 : node42431;
														assign node42431 = (inp[14]) ? node42433 : 4'b0100;
															assign node42433 = (inp[0]) ? node42437 : node42434;
																assign node42434 = (inp[15]) ? 4'b0100 : 4'b0110;
																assign node42437 = (inp[15]) ? 4'b0110 : 4'b0100;
														assign node42440 = (inp[0]) ? node42444 : node42441;
															assign node42441 = (inp[15]) ? 4'b0110 : 4'b0100;
															assign node42444 = (inp[15]) ? 4'b0100 : 4'b0110;
													assign node42447 = (inp[0]) ? node42451 : node42448;
														assign node42448 = (inp[15]) ? 4'b0110 : 4'b0100;
														assign node42451 = (inp[15]) ? 4'b0100 : 4'b0110;
										assign node42454 = (inp[12]) ? node42510 : node42455;
											assign node42455 = (inp[14]) ? node42487 : node42456;
												assign node42456 = (inp[10]) ? node42474 : node42457;
													assign node42457 = (inp[3]) ? node42467 : node42458;
														assign node42458 = (inp[15]) ? 4'b0110 : node42459;
															assign node42459 = (inp[5]) ? node42463 : node42460;
																assign node42460 = (inp[0]) ? 4'b0100 : 4'b0110;
																assign node42463 = (inp[0]) ? 4'b0110 : 4'b0100;
														assign node42467 = (inp[0]) ? node42471 : node42468;
															assign node42468 = (inp[15]) ? 4'b0110 : 4'b0100;
															assign node42471 = (inp[15]) ? 4'b0100 : 4'b0110;
													assign node42474 = (inp[3]) ? node42476 : 4'b0100;
														assign node42476 = (inp[5]) ? node42482 : node42477;
															assign node42477 = (inp[0]) ? node42479 : 4'b0100;
																assign node42479 = (inp[15]) ? 4'b0100 : 4'b0110;
															assign node42482 = (inp[15]) ? 4'b0110 : node42483;
																assign node42483 = (inp[0]) ? 4'b0110 : 4'b0100;
												assign node42487 = (inp[15]) ? node42499 : node42488;
													assign node42488 = (inp[0]) ? node42494 : node42489;
														assign node42489 = (inp[5]) ? 4'b0100 : node42490;
															assign node42490 = (inp[3]) ? 4'b0100 : 4'b0110;
														assign node42494 = (inp[3]) ? 4'b0110 : node42495;
															assign node42495 = (inp[5]) ? 4'b0110 : 4'b0100;
													assign node42499 = (inp[0]) ? node42505 : node42500;
														assign node42500 = (inp[5]) ? 4'b0110 : node42501;
															assign node42501 = (inp[3]) ? 4'b0110 : 4'b0100;
														assign node42505 = (inp[5]) ? 4'b0100 : node42506;
															assign node42506 = (inp[3]) ? 4'b0100 : 4'b0110;
											assign node42510 = (inp[10]) ? node42534 : node42511;
												assign node42511 = (inp[0]) ? node42523 : node42512;
													assign node42512 = (inp[15]) ? node42518 : node42513;
														assign node42513 = (inp[3]) ? 4'b0100 : node42514;
															assign node42514 = (inp[5]) ? 4'b0100 : 4'b0110;
														assign node42518 = (inp[14]) ? node42520 : 4'b0110;
															assign node42520 = (inp[3]) ? 4'b0110 : 4'b0100;
													assign node42523 = (inp[15]) ? node42529 : node42524;
														assign node42524 = (inp[5]) ? 4'b0110 : node42525;
															assign node42525 = (inp[3]) ? 4'b0110 : 4'b0100;
														assign node42529 = (inp[5]) ? 4'b0100 : node42530;
															assign node42530 = (inp[3]) ? 4'b0100 : 4'b0110;
												assign node42534 = (inp[0]) ? node42546 : node42535;
													assign node42535 = (inp[15]) ? node42541 : node42536;
														assign node42536 = (inp[3]) ? 4'b0000 : node42537;
															assign node42537 = (inp[14]) ? 4'b0000 : 4'b0010;
														assign node42541 = (inp[5]) ? 4'b0010 : node42542;
															assign node42542 = (inp[14]) ? 4'b0000 : 4'b0010;
													assign node42546 = (inp[15]) ? node42550 : node42547;
														assign node42547 = (inp[3]) ? 4'b0010 : 4'b0000;
														assign node42550 = (inp[3]) ? 4'b0000 : node42551;
															assign node42551 = (inp[14]) ? 4'b0010 : 4'b0000;
							assign node42555 = (inp[2]) ? node43145 : node42556;
								assign node42556 = (inp[14]) ? node42892 : node42557;
									assign node42557 = (inp[10]) ? node42687 : node42558;
										assign node42558 = (inp[4]) ? node42624 : node42559;
											assign node42559 = (inp[9]) ? node42587 : node42560;
												assign node42560 = (inp[5]) ? node42570 : node42561;
													assign node42561 = (inp[3]) ? node42563 : 4'b0100;
														assign node42563 = (inp[15]) ? node42567 : node42564;
															assign node42564 = (inp[0]) ? 4'b0100 : 4'b0110;
															assign node42567 = (inp[0]) ? 4'b0110 : 4'b0100;
													assign node42570 = (inp[0]) ? node42578 : node42571;
														assign node42571 = (inp[3]) ? node42575 : node42572;
															assign node42572 = (inp[15]) ? 4'b0100 : 4'b0110;
															assign node42575 = (inp[15]) ? 4'b0110 : 4'b0100;
														assign node42578 = (inp[12]) ? node42584 : node42579;
															assign node42579 = (inp[3]) ? 4'b0110 : node42580;
																assign node42580 = (inp[15]) ? 4'b0110 : 4'b0100;
															assign node42584 = (inp[15]) ? 4'b0100 : 4'b0110;
												assign node42587 = (inp[12]) ? node42601 : node42588;
													assign node42588 = (inp[0]) ? node42594 : node42589;
														assign node42589 = (inp[15]) ? node42591 : 4'b0010;
															assign node42591 = (inp[3]) ? 4'b0010 : 4'b0000;
														assign node42594 = (inp[15]) ? 4'b0010 : node42595;
															assign node42595 = (inp[3]) ? node42597 : 4'b0000;
																assign node42597 = (inp[5]) ? 4'b0010 : 4'b0000;
													assign node42601 = (inp[5]) ? node42609 : node42602;
														assign node42602 = (inp[0]) ? node42606 : node42603;
															assign node42603 = (inp[15]) ? 4'b0000 : 4'b0010;
															assign node42606 = (inp[15]) ? 4'b0010 : 4'b0000;
														assign node42609 = (inp[0]) ? node42617 : node42610;
															assign node42610 = (inp[3]) ? node42614 : node42611;
																assign node42611 = (inp[15]) ? 4'b0000 : 4'b0010;
																assign node42614 = (inp[15]) ? 4'b0010 : 4'b0000;
															assign node42617 = (inp[3]) ? node42621 : node42618;
																assign node42618 = (inp[15]) ? 4'b0010 : 4'b0000;
																assign node42621 = (inp[15]) ? 4'b0000 : 4'b0010;
											assign node42624 = (inp[9]) ? node42648 : node42625;
												assign node42625 = (inp[0]) ? node42637 : node42626;
													assign node42626 = (inp[15]) ? node42632 : node42627;
														assign node42627 = (inp[5]) ? node42629 : 4'b0010;
															assign node42629 = (inp[3]) ? 4'b0000 : 4'b0010;
														assign node42632 = (inp[5]) ? node42634 : 4'b0000;
															assign node42634 = (inp[3]) ? 4'b0010 : 4'b0000;
													assign node42637 = (inp[15]) ? node42643 : node42638;
														assign node42638 = (inp[5]) ? node42640 : 4'b0000;
															assign node42640 = (inp[3]) ? 4'b0010 : 4'b0000;
														assign node42643 = (inp[5]) ? node42645 : 4'b0010;
															assign node42645 = (inp[3]) ? 4'b0000 : 4'b0010;
												assign node42648 = (inp[3]) ? node42672 : node42649;
													assign node42649 = (inp[15]) ? node42665 : node42650;
														assign node42650 = (inp[12]) ? node42658 : node42651;
															assign node42651 = (inp[5]) ? node42655 : node42652;
																assign node42652 = (inp[0]) ? 4'b0100 : 4'b0110;
																assign node42655 = (inp[0]) ? 4'b0110 : 4'b0100;
															assign node42658 = (inp[0]) ? node42662 : node42659;
																assign node42659 = (inp[5]) ? 4'b0100 : 4'b0110;
																assign node42662 = (inp[5]) ? 4'b0110 : 4'b0100;
														assign node42665 = (inp[5]) ? node42669 : node42666;
															assign node42666 = (inp[0]) ? 4'b0110 : 4'b0100;
															assign node42669 = (inp[0]) ? 4'b0100 : 4'b0110;
													assign node42672 = (inp[5]) ? node42680 : node42673;
														assign node42673 = (inp[15]) ? node42677 : node42674;
															assign node42674 = (inp[0]) ? 4'b0110 : 4'b0100;
															assign node42677 = (inp[0]) ? 4'b0100 : 4'b0110;
														assign node42680 = (inp[15]) ? node42684 : node42681;
															assign node42681 = (inp[0]) ? 4'b0110 : 4'b0100;
															assign node42684 = (inp[0]) ? 4'b0100 : 4'b0110;
										assign node42687 = (inp[15]) ? node42789 : node42688;
											assign node42688 = (inp[5]) ? node42740 : node42689;
												assign node42689 = (inp[0]) ? node42717 : node42690;
													assign node42690 = (inp[3]) ? node42704 : node42691;
														assign node42691 = (inp[9]) ? node42699 : node42692;
															assign node42692 = (inp[12]) ? node42696 : node42693;
																assign node42693 = (inp[4]) ? 4'b0010 : 4'b0110;
																assign node42696 = (inp[4]) ? 4'b0110 : 4'b0010;
															assign node42699 = (inp[4]) ? 4'b0010 : node42700;
																assign node42700 = (inp[12]) ? 4'b0110 : 4'b0010;
														assign node42704 = (inp[4]) ? node42712 : node42705;
															assign node42705 = (inp[12]) ? node42709 : node42706;
																assign node42706 = (inp[9]) ? 4'b0010 : 4'b0110;
																assign node42709 = (inp[9]) ? 4'b0100 : 4'b0010;
															assign node42712 = (inp[9]) ? 4'b0100 : node42713;
																assign node42713 = (inp[12]) ? 4'b0100 : 4'b0010;
													assign node42717 = (inp[3]) ? node42733 : node42718;
														assign node42718 = (inp[4]) ? node42726 : node42719;
															assign node42719 = (inp[12]) ? node42723 : node42720;
																assign node42720 = (inp[9]) ? 4'b0000 : 4'b0100;
																assign node42723 = (inp[9]) ? 4'b0100 : 4'b0000;
															assign node42726 = (inp[12]) ? node42730 : node42727;
																assign node42727 = (inp[9]) ? 4'b0100 : 4'b0000;
																assign node42730 = (inp[9]) ? 4'b0000 : 4'b0100;
														assign node42733 = (inp[9]) ? node42735 : 4'b0000;
															assign node42735 = (inp[12]) ? node42737 : 4'b0110;
																assign node42737 = (inp[4]) ? 4'b0010 : 4'b0110;
												assign node42740 = (inp[0]) ? node42766 : node42741;
													assign node42741 = (inp[4]) ? node42755 : node42742;
														assign node42742 = (inp[3]) ? node42748 : node42743;
															assign node42743 = (inp[12]) ? node42745 : 4'b0010;
																assign node42745 = (inp[9]) ? 4'b0100 : 4'b0010;
															assign node42748 = (inp[12]) ? node42752 : node42749;
																assign node42749 = (inp[9]) ? 4'b0000 : 4'b0100;
																assign node42752 = (inp[9]) ? 4'b0100 : 4'b0000;
														assign node42755 = (inp[3]) ? node42761 : node42756;
															assign node42756 = (inp[12]) ? node42758 : 4'b0100;
																assign node42758 = (inp[9]) ? 4'b0000 : 4'b0100;
															assign node42761 = (inp[12]) ? 4'b0100 : node42762;
																assign node42762 = (inp[9]) ? 4'b0100 : 4'b0000;
													assign node42766 = (inp[3]) ? node42782 : node42767;
														assign node42767 = (inp[12]) ? node42775 : node42768;
															assign node42768 = (inp[4]) ? node42772 : node42769;
																assign node42769 = (inp[9]) ? 4'b0000 : 4'b0100;
																assign node42772 = (inp[9]) ? 4'b0110 : 4'b0000;
															assign node42775 = (inp[4]) ? node42779 : node42776;
																assign node42776 = (inp[9]) ? 4'b0110 : 4'b0000;
																assign node42779 = (inp[9]) ? 4'b0010 : 4'b0110;
														assign node42782 = (inp[12]) ? node42784 : 4'b0110;
															assign node42784 = (inp[4]) ? node42786 : 4'b0010;
																assign node42786 = (inp[9]) ? 4'b0010 : 4'b0110;
											assign node42789 = (inp[0]) ? node42839 : node42790;
												assign node42790 = (inp[5]) ? node42816 : node42791;
													assign node42791 = (inp[3]) ? node42807 : node42792;
														assign node42792 = (inp[9]) ? node42800 : node42793;
															assign node42793 = (inp[4]) ? node42797 : node42794;
																assign node42794 = (inp[12]) ? 4'b0000 : 4'b0100;
																assign node42797 = (inp[12]) ? 4'b0100 : 4'b0000;
															assign node42800 = (inp[12]) ? node42804 : node42801;
																assign node42801 = (inp[4]) ? 4'b0100 : 4'b0000;
																assign node42804 = (inp[4]) ? 4'b0000 : 4'b0100;
														assign node42807 = (inp[4]) ? node42813 : node42808;
															assign node42808 = (inp[12]) ? 4'b0000 : node42809;
																assign node42809 = (inp[9]) ? 4'b0000 : 4'b0100;
															assign node42813 = (inp[9]) ? 4'b0110 : 4'b0000;
													assign node42816 = (inp[3]) ? node42828 : node42817;
														assign node42817 = (inp[12]) ? node42823 : node42818;
															assign node42818 = (inp[4]) ? 4'b0000 : node42819;
																assign node42819 = (inp[9]) ? 4'b0000 : 4'b0100;
															assign node42823 = (inp[4]) ? 4'b0110 : node42824;
																assign node42824 = (inp[9]) ? 4'b0110 : 4'b0000;
														assign node42828 = (inp[9]) ? node42834 : node42829;
															assign node42829 = (inp[4]) ? node42831 : 4'b0110;
																assign node42831 = (inp[12]) ? 4'b0110 : 4'b0010;
															assign node42834 = (inp[12]) ? 4'b0010 : node42835;
																assign node42835 = (inp[4]) ? 4'b0110 : 4'b0010;
												assign node42839 = (inp[5]) ? node42869 : node42840;
													assign node42840 = (inp[3]) ? node42856 : node42841;
														assign node42841 = (inp[4]) ? node42849 : node42842;
															assign node42842 = (inp[12]) ? node42846 : node42843;
																assign node42843 = (inp[9]) ? 4'b0010 : 4'b0110;
																assign node42846 = (inp[9]) ? 4'b0110 : 4'b0010;
															assign node42849 = (inp[9]) ? node42853 : node42850;
																assign node42850 = (inp[12]) ? 4'b0110 : 4'b0010;
																assign node42853 = (inp[12]) ? 4'b0010 : 4'b0110;
														assign node42856 = (inp[9]) ? node42864 : node42857;
															assign node42857 = (inp[12]) ? node42861 : node42858;
																assign node42858 = (inp[4]) ? 4'b0010 : 4'b0110;
																assign node42861 = (inp[4]) ? 4'b0100 : 4'b0010;
															assign node42864 = (inp[4]) ? node42866 : 4'b0100;
																assign node42866 = (inp[12]) ? 4'b0000 : 4'b0100;
													assign node42869 = (inp[3]) ? node42879 : node42870;
														assign node42870 = (inp[9]) ? node42872 : 4'b0010;
															assign node42872 = (inp[12]) ? node42876 : node42873;
																assign node42873 = (inp[4]) ? 4'b0100 : 4'b0010;
																assign node42876 = (inp[4]) ? 4'b0000 : 4'b0100;
														assign node42879 = (inp[9]) ? node42885 : node42880;
															assign node42880 = (inp[12]) ? 4'b0000 : node42881;
																assign node42881 = (inp[4]) ? 4'b0000 : 4'b0100;
															assign node42885 = (inp[12]) ? node42889 : node42886;
																assign node42886 = (inp[4]) ? 4'b0100 : 4'b0000;
																assign node42889 = (inp[4]) ? 4'b0000 : 4'b0100;
									assign node42892 = (inp[12]) ? node43030 : node42893;
										assign node42893 = (inp[10]) ? node42957 : node42894;
											assign node42894 = (inp[9]) ? node42924 : node42895;
												assign node42895 = (inp[4]) ? node42909 : node42896;
													assign node42896 = (inp[0]) ? 4'b1101 : node42897;
														assign node42897 = (inp[15]) ? node42903 : node42898;
															assign node42898 = (inp[3]) ? node42900 : 4'b1111;
																assign node42900 = (inp[5]) ? 4'b1101 : 4'b1111;
															assign node42903 = (inp[5]) ? node42905 : 4'b1101;
																assign node42905 = (inp[3]) ? 4'b1111 : 4'b1101;
													assign node42909 = (inp[5]) ? node42917 : node42910;
														assign node42910 = (inp[3]) ? 4'b1011 : node42911;
															assign node42911 = (inp[0]) ? node42913 : 4'b1011;
																assign node42913 = (inp[15]) ? 4'b1011 : 4'b1001;
														assign node42917 = (inp[15]) ? 4'b1001 : node42918;
															assign node42918 = (inp[3]) ? 4'b1001 : node42919;
																assign node42919 = (inp[0]) ? 4'b1001 : 4'b1011;
												assign node42924 = (inp[4]) ? node42940 : node42925;
													assign node42925 = (inp[0]) ? node42935 : node42926;
														assign node42926 = (inp[3]) ? node42930 : node42927;
															assign node42927 = (inp[15]) ? 4'b1001 : 4'b1011;
															assign node42930 = (inp[5]) ? node42932 : 4'b1011;
																assign node42932 = (inp[15]) ? 4'b1011 : 4'b1001;
														assign node42935 = (inp[3]) ? node42937 : 4'b1011;
															assign node42937 = (inp[5]) ? 4'b1011 : 4'b1001;
													assign node42940 = (inp[15]) ? node42948 : node42941;
														assign node42941 = (inp[0]) ? node42945 : node42942;
															assign node42942 = (inp[3]) ? 4'b1101 : 4'b1111;
															assign node42945 = (inp[3]) ? 4'b1111 : 4'b1101;
														assign node42948 = (inp[3]) ? 4'b1111 : node42949;
															assign node42949 = (inp[5]) ? node42953 : node42950;
																assign node42950 = (inp[0]) ? 4'b1111 : 4'b1101;
																assign node42953 = (inp[0]) ? 4'b1101 : 4'b1111;
											assign node42957 = (inp[9]) ? node42987 : node42958;
												assign node42958 = (inp[4]) ? node42974 : node42959;
													assign node42959 = (inp[15]) ? node42965 : node42960;
														assign node42960 = (inp[5]) ? 4'b1011 : node42961;
															assign node42961 = (inp[0]) ? 4'b1001 : 4'b1011;
														assign node42965 = (inp[0]) ? node42971 : node42966;
															assign node42966 = (inp[5]) ? node42968 : 4'b1001;
																assign node42968 = (inp[3]) ? 4'b1011 : 4'b1001;
															assign node42971 = (inp[3]) ? 4'b1001 : 4'b1011;
													assign node42974 = (inp[15]) ? node42978 : node42975;
														assign node42975 = (inp[5]) ? 4'b1101 : 4'b1111;
														assign node42978 = (inp[0]) ? node42984 : node42979;
															assign node42979 = (inp[3]) ? 4'b1111 : node42980;
																assign node42980 = (inp[5]) ? 4'b1111 : 4'b1101;
															assign node42984 = (inp[3]) ? 4'b1101 : 4'b1111;
												assign node42987 = (inp[4]) ? node43009 : node42988;
													assign node42988 = (inp[0]) ? node42998 : node42989;
														assign node42989 = (inp[3]) ? 4'b1101 : node42990;
															assign node42990 = (inp[5]) ? node42994 : node42991;
																assign node42991 = (inp[15]) ? 4'b1101 : 4'b1111;
																assign node42994 = (inp[15]) ? 4'b1111 : 4'b1101;
														assign node42998 = (inp[15]) ? node43004 : node42999;
															assign node42999 = (inp[3]) ? 4'b1111 : node43000;
																assign node43000 = (inp[5]) ? 4'b1111 : 4'b1101;
															assign node43004 = (inp[3]) ? 4'b1101 : node43005;
																assign node43005 = (inp[5]) ? 4'b1101 : 4'b1111;
													assign node43009 = (inp[5]) ? node43023 : node43010;
														assign node43010 = (inp[0]) ? node43018 : node43011;
															assign node43011 = (inp[15]) ? node43015 : node43012;
																assign node43012 = (inp[3]) ? 4'b1001 : 4'b1011;
																assign node43015 = (inp[3]) ? 4'b1011 : 4'b1001;
															assign node43018 = (inp[15]) ? 4'b1001 : node43019;
																assign node43019 = (inp[3]) ? 4'b1011 : 4'b1001;
														assign node43023 = (inp[3]) ? node43025 : 4'b1001;
															assign node43025 = (inp[15]) ? node43027 : 4'b1001;
																assign node43027 = (inp[0]) ? 4'b1001 : 4'b1011;
										assign node43030 = (inp[3]) ? node43096 : node43031;
											assign node43031 = (inp[5]) ? node43065 : node43032;
												assign node43032 = (inp[4]) ? node43044 : node43033;
													assign node43033 = (inp[9]) ? node43041 : node43034;
														assign node43034 = (inp[15]) ? node43038 : node43035;
															assign node43035 = (inp[0]) ? 4'b1001 : 4'b1011;
															assign node43038 = (inp[0]) ? 4'b1011 : 4'b1001;
														assign node43041 = (inp[0]) ? 4'b1111 : 4'b1101;
													assign node43044 = (inp[9]) ? node43054 : node43045;
														assign node43045 = (inp[10]) ? node43051 : node43046;
															assign node43046 = (inp[15]) ? 4'b1101 : node43047;
																assign node43047 = (inp[0]) ? 4'b1101 : 4'b1111;
															assign node43051 = (inp[15]) ? 4'b1111 : 4'b1101;
														assign node43054 = (inp[10]) ? node43060 : node43055;
															assign node43055 = (inp[15]) ? 4'b1011 : node43056;
																assign node43056 = (inp[0]) ? 4'b1001 : 4'b1011;
															assign node43060 = (inp[0]) ? 4'b1011 : node43061;
																assign node43061 = (inp[15]) ? 4'b1001 : 4'b1011;
												assign node43065 = (inp[0]) ? node43081 : node43066;
													assign node43066 = (inp[15]) ? node43074 : node43067;
														assign node43067 = (inp[4]) ? node43071 : node43068;
															assign node43068 = (inp[9]) ? 4'b1101 : 4'b1011;
															assign node43071 = (inp[9]) ? 4'b1001 : 4'b1101;
														assign node43074 = (inp[9]) ? node43078 : node43075;
															assign node43075 = (inp[4]) ? 4'b1111 : 4'b1001;
															assign node43078 = (inp[4]) ? 4'b1011 : 4'b1111;
													assign node43081 = (inp[15]) ? node43089 : node43082;
														assign node43082 = (inp[9]) ? node43086 : node43083;
															assign node43083 = (inp[4]) ? 4'b1111 : 4'b1001;
															assign node43086 = (inp[4]) ? 4'b1011 : 4'b1111;
														assign node43089 = (inp[4]) ? node43093 : node43090;
															assign node43090 = (inp[9]) ? 4'b1101 : 4'b1011;
															assign node43093 = (inp[9]) ? 4'b1001 : 4'b1101;
											assign node43096 = (inp[15]) ? node43126 : node43097;
												assign node43097 = (inp[0]) ? node43111 : node43098;
													assign node43098 = (inp[5]) ? node43104 : node43099;
														assign node43099 = (inp[4]) ? node43101 : 4'b1101;
															assign node43101 = (inp[9]) ? 4'b1001 : 4'b1101;
														assign node43104 = (inp[4]) ? node43108 : node43105;
															assign node43105 = (inp[9]) ? 4'b1101 : 4'b1001;
															assign node43108 = (inp[9]) ? 4'b1001 : 4'b1101;
													assign node43111 = (inp[5]) ? node43119 : node43112;
														assign node43112 = (inp[9]) ? node43116 : node43113;
															assign node43113 = (inp[4]) ? 4'b1111 : 4'b1001;
															assign node43116 = (inp[4]) ? 4'b1011 : 4'b1111;
														assign node43119 = (inp[9]) ? node43123 : node43120;
															assign node43120 = (inp[4]) ? 4'b1111 : 4'b1011;
															assign node43123 = (inp[4]) ? 4'b1011 : 4'b1111;
												assign node43126 = (inp[0]) ? node43136 : node43127;
													assign node43127 = (inp[9]) ? node43133 : node43128;
														assign node43128 = (inp[4]) ? 4'b1111 : node43129;
															assign node43129 = (inp[5]) ? 4'b1011 : 4'b1001;
														assign node43133 = (inp[4]) ? 4'b1011 : 4'b1111;
													assign node43136 = (inp[4]) ? node43142 : node43137;
														assign node43137 = (inp[9]) ? 4'b1101 : node43138;
															assign node43138 = (inp[5]) ? 4'b1001 : 4'b1011;
														assign node43142 = (inp[9]) ? 4'b1001 : 4'b1101;
								assign node43145 = (inp[9]) ? node43365 : node43146;
									assign node43146 = (inp[4]) ? node43252 : node43147;
										assign node43147 = (inp[12]) ? node43197 : node43148;
											assign node43148 = (inp[10]) ? node43172 : node43149;
												assign node43149 = (inp[0]) ? node43161 : node43150;
													assign node43150 = (inp[15]) ? node43156 : node43151;
														assign node43151 = (inp[3]) ? node43153 : 4'b1111;
															assign node43153 = (inp[5]) ? 4'b1101 : 4'b1111;
														assign node43156 = (inp[5]) ? node43158 : 4'b1101;
															assign node43158 = (inp[3]) ? 4'b1111 : 4'b1101;
													assign node43161 = (inp[15]) ? node43167 : node43162;
														assign node43162 = (inp[5]) ? node43164 : 4'b1101;
															assign node43164 = (inp[3]) ? 4'b1111 : 4'b1101;
														assign node43167 = (inp[5]) ? node43169 : 4'b1111;
															assign node43169 = (inp[3]) ? 4'b1101 : 4'b1111;
												assign node43172 = (inp[3]) ? node43186 : node43173;
													assign node43173 = (inp[14]) ? node43181 : node43174;
														assign node43174 = (inp[0]) ? node43178 : node43175;
															assign node43175 = (inp[15]) ? 4'b1001 : 4'b1011;
															assign node43178 = (inp[15]) ? 4'b1011 : 4'b1001;
														assign node43181 = (inp[5]) ? node43183 : 4'b1001;
															assign node43183 = (inp[0]) ? 4'b1001 : 4'b1011;
													assign node43186 = (inp[14]) ? node43188 : 4'b1001;
														assign node43188 = (inp[5]) ? node43190 : 4'b1001;
															assign node43190 = (inp[15]) ? node43194 : node43191;
																assign node43191 = (inp[0]) ? 4'b1011 : 4'b1001;
																assign node43194 = (inp[0]) ? 4'b1001 : 4'b1011;
											assign node43197 = (inp[5]) ? node43225 : node43198;
												assign node43198 = (inp[14]) ? node43206 : node43199;
													assign node43199 = (inp[15]) ? node43203 : node43200;
														assign node43200 = (inp[0]) ? 4'b1001 : 4'b1011;
														assign node43203 = (inp[0]) ? 4'b1011 : 4'b1001;
													assign node43206 = (inp[3]) ? node43212 : node43207;
														assign node43207 = (inp[15]) ? node43209 : 4'b1011;
															assign node43209 = (inp[10]) ? 4'b1001 : 4'b1011;
														assign node43212 = (inp[10]) ? node43220 : node43213;
															assign node43213 = (inp[15]) ? node43217 : node43214;
																assign node43214 = (inp[0]) ? 4'b1001 : 4'b1011;
																assign node43217 = (inp[0]) ? 4'b1011 : 4'b1001;
															assign node43220 = (inp[0]) ? node43222 : 4'b1011;
																assign node43222 = (inp[15]) ? 4'b1011 : 4'b1001;
												assign node43225 = (inp[14]) ? node43241 : node43226;
													assign node43226 = (inp[3]) ? node43232 : node43227;
														assign node43227 = (inp[0]) ? 4'b1011 : node43228;
															assign node43228 = (inp[15]) ? 4'b1001 : 4'b1011;
														assign node43232 = (inp[10]) ? 4'b1001 : node43233;
															assign node43233 = (inp[0]) ? node43237 : node43234;
																assign node43234 = (inp[15]) ? 4'b1011 : 4'b1001;
																assign node43237 = (inp[15]) ? 4'b1001 : 4'b1011;
													assign node43241 = (inp[15]) ? 4'b1001 : node43242;
														assign node43242 = (inp[10]) ? 4'b1001 : node43243;
															assign node43243 = (inp[3]) ? node43247 : node43244;
																assign node43244 = (inp[0]) ? 4'b1001 : 4'b1011;
																assign node43247 = (inp[0]) ? 4'b1011 : 4'b1001;
										assign node43252 = (inp[12]) ? node43296 : node43253;
											assign node43253 = (inp[10]) ? node43273 : node43254;
												assign node43254 = (inp[15]) ? node43262 : node43255;
													assign node43255 = (inp[0]) ? 4'b1001 : node43256;
														assign node43256 = (inp[5]) ? node43258 : 4'b1011;
															assign node43258 = (inp[3]) ? 4'b1001 : 4'b1011;
													assign node43262 = (inp[0]) ? node43268 : node43263;
														assign node43263 = (inp[5]) ? node43265 : 4'b1001;
															assign node43265 = (inp[3]) ? 4'b1011 : 4'b1001;
														assign node43268 = (inp[5]) ? node43270 : 4'b1011;
															assign node43270 = (inp[3]) ? 4'b1001 : 4'b1011;
												assign node43273 = (inp[0]) ? node43285 : node43274;
													assign node43274 = (inp[15]) ? node43280 : node43275;
														assign node43275 = (inp[5]) ? 4'b1101 : node43276;
															assign node43276 = (inp[3]) ? 4'b1101 : 4'b1111;
														assign node43280 = (inp[3]) ? 4'b1111 : node43281;
															assign node43281 = (inp[5]) ? 4'b1111 : 4'b1101;
													assign node43285 = (inp[15]) ? node43291 : node43286;
														assign node43286 = (inp[5]) ? 4'b1111 : node43287;
															assign node43287 = (inp[3]) ? 4'b1111 : 4'b1101;
														assign node43291 = (inp[3]) ? 4'b1101 : node43292;
															assign node43292 = (inp[5]) ? 4'b1101 : 4'b1111;
											assign node43296 = (inp[10]) ? node43336 : node43297;
												assign node43297 = (inp[14]) ? node43321 : node43298;
													assign node43298 = (inp[15]) ? node43310 : node43299;
														assign node43299 = (inp[0]) ? node43305 : node43300;
															assign node43300 = (inp[5]) ? 4'b1101 : node43301;
																assign node43301 = (inp[3]) ? 4'b1101 : 4'b1111;
															assign node43305 = (inp[5]) ? 4'b1111 : node43306;
																assign node43306 = (inp[3]) ? 4'b1111 : 4'b1101;
														assign node43310 = (inp[0]) ? node43316 : node43311;
															assign node43311 = (inp[5]) ? 4'b1111 : node43312;
																assign node43312 = (inp[3]) ? 4'b1111 : 4'b1101;
															assign node43316 = (inp[5]) ? 4'b1101 : node43317;
																assign node43317 = (inp[3]) ? 4'b1101 : 4'b1111;
													assign node43321 = (inp[0]) ? node43329 : node43322;
														assign node43322 = (inp[15]) ? node43324 : 4'b1101;
															assign node43324 = (inp[3]) ? 4'b1111 : node43325;
																assign node43325 = (inp[5]) ? 4'b1111 : 4'b1101;
														assign node43329 = (inp[15]) ? 4'b1101 : node43330;
															assign node43330 = (inp[3]) ? 4'b1111 : node43331;
																assign node43331 = (inp[5]) ? 4'b1111 : 4'b1101;
												assign node43336 = (inp[5]) ? node43358 : node43337;
													assign node43337 = (inp[0]) ? node43351 : node43338;
														assign node43338 = (inp[14]) ? node43344 : node43339;
															assign node43339 = (inp[15]) ? 4'b1101 : node43340;
																assign node43340 = (inp[3]) ? 4'b1101 : 4'b1111;
															assign node43344 = (inp[15]) ? node43348 : node43345;
																assign node43345 = (inp[3]) ? 4'b1101 : 4'b1111;
																assign node43348 = (inp[3]) ? 4'b1111 : 4'b1101;
														assign node43351 = (inp[3]) ? node43355 : node43352;
															assign node43352 = (inp[15]) ? 4'b1111 : 4'b1101;
															assign node43355 = (inp[15]) ? 4'b1101 : 4'b1111;
													assign node43358 = (inp[0]) ? node43362 : node43359;
														assign node43359 = (inp[15]) ? 4'b1111 : 4'b1101;
														assign node43362 = (inp[15]) ? 4'b1101 : 4'b1111;
									assign node43365 = (inp[4]) ? node43491 : node43366;
										assign node43366 = (inp[10]) ? node43436 : node43367;
											assign node43367 = (inp[12]) ? node43409 : node43368;
												assign node43368 = (inp[14]) ? node43392 : node43369;
													assign node43369 = (inp[0]) ? node43381 : node43370;
														assign node43370 = (inp[15]) ? node43376 : node43371;
															assign node43371 = (inp[3]) ? node43373 : 4'b1011;
																assign node43373 = (inp[5]) ? 4'b1001 : 4'b1011;
															assign node43376 = (inp[3]) ? node43378 : 4'b1001;
																assign node43378 = (inp[5]) ? 4'b1011 : 4'b1001;
														assign node43381 = (inp[15]) ? node43387 : node43382;
															assign node43382 = (inp[3]) ? node43384 : 4'b1001;
																assign node43384 = (inp[5]) ? 4'b1011 : 4'b1001;
															assign node43387 = (inp[5]) ? node43389 : 4'b1011;
																assign node43389 = (inp[3]) ? 4'b1001 : 4'b1011;
													assign node43392 = (inp[5]) ? node43398 : node43393;
														assign node43393 = (inp[3]) ? 4'b1001 : node43394;
															assign node43394 = (inp[0]) ? 4'b1001 : 4'b1011;
														assign node43398 = (inp[0]) ? node43404 : node43399;
															assign node43399 = (inp[15]) ? 4'b1001 : node43400;
																assign node43400 = (inp[3]) ? 4'b1001 : 4'b1011;
															assign node43404 = (inp[3]) ? 4'b1011 : node43405;
																assign node43405 = (inp[15]) ? 4'b1011 : 4'b1001;
												assign node43409 = (inp[5]) ? node43429 : node43410;
													assign node43410 = (inp[14]) ? node43422 : node43411;
														assign node43411 = (inp[15]) ? node43417 : node43412;
															assign node43412 = (inp[3]) ? node43414 : 4'b1101;
																assign node43414 = (inp[0]) ? 4'b1111 : 4'b1101;
															assign node43417 = (inp[0]) ? node43419 : 4'b1111;
																assign node43419 = (inp[3]) ? 4'b1101 : 4'b1111;
														assign node43422 = (inp[15]) ? 4'b1111 : node43423;
															assign node43423 = (inp[3]) ? node43425 : 4'b1111;
																assign node43425 = (inp[0]) ? 4'b1111 : 4'b1101;
													assign node43429 = (inp[0]) ? node43433 : node43430;
														assign node43430 = (inp[15]) ? 4'b1111 : 4'b1101;
														assign node43433 = (inp[15]) ? 4'b1101 : 4'b1111;
											assign node43436 = (inp[3]) ? node43476 : node43437;
												assign node43437 = (inp[5]) ? node43453 : node43438;
													assign node43438 = (inp[14]) ? node43446 : node43439;
														assign node43439 = (inp[0]) ? node43443 : node43440;
															assign node43440 = (inp[15]) ? 4'b1101 : 4'b1111;
															assign node43443 = (inp[15]) ? 4'b1111 : 4'b1101;
														assign node43446 = (inp[12]) ? node43448 : 4'b1101;
															assign node43448 = (inp[0]) ? 4'b1101 : node43449;
																assign node43449 = (inp[15]) ? 4'b1101 : 4'b1111;
													assign node43453 = (inp[14]) ? node43461 : node43454;
														assign node43454 = (inp[15]) ? node43458 : node43455;
															assign node43455 = (inp[0]) ? 4'b1111 : 4'b1101;
															assign node43458 = (inp[0]) ? 4'b1101 : 4'b1111;
														assign node43461 = (inp[12]) ? node43469 : node43462;
															assign node43462 = (inp[0]) ? node43466 : node43463;
																assign node43463 = (inp[15]) ? 4'b1111 : 4'b1101;
																assign node43466 = (inp[15]) ? 4'b1101 : 4'b1111;
															assign node43469 = (inp[0]) ? node43473 : node43470;
																assign node43470 = (inp[15]) ? 4'b1111 : 4'b1101;
																assign node43473 = (inp[15]) ? 4'b1101 : 4'b1111;
												assign node43476 = (inp[5]) ? node43484 : node43477;
													assign node43477 = (inp[15]) ? node43481 : node43478;
														assign node43478 = (inp[0]) ? 4'b1111 : 4'b1101;
														assign node43481 = (inp[0]) ? 4'b1101 : 4'b1111;
													assign node43484 = (inp[0]) ? node43488 : node43485;
														assign node43485 = (inp[15]) ? 4'b1111 : 4'b1101;
														assign node43488 = (inp[15]) ? 4'b1101 : 4'b1111;
										assign node43491 = (inp[10]) ? node43553 : node43492;
											assign node43492 = (inp[12]) ? node43514 : node43493;
												assign node43493 = (inp[15]) ? node43503 : node43494;
													assign node43494 = (inp[0]) ? node43500 : node43495;
														assign node43495 = (inp[3]) ? 4'b1101 : node43496;
															assign node43496 = (inp[5]) ? 4'b1101 : 4'b1111;
														assign node43500 = (inp[5]) ? 4'b1111 : 4'b1101;
													assign node43503 = (inp[0]) ? node43509 : node43504;
														assign node43504 = (inp[3]) ? 4'b1111 : node43505;
															assign node43505 = (inp[5]) ? 4'b1111 : 4'b1101;
														assign node43509 = (inp[3]) ? 4'b1101 : node43510;
															assign node43510 = (inp[5]) ? 4'b1101 : 4'b1111;
												assign node43514 = (inp[14]) ? node43538 : node43515;
													assign node43515 = (inp[5]) ? node43531 : node43516;
														assign node43516 = (inp[3]) ? node43524 : node43517;
															assign node43517 = (inp[0]) ? node43521 : node43518;
																assign node43518 = (inp[15]) ? 4'b1001 : 4'b1011;
																assign node43521 = (inp[15]) ? 4'b1011 : 4'b1001;
															assign node43524 = (inp[15]) ? node43528 : node43525;
																assign node43525 = (inp[0]) ? 4'b1011 : 4'b1001;
																assign node43528 = (inp[0]) ? 4'b1001 : 4'b1011;
														assign node43531 = (inp[15]) ? node43535 : node43532;
															assign node43532 = (inp[0]) ? 4'b1011 : 4'b1001;
															assign node43535 = (inp[0]) ? 4'b1001 : 4'b1011;
													assign node43538 = (inp[5]) ? node43546 : node43539;
														assign node43539 = (inp[0]) ? node43541 : 4'b1001;
															assign node43541 = (inp[3]) ? 4'b1001 : node43542;
																assign node43542 = (inp[15]) ? 4'b1011 : 4'b1001;
														assign node43546 = (inp[15]) ? node43550 : node43547;
															assign node43547 = (inp[0]) ? 4'b1011 : 4'b1001;
															assign node43550 = (inp[0]) ? 4'b1001 : 4'b1011;
											assign node43553 = (inp[3]) ? node43595 : node43554;
												assign node43554 = (inp[14]) ? node43574 : node43555;
													assign node43555 = (inp[12]) ? node43565 : node43556;
														assign node43556 = (inp[0]) ? 4'b1001 : node43557;
															assign node43557 = (inp[5]) ? node43561 : node43558;
																assign node43558 = (inp[15]) ? 4'b1001 : 4'b1011;
																assign node43561 = (inp[15]) ? 4'b1011 : 4'b1001;
														assign node43565 = (inp[5]) ? 4'b1011 : node43566;
															assign node43566 = (inp[0]) ? node43570 : node43567;
																assign node43567 = (inp[15]) ? 4'b1001 : 4'b1011;
																assign node43570 = (inp[15]) ? 4'b1011 : 4'b1001;
													assign node43574 = (inp[12]) ? node43586 : node43575;
														assign node43575 = (inp[5]) ? node43581 : node43576;
															assign node43576 = (inp[15]) ? node43578 : 4'b1011;
																assign node43578 = (inp[0]) ? 4'b1011 : 4'b1001;
															assign node43581 = (inp[15]) ? node43583 : 4'b1001;
																assign node43583 = (inp[0]) ? 4'b1001 : 4'b1011;
														assign node43586 = (inp[0]) ? node43588 : 4'b1001;
															assign node43588 = (inp[5]) ? node43592 : node43589;
																assign node43589 = (inp[15]) ? 4'b1011 : 4'b1001;
																assign node43592 = (inp[15]) ? 4'b1001 : 4'b1011;
												assign node43595 = (inp[0]) ? node43599 : node43596;
													assign node43596 = (inp[15]) ? 4'b1011 : 4'b1001;
													assign node43599 = (inp[15]) ? 4'b1001 : 4'b1011;
						assign node43602 = (inp[7]) ? node44512 : node43603;
							assign node43603 = (inp[2]) ? node44163 : node43604;
								assign node43604 = (inp[14]) ? node43910 : node43605;
									assign node43605 = (inp[15]) ? node43777 : node43606;
										assign node43606 = (inp[12]) ? node43684 : node43607;
											assign node43607 = (inp[10]) ? node43659 : node43608;
												assign node43608 = (inp[0]) ? node43636 : node43609;
													assign node43609 = (inp[3]) ? node43623 : node43610;
														assign node43610 = (inp[5]) ? node43618 : node43611;
															assign node43611 = (inp[4]) ? node43615 : node43612;
																assign node43612 = (inp[9]) ? 4'b0010 : 4'b0110;
																assign node43615 = (inp[9]) ? 4'b0110 : 4'b0010;
															assign node43618 = (inp[9]) ? 4'b0010 : node43619;
																assign node43619 = (inp[4]) ? 4'b0010 : 4'b0110;
														assign node43623 = (inp[5]) ? node43631 : node43624;
															assign node43624 = (inp[4]) ? node43628 : node43625;
																assign node43625 = (inp[9]) ? 4'b0010 : 4'b0110;
																assign node43628 = (inp[9]) ? 4'b0100 : 4'b0010;
															assign node43631 = (inp[4]) ? node43633 : 4'b0000;
																assign node43633 = (inp[9]) ? 4'b0100 : 4'b0000;
													assign node43636 = (inp[3]) ? node43646 : node43637;
														assign node43637 = (inp[5]) ? node43639 : 4'b0100;
															assign node43639 = (inp[4]) ? node43643 : node43640;
																assign node43640 = (inp[9]) ? 4'b0000 : 4'b0100;
																assign node43643 = (inp[9]) ? 4'b0110 : 4'b0000;
														assign node43646 = (inp[5]) ? node43652 : node43647;
															assign node43647 = (inp[4]) ? node43649 : 4'b0000;
																assign node43649 = (inp[9]) ? 4'b0110 : 4'b0000;
															assign node43652 = (inp[4]) ? node43656 : node43653;
																assign node43653 = (inp[9]) ? 4'b0010 : 4'b0110;
																assign node43656 = (inp[9]) ? 4'b0110 : 4'b0010;
												assign node43659 = (inp[4]) ? node43675 : node43660;
													assign node43660 = (inp[9]) ? node43668 : node43661;
														assign node43661 = (inp[0]) ? node43663 : 4'b0110;
															assign node43663 = (inp[3]) ? node43665 : 4'b0100;
																assign node43665 = (inp[5]) ? 4'b0110 : 4'b0100;
														assign node43668 = (inp[5]) ? node43670 : 4'b0000;
															assign node43670 = (inp[3]) ? node43672 : 4'b0010;
																assign node43672 = (inp[0]) ? 4'b0010 : 4'b0000;
													assign node43675 = (inp[9]) ? node43681 : node43676;
														assign node43676 = (inp[0]) ? 4'b0000 : node43677;
															assign node43677 = (inp[5]) ? 4'b0000 : 4'b0010;
														assign node43681 = (inp[0]) ? 4'b0110 : 4'b0100;
											assign node43684 = (inp[3]) ? node43738 : node43685;
												assign node43685 = (inp[0]) ? node43713 : node43686;
													assign node43686 = (inp[5]) ? node43702 : node43687;
														assign node43687 = (inp[9]) ? node43695 : node43688;
															assign node43688 = (inp[4]) ? node43692 : node43689;
																assign node43689 = (inp[10]) ? 4'b0010 : 4'b0110;
																assign node43692 = (inp[10]) ? 4'b0110 : 4'b0010;
															assign node43695 = (inp[4]) ? node43699 : node43696;
																assign node43696 = (inp[10]) ? 4'b0110 : 4'b0010;
																assign node43699 = (inp[10]) ? 4'b0010 : 4'b0110;
														assign node43702 = (inp[4]) ? node43708 : node43703;
															assign node43703 = (inp[10]) ? 4'b0010 : node43704;
																assign node43704 = (inp[9]) ? 4'b0010 : 4'b0110;
															assign node43708 = (inp[9]) ? node43710 : 4'b0100;
																assign node43710 = (inp[10]) ? 4'b0000 : 4'b0100;
													assign node43713 = (inp[5]) ? node43725 : node43714;
														assign node43714 = (inp[4]) ? node43720 : node43715;
															assign node43715 = (inp[10]) ? 4'b0100 : node43716;
																assign node43716 = (inp[9]) ? 4'b0000 : 4'b0100;
															assign node43720 = (inp[9]) ? 4'b0000 : node43721;
																assign node43721 = (inp[10]) ? 4'b0100 : 4'b0000;
														assign node43725 = (inp[4]) ? node43733 : node43726;
															assign node43726 = (inp[10]) ? node43730 : node43727;
																assign node43727 = (inp[9]) ? 4'b0000 : 4'b0100;
																assign node43730 = (inp[9]) ? 4'b0110 : 4'b0000;
															assign node43733 = (inp[9]) ? node43735 : 4'b0110;
																assign node43735 = (inp[10]) ? 4'b0010 : 4'b0110;
												assign node43738 = (inp[0]) ? node43752 : node43739;
													assign node43739 = (inp[4]) ? 4'b0100 : node43740;
														assign node43740 = (inp[5]) ? node43746 : node43741;
															assign node43741 = (inp[9]) ? 4'b0100 : node43742;
																assign node43742 = (inp[10]) ? 4'b0010 : 4'b0110;
															assign node43746 = (inp[9]) ? node43748 : 4'b0000;
																assign node43748 = (inp[10]) ? 4'b0100 : 4'b0000;
													assign node43752 = (inp[5]) ? node43762 : node43753;
														assign node43753 = (inp[9]) ? node43757 : node43754;
															assign node43754 = (inp[10]) ? 4'b0110 : 4'b0100;
															assign node43757 = (inp[4]) ? node43759 : 4'b0110;
																assign node43759 = (inp[10]) ? 4'b0010 : 4'b0110;
														assign node43762 = (inp[9]) ? node43770 : node43763;
															assign node43763 = (inp[4]) ? node43767 : node43764;
																assign node43764 = (inp[10]) ? 4'b0010 : 4'b0110;
																assign node43767 = (inp[10]) ? 4'b0110 : 4'b0010;
															assign node43770 = (inp[10]) ? node43774 : node43771;
																assign node43771 = (inp[4]) ? 4'b0110 : 4'b0010;
																assign node43774 = (inp[4]) ? 4'b0010 : 4'b0110;
										assign node43777 = (inp[0]) ? node43845 : node43778;
											assign node43778 = (inp[3]) ? node43816 : node43779;
												assign node43779 = (inp[5]) ? node43799 : node43780;
													assign node43780 = (inp[9]) ? node43792 : node43781;
														assign node43781 = (inp[4]) ? node43787 : node43782;
															assign node43782 = (inp[10]) ? node43784 : 4'b0100;
																assign node43784 = (inp[12]) ? 4'b0000 : 4'b0100;
															assign node43787 = (inp[12]) ? node43789 : 4'b0000;
																assign node43789 = (inp[10]) ? 4'b0100 : 4'b0000;
														assign node43792 = (inp[4]) ? 4'b0100 : node43793;
															assign node43793 = (inp[12]) ? node43795 : 4'b0000;
																assign node43795 = (inp[10]) ? 4'b0100 : 4'b0000;
													assign node43799 = (inp[4]) ? node43811 : node43800;
														assign node43800 = (inp[9]) ? node43806 : node43801;
															assign node43801 = (inp[10]) ? node43803 : 4'b0100;
																assign node43803 = (inp[12]) ? 4'b0000 : 4'b0100;
															assign node43806 = (inp[12]) ? node43808 : 4'b0000;
																assign node43808 = (inp[10]) ? 4'b0110 : 4'b0000;
														assign node43811 = (inp[12]) ? 4'b0110 : node43812;
															assign node43812 = (inp[9]) ? 4'b0110 : 4'b0000;
												assign node43816 = (inp[5]) ? node43834 : node43817;
													assign node43817 = (inp[9]) ? node43825 : node43818;
														assign node43818 = (inp[4]) ? 4'b0000 : node43819;
															assign node43819 = (inp[10]) ? node43821 : 4'b0100;
																assign node43821 = (inp[12]) ? 4'b0000 : 4'b0100;
														assign node43825 = (inp[4]) ? node43829 : node43826;
															assign node43826 = (inp[10]) ? 4'b0110 : 4'b0000;
															assign node43829 = (inp[10]) ? node43831 : 4'b0110;
																assign node43831 = (inp[12]) ? 4'b0010 : 4'b0110;
													assign node43834 = (inp[9]) ? node43840 : node43835;
														assign node43835 = (inp[12]) ? node43837 : 4'b0010;
															assign node43837 = (inp[4]) ? 4'b0110 : 4'b0010;
														assign node43840 = (inp[10]) ? 4'b0110 : node43841;
															assign node43841 = (inp[4]) ? 4'b0110 : 4'b0010;
											assign node43845 = (inp[3]) ? node43873 : node43846;
												assign node43846 = (inp[5]) ? node43862 : node43847;
													assign node43847 = (inp[12]) ? node43855 : node43848;
														assign node43848 = (inp[9]) ? node43852 : node43849;
															assign node43849 = (inp[4]) ? 4'b0010 : 4'b0110;
															assign node43852 = (inp[4]) ? 4'b0110 : 4'b0010;
														assign node43855 = (inp[10]) ? node43857 : 4'b0010;
															assign node43857 = (inp[4]) ? 4'b0010 : node43858;
																assign node43858 = (inp[9]) ? 4'b0110 : 4'b0010;
													assign node43862 = (inp[9]) ? node43866 : node43863;
														assign node43863 = (inp[4]) ? 4'b0010 : 4'b0110;
														assign node43866 = (inp[4]) ? node43870 : node43867;
															assign node43867 = (inp[12]) ? 4'b0100 : 4'b0010;
															assign node43870 = (inp[10]) ? 4'b0000 : 4'b0100;
												assign node43873 = (inp[5]) ? node43891 : node43874;
													assign node43874 = (inp[9]) ? node43882 : node43875;
														assign node43875 = (inp[10]) ? node43877 : 4'b0010;
															assign node43877 = (inp[4]) ? 4'b0100 : node43878;
																assign node43878 = (inp[12]) ? 4'b0010 : 4'b0110;
														assign node43882 = (inp[4]) ? node43886 : node43883;
															assign node43883 = (inp[10]) ? 4'b0100 : 4'b0010;
															assign node43886 = (inp[12]) ? node43888 : 4'b0100;
																assign node43888 = (inp[10]) ? 4'b0000 : 4'b0100;
													assign node43891 = (inp[10]) ? node43899 : node43892;
														assign node43892 = (inp[9]) ? node43896 : node43893;
															assign node43893 = (inp[4]) ? 4'b0000 : 4'b0100;
															assign node43896 = (inp[4]) ? 4'b0100 : 4'b0000;
														assign node43899 = (inp[12]) ? node43905 : node43900;
															assign node43900 = (inp[9]) ? 4'b0000 : node43901;
																assign node43901 = (inp[4]) ? 4'b0000 : 4'b0100;
															assign node43905 = (inp[9]) ? node43907 : 4'b0100;
																assign node43907 = (inp[4]) ? 4'b0000 : 4'b0100;
									assign node43910 = (inp[4]) ? node44030 : node43911;
										assign node43911 = (inp[9]) ? node43973 : node43912;
											assign node43912 = (inp[10]) ? node43942 : node43913;
												assign node43913 = (inp[12]) ? node43927 : node43914;
													assign node43914 = (inp[5]) ? node43920 : node43915;
														assign node43915 = (inp[0]) ? node43917 : 4'b1111;
															assign node43917 = (inp[15]) ? 4'b1111 : 4'b1101;
														assign node43920 = (inp[15]) ? 4'b1101 : node43921;
															assign node43921 = (inp[0]) ? 4'b1111 : node43922;
																assign node43922 = (inp[3]) ? 4'b1101 : 4'b1111;
													assign node43927 = (inp[0]) ? node43933 : node43928;
														assign node43928 = (inp[15]) ? node43930 : 4'b1011;
															assign node43930 = (inp[3]) ? 4'b1011 : 4'b1001;
														assign node43933 = (inp[15]) ? node43939 : node43934;
															assign node43934 = (inp[5]) ? node43936 : 4'b1001;
																assign node43936 = (inp[3]) ? 4'b1011 : 4'b1001;
															assign node43939 = (inp[3]) ? 4'b1001 : 4'b1011;
												assign node43942 = (inp[12]) ? node43956 : node43943;
													assign node43943 = (inp[0]) ? node43945 : 4'b1011;
														assign node43945 = (inp[15]) ? node43951 : node43946;
															assign node43946 = (inp[5]) ? node43948 : 4'b1001;
																assign node43948 = (inp[3]) ? 4'b1011 : 4'b1001;
															assign node43951 = (inp[3]) ? node43953 : 4'b1011;
																assign node43953 = (inp[5]) ? 4'b1001 : 4'b1011;
													assign node43956 = (inp[15]) ? node43964 : node43957;
														assign node43957 = (inp[0]) ? 4'b1001 : node43958;
															assign node43958 = (inp[5]) ? node43960 : 4'b1011;
																assign node43960 = (inp[3]) ? 4'b1001 : 4'b1011;
														assign node43964 = (inp[0]) ? node43970 : node43965;
															assign node43965 = (inp[5]) ? node43967 : 4'b1001;
																assign node43967 = (inp[3]) ? 4'b1011 : 4'b1001;
															assign node43970 = (inp[3]) ? 4'b1001 : 4'b1011;
											assign node43973 = (inp[10]) ? node44001 : node43974;
												assign node43974 = (inp[12]) ? node43984 : node43975;
													assign node43975 = (inp[15]) ? 4'b1011 : node43976;
														assign node43976 = (inp[0]) ? node43978 : 4'b1011;
															assign node43978 = (inp[3]) ? node43980 : 4'b1001;
																assign node43980 = (inp[5]) ? 4'b1011 : 4'b1001;
													assign node43984 = (inp[3]) ? node43994 : node43985;
														assign node43985 = (inp[15]) ? node43987 : 4'b1111;
															assign node43987 = (inp[0]) ? node43991 : node43988;
																assign node43988 = (inp[5]) ? 4'b1111 : 4'b1101;
																assign node43991 = (inp[5]) ? 4'b1101 : 4'b1111;
														assign node43994 = (inp[0]) ? node43998 : node43995;
															assign node43995 = (inp[15]) ? 4'b1111 : 4'b1101;
															assign node43998 = (inp[15]) ? 4'b1101 : 4'b1111;
												assign node44001 = (inp[3]) ? node44023 : node44002;
													assign node44002 = (inp[0]) ? node44010 : node44003;
														assign node44003 = (inp[5]) ? node44007 : node44004;
															assign node44004 = (inp[15]) ? 4'b1101 : 4'b1111;
															assign node44007 = (inp[15]) ? 4'b1111 : 4'b1101;
														assign node44010 = (inp[12]) ? node44016 : node44011;
															assign node44011 = (inp[15]) ? 4'b1111 : node44012;
																assign node44012 = (inp[5]) ? 4'b1111 : 4'b1101;
															assign node44016 = (inp[5]) ? node44020 : node44017;
																assign node44017 = (inp[15]) ? 4'b1111 : 4'b1101;
																assign node44020 = (inp[15]) ? 4'b1101 : 4'b1111;
													assign node44023 = (inp[0]) ? node44027 : node44024;
														assign node44024 = (inp[15]) ? 4'b1111 : 4'b1101;
														assign node44027 = (inp[15]) ? 4'b1101 : 4'b1111;
										assign node44030 = (inp[9]) ? node44092 : node44031;
											assign node44031 = (inp[10]) ? node44067 : node44032;
												assign node44032 = (inp[12]) ? node44056 : node44033;
													assign node44033 = (inp[3]) ? node44047 : node44034;
														assign node44034 = (inp[5]) ? node44040 : node44035;
															assign node44035 = (inp[15]) ? node44037 : 4'b1001;
																assign node44037 = (inp[0]) ? 4'b1011 : 4'b1001;
															assign node44040 = (inp[15]) ? node44044 : node44041;
																assign node44041 = (inp[0]) ? 4'b1001 : 4'b1011;
																assign node44044 = (inp[0]) ? 4'b1011 : 4'b1001;
														assign node44047 = (inp[0]) ? 4'b1011 : node44048;
															assign node44048 = (inp[15]) ? node44052 : node44049;
																assign node44049 = (inp[5]) ? 4'b1001 : 4'b1011;
																assign node44052 = (inp[5]) ? 4'b1011 : 4'b1001;
													assign node44056 = (inp[5]) ? node44060 : node44057;
														assign node44057 = (inp[3]) ? 4'b1111 : 4'b1101;
														assign node44060 = (inp[0]) ? node44064 : node44061;
															assign node44061 = (inp[15]) ? 4'b1111 : 4'b1101;
															assign node44064 = (inp[15]) ? 4'b1101 : 4'b1111;
												assign node44067 = (inp[5]) ? node44085 : node44068;
													assign node44068 = (inp[3]) ? node44078 : node44069;
														assign node44069 = (inp[12]) ? node44075 : node44070;
															assign node44070 = (inp[15]) ? node44072 : 4'b1111;
																assign node44072 = (inp[0]) ? 4'b1111 : 4'b1101;
															assign node44075 = (inp[15]) ? 4'b1111 : 4'b1101;
														assign node44078 = (inp[15]) ? node44082 : node44079;
															assign node44079 = (inp[0]) ? 4'b1111 : 4'b1101;
															assign node44082 = (inp[0]) ? 4'b1101 : 4'b1111;
													assign node44085 = (inp[15]) ? node44089 : node44086;
														assign node44086 = (inp[0]) ? 4'b1111 : 4'b1101;
														assign node44089 = (inp[0]) ? 4'b1101 : 4'b1111;
											assign node44092 = (inp[12]) ? node44128 : node44093;
												assign node44093 = (inp[10]) ? node44107 : node44094;
													assign node44094 = (inp[3]) ? node44100 : node44095;
														assign node44095 = (inp[15]) ? node44097 : 4'b1111;
															assign node44097 = (inp[5]) ? 4'b1101 : 4'b1111;
														assign node44100 = (inp[15]) ? node44104 : node44101;
															assign node44101 = (inp[0]) ? 4'b1111 : 4'b1101;
															assign node44104 = (inp[0]) ? 4'b1101 : 4'b1111;
													assign node44107 = (inp[15]) ? node44119 : node44108;
														assign node44108 = (inp[0]) ? node44114 : node44109;
															assign node44109 = (inp[3]) ? 4'b1001 : node44110;
																assign node44110 = (inp[5]) ? 4'b1001 : 4'b1011;
															assign node44114 = (inp[3]) ? 4'b1011 : node44115;
																assign node44115 = (inp[5]) ? 4'b1011 : 4'b1001;
														assign node44119 = (inp[0]) ? node44125 : node44120;
															assign node44120 = (inp[5]) ? 4'b1011 : node44121;
																assign node44121 = (inp[3]) ? 4'b1011 : 4'b1001;
															assign node44125 = (inp[5]) ? 4'b1001 : 4'b1011;
												assign node44128 = (inp[10]) ? node44150 : node44129;
													assign node44129 = (inp[0]) ? node44139 : node44130;
														assign node44130 = (inp[15]) ? node44134 : node44131;
															assign node44131 = (inp[5]) ? 4'b1001 : 4'b1011;
															assign node44134 = (inp[3]) ? 4'b1011 : node44135;
																assign node44135 = (inp[5]) ? 4'b1011 : 4'b1001;
														assign node44139 = (inp[15]) ? node44145 : node44140;
															assign node44140 = (inp[3]) ? 4'b1011 : node44141;
																assign node44141 = (inp[5]) ? 4'b1011 : 4'b1001;
															assign node44145 = (inp[3]) ? 4'b1001 : node44146;
																assign node44146 = (inp[5]) ? 4'b1001 : 4'b1011;
													assign node44150 = (inp[15]) ? node44158 : node44151;
														assign node44151 = (inp[0]) ? node44153 : 4'b1001;
															assign node44153 = (inp[3]) ? 4'b1011 : node44154;
																assign node44154 = (inp[5]) ? 4'b1011 : 4'b1001;
														assign node44158 = (inp[0]) ? node44160 : 4'b1011;
															assign node44160 = (inp[5]) ? 4'b1001 : 4'b1011;
								assign node44163 = (inp[15]) ? node44305 : node44164;
									assign node44164 = (inp[4]) ? node44232 : node44165;
										assign node44165 = (inp[9]) ? node44197 : node44166;
											assign node44166 = (inp[10]) ? node44186 : node44167;
												assign node44167 = (inp[12]) ? node44179 : node44168;
													assign node44168 = (inp[0]) ? node44174 : node44169;
														assign node44169 = (inp[3]) ? node44171 : 4'b1111;
															assign node44171 = (inp[5]) ? 4'b1101 : 4'b1111;
														assign node44174 = (inp[3]) ? node44176 : 4'b1101;
															assign node44176 = (inp[5]) ? 4'b1111 : 4'b1101;
													assign node44179 = (inp[0]) ? 4'b1001 : node44180;
														assign node44180 = (inp[3]) ? node44182 : 4'b1011;
															assign node44182 = (inp[5]) ? 4'b1001 : 4'b1011;
												assign node44186 = (inp[0]) ? node44192 : node44187;
													assign node44187 = (inp[5]) ? node44189 : 4'b1011;
														assign node44189 = (inp[3]) ? 4'b1001 : 4'b1011;
													assign node44192 = (inp[5]) ? node44194 : 4'b1001;
														assign node44194 = (inp[3]) ? 4'b1011 : 4'b1001;
											assign node44197 = (inp[10]) ? node44221 : node44198;
												assign node44198 = (inp[12]) ? node44210 : node44199;
													assign node44199 = (inp[0]) ? node44205 : node44200;
														assign node44200 = (inp[3]) ? node44202 : 4'b1011;
															assign node44202 = (inp[5]) ? 4'b1001 : 4'b1011;
														assign node44205 = (inp[5]) ? node44207 : 4'b1001;
															assign node44207 = (inp[3]) ? 4'b1011 : 4'b1001;
													assign node44210 = (inp[0]) ? node44216 : node44211;
														assign node44211 = (inp[5]) ? 4'b1101 : node44212;
															assign node44212 = (inp[3]) ? 4'b1101 : 4'b1111;
														assign node44216 = (inp[5]) ? 4'b1111 : node44217;
															assign node44217 = (inp[3]) ? 4'b1111 : 4'b1101;
												assign node44221 = (inp[0]) ? node44227 : node44222;
													assign node44222 = (inp[3]) ? 4'b1101 : node44223;
														assign node44223 = (inp[5]) ? 4'b1101 : 4'b1111;
													assign node44227 = (inp[5]) ? 4'b1111 : node44228;
														assign node44228 = (inp[3]) ? 4'b1111 : 4'b1101;
										assign node44232 = (inp[9]) ? node44270 : node44233;
											assign node44233 = (inp[12]) ? node44259 : node44234;
												assign node44234 = (inp[10]) ? node44242 : node44235;
													assign node44235 = (inp[0]) ? node44237 : 4'b1011;
														assign node44237 = (inp[5]) ? node44239 : 4'b1001;
															assign node44239 = (inp[3]) ? 4'b1011 : 4'b1001;
													assign node44242 = (inp[14]) ? node44248 : node44243;
														assign node44243 = (inp[0]) ? 4'b1101 : node44244;
															assign node44244 = (inp[5]) ? 4'b1101 : 4'b1111;
														assign node44248 = (inp[0]) ? node44254 : node44249;
															assign node44249 = (inp[3]) ? 4'b1101 : node44250;
																assign node44250 = (inp[5]) ? 4'b1101 : 4'b1111;
															assign node44254 = (inp[3]) ? 4'b1111 : node44255;
																assign node44255 = (inp[5]) ? 4'b1111 : 4'b1101;
												assign node44259 = (inp[0]) ? node44265 : node44260;
													assign node44260 = (inp[3]) ? 4'b1101 : node44261;
														assign node44261 = (inp[5]) ? 4'b1101 : 4'b1111;
													assign node44265 = (inp[3]) ? 4'b1111 : node44266;
														assign node44266 = (inp[5]) ? 4'b1111 : 4'b1101;
											assign node44270 = (inp[10]) ? node44294 : node44271;
												assign node44271 = (inp[12]) ? node44281 : node44272;
													assign node44272 = (inp[0]) ? node44276 : node44273;
														assign node44273 = (inp[5]) ? 4'b1101 : 4'b1111;
														assign node44276 = (inp[5]) ? 4'b1111 : node44277;
															assign node44277 = (inp[3]) ? 4'b1111 : 4'b1101;
													assign node44281 = (inp[14]) ? node44289 : node44282;
														assign node44282 = (inp[5]) ? node44286 : node44283;
															assign node44283 = (inp[0]) ? 4'b1001 : 4'b1011;
															assign node44286 = (inp[0]) ? 4'b1011 : 4'b1001;
														assign node44289 = (inp[0]) ? 4'b1011 : node44290;
															assign node44290 = (inp[5]) ? 4'b1001 : 4'b1011;
												assign node44294 = (inp[0]) ? node44300 : node44295;
													assign node44295 = (inp[5]) ? 4'b1001 : node44296;
														assign node44296 = (inp[3]) ? 4'b1001 : 4'b1011;
													assign node44300 = (inp[5]) ? 4'b1011 : node44301;
														assign node44301 = (inp[3]) ? 4'b1011 : 4'b1001;
									assign node44305 = (inp[0]) ? node44407 : node44306;
										assign node44306 = (inp[3]) ? node44354 : node44307;
											assign node44307 = (inp[5]) ? node44331 : node44308;
												assign node44308 = (inp[12]) ? node44324 : node44309;
													assign node44309 = (inp[4]) ? node44317 : node44310;
														assign node44310 = (inp[9]) ? node44314 : node44311;
															assign node44311 = (inp[10]) ? 4'b1001 : 4'b1101;
															assign node44314 = (inp[10]) ? 4'b1101 : 4'b1001;
														assign node44317 = (inp[10]) ? node44321 : node44318;
															assign node44318 = (inp[9]) ? 4'b1101 : 4'b1001;
															assign node44321 = (inp[9]) ? 4'b1001 : 4'b1101;
													assign node44324 = (inp[9]) ? node44328 : node44325;
														assign node44325 = (inp[4]) ? 4'b1101 : 4'b1001;
														assign node44328 = (inp[4]) ? 4'b1001 : 4'b1101;
												assign node44331 = (inp[9]) ? node44343 : node44332;
													assign node44332 = (inp[4]) ? node44338 : node44333;
														assign node44333 = (inp[10]) ? 4'b1001 : node44334;
															assign node44334 = (inp[12]) ? 4'b1001 : 4'b1101;
														assign node44338 = (inp[12]) ? 4'b1111 : node44339;
															assign node44339 = (inp[10]) ? 4'b1111 : 4'b1001;
													assign node44343 = (inp[4]) ? node44349 : node44344;
														assign node44344 = (inp[12]) ? 4'b1111 : node44345;
															assign node44345 = (inp[10]) ? 4'b1111 : 4'b1001;
														assign node44349 = (inp[12]) ? 4'b1011 : node44350;
															assign node44350 = (inp[10]) ? 4'b1011 : 4'b1111;
											assign node44354 = (inp[5]) ? node44374 : node44355;
												assign node44355 = (inp[9]) ? node44367 : node44356;
													assign node44356 = (inp[4]) ? node44362 : node44357;
														assign node44357 = (inp[10]) ? 4'b1001 : node44358;
															assign node44358 = (inp[12]) ? 4'b1001 : 4'b1101;
														assign node44362 = (inp[10]) ? 4'b1111 : node44363;
															assign node44363 = (inp[12]) ? 4'b1111 : 4'b1001;
													assign node44367 = (inp[4]) ? node44369 : 4'b1111;
														assign node44369 = (inp[10]) ? 4'b1011 : node44370;
															assign node44370 = (inp[12]) ? 4'b1011 : 4'b1111;
												assign node44374 = (inp[12]) ? node44394 : node44375;
													assign node44375 = (inp[10]) ? node44389 : node44376;
														assign node44376 = (inp[14]) ? node44382 : node44377;
															assign node44377 = (inp[4]) ? node44379 : 4'b1111;
																assign node44379 = (inp[9]) ? 4'b1111 : 4'b1011;
															assign node44382 = (inp[9]) ? node44386 : node44383;
																assign node44383 = (inp[4]) ? 4'b1011 : 4'b1111;
																assign node44386 = (inp[4]) ? 4'b1111 : 4'b1011;
														assign node44389 = (inp[4]) ? 4'b1111 : node44390;
															assign node44390 = (inp[9]) ? 4'b1111 : 4'b1011;
													assign node44394 = (inp[14]) ? node44402 : node44395;
														assign node44395 = (inp[10]) ? node44397 : 4'b1011;
															assign node44397 = (inp[9]) ? 4'b1011 : node44398;
																assign node44398 = (inp[4]) ? 4'b1111 : 4'b1011;
														assign node44402 = (inp[9]) ? 4'b1111 : node44403;
															assign node44403 = (inp[4]) ? 4'b1111 : 4'b1011;
										assign node44407 = (inp[5]) ? node44459 : node44408;
											assign node44408 = (inp[3]) ? node44442 : node44409;
												assign node44409 = (inp[14]) ? node44423 : node44410;
													assign node44410 = (inp[9]) ? node44418 : node44411;
														assign node44411 = (inp[4]) ? node44413 : 4'b1011;
															assign node44413 = (inp[10]) ? 4'b1111 : node44414;
																assign node44414 = (inp[12]) ? 4'b1111 : 4'b1011;
														assign node44418 = (inp[4]) ? node44420 : 4'b1111;
															assign node44420 = (inp[12]) ? 4'b1011 : 4'b1111;
													assign node44423 = (inp[9]) ? node44433 : node44424;
														assign node44424 = (inp[4]) ? node44428 : node44425;
															assign node44425 = (inp[10]) ? 4'b1011 : 4'b1111;
															assign node44428 = (inp[12]) ? 4'b1111 : node44429;
																assign node44429 = (inp[10]) ? 4'b1111 : 4'b1011;
														assign node44433 = (inp[12]) ? 4'b1011 : node44434;
															assign node44434 = (inp[4]) ? node44438 : node44435;
																assign node44435 = (inp[10]) ? 4'b1111 : 4'b1011;
																assign node44438 = (inp[10]) ? 4'b1011 : 4'b1111;
												assign node44442 = (inp[9]) ? node44452 : node44443;
													assign node44443 = (inp[4]) ? node44449 : node44444;
														assign node44444 = (inp[12]) ? 4'b1011 : node44445;
															assign node44445 = (inp[10]) ? 4'b1011 : 4'b1111;
														assign node44449 = (inp[12]) ? 4'b1101 : 4'b1011;
													assign node44452 = (inp[4]) ? 4'b1001 : node44453;
														assign node44453 = (inp[10]) ? 4'b1101 : node44454;
															assign node44454 = (inp[12]) ? 4'b1101 : 4'b1011;
											assign node44459 = (inp[3]) ? node44481 : node44460;
												assign node44460 = (inp[4]) ? node44470 : node44461;
													assign node44461 = (inp[9]) ? node44467 : node44462;
														assign node44462 = (inp[10]) ? 4'b1011 : node44463;
															assign node44463 = (inp[12]) ? 4'b1011 : 4'b1111;
														assign node44467 = (inp[12]) ? 4'b1101 : 4'b1011;
													assign node44470 = (inp[9]) ? node44476 : node44471;
														assign node44471 = (inp[12]) ? 4'b1101 : node44472;
															assign node44472 = (inp[10]) ? 4'b1101 : 4'b1011;
														assign node44476 = (inp[12]) ? 4'b1001 : node44477;
															assign node44477 = (inp[14]) ? 4'b1101 : 4'b1001;
												assign node44481 = (inp[14]) ? node44497 : node44482;
													assign node44482 = (inp[4]) ? node44486 : node44483;
														assign node44483 = (inp[9]) ? 4'b1101 : 4'b1001;
														assign node44486 = (inp[9]) ? node44492 : node44487;
															assign node44487 = (inp[10]) ? 4'b1101 : node44488;
																assign node44488 = (inp[12]) ? 4'b1101 : 4'b1001;
															assign node44492 = (inp[12]) ? 4'b1001 : node44493;
																assign node44493 = (inp[10]) ? 4'b1001 : 4'b1101;
													assign node44497 = (inp[10]) ? 4'b1001 : node44498;
														assign node44498 = (inp[9]) ? node44506 : node44499;
															assign node44499 = (inp[12]) ? node44503 : node44500;
																assign node44500 = (inp[4]) ? 4'b1001 : 4'b1101;
																assign node44503 = (inp[4]) ? 4'b1101 : 4'b1001;
															assign node44506 = (inp[12]) ? node44508 : 4'b1101;
																assign node44508 = (inp[4]) ? 4'b1001 : 4'b1101;
							assign node44512 = (inp[14]) ? node45050 : node44513;
								assign node44513 = (inp[2]) ? node44783 : node44514;
									assign node44514 = (inp[0]) ? node44630 : node44515;
										assign node44515 = (inp[10]) ? node44589 : node44516;
											assign node44516 = (inp[4]) ? node44564 : node44517;
												assign node44517 = (inp[15]) ? node44539 : node44518;
													assign node44518 = (inp[3]) ? node44532 : node44519;
														assign node44519 = (inp[5]) ? node44527 : node44520;
															assign node44520 = (inp[12]) ? node44524 : node44521;
																assign node44521 = (inp[9]) ? 4'b1011 : 4'b1111;
																assign node44524 = (inp[9]) ? 4'b1111 : 4'b1011;
															assign node44527 = (inp[9]) ? 4'b1101 : node44528;
																assign node44528 = (inp[12]) ? 4'b1011 : 4'b1111;
														assign node44532 = (inp[12]) ? node44536 : node44533;
															assign node44533 = (inp[5]) ? 4'b1001 : 4'b1011;
															assign node44536 = (inp[9]) ? 4'b1101 : 4'b1001;
													assign node44539 = (inp[5]) ? node44549 : node44540;
														assign node44540 = (inp[3]) ? node44546 : node44541;
															assign node44541 = (inp[9]) ? 4'b1101 : node44542;
																assign node44542 = (inp[12]) ? 4'b1001 : 4'b1101;
															assign node44546 = (inp[9]) ? 4'b1001 : 4'b1101;
														assign node44549 = (inp[3]) ? node44557 : node44550;
															assign node44550 = (inp[9]) ? node44554 : node44551;
																assign node44551 = (inp[12]) ? 4'b1001 : 4'b1101;
																assign node44554 = (inp[12]) ? 4'b1111 : 4'b1001;
															assign node44557 = (inp[12]) ? node44561 : node44558;
																assign node44558 = (inp[9]) ? 4'b1011 : 4'b1111;
																assign node44561 = (inp[9]) ? 4'b1111 : 4'b1011;
												assign node44564 = (inp[12]) ? node44572 : node44565;
													assign node44565 = (inp[9]) ? 4'b1101 : node44566;
														assign node44566 = (inp[15]) ? 4'b1001 : node44567;
															assign node44567 = (inp[5]) ? 4'b1001 : 4'b1011;
													assign node44572 = (inp[9]) ? node44582 : node44573;
														assign node44573 = (inp[5]) ? node44579 : node44574;
															assign node44574 = (inp[3]) ? 4'b1101 : node44575;
																assign node44575 = (inp[15]) ? 4'b1101 : 4'b1111;
															assign node44579 = (inp[15]) ? 4'b1111 : 4'b1101;
														assign node44582 = (inp[15]) ? 4'b1011 : node44583;
															assign node44583 = (inp[3]) ? 4'b1001 : node44584;
																assign node44584 = (inp[5]) ? 4'b1001 : 4'b1011;
											assign node44589 = (inp[15]) ? node44613 : node44590;
												assign node44590 = (inp[3]) ? node44600 : node44591;
													assign node44591 = (inp[9]) ? node44595 : node44592;
														assign node44592 = (inp[4]) ? 4'b1111 : 4'b1011;
														assign node44595 = (inp[5]) ? 4'b1101 : node44596;
															assign node44596 = (inp[4]) ? 4'b1011 : 4'b1111;
													assign node44600 = (inp[5]) ? node44606 : node44601;
														assign node44601 = (inp[4]) ? node44603 : 4'b1011;
															assign node44603 = (inp[9]) ? 4'b1001 : 4'b1101;
														assign node44606 = (inp[4]) ? node44610 : node44607;
															assign node44607 = (inp[9]) ? 4'b1101 : 4'b1001;
															assign node44610 = (inp[9]) ? 4'b1001 : 4'b1101;
												assign node44613 = (inp[9]) ? node44625 : node44614;
													assign node44614 = (inp[4]) ? node44620 : node44615;
														assign node44615 = (inp[3]) ? node44617 : 4'b1001;
															assign node44617 = (inp[5]) ? 4'b1011 : 4'b1001;
														assign node44620 = (inp[5]) ? 4'b1111 : node44621;
															assign node44621 = (inp[3]) ? 4'b1111 : 4'b1101;
													assign node44625 = (inp[4]) ? 4'b1011 : node44626;
														assign node44626 = (inp[3]) ? 4'b1111 : 4'b1101;
										assign node44630 = (inp[15]) ? node44706 : node44631;
											assign node44631 = (inp[3]) ? node44667 : node44632;
												assign node44632 = (inp[5]) ? node44652 : node44633;
													assign node44633 = (inp[9]) ? node44643 : node44634;
														assign node44634 = (inp[4]) ? node44640 : node44635;
															assign node44635 = (inp[12]) ? 4'b1001 : node44636;
																assign node44636 = (inp[10]) ? 4'b1001 : 4'b1101;
															assign node44640 = (inp[12]) ? 4'b1101 : 4'b1001;
														assign node44643 = (inp[12]) ? 4'b1101 : node44644;
															assign node44644 = (inp[4]) ? node44648 : node44645;
																assign node44645 = (inp[10]) ? 4'b1101 : 4'b1001;
																assign node44648 = (inp[10]) ? 4'b1001 : 4'b1101;
													assign node44652 = (inp[9]) ? node44660 : node44653;
														assign node44653 = (inp[4]) ? 4'b1111 : node44654;
															assign node44654 = (inp[12]) ? 4'b1001 : node44655;
																assign node44655 = (inp[10]) ? 4'b1001 : 4'b1101;
														assign node44660 = (inp[4]) ? node44662 : 4'b1111;
															assign node44662 = (inp[10]) ? 4'b1011 : node44663;
																assign node44663 = (inp[12]) ? 4'b1011 : 4'b1111;
												assign node44667 = (inp[5]) ? node44687 : node44668;
													assign node44668 = (inp[4]) ? node44676 : node44669;
														assign node44669 = (inp[9]) ? node44671 : 4'b1001;
															assign node44671 = (inp[10]) ? 4'b1111 : node44672;
																assign node44672 = (inp[12]) ? 4'b1111 : 4'b1001;
														assign node44676 = (inp[9]) ? node44682 : node44677;
															assign node44677 = (inp[10]) ? 4'b1111 : node44678;
																assign node44678 = (inp[12]) ? 4'b1111 : 4'b1001;
															assign node44682 = (inp[12]) ? 4'b1011 : node44683;
																assign node44683 = (inp[10]) ? 4'b1011 : 4'b1111;
													assign node44687 = (inp[9]) ? node44697 : node44688;
														assign node44688 = (inp[4]) ? node44694 : node44689;
															assign node44689 = (inp[12]) ? 4'b1011 : node44690;
																assign node44690 = (inp[10]) ? 4'b1011 : 4'b1111;
															assign node44694 = (inp[12]) ? 4'b1111 : 4'b1011;
														assign node44697 = (inp[10]) ? 4'b1111 : node44698;
															assign node44698 = (inp[4]) ? node44702 : node44699;
																assign node44699 = (inp[12]) ? 4'b1111 : 4'b1011;
																assign node44702 = (inp[12]) ? 4'b1011 : 4'b1111;
											assign node44706 = (inp[5]) ? node44746 : node44707;
												assign node44707 = (inp[3]) ? node44731 : node44708;
													assign node44708 = (inp[12]) ? node44718 : node44709;
														assign node44709 = (inp[9]) ? node44711 : 4'b1111;
															assign node44711 = (inp[10]) ? node44715 : node44712;
																assign node44712 = (inp[4]) ? 4'b1111 : 4'b1011;
																assign node44715 = (inp[4]) ? 4'b1011 : 4'b1111;
														assign node44718 = (inp[10]) ? node44726 : node44719;
															assign node44719 = (inp[9]) ? node44723 : node44720;
																assign node44720 = (inp[4]) ? 4'b1111 : 4'b1011;
																assign node44723 = (inp[4]) ? 4'b1011 : 4'b1111;
															assign node44726 = (inp[9]) ? 4'b1011 : node44727;
																assign node44727 = (inp[4]) ? 4'b1111 : 4'b1011;
													assign node44731 = (inp[4]) ? node44741 : node44732;
														assign node44732 = (inp[9]) ? node44738 : node44733;
															assign node44733 = (inp[10]) ? 4'b1011 : node44734;
																assign node44734 = (inp[12]) ? 4'b1011 : 4'b1111;
															assign node44738 = (inp[12]) ? 4'b1101 : 4'b1011;
														assign node44741 = (inp[10]) ? node44743 : 4'b1101;
															assign node44743 = (inp[9]) ? 4'b1001 : 4'b1101;
												assign node44746 = (inp[3]) ? node44768 : node44747;
													assign node44747 = (inp[12]) ? node44761 : node44748;
														assign node44748 = (inp[10]) ? node44754 : node44749;
															assign node44749 = (inp[4]) ? 4'b1011 : node44750;
																assign node44750 = (inp[9]) ? 4'b1011 : 4'b1111;
															assign node44754 = (inp[9]) ? node44758 : node44755;
																assign node44755 = (inp[4]) ? 4'b1101 : 4'b1011;
																assign node44758 = (inp[4]) ? 4'b1001 : 4'b1101;
														assign node44761 = (inp[9]) ? node44765 : node44762;
															assign node44762 = (inp[4]) ? 4'b1101 : 4'b1011;
															assign node44765 = (inp[4]) ? 4'b1001 : 4'b1101;
													assign node44768 = (inp[9]) ? node44772 : node44769;
														assign node44769 = (inp[4]) ? 4'b1101 : 4'b1001;
														assign node44772 = (inp[4]) ? node44778 : node44773;
															assign node44773 = (inp[10]) ? 4'b1101 : node44774;
																assign node44774 = (inp[12]) ? 4'b1101 : 4'b1001;
															assign node44778 = (inp[10]) ? 4'b1001 : node44779;
																assign node44779 = (inp[12]) ? 4'b1001 : 4'b1101;
									assign node44783 = (inp[9]) ? node44925 : node44784;
										assign node44784 = (inp[4]) ? node44848 : node44785;
											assign node44785 = (inp[10]) ? node44823 : node44786;
												assign node44786 = (inp[12]) ? node44808 : node44787;
													assign node44787 = (inp[0]) ? node44797 : node44788;
														assign node44788 = (inp[5]) ? node44790 : 4'b1110;
															assign node44790 = (inp[3]) ? node44794 : node44791;
																assign node44791 = (inp[15]) ? 4'b1100 : 4'b1110;
																assign node44794 = (inp[15]) ? 4'b1110 : 4'b1100;
														assign node44797 = (inp[15]) ? node44803 : node44798;
															assign node44798 = (inp[3]) ? node44800 : 4'b1100;
																assign node44800 = (inp[5]) ? 4'b1110 : 4'b1100;
															assign node44803 = (inp[3]) ? node44805 : 4'b1110;
																assign node44805 = (inp[5]) ? 4'b1100 : 4'b1110;
													assign node44808 = (inp[15]) ? node44818 : node44809;
														assign node44809 = (inp[5]) ? node44811 : 4'b1010;
															assign node44811 = (inp[3]) ? node44815 : node44812;
																assign node44812 = (inp[0]) ? 4'b1000 : 4'b1010;
																assign node44815 = (inp[0]) ? 4'b1010 : 4'b1000;
														assign node44818 = (inp[5]) ? node44820 : 4'b1000;
															assign node44820 = (inp[3]) ? 4'b1010 : 4'b1000;
												assign node44823 = (inp[12]) ? node44833 : node44824;
													assign node44824 = (inp[15]) ? node44826 : 4'b1010;
														assign node44826 = (inp[0]) ? node44828 : 4'b1000;
															assign node44828 = (inp[3]) ? node44830 : 4'b1010;
																assign node44830 = (inp[5]) ? 4'b1000 : 4'b1010;
													assign node44833 = (inp[3]) ? node44841 : node44834;
														assign node44834 = (inp[15]) ? node44838 : node44835;
															assign node44835 = (inp[0]) ? 4'b1000 : 4'b1010;
															assign node44838 = (inp[0]) ? 4'b1010 : 4'b1000;
														assign node44841 = (inp[5]) ? 4'b1010 : node44842;
															assign node44842 = (inp[15]) ? node44844 : 4'b1010;
																assign node44844 = (inp[0]) ? 4'b1010 : 4'b1000;
											assign node44848 = (inp[10]) ? node44888 : node44849;
												assign node44849 = (inp[12]) ? node44871 : node44850;
													assign node44850 = (inp[5]) ? node44858 : node44851;
														assign node44851 = (inp[3]) ? node44853 : 4'b1010;
															assign node44853 = (inp[15]) ? node44855 : 4'b1000;
																assign node44855 = (inp[0]) ? 4'b1010 : 4'b1000;
														assign node44858 = (inp[0]) ? node44866 : node44859;
															assign node44859 = (inp[15]) ? node44863 : node44860;
																assign node44860 = (inp[3]) ? 4'b1000 : 4'b1010;
																assign node44863 = (inp[3]) ? 4'b1010 : 4'b1000;
															assign node44866 = (inp[15]) ? 4'b1000 : node44867;
																assign node44867 = (inp[3]) ? 4'b1010 : 4'b1000;
													assign node44871 = (inp[15]) ? node44879 : node44872;
														assign node44872 = (inp[0]) ? 4'b1110 : node44873;
															assign node44873 = (inp[3]) ? 4'b1100 : node44874;
																assign node44874 = (inp[5]) ? 4'b1100 : 4'b1110;
														assign node44879 = (inp[3]) ? 4'b1100 : node44880;
															assign node44880 = (inp[0]) ? node44884 : node44881;
																assign node44881 = (inp[5]) ? 4'b1110 : 4'b1100;
																assign node44884 = (inp[5]) ? 4'b1100 : 4'b1110;
												assign node44888 = (inp[3]) ? node44912 : node44889;
													assign node44889 = (inp[0]) ? node44905 : node44890;
														assign node44890 = (inp[12]) ? node44898 : node44891;
															assign node44891 = (inp[15]) ? node44895 : node44892;
																assign node44892 = (inp[5]) ? 4'b1100 : 4'b1110;
																assign node44895 = (inp[5]) ? 4'b1110 : 4'b1100;
															assign node44898 = (inp[5]) ? node44902 : node44899;
																assign node44899 = (inp[15]) ? 4'b1100 : 4'b1110;
																assign node44902 = (inp[15]) ? 4'b1110 : 4'b1100;
														assign node44905 = (inp[15]) ? node44909 : node44906;
															assign node44906 = (inp[5]) ? 4'b1110 : 4'b1100;
															assign node44909 = (inp[5]) ? 4'b1100 : 4'b1110;
													assign node44912 = (inp[5]) ? node44920 : node44913;
														assign node44913 = (inp[0]) ? node44917 : node44914;
															assign node44914 = (inp[15]) ? 4'b1110 : 4'b1100;
															assign node44917 = (inp[15]) ? 4'b1100 : 4'b1110;
														assign node44920 = (inp[0]) ? 4'b1110 : node44921;
															assign node44921 = (inp[15]) ? 4'b1110 : 4'b1100;
										assign node44925 = (inp[4]) ? node44999 : node44926;
											assign node44926 = (inp[12]) ? node44964 : node44927;
												assign node44927 = (inp[10]) ? node44949 : node44928;
													assign node44928 = (inp[3]) ? node44938 : node44929;
														assign node44929 = (inp[5]) ? 4'b1000 : node44930;
															assign node44930 = (inp[0]) ? node44934 : node44931;
																assign node44931 = (inp[15]) ? 4'b1000 : 4'b1010;
																assign node44934 = (inp[15]) ? 4'b1010 : 4'b1000;
														assign node44938 = (inp[5]) ? node44944 : node44939;
															assign node44939 = (inp[0]) ? 4'b1000 : node44940;
																assign node44940 = (inp[15]) ? 4'b1000 : 4'b1010;
															assign node44944 = (inp[0]) ? 4'b1010 : node44945;
																assign node44945 = (inp[15]) ? 4'b1010 : 4'b1000;
													assign node44949 = (inp[0]) ? node44959 : node44950;
														assign node44950 = (inp[15]) ? node44954 : node44951;
															assign node44951 = (inp[5]) ? 4'b1100 : 4'b1110;
															assign node44954 = (inp[5]) ? 4'b1110 : node44955;
																assign node44955 = (inp[3]) ? 4'b1110 : 4'b1100;
														assign node44959 = (inp[15]) ? node44961 : 4'b1110;
															assign node44961 = (inp[3]) ? 4'b1100 : 4'b1110;
												assign node44964 = (inp[10]) ? node44986 : node44965;
													assign node44965 = (inp[15]) ? node44977 : node44966;
														assign node44966 = (inp[0]) ? node44972 : node44967;
															assign node44967 = (inp[5]) ? 4'b1100 : node44968;
																assign node44968 = (inp[3]) ? 4'b1100 : 4'b1110;
															assign node44972 = (inp[3]) ? 4'b1110 : node44973;
																assign node44973 = (inp[5]) ? 4'b1110 : 4'b1100;
														assign node44977 = (inp[0]) ? node44981 : node44978;
															assign node44978 = (inp[5]) ? 4'b1110 : 4'b1100;
															assign node44981 = (inp[3]) ? 4'b1100 : node44982;
																assign node44982 = (inp[5]) ? 4'b1100 : 4'b1110;
													assign node44986 = (inp[5]) ? 4'b1100 : node44987;
														assign node44987 = (inp[3]) ? node44993 : node44988;
															assign node44988 = (inp[15]) ? 4'b1100 : node44989;
																assign node44989 = (inp[0]) ? 4'b1100 : 4'b1110;
															assign node44993 = (inp[15]) ? 4'b1110 : node44994;
																assign node44994 = (inp[0]) ? 4'b1110 : 4'b1100;
											assign node44999 = (inp[10]) ? node45029 : node45000;
												assign node45000 = (inp[12]) ? node45012 : node45001;
													assign node45001 = (inp[5]) ? node45007 : node45002;
														assign node45002 = (inp[0]) ? node45004 : 4'b1100;
															assign node45004 = (inp[3]) ? 4'b1100 : 4'b1110;
														assign node45007 = (inp[0]) ? node45009 : 4'b1110;
															assign node45009 = (inp[15]) ? 4'b1100 : 4'b1110;
													assign node45012 = (inp[0]) ? node45024 : node45013;
														assign node45013 = (inp[15]) ? node45019 : node45014;
															assign node45014 = (inp[3]) ? 4'b1000 : node45015;
																assign node45015 = (inp[5]) ? 4'b1000 : 4'b1010;
															assign node45019 = (inp[5]) ? 4'b1010 : node45020;
																assign node45020 = (inp[3]) ? 4'b1010 : 4'b1000;
														assign node45024 = (inp[15]) ? 4'b1000 : node45025;
															assign node45025 = (inp[3]) ? 4'b1010 : 4'b1000;
												assign node45029 = (inp[3]) ? node45043 : node45030;
													assign node45030 = (inp[5]) ? node45038 : node45031;
														assign node45031 = (inp[12]) ? 4'b1000 : node45032;
															assign node45032 = (inp[15]) ? 4'b1010 : node45033;
																assign node45033 = (inp[0]) ? 4'b1000 : 4'b1010;
														assign node45038 = (inp[0]) ? 4'b1010 : node45039;
															assign node45039 = (inp[15]) ? 4'b1010 : 4'b1000;
													assign node45043 = (inp[0]) ? node45047 : node45044;
														assign node45044 = (inp[15]) ? 4'b1010 : 4'b1000;
														assign node45047 = (inp[15]) ? 4'b1000 : 4'b1010;
								assign node45050 = (inp[15]) ? node45250 : node45051;
									assign node45051 = (inp[0]) ? node45157 : node45052;
										assign node45052 = (inp[5]) ? node45098 : node45053;
											assign node45053 = (inp[3]) ? node45079 : node45054;
												assign node45054 = (inp[12]) ? node45070 : node45055;
													assign node45055 = (inp[9]) ? node45063 : node45056;
														assign node45056 = (inp[4]) ? node45060 : node45057;
															assign node45057 = (inp[10]) ? 4'b1010 : 4'b1110;
															assign node45060 = (inp[10]) ? 4'b1110 : 4'b1010;
														assign node45063 = (inp[10]) ? node45067 : node45064;
															assign node45064 = (inp[4]) ? 4'b1110 : 4'b1010;
															assign node45067 = (inp[4]) ? 4'b1010 : 4'b1110;
													assign node45070 = (inp[10]) ? node45072 : 4'b1110;
														assign node45072 = (inp[9]) ? node45076 : node45073;
															assign node45073 = (inp[4]) ? 4'b1110 : 4'b1010;
															assign node45076 = (inp[4]) ? 4'b1010 : 4'b1110;
												assign node45079 = (inp[9]) ? node45091 : node45080;
													assign node45080 = (inp[4]) ? node45086 : node45081;
														assign node45081 = (inp[10]) ? 4'b1010 : node45082;
															assign node45082 = (inp[2]) ? 4'b1110 : 4'b1010;
														assign node45086 = (inp[12]) ? 4'b1100 : node45087;
															assign node45087 = (inp[10]) ? 4'b1100 : 4'b1010;
													assign node45091 = (inp[4]) ? node45093 : 4'b1100;
														assign node45093 = (inp[10]) ? 4'b1000 : node45094;
															assign node45094 = (inp[12]) ? 4'b1000 : 4'b1100;
											assign node45098 = (inp[3]) ? node45122 : node45099;
												assign node45099 = (inp[9]) ? node45111 : node45100;
													assign node45100 = (inp[4]) ? node45106 : node45101;
														assign node45101 = (inp[12]) ? 4'b1010 : node45102;
															assign node45102 = (inp[10]) ? 4'b1010 : 4'b1110;
														assign node45106 = (inp[12]) ? 4'b1100 : node45107;
															assign node45107 = (inp[10]) ? 4'b1100 : 4'b1010;
													assign node45111 = (inp[4]) ? node45117 : node45112;
														assign node45112 = (inp[10]) ? 4'b1100 : node45113;
															assign node45113 = (inp[12]) ? 4'b1100 : 4'b1010;
														assign node45117 = (inp[10]) ? 4'b1000 : node45118;
															assign node45118 = (inp[12]) ? 4'b1000 : 4'b1100;
												assign node45122 = (inp[2]) ? node45136 : node45123;
													assign node45123 = (inp[12]) ? node45131 : node45124;
														assign node45124 = (inp[10]) ? 4'b1100 : node45125;
															assign node45125 = (inp[4]) ? 4'b1000 : node45126;
																assign node45126 = (inp[9]) ? 4'b1000 : 4'b1100;
														assign node45131 = (inp[4]) ? node45133 : 4'b1000;
															assign node45133 = (inp[9]) ? 4'b1000 : 4'b1100;
													assign node45136 = (inp[12]) ? node45152 : node45137;
														assign node45137 = (inp[4]) ? node45145 : node45138;
															assign node45138 = (inp[10]) ? node45142 : node45139;
																assign node45139 = (inp[9]) ? 4'b1000 : 4'b1100;
																assign node45142 = (inp[9]) ? 4'b1100 : 4'b1000;
															assign node45145 = (inp[10]) ? node45149 : node45146;
																assign node45146 = (inp[9]) ? 4'b1100 : 4'b1000;
																assign node45149 = (inp[9]) ? 4'b1000 : 4'b1100;
														assign node45152 = (inp[4]) ? node45154 : 4'b1100;
															assign node45154 = (inp[9]) ? 4'b1000 : 4'b1100;
										assign node45157 = (inp[5]) ? node45203 : node45158;
											assign node45158 = (inp[3]) ? node45180 : node45159;
												assign node45159 = (inp[10]) ? node45173 : node45160;
													assign node45160 = (inp[12]) ? node45166 : node45161;
														assign node45161 = (inp[9]) ? node45163 : 4'b1100;
															assign node45163 = (inp[4]) ? 4'b1100 : 4'b1000;
														assign node45166 = (inp[9]) ? node45170 : node45167;
															assign node45167 = (inp[4]) ? 4'b1100 : 4'b1000;
															assign node45170 = (inp[4]) ? 4'b1000 : 4'b1100;
													assign node45173 = (inp[4]) ? node45177 : node45174;
														assign node45174 = (inp[9]) ? 4'b1100 : 4'b1000;
														assign node45177 = (inp[9]) ? 4'b1000 : 4'b1100;
												assign node45180 = (inp[9]) ? node45192 : node45181;
													assign node45181 = (inp[4]) ? node45187 : node45182;
														assign node45182 = (inp[10]) ? 4'b1000 : node45183;
															assign node45183 = (inp[12]) ? 4'b1000 : 4'b1100;
														assign node45187 = (inp[10]) ? 4'b1110 : node45188;
															assign node45188 = (inp[12]) ? 4'b1110 : 4'b1000;
													assign node45192 = (inp[4]) ? node45198 : node45193;
														assign node45193 = (inp[12]) ? 4'b1110 : node45194;
															assign node45194 = (inp[10]) ? 4'b1110 : 4'b1000;
														assign node45198 = (inp[12]) ? 4'b1010 : node45199;
															assign node45199 = (inp[10]) ? 4'b1010 : 4'b1110;
											assign node45203 = (inp[3]) ? node45227 : node45204;
												assign node45204 = (inp[4]) ? node45216 : node45205;
													assign node45205 = (inp[9]) ? node45211 : node45206;
														assign node45206 = (inp[12]) ? 4'b1000 : node45207;
															assign node45207 = (inp[10]) ? 4'b1000 : 4'b1100;
														assign node45211 = (inp[12]) ? 4'b1110 : node45212;
															assign node45212 = (inp[10]) ? 4'b1110 : 4'b1000;
													assign node45216 = (inp[9]) ? node45222 : node45217;
														assign node45217 = (inp[12]) ? 4'b1110 : node45218;
															assign node45218 = (inp[10]) ? 4'b1110 : 4'b1000;
														assign node45222 = (inp[12]) ? 4'b1010 : node45223;
															assign node45223 = (inp[10]) ? 4'b1010 : 4'b1110;
												assign node45227 = (inp[4]) ? node45239 : node45228;
													assign node45228 = (inp[9]) ? node45234 : node45229;
														assign node45229 = (inp[10]) ? 4'b1010 : node45230;
															assign node45230 = (inp[12]) ? 4'b1010 : 4'b1110;
														assign node45234 = (inp[12]) ? 4'b1110 : node45235;
															assign node45235 = (inp[10]) ? 4'b1110 : 4'b1010;
													assign node45239 = (inp[9]) ? node45245 : node45240;
														assign node45240 = (inp[12]) ? 4'b1110 : node45241;
															assign node45241 = (inp[10]) ? 4'b1110 : 4'b1010;
														assign node45245 = (inp[12]) ? 4'b1010 : node45246;
															assign node45246 = (inp[10]) ? 4'b1010 : 4'b1110;
									assign node45250 = (inp[2]) ? node45392 : node45251;
										assign node45251 = (inp[0]) ? node45331 : node45252;
											assign node45252 = (inp[3]) ? node45296 : node45253;
												assign node45253 = (inp[5]) ? node45279 : node45254;
													assign node45254 = (inp[10]) ? node45270 : node45255;
														assign node45255 = (inp[9]) ? node45263 : node45256;
															assign node45256 = (inp[12]) ? node45260 : node45257;
																assign node45257 = (inp[4]) ? 4'b1000 : 4'b1100;
																assign node45260 = (inp[4]) ? 4'b1100 : 4'b1000;
															assign node45263 = (inp[12]) ? node45267 : node45264;
																assign node45264 = (inp[4]) ? 4'b1100 : 4'b1000;
																assign node45267 = (inp[4]) ? 4'b1000 : 4'b1100;
														assign node45270 = (inp[12]) ? node45276 : node45271;
															assign node45271 = (inp[9]) ? 4'b1000 : node45272;
																assign node45272 = (inp[4]) ? 4'b1100 : 4'b1000;
															assign node45276 = (inp[4]) ? 4'b1000 : 4'b1100;
													assign node45279 = (inp[9]) ? node45287 : node45280;
														assign node45280 = (inp[4]) ? node45282 : 4'b1000;
															assign node45282 = (inp[10]) ? 4'b1110 : node45283;
																assign node45283 = (inp[12]) ? 4'b1110 : 4'b1000;
														assign node45287 = (inp[4]) ? node45293 : node45288;
															assign node45288 = (inp[12]) ? 4'b1110 : node45289;
																assign node45289 = (inp[10]) ? 4'b1110 : 4'b1000;
															assign node45293 = (inp[10]) ? 4'b1010 : 4'b1110;
												assign node45296 = (inp[5]) ? node45314 : node45297;
													assign node45297 = (inp[9]) ? node45303 : node45298;
														assign node45298 = (inp[12]) ? 4'b1000 : node45299;
															assign node45299 = (inp[10]) ? 4'b1110 : 4'b1100;
														assign node45303 = (inp[4]) ? node45309 : node45304;
															assign node45304 = (inp[10]) ? 4'b1110 : node45305;
																assign node45305 = (inp[12]) ? 4'b1110 : 4'b1000;
															assign node45309 = (inp[10]) ? 4'b1010 : node45310;
																assign node45310 = (inp[12]) ? 4'b1010 : 4'b1110;
													assign node45314 = (inp[10]) ? node45324 : node45315;
														assign node45315 = (inp[12]) ? 4'b1110 : node45316;
															assign node45316 = (inp[9]) ? node45320 : node45317;
																assign node45317 = (inp[4]) ? 4'b1010 : 4'b1110;
																assign node45320 = (inp[4]) ? 4'b1110 : 4'b1010;
														assign node45324 = (inp[9]) ? node45328 : node45325;
															assign node45325 = (inp[4]) ? 4'b1110 : 4'b1010;
															assign node45328 = (inp[4]) ? 4'b1010 : 4'b1110;
											assign node45331 = (inp[3]) ? node45365 : node45332;
												assign node45332 = (inp[5]) ? node45346 : node45333;
													assign node45333 = (inp[10]) ? node45341 : node45334;
														assign node45334 = (inp[4]) ? 4'b1110 : node45335;
															assign node45335 = (inp[12]) ? 4'b1010 : node45336;
																assign node45336 = (inp[9]) ? 4'b1010 : 4'b1110;
														assign node45341 = (inp[4]) ? 4'b1010 : node45342;
															assign node45342 = (inp[9]) ? 4'b1110 : 4'b1010;
													assign node45346 = (inp[4]) ? node45356 : node45347;
														assign node45347 = (inp[9]) ? node45351 : node45348;
															assign node45348 = (inp[10]) ? 4'b1010 : 4'b1110;
															assign node45351 = (inp[10]) ? 4'b1100 : node45352;
																assign node45352 = (inp[12]) ? 4'b1100 : 4'b1010;
														assign node45356 = (inp[12]) ? 4'b1100 : node45357;
															assign node45357 = (inp[10]) ? node45361 : node45358;
																assign node45358 = (inp[9]) ? 4'b1100 : 4'b1010;
																assign node45361 = (inp[9]) ? 4'b1000 : 4'b1100;
												assign node45365 = (inp[9]) ? node45381 : node45366;
													assign node45366 = (inp[4]) ? node45374 : node45367;
														assign node45367 = (inp[5]) ? 4'b1000 : node45368;
															assign node45368 = (inp[10]) ? 4'b1010 : node45369;
																assign node45369 = (inp[12]) ? 4'b1010 : 4'b1110;
														assign node45374 = (inp[10]) ? 4'b1100 : node45375;
															assign node45375 = (inp[12]) ? 4'b1100 : node45376;
																assign node45376 = (inp[5]) ? 4'b1000 : 4'b1010;
													assign node45381 = (inp[4]) ? node45387 : node45382;
														assign node45382 = (inp[10]) ? 4'b1100 : node45383;
															assign node45383 = (inp[12]) ? 4'b1100 : 4'b1000;
														assign node45387 = (inp[12]) ? 4'b1000 : node45388;
															assign node45388 = (inp[10]) ? 4'b1000 : 4'b1100;
										assign node45392 = (inp[3]) ? node45466 : node45393;
											assign node45393 = (inp[0]) ? node45433 : node45394;
												assign node45394 = (inp[5]) ? node45418 : node45395;
													assign node45395 = (inp[10]) ? node45411 : node45396;
														assign node45396 = (inp[9]) ? node45404 : node45397;
															assign node45397 = (inp[4]) ? node45401 : node45398;
																assign node45398 = (inp[12]) ? 4'b1000 : 4'b1100;
																assign node45401 = (inp[12]) ? 4'b1100 : 4'b1000;
															assign node45404 = (inp[4]) ? node45408 : node45405;
																assign node45405 = (inp[12]) ? 4'b1100 : 4'b1000;
																assign node45408 = (inp[12]) ? 4'b1000 : 4'b1100;
														assign node45411 = (inp[4]) ? node45415 : node45412;
															assign node45412 = (inp[9]) ? 4'b1100 : 4'b1000;
															assign node45415 = (inp[9]) ? 4'b1000 : 4'b1100;
													assign node45418 = (inp[12]) ? node45428 : node45419;
														assign node45419 = (inp[10]) ? node45425 : node45420;
															assign node45420 = (inp[4]) ? 4'b1000 : node45421;
																assign node45421 = (inp[9]) ? 4'b1000 : 4'b1100;
															assign node45425 = (inp[4]) ? 4'b1110 : 4'b1000;
														assign node45428 = (inp[9]) ? node45430 : 4'b1110;
															assign node45430 = (inp[4]) ? 4'b1010 : 4'b1110;
												assign node45433 = (inp[5]) ? node45453 : node45434;
													assign node45434 = (inp[9]) ? node45442 : node45435;
														assign node45435 = (inp[4]) ? node45437 : 4'b1010;
															assign node45437 = (inp[12]) ? 4'b1110 : node45438;
																assign node45438 = (inp[10]) ? 4'b1110 : 4'b1010;
														assign node45442 = (inp[4]) ? node45448 : node45443;
															assign node45443 = (inp[12]) ? 4'b1110 : node45444;
																assign node45444 = (inp[10]) ? 4'b1110 : 4'b1010;
															assign node45448 = (inp[10]) ? 4'b1010 : node45449;
																assign node45449 = (inp[12]) ? 4'b1010 : 4'b1110;
													assign node45453 = (inp[12]) ? node45461 : node45454;
														assign node45454 = (inp[10]) ? node45456 : 4'b1010;
															assign node45456 = (inp[9]) ? 4'b1100 : node45457;
																assign node45457 = (inp[4]) ? 4'b1100 : 4'b1010;
														assign node45461 = (inp[9]) ? node45463 : 4'b1100;
															assign node45463 = (inp[4]) ? 4'b1000 : 4'b1100;
											assign node45466 = (inp[0]) ? node45500 : node45467;
												assign node45467 = (inp[5]) ? node45487 : node45468;
													assign node45468 = (inp[4]) ? node45478 : node45469;
														assign node45469 = (inp[9]) ? node45475 : node45470;
															assign node45470 = (inp[10]) ? 4'b1000 : node45471;
																assign node45471 = (inp[12]) ? 4'b1000 : 4'b1100;
															assign node45475 = (inp[12]) ? 4'b1110 : 4'b1000;
														assign node45478 = (inp[9]) ? node45482 : node45479;
															assign node45479 = (inp[10]) ? 4'b1110 : 4'b1000;
															assign node45482 = (inp[12]) ? 4'b1010 : node45483;
																assign node45483 = (inp[10]) ? 4'b1010 : 4'b1110;
													assign node45487 = (inp[12]) ? node45493 : node45488;
														assign node45488 = (inp[10]) ? node45490 : 4'b1110;
															assign node45490 = (inp[4]) ? 4'b1110 : 4'b1010;
														assign node45493 = (inp[10]) ? node45495 : 4'b1010;
															assign node45495 = (inp[9]) ? 4'b1010 : node45496;
																assign node45496 = (inp[4]) ? 4'b1110 : 4'b1010;
												assign node45500 = (inp[5]) ? node45514 : node45501;
													assign node45501 = (inp[9]) ? node45507 : node45502;
														assign node45502 = (inp[4]) ? node45504 : 4'b1010;
															assign node45504 = (inp[10]) ? 4'b1100 : 4'b1010;
														assign node45507 = (inp[12]) ? 4'b1000 : node45508;
															assign node45508 = (inp[4]) ? 4'b1100 : node45509;
																assign node45509 = (inp[10]) ? 4'b1100 : 4'b1010;
													assign node45514 = (inp[10]) ? node45530 : node45515;
														assign node45515 = (inp[12]) ? node45523 : node45516;
															assign node45516 = (inp[4]) ? node45520 : node45517;
																assign node45517 = (inp[9]) ? 4'b1000 : 4'b1100;
																assign node45520 = (inp[9]) ? 4'b1100 : 4'b1000;
															assign node45523 = (inp[4]) ? node45527 : node45524;
																assign node45524 = (inp[9]) ? 4'b1100 : 4'b1000;
																assign node45527 = (inp[9]) ? 4'b1000 : 4'b1100;
														assign node45530 = (inp[12]) ? node45532 : 4'b1000;
															assign node45532 = (inp[4]) ? node45536 : node45533;
																assign node45533 = (inp[9]) ? 4'b1100 : 4'b1000;
																assign node45536 = (inp[9]) ? 4'b1000 : 4'b1100;
					assign node45539 = (inp[10]) ? node48029 : node45540;
						assign node45540 = (inp[5]) ? node46732 : node45541;
							assign node45541 = (inp[15]) ? node46139 : node45542;
								assign node45542 = (inp[0]) ? node45858 : node45543;
									assign node45543 = (inp[3]) ? node45709 : node45544;
										assign node45544 = (inp[12]) ? node45624 : node45545;
											assign node45545 = (inp[14]) ? node45593 : node45546;
												assign node45546 = (inp[9]) ? node45570 : node45547;
													assign node45547 = (inp[4]) ? node45557 : node45548;
														assign node45548 = (inp[8]) ? node45550 : 4'b1110;
															assign node45550 = (inp[7]) ? node45554 : node45551;
																assign node45551 = (inp[2]) ? 4'b1111 : 4'b1110;
																assign node45554 = (inp[2]) ? 4'b1110 : 4'b1111;
														assign node45557 = (inp[8]) ? node45563 : node45558;
															assign node45558 = (inp[2]) ? 4'b1010 : node45559;
																assign node45559 = (inp[7]) ? 4'b1010 : 4'b1011;
															assign node45563 = (inp[7]) ? node45567 : node45564;
																assign node45564 = (inp[2]) ? 4'b1011 : 4'b1010;
																assign node45567 = (inp[2]) ? 4'b1010 : 4'b1011;
													assign node45570 = (inp[4]) ? node45582 : node45571;
														assign node45571 = (inp[7]) ? node45577 : node45572;
															assign node45572 = (inp[8]) ? 4'b1010 : node45573;
																assign node45573 = (inp[2]) ? 4'b1010 : 4'b1011;
															assign node45577 = (inp[2]) ? node45579 : 4'b1011;
																assign node45579 = (inp[8]) ? 4'b1010 : 4'b1011;
														assign node45582 = (inp[2]) ? node45588 : node45583;
															assign node45583 = (inp[8]) ? 4'b1110 : node45584;
																assign node45584 = (inp[7]) ? 4'b1110 : 4'b1111;
															assign node45588 = (inp[8]) ? 4'b1111 : node45589;
																assign node45589 = (inp[7]) ? 4'b1111 : 4'b1110;
												assign node45593 = (inp[7]) ? node45609 : node45594;
													assign node45594 = (inp[8]) ? node45602 : node45595;
														assign node45595 = (inp[9]) ? node45599 : node45596;
															assign node45596 = (inp[4]) ? 4'b1010 : 4'b1110;
															assign node45599 = (inp[4]) ? 4'b1110 : 4'b1010;
														assign node45602 = (inp[4]) ? node45606 : node45603;
															assign node45603 = (inp[9]) ? 4'b1011 : 4'b1111;
															assign node45606 = (inp[9]) ? 4'b1111 : 4'b1011;
													assign node45609 = (inp[8]) ? node45617 : node45610;
														assign node45610 = (inp[4]) ? node45614 : node45611;
															assign node45611 = (inp[9]) ? 4'b1011 : 4'b1111;
															assign node45614 = (inp[9]) ? 4'b1111 : 4'b1011;
														assign node45617 = (inp[9]) ? node45621 : node45618;
															assign node45618 = (inp[4]) ? 4'b1010 : 4'b1110;
															assign node45621 = (inp[4]) ? 4'b1110 : 4'b1010;
											assign node45624 = (inp[2]) ? node45676 : node45625;
												assign node45625 = (inp[14]) ? node45649 : node45626;
													assign node45626 = (inp[9]) ? node45638 : node45627;
														assign node45627 = (inp[4]) ? node45633 : node45628;
															assign node45628 = (inp[7]) ? 4'b1011 : node45629;
																assign node45629 = (inp[8]) ? 4'b1010 : 4'b1011;
															assign node45633 = (inp[8]) ? 4'b1111 : node45634;
																assign node45634 = (inp[7]) ? 4'b1110 : 4'b1111;
														assign node45638 = (inp[4]) ? node45646 : node45639;
															assign node45639 = (inp[7]) ? node45643 : node45640;
																assign node45640 = (inp[8]) ? 4'b1110 : 4'b1111;
																assign node45643 = (inp[8]) ? 4'b1111 : 4'b1110;
															assign node45646 = (inp[7]) ? 4'b1010 : 4'b1011;
													assign node45649 = (inp[4]) ? node45663 : node45650;
														assign node45650 = (inp[9]) ? node45656 : node45651;
															assign node45651 = (inp[8]) ? node45653 : 4'b1010;
																assign node45653 = (inp[7]) ? 4'b1010 : 4'b1011;
															assign node45656 = (inp[8]) ? node45660 : node45657;
																assign node45657 = (inp[7]) ? 4'b1111 : 4'b1110;
																assign node45660 = (inp[7]) ? 4'b1110 : 4'b1111;
														assign node45663 = (inp[9]) ? node45671 : node45664;
															assign node45664 = (inp[7]) ? node45668 : node45665;
																assign node45665 = (inp[8]) ? 4'b1111 : 4'b1110;
																assign node45668 = (inp[8]) ? 4'b1110 : 4'b1111;
															assign node45671 = (inp[8]) ? 4'b1010 : node45672;
																assign node45672 = (inp[7]) ? 4'b1011 : 4'b1010;
												assign node45676 = (inp[8]) ? node45692 : node45677;
													assign node45677 = (inp[7]) ? node45685 : node45678;
														assign node45678 = (inp[9]) ? node45682 : node45679;
															assign node45679 = (inp[4]) ? 4'b1110 : 4'b1010;
															assign node45682 = (inp[4]) ? 4'b1010 : 4'b1110;
														assign node45685 = (inp[14]) ? node45687 : 4'b1111;
															assign node45687 = (inp[9]) ? 4'b1111 : node45688;
																assign node45688 = (inp[4]) ? 4'b1111 : 4'b1011;
													assign node45692 = (inp[7]) ? node45702 : node45693;
														assign node45693 = (inp[14]) ? node45697 : node45694;
															assign node45694 = (inp[4]) ? 4'b1011 : 4'b1111;
															assign node45697 = (inp[4]) ? node45699 : 4'b1011;
																assign node45699 = (inp[9]) ? 4'b1011 : 4'b1111;
														assign node45702 = (inp[4]) ? node45706 : node45703;
															assign node45703 = (inp[9]) ? 4'b1110 : 4'b1010;
															assign node45706 = (inp[9]) ? 4'b1010 : 4'b1110;
										assign node45709 = (inp[9]) ? node45791 : node45710;
											assign node45710 = (inp[4]) ? node45748 : node45711;
												assign node45711 = (inp[12]) ? node45727 : node45712;
													assign node45712 = (inp[14]) ? node45720 : node45713;
														assign node45713 = (inp[8]) ? node45715 : 4'b1111;
															assign node45715 = (inp[2]) ? 4'b1111 : node45716;
																assign node45716 = (inp[7]) ? 4'b1111 : 4'b1110;
														assign node45720 = (inp[7]) ? node45724 : node45721;
															assign node45721 = (inp[8]) ? 4'b1111 : 4'b1110;
															assign node45724 = (inp[8]) ? 4'b1110 : 4'b1111;
													assign node45727 = (inp[2]) ? node45741 : node45728;
														assign node45728 = (inp[8]) ? node45734 : node45729;
															assign node45729 = (inp[14]) ? 4'b1011 : node45730;
																assign node45730 = (inp[7]) ? 4'b1010 : 4'b1011;
															assign node45734 = (inp[14]) ? node45738 : node45735;
																assign node45735 = (inp[7]) ? 4'b1011 : 4'b1010;
																assign node45738 = (inp[7]) ? 4'b1010 : 4'b1011;
														assign node45741 = (inp[8]) ? node45745 : node45742;
															assign node45742 = (inp[7]) ? 4'b1011 : 4'b1010;
															assign node45745 = (inp[7]) ? 4'b1010 : 4'b1011;
												assign node45748 = (inp[12]) ? node45772 : node45749;
													assign node45749 = (inp[2]) ? node45765 : node45750;
														assign node45750 = (inp[8]) ? node45758 : node45751;
															assign node45751 = (inp[7]) ? node45755 : node45752;
																assign node45752 = (inp[14]) ? 4'b1010 : 4'b1011;
																assign node45755 = (inp[14]) ? 4'b1011 : 4'b1010;
															assign node45758 = (inp[14]) ? node45762 : node45759;
																assign node45759 = (inp[7]) ? 4'b1011 : 4'b1010;
																assign node45762 = (inp[7]) ? 4'b1010 : 4'b1011;
														assign node45765 = (inp[14]) ? node45769 : node45766;
															assign node45766 = (inp[8]) ? 4'b1010 : 4'b1011;
															assign node45769 = (inp[8]) ? 4'b1011 : 4'b1010;
													assign node45772 = (inp[14]) ? node45786 : node45773;
														assign node45773 = (inp[7]) ? node45781 : node45774;
															assign node45774 = (inp[8]) ? node45778 : node45775;
																assign node45775 = (inp[2]) ? 4'b1100 : 4'b1101;
																assign node45778 = (inp[2]) ? 4'b1101 : 4'b1100;
															assign node45781 = (inp[2]) ? node45783 : 4'b1100;
																assign node45783 = (inp[8]) ? 4'b1100 : 4'b1101;
														assign node45786 = (inp[7]) ? node45788 : 4'b1101;
															assign node45788 = (inp[8]) ? 4'b1100 : 4'b1101;
											assign node45791 = (inp[12]) ? node45825 : node45792;
												assign node45792 = (inp[4]) ? node45806 : node45793;
													assign node45793 = (inp[7]) ? node45801 : node45794;
														assign node45794 = (inp[8]) ? node45798 : node45795;
															assign node45795 = (inp[14]) ? 4'b1010 : 4'b1011;
															assign node45798 = (inp[14]) ? 4'b1011 : 4'b1010;
														assign node45801 = (inp[8]) ? 4'b1010 : node45802;
															assign node45802 = (inp[14]) ? 4'b1011 : 4'b1010;
													assign node45806 = (inp[2]) ? node45820 : node45807;
														assign node45807 = (inp[8]) ? node45813 : node45808;
															assign node45808 = (inp[14]) ? node45810 : 4'b1100;
																assign node45810 = (inp[7]) ? 4'b1101 : 4'b1100;
															assign node45813 = (inp[7]) ? node45817 : node45814;
																assign node45814 = (inp[14]) ? 4'b1101 : 4'b1100;
																assign node45817 = (inp[14]) ? 4'b1100 : 4'b1101;
														assign node45820 = (inp[7]) ? node45822 : 4'b1101;
															assign node45822 = (inp[8]) ? 4'b1100 : 4'b1101;
												assign node45825 = (inp[4]) ? node45847 : node45826;
													assign node45826 = (inp[14]) ? node45840 : node45827;
														assign node45827 = (inp[8]) ? node45835 : node45828;
															assign node45828 = (inp[2]) ? node45832 : node45829;
																assign node45829 = (inp[7]) ? 4'b1100 : 4'b1101;
																assign node45832 = (inp[7]) ? 4'b1101 : 4'b1100;
															assign node45835 = (inp[2]) ? 4'b1100 : node45836;
																assign node45836 = (inp[7]) ? 4'b1101 : 4'b1100;
														assign node45840 = (inp[7]) ? node45844 : node45841;
															assign node45841 = (inp[8]) ? 4'b1101 : 4'b1100;
															assign node45844 = (inp[8]) ? 4'b1100 : 4'b1101;
													assign node45847 = (inp[8]) ? node45855 : node45848;
														assign node45848 = (inp[7]) ? 4'b1001 : node45849;
															assign node45849 = (inp[2]) ? 4'b1000 : node45850;
																assign node45850 = (inp[14]) ? 4'b1000 : 4'b1001;
														assign node45855 = (inp[7]) ? 4'b1000 : 4'b1001;
									assign node45858 = (inp[3]) ? node46006 : node45859;
										assign node45859 = (inp[12]) ? node45931 : node45860;
											assign node45860 = (inp[8]) ? node45898 : node45861;
												assign node45861 = (inp[7]) ? node45883 : node45862;
													assign node45862 = (inp[2]) ? node45876 : node45863;
														assign node45863 = (inp[14]) ? node45869 : node45864;
															assign node45864 = (inp[4]) ? node45866 : 4'b1001;
																assign node45866 = (inp[9]) ? 4'b1101 : 4'b1001;
															assign node45869 = (inp[9]) ? node45873 : node45870;
																assign node45870 = (inp[4]) ? 4'b1000 : 4'b1100;
																assign node45873 = (inp[4]) ? 4'b1100 : 4'b1000;
														assign node45876 = (inp[9]) ? node45880 : node45877;
															assign node45877 = (inp[4]) ? 4'b1000 : 4'b1100;
															assign node45880 = (inp[4]) ? 4'b1100 : 4'b1000;
													assign node45883 = (inp[14]) ? node45889 : node45884;
														assign node45884 = (inp[9]) ? node45886 : 4'b1001;
															assign node45886 = (inp[4]) ? 4'b1100 : 4'b1000;
														assign node45889 = (inp[2]) ? node45895 : node45890;
															assign node45890 = (inp[9]) ? 4'b1001 : node45891;
																assign node45891 = (inp[4]) ? 4'b1001 : 4'b1101;
															assign node45895 = (inp[4]) ? 4'b1101 : 4'b1001;
												assign node45898 = (inp[7]) ? node45914 : node45899;
													assign node45899 = (inp[2]) ? node45907 : node45900;
														assign node45900 = (inp[4]) ? node45904 : node45901;
															assign node45901 = (inp[9]) ? 4'b1000 : 4'b1100;
															assign node45904 = (inp[9]) ? 4'b1100 : 4'b1000;
														assign node45907 = (inp[4]) ? node45911 : node45908;
															assign node45908 = (inp[9]) ? 4'b1001 : 4'b1101;
															assign node45911 = (inp[9]) ? 4'b1101 : 4'b1001;
													assign node45914 = (inp[2]) ? node45924 : node45915;
														assign node45915 = (inp[14]) ? 4'b1100 : node45916;
															assign node45916 = (inp[9]) ? node45920 : node45917;
																assign node45917 = (inp[4]) ? 4'b1001 : 4'b1101;
																assign node45920 = (inp[4]) ? 4'b1101 : 4'b1001;
														assign node45924 = (inp[4]) ? node45928 : node45925;
															assign node45925 = (inp[9]) ? 4'b1000 : 4'b1100;
															assign node45928 = (inp[9]) ? 4'b1100 : 4'b1000;
											assign node45931 = (inp[7]) ? node45963 : node45932;
												assign node45932 = (inp[8]) ? node45944 : node45933;
													assign node45933 = (inp[4]) ? node45941 : node45934;
														assign node45934 = (inp[9]) ? node45936 : 4'b1001;
															assign node45936 = (inp[14]) ? 4'b1100 : node45937;
																assign node45937 = (inp[2]) ? 4'b1100 : 4'b1101;
														assign node45941 = (inp[9]) ? 4'b1000 : 4'b1100;
													assign node45944 = (inp[2]) ? node45956 : node45945;
														assign node45945 = (inp[14]) ? node45951 : node45946;
															assign node45946 = (inp[4]) ? 4'b1100 : node45947;
																assign node45947 = (inp[9]) ? 4'b1100 : 4'b1000;
															assign node45951 = (inp[9]) ? node45953 : 4'b1101;
																assign node45953 = (inp[4]) ? 4'b1001 : 4'b1101;
														assign node45956 = (inp[9]) ? node45960 : node45957;
															assign node45957 = (inp[4]) ? 4'b1101 : 4'b1001;
															assign node45960 = (inp[4]) ? 4'b1001 : 4'b1101;
												assign node45963 = (inp[8]) ? node45977 : node45964;
													assign node45964 = (inp[2]) ? node45970 : node45965;
														assign node45965 = (inp[14]) ? 4'b1001 : node45966;
															assign node45966 = (inp[4]) ? 4'b1100 : 4'b1000;
														assign node45970 = (inp[9]) ? node45974 : node45971;
															assign node45971 = (inp[4]) ? 4'b1101 : 4'b1001;
															assign node45974 = (inp[4]) ? 4'b1001 : 4'b1101;
													assign node45977 = (inp[14]) ? node45991 : node45978;
														assign node45978 = (inp[2]) ? node45986 : node45979;
															assign node45979 = (inp[9]) ? node45983 : node45980;
																assign node45980 = (inp[4]) ? 4'b1101 : 4'b1001;
																assign node45983 = (inp[4]) ? 4'b1001 : 4'b1101;
															assign node45986 = (inp[9]) ? node45988 : 4'b1100;
																assign node45988 = (inp[4]) ? 4'b1000 : 4'b1100;
														assign node45991 = (inp[2]) ? node45999 : node45992;
															assign node45992 = (inp[9]) ? node45996 : node45993;
																assign node45993 = (inp[4]) ? 4'b1100 : 4'b1000;
																assign node45996 = (inp[4]) ? 4'b1000 : 4'b1100;
															assign node45999 = (inp[4]) ? node46003 : node46000;
																assign node46000 = (inp[9]) ? 4'b1100 : 4'b1000;
																assign node46003 = (inp[9]) ? 4'b1000 : 4'b1100;
										assign node46006 = (inp[12]) ? node46068 : node46007;
											assign node46007 = (inp[4]) ? node46041 : node46008;
												assign node46008 = (inp[9]) ? node46018 : node46009;
													assign node46009 = (inp[7]) ? 4'b1101 : node46010;
														assign node46010 = (inp[8]) ? node46012 : 4'b1100;
															assign node46012 = (inp[14]) ? 4'b1101 : node46013;
																assign node46013 = (inp[2]) ? 4'b1101 : 4'b1100;
													assign node46018 = (inp[8]) ? node46030 : node46019;
														assign node46019 = (inp[7]) ? node46025 : node46020;
															assign node46020 = (inp[2]) ? 4'b1000 : node46021;
																assign node46021 = (inp[14]) ? 4'b1000 : 4'b1001;
															assign node46025 = (inp[2]) ? 4'b1001 : node46026;
																assign node46026 = (inp[14]) ? 4'b1001 : 4'b1000;
														assign node46030 = (inp[7]) ? node46036 : node46031;
															assign node46031 = (inp[2]) ? 4'b1001 : node46032;
																assign node46032 = (inp[14]) ? 4'b1001 : 4'b1000;
															assign node46036 = (inp[14]) ? 4'b1000 : node46037;
																assign node46037 = (inp[2]) ? 4'b1000 : 4'b1001;
												assign node46041 = (inp[9]) ? node46053 : node46042;
													assign node46042 = (inp[8]) ? node46044 : 4'b1001;
														assign node46044 = (inp[7]) ? node46050 : node46045;
															assign node46045 = (inp[2]) ? 4'b1001 : node46046;
																assign node46046 = (inp[14]) ? 4'b1001 : 4'b1000;
															assign node46050 = (inp[2]) ? 4'b1000 : 4'b1001;
													assign node46053 = (inp[8]) ? node46061 : node46054;
														assign node46054 = (inp[7]) ? 4'b1111 : node46055;
															assign node46055 = (inp[14]) ? 4'b1110 : node46056;
																assign node46056 = (inp[2]) ? 4'b1110 : 4'b1111;
														assign node46061 = (inp[7]) ? 4'b1110 : node46062;
															assign node46062 = (inp[2]) ? 4'b1111 : node46063;
																assign node46063 = (inp[14]) ? 4'b1111 : 4'b1110;
											assign node46068 = (inp[9]) ? node46100 : node46069;
												assign node46069 = (inp[4]) ? node46083 : node46070;
													assign node46070 = (inp[7]) ? node46078 : node46071;
														assign node46071 = (inp[8]) ? 4'b1001 : node46072;
															assign node46072 = (inp[14]) ? 4'b1000 : node46073;
																assign node46073 = (inp[2]) ? 4'b1000 : 4'b1001;
														assign node46078 = (inp[8]) ? 4'b1000 : node46079;
															assign node46079 = (inp[14]) ? 4'b1001 : 4'b1000;
													assign node46083 = (inp[8]) ? node46091 : node46084;
														assign node46084 = (inp[7]) ? 4'b1111 : node46085;
															assign node46085 = (inp[2]) ? 4'b1110 : node46086;
																assign node46086 = (inp[14]) ? 4'b1110 : 4'b1111;
														assign node46091 = (inp[7]) ? node46095 : node46092;
															assign node46092 = (inp[14]) ? 4'b1111 : 4'b1110;
															assign node46095 = (inp[2]) ? 4'b1110 : node46096;
																assign node46096 = (inp[14]) ? 4'b1110 : 4'b1111;
												assign node46100 = (inp[4]) ? node46122 : node46101;
													assign node46101 = (inp[8]) ? node46111 : node46102;
														assign node46102 = (inp[7]) ? node46108 : node46103;
															assign node46103 = (inp[2]) ? 4'b1110 : node46104;
																assign node46104 = (inp[14]) ? 4'b1110 : 4'b1111;
															assign node46108 = (inp[2]) ? 4'b1111 : 4'b1110;
														assign node46111 = (inp[7]) ? node46117 : node46112;
															assign node46112 = (inp[2]) ? 4'b1111 : node46113;
																assign node46113 = (inp[14]) ? 4'b1111 : 4'b1110;
															assign node46117 = (inp[14]) ? 4'b1110 : node46118;
																assign node46118 = (inp[2]) ? 4'b1110 : 4'b1111;
													assign node46122 = (inp[8]) ? node46132 : node46123;
														assign node46123 = (inp[7]) ? node46129 : node46124;
															assign node46124 = (inp[2]) ? 4'b1010 : node46125;
																assign node46125 = (inp[14]) ? 4'b1010 : 4'b1011;
															assign node46129 = (inp[2]) ? 4'b1011 : 4'b1010;
														assign node46132 = (inp[7]) ? node46134 : 4'b1011;
															assign node46134 = (inp[14]) ? 4'b1010 : node46135;
																assign node46135 = (inp[2]) ? 4'b1010 : 4'b1011;
								assign node46139 = (inp[0]) ? node46431 : node46140;
									assign node46140 = (inp[3]) ? node46276 : node46141;
										assign node46141 = (inp[7]) ? node46203 : node46142;
											assign node46142 = (inp[8]) ? node46168 : node46143;
												assign node46143 = (inp[14]) ? node46151 : node46144;
													assign node46144 = (inp[2]) ? node46146 : 4'b1001;
														assign node46146 = (inp[4]) ? 4'b1000 : node46147;
															assign node46147 = (inp[12]) ? 4'b1000 : 4'b1100;
													assign node46151 = (inp[12]) ? node46159 : node46152;
														assign node46152 = (inp[2]) ? node46154 : 4'b1000;
															assign node46154 = (inp[4]) ? node46156 : 4'b1100;
																assign node46156 = (inp[9]) ? 4'b1100 : 4'b1000;
														assign node46159 = (inp[2]) ? node46161 : 4'b1100;
															assign node46161 = (inp[4]) ? node46165 : node46162;
																assign node46162 = (inp[9]) ? 4'b1100 : 4'b1000;
																assign node46165 = (inp[9]) ? 4'b1000 : 4'b1100;
												assign node46168 = (inp[14]) ? node46188 : node46169;
													assign node46169 = (inp[2]) ? node46183 : node46170;
														assign node46170 = (inp[12]) ? node46176 : node46171;
															assign node46171 = (inp[9]) ? node46173 : 4'b1100;
																assign node46173 = (inp[4]) ? 4'b1100 : 4'b1000;
															assign node46176 = (inp[9]) ? node46180 : node46177;
																assign node46177 = (inp[4]) ? 4'b1100 : 4'b1000;
																assign node46180 = (inp[4]) ? 4'b1000 : 4'b1100;
														assign node46183 = (inp[12]) ? 4'b1001 : node46184;
															assign node46184 = (inp[9]) ? 4'b1101 : 4'b1001;
													assign node46188 = (inp[9]) ? node46196 : node46189;
														assign node46189 = (inp[12]) ? node46193 : node46190;
															assign node46190 = (inp[4]) ? 4'b1001 : 4'b1101;
															assign node46193 = (inp[4]) ? 4'b1101 : 4'b1001;
														assign node46196 = (inp[2]) ? node46198 : 4'b1001;
															assign node46198 = (inp[4]) ? node46200 : 4'b1001;
																assign node46200 = (inp[12]) ? 4'b1001 : 4'b1101;
											assign node46203 = (inp[8]) ? node46239 : node46204;
												assign node46204 = (inp[2]) ? node46226 : node46205;
													assign node46205 = (inp[14]) ? node46215 : node46206;
														assign node46206 = (inp[12]) ? 4'b1100 : node46207;
															assign node46207 = (inp[4]) ? node46211 : node46208;
																assign node46208 = (inp[9]) ? 4'b1000 : 4'b1100;
																assign node46211 = (inp[9]) ? 4'b1100 : 4'b1000;
														assign node46215 = (inp[4]) ? node46221 : node46216;
															assign node46216 = (inp[9]) ? node46218 : 4'b1101;
																assign node46218 = (inp[12]) ? 4'b1101 : 4'b1001;
															assign node46221 = (inp[12]) ? node46223 : 4'b1001;
																assign node46223 = (inp[9]) ? 4'b1001 : 4'b1101;
													assign node46226 = (inp[12]) ? node46232 : node46227;
														assign node46227 = (inp[4]) ? 4'b1001 : node46228;
															assign node46228 = (inp[9]) ? 4'b1001 : 4'b1101;
														assign node46232 = (inp[9]) ? node46236 : node46233;
															assign node46233 = (inp[4]) ? 4'b1101 : 4'b1001;
															assign node46236 = (inp[4]) ? 4'b1001 : 4'b1101;
												assign node46239 = (inp[14]) ? node46261 : node46240;
													assign node46240 = (inp[2]) ? node46252 : node46241;
														assign node46241 = (inp[12]) ? node46247 : node46242;
															assign node46242 = (inp[9]) ? 4'b1001 : node46243;
																assign node46243 = (inp[4]) ? 4'b1001 : 4'b1101;
															assign node46247 = (inp[4]) ? 4'b1101 : node46248;
																assign node46248 = (inp[9]) ? 4'b1101 : 4'b1001;
														assign node46252 = (inp[12]) ? node46254 : 4'b1000;
															assign node46254 = (inp[9]) ? node46258 : node46255;
																assign node46255 = (inp[4]) ? 4'b1100 : 4'b1000;
																assign node46258 = (inp[4]) ? 4'b1000 : 4'b1100;
													assign node46261 = (inp[4]) ? node46269 : node46262;
														assign node46262 = (inp[9]) ? node46266 : node46263;
															assign node46263 = (inp[12]) ? 4'b1000 : 4'b1100;
															assign node46266 = (inp[12]) ? 4'b1100 : 4'b1000;
														assign node46269 = (inp[12]) ? node46273 : node46270;
															assign node46270 = (inp[9]) ? 4'b1100 : 4'b1000;
															assign node46273 = (inp[9]) ? 4'b1000 : 4'b1100;
										assign node46276 = (inp[9]) ? node46350 : node46277;
											assign node46277 = (inp[4]) ? node46325 : node46278;
												assign node46278 = (inp[12]) ? node46298 : node46279;
													assign node46279 = (inp[8]) ? node46289 : node46280;
														assign node46280 = (inp[14]) ? 4'b1100 : node46281;
															assign node46281 = (inp[7]) ? node46285 : node46282;
																assign node46282 = (inp[2]) ? 4'b1100 : 4'b1101;
																assign node46285 = (inp[2]) ? 4'b1101 : 4'b1100;
														assign node46289 = (inp[14]) ? 4'b1101 : node46290;
															assign node46290 = (inp[7]) ? node46294 : node46291;
																assign node46291 = (inp[2]) ? 4'b1101 : 4'b1100;
																assign node46294 = (inp[2]) ? 4'b1100 : 4'b1101;
													assign node46298 = (inp[14]) ? node46312 : node46299;
														assign node46299 = (inp[7]) ? node46305 : node46300;
															assign node46300 = (inp[2]) ? 4'b1000 : node46301;
																assign node46301 = (inp[8]) ? 4'b1000 : 4'b1001;
															assign node46305 = (inp[8]) ? node46309 : node46306;
																assign node46306 = (inp[2]) ? 4'b1001 : 4'b1000;
																assign node46309 = (inp[2]) ? 4'b1000 : 4'b1001;
														assign node46312 = (inp[2]) ? node46320 : node46313;
															assign node46313 = (inp[8]) ? node46317 : node46314;
																assign node46314 = (inp[7]) ? 4'b1001 : 4'b1000;
																assign node46317 = (inp[7]) ? 4'b1000 : 4'b1001;
															assign node46320 = (inp[7]) ? 4'b1001 : node46321;
																assign node46321 = (inp[8]) ? 4'b1001 : 4'b1000;
												assign node46325 = (inp[12]) ? node46341 : node46326;
													assign node46326 = (inp[2]) ? node46334 : node46327;
														assign node46327 = (inp[14]) ? node46329 : 4'b1001;
															assign node46329 = (inp[8]) ? 4'b1000 : node46330;
																assign node46330 = (inp[7]) ? 4'b1001 : 4'b1000;
														assign node46334 = (inp[7]) ? node46338 : node46335;
															assign node46335 = (inp[8]) ? 4'b1001 : 4'b1000;
															assign node46338 = (inp[8]) ? 4'b1000 : 4'b1001;
													assign node46341 = (inp[8]) ? node46343 : 4'b1110;
														assign node46343 = (inp[14]) ? 4'b1111 : node46344;
															assign node46344 = (inp[2]) ? 4'b1110 : node46345;
																assign node46345 = (inp[7]) ? 4'b1111 : 4'b1110;
											assign node46350 = (inp[12]) ? node46388 : node46351;
												assign node46351 = (inp[4]) ? node46375 : node46352;
													assign node46352 = (inp[14]) ? node46362 : node46353;
														assign node46353 = (inp[8]) ? node46355 : 4'b1001;
															assign node46355 = (inp[2]) ? node46359 : node46356;
																assign node46356 = (inp[7]) ? 4'b1001 : 4'b1000;
																assign node46359 = (inp[7]) ? 4'b1000 : 4'b1001;
														assign node46362 = (inp[2]) ? node46370 : node46363;
															assign node46363 = (inp[7]) ? node46367 : node46364;
																assign node46364 = (inp[8]) ? 4'b1001 : 4'b1000;
																assign node46367 = (inp[8]) ? 4'b1000 : 4'b1001;
															assign node46370 = (inp[7]) ? node46372 : 4'b1000;
																assign node46372 = (inp[8]) ? 4'b1000 : 4'b1001;
													assign node46375 = (inp[8]) ? node46379 : node46376;
														assign node46376 = (inp[14]) ? 4'b1111 : 4'b1110;
														assign node46379 = (inp[7]) ? node46385 : node46380;
															assign node46380 = (inp[2]) ? 4'b1111 : node46381;
																assign node46381 = (inp[14]) ? 4'b1111 : 4'b1110;
															assign node46385 = (inp[14]) ? 4'b1110 : 4'b1111;
												assign node46388 = (inp[4]) ? node46414 : node46389;
													assign node46389 = (inp[2]) ? node46401 : node46390;
														assign node46390 = (inp[14]) ? node46396 : node46391;
															assign node46391 = (inp[8]) ? 4'b1110 : node46392;
																assign node46392 = (inp[7]) ? 4'b1110 : 4'b1111;
															assign node46396 = (inp[7]) ? 4'b1111 : node46397;
																assign node46397 = (inp[8]) ? 4'b1111 : 4'b1110;
														assign node46401 = (inp[14]) ? node46407 : node46402;
															assign node46402 = (inp[8]) ? node46404 : 4'b1111;
																assign node46404 = (inp[7]) ? 4'b1110 : 4'b1111;
															assign node46407 = (inp[8]) ? node46411 : node46408;
																assign node46408 = (inp[7]) ? 4'b1111 : 4'b1110;
																assign node46411 = (inp[7]) ? 4'b1110 : 4'b1111;
													assign node46414 = (inp[8]) ? node46424 : node46415;
														assign node46415 = (inp[2]) ? 4'b1011 : node46416;
															assign node46416 = (inp[14]) ? node46420 : node46417;
																assign node46417 = (inp[7]) ? 4'b1010 : 4'b1011;
																assign node46420 = (inp[7]) ? 4'b1011 : 4'b1010;
														assign node46424 = (inp[7]) ? 4'b1010 : node46425;
															assign node46425 = (inp[2]) ? 4'b1011 : node46426;
																assign node46426 = (inp[14]) ? 4'b1011 : 4'b1010;
									assign node46431 = (inp[3]) ? node46601 : node46432;
										assign node46432 = (inp[9]) ? node46536 : node46433;
											assign node46433 = (inp[14]) ? node46485 : node46434;
												assign node46434 = (inp[7]) ? node46456 : node46435;
													assign node46435 = (inp[12]) ? node46445 : node46436;
														assign node46436 = (inp[4]) ? 4'b1011 : node46437;
															assign node46437 = (inp[8]) ? node46441 : node46438;
																assign node46438 = (inp[2]) ? 4'b1110 : 4'b1111;
																assign node46441 = (inp[2]) ? 4'b1111 : 4'b1110;
														assign node46445 = (inp[4]) ? node46451 : node46446;
															assign node46446 = (inp[2]) ? node46448 : 4'b1010;
																assign node46448 = (inp[8]) ? 4'b1011 : 4'b1010;
															assign node46451 = (inp[8]) ? 4'b1110 : node46452;
																assign node46452 = (inp[2]) ? 4'b1110 : 4'b1111;
													assign node46456 = (inp[2]) ? node46472 : node46457;
														assign node46457 = (inp[8]) ? node46465 : node46458;
															assign node46458 = (inp[12]) ? node46462 : node46459;
																assign node46459 = (inp[4]) ? 4'b1010 : 4'b1110;
																assign node46462 = (inp[4]) ? 4'b1110 : 4'b1010;
															assign node46465 = (inp[12]) ? node46469 : node46466;
																assign node46466 = (inp[4]) ? 4'b1011 : 4'b1111;
																assign node46469 = (inp[4]) ? 4'b1111 : 4'b1011;
														assign node46472 = (inp[8]) ? node46478 : node46473;
															assign node46473 = (inp[4]) ? node46475 : 4'b1011;
																assign node46475 = (inp[12]) ? 4'b1111 : 4'b1011;
															assign node46478 = (inp[12]) ? node46482 : node46479;
																assign node46479 = (inp[4]) ? 4'b1010 : 4'b1110;
																assign node46482 = (inp[4]) ? 4'b1110 : 4'b1010;
												assign node46485 = (inp[2]) ? node46509 : node46486;
													assign node46486 = (inp[4]) ? node46498 : node46487;
														assign node46487 = (inp[12]) ? node46493 : node46488;
															assign node46488 = (inp[8]) ? node46490 : 4'b1111;
																assign node46490 = (inp[7]) ? 4'b1110 : 4'b1111;
															assign node46493 = (inp[8]) ? 4'b1011 : node46494;
																assign node46494 = (inp[7]) ? 4'b1011 : 4'b1010;
														assign node46498 = (inp[12]) ? node46506 : node46499;
															assign node46499 = (inp[8]) ? node46503 : node46500;
																assign node46500 = (inp[7]) ? 4'b1011 : 4'b1010;
																assign node46503 = (inp[7]) ? 4'b1010 : 4'b1011;
															assign node46506 = (inp[7]) ? 4'b1111 : 4'b1110;
													assign node46509 = (inp[8]) ? node46521 : node46510;
														assign node46510 = (inp[7]) ? node46516 : node46511;
															assign node46511 = (inp[12]) ? 4'b1110 : node46512;
																assign node46512 = (inp[4]) ? 4'b1010 : 4'b1110;
															assign node46516 = (inp[4]) ? 4'b1111 : node46517;
																assign node46517 = (inp[12]) ? 4'b1011 : 4'b1111;
														assign node46521 = (inp[7]) ? node46529 : node46522;
															assign node46522 = (inp[4]) ? node46526 : node46523;
																assign node46523 = (inp[12]) ? 4'b1011 : 4'b1111;
																assign node46526 = (inp[12]) ? 4'b1111 : 4'b1011;
															assign node46529 = (inp[4]) ? node46533 : node46530;
																assign node46530 = (inp[12]) ? 4'b1010 : 4'b1110;
																assign node46533 = (inp[12]) ? 4'b1110 : 4'b1010;
											assign node46536 = (inp[12]) ? node46564 : node46537;
												assign node46537 = (inp[4]) ? node46549 : node46538;
													assign node46538 = (inp[8]) ? node46540 : 4'b1010;
														assign node46540 = (inp[14]) ? node46546 : node46541;
															assign node46541 = (inp[2]) ? 4'b1011 : node46542;
																assign node46542 = (inp[7]) ? 4'b1011 : 4'b1010;
															assign node46546 = (inp[7]) ? 4'b1010 : 4'b1011;
													assign node46549 = (inp[8]) ? node46555 : node46550;
														assign node46550 = (inp[7]) ? 4'b1111 : node46551;
															assign node46551 = (inp[14]) ? 4'b1110 : 4'b1111;
														assign node46555 = (inp[2]) ? 4'b1110 : node46556;
															assign node46556 = (inp[14]) ? node46560 : node46557;
																assign node46557 = (inp[7]) ? 4'b1111 : 4'b1110;
																assign node46560 = (inp[7]) ? 4'b1110 : 4'b1111;
												assign node46564 = (inp[4]) ? node46578 : node46565;
													assign node46565 = (inp[8]) ? node46571 : node46566;
														assign node46566 = (inp[14]) ? node46568 : 4'b1110;
															assign node46568 = (inp[7]) ? 4'b1111 : 4'b1110;
														assign node46571 = (inp[7]) ? node46575 : node46572;
															assign node46572 = (inp[2]) ? 4'b1111 : 4'b1110;
															assign node46575 = (inp[2]) ? 4'b1110 : 4'b1111;
													assign node46578 = (inp[14]) ? node46594 : node46579;
														assign node46579 = (inp[7]) ? node46587 : node46580;
															assign node46580 = (inp[2]) ? node46584 : node46581;
																assign node46581 = (inp[8]) ? 4'b1010 : 4'b1011;
																assign node46584 = (inp[8]) ? 4'b1011 : 4'b1010;
															assign node46587 = (inp[8]) ? node46591 : node46588;
																assign node46588 = (inp[2]) ? 4'b1011 : 4'b1010;
																assign node46591 = (inp[2]) ? 4'b1010 : 4'b1011;
														assign node46594 = (inp[8]) ? node46598 : node46595;
															assign node46595 = (inp[7]) ? 4'b1011 : 4'b1010;
															assign node46598 = (inp[7]) ? 4'b1010 : 4'b1011;
										assign node46601 = (inp[4]) ? node46685 : node46602;
											assign node46602 = (inp[9]) ? node46648 : node46603;
												assign node46603 = (inp[12]) ? node46625 : node46604;
													assign node46604 = (inp[14]) ? node46618 : node46605;
														assign node46605 = (inp[7]) ? node46613 : node46606;
															assign node46606 = (inp[8]) ? node46610 : node46607;
																assign node46607 = (inp[2]) ? 4'b1110 : 4'b1111;
																assign node46610 = (inp[2]) ? 4'b1111 : 4'b1110;
															assign node46613 = (inp[8]) ? node46615 : 4'b1110;
																assign node46615 = (inp[2]) ? 4'b1110 : 4'b1111;
														assign node46618 = (inp[8]) ? node46622 : node46619;
															assign node46619 = (inp[7]) ? 4'b1111 : 4'b1110;
															assign node46622 = (inp[7]) ? 4'b1110 : 4'b1111;
													assign node46625 = (inp[8]) ? node46637 : node46626;
														assign node46626 = (inp[7]) ? node46632 : node46627;
															assign node46627 = (inp[14]) ? 4'b1010 : node46628;
																assign node46628 = (inp[2]) ? 4'b1010 : 4'b1011;
															assign node46632 = (inp[14]) ? 4'b1011 : node46633;
																assign node46633 = (inp[2]) ? 4'b1011 : 4'b1010;
														assign node46637 = (inp[7]) ? node46643 : node46638;
															assign node46638 = (inp[2]) ? 4'b1011 : node46639;
																assign node46639 = (inp[14]) ? 4'b1011 : 4'b1010;
															assign node46643 = (inp[2]) ? 4'b1010 : node46644;
																assign node46644 = (inp[14]) ? 4'b1010 : 4'b1011;
												assign node46648 = (inp[12]) ? node46670 : node46649;
													assign node46649 = (inp[2]) ? node46663 : node46650;
														assign node46650 = (inp[14]) ? node46658 : node46651;
															assign node46651 = (inp[8]) ? node46655 : node46652;
																assign node46652 = (inp[7]) ? 4'b1010 : 4'b1011;
																assign node46655 = (inp[7]) ? 4'b1011 : 4'b1010;
															assign node46658 = (inp[7]) ? 4'b1010 : node46659;
																assign node46659 = (inp[8]) ? 4'b1011 : 4'b1010;
														assign node46663 = (inp[8]) ? node46667 : node46664;
															assign node46664 = (inp[7]) ? 4'b1011 : 4'b1010;
															assign node46667 = (inp[7]) ? 4'b1010 : 4'b1011;
													assign node46670 = (inp[14]) ? node46678 : node46671;
														assign node46671 = (inp[2]) ? node46673 : 4'b1100;
															assign node46673 = (inp[7]) ? 4'b1100 : node46674;
																assign node46674 = (inp[8]) ? 4'b1101 : 4'b1100;
														assign node46678 = (inp[8]) ? node46682 : node46679;
															assign node46679 = (inp[7]) ? 4'b1101 : 4'b1100;
															assign node46682 = (inp[7]) ? 4'b1100 : 4'b1101;
											assign node46685 = (inp[9]) ? node46701 : node46686;
												assign node46686 = (inp[12]) ? node46688 : 4'b1010;
													assign node46688 = (inp[14]) ? node46694 : node46689;
														assign node46689 = (inp[7]) ? node46691 : 4'b1100;
															assign node46691 = (inp[2]) ? 4'b1100 : 4'b1101;
														assign node46694 = (inp[7]) ? node46698 : node46695;
															assign node46695 = (inp[8]) ? 4'b1101 : 4'b1100;
															assign node46698 = (inp[8]) ? 4'b1100 : 4'b1101;
												assign node46701 = (inp[12]) ? node46717 : node46702;
													assign node46702 = (inp[7]) ? node46712 : node46703;
														assign node46703 = (inp[14]) ? 4'b1101 : node46704;
															assign node46704 = (inp[2]) ? node46708 : node46705;
																assign node46705 = (inp[8]) ? 4'b1100 : 4'b1101;
																assign node46708 = (inp[8]) ? 4'b1101 : 4'b1100;
														assign node46712 = (inp[8]) ? 4'b1100 : node46713;
															assign node46713 = (inp[2]) ? 4'b1101 : 4'b1100;
													assign node46717 = (inp[7]) ? node46723 : node46718;
														assign node46718 = (inp[2]) ? node46720 : 4'b1000;
															assign node46720 = (inp[8]) ? 4'b1001 : 4'b1000;
														assign node46723 = (inp[8]) ? node46729 : node46724;
															assign node46724 = (inp[14]) ? 4'b1001 : node46725;
																assign node46725 = (inp[2]) ? 4'b1001 : 4'b1000;
															assign node46729 = (inp[2]) ? 4'b1000 : 4'b1001;
							assign node46732 = (inp[7]) ? node47404 : node46733;
								assign node46733 = (inp[8]) ? node47071 : node46734;
									assign node46734 = (inp[14]) ? node46900 : node46735;
										assign node46735 = (inp[2]) ? node46837 : node46736;
											assign node46736 = (inp[3]) ? node46784 : node46737;
												assign node46737 = (inp[12]) ? node46757 : node46738;
													assign node46738 = (inp[4]) ? node46750 : node46739;
														assign node46739 = (inp[9]) ? node46743 : node46740;
															assign node46740 = (inp[15]) ? 4'b1101 : 4'b1111;
															assign node46743 = (inp[0]) ? node46747 : node46744;
																assign node46744 = (inp[15]) ? 4'b1001 : 4'b1011;
																assign node46747 = (inp[15]) ? 4'b1011 : 4'b1001;
														assign node46750 = (inp[9]) ? 4'b1111 : node46751;
															assign node46751 = (inp[0]) ? 4'b1011 : node46752;
																assign node46752 = (inp[15]) ? 4'b1001 : 4'b1011;
													assign node46757 = (inp[4]) ? node46771 : node46758;
														assign node46758 = (inp[9]) ? node46766 : node46759;
															assign node46759 = (inp[15]) ? node46763 : node46760;
																assign node46760 = (inp[0]) ? 4'b1001 : 4'b1011;
																assign node46763 = (inp[0]) ? 4'b1011 : 4'b1001;
															assign node46766 = (inp[0]) ? 4'b1101 : node46767;
																assign node46767 = (inp[15]) ? 4'b1111 : 4'b1101;
														assign node46771 = (inp[9]) ? node46777 : node46772;
															assign node46772 = (inp[0]) ? node46774 : 4'b1101;
																assign node46774 = (inp[15]) ? 4'b1101 : 4'b1111;
															assign node46777 = (inp[15]) ? node46781 : node46778;
																assign node46778 = (inp[0]) ? 4'b1011 : 4'b1001;
																assign node46781 = (inp[0]) ? 4'b1001 : 4'b1011;
												assign node46784 = (inp[12]) ? node46810 : node46785;
													assign node46785 = (inp[9]) ? node46795 : node46786;
														assign node46786 = (inp[4]) ? node46788 : 4'b1101;
															assign node46788 = (inp[15]) ? node46792 : node46789;
																assign node46789 = (inp[0]) ? 4'b1011 : 4'b1001;
																assign node46792 = (inp[0]) ? 4'b1001 : 4'b1011;
														assign node46795 = (inp[4]) ? node46803 : node46796;
															assign node46796 = (inp[15]) ? node46800 : node46797;
																assign node46797 = (inp[0]) ? 4'b1011 : 4'b1001;
																assign node46800 = (inp[0]) ? 4'b1001 : 4'b1011;
															assign node46803 = (inp[0]) ? node46807 : node46804;
																assign node46804 = (inp[15]) ? 4'b1111 : 4'b1101;
																assign node46807 = (inp[15]) ? 4'b1101 : 4'b1111;
													assign node46810 = (inp[15]) ? node46824 : node46811;
														assign node46811 = (inp[0]) ? node46819 : node46812;
															assign node46812 = (inp[4]) ? node46816 : node46813;
																assign node46813 = (inp[9]) ? 4'b1101 : 4'b1001;
																assign node46816 = (inp[9]) ? 4'b1001 : 4'b1101;
															assign node46819 = (inp[4]) ? node46821 : 4'b1111;
																assign node46821 = (inp[9]) ? 4'b1011 : 4'b1111;
														assign node46824 = (inp[0]) ? node46830 : node46825;
															assign node46825 = (inp[4]) ? 4'b1111 : node46826;
																assign node46826 = (inp[9]) ? 4'b1111 : 4'b1011;
															assign node46830 = (inp[9]) ? node46834 : node46831;
																assign node46831 = (inp[4]) ? 4'b1101 : 4'b1001;
																assign node46834 = (inp[4]) ? 4'b1001 : 4'b1101;
											assign node46837 = (inp[9]) ? node46873 : node46838;
												assign node46838 = (inp[3]) ? node46860 : node46839;
													assign node46839 = (inp[4]) ? node46851 : node46840;
														assign node46840 = (inp[12]) ? node46848 : node46841;
															assign node46841 = (inp[15]) ? node46845 : node46842;
																assign node46842 = (inp[0]) ? 4'b1100 : 4'b1110;
																assign node46845 = (inp[0]) ? 4'b1110 : 4'b1100;
															assign node46848 = (inp[0]) ? 4'b1000 : 4'b1010;
														assign node46851 = (inp[12]) ? node46857 : node46852;
															assign node46852 = (inp[0]) ? node46854 : 4'b1000;
																assign node46854 = (inp[15]) ? 4'b1010 : 4'b1000;
															assign node46857 = (inp[0]) ? 4'b1110 : 4'b1100;
													assign node46860 = (inp[12]) ? node46864 : node46861;
														assign node46861 = (inp[4]) ? 4'b1010 : 4'b1100;
														assign node46864 = (inp[4]) ? 4'b1100 : node46865;
															assign node46865 = (inp[0]) ? node46869 : node46866;
																assign node46866 = (inp[15]) ? 4'b1010 : 4'b1000;
																assign node46869 = (inp[15]) ? 4'b1000 : 4'b1010;
												assign node46873 = (inp[4]) ? node46885 : node46874;
													assign node46874 = (inp[12]) ? node46878 : node46875;
														assign node46875 = (inp[0]) ? 4'b1000 : 4'b1010;
														assign node46878 = (inp[0]) ? node46882 : node46879;
															assign node46879 = (inp[15]) ? 4'b1110 : 4'b1100;
															assign node46882 = (inp[15]) ? 4'b1100 : 4'b1110;
													assign node46885 = (inp[12]) ? node46893 : node46886;
														assign node46886 = (inp[0]) ? node46890 : node46887;
															assign node46887 = (inp[15]) ? 4'b1110 : 4'b1100;
															assign node46890 = (inp[15]) ? 4'b1100 : 4'b1110;
														assign node46893 = (inp[0]) ? node46897 : node46894;
															assign node46894 = (inp[15]) ? 4'b1010 : 4'b1000;
															assign node46897 = (inp[15]) ? 4'b1000 : 4'b1010;
										assign node46900 = (inp[2]) ? node46988 : node46901;
											assign node46901 = (inp[3]) ? node46943 : node46902;
												assign node46902 = (inp[4]) ? node46926 : node46903;
													assign node46903 = (inp[12]) ? node46913 : node46904;
														assign node46904 = (inp[9]) ? 4'b1000 : node46905;
															assign node46905 = (inp[0]) ? node46909 : node46906;
																assign node46906 = (inp[15]) ? 4'b1100 : 4'b1110;
																assign node46909 = (inp[15]) ? 4'b1110 : 4'b1100;
														assign node46913 = (inp[9]) ? node46919 : node46914;
															assign node46914 = (inp[15]) ? 4'b1000 : node46915;
																assign node46915 = (inp[0]) ? 4'b1000 : 4'b1010;
															assign node46919 = (inp[0]) ? node46923 : node46920;
																assign node46920 = (inp[15]) ? 4'b1110 : 4'b1100;
																assign node46923 = (inp[15]) ? 4'b1100 : 4'b1110;
													assign node46926 = (inp[15]) ? node46930 : node46927;
														assign node46927 = (inp[0]) ? 4'b1110 : 4'b1100;
														assign node46930 = (inp[0]) ? node46938 : node46931;
															assign node46931 = (inp[9]) ? node46935 : node46932;
																assign node46932 = (inp[12]) ? 4'b1110 : 4'b1000;
																assign node46935 = (inp[12]) ? 4'b1010 : 4'b1110;
															assign node46938 = (inp[12]) ? node46940 : 4'b1010;
																assign node46940 = (inp[9]) ? 4'b1000 : 4'b1100;
												assign node46943 = (inp[9]) ? node46965 : node46944;
													assign node46944 = (inp[0]) ? node46956 : node46945;
														assign node46945 = (inp[15]) ? node46953 : node46946;
															assign node46946 = (inp[4]) ? node46950 : node46947;
																assign node46947 = (inp[12]) ? 4'b1000 : 4'b1100;
																assign node46950 = (inp[12]) ? 4'b1100 : 4'b1000;
															assign node46953 = (inp[12]) ? 4'b1110 : 4'b1010;
														assign node46956 = (inp[15]) ? node46960 : node46957;
															assign node46957 = (inp[12]) ? 4'b1010 : 4'b1110;
															assign node46960 = (inp[4]) ? node46962 : 4'b1000;
																assign node46962 = (inp[12]) ? 4'b1100 : 4'b1000;
													assign node46965 = (inp[4]) ? node46979 : node46966;
														assign node46966 = (inp[12]) ? node46974 : node46967;
															assign node46967 = (inp[15]) ? node46971 : node46968;
																assign node46968 = (inp[0]) ? 4'b1010 : 4'b1000;
																assign node46971 = (inp[0]) ? 4'b1000 : 4'b1010;
															assign node46974 = (inp[15]) ? node46976 : 4'b1110;
																assign node46976 = (inp[0]) ? 4'b1100 : 4'b1110;
														assign node46979 = (inp[12]) ? node46983 : node46980;
															assign node46980 = (inp[15]) ? 4'b1110 : 4'b1100;
															assign node46983 = (inp[15]) ? 4'b1000 : node46984;
																assign node46984 = (inp[0]) ? 4'b1010 : 4'b1000;
											assign node46988 = (inp[3]) ? node47030 : node46989;
												assign node46989 = (inp[15]) ? node47009 : node46990;
													assign node46990 = (inp[0]) ? node47002 : node46991;
														assign node46991 = (inp[9]) ? node46997 : node46992;
															assign node46992 = (inp[12]) ? node46994 : 4'b1010;
																assign node46994 = (inp[4]) ? 4'b1100 : 4'b1010;
															assign node46997 = (inp[12]) ? node46999 : 4'b1100;
																assign node46999 = (inp[4]) ? 4'b1000 : 4'b1100;
														assign node47002 = (inp[4]) ? 4'b1010 : node47003;
															assign node47003 = (inp[12]) ? 4'b1000 : node47004;
																assign node47004 = (inp[9]) ? 4'b1000 : 4'b1100;
													assign node47009 = (inp[4]) ? node47021 : node47010;
														assign node47010 = (inp[0]) ? node47014 : node47011;
															assign node47011 = (inp[9]) ? 4'b1110 : 4'b1100;
															assign node47014 = (inp[12]) ? node47018 : node47015;
																assign node47015 = (inp[9]) ? 4'b1010 : 4'b1110;
																assign node47018 = (inp[9]) ? 4'b1100 : 4'b1010;
														assign node47021 = (inp[9]) ? node47027 : node47022;
															assign node47022 = (inp[12]) ? 4'b1110 : node47023;
																assign node47023 = (inp[0]) ? 4'b1010 : 4'b1000;
															assign node47027 = (inp[0]) ? 4'b1000 : 4'b1010;
												assign node47030 = (inp[9]) ? node47050 : node47031;
													assign node47031 = (inp[15]) ? node47041 : node47032;
														assign node47032 = (inp[0]) ? node47034 : 4'b1100;
															assign node47034 = (inp[4]) ? node47038 : node47035;
																assign node47035 = (inp[12]) ? 4'b1010 : 4'b1110;
																assign node47038 = (inp[12]) ? 4'b1110 : 4'b1010;
														assign node47041 = (inp[0]) ? 4'b1100 : node47042;
															assign node47042 = (inp[4]) ? node47046 : node47043;
																assign node47043 = (inp[12]) ? 4'b1010 : 4'b1110;
																assign node47046 = (inp[12]) ? 4'b1110 : 4'b1010;
													assign node47050 = (inp[12]) ? node47058 : node47051;
														assign node47051 = (inp[4]) ? node47053 : 4'b1010;
															assign node47053 = (inp[15]) ? 4'b1110 : node47054;
																assign node47054 = (inp[0]) ? 4'b1110 : 4'b1100;
														assign node47058 = (inp[4]) ? node47064 : node47059;
															assign node47059 = (inp[0]) ? node47061 : 4'b1110;
																assign node47061 = (inp[15]) ? 4'b1100 : 4'b1110;
															assign node47064 = (inp[15]) ? node47068 : node47065;
																assign node47065 = (inp[0]) ? 4'b1010 : 4'b1000;
																assign node47068 = (inp[0]) ? 4'b1000 : 4'b1010;
									assign node47071 = (inp[14]) ? node47233 : node47072;
										assign node47072 = (inp[2]) ? node47162 : node47073;
											assign node47073 = (inp[15]) ? node47121 : node47074;
												assign node47074 = (inp[0]) ? node47100 : node47075;
													assign node47075 = (inp[3]) ? node47085 : node47076;
														assign node47076 = (inp[12]) ? 4'b1000 : node47077;
															assign node47077 = (inp[4]) ? node47081 : node47078;
																assign node47078 = (inp[9]) ? 4'b1010 : 4'b1110;
																assign node47081 = (inp[9]) ? 4'b1100 : 4'b1010;
														assign node47085 = (inp[12]) ? node47093 : node47086;
															assign node47086 = (inp[4]) ? node47090 : node47087;
																assign node47087 = (inp[9]) ? 4'b1000 : 4'b1100;
																assign node47090 = (inp[9]) ? 4'b1100 : 4'b1000;
															assign node47093 = (inp[9]) ? node47097 : node47094;
																assign node47094 = (inp[4]) ? 4'b1100 : 4'b1000;
																assign node47097 = (inp[4]) ? 4'b1000 : 4'b1100;
													assign node47100 = (inp[3]) ? node47108 : node47101;
														assign node47101 = (inp[9]) ? 4'b1110 : node47102;
															assign node47102 = (inp[4]) ? node47104 : 4'b1000;
																assign node47104 = (inp[12]) ? 4'b1110 : 4'b1000;
														assign node47108 = (inp[12]) ? node47114 : node47109;
															assign node47109 = (inp[9]) ? node47111 : 4'b1110;
																assign node47111 = (inp[4]) ? 4'b1110 : 4'b1010;
															assign node47114 = (inp[9]) ? node47118 : node47115;
																assign node47115 = (inp[4]) ? 4'b1110 : 4'b1010;
																assign node47118 = (inp[4]) ? 4'b1010 : 4'b1110;
												assign node47121 = (inp[0]) ? node47145 : node47122;
													assign node47122 = (inp[3]) ? node47132 : node47123;
														assign node47123 = (inp[12]) ? node47125 : 4'b1100;
															assign node47125 = (inp[9]) ? node47129 : node47126;
																assign node47126 = (inp[4]) ? 4'b1110 : 4'b1000;
																assign node47129 = (inp[4]) ? 4'b1010 : 4'b1110;
														assign node47132 = (inp[12]) ? node47140 : node47133;
															assign node47133 = (inp[9]) ? node47137 : node47134;
																assign node47134 = (inp[4]) ? 4'b1010 : 4'b1110;
																assign node47137 = (inp[4]) ? 4'b1110 : 4'b1010;
															assign node47140 = (inp[9]) ? node47142 : 4'b1010;
																assign node47142 = (inp[4]) ? 4'b1010 : 4'b1110;
													assign node47145 = (inp[3]) ? node47155 : node47146;
														assign node47146 = (inp[4]) ? node47148 : 4'b1010;
															assign node47148 = (inp[9]) ? node47152 : node47149;
																assign node47149 = (inp[12]) ? 4'b1100 : 4'b1010;
																assign node47152 = (inp[12]) ? 4'b1000 : 4'b1100;
														assign node47155 = (inp[9]) ? 4'b1000 : node47156;
															assign node47156 = (inp[4]) ? 4'b1100 : node47157;
																assign node47157 = (inp[12]) ? 4'b1000 : 4'b1100;
											assign node47162 = (inp[12]) ? node47204 : node47163;
												assign node47163 = (inp[9]) ? node47187 : node47164;
													assign node47164 = (inp[4]) ? node47172 : node47165;
														assign node47165 = (inp[15]) ? node47167 : 4'b1111;
															assign node47167 = (inp[0]) ? 4'b1101 : node47168;
																assign node47168 = (inp[3]) ? 4'b1111 : 4'b1101;
														assign node47172 = (inp[0]) ? node47180 : node47173;
															assign node47173 = (inp[3]) ? node47177 : node47174;
																assign node47174 = (inp[15]) ? 4'b1001 : 4'b1011;
																assign node47177 = (inp[15]) ? 4'b1011 : 4'b1001;
															assign node47180 = (inp[3]) ? node47184 : node47181;
																assign node47181 = (inp[15]) ? 4'b1011 : 4'b1001;
																assign node47184 = (inp[15]) ? 4'b1001 : 4'b1011;
													assign node47187 = (inp[4]) ? node47197 : node47188;
														assign node47188 = (inp[3]) ? node47190 : 4'b1001;
															assign node47190 = (inp[0]) ? node47194 : node47191;
																assign node47191 = (inp[15]) ? 4'b1011 : 4'b1001;
																assign node47194 = (inp[15]) ? 4'b1001 : 4'b1011;
														assign node47197 = (inp[15]) ? node47201 : node47198;
															assign node47198 = (inp[0]) ? 4'b1111 : 4'b1101;
															assign node47201 = (inp[0]) ? 4'b1101 : 4'b1111;
												assign node47204 = (inp[0]) ? node47224 : node47205;
													assign node47205 = (inp[15]) ? node47215 : node47206;
														assign node47206 = (inp[9]) ? node47212 : node47207;
															assign node47207 = (inp[4]) ? 4'b1101 : node47208;
																assign node47208 = (inp[3]) ? 4'b1001 : 4'b1011;
															assign node47212 = (inp[4]) ? 4'b1001 : 4'b1101;
														assign node47215 = (inp[3]) ? 4'b1011 : node47216;
															assign node47216 = (inp[9]) ? node47220 : node47217;
																assign node47217 = (inp[4]) ? 4'b1111 : 4'b1001;
																assign node47220 = (inp[4]) ? 4'b1011 : 4'b1111;
													assign node47224 = (inp[15]) ? node47228 : node47225;
														assign node47225 = (inp[4]) ? 4'b1011 : 4'b1111;
														assign node47228 = (inp[4]) ? node47230 : 4'b1101;
															assign node47230 = (inp[9]) ? 4'b1001 : 4'b1101;
										assign node47233 = (inp[9]) ? node47315 : node47234;
											assign node47234 = (inp[3]) ? node47270 : node47235;
												assign node47235 = (inp[4]) ? node47253 : node47236;
													assign node47236 = (inp[12]) ? node47246 : node47237;
														assign node47237 = (inp[2]) ? node47239 : 4'b1111;
															assign node47239 = (inp[15]) ? node47243 : node47240;
																assign node47240 = (inp[0]) ? 4'b1101 : 4'b1111;
																assign node47243 = (inp[0]) ? 4'b1111 : 4'b1101;
														assign node47246 = (inp[15]) ? node47250 : node47247;
															assign node47247 = (inp[0]) ? 4'b1001 : 4'b1011;
															assign node47250 = (inp[0]) ? 4'b1011 : 4'b1001;
													assign node47253 = (inp[12]) ? node47263 : node47254;
														assign node47254 = (inp[2]) ? node47256 : 4'b1001;
															assign node47256 = (inp[15]) ? node47260 : node47257;
																assign node47257 = (inp[0]) ? 4'b1001 : 4'b1011;
																assign node47260 = (inp[0]) ? 4'b1011 : 4'b1001;
														assign node47263 = (inp[0]) ? node47267 : node47264;
															assign node47264 = (inp[15]) ? 4'b1111 : 4'b1101;
															assign node47267 = (inp[15]) ? 4'b1101 : 4'b1111;
												assign node47270 = (inp[2]) ? node47294 : node47271;
													assign node47271 = (inp[0]) ? node47285 : node47272;
														assign node47272 = (inp[15]) ? node47278 : node47273;
															assign node47273 = (inp[12]) ? node47275 : 4'b1101;
																assign node47275 = (inp[4]) ? 4'b1101 : 4'b1001;
															assign node47278 = (inp[12]) ? node47282 : node47279;
																assign node47279 = (inp[4]) ? 4'b1011 : 4'b1111;
																assign node47282 = (inp[4]) ? 4'b1111 : 4'b1011;
														assign node47285 = (inp[15]) ? 4'b1101 : node47286;
															assign node47286 = (inp[4]) ? node47290 : node47287;
																assign node47287 = (inp[12]) ? 4'b1011 : 4'b1111;
																assign node47290 = (inp[12]) ? 4'b1111 : 4'b1011;
													assign node47294 = (inp[4]) ? node47304 : node47295;
														assign node47295 = (inp[12]) ? 4'b1001 : node47296;
															assign node47296 = (inp[0]) ? node47300 : node47297;
																assign node47297 = (inp[15]) ? 4'b1111 : 4'b1101;
																assign node47300 = (inp[15]) ? 4'b1101 : 4'b1111;
														assign node47304 = (inp[12]) ? node47310 : node47305;
															assign node47305 = (inp[0]) ? node47307 : 4'b1001;
																assign node47307 = (inp[15]) ? 4'b1001 : 4'b1011;
															assign node47310 = (inp[0]) ? node47312 : 4'b1101;
																assign node47312 = (inp[15]) ? 4'b1101 : 4'b1111;
											assign node47315 = (inp[2]) ? node47367 : node47316;
												assign node47316 = (inp[0]) ? node47344 : node47317;
													assign node47317 = (inp[15]) ? node47329 : node47318;
														assign node47318 = (inp[3]) ? node47324 : node47319;
															assign node47319 = (inp[4]) ? node47321 : 4'b1011;
																assign node47321 = (inp[12]) ? 4'b1001 : 4'b1101;
															assign node47324 = (inp[4]) ? 4'b1001 : node47325;
																assign node47325 = (inp[12]) ? 4'b1101 : 4'b1001;
														assign node47329 = (inp[3]) ? node47337 : node47330;
															assign node47330 = (inp[4]) ? node47334 : node47331;
																assign node47331 = (inp[12]) ? 4'b1111 : 4'b1001;
																assign node47334 = (inp[12]) ? 4'b1011 : 4'b1111;
															assign node47337 = (inp[12]) ? node47341 : node47338;
																assign node47338 = (inp[4]) ? 4'b1111 : 4'b1011;
																assign node47341 = (inp[4]) ? 4'b1011 : 4'b1111;
													assign node47344 = (inp[15]) ? node47358 : node47345;
														assign node47345 = (inp[3]) ? node47351 : node47346;
															assign node47346 = (inp[4]) ? 4'b1111 : node47347;
																assign node47347 = (inp[12]) ? 4'b1111 : 4'b1001;
															assign node47351 = (inp[12]) ? node47355 : node47352;
																assign node47352 = (inp[4]) ? 4'b1111 : 4'b1011;
																assign node47355 = (inp[4]) ? 4'b1011 : 4'b1111;
														assign node47358 = (inp[4]) ? node47364 : node47359;
															assign node47359 = (inp[12]) ? 4'b1101 : node47360;
																assign node47360 = (inp[3]) ? 4'b1001 : 4'b1011;
															assign node47364 = (inp[12]) ? 4'b1001 : 4'b1101;
												assign node47367 = (inp[12]) ? node47389 : node47368;
													assign node47368 = (inp[4]) ? node47382 : node47369;
														assign node47369 = (inp[3]) ? node47375 : node47370;
															assign node47370 = (inp[0]) ? node47372 : 4'b1001;
																assign node47372 = (inp[15]) ? 4'b1011 : 4'b1001;
															assign node47375 = (inp[15]) ? node47379 : node47376;
																assign node47376 = (inp[0]) ? 4'b1011 : 4'b1001;
																assign node47379 = (inp[0]) ? 4'b1001 : 4'b1011;
														assign node47382 = (inp[0]) ? node47386 : node47383;
															assign node47383 = (inp[15]) ? 4'b1111 : 4'b1101;
															assign node47386 = (inp[15]) ? 4'b1101 : 4'b1111;
													assign node47389 = (inp[4]) ? node47397 : node47390;
														assign node47390 = (inp[15]) ? node47394 : node47391;
															assign node47391 = (inp[0]) ? 4'b1111 : 4'b1101;
															assign node47394 = (inp[0]) ? 4'b1101 : 4'b1111;
														assign node47397 = (inp[15]) ? node47401 : node47398;
															assign node47398 = (inp[0]) ? 4'b1011 : 4'b1001;
															assign node47401 = (inp[0]) ? 4'b1001 : 4'b1011;
								assign node47404 = (inp[8]) ? node47700 : node47405;
									assign node47405 = (inp[14]) ? node47559 : node47406;
										assign node47406 = (inp[2]) ? node47490 : node47407;
											assign node47407 = (inp[0]) ? node47447 : node47408;
												assign node47408 = (inp[15]) ? node47424 : node47409;
													assign node47409 = (inp[3]) ? node47415 : node47410;
														assign node47410 = (inp[9]) ? node47412 : 4'b1010;
															assign node47412 = (inp[4]) ? 4'b1000 : 4'b1100;
														assign node47415 = (inp[9]) ? node47417 : 4'b1100;
															assign node47417 = (inp[4]) ? node47421 : node47418;
																assign node47418 = (inp[12]) ? 4'b1100 : 4'b1000;
																assign node47421 = (inp[12]) ? 4'b1000 : 4'b1100;
													assign node47424 = (inp[3]) ? node47440 : node47425;
														assign node47425 = (inp[12]) ? node47433 : node47426;
															assign node47426 = (inp[9]) ? node47430 : node47427;
																assign node47427 = (inp[4]) ? 4'b1000 : 4'b1100;
																assign node47430 = (inp[4]) ? 4'b1110 : 4'b1000;
															assign node47433 = (inp[4]) ? node47437 : node47434;
																assign node47434 = (inp[9]) ? 4'b1110 : 4'b1000;
																assign node47437 = (inp[9]) ? 4'b1010 : 4'b1110;
														assign node47440 = (inp[4]) ? node47442 : 4'b1010;
															assign node47442 = (inp[12]) ? 4'b1110 : node47443;
																assign node47443 = (inp[9]) ? 4'b1110 : 4'b1010;
												assign node47447 = (inp[15]) ? node47473 : node47448;
													assign node47448 = (inp[3]) ? node47458 : node47449;
														assign node47449 = (inp[4]) ? node47453 : node47450;
															assign node47450 = (inp[9]) ? 4'b1110 : 4'b1000;
															assign node47453 = (inp[12]) ? node47455 : 4'b1110;
																assign node47455 = (inp[9]) ? 4'b1010 : 4'b1110;
														assign node47458 = (inp[12]) ? node47466 : node47459;
															assign node47459 = (inp[9]) ? node47463 : node47460;
																assign node47460 = (inp[4]) ? 4'b1010 : 4'b1110;
																assign node47463 = (inp[4]) ? 4'b1110 : 4'b1010;
															assign node47466 = (inp[9]) ? node47470 : node47467;
																assign node47467 = (inp[4]) ? 4'b1110 : 4'b1010;
																assign node47470 = (inp[4]) ? 4'b1010 : 4'b1110;
													assign node47473 = (inp[3]) ? node47483 : node47474;
														assign node47474 = (inp[4]) ? node47480 : node47475;
															assign node47475 = (inp[12]) ? 4'b1010 : node47476;
																assign node47476 = (inp[9]) ? 4'b1010 : 4'b1110;
															assign node47480 = (inp[12]) ? 4'b1000 : 4'b1100;
														assign node47483 = (inp[9]) ? node47485 : 4'b1100;
															assign node47485 = (inp[4]) ? 4'b1000 : node47486;
																assign node47486 = (inp[12]) ? 4'b1100 : 4'b1000;
											assign node47490 = (inp[12]) ? node47530 : node47491;
												assign node47491 = (inp[0]) ? node47513 : node47492;
													assign node47492 = (inp[15]) ? node47500 : node47493;
														assign node47493 = (inp[9]) ? node47497 : node47494;
															assign node47494 = (inp[3]) ? 4'b1001 : 4'b1011;
															assign node47497 = (inp[4]) ? 4'b1101 : 4'b1001;
														assign node47500 = (inp[3]) ? node47506 : node47501;
															assign node47501 = (inp[4]) ? node47503 : 4'b1001;
																assign node47503 = (inp[9]) ? 4'b1111 : 4'b1001;
															assign node47506 = (inp[4]) ? node47510 : node47507;
																assign node47507 = (inp[9]) ? 4'b1011 : 4'b1111;
																assign node47510 = (inp[9]) ? 4'b1111 : 4'b1011;
													assign node47513 = (inp[15]) ? node47519 : node47514;
														assign node47514 = (inp[3]) ? 4'b1111 : node47515;
															assign node47515 = (inp[4]) ? 4'b1001 : 4'b1101;
														assign node47519 = (inp[3]) ? node47523 : node47520;
															assign node47520 = (inp[9]) ? 4'b1101 : 4'b1111;
															assign node47523 = (inp[9]) ? node47527 : node47524;
																assign node47524 = (inp[4]) ? 4'b1001 : 4'b1101;
																assign node47527 = (inp[4]) ? 4'b1101 : 4'b1001;
												assign node47530 = (inp[9]) ? node47548 : node47531;
													assign node47531 = (inp[4]) ? node47541 : node47532;
														assign node47532 = (inp[0]) ? node47534 : 4'b1011;
															assign node47534 = (inp[3]) ? node47538 : node47535;
																assign node47535 = (inp[15]) ? 4'b1011 : 4'b1001;
																assign node47538 = (inp[15]) ? 4'b1001 : 4'b1011;
														assign node47541 = (inp[15]) ? node47545 : node47542;
															assign node47542 = (inp[3]) ? 4'b1111 : 4'b1101;
															assign node47545 = (inp[0]) ? 4'b1101 : 4'b1111;
													assign node47548 = (inp[4]) ? node47554 : node47549;
														assign node47549 = (inp[15]) ? 4'b1111 : node47550;
															assign node47550 = (inp[0]) ? 4'b1111 : 4'b1101;
														assign node47554 = (inp[0]) ? 4'b1011 : node47555;
															assign node47555 = (inp[15]) ? 4'b1011 : 4'b1001;
										assign node47559 = (inp[0]) ? node47639 : node47560;
											assign node47560 = (inp[15]) ? node47600 : node47561;
												assign node47561 = (inp[3]) ? node47577 : node47562;
													assign node47562 = (inp[9]) ? node47570 : node47563;
														assign node47563 = (inp[4]) ? node47567 : node47564;
															assign node47564 = (inp[12]) ? 4'b1011 : 4'b1111;
															assign node47567 = (inp[12]) ? 4'b1101 : 4'b1011;
														assign node47570 = (inp[4]) ? node47574 : node47571;
															assign node47571 = (inp[12]) ? 4'b1101 : 4'b1011;
															assign node47574 = (inp[12]) ? 4'b1001 : 4'b1101;
													assign node47577 = (inp[9]) ? node47591 : node47578;
														assign node47578 = (inp[2]) ? node47584 : node47579;
															assign node47579 = (inp[4]) ? 4'b1101 : node47580;
																assign node47580 = (inp[12]) ? 4'b1001 : 4'b1101;
															assign node47584 = (inp[12]) ? node47588 : node47585;
																assign node47585 = (inp[4]) ? 4'b1001 : 4'b1101;
																assign node47588 = (inp[4]) ? 4'b1101 : 4'b1001;
														assign node47591 = (inp[2]) ? node47593 : 4'b1001;
															assign node47593 = (inp[12]) ? node47597 : node47594;
																assign node47594 = (inp[4]) ? 4'b1101 : 4'b1001;
																assign node47597 = (inp[4]) ? 4'b1001 : 4'b1101;
												assign node47600 = (inp[3]) ? node47620 : node47601;
													assign node47601 = (inp[4]) ? node47609 : node47602;
														assign node47602 = (inp[9]) ? node47606 : node47603;
															assign node47603 = (inp[12]) ? 4'b1001 : 4'b1101;
															assign node47606 = (inp[12]) ? 4'b1111 : 4'b1001;
														assign node47609 = (inp[2]) ? node47615 : node47610;
															assign node47610 = (inp[9]) ? node47612 : 4'b1111;
																assign node47612 = (inp[12]) ? 4'b1011 : 4'b1111;
															assign node47615 = (inp[12]) ? node47617 : 4'b1001;
																assign node47617 = (inp[9]) ? 4'b1011 : 4'b1111;
													assign node47620 = (inp[4]) ? node47634 : node47621;
														assign node47621 = (inp[2]) ? node47629 : node47622;
															assign node47622 = (inp[12]) ? node47626 : node47623;
																assign node47623 = (inp[9]) ? 4'b1011 : 4'b1111;
																assign node47626 = (inp[9]) ? 4'b1111 : 4'b1011;
															assign node47629 = (inp[12]) ? node47631 : 4'b1111;
																assign node47631 = (inp[9]) ? 4'b1111 : 4'b1011;
														assign node47634 = (inp[9]) ? 4'b1011 : node47635;
															assign node47635 = (inp[12]) ? 4'b1111 : 4'b1011;
											assign node47639 = (inp[15]) ? node47673 : node47640;
												assign node47640 = (inp[3]) ? node47656 : node47641;
													assign node47641 = (inp[12]) ? node47649 : node47642;
														assign node47642 = (inp[4]) ? node47646 : node47643;
															assign node47643 = (inp[9]) ? 4'b1001 : 4'b1101;
															assign node47646 = (inp[9]) ? 4'b1111 : 4'b1001;
														assign node47649 = (inp[2]) ? node47651 : 4'b1111;
															assign node47651 = (inp[9]) ? node47653 : 4'b1001;
																assign node47653 = (inp[4]) ? 4'b1011 : 4'b1111;
													assign node47656 = (inp[9]) ? node47666 : node47657;
														assign node47657 = (inp[2]) ? node47659 : 4'b1011;
															assign node47659 = (inp[4]) ? node47663 : node47660;
																assign node47660 = (inp[12]) ? 4'b1011 : 4'b1111;
																assign node47663 = (inp[12]) ? 4'b1111 : 4'b1011;
														assign node47666 = (inp[4]) ? node47670 : node47667;
															assign node47667 = (inp[12]) ? 4'b1111 : 4'b1011;
															assign node47670 = (inp[12]) ? 4'b1011 : 4'b1111;
												assign node47673 = (inp[3]) ? node47683 : node47674;
													assign node47674 = (inp[4]) ? 4'b1101 : node47675;
														assign node47675 = (inp[12]) ? node47679 : node47676;
															assign node47676 = (inp[9]) ? 4'b1011 : 4'b1111;
															assign node47679 = (inp[9]) ? 4'b1101 : 4'b1011;
													assign node47683 = (inp[2]) ? node47691 : node47684;
														assign node47684 = (inp[12]) ? 4'b1101 : node47685;
															assign node47685 = (inp[9]) ? node47687 : 4'b1101;
																assign node47687 = (inp[4]) ? 4'b1101 : 4'b1001;
														assign node47691 = (inp[9]) ? node47693 : 4'b1001;
															assign node47693 = (inp[4]) ? node47697 : node47694;
																assign node47694 = (inp[12]) ? 4'b1101 : 4'b1001;
																assign node47697 = (inp[12]) ? 4'b1001 : 4'b1101;
									assign node47700 = (inp[14]) ? node47886 : node47701;
										assign node47701 = (inp[2]) ? node47803 : node47702;
											assign node47702 = (inp[15]) ? node47758 : node47703;
												assign node47703 = (inp[0]) ? node47729 : node47704;
													assign node47704 = (inp[3]) ? node47718 : node47705;
														assign node47705 = (inp[9]) ? node47713 : node47706;
															assign node47706 = (inp[12]) ? node47710 : node47707;
																assign node47707 = (inp[4]) ? 4'b1011 : 4'b1111;
																assign node47710 = (inp[4]) ? 4'b1101 : 4'b1011;
															assign node47713 = (inp[4]) ? 4'b1101 : node47714;
																assign node47714 = (inp[12]) ? 4'b1101 : 4'b1011;
														assign node47718 = (inp[12]) ? node47724 : node47719;
															assign node47719 = (inp[9]) ? 4'b1101 : node47720;
																assign node47720 = (inp[4]) ? 4'b1001 : 4'b1101;
															assign node47724 = (inp[9]) ? node47726 : 4'b1001;
																assign node47726 = (inp[4]) ? 4'b1001 : 4'b1101;
													assign node47729 = (inp[3]) ? node47745 : node47730;
														assign node47730 = (inp[4]) ? node47738 : node47731;
															assign node47731 = (inp[12]) ? node47735 : node47732;
																assign node47732 = (inp[9]) ? 4'b1001 : 4'b1101;
																assign node47735 = (inp[9]) ? 4'b1111 : 4'b1001;
															assign node47738 = (inp[12]) ? node47742 : node47739;
																assign node47739 = (inp[9]) ? 4'b1111 : 4'b1001;
																assign node47742 = (inp[9]) ? 4'b1011 : 4'b1111;
														assign node47745 = (inp[12]) ? node47751 : node47746;
															assign node47746 = (inp[9]) ? node47748 : 4'b1011;
																assign node47748 = (inp[4]) ? 4'b1111 : 4'b1011;
															assign node47751 = (inp[4]) ? node47755 : node47752;
																assign node47752 = (inp[9]) ? 4'b1111 : 4'b1011;
																assign node47755 = (inp[9]) ? 4'b1011 : 4'b1111;
												assign node47758 = (inp[0]) ? node47776 : node47759;
													assign node47759 = (inp[3]) ? node47769 : node47760;
														assign node47760 = (inp[12]) ? node47766 : node47761;
															assign node47761 = (inp[4]) ? 4'b1001 : node47762;
																assign node47762 = (inp[9]) ? 4'b1001 : 4'b1101;
															assign node47766 = (inp[4]) ? 4'b1011 : 4'b1001;
														assign node47769 = (inp[12]) ? 4'b1111 : node47770;
															assign node47770 = (inp[4]) ? 4'b1011 : node47771;
																assign node47771 = (inp[9]) ? 4'b1011 : 4'b1111;
													assign node47776 = (inp[3]) ? node47790 : node47777;
														assign node47777 = (inp[9]) ? node47783 : node47778;
															assign node47778 = (inp[4]) ? 4'b1011 : node47779;
																assign node47779 = (inp[12]) ? 4'b1011 : 4'b1111;
															assign node47783 = (inp[12]) ? node47787 : node47784;
																assign node47784 = (inp[4]) ? 4'b1101 : 4'b1011;
																assign node47787 = (inp[4]) ? 4'b1001 : 4'b1101;
														assign node47790 = (inp[4]) ? node47798 : node47791;
															assign node47791 = (inp[12]) ? node47795 : node47792;
																assign node47792 = (inp[9]) ? 4'b1001 : 4'b1101;
																assign node47795 = (inp[9]) ? 4'b1101 : 4'b1001;
															assign node47798 = (inp[12]) ? 4'b1001 : node47799;
																assign node47799 = (inp[9]) ? 4'b1101 : 4'b1001;
											assign node47803 = (inp[3]) ? node47841 : node47804;
												assign node47804 = (inp[0]) ? node47822 : node47805;
													assign node47805 = (inp[12]) ? node47809 : node47806;
														assign node47806 = (inp[15]) ? 4'b1000 : 4'b1010;
														assign node47809 = (inp[15]) ? node47817 : node47810;
															assign node47810 = (inp[9]) ? node47814 : node47811;
																assign node47811 = (inp[4]) ? 4'b1100 : 4'b1010;
																assign node47814 = (inp[4]) ? 4'b1000 : 4'b1100;
															assign node47817 = (inp[4]) ? node47819 : 4'b1000;
																assign node47819 = (inp[9]) ? 4'b1010 : 4'b1110;
													assign node47822 = (inp[9]) ? node47828 : node47823;
														assign node47823 = (inp[15]) ? 4'b1100 : node47824;
															assign node47824 = (inp[12]) ? 4'b1000 : 4'b1100;
														assign node47828 = (inp[15]) ? node47834 : node47829;
															assign node47829 = (inp[4]) ? node47831 : 4'b1000;
																assign node47831 = (inp[12]) ? 4'b1010 : 4'b1110;
															assign node47834 = (inp[12]) ? node47838 : node47835;
																assign node47835 = (inp[4]) ? 4'b1100 : 4'b1010;
																assign node47838 = (inp[4]) ? 4'b1000 : 4'b1100;
												assign node47841 = (inp[12]) ? node47859 : node47842;
													assign node47842 = (inp[0]) ? node47850 : node47843;
														assign node47843 = (inp[15]) ? node47845 : 4'b1100;
															assign node47845 = (inp[9]) ? node47847 : 4'b1110;
																assign node47847 = (inp[4]) ? 4'b1110 : 4'b1010;
														assign node47850 = (inp[15]) ? node47856 : node47851;
															assign node47851 = (inp[4]) ? 4'b1010 : node47852;
																assign node47852 = (inp[9]) ? 4'b1010 : 4'b1110;
															assign node47856 = (inp[9]) ? 4'b1000 : 4'b1100;
													assign node47859 = (inp[15]) ? node47873 : node47860;
														assign node47860 = (inp[0]) ? node47866 : node47861;
															assign node47861 = (inp[4]) ? 4'b1000 : node47862;
																assign node47862 = (inp[9]) ? 4'b1100 : 4'b1000;
															assign node47866 = (inp[9]) ? node47870 : node47867;
																assign node47867 = (inp[4]) ? 4'b1110 : 4'b1010;
																assign node47870 = (inp[4]) ? 4'b1010 : 4'b1110;
														assign node47873 = (inp[0]) ? node47881 : node47874;
															assign node47874 = (inp[9]) ? node47878 : node47875;
																assign node47875 = (inp[4]) ? 4'b1110 : 4'b1010;
																assign node47878 = (inp[4]) ? 4'b1010 : 4'b1110;
															assign node47881 = (inp[4]) ? node47883 : 4'b1000;
																assign node47883 = (inp[9]) ? 4'b1000 : 4'b1100;
										assign node47886 = (inp[0]) ? node47958 : node47887;
											assign node47887 = (inp[15]) ? node47921 : node47888;
												assign node47888 = (inp[3]) ? node47904 : node47889;
													assign node47889 = (inp[12]) ? node47897 : node47890;
														assign node47890 = (inp[2]) ? 4'b1010 : node47891;
															assign node47891 = (inp[9]) ? 4'b1010 : node47892;
																assign node47892 = (inp[4]) ? 4'b1010 : 4'b1110;
														assign node47897 = (inp[9]) ? node47901 : node47898;
															assign node47898 = (inp[4]) ? 4'b1100 : 4'b1010;
															assign node47901 = (inp[4]) ? 4'b1000 : 4'b1100;
													assign node47904 = (inp[9]) ? node47912 : node47905;
														assign node47905 = (inp[4]) ? node47909 : node47906;
															assign node47906 = (inp[12]) ? 4'b1000 : 4'b1100;
															assign node47909 = (inp[12]) ? 4'b1100 : 4'b1000;
														assign node47912 = (inp[2]) ? node47914 : 4'b1000;
															assign node47914 = (inp[12]) ? node47918 : node47915;
																assign node47915 = (inp[4]) ? 4'b1100 : 4'b1000;
																assign node47918 = (inp[4]) ? 4'b1000 : 4'b1100;
												assign node47921 = (inp[3]) ? node47935 : node47922;
													assign node47922 = (inp[12]) ? node47928 : node47923;
														assign node47923 = (inp[4]) ? 4'b1000 : node47924;
															assign node47924 = (inp[9]) ? 4'b1000 : 4'b1100;
														assign node47928 = (inp[9]) ? node47932 : node47929;
															assign node47929 = (inp[4]) ? 4'b1110 : 4'b1000;
															assign node47932 = (inp[4]) ? 4'b1010 : 4'b1110;
													assign node47935 = (inp[2]) ? node47949 : node47936;
														assign node47936 = (inp[9]) ? node47942 : node47937;
															assign node47937 = (inp[12]) ? node47939 : 4'b1010;
																assign node47939 = (inp[4]) ? 4'b1110 : 4'b1010;
															assign node47942 = (inp[4]) ? node47946 : node47943;
																assign node47943 = (inp[12]) ? 4'b1110 : 4'b1010;
																assign node47946 = (inp[12]) ? 4'b1010 : 4'b1110;
														assign node47949 = (inp[4]) ? node47951 : 4'b1110;
															assign node47951 = (inp[12]) ? node47955 : node47952;
																assign node47952 = (inp[9]) ? 4'b1110 : 4'b1010;
																assign node47955 = (inp[9]) ? 4'b1010 : 4'b1110;
											assign node47958 = (inp[15]) ? node47990 : node47959;
												assign node47959 = (inp[3]) ? node47975 : node47960;
													assign node47960 = (inp[9]) ? node47968 : node47961;
														assign node47961 = (inp[12]) ? node47965 : node47962;
															assign node47962 = (inp[4]) ? 4'b1000 : 4'b1100;
															assign node47965 = (inp[4]) ? 4'b1110 : 4'b1000;
														assign node47968 = (inp[4]) ? node47972 : node47969;
															assign node47969 = (inp[12]) ? 4'b1110 : 4'b1000;
															assign node47972 = (inp[12]) ? 4'b1010 : 4'b1110;
													assign node47975 = (inp[4]) ? node47983 : node47976;
														assign node47976 = (inp[9]) ? node47980 : node47977;
															assign node47977 = (inp[12]) ? 4'b1010 : 4'b1110;
															assign node47980 = (inp[12]) ? 4'b1110 : 4'b1010;
														assign node47983 = (inp[9]) ? node47987 : node47984;
															assign node47984 = (inp[12]) ? 4'b1110 : 4'b1010;
															assign node47987 = (inp[12]) ? 4'b1010 : 4'b1110;
												assign node47990 = (inp[3]) ? node48006 : node47991;
													assign node47991 = (inp[12]) ? node47999 : node47992;
														assign node47992 = (inp[4]) ? node47996 : node47993;
															assign node47993 = (inp[9]) ? 4'b1010 : 4'b1110;
															assign node47996 = (inp[9]) ? 4'b1100 : 4'b1010;
														assign node47999 = (inp[9]) ? node48003 : node48000;
															assign node48000 = (inp[4]) ? 4'b1100 : 4'b1010;
															assign node48003 = (inp[4]) ? 4'b1000 : 4'b1100;
													assign node48006 = (inp[9]) ? node48016 : node48007;
														assign node48007 = (inp[2]) ? 4'b1000 : node48008;
															assign node48008 = (inp[4]) ? node48012 : node48009;
																assign node48009 = (inp[12]) ? 4'b1000 : 4'b1100;
																assign node48012 = (inp[12]) ? 4'b1100 : 4'b1000;
														assign node48016 = (inp[2]) ? node48022 : node48017;
															assign node48017 = (inp[12]) ? 4'b1100 : node48018;
																assign node48018 = (inp[4]) ? 4'b1100 : 4'b1000;
															assign node48022 = (inp[12]) ? node48026 : node48023;
																assign node48023 = (inp[4]) ? 4'b1100 : 4'b1000;
																assign node48026 = (inp[4]) ? 4'b1000 : 4'b1100;
						assign node48029 = (inp[3]) ? node49059 : node48030;
							assign node48030 = (inp[2]) ? node48658 : node48031;
								assign node48031 = (inp[5]) ? node48353 : node48032;
									assign node48032 = (inp[0]) ? node48190 : node48033;
										assign node48033 = (inp[15]) ? node48113 : node48034;
											assign node48034 = (inp[9]) ? node48082 : node48035;
												assign node48035 = (inp[4]) ? node48059 : node48036;
													assign node48036 = (inp[7]) ? node48050 : node48037;
														assign node48037 = (inp[12]) ? node48045 : node48038;
															assign node48038 = (inp[14]) ? node48042 : node48039;
																assign node48039 = (inp[8]) ? 4'b1010 : 4'b1011;
																assign node48042 = (inp[8]) ? 4'b1011 : 4'b1010;
															assign node48045 = (inp[14]) ? node48047 : 4'b1010;
																assign node48047 = (inp[8]) ? 4'b1011 : 4'b1010;
														assign node48050 = (inp[12]) ? 4'b1011 : node48051;
															assign node48051 = (inp[8]) ? node48055 : node48052;
																assign node48052 = (inp[14]) ? 4'b1011 : 4'b1010;
																assign node48055 = (inp[14]) ? 4'b1010 : 4'b1011;
													assign node48059 = (inp[8]) ? node48067 : node48060;
														assign node48060 = (inp[7]) ? node48064 : node48061;
															assign node48061 = (inp[14]) ? 4'b1110 : 4'b1111;
															assign node48064 = (inp[14]) ? 4'b1111 : 4'b1110;
														assign node48067 = (inp[12]) ? node48075 : node48068;
															assign node48068 = (inp[14]) ? node48072 : node48069;
																assign node48069 = (inp[7]) ? 4'b1111 : 4'b1110;
																assign node48072 = (inp[7]) ? 4'b1110 : 4'b1111;
															assign node48075 = (inp[14]) ? node48079 : node48076;
																assign node48076 = (inp[7]) ? 4'b1111 : 4'b1110;
																assign node48079 = (inp[7]) ? 4'b1110 : 4'b1111;
												assign node48082 = (inp[4]) ? node48098 : node48083;
													assign node48083 = (inp[7]) ? node48091 : node48084;
														assign node48084 = (inp[14]) ? node48088 : node48085;
															assign node48085 = (inp[8]) ? 4'b1110 : 4'b1111;
															assign node48088 = (inp[8]) ? 4'b1111 : 4'b1110;
														assign node48091 = (inp[8]) ? node48095 : node48092;
															assign node48092 = (inp[14]) ? 4'b1111 : 4'b1110;
															assign node48095 = (inp[14]) ? 4'b1110 : 4'b1111;
													assign node48098 = (inp[7]) ? node48106 : node48099;
														assign node48099 = (inp[14]) ? node48103 : node48100;
															assign node48100 = (inp[8]) ? 4'b1010 : 4'b1011;
															assign node48103 = (inp[8]) ? 4'b1011 : 4'b1010;
														assign node48106 = (inp[14]) ? node48110 : node48107;
															assign node48107 = (inp[8]) ? 4'b1011 : 4'b1010;
															assign node48110 = (inp[8]) ? 4'b1010 : 4'b1011;
											assign node48113 = (inp[9]) ? node48153 : node48114;
												assign node48114 = (inp[4]) ? node48140 : node48115;
													assign node48115 = (inp[12]) ? node48125 : node48116;
														assign node48116 = (inp[7]) ? node48118 : 4'b1001;
															assign node48118 = (inp[8]) ? node48122 : node48119;
																assign node48119 = (inp[14]) ? 4'b1001 : 4'b1000;
																assign node48122 = (inp[14]) ? 4'b1000 : 4'b1001;
														assign node48125 = (inp[14]) ? node48133 : node48126;
															assign node48126 = (inp[8]) ? node48130 : node48127;
																assign node48127 = (inp[7]) ? 4'b1000 : 4'b1001;
																assign node48130 = (inp[7]) ? 4'b1001 : 4'b1000;
															assign node48133 = (inp[7]) ? node48137 : node48134;
																assign node48134 = (inp[8]) ? 4'b1001 : 4'b1000;
																assign node48137 = (inp[8]) ? 4'b1000 : 4'b1001;
													assign node48140 = (inp[8]) ? node48148 : node48141;
														assign node48141 = (inp[7]) ? node48145 : node48142;
															assign node48142 = (inp[12]) ? 4'b1101 : 4'b1100;
															assign node48145 = (inp[14]) ? 4'b1101 : 4'b1100;
														assign node48148 = (inp[14]) ? 4'b1100 : node48149;
															assign node48149 = (inp[7]) ? 4'b1101 : 4'b1100;
												assign node48153 = (inp[4]) ? node48171 : node48154;
													assign node48154 = (inp[12]) ? node48156 : 4'b1101;
														assign node48156 = (inp[7]) ? node48164 : node48157;
															assign node48157 = (inp[14]) ? node48161 : node48158;
																assign node48158 = (inp[8]) ? 4'b1100 : 4'b1101;
																assign node48161 = (inp[8]) ? 4'b1101 : 4'b1100;
															assign node48164 = (inp[14]) ? node48168 : node48165;
																assign node48165 = (inp[8]) ? 4'b1101 : 4'b1100;
																assign node48168 = (inp[8]) ? 4'b1100 : 4'b1101;
													assign node48171 = (inp[14]) ? node48183 : node48172;
														assign node48172 = (inp[12]) ? node48178 : node48173;
															assign node48173 = (inp[8]) ? 4'b1000 : node48174;
																assign node48174 = (inp[7]) ? 4'b1000 : 4'b1001;
															assign node48178 = (inp[8]) ? node48180 : 4'b1001;
																assign node48180 = (inp[7]) ? 4'b1001 : 4'b1000;
														assign node48183 = (inp[8]) ? node48187 : node48184;
															assign node48184 = (inp[7]) ? 4'b1001 : 4'b1000;
															assign node48187 = (inp[7]) ? 4'b1000 : 4'b1001;
										assign node48190 = (inp[15]) ? node48278 : node48191;
											assign node48191 = (inp[8]) ? node48235 : node48192;
												assign node48192 = (inp[12]) ? node48222 : node48193;
													assign node48193 = (inp[4]) ? node48207 : node48194;
														assign node48194 = (inp[9]) ? node48200 : node48195;
															assign node48195 = (inp[14]) ? 4'b1000 : node48196;
																assign node48196 = (inp[7]) ? 4'b1000 : 4'b1001;
															assign node48200 = (inp[14]) ? node48204 : node48201;
																assign node48201 = (inp[7]) ? 4'b1100 : 4'b1101;
																assign node48204 = (inp[7]) ? 4'b1101 : 4'b1100;
														assign node48207 = (inp[9]) ? node48215 : node48208;
															assign node48208 = (inp[14]) ? node48212 : node48209;
																assign node48209 = (inp[7]) ? 4'b1100 : 4'b1101;
																assign node48212 = (inp[7]) ? 4'b1101 : 4'b1100;
															assign node48215 = (inp[14]) ? node48219 : node48216;
																assign node48216 = (inp[7]) ? 4'b1000 : 4'b1001;
																assign node48219 = (inp[7]) ? 4'b1001 : 4'b1000;
													assign node48222 = (inp[14]) ? node48232 : node48223;
														assign node48223 = (inp[7]) ? node48227 : node48224;
															assign node48224 = (inp[4]) ? 4'b1001 : 4'b1101;
															assign node48227 = (inp[4]) ? 4'b1100 : node48228;
																assign node48228 = (inp[9]) ? 4'b1100 : 4'b1000;
														assign node48232 = (inp[7]) ? 4'b1101 : 4'b1100;
												assign node48235 = (inp[12]) ? node48261 : node48236;
													assign node48236 = (inp[9]) ? node48248 : node48237;
														assign node48237 = (inp[4]) ? node48243 : node48238;
															assign node48238 = (inp[7]) ? node48240 : 4'b1001;
																assign node48240 = (inp[14]) ? 4'b1000 : 4'b1001;
															assign node48243 = (inp[7]) ? 4'b1101 : node48244;
																assign node48244 = (inp[14]) ? 4'b1101 : 4'b1100;
														assign node48248 = (inp[4]) ? node48254 : node48249;
															assign node48249 = (inp[14]) ? 4'b1100 : node48250;
																assign node48250 = (inp[7]) ? 4'b1101 : 4'b1100;
															assign node48254 = (inp[14]) ? node48258 : node48255;
																assign node48255 = (inp[7]) ? 4'b1001 : 4'b1000;
																assign node48258 = (inp[7]) ? 4'b1000 : 4'b1001;
													assign node48261 = (inp[9]) ? node48265 : node48262;
														assign node48262 = (inp[4]) ? 4'b1100 : 4'b1000;
														assign node48265 = (inp[4]) ? node48271 : node48266;
															assign node48266 = (inp[14]) ? node48268 : 4'b1101;
																assign node48268 = (inp[7]) ? 4'b1100 : 4'b1101;
															assign node48271 = (inp[14]) ? node48275 : node48272;
																assign node48272 = (inp[7]) ? 4'b1001 : 4'b1000;
																assign node48275 = (inp[7]) ? 4'b1000 : 4'b1001;
											assign node48278 = (inp[8]) ? node48322 : node48279;
												assign node48279 = (inp[4]) ? node48301 : node48280;
													assign node48280 = (inp[9]) ? node48288 : node48281;
														assign node48281 = (inp[14]) ? node48285 : node48282;
															assign node48282 = (inp[7]) ? 4'b1010 : 4'b1011;
															assign node48285 = (inp[7]) ? 4'b1011 : 4'b1010;
														assign node48288 = (inp[12]) ? node48294 : node48289;
															assign node48289 = (inp[7]) ? node48291 : 4'b1110;
																assign node48291 = (inp[14]) ? 4'b1111 : 4'b1110;
															assign node48294 = (inp[7]) ? node48298 : node48295;
																assign node48295 = (inp[14]) ? 4'b1110 : 4'b1111;
																assign node48298 = (inp[14]) ? 4'b1111 : 4'b1110;
													assign node48301 = (inp[9]) ? node48317 : node48302;
														assign node48302 = (inp[12]) ? node48310 : node48303;
															assign node48303 = (inp[14]) ? node48307 : node48304;
																assign node48304 = (inp[7]) ? 4'b1110 : 4'b1111;
																assign node48307 = (inp[7]) ? 4'b1111 : 4'b1110;
															assign node48310 = (inp[14]) ? node48314 : node48311;
																assign node48311 = (inp[7]) ? 4'b1110 : 4'b1111;
																assign node48314 = (inp[7]) ? 4'b1111 : 4'b1110;
														assign node48317 = (inp[14]) ? 4'b1011 : node48318;
															assign node48318 = (inp[7]) ? 4'b1010 : 4'b1011;
												assign node48322 = (inp[9]) ? node48338 : node48323;
													assign node48323 = (inp[4]) ? node48331 : node48324;
														assign node48324 = (inp[14]) ? node48328 : node48325;
															assign node48325 = (inp[7]) ? 4'b1011 : 4'b1010;
															assign node48328 = (inp[7]) ? 4'b1010 : 4'b1011;
														assign node48331 = (inp[7]) ? node48335 : node48332;
															assign node48332 = (inp[14]) ? 4'b1111 : 4'b1110;
															assign node48335 = (inp[14]) ? 4'b1110 : 4'b1111;
													assign node48338 = (inp[4]) ? node48346 : node48339;
														assign node48339 = (inp[14]) ? node48343 : node48340;
															assign node48340 = (inp[7]) ? 4'b1111 : 4'b1110;
															assign node48343 = (inp[7]) ? 4'b1110 : 4'b1111;
														assign node48346 = (inp[14]) ? node48350 : node48347;
															assign node48347 = (inp[7]) ? 4'b1011 : 4'b1010;
															assign node48350 = (inp[7]) ? 4'b1010 : 4'b1011;
									assign node48353 = (inp[9]) ? node48517 : node48354;
										assign node48354 = (inp[4]) ? node48430 : node48355;
											assign node48355 = (inp[8]) ? node48401 : node48356;
												assign node48356 = (inp[12]) ? node48376 : node48357;
													assign node48357 = (inp[7]) ? node48367 : node48358;
														assign node48358 = (inp[14]) ? node48360 : 4'b1011;
															assign node48360 = (inp[0]) ? node48364 : node48361;
																assign node48361 = (inp[15]) ? 4'b1000 : 4'b1010;
																assign node48364 = (inp[15]) ? 4'b1010 : 4'b1000;
														assign node48367 = (inp[14]) ? 4'b1011 : node48368;
															assign node48368 = (inp[15]) ? node48372 : node48369;
																assign node48369 = (inp[0]) ? 4'b1000 : 4'b1010;
																assign node48372 = (inp[0]) ? 4'b1010 : 4'b1000;
													assign node48376 = (inp[7]) ? node48390 : node48377;
														assign node48377 = (inp[14]) ? node48383 : node48378;
															assign node48378 = (inp[15]) ? 4'b1001 : node48379;
																assign node48379 = (inp[0]) ? 4'b1001 : 4'b1011;
															assign node48383 = (inp[15]) ? node48387 : node48384;
																assign node48384 = (inp[0]) ? 4'b1000 : 4'b1010;
																assign node48387 = (inp[0]) ? 4'b1010 : 4'b1000;
														assign node48390 = (inp[14]) ? node48394 : node48391;
															assign node48391 = (inp[15]) ? 4'b1010 : 4'b1000;
															assign node48394 = (inp[15]) ? node48398 : node48395;
																assign node48395 = (inp[0]) ? 4'b1001 : 4'b1011;
																assign node48398 = (inp[0]) ? 4'b1011 : 4'b1001;
												assign node48401 = (inp[7]) ? node48417 : node48402;
													assign node48402 = (inp[14]) ? node48410 : node48403;
														assign node48403 = (inp[15]) ? node48407 : node48404;
															assign node48404 = (inp[0]) ? 4'b1000 : 4'b1010;
															assign node48407 = (inp[0]) ? 4'b1010 : 4'b1000;
														assign node48410 = (inp[15]) ? node48414 : node48411;
															assign node48411 = (inp[0]) ? 4'b1001 : 4'b1011;
															assign node48414 = (inp[0]) ? 4'b1011 : 4'b1001;
													assign node48417 = (inp[14]) ? node48425 : node48418;
														assign node48418 = (inp[15]) ? node48422 : node48419;
															assign node48419 = (inp[0]) ? 4'b1001 : 4'b1011;
															assign node48422 = (inp[0]) ? 4'b1011 : 4'b1001;
														assign node48425 = (inp[15]) ? 4'b1000 : node48426;
															assign node48426 = (inp[0]) ? 4'b1000 : 4'b1010;
											assign node48430 = (inp[8]) ? node48470 : node48431;
												assign node48431 = (inp[7]) ? node48453 : node48432;
													assign node48432 = (inp[14]) ? node48440 : node48433;
														assign node48433 = (inp[15]) ? node48437 : node48434;
															assign node48434 = (inp[0]) ? 4'b1111 : 4'b1101;
															assign node48437 = (inp[0]) ? 4'b1101 : 4'b1111;
														assign node48440 = (inp[12]) ? node48446 : node48441;
															assign node48441 = (inp[0]) ? 4'b1100 : node48442;
																assign node48442 = (inp[15]) ? 4'b1110 : 4'b1100;
															assign node48446 = (inp[15]) ? node48450 : node48447;
																assign node48447 = (inp[0]) ? 4'b1110 : 4'b1100;
																assign node48450 = (inp[0]) ? 4'b1100 : 4'b1110;
													assign node48453 = (inp[14]) ? node48465 : node48454;
														assign node48454 = (inp[12]) ? node48460 : node48455;
															assign node48455 = (inp[15]) ? 4'b1100 : node48456;
																assign node48456 = (inp[0]) ? 4'b1110 : 4'b1100;
															assign node48460 = (inp[0]) ? 4'b1100 : node48461;
																assign node48461 = (inp[15]) ? 4'b1110 : 4'b1100;
														assign node48465 = (inp[0]) ? node48467 : 4'b1101;
															assign node48467 = (inp[15]) ? 4'b1101 : 4'b1111;
												assign node48470 = (inp[12]) ? node48492 : node48471;
													assign node48471 = (inp[14]) ? node48481 : node48472;
														assign node48472 = (inp[7]) ? node48474 : 4'b1100;
															assign node48474 = (inp[15]) ? node48478 : node48475;
																assign node48475 = (inp[0]) ? 4'b1111 : 4'b1101;
																assign node48478 = (inp[0]) ? 4'b1101 : 4'b1111;
														assign node48481 = (inp[7]) ? node48487 : node48482;
															assign node48482 = (inp[15]) ? node48484 : 4'b1111;
																assign node48484 = (inp[0]) ? 4'b1101 : 4'b1111;
															assign node48487 = (inp[15]) ? 4'b1100 : node48488;
																assign node48488 = (inp[0]) ? 4'b1110 : 4'b1100;
													assign node48492 = (inp[0]) ? node48504 : node48493;
														assign node48493 = (inp[15]) ? node48497 : node48494;
															assign node48494 = (inp[7]) ? 4'b1101 : 4'b1100;
															assign node48497 = (inp[14]) ? node48501 : node48498;
																assign node48498 = (inp[7]) ? 4'b1111 : 4'b1110;
																assign node48501 = (inp[7]) ? 4'b1110 : 4'b1111;
														assign node48504 = (inp[15]) ? node48510 : node48505;
															assign node48505 = (inp[7]) ? 4'b1111 : node48506;
																assign node48506 = (inp[14]) ? 4'b1111 : 4'b1110;
															assign node48510 = (inp[14]) ? node48514 : node48511;
																assign node48511 = (inp[7]) ? 4'b1101 : 4'b1100;
																assign node48514 = (inp[7]) ? 4'b1100 : 4'b1101;
										assign node48517 = (inp[4]) ? node48593 : node48518;
											assign node48518 = (inp[15]) ? node48556 : node48519;
												assign node48519 = (inp[0]) ? node48533 : node48520;
													assign node48520 = (inp[14]) ? node48526 : node48521;
														assign node48521 = (inp[7]) ? node48523 : 4'b1101;
															assign node48523 = (inp[8]) ? 4'b1101 : 4'b1100;
														assign node48526 = (inp[8]) ? node48530 : node48527;
															assign node48527 = (inp[7]) ? 4'b1101 : 4'b1100;
															assign node48530 = (inp[7]) ? 4'b1100 : 4'b1101;
													assign node48533 = (inp[7]) ? node48541 : node48534;
														assign node48534 = (inp[8]) ? node48538 : node48535;
															assign node48535 = (inp[14]) ? 4'b1110 : 4'b1111;
															assign node48538 = (inp[14]) ? 4'b1111 : 4'b1110;
														assign node48541 = (inp[12]) ? node48549 : node48542;
															assign node48542 = (inp[8]) ? node48546 : node48543;
																assign node48543 = (inp[14]) ? 4'b1111 : 4'b1110;
																assign node48546 = (inp[14]) ? 4'b1110 : 4'b1111;
															assign node48549 = (inp[14]) ? node48553 : node48550;
																assign node48550 = (inp[8]) ? 4'b1111 : 4'b1110;
																assign node48553 = (inp[8]) ? 4'b1110 : 4'b1111;
												assign node48556 = (inp[0]) ? node48572 : node48557;
													assign node48557 = (inp[14]) ? node48565 : node48558;
														assign node48558 = (inp[8]) ? node48562 : node48559;
															assign node48559 = (inp[7]) ? 4'b1110 : 4'b1111;
															assign node48562 = (inp[7]) ? 4'b1111 : 4'b1110;
														assign node48565 = (inp[7]) ? node48569 : node48566;
															assign node48566 = (inp[8]) ? 4'b1111 : 4'b1110;
															assign node48569 = (inp[8]) ? 4'b1110 : 4'b1111;
													assign node48572 = (inp[8]) ? node48586 : node48573;
														assign node48573 = (inp[12]) ? node48581 : node48574;
															assign node48574 = (inp[7]) ? node48578 : node48575;
																assign node48575 = (inp[14]) ? 4'b1100 : 4'b1101;
																assign node48578 = (inp[14]) ? 4'b1101 : 4'b1100;
															assign node48581 = (inp[14]) ? 4'b1101 : node48582;
																assign node48582 = (inp[7]) ? 4'b1100 : 4'b1101;
														assign node48586 = (inp[7]) ? node48590 : node48587;
															assign node48587 = (inp[14]) ? 4'b1101 : 4'b1100;
															assign node48590 = (inp[14]) ? 4'b1100 : 4'b1101;
											assign node48593 = (inp[8]) ? node48631 : node48594;
												assign node48594 = (inp[12]) ? node48616 : node48595;
													assign node48595 = (inp[15]) ? node48609 : node48596;
														assign node48596 = (inp[0]) ? node48602 : node48597;
															assign node48597 = (inp[14]) ? node48599 : 4'b1001;
																assign node48599 = (inp[7]) ? 4'b1001 : 4'b1000;
															assign node48602 = (inp[14]) ? node48606 : node48603;
																assign node48603 = (inp[7]) ? 4'b1010 : 4'b1011;
																assign node48606 = (inp[7]) ? 4'b1011 : 4'b1010;
														assign node48609 = (inp[0]) ? 4'b1000 : node48610;
															assign node48610 = (inp[7]) ? 4'b1010 : node48611;
																assign node48611 = (inp[14]) ? 4'b1010 : 4'b1011;
													assign node48616 = (inp[0]) ? node48626 : node48617;
														assign node48617 = (inp[15]) ? node48619 : 4'b1001;
															assign node48619 = (inp[7]) ? node48623 : node48620;
																assign node48620 = (inp[14]) ? 4'b1010 : 4'b1011;
																assign node48623 = (inp[14]) ? 4'b1011 : 4'b1010;
														assign node48626 = (inp[15]) ? 4'b1001 : node48627;
															assign node48627 = (inp[14]) ? 4'b1010 : 4'b1011;
												assign node48631 = (inp[15]) ? node48647 : node48632;
													assign node48632 = (inp[0]) ? node48642 : node48633;
														assign node48633 = (inp[12]) ? node48635 : 4'b1001;
															assign node48635 = (inp[14]) ? node48639 : node48636;
																assign node48636 = (inp[7]) ? 4'b1001 : 4'b1000;
																assign node48639 = (inp[7]) ? 4'b1000 : 4'b1001;
														assign node48642 = (inp[7]) ? node48644 : 4'b1010;
															assign node48644 = (inp[14]) ? 4'b1010 : 4'b1011;
													assign node48647 = (inp[0]) ? node48651 : node48648;
														assign node48648 = (inp[14]) ? 4'b1011 : 4'b1010;
														assign node48651 = (inp[7]) ? node48655 : node48652;
															assign node48652 = (inp[14]) ? 4'b1001 : 4'b1000;
															assign node48655 = (inp[14]) ? 4'b1000 : 4'b1001;
								assign node48658 = (inp[0]) ? node48866 : node48659;
									assign node48659 = (inp[15]) ? node48765 : node48660;
										assign node48660 = (inp[5]) ? node48706 : node48661;
											assign node48661 = (inp[7]) ? node48683 : node48662;
												assign node48662 = (inp[8]) ? node48670 : node48663;
													assign node48663 = (inp[9]) ? node48667 : node48664;
														assign node48664 = (inp[4]) ? 4'b1110 : 4'b1010;
														assign node48667 = (inp[4]) ? 4'b1010 : 4'b1110;
													assign node48670 = (inp[14]) ? node48676 : node48671;
														assign node48671 = (inp[4]) ? 4'b1111 : node48672;
															assign node48672 = (inp[9]) ? 4'b1111 : 4'b1011;
														assign node48676 = (inp[9]) ? node48680 : node48677;
															assign node48677 = (inp[4]) ? 4'b1111 : 4'b1011;
															assign node48680 = (inp[4]) ? 4'b1011 : 4'b1111;
												assign node48683 = (inp[8]) ? node48699 : node48684;
													assign node48684 = (inp[12]) ? node48692 : node48685;
														assign node48685 = (inp[9]) ? node48689 : node48686;
															assign node48686 = (inp[4]) ? 4'b1111 : 4'b1011;
															assign node48689 = (inp[4]) ? 4'b1011 : 4'b1111;
														assign node48692 = (inp[9]) ? node48696 : node48693;
															assign node48693 = (inp[4]) ? 4'b1111 : 4'b1011;
															assign node48696 = (inp[4]) ? 4'b1011 : 4'b1111;
													assign node48699 = (inp[9]) ? node48703 : node48700;
														assign node48700 = (inp[4]) ? 4'b1110 : 4'b1010;
														assign node48703 = (inp[4]) ? 4'b1010 : 4'b1110;
											assign node48706 = (inp[4]) ? node48736 : node48707;
												assign node48707 = (inp[9]) ? node48729 : node48708;
													assign node48708 = (inp[12]) ? node48716 : node48709;
														assign node48709 = (inp[14]) ? node48711 : 4'b1011;
															assign node48711 = (inp[8]) ? node48713 : 4'b1011;
																assign node48713 = (inp[7]) ? 4'b1010 : 4'b1011;
														assign node48716 = (inp[14]) ? node48722 : node48717;
															assign node48717 = (inp[7]) ? node48719 : 4'b1010;
																assign node48719 = (inp[8]) ? 4'b1010 : 4'b1011;
															assign node48722 = (inp[8]) ? node48726 : node48723;
																assign node48723 = (inp[7]) ? 4'b1011 : 4'b1010;
																assign node48726 = (inp[7]) ? 4'b1010 : 4'b1011;
													assign node48729 = (inp[7]) ? node48733 : node48730;
														assign node48730 = (inp[8]) ? 4'b1101 : 4'b1100;
														assign node48733 = (inp[8]) ? 4'b1100 : 4'b1101;
												assign node48736 = (inp[9]) ? node48752 : node48737;
													assign node48737 = (inp[14]) ? node48745 : node48738;
														assign node48738 = (inp[8]) ? node48742 : node48739;
															assign node48739 = (inp[7]) ? 4'b1101 : 4'b1100;
															assign node48742 = (inp[7]) ? 4'b1100 : 4'b1101;
														assign node48745 = (inp[7]) ? node48749 : node48746;
															assign node48746 = (inp[8]) ? 4'b1101 : 4'b1100;
															assign node48749 = (inp[8]) ? 4'b1100 : 4'b1101;
													assign node48752 = (inp[14]) ? node48758 : node48753;
														assign node48753 = (inp[8]) ? 4'b1001 : node48754;
															assign node48754 = (inp[7]) ? 4'b1001 : 4'b1000;
														assign node48758 = (inp[8]) ? node48762 : node48759;
															assign node48759 = (inp[7]) ? 4'b1001 : 4'b1000;
															assign node48762 = (inp[7]) ? 4'b1000 : 4'b1001;
										assign node48765 = (inp[5]) ? node48811 : node48766;
											assign node48766 = (inp[8]) ? node48790 : node48767;
												assign node48767 = (inp[7]) ? node48783 : node48768;
													assign node48768 = (inp[12]) ? node48776 : node48769;
														assign node48769 = (inp[4]) ? node48773 : node48770;
															assign node48770 = (inp[9]) ? 4'b1100 : 4'b1000;
															assign node48773 = (inp[9]) ? 4'b1000 : 4'b1100;
														assign node48776 = (inp[4]) ? node48780 : node48777;
															assign node48777 = (inp[9]) ? 4'b1100 : 4'b1000;
															assign node48780 = (inp[9]) ? 4'b1000 : 4'b1100;
													assign node48783 = (inp[4]) ? node48787 : node48784;
														assign node48784 = (inp[9]) ? 4'b1101 : 4'b1001;
														assign node48787 = (inp[9]) ? 4'b1001 : 4'b1101;
												assign node48790 = (inp[7]) ? node48798 : node48791;
													assign node48791 = (inp[9]) ? node48795 : node48792;
														assign node48792 = (inp[4]) ? 4'b1101 : 4'b1001;
														assign node48795 = (inp[4]) ? 4'b1001 : 4'b1101;
													assign node48798 = (inp[12]) ? node48804 : node48799;
														assign node48799 = (inp[4]) ? node48801 : 4'b1100;
															assign node48801 = (inp[9]) ? 4'b1000 : 4'b1100;
														assign node48804 = (inp[9]) ? node48808 : node48805;
															assign node48805 = (inp[4]) ? 4'b1100 : 4'b1000;
															assign node48808 = (inp[4]) ? 4'b1000 : 4'b1100;
											assign node48811 = (inp[9]) ? node48835 : node48812;
												assign node48812 = (inp[4]) ? node48820 : node48813;
													assign node48813 = (inp[8]) ? node48817 : node48814;
														assign node48814 = (inp[7]) ? 4'b1001 : 4'b1000;
														assign node48817 = (inp[7]) ? 4'b1000 : 4'b1001;
													assign node48820 = (inp[12]) ? node48828 : node48821;
														assign node48821 = (inp[8]) ? node48825 : node48822;
															assign node48822 = (inp[7]) ? 4'b1111 : 4'b1110;
															assign node48825 = (inp[7]) ? 4'b1110 : 4'b1111;
														assign node48828 = (inp[8]) ? node48832 : node48829;
															assign node48829 = (inp[7]) ? 4'b1111 : 4'b1110;
															assign node48832 = (inp[7]) ? 4'b1110 : 4'b1111;
												assign node48835 = (inp[4]) ? node48851 : node48836;
													assign node48836 = (inp[12]) ? node48844 : node48837;
														assign node48837 = (inp[7]) ? node48841 : node48838;
															assign node48838 = (inp[8]) ? 4'b1111 : 4'b1110;
															assign node48841 = (inp[8]) ? 4'b1110 : 4'b1111;
														assign node48844 = (inp[8]) ? node48848 : node48845;
															assign node48845 = (inp[7]) ? 4'b1111 : 4'b1110;
															assign node48848 = (inp[7]) ? 4'b1110 : 4'b1111;
													assign node48851 = (inp[12]) ? node48859 : node48852;
														assign node48852 = (inp[8]) ? node48856 : node48853;
															assign node48853 = (inp[7]) ? 4'b1011 : 4'b1010;
															assign node48856 = (inp[7]) ? 4'b1010 : 4'b1011;
														assign node48859 = (inp[14]) ? 4'b1011 : node48860;
															assign node48860 = (inp[7]) ? 4'b1011 : node48861;
																assign node48861 = (inp[8]) ? 4'b1011 : 4'b1010;
									assign node48866 = (inp[15]) ? node48970 : node48867;
										assign node48867 = (inp[5]) ? node48909 : node48868;
											assign node48868 = (inp[8]) ? node48886 : node48869;
												assign node48869 = (inp[7]) ? node48879 : node48870;
													assign node48870 = (inp[14]) ? node48872 : 4'b1000;
														assign node48872 = (inp[4]) ? node48876 : node48873;
															assign node48873 = (inp[9]) ? 4'b1100 : 4'b1000;
															assign node48876 = (inp[9]) ? 4'b1000 : 4'b1100;
													assign node48879 = (inp[4]) ? node48883 : node48880;
														assign node48880 = (inp[9]) ? 4'b1101 : 4'b1001;
														assign node48883 = (inp[9]) ? 4'b1001 : 4'b1101;
												assign node48886 = (inp[7]) ? node48902 : node48887;
													assign node48887 = (inp[14]) ? node48895 : node48888;
														assign node48888 = (inp[12]) ? 4'b1101 : node48889;
															assign node48889 = (inp[4]) ? node48891 : 4'b1101;
																assign node48891 = (inp[9]) ? 4'b1001 : 4'b1101;
														assign node48895 = (inp[4]) ? node48899 : node48896;
															assign node48896 = (inp[9]) ? 4'b1101 : 4'b1001;
															assign node48899 = (inp[9]) ? 4'b1001 : 4'b1101;
													assign node48902 = (inp[9]) ? node48906 : node48903;
														assign node48903 = (inp[4]) ? 4'b1100 : 4'b1000;
														assign node48906 = (inp[4]) ? 4'b1000 : 4'b1100;
											assign node48909 = (inp[4]) ? node48931 : node48910;
												assign node48910 = (inp[9]) ? node48918 : node48911;
													assign node48911 = (inp[7]) ? node48915 : node48912;
														assign node48912 = (inp[8]) ? 4'b1001 : 4'b1000;
														assign node48915 = (inp[8]) ? 4'b1000 : 4'b1001;
													assign node48918 = (inp[12]) ? node48926 : node48919;
														assign node48919 = (inp[8]) ? node48923 : node48920;
															assign node48920 = (inp[7]) ? 4'b1111 : 4'b1110;
															assign node48923 = (inp[7]) ? 4'b1110 : 4'b1111;
														assign node48926 = (inp[7]) ? 4'b1111 : node48927;
															assign node48927 = (inp[8]) ? 4'b1111 : 4'b1110;
												assign node48931 = (inp[9]) ? node48951 : node48932;
													assign node48932 = (inp[12]) ? node48942 : node48933;
														assign node48933 = (inp[14]) ? 4'b1111 : node48934;
															assign node48934 = (inp[7]) ? node48938 : node48935;
																assign node48935 = (inp[8]) ? 4'b1111 : 4'b1110;
																assign node48938 = (inp[8]) ? 4'b1110 : 4'b1111;
														assign node48942 = (inp[14]) ? node48944 : 4'b1111;
															assign node48944 = (inp[7]) ? node48948 : node48945;
																assign node48945 = (inp[8]) ? 4'b1111 : 4'b1110;
																assign node48948 = (inp[8]) ? 4'b1110 : 4'b1111;
													assign node48951 = (inp[12]) ? node48957 : node48952;
														assign node48952 = (inp[8]) ? 4'b1010 : node48953;
															assign node48953 = (inp[7]) ? 4'b1011 : 4'b1010;
														assign node48957 = (inp[14]) ? node48965 : node48958;
															assign node48958 = (inp[7]) ? node48962 : node48959;
																assign node48959 = (inp[8]) ? 4'b1011 : 4'b1010;
																assign node48962 = (inp[8]) ? 4'b1010 : 4'b1011;
															assign node48965 = (inp[8]) ? node48967 : 4'b1011;
																assign node48967 = (inp[7]) ? 4'b1010 : 4'b1011;
										assign node48970 = (inp[5]) ? node49012 : node48971;
											assign node48971 = (inp[8]) ? node48993 : node48972;
												assign node48972 = (inp[7]) ? node48986 : node48973;
													assign node48973 = (inp[14]) ? node48981 : node48974;
														assign node48974 = (inp[4]) ? node48978 : node48975;
															assign node48975 = (inp[9]) ? 4'b1110 : 4'b1010;
															assign node48978 = (inp[9]) ? 4'b1010 : 4'b1110;
														assign node48981 = (inp[9]) ? 4'b1110 : node48982;
															assign node48982 = (inp[4]) ? 4'b1110 : 4'b1010;
													assign node48986 = (inp[9]) ? node48990 : node48987;
														assign node48987 = (inp[4]) ? 4'b1111 : 4'b1011;
														assign node48990 = (inp[4]) ? 4'b1011 : 4'b1111;
												assign node48993 = (inp[7]) ? node49001 : node48994;
													assign node48994 = (inp[4]) ? node48998 : node48995;
														assign node48995 = (inp[9]) ? 4'b1111 : 4'b1011;
														assign node48998 = (inp[9]) ? 4'b1011 : 4'b1111;
													assign node49001 = (inp[14]) ? node49007 : node49002;
														assign node49002 = (inp[4]) ? 4'b1110 : node49003;
															assign node49003 = (inp[9]) ? 4'b1110 : 4'b1010;
														assign node49007 = (inp[4]) ? 4'b1010 : node49008;
															assign node49008 = (inp[12]) ? 4'b1010 : 4'b1110;
											assign node49012 = (inp[4]) ? node49034 : node49013;
												assign node49013 = (inp[9]) ? node49021 : node49014;
													assign node49014 = (inp[7]) ? node49018 : node49015;
														assign node49015 = (inp[8]) ? 4'b1011 : 4'b1010;
														assign node49018 = (inp[8]) ? 4'b1010 : 4'b1011;
													assign node49021 = (inp[14]) ? node49027 : node49022;
														assign node49022 = (inp[8]) ? node49024 : 4'b1101;
															assign node49024 = (inp[7]) ? 4'b1100 : 4'b1101;
														assign node49027 = (inp[8]) ? node49031 : node49028;
															assign node49028 = (inp[7]) ? 4'b1101 : 4'b1100;
															assign node49031 = (inp[7]) ? 4'b1100 : 4'b1101;
												assign node49034 = (inp[9]) ? node49042 : node49035;
													assign node49035 = (inp[8]) ? node49039 : node49036;
														assign node49036 = (inp[7]) ? 4'b1101 : 4'b1100;
														assign node49039 = (inp[7]) ? 4'b1100 : 4'b1101;
													assign node49042 = (inp[14]) ? node49050 : node49043;
														assign node49043 = (inp[7]) ? node49047 : node49044;
															assign node49044 = (inp[8]) ? 4'b1001 : 4'b1000;
															assign node49047 = (inp[8]) ? 4'b1000 : 4'b1001;
														assign node49050 = (inp[12]) ? node49052 : 4'b1001;
															assign node49052 = (inp[8]) ? node49056 : node49053;
																assign node49053 = (inp[7]) ? 4'b1001 : 4'b1000;
																assign node49056 = (inp[7]) ? 4'b1000 : 4'b1001;
							assign node49059 = (inp[8]) ? node49511 : node49060;
								assign node49060 = (inp[7]) ? node49292 : node49061;
									assign node49061 = (inp[2]) ? node49177 : node49062;
										assign node49062 = (inp[14]) ? node49130 : node49063;
											assign node49063 = (inp[12]) ? node49091 : node49064;
												assign node49064 = (inp[4]) ? node49078 : node49065;
													assign node49065 = (inp[9]) ? node49071 : node49066;
														assign node49066 = (inp[0]) ? 4'b1011 : node49067;
															assign node49067 = (inp[15]) ? 4'b1011 : 4'b1001;
														assign node49071 = (inp[0]) ? node49075 : node49072;
															assign node49072 = (inp[15]) ? 4'b1111 : 4'b1101;
															assign node49075 = (inp[15]) ? 4'b1101 : 4'b1111;
													assign node49078 = (inp[9]) ? node49086 : node49079;
														assign node49079 = (inp[0]) ? node49083 : node49080;
															assign node49080 = (inp[15]) ? 4'b1111 : 4'b1101;
															assign node49083 = (inp[15]) ? 4'b1101 : 4'b1111;
														assign node49086 = (inp[15]) ? node49088 : 4'b1001;
															assign node49088 = (inp[5]) ? 4'b1011 : 4'b1001;
												assign node49091 = (inp[15]) ? node49111 : node49092;
													assign node49092 = (inp[0]) ? node49102 : node49093;
														assign node49093 = (inp[9]) ? node49099 : node49094;
															assign node49094 = (inp[4]) ? 4'b1101 : node49095;
																assign node49095 = (inp[5]) ? 4'b1001 : 4'b1011;
															assign node49099 = (inp[4]) ? 4'b1001 : 4'b1101;
														assign node49102 = (inp[4]) ? node49108 : node49103;
															assign node49103 = (inp[9]) ? 4'b1111 : node49104;
																assign node49104 = (inp[5]) ? 4'b1011 : 4'b1001;
															assign node49108 = (inp[9]) ? 4'b1011 : 4'b1111;
													assign node49111 = (inp[0]) ? node49121 : node49112;
														assign node49112 = (inp[4]) ? node49118 : node49113;
															assign node49113 = (inp[9]) ? 4'b1111 : node49114;
																assign node49114 = (inp[5]) ? 4'b1011 : 4'b1001;
															assign node49118 = (inp[9]) ? 4'b1011 : 4'b1111;
														assign node49121 = (inp[5]) ? node49125 : node49122;
															assign node49122 = (inp[9]) ? 4'b1001 : 4'b1101;
															assign node49125 = (inp[4]) ? 4'b1001 : node49126;
																assign node49126 = (inp[9]) ? 4'b1101 : 4'b1001;
											assign node49130 = (inp[9]) ? node49154 : node49131;
												assign node49131 = (inp[4]) ? node49147 : node49132;
													assign node49132 = (inp[15]) ? 4'b1000 : node49133;
														assign node49133 = (inp[12]) ? node49139 : node49134;
															assign node49134 = (inp[5]) ? node49136 : 4'b1000;
																assign node49136 = (inp[0]) ? 4'b1010 : 4'b1000;
															assign node49139 = (inp[5]) ? node49143 : node49140;
																assign node49140 = (inp[0]) ? 4'b1000 : 4'b1010;
																assign node49143 = (inp[0]) ? 4'b1010 : 4'b1000;
													assign node49147 = (inp[0]) ? node49151 : node49148;
														assign node49148 = (inp[15]) ? 4'b1110 : 4'b1100;
														assign node49151 = (inp[15]) ? 4'b1100 : 4'b1110;
												assign node49154 = (inp[4]) ? node49162 : node49155;
													assign node49155 = (inp[0]) ? node49159 : node49156;
														assign node49156 = (inp[15]) ? 4'b1110 : 4'b1100;
														assign node49159 = (inp[15]) ? 4'b1100 : 4'b1110;
													assign node49162 = (inp[5]) ? node49170 : node49163;
														assign node49163 = (inp[0]) ? node49167 : node49164;
															assign node49164 = (inp[15]) ? 4'b1010 : 4'b1000;
															assign node49167 = (inp[15]) ? 4'b1000 : 4'b1010;
														assign node49170 = (inp[0]) ? node49174 : node49171;
															assign node49171 = (inp[15]) ? 4'b1010 : 4'b1000;
															assign node49174 = (inp[15]) ? 4'b1000 : 4'b1010;
										assign node49177 = (inp[5]) ? node49237 : node49178;
											assign node49178 = (inp[14]) ? node49208 : node49179;
												assign node49179 = (inp[0]) ? node49195 : node49180;
													assign node49180 = (inp[15]) ? node49188 : node49181;
														assign node49181 = (inp[9]) ? node49185 : node49182;
															assign node49182 = (inp[4]) ? 4'b1100 : 4'b1010;
															assign node49185 = (inp[4]) ? 4'b1000 : 4'b1100;
														assign node49188 = (inp[4]) ? node49192 : node49189;
															assign node49189 = (inp[9]) ? 4'b1110 : 4'b1000;
															assign node49192 = (inp[9]) ? 4'b1010 : 4'b1110;
													assign node49195 = (inp[15]) ? node49201 : node49196;
														assign node49196 = (inp[9]) ? node49198 : 4'b1110;
															assign node49198 = (inp[4]) ? 4'b1010 : 4'b1110;
														assign node49201 = (inp[4]) ? node49205 : node49202;
															assign node49202 = (inp[9]) ? 4'b1100 : 4'b1010;
															assign node49205 = (inp[9]) ? 4'b1000 : 4'b1100;
												assign node49208 = (inp[0]) ? node49222 : node49209;
													assign node49209 = (inp[15]) ? node49215 : node49210;
														assign node49210 = (inp[4]) ? node49212 : 4'b1010;
															assign node49212 = (inp[9]) ? 4'b1000 : 4'b1100;
														assign node49215 = (inp[9]) ? node49219 : node49216;
															assign node49216 = (inp[4]) ? 4'b1110 : 4'b1000;
															assign node49219 = (inp[4]) ? 4'b1010 : 4'b1110;
													assign node49222 = (inp[15]) ? node49230 : node49223;
														assign node49223 = (inp[4]) ? node49227 : node49224;
															assign node49224 = (inp[9]) ? 4'b1110 : 4'b1000;
															assign node49227 = (inp[9]) ? 4'b1010 : 4'b1110;
														assign node49230 = (inp[4]) ? node49234 : node49231;
															assign node49231 = (inp[9]) ? 4'b1100 : 4'b1010;
															assign node49234 = (inp[9]) ? 4'b1000 : 4'b1100;
											assign node49237 = (inp[4]) ? node49277 : node49238;
												assign node49238 = (inp[9]) ? node49258 : node49239;
													assign node49239 = (inp[14]) ? node49251 : node49240;
														assign node49240 = (inp[12]) ? node49246 : node49241;
															assign node49241 = (inp[15]) ? 4'b1010 : node49242;
																assign node49242 = (inp[0]) ? 4'b1010 : 4'b1000;
															assign node49246 = (inp[15]) ? 4'b1000 : node49247;
																assign node49247 = (inp[0]) ? 4'b1010 : 4'b1000;
														assign node49251 = (inp[0]) ? node49255 : node49252;
															assign node49252 = (inp[15]) ? 4'b1010 : 4'b1000;
															assign node49255 = (inp[15]) ? 4'b1000 : 4'b1010;
													assign node49258 = (inp[12]) ? node49270 : node49259;
														assign node49259 = (inp[14]) ? node49265 : node49260;
															assign node49260 = (inp[0]) ? 4'b1100 : node49261;
																assign node49261 = (inp[15]) ? 4'b1110 : 4'b1100;
															assign node49265 = (inp[15]) ? 4'b1100 : node49266;
																assign node49266 = (inp[0]) ? 4'b1110 : 4'b1100;
														assign node49270 = (inp[0]) ? node49274 : node49271;
															assign node49271 = (inp[15]) ? 4'b1110 : 4'b1100;
															assign node49274 = (inp[15]) ? 4'b1100 : 4'b1110;
												assign node49277 = (inp[9]) ? node49285 : node49278;
													assign node49278 = (inp[0]) ? node49282 : node49279;
														assign node49279 = (inp[15]) ? 4'b1110 : 4'b1100;
														assign node49282 = (inp[15]) ? 4'b1100 : 4'b1110;
													assign node49285 = (inp[0]) ? node49289 : node49286;
														assign node49286 = (inp[15]) ? 4'b1010 : 4'b1000;
														assign node49289 = (inp[15]) ? 4'b1000 : 4'b1010;
									assign node49292 = (inp[2]) ? node49404 : node49293;
										assign node49293 = (inp[14]) ? node49351 : node49294;
											assign node49294 = (inp[0]) ? node49314 : node49295;
												assign node49295 = (inp[15]) ? node49305 : node49296;
													assign node49296 = (inp[4]) ? node49302 : node49297;
														assign node49297 = (inp[9]) ? 4'b1100 : node49298;
															assign node49298 = (inp[5]) ? 4'b1000 : 4'b1010;
														assign node49302 = (inp[9]) ? 4'b1000 : 4'b1100;
													assign node49305 = (inp[4]) ? node49311 : node49306;
														assign node49306 = (inp[9]) ? 4'b1110 : node49307;
															assign node49307 = (inp[5]) ? 4'b1010 : 4'b1000;
														assign node49311 = (inp[9]) ? 4'b1010 : 4'b1110;
												assign node49314 = (inp[15]) ? node49330 : node49315;
													assign node49315 = (inp[5]) ? node49323 : node49316;
														assign node49316 = (inp[9]) ? node49320 : node49317;
															assign node49317 = (inp[12]) ? 4'b1110 : 4'b1000;
															assign node49320 = (inp[4]) ? 4'b1010 : 4'b1110;
														assign node49323 = (inp[9]) ? node49327 : node49324;
															assign node49324 = (inp[4]) ? 4'b1110 : 4'b1010;
															assign node49327 = (inp[4]) ? 4'b1010 : 4'b1110;
													assign node49330 = (inp[12]) ? node49342 : node49331;
														assign node49331 = (inp[5]) ? node49337 : node49332;
															assign node49332 = (inp[9]) ? node49334 : 4'b1100;
																assign node49334 = (inp[4]) ? 4'b1000 : 4'b1100;
															assign node49337 = (inp[4]) ? 4'b1100 : node49338;
																assign node49338 = (inp[9]) ? 4'b1100 : 4'b1000;
														assign node49342 = (inp[9]) ? node49348 : node49343;
															assign node49343 = (inp[4]) ? 4'b1100 : node49344;
																assign node49344 = (inp[5]) ? 4'b1000 : 4'b1010;
															assign node49348 = (inp[4]) ? 4'b1000 : 4'b1100;
											assign node49351 = (inp[15]) ? node49381 : node49352;
												assign node49352 = (inp[0]) ? node49366 : node49353;
													assign node49353 = (inp[5]) ? node49359 : node49354;
														assign node49354 = (inp[4]) ? node49356 : 4'b1011;
															assign node49356 = (inp[9]) ? 4'b1001 : 4'b1101;
														assign node49359 = (inp[4]) ? node49363 : node49360;
															assign node49360 = (inp[9]) ? 4'b1101 : 4'b1001;
															assign node49363 = (inp[9]) ? 4'b1001 : 4'b1101;
													assign node49366 = (inp[5]) ? node49374 : node49367;
														assign node49367 = (inp[9]) ? node49371 : node49368;
															assign node49368 = (inp[4]) ? 4'b1111 : 4'b1001;
															assign node49371 = (inp[4]) ? 4'b1011 : 4'b1111;
														assign node49374 = (inp[9]) ? node49378 : node49375;
															assign node49375 = (inp[4]) ? 4'b1111 : 4'b1011;
															assign node49378 = (inp[4]) ? 4'b1011 : 4'b1111;
												assign node49381 = (inp[0]) ? node49391 : node49382;
													assign node49382 = (inp[9]) ? node49388 : node49383;
														assign node49383 = (inp[4]) ? 4'b1111 : node49384;
															assign node49384 = (inp[5]) ? 4'b1011 : 4'b1001;
														assign node49388 = (inp[4]) ? 4'b1011 : 4'b1111;
													assign node49391 = (inp[12]) ? node49399 : node49392;
														assign node49392 = (inp[4]) ? 4'b1101 : node49393;
															assign node49393 = (inp[9]) ? 4'b1101 : node49394;
																assign node49394 = (inp[5]) ? 4'b1001 : 4'b1011;
														assign node49399 = (inp[5]) ? 4'b1001 : node49400;
															assign node49400 = (inp[4]) ? 4'b1001 : 4'b1101;
										assign node49404 = (inp[12]) ? node49454 : node49405;
											assign node49405 = (inp[15]) ? node49427 : node49406;
												assign node49406 = (inp[0]) ? node49418 : node49407;
													assign node49407 = (inp[14]) ? 4'b1001 : node49408;
														assign node49408 = (inp[4]) ? node49414 : node49409;
															assign node49409 = (inp[9]) ? 4'b1101 : node49410;
																assign node49410 = (inp[5]) ? 4'b1001 : 4'b1011;
															assign node49414 = (inp[9]) ? 4'b1001 : 4'b1101;
													assign node49418 = (inp[4]) ? node49424 : node49419;
														assign node49419 = (inp[9]) ? 4'b1111 : node49420;
															assign node49420 = (inp[5]) ? 4'b1011 : 4'b1001;
														assign node49424 = (inp[9]) ? 4'b1011 : 4'b1111;
												assign node49427 = (inp[0]) ? node49445 : node49428;
													assign node49428 = (inp[5]) ? node49438 : node49429;
														assign node49429 = (inp[14]) ? 4'b1111 : node49430;
															assign node49430 = (inp[4]) ? node49434 : node49431;
																assign node49431 = (inp[9]) ? 4'b1111 : 4'b1001;
																assign node49434 = (inp[9]) ? 4'b1011 : 4'b1111;
														assign node49438 = (inp[9]) ? node49442 : node49439;
															assign node49439 = (inp[4]) ? 4'b1111 : 4'b1011;
															assign node49442 = (inp[4]) ? 4'b1011 : 4'b1111;
													assign node49445 = (inp[9]) ? node49451 : node49446;
														assign node49446 = (inp[4]) ? 4'b1101 : node49447;
															assign node49447 = (inp[5]) ? 4'b1001 : 4'b1011;
														assign node49451 = (inp[4]) ? 4'b1001 : 4'b1101;
											assign node49454 = (inp[5]) ? node49486 : node49455;
												assign node49455 = (inp[15]) ? node49471 : node49456;
													assign node49456 = (inp[0]) ? node49464 : node49457;
														assign node49457 = (inp[9]) ? node49461 : node49458;
															assign node49458 = (inp[4]) ? 4'b1101 : 4'b1011;
															assign node49461 = (inp[4]) ? 4'b1001 : 4'b1101;
														assign node49464 = (inp[9]) ? node49468 : node49465;
															assign node49465 = (inp[4]) ? 4'b1111 : 4'b1001;
															assign node49468 = (inp[4]) ? 4'b1011 : 4'b1111;
													assign node49471 = (inp[0]) ? node49479 : node49472;
														assign node49472 = (inp[9]) ? node49476 : node49473;
															assign node49473 = (inp[4]) ? 4'b1111 : 4'b1001;
															assign node49476 = (inp[4]) ? 4'b1011 : 4'b1111;
														assign node49479 = (inp[9]) ? node49483 : node49480;
															assign node49480 = (inp[4]) ? 4'b1101 : 4'b1011;
															assign node49483 = (inp[4]) ? 4'b1001 : 4'b1101;
												assign node49486 = (inp[0]) ? node49500 : node49487;
													assign node49487 = (inp[15]) ? node49495 : node49488;
														assign node49488 = (inp[4]) ? node49492 : node49489;
															assign node49489 = (inp[9]) ? 4'b1101 : 4'b1001;
															assign node49492 = (inp[9]) ? 4'b1001 : 4'b1101;
														assign node49495 = (inp[4]) ? node49497 : 4'b1111;
															assign node49497 = (inp[9]) ? 4'b1011 : 4'b1111;
													assign node49500 = (inp[15]) ? node49506 : node49501;
														assign node49501 = (inp[4]) ? 4'b1111 : node49502;
															assign node49502 = (inp[14]) ? 4'b1111 : 4'b1011;
														assign node49506 = (inp[4]) ? 4'b1101 : node49507;
															assign node49507 = (inp[9]) ? 4'b1101 : 4'b1001;
								assign node49511 = (inp[7]) ? node49643 : node49512;
									assign node49512 = (inp[14]) ? node49604 : node49513;
										assign node49513 = (inp[2]) ? node49557 : node49514;
											assign node49514 = (inp[0]) ? node49538 : node49515;
												assign node49515 = (inp[15]) ? node49531 : node49516;
													assign node49516 = (inp[12]) ? node49522 : node49517;
														assign node49517 = (inp[4]) ? 4'b1100 : node49518;
															assign node49518 = (inp[9]) ? 4'b1100 : 4'b1010;
														assign node49522 = (inp[5]) ? node49526 : node49523;
															assign node49523 = (inp[4]) ? 4'b1000 : 4'b1100;
															assign node49526 = (inp[9]) ? 4'b1100 : node49527;
																assign node49527 = (inp[4]) ? 4'b1100 : 4'b1000;
													assign node49531 = (inp[4]) ? node49535 : node49532;
														assign node49532 = (inp[9]) ? 4'b1110 : 4'b1000;
														assign node49535 = (inp[9]) ? 4'b1010 : 4'b1110;
												assign node49538 = (inp[15]) ? node49548 : node49539;
													assign node49539 = (inp[4]) ? node49545 : node49540;
														assign node49540 = (inp[9]) ? 4'b1110 : node49541;
															assign node49541 = (inp[5]) ? 4'b1010 : 4'b1000;
														assign node49545 = (inp[9]) ? 4'b1010 : 4'b1110;
													assign node49548 = (inp[4]) ? node49554 : node49549;
														assign node49549 = (inp[9]) ? 4'b1100 : node49550;
															assign node49550 = (inp[5]) ? 4'b1000 : 4'b1010;
														assign node49554 = (inp[9]) ? 4'b1000 : 4'b1100;
											assign node49557 = (inp[9]) ? node49583 : node49558;
												assign node49558 = (inp[4]) ? node49574 : node49559;
													assign node49559 = (inp[15]) ? node49567 : node49560;
														assign node49560 = (inp[0]) ? node49564 : node49561;
															assign node49561 = (inp[5]) ? 4'b1001 : 4'b1011;
															assign node49564 = (inp[5]) ? 4'b1011 : 4'b1001;
														assign node49567 = (inp[0]) ? node49571 : node49568;
															assign node49568 = (inp[5]) ? 4'b1011 : 4'b1001;
															assign node49571 = (inp[5]) ? 4'b1001 : 4'b1011;
													assign node49574 = (inp[5]) ? 4'b1101 : node49575;
														assign node49575 = (inp[15]) ? node49579 : node49576;
															assign node49576 = (inp[0]) ? 4'b1111 : 4'b1101;
															assign node49579 = (inp[0]) ? 4'b1101 : 4'b1111;
												assign node49583 = (inp[4]) ? node49591 : node49584;
													assign node49584 = (inp[15]) ? node49588 : node49585;
														assign node49585 = (inp[0]) ? 4'b1111 : 4'b1101;
														assign node49588 = (inp[0]) ? 4'b1101 : 4'b1111;
													assign node49591 = (inp[12]) ? node49597 : node49592;
														assign node49592 = (inp[15]) ? node49594 : 4'b1001;
															assign node49594 = (inp[0]) ? 4'b1001 : 4'b1011;
														assign node49597 = (inp[0]) ? node49601 : node49598;
															assign node49598 = (inp[15]) ? 4'b1011 : 4'b1001;
															assign node49601 = (inp[15]) ? 4'b1001 : 4'b1011;
										assign node49604 = (inp[15]) ? node49624 : node49605;
											assign node49605 = (inp[0]) ? node49615 : node49606;
												assign node49606 = (inp[9]) ? node49612 : node49607;
													assign node49607 = (inp[4]) ? 4'b1101 : node49608;
														assign node49608 = (inp[12]) ? 4'b1011 : 4'b1001;
													assign node49612 = (inp[4]) ? 4'b1001 : 4'b1101;
												assign node49615 = (inp[9]) ? node49621 : node49616;
													assign node49616 = (inp[4]) ? 4'b1111 : node49617;
														assign node49617 = (inp[5]) ? 4'b1011 : 4'b1001;
													assign node49621 = (inp[4]) ? 4'b1011 : 4'b1111;
											assign node49624 = (inp[0]) ? node49634 : node49625;
												assign node49625 = (inp[9]) ? node49631 : node49626;
													assign node49626 = (inp[4]) ? 4'b1111 : node49627;
														assign node49627 = (inp[5]) ? 4'b1011 : 4'b1001;
													assign node49631 = (inp[4]) ? 4'b1011 : 4'b1111;
												assign node49634 = (inp[4]) ? node49640 : node49635;
													assign node49635 = (inp[9]) ? 4'b1101 : node49636;
														assign node49636 = (inp[5]) ? 4'b1001 : 4'b1011;
													assign node49640 = (inp[9]) ? 4'b1001 : 4'b1101;
									assign node49643 = (inp[2]) ? node49777 : node49644;
										assign node49644 = (inp[14]) ? node49702 : node49645;
											assign node49645 = (inp[4]) ? node49679 : node49646;
												assign node49646 = (inp[9]) ? node49656 : node49647;
													assign node49647 = (inp[5]) ? node49649 : 4'b1001;
														assign node49649 = (inp[15]) ? node49653 : node49650;
															assign node49650 = (inp[0]) ? 4'b1011 : 4'b1001;
															assign node49653 = (inp[0]) ? 4'b1001 : 4'b1011;
													assign node49656 = (inp[5]) ? node49672 : node49657;
														assign node49657 = (inp[12]) ? node49665 : node49658;
															assign node49658 = (inp[0]) ? node49662 : node49659;
																assign node49659 = (inp[15]) ? 4'b1111 : 4'b1101;
																assign node49662 = (inp[15]) ? 4'b1101 : 4'b1111;
															assign node49665 = (inp[0]) ? node49669 : node49666;
																assign node49666 = (inp[15]) ? 4'b1111 : 4'b1101;
																assign node49669 = (inp[15]) ? 4'b1101 : 4'b1111;
														assign node49672 = (inp[0]) ? node49676 : node49673;
															assign node49673 = (inp[15]) ? 4'b1111 : 4'b1101;
															assign node49676 = (inp[15]) ? 4'b1101 : 4'b1111;
												assign node49679 = (inp[9]) ? node49687 : node49680;
													assign node49680 = (inp[0]) ? node49684 : node49681;
														assign node49681 = (inp[15]) ? 4'b1111 : 4'b1101;
														assign node49684 = (inp[15]) ? 4'b1101 : 4'b1111;
													assign node49687 = (inp[12]) ? node49695 : node49688;
														assign node49688 = (inp[0]) ? node49692 : node49689;
															assign node49689 = (inp[15]) ? 4'b1011 : 4'b1001;
															assign node49692 = (inp[15]) ? 4'b1001 : 4'b1011;
														assign node49695 = (inp[0]) ? node49699 : node49696;
															assign node49696 = (inp[15]) ? 4'b1011 : 4'b1001;
															assign node49699 = (inp[15]) ? 4'b1001 : 4'b1011;
											assign node49702 = (inp[4]) ? node49744 : node49703;
												assign node49703 = (inp[9]) ? node49721 : node49704;
													assign node49704 = (inp[5]) ? node49716 : node49705;
														assign node49705 = (inp[12]) ? node49711 : node49706;
															assign node49706 = (inp[15]) ? node49708 : 4'b1010;
																assign node49708 = (inp[0]) ? 4'b1010 : 4'b1000;
															assign node49711 = (inp[15]) ? 4'b1010 : node49712;
																assign node49712 = (inp[0]) ? 4'b1000 : 4'b1010;
														assign node49716 = (inp[15]) ? 4'b1000 : node49717;
															assign node49717 = (inp[0]) ? 4'b1010 : 4'b1000;
													assign node49721 = (inp[12]) ? node49731 : node49722;
														assign node49722 = (inp[5]) ? 4'b1100 : node49723;
															assign node49723 = (inp[15]) ? node49727 : node49724;
																assign node49724 = (inp[0]) ? 4'b1110 : 4'b1100;
																assign node49727 = (inp[0]) ? 4'b1100 : 4'b1110;
														assign node49731 = (inp[5]) ? node49737 : node49732;
															assign node49732 = (inp[0]) ? 4'b1100 : node49733;
																assign node49733 = (inp[15]) ? 4'b1110 : 4'b1100;
															assign node49737 = (inp[15]) ? node49741 : node49738;
																assign node49738 = (inp[0]) ? 4'b1110 : 4'b1100;
																assign node49741 = (inp[0]) ? 4'b1100 : 4'b1110;
												assign node49744 = (inp[9]) ? node49760 : node49745;
													assign node49745 = (inp[12]) ? node49755 : node49746;
														assign node49746 = (inp[5]) ? node49748 : 4'b1110;
															assign node49748 = (inp[15]) ? node49752 : node49749;
																assign node49749 = (inp[0]) ? 4'b1110 : 4'b1100;
																assign node49752 = (inp[0]) ? 4'b1100 : 4'b1110;
														assign node49755 = (inp[15]) ? 4'b1100 : node49756;
															assign node49756 = (inp[0]) ? 4'b1110 : 4'b1100;
													assign node49760 = (inp[5]) ? node49772 : node49761;
														assign node49761 = (inp[12]) ? node49767 : node49762;
															assign node49762 = (inp[0]) ? node49764 : 4'b1000;
																assign node49764 = (inp[15]) ? 4'b1000 : 4'b1010;
															assign node49767 = (inp[15]) ? node49769 : 4'b1000;
																assign node49769 = (inp[0]) ? 4'b1000 : 4'b1010;
														assign node49772 = (inp[15]) ? 4'b1010 : node49773;
															assign node49773 = (inp[0]) ? 4'b1010 : 4'b1000;
										assign node49777 = (inp[9]) ? node49829 : node49778;
											assign node49778 = (inp[4]) ? node49822 : node49779;
												assign node49779 = (inp[5]) ? node49807 : node49780;
													assign node49780 = (inp[12]) ? node49792 : node49781;
														assign node49781 = (inp[14]) ? node49787 : node49782;
															assign node49782 = (inp[15]) ? node49784 : 4'b1000;
																assign node49784 = (inp[0]) ? 4'b1010 : 4'b1000;
															assign node49787 = (inp[15]) ? 4'b1000 : node49788;
																assign node49788 = (inp[0]) ? 4'b1000 : 4'b1010;
														assign node49792 = (inp[14]) ? node49800 : node49793;
															assign node49793 = (inp[0]) ? node49797 : node49794;
																assign node49794 = (inp[15]) ? 4'b1000 : 4'b1010;
																assign node49797 = (inp[15]) ? 4'b1010 : 4'b1000;
															assign node49800 = (inp[15]) ? node49804 : node49801;
																assign node49801 = (inp[0]) ? 4'b1000 : 4'b1010;
																assign node49804 = (inp[0]) ? 4'b1010 : 4'b1000;
													assign node49807 = (inp[14]) ? node49815 : node49808;
														assign node49808 = (inp[15]) ? node49812 : node49809;
															assign node49809 = (inp[0]) ? 4'b1010 : 4'b1000;
															assign node49812 = (inp[0]) ? 4'b1000 : 4'b1010;
														assign node49815 = (inp[0]) ? node49819 : node49816;
															assign node49816 = (inp[15]) ? 4'b1010 : 4'b1000;
															assign node49819 = (inp[15]) ? 4'b1000 : 4'b1010;
												assign node49822 = (inp[15]) ? node49826 : node49823;
													assign node49823 = (inp[0]) ? 4'b1110 : 4'b1100;
													assign node49826 = (inp[0]) ? 4'b1100 : 4'b1110;
											assign node49829 = (inp[4]) ? node49845 : node49830;
												assign node49830 = (inp[5]) ? node49838 : node49831;
													assign node49831 = (inp[15]) ? node49835 : node49832;
														assign node49832 = (inp[0]) ? 4'b1110 : 4'b1100;
														assign node49835 = (inp[0]) ? 4'b1100 : 4'b1110;
													assign node49838 = (inp[15]) ? node49842 : node49839;
														assign node49839 = (inp[0]) ? 4'b1110 : 4'b1100;
														assign node49842 = (inp[0]) ? 4'b1100 : 4'b1110;
												assign node49845 = (inp[0]) ? node49849 : node49846;
													assign node49846 = (inp[15]) ? 4'b1010 : 4'b1000;
													assign node49849 = (inp[15]) ? 4'b1000 : 4'b1010;
			assign node49852 = (inp[1]) ? node58052 : node49853;
				assign node49853 = (inp[13]) ? node54113 : node49854;
					assign node49854 = (inp[5]) ? node52070 : node49855;
						assign node49855 = (inp[12]) ? node51149 : node49856;
							assign node49856 = (inp[7]) ? node50530 : node49857;
								assign node49857 = (inp[8]) ? node50181 : node49858;
									assign node49858 = (inp[14]) ? node50052 : node49859;
										assign node49859 = (inp[2]) ? node49963 : node49860;
											assign node49860 = (inp[0]) ? node49914 : node49861;
												assign node49861 = (inp[15]) ? node49889 : node49862;
													assign node49862 = (inp[3]) ? node49878 : node49863;
														assign node49863 = (inp[4]) ? node49871 : node49864;
															assign node49864 = (inp[9]) ? node49868 : node49865;
																assign node49865 = (inp[10]) ? 4'b1011 : 4'b1111;
																assign node49868 = (inp[10]) ? 4'b1111 : 4'b1011;
															assign node49871 = (inp[9]) ? node49875 : node49872;
																assign node49872 = (inp[10]) ? 4'b1111 : 4'b1011;
																assign node49875 = (inp[10]) ? 4'b1011 : 4'b1111;
														assign node49878 = (inp[4]) ? node49884 : node49879;
															assign node49879 = (inp[10]) ? node49881 : 4'b1011;
																assign node49881 = (inp[9]) ? 4'b1101 : 4'b1011;
															assign node49884 = (inp[10]) ? node49886 : 4'b1101;
																assign node49886 = (inp[9]) ? 4'b1001 : 4'b1101;
													assign node49889 = (inp[3]) ? node49905 : node49890;
														assign node49890 = (inp[4]) ? node49898 : node49891;
															assign node49891 = (inp[9]) ? node49895 : node49892;
																assign node49892 = (inp[10]) ? 4'b1001 : 4'b1101;
																assign node49895 = (inp[10]) ? 4'b1101 : 4'b1001;
															assign node49898 = (inp[9]) ? node49902 : node49899;
																assign node49899 = (inp[10]) ? 4'b1101 : 4'b1001;
																assign node49902 = (inp[10]) ? 4'b1001 : 4'b1101;
														assign node49905 = (inp[4]) ? node49911 : node49906;
															assign node49906 = (inp[9]) ? 4'b1001 : node49907;
																assign node49907 = (inp[10]) ? 4'b1001 : 4'b1101;
															assign node49911 = (inp[10]) ? 4'b1111 : 4'b1001;
												assign node49914 = (inp[15]) ? node49936 : node49915;
													assign node49915 = (inp[4]) ? node49923 : node49916;
														assign node49916 = (inp[9]) ? node49920 : node49917;
															assign node49917 = (inp[10]) ? 4'b1001 : 4'b1101;
															assign node49920 = (inp[10]) ? 4'b1101 : 4'b1001;
														assign node49923 = (inp[3]) ? node49929 : node49924;
															assign node49924 = (inp[9]) ? node49926 : 4'b1001;
																assign node49926 = (inp[10]) ? 4'b1001 : 4'b1101;
															assign node49929 = (inp[9]) ? node49933 : node49930;
																assign node49930 = (inp[10]) ? 4'b1111 : 4'b1001;
																assign node49933 = (inp[10]) ? 4'b1011 : 4'b1111;
													assign node49936 = (inp[3]) ? node49950 : node49937;
														assign node49937 = (inp[9]) ? node49943 : node49938;
															assign node49938 = (inp[10]) ? 4'b1011 : node49939;
																assign node49939 = (inp[4]) ? 4'b1011 : 4'b1111;
															assign node49943 = (inp[10]) ? node49947 : node49944;
																assign node49944 = (inp[4]) ? 4'b1111 : 4'b1011;
																assign node49947 = (inp[4]) ? 4'b1011 : 4'b1111;
														assign node49950 = (inp[9]) ? node49956 : node49951;
															assign node49951 = (inp[10]) ? 4'b1011 : node49952;
																assign node49952 = (inp[4]) ? 4'b1011 : 4'b1111;
															assign node49956 = (inp[10]) ? node49960 : node49957;
																assign node49957 = (inp[4]) ? 4'b1101 : 4'b1011;
																assign node49960 = (inp[4]) ? 4'b1001 : 4'b1101;
											assign node49963 = (inp[15]) ? node50017 : node49964;
												assign node49964 = (inp[0]) ? node49990 : node49965;
													assign node49965 = (inp[3]) ? node49979 : node49966;
														assign node49966 = (inp[9]) ? node49972 : node49967;
															assign node49967 = (inp[10]) ? 4'b1110 : node49968;
																assign node49968 = (inp[4]) ? 4'b1010 : 4'b1110;
															assign node49972 = (inp[10]) ? node49976 : node49973;
																assign node49973 = (inp[4]) ? 4'b1110 : 4'b1010;
																assign node49976 = (inp[4]) ? 4'b1010 : 4'b1110;
														assign node49979 = (inp[4]) ? node49985 : node49980;
															assign node49980 = (inp[10]) ? 4'b1010 : node49981;
																assign node49981 = (inp[9]) ? 4'b1010 : 4'b1110;
															assign node49985 = (inp[9]) ? node49987 : 4'b1100;
																assign node49987 = (inp[10]) ? 4'b1000 : 4'b1100;
													assign node49990 = (inp[3]) ? node50004 : node49991;
														assign node49991 = (inp[10]) ? node49997 : node49992;
															assign node49992 = (inp[9]) ? 4'b1000 : node49993;
																assign node49993 = (inp[4]) ? 4'b1000 : 4'b1100;
															assign node49997 = (inp[4]) ? node50001 : node49998;
																assign node49998 = (inp[9]) ? 4'b1100 : 4'b1000;
																assign node50001 = (inp[9]) ? 4'b1000 : 4'b1100;
														assign node50004 = (inp[10]) ? node50010 : node50005;
															assign node50005 = (inp[9]) ? node50007 : 4'b1000;
																assign node50007 = (inp[4]) ? 4'b1110 : 4'b1000;
															assign node50010 = (inp[4]) ? node50014 : node50011;
																assign node50011 = (inp[9]) ? 4'b1110 : 4'b1000;
																assign node50014 = (inp[9]) ? 4'b1010 : 4'b1110;
												assign node50017 = (inp[0]) ? node50033 : node50018;
													assign node50018 = (inp[3]) ? node50026 : node50019;
														assign node50019 = (inp[4]) ? node50021 : 4'b1000;
															assign node50021 = (inp[9]) ? node50023 : 4'b1000;
																assign node50023 = (inp[10]) ? 4'b1000 : 4'b1100;
														assign node50026 = (inp[4]) ? node50030 : node50027;
															assign node50027 = (inp[9]) ? 4'b1000 : 4'b1100;
															assign node50030 = (inp[10]) ? 4'b1010 : 4'b1110;
													assign node50033 = (inp[3]) ? node50045 : node50034;
														assign node50034 = (inp[4]) ? node50040 : node50035;
															assign node50035 = (inp[10]) ? node50037 : 4'b1010;
																assign node50037 = (inp[9]) ? 4'b1110 : 4'b1010;
															assign node50040 = (inp[10]) ? node50042 : 4'b1110;
																assign node50042 = (inp[9]) ? 4'b1010 : 4'b1110;
														assign node50045 = (inp[9]) ? 4'b1000 : node50046;
															assign node50046 = (inp[4]) ? 4'b1010 : node50047;
																assign node50047 = (inp[10]) ? 4'b1010 : 4'b1110;
										assign node50052 = (inp[0]) ? node50124 : node50053;
											assign node50053 = (inp[15]) ? node50091 : node50054;
												assign node50054 = (inp[3]) ? node50074 : node50055;
													assign node50055 = (inp[2]) ? node50067 : node50056;
														assign node50056 = (inp[4]) ? node50062 : node50057;
															assign node50057 = (inp[9]) ? node50059 : 4'b1010;
																assign node50059 = (inp[10]) ? 4'b1110 : 4'b1010;
															assign node50062 = (inp[10]) ? node50064 : 4'b1110;
																assign node50064 = (inp[9]) ? 4'b1010 : 4'b1110;
														assign node50067 = (inp[4]) ? 4'b1010 : node50068;
															assign node50068 = (inp[10]) ? 4'b1010 : node50069;
																assign node50069 = (inp[9]) ? 4'b1010 : 4'b1110;
													assign node50074 = (inp[10]) ? node50084 : node50075;
														assign node50075 = (inp[2]) ? node50077 : 4'b1010;
															assign node50077 = (inp[9]) ? node50081 : node50078;
																assign node50078 = (inp[4]) ? 4'b1010 : 4'b1110;
																assign node50081 = (inp[4]) ? 4'b1100 : 4'b1010;
														assign node50084 = (inp[4]) ? node50088 : node50085;
															assign node50085 = (inp[9]) ? 4'b1100 : 4'b1010;
															assign node50088 = (inp[9]) ? 4'b1000 : 4'b1100;
												assign node50091 = (inp[3]) ? node50109 : node50092;
													assign node50092 = (inp[9]) ? node50100 : node50093;
														assign node50093 = (inp[2]) ? node50095 : 4'b1000;
															assign node50095 = (inp[4]) ? node50097 : 4'b1000;
																assign node50097 = (inp[10]) ? 4'b1100 : 4'b1000;
														assign node50100 = (inp[2]) ? 4'b1100 : node50101;
															assign node50101 = (inp[10]) ? node50105 : node50102;
																assign node50102 = (inp[4]) ? 4'b1100 : 4'b1000;
																assign node50105 = (inp[4]) ? 4'b1000 : 4'b1100;
													assign node50109 = (inp[10]) ? node50119 : node50110;
														assign node50110 = (inp[2]) ? node50112 : 4'b1000;
															assign node50112 = (inp[4]) ? node50116 : node50113;
																assign node50113 = (inp[9]) ? 4'b1000 : 4'b1100;
																assign node50116 = (inp[9]) ? 4'b1110 : 4'b1000;
														assign node50119 = (inp[9]) ? node50121 : 4'b1110;
															assign node50121 = (inp[4]) ? 4'b1010 : 4'b1110;
											assign node50124 = (inp[15]) ? node50150 : node50125;
												assign node50125 = (inp[3]) ? node50135 : node50126;
													assign node50126 = (inp[9]) ? 4'b1000 : node50127;
														assign node50127 = (inp[10]) ? node50131 : node50128;
															assign node50128 = (inp[4]) ? 4'b1000 : 4'b1100;
															assign node50131 = (inp[4]) ? 4'b1100 : 4'b1000;
													assign node50135 = (inp[9]) ? node50143 : node50136;
														assign node50136 = (inp[10]) ? node50140 : node50137;
															assign node50137 = (inp[4]) ? 4'b1000 : 4'b1100;
															assign node50140 = (inp[4]) ? 4'b1110 : 4'b1000;
														assign node50143 = (inp[10]) ? node50147 : node50144;
															assign node50144 = (inp[4]) ? 4'b1110 : 4'b1000;
															assign node50147 = (inp[4]) ? 4'b1010 : 4'b1110;
												assign node50150 = (inp[3]) ? node50166 : node50151;
													assign node50151 = (inp[4]) ? node50159 : node50152;
														assign node50152 = (inp[10]) ? node50156 : node50153;
															assign node50153 = (inp[9]) ? 4'b1010 : 4'b1110;
															assign node50156 = (inp[9]) ? 4'b1110 : 4'b1010;
														assign node50159 = (inp[10]) ? node50163 : node50160;
															assign node50160 = (inp[9]) ? 4'b1110 : 4'b1010;
															assign node50163 = (inp[9]) ? 4'b1010 : 4'b1110;
													assign node50166 = (inp[4]) ? node50172 : node50167;
														assign node50167 = (inp[10]) ? node50169 : 4'b1010;
															assign node50169 = (inp[9]) ? 4'b1100 : 4'b1010;
														assign node50172 = (inp[2]) ? node50174 : 4'b1100;
															assign node50174 = (inp[9]) ? node50178 : node50175;
																assign node50175 = (inp[10]) ? 4'b1100 : 4'b1010;
																assign node50178 = (inp[10]) ? 4'b1000 : 4'b1100;
									assign node50181 = (inp[2]) ? node50353 : node50182;
										assign node50182 = (inp[14]) ? node50266 : node50183;
											assign node50183 = (inp[10]) ? node50213 : node50184;
												assign node50184 = (inp[0]) ? node50202 : node50185;
													assign node50185 = (inp[15]) ? node50195 : node50186;
														assign node50186 = (inp[9]) ? node50190 : node50187;
															assign node50187 = (inp[4]) ? 4'b1010 : 4'b1110;
															assign node50190 = (inp[4]) ? node50192 : 4'b1010;
																assign node50192 = (inp[3]) ? 4'b1100 : 4'b1110;
														assign node50195 = (inp[4]) ? node50199 : node50196;
															assign node50196 = (inp[9]) ? 4'b1000 : 4'b1100;
															assign node50199 = (inp[9]) ? 4'b1110 : 4'b1000;
													assign node50202 = (inp[15]) ? node50204 : 4'b1000;
														assign node50204 = (inp[3]) ? node50210 : node50205;
															assign node50205 = (inp[9]) ? 4'b1010 : node50206;
																assign node50206 = (inp[4]) ? 4'b1010 : 4'b1110;
															assign node50210 = (inp[4]) ? 4'b1100 : 4'b1010;
												assign node50213 = (inp[0]) ? node50237 : node50214;
													assign node50214 = (inp[15]) ? node50224 : node50215;
														assign node50215 = (inp[3]) ? node50221 : node50216;
															assign node50216 = (inp[4]) ? 4'b1110 : node50217;
																assign node50217 = (inp[9]) ? 4'b1110 : 4'b1010;
															assign node50221 = (inp[9]) ? 4'b1000 : 4'b1100;
														assign node50224 = (inp[3]) ? node50232 : node50225;
															assign node50225 = (inp[9]) ? node50229 : node50226;
																assign node50226 = (inp[4]) ? 4'b1100 : 4'b1000;
																assign node50229 = (inp[4]) ? 4'b1000 : 4'b1100;
															assign node50232 = (inp[9]) ? 4'b1110 : node50233;
																assign node50233 = (inp[4]) ? 4'b1110 : 4'b1000;
													assign node50237 = (inp[15]) ? node50253 : node50238;
														assign node50238 = (inp[3]) ? node50246 : node50239;
															assign node50239 = (inp[9]) ? node50243 : node50240;
																assign node50240 = (inp[4]) ? 4'b1100 : 4'b1000;
																assign node50243 = (inp[4]) ? 4'b1000 : 4'b1100;
															assign node50246 = (inp[4]) ? node50250 : node50247;
																assign node50247 = (inp[9]) ? 4'b1110 : 4'b1000;
																assign node50250 = (inp[9]) ? 4'b1010 : 4'b1110;
														assign node50253 = (inp[3]) ? node50259 : node50254;
															assign node50254 = (inp[4]) ? 4'b1010 : node50255;
																assign node50255 = (inp[9]) ? 4'b1110 : 4'b1010;
															assign node50259 = (inp[4]) ? node50263 : node50260;
																assign node50260 = (inp[9]) ? 4'b1100 : 4'b1010;
																assign node50263 = (inp[9]) ? 4'b1000 : 4'b1100;
											assign node50266 = (inp[4]) ? node50306 : node50267;
												assign node50267 = (inp[9]) ? node50281 : node50268;
													assign node50268 = (inp[10]) ? node50274 : node50269;
														assign node50269 = (inp[15]) ? node50271 : 4'b1111;
															assign node50271 = (inp[0]) ? 4'b1111 : 4'b1101;
														assign node50274 = (inp[15]) ? node50278 : node50275;
															assign node50275 = (inp[0]) ? 4'b1001 : 4'b1011;
															assign node50278 = (inp[0]) ? 4'b1011 : 4'b1001;
													assign node50281 = (inp[10]) ? node50293 : node50282;
														assign node50282 = (inp[3]) ? node50288 : node50283;
															assign node50283 = (inp[0]) ? node50285 : 4'b1011;
																assign node50285 = (inp[15]) ? 4'b1011 : 4'b1001;
															assign node50288 = (inp[15]) ? node50290 : 4'b1001;
																assign node50290 = (inp[0]) ? 4'b1011 : 4'b1001;
														assign node50293 = (inp[0]) ? node50301 : node50294;
															assign node50294 = (inp[3]) ? node50298 : node50295;
																assign node50295 = (inp[15]) ? 4'b1101 : 4'b1111;
																assign node50298 = (inp[15]) ? 4'b1111 : 4'b1101;
															assign node50301 = (inp[15]) ? node50303 : 4'b1111;
																assign node50303 = (inp[3]) ? 4'b1101 : 4'b1111;
												assign node50306 = (inp[0]) ? node50324 : node50307;
													assign node50307 = (inp[15]) ? node50315 : node50308;
														assign node50308 = (inp[3]) ? node50310 : 4'b1011;
															assign node50310 = (inp[10]) ? node50312 : 4'b1011;
																assign node50312 = (inp[9]) ? 4'b1001 : 4'b1101;
														assign node50315 = (inp[3]) ? node50321 : node50316;
															assign node50316 = (inp[10]) ? node50318 : 4'b1101;
																assign node50318 = (inp[9]) ? 4'b1001 : 4'b1101;
															assign node50321 = (inp[9]) ? 4'b1011 : 4'b1001;
													assign node50324 = (inp[15]) ? node50338 : node50325;
														assign node50325 = (inp[3]) ? node50333 : node50326;
															assign node50326 = (inp[9]) ? node50330 : node50327;
																assign node50327 = (inp[10]) ? 4'b1101 : 4'b1001;
																assign node50330 = (inp[10]) ? 4'b1001 : 4'b1101;
															assign node50333 = (inp[9]) ? node50335 : 4'b1001;
																assign node50335 = (inp[10]) ? 4'b1011 : 4'b1111;
														assign node50338 = (inp[3]) ? node50346 : node50339;
															assign node50339 = (inp[9]) ? node50343 : node50340;
																assign node50340 = (inp[10]) ? 4'b1111 : 4'b1011;
																assign node50343 = (inp[10]) ? 4'b1011 : 4'b1111;
															assign node50346 = (inp[10]) ? node50350 : node50347;
																assign node50347 = (inp[9]) ? 4'b1101 : 4'b1011;
																assign node50350 = (inp[9]) ? 4'b1001 : 4'b1101;
										assign node50353 = (inp[14]) ? node50449 : node50354;
											assign node50354 = (inp[3]) ? node50398 : node50355;
												assign node50355 = (inp[15]) ? node50375 : node50356;
													assign node50356 = (inp[0]) ? node50366 : node50357;
														assign node50357 = (inp[4]) ? 4'b1111 : node50358;
															assign node50358 = (inp[9]) ? node50362 : node50359;
																assign node50359 = (inp[10]) ? 4'b1011 : 4'b1111;
																assign node50362 = (inp[10]) ? 4'b1111 : 4'b1011;
														assign node50366 = (inp[10]) ? 4'b1101 : node50367;
															assign node50367 = (inp[4]) ? node50371 : node50368;
																assign node50368 = (inp[9]) ? 4'b1001 : 4'b1101;
																assign node50371 = (inp[9]) ? 4'b1101 : 4'b1001;
													assign node50375 = (inp[0]) ? node50383 : node50376;
														assign node50376 = (inp[9]) ? 4'b1101 : node50377;
															assign node50377 = (inp[4]) ? 4'b1001 : node50378;
																assign node50378 = (inp[10]) ? 4'b1001 : 4'b1101;
														assign node50383 = (inp[9]) ? node50391 : node50384;
															assign node50384 = (inp[10]) ? node50388 : node50385;
																assign node50385 = (inp[4]) ? 4'b1011 : 4'b1111;
																assign node50388 = (inp[4]) ? 4'b1111 : 4'b1011;
															assign node50391 = (inp[10]) ? node50395 : node50392;
																assign node50392 = (inp[4]) ? 4'b1111 : 4'b1011;
																assign node50395 = (inp[4]) ? 4'b1011 : 4'b1111;
												assign node50398 = (inp[0]) ? node50428 : node50399;
													assign node50399 = (inp[10]) ? node50415 : node50400;
														assign node50400 = (inp[15]) ? node50408 : node50401;
															assign node50401 = (inp[4]) ? node50405 : node50402;
																assign node50402 = (inp[9]) ? 4'b1011 : 4'b1111;
																assign node50405 = (inp[9]) ? 4'b1101 : 4'b1011;
															assign node50408 = (inp[9]) ? node50412 : node50409;
																assign node50409 = (inp[4]) ? 4'b1001 : 4'b1101;
																assign node50412 = (inp[4]) ? 4'b1111 : 4'b1001;
														assign node50415 = (inp[15]) ? node50423 : node50416;
															assign node50416 = (inp[9]) ? node50420 : node50417;
																assign node50417 = (inp[4]) ? 4'b1101 : 4'b1011;
																assign node50420 = (inp[4]) ? 4'b1001 : 4'b1101;
															assign node50423 = (inp[4]) ? node50425 : 4'b1001;
																assign node50425 = (inp[9]) ? 4'b1011 : 4'b1111;
													assign node50428 = (inp[10]) ? node50442 : node50429;
														assign node50429 = (inp[15]) ? node50437 : node50430;
															assign node50430 = (inp[4]) ? node50434 : node50431;
																assign node50431 = (inp[9]) ? 4'b1001 : 4'b1101;
																assign node50434 = (inp[9]) ? 4'b1111 : 4'b1001;
															assign node50437 = (inp[9]) ? 4'b1101 : node50438;
																assign node50438 = (inp[4]) ? 4'b1011 : 4'b1111;
														assign node50442 = (inp[15]) ? 4'b1101 : node50443;
															assign node50443 = (inp[4]) ? 4'b1111 : node50444;
																assign node50444 = (inp[9]) ? 4'b1111 : 4'b1001;
											assign node50449 = (inp[15]) ? node50489 : node50450;
												assign node50450 = (inp[0]) ? node50468 : node50451;
													assign node50451 = (inp[10]) ? node50459 : node50452;
														assign node50452 = (inp[4]) ? node50456 : node50453;
															assign node50453 = (inp[9]) ? 4'b1011 : 4'b1111;
															assign node50456 = (inp[9]) ? 4'b1111 : 4'b1011;
														assign node50459 = (inp[3]) ? node50463 : node50460;
															assign node50460 = (inp[9]) ? 4'b1011 : 4'b1111;
															assign node50463 = (inp[9]) ? node50465 : 4'b1011;
																assign node50465 = (inp[4]) ? 4'b1001 : 4'b1101;
													assign node50468 = (inp[3]) ? node50474 : node50469;
														assign node50469 = (inp[4]) ? 4'b1001 : node50470;
															assign node50470 = (inp[9]) ? 4'b1101 : 4'b1001;
														assign node50474 = (inp[4]) ? node50482 : node50475;
															assign node50475 = (inp[10]) ? node50479 : node50476;
																assign node50476 = (inp[9]) ? 4'b1001 : 4'b1101;
																assign node50479 = (inp[9]) ? 4'b1111 : 4'b1001;
															assign node50482 = (inp[9]) ? node50486 : node50483;
																assign node50483 = (inp[10]) ? 4'b1111 : 4'b1001;
																assign node50486 = (inp[10]) ? 4'b1011 : 4'b1111;
												assign node50489 = (inp[0]) ? node50513 : node50490;
													assign node50490 = (inp[3]) ? node50500 : node50491;
														assign node50491 = (inp[9]) ? 4'b1001 : node50492;
															assign node50492 = (inp[10]) ? node50496 : node50493;
																assign node50493 = (inp[4]) ? 4'b1001 : 4'b1101;
																assign node50496 = (inp[4]) ? 4'b1101 : 4'b1001;
														assign node50500 = (inp[9]) ? node50506 : node50501;
															assign node50501 = (inp[4]) ? node50503 : 4'b1001;
																assign node50503 = (inp[10]) ? 4'b1111 : 4'b1001;
															assign node50506 = (inp[4]) ? node50510 : node50507;
																assign node50507 = (inp[10]) ? 4'b1111 : 4'b1001;
																assign node50510 = (inp[10]) ? 4'b1011 : 4'b1111;
													assign node50513 = (inp[4]) ? node50523 : node50514;
														assign node50514 = (inp[9]) ? node50518 : node50515;
															assign node50515 = (inp[10]) ? 4'b1011 : 4'b1111;
															assign node50518 = (inp[10]) ? node50520 : 4'b1011;
																assign node50520 = (inp[3]) ? 4'b1101 : 4'b1111;
														assign node50523 = (inp[3]) ? node50525 : 4'b1111;
															assign node50525 = (inp[10]) ? node50527 : 4'b1101;
																assign node50527 = (inp[9]) ? 4'b1001 : 4'b1101;
								assign node50530 = (inp[8]) ? node50826 : node50531;
									assign node50531 = (inp[2]) ? node50709 : node50532;
										assign node50532 = (inp[14]) ? node50632 : node50533;
											assign node50533 = (inp[4]) ? node50583 : node50534;
												assign node50534 = (inp[3]) ? node50556 : node50535;
													assign node50535 = (inp[0]) ? node50549 : node50536;
														assign node50536 = (inp[15]) ? node50542 : node50537;
															assign node50537 = (inp[10]) ? 4'b1010 : node50538;
																assign node50538 = (inp[9]) ? 4'b1010 : 4'b1110;
															assign node50542 = (inp[9]) ? node50546 : node50543;
																assign node50543 = (inp[10]) ? 4'b1000 : 4'b1100;
																assign node50546 = (inp[10]) ? 4'b1100 : 4'b1000;
														assign node50549 = (inp[15]) ? node50551 : 4'b1000;
															assign node50551 = (inp[9]) ? 4'b1010 : node50552;
																assign node50552 = (inp[10]) ? 4'b1010 : 4'b1110;
													assign node50556 = (inp[0]) ? node50570 : node50557;
														assign node50557 = (inp[15]) ? node50565 : node50558;
															assign node50558 = (inp[10]) ? node50562 : node50559;
																assign node50559 = (inp[9]) ? 4'b1010 : 4'b1110;
																assign node50562 = (inp[9]) ? 4'b1100 : 4'b1010;
															assign node50565 = (inp[9]) ? node50567 : 4'b1000;
																assign node50567 = (inp[10]) ? 4'b1110 : 4'b1000;
														assign node50570 = (inp[15]) ? node50578 : node50571;
															assign node50571 = (inp[9]) ? node50575 : node50572;
																assign node50572 = (inp[10]) ? 4'b1000 : 4'b1100;
																assign node50575 = (inp[10]) ? 4'b1110 : 4'b1000;
															assign node50578 = (inp[9]) ? 4'b1100 : node50579;
																assign node50579 = (inp[10]) ? 4'b1010 : 4'b1110;
												assign node50583 = (inp[3]) ? node50607 : node50584;
													assign node50584 = (inp[0]) ? node50594 : node50585;
														assign node50585 = (inp[15]) ? node50587 : 4'b1110;
															assign node50587 = (inp[10]) ? node50591 : node50588;
																assign node50588 = (inp[9]) ? 4'b1100 : 4'b1000;
																assign node50591 = (inp[9]) ? 4'b1000 : 4'b1100;
														assign node50594 = (inp[15]) ? node50602 : node50595;
															assign node50595 = (inp[10]) ? node50599 : node50596;
																assign node50596 = (inp[9]) ? 4'b1100 : 4'b1000;
																assign node50599 = (inp[9]) ? 4'b1000 : 4'b1100;
															assign node50602 = (inp[10]) ? node50604 : 4'b1110;
																assign node50604 = (inp[9]) ? 4'b1010 : 4'b1110;
													assign node50607 = (inp[10]) ? node50617 : node50608;
														assign node50608 = (inp[9]) ? node50610 : 4'b1010;
															assign node50610 = (inp[15]) ? node50614 : node50611;
																assign node50611 = (inp[0]) ? 4'b1110 : 4'b1100;
																assign node50614 = (inp[0]) ? 4'b1100 : 4'b1110;
														assign node50617 = (inp[9]) ? node50625 : node50618;
															assign node50618 = (inp[15]) ? node50622 : node50619;
																assign node50619 = (inp[0]) ? 4'b1110 : 4'b1100;
																assign node50622 = (inp[0]) ? 4'b1100 : 4'b1110;
															assign node50625 = (inp[15]) ? node50629 : node50626;
																assign node50626 = (inp[0]) ? 4'b1010 : 4'b1000;
																assign node50629 = (inp[0]) ? 4'b1000 : 4'b1010;
											assign node50632 = (inp[10]) ? node50668 : node50633;
												assign node50633 = (inp[0]) ? node50655 : node50634;
													assign node50634 = (inp[15]) ? node50646 : node50635;
														assign node50635 = (inp[3]) ? node50641 : node50636;
															assign node50636 = (inp[4]) ? 4'b1111 : node50637;
																assign node50637 = (inp[9]) ? 4'b1011 : 4'b1111;
															assign node50641 = (inp[9]) ? 4'b1011 : node50642;
																assign node50642 = (inp[4]) ? 4'b1011 : 4'b1111;
														assign node50646 = (inp[9]) ? node50650 : node50647;
															assign node50647 = (inp[4]) ? 4'b1001 : 4'b1101;
															assign node50650 = (inp[4]) ? node50652 : 4'b1001;
																assign node50652 = (inp[3]) ? 4'b1111 : 4'b1101;
													assign node50655 = (inp[15]) ? node50661 : node50656;
														assign node50656 = (inp[9]) ? node50658 : 4'b1001;
															assign node50658 = (inp[4]) ? 4'b1111 : 4'b1001;
														assign node50661 = (inp[9]) ? node50665 : node50662;
															assign node50662 = (inp[4]) ? 4'b1011 : 4'b1111;
															assign node50665 = (inp[4]) ? 4'b1111 : 4'b1011;
												assign node50668 = (inp[3]) ? node50694 : node50669;
													assign node50669 = (inp[4]) ? node50685 : node50670;
														assign node50670 = (inp[9]) ? node50678 : node50671;
															assign node50671 = (inp[0]) ? node50675 : node50672;
																assign node50672 = (inp[15]) ? 4'b1001 : 4'b1011;
																assign node50675 = (inp[15]) ? 4'b1011 : 4'b1001;
															assign node50678 = (inp[0]) ? node50682 : node50679;
																assign node50679 = (inp[15]) ? 4'b1101 : 4'b1111;
																assign node50682 = (inp[15]) ? 4'b1111 : 4'b1101;
														assign node50685 = (inp[9]) ? node50687 : 4'b1101;
															assign node50687 = (inp[0]) ? node50691 : node50688;
																assign node50688 = (inp[15]) ? 4'b1001 : 4'b1011;
																assign node50691 = (inp[15]) ? 4'b1011 : 4'b1001;
													assign node50694 = (inp[9]) ? node50706 : node50695;
														assign node50695 = (inp[4]) ? node50701 : node50696;
															assign node50696 = (inp[15]) ? 4'b1001 : node50697;
																assign node50697 = (inp[0]) ? 4'b1001 : 4'b1011;
															assign node50701 = (inp[0]) ? 4'b1111 : node50702;
																assign node50702 = (inp[15]) ? 4'b1111 : 4'b1101;
														assign node50706 = (inp[4]) ? 4'b1001 : 4'b1101;
										assign node50709 = (inp[4]) ? node50761 : node50710;
											assign node50710 = (inp[0]) ? node50736 : node50711;
												assign node50711 = (inp[15]) ? node50727 : node50712;
													assign node50712 = (inp[3]) ? node50720 : node50713;
														assign node50713 = (inp[9]) ? node50717 : node50714;
															assign node50714 = (inp[10]) ? 4'b1011 : 4'b1111;
															assign node50717 = (inp[10]) ? 4'b1111 : 4'b1011;
														assign node50720 = (inp[9]) ? node50724 : node50721;
															assign node50721 = (inp[10]) ? 4'b1011 : 4'b1111;
															assign node50724 = (inp[10]) ? 4'b1101 : 4'b1011;
													assign node50727 = (inp[10]) ? node50731 : node50728;
														assign node50728 = (inp[9]) ? 4'b1001 : 4'b1101;
														assign node50731 = (inp[9]) ? node50733 : 4'b1001;
															assign node50733 = (inp[14]) ? 4'b1111 : 4'b1101;
												assign node50736 = (inp[15]) ? node50746 : node50737;
													assign node50737 = (inp[9]) ? node50741 : node50738;
														assign node50738 = (inp[10]) ? 4'b1001 : 4'b1101;
														assign node50741 = (inp[10]) ? node50743 : 4'b1001;
															assign node50743 = (inp[3]) ? 4'b1111 : 4'b1101;
													assign node50746 = (inp[3]) ? node50754 : node50747;
														assign node50747 = (inp[9]) ? node50751 : node50748;
															assign node50748 = (inp[10]) ? 4'b1011 : 4'b1111;
															assign node50751 = (inp[10]) ? 4'b1111 : 4'b1011;
														assign node50754 = (inp[10]) ? node50758 : node50755;
															assign node50755 = (inp[9]) ? 4'b1011 : 4'b1111;
															assign node50758 = (inp[9]) ? 4'b1101 : 4'b1011;
											assign node50761 = (inp[15]) ? node50793 : node50762;
												assign node50762 = (inp[0]) ? node50778 : node50763;
													assign node50763 = (inp[3]) ? node50771 : node50764;
														assign node50764 = (inp[10]) ? node50768 : node50765;
															assign node50765 = (inp[9]) ? 4'b1111 : 4'b1011;
															assign node50768 = (inp[9]) ? 4'b1011 : 4'b1111;
														assign node50771 = (inp[9]) ? node50775 : node50772;
															assign node50772 = (inp[10]) ? 4'b1101 : 4'b1011;
															assign node50775 = (inp[10]) ? 4'b1001 : 4'b1101;
													assign node50778 = (inp[3]) ? node50786 : node50779;
														assign node50779 = (inp[14]) ? 4'b1001 : node50780;
															assign node50780 = (inp[10]) ? node50782 : 4'b1101;
																assign node50782 = (inp[9]) ? 4'b1001 : 4'b1101;
														assign node50786 = (inp[10]) ? node50790 : node50787;
															assign node50787 = (inp[14]) ? 4'b1111 : 4'b1001;
															assign node50790 = (inp[9]) ? 4'b1011 : 4'b1111;
												assign node50793 = (inp[0]) ? node50809 : node50794;
													assign node50794 = (inp[3]) ? node50802 : node50795;
														assign node50795 = (inp[9]) ? node50799 : node50796;
															assign node50796 = (inp[10]) ? 4'b1101 : 4'b1001;
															assign node50799 = (inp[10]) ? 4'b1001 : 4'b1101;
														assign node50802 = (inp[10]) ? node50806 : node50803;
															assign node50803 = (inp[9]) ? 4'b1111 : 4'b1001;
															assign node50806 = (inp[9]) ? 4'b1011 : 4'b1111;
													assign node50809 = (inp[3]) ? node50819 : node50810;
														assign node50810 = (inp[14]) ? node50812 : 4'b1011;
															assign node50812 = (inp[10]) ? node50816 : node50813;
																assign node50813 = (inp[9]) ? 4'b1111 : 4'b1011;
																assign node50816 = (inp[9]) ? 4'b1011 : 4'b1111;
														assign node50819 = (inp[10]) ? node50823 : node50820;
															assign node50820 = (inp[9]) ? 4'b1101 : 4'b1011;
															assign node50823 = (inp[9]) ? 4'b1001 : 4'b1101;
									assign node50826 = (inp[2]) ? node51016 : node50827;
										assign node50827 = (inp[14]) ? node50921 : node50828;
											assign node50828 = (inp[3]) ? node50874 : node50829;
												assign node50829 = (inp[15]) ? node50853 : node50830;
													assign node50830 = (inp[0]) ? node50844 : node50831;
														assign node50831 = (inp[9]) ? node50839 : node50832;
															assign node50832 = (inp[10]) ? node50836 : node50833;
																assign node50833 = (inp[4]) ? 4'b1011 : 4'b1111;
																assign node50836 = (inp[4]) ? 4'b1111 : 4'b1011;
															assign node50839 = (inp[10]) ? 4'b1111 : node50840;
																assign node50840 = (inp[4]) ? 4'b1111 : 4'b1011;
														assign node50844 = (inp[10]) ? 4'b1101 : node50845;
															assign node50845 = (inp[4]) ? node50849 : node50846;
																assign node50846 = (inp[9]) ? 4'b1001 : 4'b1101;
																assign node50849 = (inp[9]) ? 4'b1101 : 4'b1001;
													assign node50853 = (inp[0]) ? node50867 : node50854;
														assign node50854 = (inp[9]) ? node50862 : node50855;
															assign node50855 = (inp[4]) ? node50859 : node50856;
																assign node50856 = (inp[10]) ? 4'b1001 : 4'b1101;
																assign node50859 = (inp[10]) ? 4'b1101 : 4'b1001;
															assign node50862 = (inp[10]) ? node50864 : 4'b1101;
																assign node50864 = (inp[4]) ? 4'b1001 : 4'b1101;
														assign node50867 = (inp[4]) ? node50869 : 4'b1011;
															assign node50869 = (inp[10]) ? 4'b1111 : node50870;
																assign node50870 = (inp[9]) ? 4'b1111 : 4'b1011;
												assign node50874 = (inp[0]) ? node50894 : node50875;
													assign node50875 = (inp[15]) ? node50883 : node50876;
														assign node50876 = (inp[9]) ? node50878 : 4'b1011;
															assign node50878 = (inp[10]) ? node50880 : 4'b1011;
																assign node50880 = (inp[4]) ? 4'b1001 : 4'b1101;
														assign node50883 = (inp[4]) ? node50889 : node50884;
															assign node50884 = (inp[9]) ? 4'b1001 : node50885;
																assign node50885 = (inp[10]) ? 4'b1001 : 4'b1101;
															assign node50889 = (inp[10]) ? 4'b1111 : node50890;
																assign node50890 = (inp[9]) ? 4'b1111 : 4'b1001;
													assign node50894 = (inp[15]) ? node50910 : node50895;
														assign node50895 = (inp[10]) ? node50903 : node50896;
															assign node50896 = (inp[4]) ? node50900 : node50897;
																assign node50897 = (inp[9]) ? 4'b1001 : 4'b1101;
																assign node50900 = (inp[9]) ? 4'b1111 : 4'b1001;
															assign node50903 = (inp[4]) ? node50907 : node50904;
																assign node50904 = (inp[9]) ? 4'b1111 : 4'b1001;
																assign node50907 = (inp[9]) ? 4'b1011 : 4'b1111;
														assign node50910 = (inp[10]) ? node50916 : node50911;
															assign node50911 = (inp[4]) ? 4'b1011 : node50912;
																assign node50912 = (inp[9]) ? 4'b1011 : 4'b1111;
															assign node50916 = (inp[4]) ? node50918 : 4'b1011;
																assign node50918 = (inp[9]) ? 4'b1001 : 4'b1101;
											assign node50921 = (inp[3]) ? node50971 : node50922;
												assign node50922 = (inp[4]) ? node50952 : node50923;
													assign node50923 = (inp[0]) ? node50937 : node50924;
														assign node50924 = (inp[15]) ? node50932 : node50925;
															assign node50925 = (inp[10]) ? node50929 : node50926;
																assign node50926 = (inp[9]) ? 4'b1010 : 4'b1110;
																assign node50929 = (inp[9]) ? 4'b1110 : 4'b1010;
															assign node50932 = (inp[10]) ? 4'b1000 : node50933;
																assign node50933 = (inp[9]) ? 4'b1000 : 4'b1100;
														assign node50937 = (inp[15]) ? node50945 : node50938;
															assign node50938 = (inp[10]) ? node50942 : node50939;
																assign node50939 = (inp[9]) ? 4'b1000 : 4'b1100;
																assign node50942 = (inp[9]) ? 4'b1100 : 4'b1000;
															assign node50945 = (inp[10]) ? node50949 : node50946;
																assign node50946 = (inp[9]) ? 4'b1010 : 4'b1110;
																assign node50949 = (inp[9]) ? 4'b1110 : 4'b1010;
													assign node50952 = (inp[15]) ? node50964 : node50953;
														assign node50953 = (inp[0]) ? node50961 : node50954;
															assign node50954 = (inp[10]) ? node50958 : node50955;
																assign node50955 = (inp[9]) ? 4'b1110 : 4'b1010;
																assign node50958 = (inp[9]) ? 4'b1010 : 4'b1110;
															assign node50961 = (inp[9]) ? 4'b1100 : 4'b1000;
														assign node50964 = (inp[0]) ? 4'b1110 : node50965;
															assign node50965 = (inp[10]) ? node50967 : 4'b1100;
																assign node50967 = (inp[9]) ? 4'b1000 : 4'b1100;
												assign node50971 = (inp[15]) ? node50993 : node50972;
													assign node50972 = (inp[4]) ? node50984 : node50973;
														assign node50973 = (inp[0]) ? node50981 : node50974;
															assign node50974 = (inp[9]) ? node50978 : node50975;
																assign node50975 = (inp[10]) ? 4'b1010 : 4'b1110;
																assign node50978 = (inp[10]) ? 4'b1100 : 4'b1010;
															assign node50981 = (inp[9]) ? 4'b1000 : 4'b1100;
														assign node50984 = (inp[0]) ? node50988 : node50985;
															assign node50985 = (inp[9]) ? 4'b1100 : 4'b1010;
															assign node50988 = (inp[9]) ? node50990 : 4'b1110;
																assign node50990 = (inp[10]) ? 4'b1010 : 4'b1110;
													assign node50993 = (inp[9]) ? node51009 : node50994;
														assign node50994 = (inp[0]) ? node51002 : node50995;
															assign node50995 = (inp[10]) ? node50999 : node50996;
																assign node50996 = (inp[4]) ? 4'b1000 : 4'b1100;
																assign node50999 = (inp[4]) ? 4'b1110 : 4'b1000;
															assign node51002 = (inp[4]) ? node51006 : node51003;
																assign node51003 = (inp[10]) ? 4'b1010 : 4'b1110;
																assign node51006 = (inp[10]) ? 4'b1100 : 4'b1010;
														assign node51009 = (inp[4]) ? node51013 : node51010;
															assign node51010 = (inp[0]) ? 4'b1010 : 4'b1110;
															assign node51013 = (inp[0]) ? 4'b1000 : 4'b1010;
										assign node51016 = (inp[9]) ? node51080 : node51017;
											assign node51017 = (inp[15]) ? node51053 : node51018;
												assign node51018 = (inp[0]) ? node51036 : node51019;
													assign node51019 = (inp[3]) ? node51029 : node51020;
														assign node51020 = (inp[14]) ? 4'b1010 : node51021;
															assign node51021 = (inp[10]) ? node51025 : node51022;
																assign node51022 = (inp[4]) ? 4'b1010 : 4'b1110;
																assign node51025 = (inp[4]) ? 4'b1110 : 4'b1010;
														assign node51029 = (inp[10]) ? node51033 : node51030;
															assign node51030 = (inp[4]) ? 4'b1010 : 4'b1110;
															assign node51033 = (inp[4]) ? 4'b1100 : 4'b1010;
													assign node51036 = (inp[14]) ? node51046 : node51037;
														assign node51037 = (inp[4]) ? node51041 : node51038;
															assign node51038 = (inp[10]) ? 4'b1000 : 4'b1100;
															assign node51041 = (inp[10]) ? node51043 : 4'b1000;
																assign node51043 = (inp[3]) ? 4'b1110 : 4'b1100;
														assign node51046 = (inp[4]) ? node51050 : node51047;
															assign node51047 = (inp[10]) ? 4'b1000 : 4'b1100;
															assign node51050 = (inp[10]) ? 4'b1100 : 4'b1000;
												assign node51053 = (inp[0]) ? node51063 : node51054;
													assign node51054 = (inp[10]) ? node51058 : node51055;
														assign node51055 = (inp[4]) ? 4'b1000 : 4'b1100;
														assign node51058 = (inp[4]) ? node51060 : 4'b1000;
															assign node51060 = (inp[3]) ? 4'b1110 : 4'b1100;
													assign node51063 = (inp[14]) ? node51073 : node51064;
														assign node51064 = (inp[3]) ? node51066 : 4'b1110;
															assign node51066 = (inp[4]) ? node51070 : node51067;
																assign node51067 = (inp[10]) ? 4'b1010 : 4'b1110;
																assign node51070 = (inp[10]) ? 4'b1100 : 4'b1010;
														assign node51073 = (inp[4]) ? node51077 : node51074;
															assign node51074 = (inp[10]) ? 4'b1010 : 4'b1110;
															assign node51077 = (inp[10]) ? 4'b1110 : 4'b1010;
											assign node51080 = (inp[0]) ? node51114 : node51081;
												assign node51081 = (inp[3]) ? node51099 : node51082;
													assign node51082 = (inp[15]) ? node51090 : node51083;
														assign node51083 = (inp[14]) ? node51085 : 4'b1010;
															assign node51085 = (inp[4]) ? 4'b1110 : node51086;
																assign node51086 = (inp[10]) ? 4'b1110 : 4'b1010;
														assign node51090 = (inp[14]) ? 4'b1000 : node51091;
															assign node51091 = (inp[10]) ? node51095 : node51092;
																assign node51092 = (inp[4]) ? 4'b1100 : 4'b1000;
																assign node51095 = (inp[4]) ? 4'b1000 : 4'b1100;
													assign node51099 = (inp[15]) ? node51107 : node51100;
														assign node51100 = (inp[10]) ? node51104 : node51101;
															assign node51101 = (inp[4]) ? 4'b1100 : 4'b1010;
															assign node51104 = (inp[4]) ? 4'b1000 : 4'b1100;
														assign node51107 = (inp[4]) ? node51111 : node51108;
															assign node51108 = (inp[10]) ? 4'b1110 : 4'b1000;
															assign node51111 = (inp[10]) ? 4'b1010 : 4'b1110;
												assign node51114 = (inp[14]) ? node51136 : node51115;
													assign node51115 = (inp[4]) ? node51127 : node51116;
														assign node51116 = (inp[10]) ? node51120 : node51117;
															assign node51117 = (inp[15]) ? 4'b1010 : 4'b1000;
															assign node51120 = (inp[3]) ? node51124 : node51121;
																assign node51121 = (inp[15]) ? 4'b1110 : 4'b1100;
																assign node51124 = (inp[15]) ? 4'b1100 : 4'b1110;
														assign node51127 = (inp[10]) ? node51129 : 4'b1110;
															assign node51129 = (inp[3]) ? node51133 : node51130;
																assign node51130 = (inp[15]) ? 4'b1010 : 4'b1000;
																assign node51133 = (inp[15]) ? 4'b1000 : 4'b1010;
													assign node51136 = (inp[4]) ? node51140 : node51137;
														assign node51137 = (inp[10]) ? 4'b1110 : 4'b1010;
														assign node51140 = (inp[10]) ? 4'b1010 : node51141;
															assign node51141 = (inp[15]) ? node51145 : node51142;
																assign node51142 = (inp[3]) ? 4'b1110 : 4'b1100;
																assign node51145 = (inp[3]) ? 4'b1100 : 4'b1110;
							assign node51149 = (inp[7]) ? node51583 : node51150;
								assign node51150 = (inp[8]) ? node51364 : node51151;
									assign node51151 = (inp[2]) ? node51291 : node51152;
										assign node51152 = (inp[14]) ? node51222 : node51153;
											assign node51153 = (inp[3]) ? node51195 : node51154;
												assign node51154 = (inp[10]) ? node51180 : node51155;
													assign node51155 = (inp[0]) ? node51169 : node51156;
														assign node51156 = (inp[15]) ? node51162 : node51157;
															assign node51157 = (inp[9]) ? 4'b1011 : node51158;
																assign node51158 = (inp[4]) ? 4'b1111 : 4'b1011;
															assign node51162 = (inp[4]) ? node51166 : node51163;
																assign node51163 = (inp[9]) ? 4'b1101 : 4'b1001;
																assign node51166 = (inp[9]) ? 4'b1001 : 4'b1101;
														assign node51169 = (inp[15]) ? node51175 : node51170;
															assign node51170 = (inp[4]) ? node51172 : 4'b1101;
																assign node51172 = (inp[9]) ? 4'b1001 : 4'b1101;
															assign node51175 = (inp[9]) ? 4'b1111 : node51176;
																assign node51176 = (inp[4]) ? 4'b1111 : 4'b1011;
													assign node51180 = (inp[15]) ? node51188 : node51181;
														assign node51181 = (inp[0]) ? node51183 : 4'b1011;
															assign node51183 = (inp[4]) ? node51185 : 4'b1001;
																assign node51185 = (inp[9]) ? 4'b1001 : 4'b1101;
														assign node51188 = (inp[0]) ? 4'b1011 : node51189;
															assign node51189 = (inp[4]) ? node51191 : 4'b1101;
																assign node51191 = (inp[9]) ? 4'b1001 : 4'b1101;
												assign node51195 = (inp[0]) ? node51211 : node51196;
													assign node51196 = (inp[15]) ? node51204 : node51197;
														assign node51197 = (inp[4]) ? node51201 : node51198;
															assign node51198 = (inp[9]) ? 4'b1101 : 4'b1011;
															assign node51201 = (inp[9]) ? 4'b1001 : 4'b1101;
														assign node51204 = (inp[9]) ? node51208 : node51205;
															assign node51205 = (inp[4]) ? 4'b1111 : 4'b1001;
															assign node51208 = (inp[4]) ? 4'b1011 : 4'b1111;
													assign node51211 = (inp[15]) ? node51217 : node51212;
														assign node51212 = (inp[4]) ? node51214 : 4'b1111;
															assign node51214 = (inp[9]) ? 4'b1011 : 4'b1111;
														assign node51217 = (inp[9]) ? 4'b1101 : node51218;
															assign node51218 = (inp[4]) ? 4'b1101 : 4'b1011;
											assign node51222 = (inp[15]) ? node51256 : node51223;
												assign node51223 = (inp[0]) ? node51241 : node51224;
													assign node51224 = (inp[3]) ? node51232 : node51225;
														assign node51225 = (inp[9]) ? node51229 : node51226;
															assign node51226 = (inp[4]) ? 4'b1110 : 4'b1010;
															assign node51229 = (inp[4]) ? 4'b1010 : 4'b1110;
														assign node51232 = (inp[10]) ? node51236 : node51233;
															assign node51233 = (inp[4]) ? 4'b1100 : 4'b1010;
															assign node51236 = (inp[4]) ? node51238 : 4'b1100;
																assign node51238 = (inp[9]) ? 4'b1000 : 4'b1100;
													assign node51241 = (inp[3]) ? node51249 : node51242;
														assign node51242 = (inp[9]) ? node51246 : node51243;
															assign node51243 = (inp[4]) ? 4'b1100 : 4'b1000;
															assign node51246 = (inp[4]) ? 4'b1000 : 4'b1100;
														assign node51249 = (inp[9]) ? node51253 : node51250;
															assign node51250 = (inp[4]) ? 4'b1110 : 4'b1000;
															assign node51253 = (inp[4]) ? 4'b1010 : 4'b1110;
												assign node51256 = (inp[0]) ? node51272 : node51257;
													assign node51257 = (inp[3]) ? node51265 : node51258;
														assign node51258 = (inp[9]) ? node51262 : node51259;
															assign node51259 = (inp[4]) ? 4'b1100 : 4'b1000;
															assign node51262 = (inp[4]) ? 4'b1000 : 4'b1100;
														assign node51265 = (inp[9]) ? node51269 : node51266;
															assign node51266 = (inp[4]) ? 4'b1110 : 4'b1000;
															assign node51269 = (inp[4]) ? 4'b1010 : 4'b1110;
													assign node51272 = (inp[3]) ? node51280 : node51273;
														assign node51273 = (inp[9]) ? node51277 : node51274;
															assign node51274 = (inp[4]) ? 4'b1110 : 4'b1010;
															assign node51277 = (inp[4]) ? 4'b1010 : 4'b1110;
														assign node51280 = (inp[10]) ? node51286 : node51281;
															assign node51281 = (inp[4]) ? node51283 : 4'b1100;
																assign node51283 = (inp[9]) ? 4'b1000 : 4'b1100;
															assign node51286 = (inp[9]) ? node51288 : 4'b1010;
																assign node51288 = (inp[4]) ? 4'b1000 : 4'b1100;
										assign node51291 = (inp[3]) ? node51333 : node51292;
											assign node51292 = (inp[0]) ? node51318 : node51293;
												assign node51293 = (inp[15]) ? node51301 : node51294;
													assign node51294 = (inp[9]) ? node51298 : node51295;
														assign node51295 = (inp[4]) ? 4'b1110 : 4'b1010;
														assign node51298 = (inp[4]) ? 4'b1010 : 4'b1110;
													assign node51301 = (inp[10]) ? node51309 : node51302;
														assign node51302 = (inp[9]) ? node51306 : node51303;
															assign node51303 = (inp[4]) ? 4'b1100 : 4'b1000;
															assign node51306 = (inp[4]) ? 4'b1000 : 4'b1100;
														assign node51309 = (inp[14]) ? node51311 : 4'b1100;
															assign node51311 = (inp[9]) ? node51315 : node51312;
																assign node51312 = (inp[4]) ? 4'b1100 : 4'b1000;
																assign node51315 = (inp[4]) ? 4'b1000 : 4'b1100;
												assign node51318 = (inp[15]) ? node51326 : node51319;
													assign node51319 = (inp[4]) ? node51323 : node51320;
														assign node51320 = (inp[9]) ? 4'b1100 : 4'b1000;
														assign node51323 = (inp[9]) ? 4'b1000 : 4'b1100;
													assign node51326 = (inp[9]) ? node51330 : node51327;
														assign node51327 = (inp[4]) ? 4'b1110 : 4'b1010;
														assign node51330 = (inp[4]) ? 4'b1010 : 4'b1110;
											assign node51333 = (inp[0]) ? node51349 : node51334;
												assign node51334 = (inp[15]) ? node51342 : node51335;
													assign node51335 = (inp[4]) ? node51339 : node51336;
														assign node51336 = (inp[9]) ? 4'b1100 : 4'b1010;
														assign node51339 = (inp[9]) ? 4'b1000 : 4'b1100;
													assign node51342 = (inp[9]) ? node51346 : node51343;
														assign node51343 = (inp[4]) ? 4'b1110 : 4'b1000;
														assign node51346 = (inp[4]) ? 4'b1010 : 4'b1110;
												assign node51349 = (inp[15]) ? node51357 : node51350;
													assign node51350 = (inp[9]) ? node51354 : node51351;
														assign node51351 = (inp[4]) ? 4'b1110 : 4'b1000;
														assign node51354 = (inp[4]) ? 4'b1010 : 4'b1110;
													assign node51357 = (inp[9]) ? node51361 : node51358;
														assign node51358 = (inp[4]) ? 4'b1100 : 4'b1010;
														assign node51361 = (inp[4]) ? 4'b1000 : 4'b1100;
									assign node51364 = (inp[14]) ? node51470 : node51365;
										assign node51365 = (inp[2]) ? node51427 : node51366;
											assign node51366 = (inp[4]) ? node51396 : node51367;
												assign node51367 = (inp[9]) ? node51381 : node51368;
													assign node51368 = (inp[10]) ? node51370 : 4'b1000;
														assign node51370 = (inp[3]) ? node51376 : node51371;
															assign node51371 = (inp[15]) ? 4'b1000 : node51372;
																assign node51372 = (inp[0]) ? 4'b1000 : 4'b1010;
															assign node51376 = (inp[0]) ? node51378 : 4'b1010;
																assign node51378 = (inp[15]) ? 4'b1010 : 4'b1000;
													assign node51381 = (inp[15]) ? node51389 : node51382;
														assign node51382 = (inp[3]) ? node51386 : node51383;
															assign node51383 = (inp[0]) ? 4'b1100 : 4'b1110;
															assign node51386 = (inp[0]) ? 4'b1110 : 4'b1100;
														assign node51389 = (inp[10]) ? 4'b1110 : node51390;
															assign node51390 = (inp[3]) ? node51392 : 4'b1100;
																assign node51392 = (inp[0]) ? 4'b1100 : 4'b1110;
												assign node51396 = (inp[9]) ? node51410 : node51397;
													assign node51397 = (inp[3]) ? node51405 : node51398;
														assign node51398 = (inp[15]) ? node51402 : node51399;
															assign node51399 = (inp[0]) ? 4'b1100 : 4'b1110;
															assign node51402 = (inp[0]) ? 4'b1110 : 4'b1100;
														assign node51405 = (inp[10]) ? node51407 : 4'b1110;
															assign node51407 = (inp[0]) ? 4'b1100 : 4'b1110;
													assign node51410 = (inp[3]) ? node51420 : node51411;
														assign node51411 = (inp[10]) ? node51413 : 4'b1010;
															assign node51413 = (inp[15]) ? node51417 : node51414;
																assign node51414 = (inp[0]) ? 4'b1000 : 4'b1010;
																assign node51417 = (inp[0]) ? 4'b1010 : 4'b1000;
														assign node51420 = (inp[0]) ? node51424 : node51421;
															assign node51421 = (inp[15]) ? 4'b1010 : 4'b1000;
															assign node51424 = (inp[15]) ? 4'b1000 : 4'b1010;
											assign node51427 = (inp[9]) ? node51447 : node51428;
												assign node51428 = (inp[4]) ? node51436 : node51429;
													assign node51429 = (inp[0]) ? node51433 : node51430;
														assign node51430 = (inp[15]) ? 4'b1001 : 4'b1011;
														assign node51433 = (inp[15]) ? 4'b1011 : 4'b1001;
													assign node51436 = (inp[15]) ? 4'b1111 : node51437;
														assign node51437 = (inp[10]) ? node51439 : 4'b1101;
															assign node51439 = (inp[0]) ? node51443 : node51440;
																assign node51440 = (inp[3]) ? 4'b1101 : 4'b1111;
																assign node51443 = (inp[3]) ? 4'b1111 : 4'b1101;
												assign node51447 = (inp[4]) ? node51459 : node51448;
													assign node51448 = (inp[15]) ? node51450 : 4'b1111;
														assign node51450 = (inp[10]) ? node51456 : node51451;
															assign node51451 = (inp[0]) ? node51453 : 4'b1101;
																assign node51453 = (inp[3]) ? 4'b1101 : 4'b1111;
															assign node51456 = (inp[0]) ? 4'b1101 : 4'b1111;
													assign node51459 = (inp[10]) ? node51465 : node51460;
														assign node51460 = (inp[0]) ? node51462 : 4'b1011;
															assign node51462 = (inp[3]) ? 4'b1011 : 4'b1001;
														assign node51465 = (inp[15]) ? 4'b1001 : node51466;
															assign node51466 = (inp[0]) ? 4'b1011 : 4'b1001;
										assign node51470 = (inp[10]) ? node51528 : node51471;
											assign node51471 = (inp[15]) ? node51493 : node51472;
												assign node51472 = (inp[4]) ? node51484 : node51473;
													assign node51473 = (inp[9]) ? node51477 : node51474;
														assign node51474 = (inp[0]) ? 4'b1001 : 4'b1011;
														assign node51477 = (inp[3]) ? node51481 : node51478;
															assign node51478 = (inp[0]) ? 4'b1101 : 4'b1111;
															assign node51481 = (inp[0]) ? 4'b1111 : 4'b1101;
													assign node51484 = (inp[9]) ? node51486 : 4'b1111;
														assign node51486 = (inp[0]) ? node51490 : node51487;
															assign node51487 = (inp[3]) ? 4'b1001 : 4'b1011;
															assign node51490 = (inp[3]) ? 4'b1011 : 4'b1001;
												assign node51493 = (inp[0]) ? node51515 : node51494;
													assign node51494 = (inp[3]) ? node51508 : node51495;
														assign node51495 = (inp[2]) ? node51501 : node51496;
															assign node51496 = (inp[4]) ? node51498 : 4'b1001;
																assign node51498 = (inp[9]) ? 4'b1001 : 4'b1101;
															assign node51501 = (inp[4]) ? node51505 : node51502;
																assign node51502 = (inp[9]) ? 4'b1101 : 4'b1001;
																assign node51505 = (inp[9]) ? 4'b1001 : 4'b1101;
														assign node51508 = (inp[9]) ? node51512 : node51509;
															assign node51509 = (inp[4]) ? 4'b1111 : 4'b1001;
															assign node51512 = (inp[4]) ? 4'b1011 : 4'b1111;
													assign node51515 = (inp[3]) ? node51521 : node51516;
														assign node51516 = (inp[9]) ? 4'b1011 : node51517;
															assign node51517 = (inp[4]) ? 4'b1111 : 4'b1011;
														assign node51521 = (inp[4]) ? node51525 : node51522;
															assign node51522 = (inp[9]) ? 4'b1101 : 4'b1011;
															assign node51525 = (inp[9]) ? 4'b1001 : 4'b1101;
											assign node51528 = (inp[3]) ? node51552 : node51529;
												assign node51529 = (inp[4]) ? node51539 : node51530;
													assign node51530 = (inp[9]) ? node51532 : 4'b1001;
														assign node51532 = (inp[15]) ? node51536 : node51533;
															assign node51533 = (inp[0]) ? 4'b1101 : 4'b1111;
															assign node51536 = (inp[0]) ? 4'b1111 : 4'b1101;
													assign node51539 = (inp[9]) ? node51547 : node51540;
														assign node51540 = (inp[0]) ? node51544 : node51541;
															assign node51541 = (inp[15]) ? 4'b1101 : 4'b1111;
															assign node51544 = (inp[15]) ? 4'b1111 : 4'b1101;
														assign node51547 = (inp[2]) ? node51549 : 4'b1001;
															assign node51549 = (inp[15]) ? 4'b1011 : 4'b1001;
												assign node51552 = (inp[15]) ? node51570 : node51553;
													assign node51553 = (inp[0]) ? node51559 : node51554;
														assign node51554 = (inp[4]) ? node51556 : 4'b1011;
															assign node51556 = (inp[9]) ? 4'b1001 : 4'b1101;
														assign node51559 = (inp[2]) ? node51565 : node51560;
															assign node51560 = (inp[9]) ? node51562 : 4'b1111;
																assign node51562 = (inp[4]) ? 4'b1011 : 4'b1111;
															assign node51565 = (inp[4]) ? node51567 : 4'b1001;
																assign node51567 = (inp[9]) ? 4'b1011 : 4'b1111;
													assign node51570 = (inp[0]) ? node51576 : node51571;
														assign node51571 = (inp[9]) ? node51573 : 4'b1001;
															assign node51573 = (inp[4]) ? 4'b1011 : 4'b1111;
														assign node51576 = (inp[9]) ? node51580 : node51577;
															assign node51577 = (inp[4]) ? 4'b1101 : 4'b1011;
															assign node51580 = (inp[4]) ? 4'b1001 : 4'b1101;
								assign node51583 = (inp[8]) ? node51859 : node51584;
									assign node51584 = (inp[14]) ? node51730 : node51585;
										assign node51585 = (inp[2]) ? node51647 : node51586;
											assign node51586 = (inp[3]) ? node51620 : node51587;
												assign node51587 = (inp[0]) ? node51605 : node51588;
													assign node51588 = (inp[15]) ? 4'b1000 : node51589;
														assign node51589 = (inp[10]) ? node51597 : node51590;
															assign node51590 = (inp[4]) ? node51594 : node51591;
																assign node51591 = (inp[9]) ? 4'b1110 : 4'b1010;
																assign node51594 = (inp[9]) ? 4'b1010 : 4'b1110;
															assign node51597 = (inp[9]) ? node51601 : node51598;
																assign node51598 = (inp[4]) ? 4'b1110 : 4'b1010;
																assign node51601 = (inp[4]) ? 4'b1010 : 4'b1110;
													assign node51605 = (inp[15]) ? node51613 : node51606;
														assign node51606 = (inp[4]) ? node51610 : node51607;
															assign node51607 = (inp[9]) ? 4'b1100 : 4'b1000;
															assign node51610 = (inp[9]) ? 4'b1000 : 4'b1100;
														assign node51613 = (inp[9]) ? node51617 : node51614;
															assign node51614 = (inp[4]) ? 4'b1110 : 4'b1010;
															assign node51617 = (inp[4]) ? 4'b1010 : 4'b1110;
												assign node51620 = (inp[15]) ? node51630 : node51621;
													assign node51621 = (inp[0]) ? node51627 : node51622;
														assign node51622 = (inp[9]) ? node51624 : 4'b1100;
															assign node51624 = (inp[4]) ? 4'b1000 : 4'b1100;
														assign node51627 = (inp[4]) ? 4'b1110 : 4'b1000;
													assign node51630 = (inp[0]) ? node51640 : node51631;
														assign node51631 = (inp[10]) ? node51637 : node51632;
															assign node51632 = (inp[9]) ? node51634 : 4'b1110;
																assign node51634 = (inp[4]) ? 4'b1010 : 4'b1110;
															assign node51637 = (inp[9]) ? 4'b1110 : 4'b1000;
														assign node51640 = (inp[9]) ? node51644 : node51641;
															assign node51641 = (inp[4]) ? 4'b1100 : 4'b1010;
															assign node51644 = (inp[4]) ? 4'b1000 : 4'b1100;
											assign node51647 = (inp[4]) ? node51693 : node51648;
												assign node51648 = (inp[9]) ? node51668 : node51649;
													assign node51649 = (inp[3]) ? node51655 : node51650;
														assign node51650 = (inp[0]) ? node51652 : 4'b1011;
															assign node51652 = (inp[15]) ? 4'b1011 : 4'b1001;
														assign node51655 = (inp[10]) ? node51663 : node51656;
															assign node51656 = (inp[0]) ? node51660 : node51657;
																assign node51657 = (inp[15]) ? 4'b1001 : 4'b1011;
																assign node51660 = (inp[15]) ? 4'b1011 : 4'b1001;
															assign node51663 = (inp[15]) ? node51665 : 4'b1001;
																assign node51665 = (inp[0]) ? 4'b1011 : 4'b1001;
													assign node51668 = (inp[15]) ? node51680 : node51669;
														assign node51669 = (inp[10]) ? node51675 : node51670;
															assign node51670 = (inp[3]) ? 4'b1111 : node51671;
																assign node51671 = (inp[0]) ? 4'b1101 : 4'b1111;
															assign node51675 = (inp[0]) ? 4'b1111 : node51676;
																assign node51676 = (inp[3]) ? 4'b1101 : 4'b1111;
														assign node51680 = (inp[10]) ? node51686 : node51681;
															assign node51681 = (inp[0]) ? 4'b1101 : node51682;
																assign node51682 = (inp[3]) ? 4'b1111 : 4'b1101;
															assign node51686 = (inp[3]) ? node51690 : node51687;
																assign node51687 = (inp[0]) ? 4'b1111 : 4'b1101;
																assign node51690 = (inp[0]) ? 4'b1101 : 4'b1111;
												assign node51693 = (inp[9]) ? node51711 : node51694;
													assign node51694 = (inp[15]) ? node51702 : node51695;
														assign node51695 = (inp[0]) ? node51699 : node51696;
															assign node51696 = (inp[3]) ? 4'b1101 : 4'b1111;
															assign node51699 = (inp[3]) ? 4'b1111 : 4'b1101;
														assign node51702 = (inp[10]) ? 4'b1101 : node51703;
															assign node51703 = (inp[3]) ? node51707 : node51704;
																assign node51704 = (inp[0]) ? 4'b1111 : 4'b1101;
																assign node51707 = (inp[0]) ? 4'b1101 : 4'b1111;
													assign node51711 = (inp[3]) ? node51723 : node51712;
														assign node51712 = (inp[10]) ? node51718 : node51713;
															assign node51713 = (inp[0]) ? 4'b1011 : node51714;
																assign node51714 = (inp[15]) ? 4'b1001 : 4'b1011;
															assign node51718 = (inp[0]) ? 4'b1001 : node51719;
																assign node51719 = (inp[15]) ? 4'b1001 : 4'b1011;
														assign node51723 = (inp[15]) ? node51727 : node51724;
															assign node51724 = (inp[0]) ? 4'b1011 : 4'b1001;
															assign node51727 = (inp[0]) ? 4'b1001 : 4'b1011;
										assign node51730 = (inp[3]) ? node51768 : node51731;
											assign node51731 = (inp[4]) ? node51753 : node51732;
												assign node51732 = (inp[9]) ? node51746 : node51733;
													assign node51733 = (inp[10]) ? node51741 : node51734;
														assign node51734 = (inp[0]) ? node51738 : node51735;
															assign node51735 = (inp[15]) ? 4'b1001 : 4'b1011;
															assign node51738 = (inp[15]) ? 4'b1011 : 4'b1001;
														assign node51741 = (inp[15]) ? node51743 : 4'b1011;
															assign node51743 = (inp[0]) ? 4'b1011 : 4'b1001;
													assign node51746 = (inp[0]) ? node51750 : node51747;
														assign node51747 = (inp[15]) ? 4'b1101 : 4'b1111;
														assign node51750 = (inp[15]) ? 4'b1111 : 4'b1101;
												assign node51753 = (inp[9]) ? node51761 : node51754;
													assign node51754 = (inp[15]) ? node51758 : node51755;
														assign node51755 = (inp[0]) ? 4'b1101 : 4'b1111;
														assign node51758 = (inp[0]) ? 4'b1111 : 4'b1101;
													assign node51761 = (inp[15]) ? node51765 : node51762;
														assign node51762 = (inp[0]) ? 4'b1001 : 4'b1011;
														assign node51765 = (inp[0]) ? 4'b1011 : 4'b1001;
											assign node51768 = (inp[2]) ? node51814 : node51769;
												assign node51769 = (inp[10]) ? node51789 : node51770;
													assign node51770 = (inp[0]) ? node51780 : node51771;
														assign node51771 = (inp[4]) ? node51775 : node51772;
															assign node51772 = (inp[15]) ? 4'b1001 : 4'b1011;
															assign node51775 = (inp[15]) ? 4'b1011 : node51776;
																assign node51776 = (inp[9]) ? 4'b1001 : 4'b1101;
														assign node51780 = (inp[15]) ? node51784 : node51781;
															assign node51781 = (inp[9]) ? 4'b1111 : 4'b1001;
															assign node51784 = (inp[9]) ? node51786 : 4'b1101;
																assign node51786 = (inp[4]) ? 4'b1001 : 4'b1101;
													assign node51789 = (inp[9]) ? node51803 : node51790;
														assign node51790 = (inp[4]) ? node51796 : node51791;
															assign node51791 = (inp[15]) ? 4'b1011 : node51792;
																assign node51792 = (inp[0]) ? 4'b1001 : 4'b1011;
															assign node51796 = (inp[0]) ? node51800 : node51797;
																assign node51797 = (inp[15]) ? 4'b1111 : 4'b1101;
																assign node51800 = (inp[15]) ? 4'b1101 : 4'b1111;
														assign node51803 = (inp[4]) ? node51809 : node51804;
															assign node51804 = (inp[15]) ? 4'b1101 : node51805;
																assign node51805 = (inp[0]) ? 4'b1111 : 4'b1101;
															assign node51809 = (inp[0]) ? node51811 : 4'b1001;
																assign node51811 = (inp[15]) ? 4'b1001 : 4'b1011;
												assign node51814 = (inp[10]) ? node51842 : node51815;
													assign node51815 = (inp[15]) ? node51831 : node51816;
														assign node51816 = (inp[0]) ? node51824 : node51817;
															assign node51817 = (inp[4]) ? node51821 : node51818;
																assign node51818 = (inp[9]) ? 4'b1101 : 4'b1011;
																assign node51821 = (inp[9]) ? 4'b1001 : 4'b1101;
															assign node51824 = (inp[4]) ? node51828 : node51825;
																assign node51825 = (inp[9]) ? 4'b1111 : 4'b1001;
																assign node51828 = (inp[9]) ? 4'b1011 : 4'b1111;
														assign node51831 = (inp[0]) ? node51837 : node51832;
															assign node51832 = (inp[4]) ? node51834 : 4'b1111;
																assign node51834 = (inp[9]) ? 4'b1011 : 4'b1111;
															assign node51837 = (inp[9]) ? node51839 : 4'b1011;
																assign node51839 = (inp[4]) ? 4'b1001 : 4'b1101;
													assign node51842 = (inp[4]) ? node51850 : node51843;
														assign node51843 = (inp[9]) ? 4'b1101 : node51844;
															assign node51844 = (inp[15]) ? 4'b1001 : node51845;
																assign node51845 = (inp[0]) ? 4'b1001 : 4'b1011;
														assign node51850 = (inp[9]) ? node51856 : node51851;
															assign node51851 = (inp[15]) ? 4'b1111 : node51852;
																assign node51852 = (inp[0]) ? 4'b1111 : 4'b1101;
															assign node51856 = (inp[0]) ? 4'b1011 : 4'b1001;
									assign node51859 = (inp[14]) ? node51973 : node51860;
										assign node51860 = (inp[2]) ? node51918 : node51861;
											assign node51861 = (inp[0]) ? node51891 : node51862;
												assign node51862 = (inp[3]) ? node51880 : node51863;
													assign node51863 = (inp[15]) ? node51873 : node51864;
														assign node51864 = (inp[10]) ? 4'b1011 : node51865;
															assign node51865 = (inp[4]) ? node51869 : node51866;
																assign node51866 = (inp[9]) ? 4'b1111 : 4'b1011;
																assign node51869 = (inp[9]) ? 4'b1011 : 4'b1111;
														assign node51873 = (inp[10]) ? 4'b1101 : node51874;
															assign node51874 = (inp[4]) ? 4'b1001 : node51875;
																assign node51875 = (inp[9]) ? 4'b1101 : 4'b1001;
													assign node51880 = (inp[15]) ? node51886 : node51881;
														assign node51881 = (inp[9]) ? 4'b1101 : node51882;
															assign node51882 = (inp[4]) ? 4'b1101 : 4'b1011;
														assign node51886 = (inp[9]) ? node51888 : 4'b1111;
															assign node51888 = (inp[4]) ? 4'b1011 : 4'b1111;
												assign node51891 = (inp[15]) ? node51905 : node51892;
													assign node51892 = (inp[3]) ? node51900 : node51893;
														assign node51893 = (inp[9]) ? node51897 : node51894;
															assign node51894 = (inp[4]) ? 4'b1101 : 4'b1001;
															assign node51897 = (inp[4]) ? 4'b1001 : 4'b1101;
														assign node51900 = (inp[9]) ? node51902 : 4'b1111;
															assign node51902 = (inp[4]) ? 4'b1011 : 4'b1111;
													assign node51905 = (inp[3]) ? node51911 : node51906;
														assign node51906 = (inp[9]) ? node51908 : 4'b1111;
															assign node51908 = (inp[4]) ? 4'b1011 : 4'b1111;
														assign node51911 = (inp[9]) ? node51915 : node51912;
															assign node51912 = (inp[4]) ? 4'b1101 : 4'b1011;
															assign node51915 = (inp[4]) ? 4'b1001 : 4'b1101;
											assign node51918 = (inp[4]) ? node51940 : node51919;
												assign node51919 = (inp[9]) ? node51927 : node51920;
													assign node51920 = (inp[0]) ? node51924 : node51921;
														assign node51921 = (inp[15]) ? 4'b1000 : 4'b1010;
														assign node51924 = (inp[15]) ? 4'b1010 : 4'b1000;
													assign node51927 = (inp[0]) ? node51935 : node51928;
														assign node51928 = (inp[3]) ? node51932 : node51929;
															assign node51929 = (inp[15]) ? 4'b1100 : 4'b1110;
															assign node51932 = (inp[15]) ? 4'b1110 : 4'b1100;
														assign node51935 = (inp[15]) ? node51937 : 4'b1110;
															assign node51937 = (inp[3]) ? 4'b1100 : 4'b1110;
												assign node51940 = (inp[9]) ? node51958 : node51941;
													assign node51941 = (inp[3]) ? node51951 : node51942;
														assign node51942 = (inp[10]) ? 4'b1100 : node51943;
															assign node51943 = (inp[15]) ? node51947 : node51944;
																assign node51944 = (inp[0]) ? 4'b1100 : 4'b1110;
																assign node51947 = (inp[0]) ? 4'b1110 : 4'b1100;
														assign node51951 = (inp[10]) ? 4'b1110 : node51952;
															assign node51952 = (inp[0]) ? 4'b1100 : node51953;
																assign node51953 = (inp[15]) ? 4'b1110 : 4'b1100;
													assign node51958 = (inp[10]) ? node51966 : node51959;
														assign node51959 = (inp[3]) ? node51961 : 4'b1010;
															assign node51961 = (inp[0]) ? 4'b1000 : node51962;
																assign node51962 = (inp[15]) ? 4'b1010 : 4'b1000;
														assign node51966 = (inp[0]) ? 4'b1000 : node51967;
															assign node51967 = (inp[15]) ? 4'b1000 : node51968;
																assign node51968 = (inp[3]) ? 4'b1000 : 4'b1010;
										assign node51973 = (inp[0]) ? node52011 : node51974;
											assign node51974 = (inp[15]) ? node51990 : node51975;
												assign node51975 = (inp[3]) ? node51983 : node51976;
													assign node51976 = (inp[4]) ? node51980 : node51977;
														assign node51977 = (inp[9]) ? 4'b1110 : 4'b1010;
														assign node51980 = (inp[9]) ? 4'b1010 : 4'b1110;
													assign node51983 = (inp[4]) ? node51987 : node51984;
														assign node51984 = (inp[9]) ? 4'b1100 : 4'b1010;
														assign node51987 = (inp[9]) ? 4'b1000 : 4'b1100;
												assign node51990 = (inp[3]) ? node52004 : node51991;
													assign node51991 = (inp[10]) ? node51999 : node51992;
														assign node51992 = (inp[4]) ? node51996 : node51993;
															assign node51993 = (inp[9]) ? 4'b1100 : 4'b1000;
															assign node51996 = (inp[9]) ? 4'b1000 : 4'b1100;
														assign node51999 = (inp[9]) ? node52001 : 4'b1100;
															assign node52001 = (inp[4]) ? 4'b1000 : 4'b1100;
													assign node52004 = (inp[9]) ? node52008 : node52005;
														assign node52005 = (inp[4]) ? 4'b1110 : 4'b1000;
														assign node52008 = (inp[4]) ? 4'b1010 : 4'b1110;
											assign node52011 = (inp[15]) ? node52049 : node52012;
												assign node52012 = (inp[3]) ? node52042 : node52013;
													assign node52013 = (inp[10]) ? node52027 : node52014;
														assign node52014 = (inp[2]) ? node52020 : node52015;
															assign node52015 = (inp[4]) ? 4'b1100 : node52016;
																assign node52016 = (inp[9]) ? 4'b1100 : 4'b1000;
															assign node52020 = (inp[4]) ? node52024 : node52021;
																assign node52021 = (inp[9]) ? 4'b1100 : 4'b1000;
																assign node52024 = (inp[9]) ? 4'b1000 : 4'b1100;
														assign node52027 = (inp[2]) ? node52035 : node52028;
															assign node52028 = (inp[4]) ? node52032 : node52029;
																assign node52029 = (inp[9]) ? 4'b1100 : 4'b1000;
																assign node52032 = (inp[9]) ? 4'b1000 : 4'b1100;
															assign node52035 = (inp[4]) ? node52039 : node52036;
																assign node52036 = (inp[9]) ? 4'b1100 : 4'b1000;
																assign node52039 = (inp[9]) ? 4'b1000 : 4'b1100;
													assign node52042 = (inp[4]) ? node52046 : node52043;
														assign node52043 = (inp[9]) ? 4'b1110 : 4'b1000;
														assign node52046 = (inp[9]) ? 4'b1010 : 4'b1110;
												assign node52049 = (inp[3]) ? node52063 : node52050;
													assign node52050 = (inp[2]) ? node52058 : node52051;
														assign node52051 = (inp[4]) ? node52055 : node52052;
															assign node52052 = (inp[9]) ? 4'b1110 : 4'b1010;
															assign node52055 = (inp[9]) ? 4'b1010 : 4'b1110;
														assign node52058 = (inp[4]) ? node52060 : 4'b1110;
															assign node52060 = (inp[9]) ? 4'b1010 : 4'b1110;
													assign node52063 = (inp[4]) ? node52067 : node52064;
														assign node52064 = (inp[9]) ? 4'b1100 : 4'b1010;
														assign node52067 = (inp[9]) ? 4'b1000 : 4'b1100;
						assign node52070 = (inp[7]) ? node53068 : node52071;
							assign node52071 = (inp[8]) ? node52581 : node52072;
								assign node52072 = (inp[14]) ? node52380 : node52073;
									assign node52073 = (inp[2]) ? node52245 : node52074;
										assign node52074 = (inp[10]) ? node52170 : node52075;
											assign node52075 = (inp[15]) ? node52121 : node52076;
												assign node52076 = (inp[0]) ? node52096 : node52077;
													assign node52077 = (inp[3]) ? node52087 : node52078;
														assign node52078 = (inp[12]) ? node52084 : node52079;
															assign node52079 = (inp[9]) ? 4'b1011 : node52080;
																assign node52080 = (inp[4]) ? 4'b1011 : 4'b1111;
															assign node52084 = (inp[4]) ? 4'b1001 : 4'b1101;
														assign node52087 = (inp[9]) ? node52089 : 4'b1001;
															assign node52089 = (inp[12]) ? node52093 : node52090;
																assign node52090 = (inp[4]) ? 4'b1101 : 4'b1001;
																assign node52093 = (inp[4]) ? 4'b1001 : 4'b1101;
													assign node52096 = (inp[3]) ? node52108 : node52097;
														assign node52097 = (inp[12]) ? node52103 : node52098;
															assign node52098 = (inp[9]) ? 4'b1001 : node52099;
																assign node52099 = (inp[4]) ? 4'b1001 : 4'b1101;
															assign node52103 = (inp[4]) ? node52105 : 4'b1001;
																assign node52105 = (inp[9]) ? 4'b1011 : 4'b1111;
														assign node52108 = (inp[12]) ? node52114 : node52109;
															assign node52109 = (inp[4]) ? 4'b1111 : node52110;
																assign node52110 = (inp[9]) ? 4'b1011 : 4'b1111;
															assign node52114 = (inp[4]) ? node52118 : node52115;
																assign node52115 = (inp[9]) ? 4'b1111 : 4'b1011;
																assign node52118 = (inp[9]) ? 4'b1011 : 4'b1111;
												assign node52121 = (inp[0]) ? node52145 : node52122;
													assign node52122 = (inp[3]) ? node52132 : node52123;
														assign node52123 = (inp[12]) ? node52127 : node52124;
															assign node52124 = (inp[4]) ? 4'b1001 : 4'b1101;
															assign node52127 = (inp[4]) ? node52129 : 4'b1111;
																assign node52129 = (inp[9]) ? 4'b1011 : 4'b1111;
														assign node52132 = (inp[12]) ? node52140 : node52133;
															assign node52133 = (inp[4]) ? node52137 : node52134;
																assign node52134 = (inp[9]) ? 4'b1011 : 4'b1111;
																assign node52137 = (inp[9]) ? 4'b1111 : 4'b1011;
															assign node52140 = (inp[9]) ? node52142 : 4'b1111;
																assign node52142 = (inp[4]) ? 4'b1011 : 4'b1111;
													assign node52145 = (inp[3]) ? node52161 : node52146;
														assign node52146 = (inp[9]) ? node52154 : node52147;
															assign node52147 = (inp[12]) ? node52151 : node52148;
																assign node52148 = (inp[4]) ? 4'b1011 : 4'b1111;
																assign node52151 = (inp[4]) ? 4'b1101 : 4'b1011;
															assign node52154 = (inp[12]) ? node52158 : node52155;
																assign node52155 = (inp[4]) ? 4'b1101 : 4'b1011;
																assign node52158 = (inp[4]) ? 4'b1001 : 4'b1101;
														assign node52161 = (inp[12]) ? 4'b1001 : node52162;
															assign node52162 = (inp[4]) ? node52166 : node52163;
																assign node52163 = (inp[9]) ? 4'b1001 : 4'b1101;
																assign node52166 = (inp[9]) ? 4'b1101 : 4'b1001;
											assign node52170 = (inp[12]) ? node52208 : node52171;
												assign node52171 = (inp[9]) ? node52195 : node52172;
													assign node52172 = (inp[4]) ? node52182 : node52173;
														assign node52173 = (inp[0]) ? 4'b1001 : node52174;
															assign node52174 = (inp[3]) ? node52178 : node52175;
																assign node52175 = (inp[15]) ? 4'b1001 : 4'b1011;
																assign node52178 = (inp[15]) ? 4'b1011 : 4'b1001;
														assign node52182 = (inp[3]) ? node52188 : node52183;
															assign node52183 = (inp[0]) ? 4'b1101 : node52184;
																assign node52184 = (inp[15]) ? 4'b1111 : 4'b1101;
															assign node52188 = (inp[0]) ? node52192 : node52189;
																assign node52189 = (inp[15]) ? 4'b1111 : 4'b1101;
																assign node52192 = (inp[15]) ? 4'b1101 : 4'b1111;
													assign node52195 = (inp[4]) ? node52201 : node52196;
														assign node52196 = (inp[15]) ? 4'b1111 : node52197;
															assign node52197 = (inp[0]) ? 4'b1111 : 4'b1101;
														assign node52201 = (inp[15]) ? node52205 : node52202;
															assign node52202 = (inp[0]) ? 4'b1011 : 4'b1001;
															assign node52205 = (inp[0]) ? 4'b1001 : 4'b1011;
												assign node52208 = (inp[0]) ? node52228 : node52209;
													assign node52209 = (inp[15]) ? node52219 : node52210;
														assign node52210 = (inp[4]) ? node52216 : node52211;
															assign node52211 = (inp[9]) ? 4'b1101 : node52212;
																assign node52212 = (inp[3]) ? 4'b1001 : 4'b1011;
															assign node52216 = (inp[9]) ? 4'b1001 : 4'b1101;
														assign node52219 = (inp[3]) ? node52223 : node52220;
															assign node52220 = (inp[4]) ? 4'b1111 : 4'b1001;
															assign node52223 = (inp[9]) ? node52225 : 4'b1011;
																assign node52225 = (inp[4]) ? 4'b1011 : 4'b1111;
													assign node52228 = (inp[15]) ? node52238 : node52229;
														assign node52229 = (inp[9]) ? node52235 : node52230;
															assign node52230 = (inp[4]) ? 4'b1111 : node52231;
																assign node52231 = (inp[3]) ? 4'b1011 : 4'b1001;
															assign node52235 = (inp[4]) ? 4'b1011 : 4'b1111;
														assign node52238 = (inp[4]) ? node52242 : node52239;
															assign node52239 = (inp[9]) ? 4'b1101 : 4'b1011;
															assign node52242 = (inp[9]) ? 4'b1001 : 4'b1101;
										assign node52245 = (inp[15]) ? node52315 : node52246;
											assign node52246 = (inp[0]) ? node52278 : node52247;
												assign node52247 = (inp[3]) ? node52263 : node52248;
													assign node52248 = (inp[4]) ? node52256 : node52249;
														assign node52249 = (inp[9]) ? node52253 : node52250;
															assign node52250 = (inp[12]) ? 4'b1010 : 4'b1110;
															assign node52253 = (inp[12]) ? 4'b1100 : 4'b1010;
														assign node52256 = (inp[9]) ? 4'b1000 : node52257;
															assign node52257 = (inp[10]) ? 4'b1100 : node52258;
																assign node52258 = (inp[12]) ? 4'b1100 : 4'b1010;
													assign node52263 = (inp[10]) ? node52271 : node52264;
														assign node52264 = (inp[4]) ? node52266 : 4'b1000;
															assign node52266 = (inp[12]) ? node52268 : 4'b1000;
																assign node52268 = (inp[9]) ? 4'b1000 : 4'b1100;
														assign node52271 = (inp[9]) ? node52275 : node52272;
															assign node52272 = (inp[4]) ? 4'b1100 : 4'b1000;
															assign node52275 = (inp[4]) ? 4'b1000 : 4'b1100;
												assign node52278 = (inp[3]) ? node52300 : node52279;
													assign node52279 = (inp[12]) ? node52295 : node52280;
														assign node52280 = (inp[9]) ? node52288 : node52281;
															assign node52281 = (inp[10]) ? node52285 : node52282;
																assign node52282 = (inp[4]) ? 4'b1000 : 4'b1100;
																assign node52285 = (inp[4]) ? 4'b1110 : 4'b1000;
															assign node52288 = (inp[10]) ? node52292 : node52289;
																assign node52289 = (inp[4]) ? 4'b1110 : 4'b1000;
																assign node52292 = (inp[4]) ? 4'b1010 : 4'b1110;
														assign node52295 = (inp[4]) ? node52297 : 4'b1110;
															assign node52297 = (inp[9]) ? 4'b1010 : 4'b1110;
													assign node52300 = (inp[10]) ? node52310 : node52301;
														assign node52301 = (inp[9]) ? node52303 : 4'b1110;
															assign node52303 = (inp[12]) ? node52307 : node52304;
																assign node52304 = (inp[4]) ? 4'b1110 : 4'b1010;
																assign node52307 = (inp[4]) ? 4'b1010 : 4'b1110;
														assign node52310 = (inp[4]) ? 4'b1010 : node52311;
															assign node52311 = (inp[9]) ? 4'b1110 : 4'b1010;
											assign node52315 = (inp[0]) ? node52347 : node52316;
												assign node52316 = (inp[3]) ? node52332 : node52317;
													assign node52317 = (inp[4]) ? node52323 : node52318;
														assign node52318 = (inp[9]) ? node52320 : 4'b1000;
															assign node52320 = (inp[10]) ? 4'b1110 : 4'b1000;
														assign node52323 = (inp[12]) ? node52329 : node52324;
															assign node52324 = (inp[9]) ? node52326 : 4'b1000;
																assign node52326 = (inp[10]) ? 4'b1010 : 4'b1110;
															assign node52329 = (inp[9]) ? 4'b1010 : 4'b1110;
													assign node52332 = (inp[9]) ? node52338 : node52333;
														assign node52333 = (inp[4]) ? 4'b1110 : node52334;
															assign node52334 = (inp[12]) ? 4'b1010 : 4'b1110;
														assign node52338 = (inp[4]) ? node52342 : node52339;
															assign node52339 = (inp[10]) ? 4'b1110 : 4'b1010;
															assign node52342 = (inp[10]) ? 4'b1010 : node52343;
																assign node52343 = (inp[12]) ? 4'b1010 : 4'b1110;
												assign node52347 = (inp[3]) ? node52367 : node52348;
													assign node52348 = (inp[12]) ? node52362 : node52349;
														assign node52349 = (inp[10]) ? node52357 : node52350;
															assign node52350 = (inp[4]) ? node52354 : node52351;
																assign node52351 = (inp[9]) ? 4'b1010 : 4'b1110;
																assign node52354 = (inp[9]) ? 4'b1100 : 4'b1010;
															assign node52357 = (inp[4]) ? 4'b1100 : node52358;
																assign node52358 = (inp[9]) ? 4'b1100 : 4'b1010;
														assign node52362 = (inp[9]) ? node52364 : 4'b1100;
															assign node52364 = (inp[4]) ? 4'b1000 : 4'b1100;
													assign node52367 = (inp[9]) ? node52375 : node52368;
														assign node52368 = (inp[4]) ? node52370 : 4'b1000;
															assign node52370 = (inp[12]) ? 4'b1100 : node52371;
																assign node52371 = (inp[10]) ? 4'b1100 : 4'b1000;
														assign node52375 = (inp[4]) ? node52377 : 4'b1100;
															assign node52377 = (inp[10]) ? 4'b1000 : 4'b1100;
									assign node52380 = (inp[10]) ? node52516 : node52381;
										assign node52381 = (inp[12]) ? node52451 : node52382;
											assign node52382 = (inp[2]) ? node52420 : node52383;
												assign node52383 = (inp[9]) ? node52401 : node52384;
													assign node52384 = (inp[4]) ? node52394 : node52385;
														assign node52385 = (inp[0]) ? node52387 : 4'b1100;
															assign node52387 = (inp[15]) ? node52391 : node52388;
																assign node52388 = (inp[3]) ? 4'b1110 : 4'b1100;
																assign node52391 = (inp[3]) ? 4'b1100 : 4'b1110;
														assign node52394 = (inp[3]) ? node52396 : 4'b1000;
															assign node52396 = (inp[15]) ? 4'b1010 : node52397;
																assign node52397 = (inp[0]) ? 4'b1010 : 4'b1000;
													assign node52401 = (inp[4]) ? node52411 : node52402;
														assign node52402 = (inp[3]) ? 4'b1010 : node52403;
															assign node52403 = (inp[15]) ? node52407 : node52404;
																assign node52404 = (inp[0]) ? 4'b1000 : 4'b1010;
																assign node52407 = (inp[0]) ? 4'b1010 : 4'b1000;
														assign node52411 = (inp[3]) ? node52413 : 4'b1110;
															assign node52413 = (inp[0]) ? node52417 : node52414;
																assign node52414 = (inp[15]) ? 4'b1110 : 4'b1100;
																assign node52417 = (inp[15]) ? 4'b1100 : 4'b1110;
												assign node52420 = (inp[3]) ? node52438 : node52421;
													assign node52421 = (inp[15]) ? node52431 : node52422;
														assign node52422 = (inp[9]) ? node52426 : node52423;
															assign node52423 = (inp[0]) ? 4'b1100 : 4'b1110;
															assign node52426 = (inp[4]) ? node52428 : 4'b1010;
																assign node52428 = (inp[0]) ? 4'b1110 : 4'b1100;
														assign node52431 = (inp[0]) ? node52433 : 4'b1100;
															assign node52433 = (inp[9]) ? 4'b1100 : node52434;
																assign node52434 = (inp[4]) ? 4'b1010 : 4'b1110;
													assign node52438 = (inp[9]) ? node52442 : node52439;
														assign node52439 = (inp[4]) ? 4'b1010 : 4'b1110;
														assign node52442 = (inp[4]) ? node52446 : node52443;
															assign node52443 = (inp[0]) ? 4'b1000 : 4'b1010;
															assign node52446 = (inp[0]) ? node52448 : 4'b1110;
																assign node52448 = (inp[15]) ? 4'b1100 : 4'b1110;
											assign node52451 = (inp[3]) ? node52479 : node52452;
												assign node52452 = (inp[0]) ? node52466 : node52453;
													assign node52453 = (inp[15]) ? node52459 : node52454;
														assign node52454 = (inp[4]) ? node52456 : 4'b1010;
															assign node52456 = (inp[9]) ? 4'b1000 : 4'b1100;
														assign node52459 = (inp[4]) ? node52463 : node52460;
															assign node52460 = (inp[9]) ? 4'b1110 : 4'b1000;
															assign node52463 = (inp[9]) ? 4'b1010 : 4'b1110;
													assign node52466 = (inp[9]) ? node52474 : node52467;
														assign node52467 = (inp[4]) ? node52471 : node52468;
															assign node52468 = (inp[15]) ? 4'b1010 : 4'b1000;
															assign node52471 = (inp[2]) ? 4'b1110 : 4'b1100;
														assign node52474 = (inp[15]) ? 4'b1100 : node52475;
															assign node52475 = (inp[4]) ? 4'b1010 : 4'b1110;
												assign node52479 = (inp[4]) ? node52499 : node52480;
													assign node52480 = (inp[9]) ? node52494 : node52481;
														assign node52481 = (inp[2]) ? node52489 : node52482;
															assign node52482 = (inp[15]) ? node52486 : node52483;
																assign node52483 = (inp[0]) ? 4'b1010 : 4'b1000;
																assign node52486 = (inp[0]) ? 4'b1000 : 4'b1010;
															assign node52489 = (inp[0]) ? 4'b1010 : node52490;
																assign node52490 = (inp[15]) ? 4'b1010 : 4'b1000;
														assign node52494 = (inp[0]) ? 4'b1100 : node52495;
															assign node52495 = (inp[15]) ? 4'b1110 : 4'b1100;
													assign node52499 = (inp[9]) ? node52507 : node52500;
														assign node52500 = (inp[0]) ? node52504 : node52501;
															assign node52501 = (inp[15]) ? 4'b1110 : 4'b1100;
															assign node52504 = (inp[15]) ? 4'b1100 : 4'b1110;
														assign node52507 = (inp[2]) ? 4'b1010 : node52508;
															assign node52508 = (inp[0]) ? node52512 : node52509;
																assign node52509 = (inp[15]) ? 4'b1010 : 4'b1000;
																assign node52512 = (inp[15]) ? 4'b1000 : 4'b1010;
										assign node52516 = (inp[15]) ? node52558 : node52517;
											assign node52517 = (inp[0]) ? node52533 : node52518;
												assign node52518 = (inp[3]) ? node52526 : node52519;
													assign node52519 = (inp[9]) ? node52523 : node52520;
														assign node52520 = (inp[4]) ? 4'b1100 : 4'b1010;
														assign node52523 = (inp[4]) ? 4'b1000 : 4'b1100;
													assign node52526 = (inp[9]) ? node52530 : node52527;
														assign node52527 = (inp[4]) ? 4'b1100 : 4'b1000;
														assign node52530 = (inp[4]) ? 4'b1000 : 4'b1100;
												assign node52533 = (inp[12]) ? node52549 : node52534;
													assign node52534 = (inp[2]) ? node52542 : node52535;
														assign node52535 = (inp[9]) ? node52539 : node52536;
															assign node52536 = (inp[4]) ? 4'b1110 : 4'b1010;
															assign node52539 = (inp[4]) ? 4'b1010 : 4'b1110;
														assign node52542 = (inp[9]) ? node52546 : node52543;
															assign node52543 = (inp[3]) ? 4'b1010 : 4'b1000;
															assign node52546 = (inp[4]) ? 4'b1010 : 4'b1110;
													assign node52549 = (inp[9]) ? node52555 : node52550;
														assign node52550 = (inp[4]) ? 4'b1110 : node52551;
															assign node52551 = (inp[3]) ? 4'b1010 : 4'b1000;
														assign node52555 = (inp[4]) ? 4'b1010 : 4'b1110;
											assign node52558 = (inp[0]) ? node52572 : node52559;
												assign node52559 = (inp[3]) ? node52567 : node52560;
													assign node52560 = (inp[4]) ? node52564 : node52561;
														assign node52561 = (inp[9]) ? 4'b1110 : 4'b1000;
														assign node52564 = (inp[9]) ? 4'b1010 : 4'b1110;
													assign node52567 = (inp[4]) ? node52569 : 4'b1110;
														assign node52569 = (inp[9]) ? 4'b1010 : 4'b1110;
												assign node52572 = (inp[4]) ? node52578 : node52573;
													assign node52573 = (inp[9]) ? 4'b1100 : node52574;
														assign node52574 = (inp[3]) ? 4'b1000 : 4'b1010;
													assign node52578 = (inp[9]) ? 4'b1000 : 4'b1100;
								assign node52581 = (inp[14]) ? node52863 : node52582;
									assign node52582 = (inp[2]) ? node52702 : node52583;
										assign node52583 = (inp[9]) ? node52655 : node52584;
											assign node52584 = (inp[4]) ? node52626 : node52585;
												assign node52585 = (inp[10]) ? node52611 : node52586;
													assign node52586 = (inp[12]) ? node52600 : node52587;
														assign node52587 = (inp[0]) ? node52593 : node52588;
															assign node52588 = (inp[15]) ? 4'b1110 : node52589;
																assign node52589 = (inp[3]) ? 4'b1100 : 4'b1110;
															assign node52593 = (inp[3]) ? node52597 : node52594;
																assign node52594 = (inp[15]) ? 4'b1110 : 4'b1100;
																assign node52597 = (inp[15]) ? 4'b1100 : 4'b1110;
														assign node52600 = (inp[0]) ? node52606 : node52601;
															assign node52601 = (inp[3]) ? node52603 : 4'b1010;
																assign node52603 = (inp[15]) ? 4'b1010 : 4'b1000;
															assign node52606 = (inp[15]) ? node52608 : 4'b1000;
																assign node52608 = (inp[3]) ? 4'b1000 : 4'b1010;
													assign node52611 = (inp[0]) ? node52619 : node52612;
														assign node52612 = (inp[3]) ? node52616 : node52613;
															assign node52613 = (inp[15]) ? 4'b1000 : 4'b1010;
															assign node52616 = (inp[15]) ? 4'b1010 : 4'b1000;
														assign node52619 = (inp[3]) ? node52623 : node52620;
															assign node52620 = (inp[15]) ? 4'b1010 : 4'b1000;
															assign node52623 = (inp[15]) ? 4'b1000 : 4'b1010;
												assign node52626 = (inp[12]) ? node52648 : node52627;
													assign node52627 = (inp[10]) ? node52641 : node52628;
														assign node52628 = (inp[3]) ? node52634 : node52629;
															assign node52629 = (inp[15]) ? node52631 : 4'b1000;
																assign node52631 = (inp[0]) ? 4'b1010 : 4'b1000;
															assign node52634 = (inp[15]) ? node52638 : node52635;
																assign node52635 = (inp[0]) ? 4'b1010 : 4'b1000;
																assign node52638 = (inp[0]) ? 4'b1000 : 4'b1010;
														assign node52641 = (inp[0]) ? node52645 : node52642;
															assign node52642 = (inp[15]) ? 4'b1110 : 4'b1100;
															assign node52645 = (inp[15]) ? 4'b1100 : 4'b1110;
													assign node52648 = (inp[15]) ? node52652 : node52649;
														assign node52649 = (inp[0]) ? 4'b1110 : 4'b1100;
														assign node52652 = (inp[0]) ? 4'b1100 : 4'b1110;
											assign node52655 = (inp[4]) ? node52679 : node52656;
												assign node52656 = (inp[12]) ? node52672 : node52657;
													assign node52657 = (inp[10]) ? node52665 : node52658;
														assign node52658 = (inp[3]) ? 4'b1000 : node52659;
															assign node52659 = (inp[15]) ? node52661 : 4'b1000;
																assign node52661 = (inp[0]) ? 4'b1010 : 4'b1000;
														assign node52665 = (inp[15]) ? node52669 : node52666;
															assign node52666 = (inp[0]) ? 4'b1110 : 4'b1100;
															assign node52669 = (inp[0]) ? 4'b1100 : 4'b1110;
													assign node52672 = (inp[0]) ? node52676 : node52673;
														assign node52673 = (inp[15]) ? 4'b1110 : 4'b1100;
														assign node52676 = (inp[15]) ? 4'b1100 : 4'b1110;
												assign node52679 = (inp[10]) ? node52695 : node52680;
													assign node52680 = (inp[12]) ? node52688 : node52681;
														assign node52681 = (inp[15]) ? node52685 : node52682;
															assign node52682 = (inp[0]) ? 4'b1110 : 4'b1100;
															assign node52685 = (inp[0]) ? 4'b1100 : 4'b1110;
														assign node52688 = (inp[15]) ? node52692 : node52689;
															assign node52689 = (inp[0]) ? 4'b1010 : 4'b1000;
															assign node52692 = (inp[0]) ? 4'b1000 : 4'b1010;
													assign node52695 = (inp[15]) ? node52699 : node52696;
														assign node52696 = (inp[0]) ? 4'b1010 : 4'b1000;
														assign node52699 = (inp[0]) ? 4'b1000 : 4'b1010;
										assign node52702 = (inp[4]) ? node52786 : node52703;
											assign node52703 = (inp[9]) ? node52761 : node52704;
												assign node52704 = (inp[12]) ? node52734 : node52705;
													assign node52705 = (inp[10]) ? node52721 : node52706;
														assign node52706 = (inp[3]) ? node52714 : node52707;
															assign node52707 = (inp[0]) ? node52711 : node52708;
																assign node52708 = (inp[15]) ? 4'b1101 : 4'b1111;
																assign node52711 = (inp[15]) ? 4'b1111 : 4'b1101;
															assign node52714 = (inp[0]) ? node52718 : node52715;
																assign node52715 = (inp[15]) ? 4'b1111 : 4'b1101;
																assign node52718 = (inp[15]) ? 4'b1101 : 4'b1111;
														assign node52721 = (inp[3]) ? node52729 : node52722;
															assign node52722 = (inp[0]) ? node52726 : node52723;
																assign node52723 = (inp[15]) ? 4'b1001 : 4'b1011;
																assign node52726 = (inp[15]) ? 4'b1011 : 4'b1001;
															assign node52729 = (inp[15]) ? 4'b1011 : node52730;
																assign node52730 = (inp[0]) ? 4'b1011 : 4'b1001;
													assign node52734 = (inp[10]) ? node52748 : node52735;
														assign node52735 = (inp[3]) ? node52741 : node52736;
															assign node52736 = (inp[15]) ? node52738 : 4'b1011;
																assign node52738 = (inp[0]) ? 4'b1011 : 4'b1001;
															assign node52741 = (inp[15]) ? node52745 : node52742;
																assign node52742 = (inp[0]) ? 4'b1011 : 4'b1001;
																assign node52745 = (inp[0]) ? 4'b1001 : 4'b1011;
														assign node52748 = (inp[0]) ? node52756 : node52749;
															assign node52749 = (inp[3]) ? node52753 : node52750;
																assign node52750 = (inp[15]) ? 4'b1001 : 4'b1011;
																assign node52753 = (inp[15]) ? 4'b1011 : 4'b1001;
															assign node52756 = (inp[15]) ? 4'b1001 : node52757;
																assign node52757 = (inp[3]) ? 4'b1011 : 4'b1001;
												assign node52761 = (inp[10]) ? node52779 : node52762;
													assign node52762 = (inp[12]) ? node52772 : node52763;
														assign node52763 = (inp[3]) ? 4'b1011 : node52764;
															assign node52764 = (inp[0]) ? node52768 : node52765;
																assign node52765 = (inp[15]) ? 4'b1001 : 4'b1011;
																assign node52768 = (inp[15]) ? 4'b1011 : 4'b1001;
														assign node52772 = (inp[3]) ? node52774 : 4'b1101;
															assign node52774 = (inp[15]) ? node52776 : 4'b1111;
																assign node52776 = (inp[0]) ? 4'b1101 : 4'b1111;
													assign node52779 = (inp[15]) ? node52783 : node52780;
														assign node52780 = (inp[0]) ? 4'b1111 : 4'b1101;
														assign node52783 = (inp[0]) ? 4'b1101 : 4'b1111;
											assign node52786 = (inp[9]) ? node52836 : node52787;
												assign node52787 = (inp[12]) ? node52809 : node52788;
													assign node52788 = (inp[10]) ? node52798 : node52789;
														assign node52789 = (inp[3]) ? 4'b1011 : node52790;
															assign node52790 = (inp[0]) ? node52794 : node52791;
																assign node52791 = (inp[15]) ? 4'b1001 : 4'b1011;
																assign node52794 = (inp[15]) ? 4'b1011 : 4'b1001;
														assign node52798 = (inp[3]) ? node52804 : node52799;
															assign node52799 = (inp[0]) ? 4'b1111 : node52800;
																assign node52800 = (inp[15]) ? 4'b1111 : 4'b1101;
															assign node52804 = (inp[0]) ? node52806 : 4'b1101;
																assign node52806 = (inp[15]) ? 4'b1101 : 4'b1111;
													assign node52809 = (inp[3]) ? node52825 : node52810;
														assign node52810 = (inp[10]) ? node52818 : node52811;
															assign node52811 = (inp[0]) ? node52815 : node52812;
																assign node52812 = (inp[15]) ? 4'b1111 : 4'b1101;
																assign node52815 = (inp[15]) ? 4'b1101 : 4'b1111;
															assign node52818 = (inp[15]) ? node52822 : node52819;
																assign node52819 = (inp[0]) ? 4'b1111 : 4'b1101;
																assign node52822 = (inp[0]) ? 4'b1101 : 4'b1111;
														assign node52825 = (inp[10]) ? node52831 : node52826;
															assign node52826 = (inp[15]) ? node52828 : 4'b1111;
																assign node52828 = (inp[0]) ? 4'b1101 : 4'b1111;
															assign node52831 = (inp[15]) ? 4'b1111 : node52832;
																assign node52832 = (inp[0]) ? 4'b1111 : 4'b1101;
												assign node52836 = (inp[10]) ? node52856 : node52837;
													assign node52837 = (inp[12]) ? node52851 : node52838;
														assign node52838 = (inp[3]) ? node52846 : node52839;
															assign node52839 = (inp[15]) ? node52843 : node52840;
																assign node52840 = (inp[0]) ? 4'b1111 : 4'b1101;
																assign node52843 = (inp[0]) ? 4'b1101 : 4'b1111;
															assign node52846 = (inp[0]) ? 4'b1111 : node52847;
																assign node52847 = (inp[15]) ? 4'b1111 : 4'b1101;
														assign node52851 = (inp[0]) ? 4'b1011 : node52852;
															assign node52852 = (inp[15]) ? 4'b1011 : 4'b1001;
													assign node52856 = (inp[0]) ? node52860 : node52857;
														assign node52857 = (inp[15]) ? 4'b1011 : 4'b1001;
														assign node52860 = (inp[15]) ? 4'b1001 : 4'b1011;
									assign node52863 = (inp[15]) ? node52967 : node52864;
										assign node52864 = (inp[0]) ? node52910 : node52865;
											assign node52865 = (inp[3]) ? node52889 : node52866;
												assign node52866 = (inp[4]) ? node52878 : node52867;
													assign node52867 = (inp[9]) ? node52873 : node52868;
														assign node52868 = (inp[10]) ? 4'b1011 : node52869;
															assign node52869 = (inp[12]) ? 4'b1011 : 4'b1111;
														assign node52873 = (inp[10]) ? 4'b1101 : node52874;
															assign node52874 = (inp[12]) ? 4'b1101 : 4'b1011;
													assign node52878 = (inp[9]) ? node52884 : node52879;
														assign node52879 = (inp[12]) ? 4'b1101 : node52880;
															assign node52880 = (inp[10]) ? 4'b1101 : 4'b1011;
														assign node52884 = (inp[12]) ? 4'b1001 : node52885;
															assign node52885 = (inp[10]) ? 4'b1001 : 4'b1101;
												assign node52889 = (inp[12]) ? node52903 : node52890;
													assign node52890 = (inp[9]) ? node52898 : node52891;
														assign node52891 = (inp[2]) ? node52893 : 4'b1101;
															assign node52893 = (inp[4]) ? node52895 : 4'b1001;
																assign node52895 = (inp[10]) ? 4'b1101 : 4'b1001;
														assign node52898 = (inp[4]) ? node52900 : 4'b1101;
															assign node52900 = (inp[10]) ? 4'b1001 : 4'b1101;
													assign node52903 = (inp[4]) ? node52907 : node52904;
														assign node52904 = (inp[9]) ? 4'b1101 : 4'b1001;
														assign node52907 = (inp[9]) ? 4'b1001 : 4'b1101;
											assign node52910 = (inp[3]) ? node52936 : node52911;
												assign node52911 = (inp[4]) ? node52923 : node52912;
													assign node52912 = (inp[9]) ? node52918 : node52913;
														assign node52913 = (inp[12]) ? 4'b1001 : node52914;
															assign node52914 = (inp[10]) ? 4'b1001 : 4'b1101;
														assign node52918 = (inp[12]) ? 4'b1111 : node52919;
															assign node52919 = (inp[10]) ? 4'b1111 : 4'b1001;
													assign node52923 = (inp[9]) ? node52931 : node52924;
														assign node52924 = (inp[2]) ? 4'b1111 : node52925;
															assign node52925 = (inp[12]) ? 4'b1111 : node52926;
																assign node52926 = (inp[10]) ? 4'b1111 : 4'b1001;
														assign node52931 = (inp[12]) ? 4'b1011 : node52932;
															assign node52932 = (inp[10]) ? 4'b1011 : 4'b1111;
												assign node52936 = (inp[2]) ? node52960 : node52937;
													assign node52937 = (inp[12]) ? node52953 : node52938;
														assign node52938 = (inp[4]) ? node52946 : node52939;
															assign node52939 = (inp[10]) ? node52943 : node52940;
																assign node52940 = (inp[9]) ? 4'b1011 : 4'b1111;
																assign node52943 = (inp[9]) ? 4'b1111 : 4'b1011;
															assign node52946 = (inp[10]) ? node52950 : node52947;
																assign node52947 = (inp[9]) ? 4'b1111 : 4'b1011;
																assign node52950 = (inp[9]) ? 4'b1011 : 4'b1111;
														assign node52953 = (inp[4]) ? node52957 : node52954;
															assign node52954 = (inp[9]) ? 4'b1111 : 4'b1011;
															assign node52957 = (inp[9]) ? 4'b1011 : 4'b1111;
													assign node52960 = (inp[9]) ? node52964 : node52961;
														assign node52961 = (inp[4]) ? 4'b1111 : 4'b1011;
														assign node52964 = (inp[4]) ? 4'b1011 : 4'b1111;
										assign node52967 = (inp[0]) ? node53021 : node52968;
											assign node52968 = (inp[3]) ? node52992 : node52969;
												assign node52969 = (inp[4]) ? node52981 : node52970;
													assign node52970 = (inp[9]) ? node52976 : node52971;
														assign node52971 = (inp[10]) ? 4'b1001 : node52972;
															assign node52972 = (inp[12]) ? 4'b1001 : 4'b1101;
														assign node52976 = (inp[12]) ? 4'b1111 : node52977;
															assign node52977 = (inp[10]) ? 4'b1111 : 4'b1001;
													assign node52981 = (inp[9]) ? node52987 : node52982;
														assign node52982 = (inp[10]) ? 4'b1111 : node52983;
															assign node52983 = (inp[12]) ? 4'b1111 : 4'b1001;
														assign node52987 = (inp[10]) ? 4'b1011 : node52988;
															assign node52988 = (inp[12]) ? 4'b1011 : 4'b1111;
												assign node52992 = (inp[2]) ? node53006 : node52993;
													assign node52993 = (inp[4]) ? node52999 : node52994;
														assign node52994 = (inp[9]) ? node52996 : 4'b1011;
															assign node52996 = (inp[10]) ? 4'b1111 : 4'b1011;
														assign node52999 = (inp[9]) ? node53001 : 4'b1111;
															assign node53001 = (inp[10]) ? 4'b1011 : node53002;
																assign node53002 = (inp[12]) ? 4'b1011 : 4'b1111;
													assign node53006 = (inp[12]) ? node53014 : node53007;
														assign node53007 = (inp[10]) ? node53009 : 4'b1011;
															assign node53009 = (inp[4]) ? node53011 : 4'b1011;
																assign node53011 = (inp[9]) ? 4'b1011 : 4'b1111;
														assign node53014 = (inp[4]) ? node53018 : node53015;
															assign node53015 = (inp[9]) ? 4'b1111 : 4'b1011;
															assign node53018 = (inp[9]) ? 4'b1011 : 4'b1111;
											assign node53021 = (inp[3]) ? node53045 : node53022;
												assign node53022 = (inp[9]) ? node53034 : node53023;
													assign node53023 = (inp[4]) ? node53029 : node53024;
														assign node53024 = (inp[10]) ? 4'b1011 : node53025;
															assign node53025 = (inp[12]) ? 4'b1011 : 4'b1111;
														assign node53029 = (inp[12]) ? 4'b1101 : node53030;
															assign node53030 = (inp[10]) ? 4'b1101 : 4'b1011;
													assign node53034 = (inp[4]) ? node53040 : node53035;
														assign node53035 = (inp[10]) ? 4'b1101 : node53036;
															assign node53036 = (inp[2]) ? 4'b1011 : 4'b1101;
														assign node53040 = (inp[10]) ? 4'b1001 : node53041;
															assign node53041 = (inp[12]) ? 4'b1001 : 4'b1101;
												assign node53045 = (inp[9]) ? node53057 : node53046;
													assign node53046 = (inp[4]) ? node53052 : node53047;
														assign node53047 = (inp[12]) ? 4'b1001 : node53048;
															assign node53048 = (inp[10]) ? 4'b1001 : 4'b1101;
														assign node53052 = (inp[10]) ? 4'b1101 : node53053;
															assign node53053 = (inp[12]) ? 4'b1101 : 4'b1001;
													assign node53057 = (inp[4]) ? node53063 : node53058;
														assign node53058 = (inp[10]) ? 4'b1101 : node53059;
															assign node53059 = (inp[12]) ? 4'b1101 : 4'b1001;
														assign node53063 = (inp[10]) ? 4'b1001 : node53064;
															assign node53064 = (inp[12]) ? 4'b1001 : 4'b1101;
							assign node53068 = (inp[8]) ? node53504 : node53069;
								assign node53069 = (inp[14]) ? node53317 : node53070;
									assign node53070 = (inp[2]) ? node53218 : node53071;
										assign node53071 = (inp[3]) ? node53151 : node53072;
											assign node53072 = (inp[10]) ? node53120 : node53073;
												assign node53073 = (inp[4]) ? node53099 : node53074;
													assign node53074 = (inp[0]) ? node53088 : node53075;
														assign node53075 = (inp[15]) ? node53083 : node53076;
															assign node53076 = (inp[12]) ? node53080 : node53077;
																assign node53077 = (inp[9]) ? 4'b1010 : 4'b1110;
																assign node53080 = (inp[9]) ? 4'b1100 : 4'b1010;
															assign node53083 = (inp[9]) ? node53085 : 4'b1000;
																assign node53085 = (inp[12]) ? 4'b1110 : 4'b1000;
														assign node53088 = (inp[15]) ? node53094 : node53089;
															assign node53089 = (inp[12]) ? 4'b1000 : node53090;
																assign node53090 = (inp[9]) ? 4'b1000 : 4'b1100;
															assign node53094 = (inp[9]) ? node53096 : 4'b1010;
																assign node53096 = (inp[12]) ? 4'b1100 : 4'b1010;
													assign node53099 = (inp[9]) ? node53109 : node53100;
														assign node53100 = (inp[12]) ? node53102 : 4'b1000;
															assign node53102 = (inp[15]) ? node53106 : node53103;
																assign node53103 = (inp[0]) ? 4'b1110 : 4'b1100;
																assign node53106 = (inp[0]) ? 4'b1100 : 4'b1110;
														assign node53109 = (inp[12]) ? node53115 : node53110;
															assign node53110 = (inp[15]) ? 4'b1110 : node53111;
																assign node53111 = (inp[0]) ? 4'b1110 : 4'b1100;
															assign node53115 = (inp[15]) ? 4'b1000 : node53116;
																assign node53116 = (inp[0]) ? 4'b1010 : 4'b1000;
												assign node53120 = (inp[4]) ? node53136 : node53121;
													assign node53121 = (inp[9]) ? node53123 : 4'b1000;
														assign node53123 = (inp[12]) ? node53131 : node53124;
															assign node53124 = (inp[0]) ? node53128 : node53125;
																assign node53125 = (inp[15]) ? 4'b1110 : 4'b1100;
																assign node53128 = (inp[15]) ? 4'b1100 : 4'b1110;
															assign node53131 = (inp[0]) ? node53133 : 4'b1100;
																assign node53133 = (inp[15]) ? 4'b1100 : 4'b1110;
													assign node53136 = (inp[9]) ? node53146 : node53137;
														assign node53137 = (inp[12]) ? 4'b1110 : node53138;
															assign node53138 = (inp[0]) ? node53142 : node53139;
																assign node53139 = (inp[15]) ? 4'b1110 : 4'b1100;
																assign node53142 = (inp[15]) ? 4'b1100 : 4'b1110;
														assign node53146 = (inp[0]) ? 4'b1000 : node53147;
															assign node53147 = (inp[15]) ? 4'b1010 : 4'b1000;
											assign node53151 = (inp[10]) ? node53185 : node53152;
												assign node53152 = (inp[15]) ? node53164 : node53153;
													assign node53153 = (inp[0]) ? node53159 : node53154;
														assign node53154 = (inp[4]) ? node53156 : 4'b1000;
															assign node53156 = (inp[9]) ? 4'b1000 : 4'b1100;
														assign node53159 = (inp[12]) ? 4'b1010 : node53160;
															assign node53160 = (inp[9]) ? 4'b1110 : 4'b1010;
													assign node53164 = (inp[0]) ? node53170 : node53165;
														assign node53165 = (inp[12]) ? node53167 : 4'b1110;
															assign node53167 = (inp[4]) ? 4'b1010 : 4'b1110;
														assign node53170 = (inp[4]) ? node53178 : node53171;
															assign node53171 = (inp[12]) ? node53175 : node53172;
																assign node53172 = (inp[9]) ? 4'b1000 : 4'b1100;
																assign node53175 = (inp[9]) ? 4'b1100 : 4'b1000;
															assign node53178 = (inp[9]) ? node53182 : node53179;
																assign node53179 = (inp[12]) ? 4'b1100 : 4'b1000;
																assign node53182 = (inp[12]) ? 4'b1000 : 4'b1100;
												assign node53185 = (inp[4]) ? node53201 : node53186;
													assign node53186 = (inp[9]) ? node53194 : node53187;
														assign node53187 = (inp[15]) ? node53191 : node53188;
															assign node53188 = (inp[0]) ? 4'b1010 : 4'b1000;
															assign node53191 = (inp[0]) ? 4'b1000 : 4'b1010;
														assign node53194 = (inp[12]) ? node53196 : 4'b1110;
															assign node53196 = (inp[0]) ? node53198 : 4'b1110;
																assign node53198 = (inp[15]) ? 4'b1100 : 4'b1110;
													assign node53201 = (inp[9]) ? node53207 : node53202;
														assign node53202 = (inp[15]) ? 4'b1110 : node53203;
															assign node53203 = (inp[0]) ? 4'b1110 : 4'b1100;
														assign node53207 = (inp[12]) ? node53213 : node53208;
															assign node53208 = (inp[0]) ? node53210 : 4'b1000;
																assign node53210 = (inp[15]) ? 4'b1000 : 4'b1010;
															assign node53213 = (inp[15]) ? node53215 : 4'b1000;
																assign node53215 = (inp[0]) ? 4'b1000 : 4'b1010;
										assign node53218 = (inp[9]) ? node53266 : node53219;
											assign node53219 = (inp[4]) ? node53249 : node53220;
												assign node53220 = (inp[12]) ? node53240 : node53221;
													assign node53221 = (inp[10]) ? node53235 : node53222;
														assign node53222 = (inp[15]) ? node53228 : node53223;
															assign node53223 = (inp[0]) ? 4'b1111 : node53224;
																assign node53224 = (inp[3]) ? 4'b1101 : 4'b1111;
															assign node53228 = (inp[0]) ? node53232 : node53229;
																assign node53229 = (inp[3]) ? 4'b1111 : 4'b1101;
																assign node53232 = (inp[3]) ? 4'b1101 : 4'b1111;
														assign node53235 = (inp[15]) ? 4'b1011 : node53236;
															assign node53236 = (inp[0]) ? 4'b1001 : 4'b1011;
													assign node53240 = (inp[0]) ? 4'b1001 : node53241;
														assign node53241 = (inp[3]) ? node53245 : node53242;
															assign node53242 = (inp[15]) ? 4'b1001 : 4'b1011;
															assign node53245 = (inp[15]) ? 4'b1011 : 4'b1001;
												assign node53249 = (inp[12]) ? node53259 : node53250;
													assign node53250 = (inp[10]) ? 4'b1111 : node53251;
														assign node53251 = (inp[0]) ? 4'b1001 : node53252;
															assign node53252 = (inp[15]) ? node53254 : 4'b1001;
																assign node53254 = (inp[3]) ? 4'b1011 : 4'b1001;
													assign node53259 = (inp[15]) ? node53263 : node53260;
														assign node53260 = (inp[0]) ? 4'b1111 : 4'b1101;
														assign node53263 = (inp[0]) ? 4'b1101 : 4'b1111;
											assign node53266 = (inp[4]) ? node53292 : node53267;
												assign node53267 = (inp[12]) ? node53275 : node53268;
													assign node53268 = (inp[10]) ? node53270 : 4'b1001;
														assign node53270 = (inp[15]) ? node53272 : 4'b1101;
															assign node53272 = (inp[0]) ? 4'b1101 : 4'b1111;
													assign node53275 = (inp[10]) ? node53283 : node53276;
														assign node53276 = (inp[0]) ? node53280 : node53277;
															assign node53277 = (inp[15]) ? 4'b1111 : 4'b1101;
															assign node53280 = (inp[15]) ? 4'b1101 : 4'b1111;
														assign node53283 = (inp[3]) ? node53285 : 4'b1101;
															assign node53285 = (inp[0]) ? node53289 : node53286;
																assign node53286 = (inp[15]) ? 4'b1111 : 4'b1101;
																assign node53289 = (inp[15]) ? 4'b1101 : 4'b1111;
												assign node53292 = (inp[10]) ? node53306 : node53293;
													assign node53293 = (inp[12]) ? node53301 : node53294;
														assign node53294 = (inp[0]) ? node53298 : node53295;
															assign node53295 = (inp[15]) ? 4'b1111 : 4'b1101;
															assign node53298 = (inp[15]) ? 4'b1101 : 4'b1111;
														assign node53301 = (inp[15]) ? 4'b1011 : node53302;
															assign node53302 = (inp[0]) ? 4'b1011 : 4'b1001;
													assign node53306 = (inp[12]) ? node53312 : node53307;
														assign node53307 = (inp[0]) ? node53309 : 4'b1001;
															assign node53309 = (inp[15]) ? 4'b1001 : 4'b1011;
														assign node53312 = (inp[0]) ? 4'b1001 : node53313;
															assign node53313 = (inp[15]) ? 4'b1011 : 4'b1001;
									assign node53317 = (inp[0]) ? node53397 : node53318;
										assign node53318 = (inp[15]) ? node53350 : node53319;
											assign node53319 = (inp[9]) ? node53339 : node53320;
												assign node53320 = (inp[4]) ? node53332 : node53321;
													assign node53321 = (inp[3]) ? node53327 : node53322;
														assign node53322 = (inp[12]) ? 4'b1011 : node53323;
															assign node53323 = (inp[10]) ? 4'b1011 : 4'b1111;
														assign node53327 = (inp[10]) ? 4'b1001 : node53328;
															assign node53328 = (inp[12]) ? 4'b1001 : 4'b1101;
													assign node53332 = (inp[10]) ? 4'b1101 : node53333;
														assign node53333 = (inp[12]) ? 4'b1101 : node53334;
															assign node53334 = (inp[3]) ? 4'b1001 : 4'b1011;
												assign node53339 = (inp[4]) ? node53345 : node53340;
													assign node53340 = (inp[10]) ? 4'b1101 : node53341;
														assign node53341 = (inp[12]) ? 4'b1101 : 4'b1001;
													assign node53345 = (inp[10]) ? 4'b1001 : node53346;
														assign node53346 = (inp[12]) ? 4'b1001 : 4'b1101;
											assign node53350 = (inp[3]) ? node53370 : node53351;
												assign node53351 = (inp[9]) ? node53359 : node53352;
													assign node53352 = (inp[4]) ? node53354 : 4'b1001;
														assign node53354 = (inp[12]) ? 4'b1111 : node53355;
															assign node53355 = (inp[10]) ? 4'b1111 : 4'b1001;
													assign node53359 = (inp[4]) ? node53365 : node53360;
														assign node53360 = (inp[10]) ? 4'b1111 : node53361;
															assign node53361 = (inp[12]) ? 4'b1111 : 4'b1001;
														assign node53365 = (inp[10]) ? 4'b1011 : node53366;
															assign node53366 = (inp[12]) ? 4'b1011 : 4'b1111;
												assign node53370 = (inp[2]) ? node53384 : node53371;
													assign node53371 = (inp[9]) ? node53377 : node53372;
														assign node53372 = (inp[4]) ? node53374 : 4'b1011;
															assign node53374 = (inp[12]) ? 4'b1111 : 4'b1011;
														assign node53377 = (inp[4]) ? node53381 : node53378;
															assign node53378 = (inp[12]) ? 4'b1111 : 4'b1011;
															assign node53381 = (inp[12]) ? 4'b1011 : 4'b1111;
													assign node53384 = (inp[4]) ? node53386 : 4'b1111;
														assign node53386 = (inp[9]) ? node53392 : node53387;
															assign node53387 = (inp[10]) ? 4'b1111 : node53388;
																assign node53388 = (inp[12]) ? 4'b1111 : 4'b1011;
															assign node53392 = (inp[10]) ? 4'b1011 : node53393;
																assign node53393 = (inp[12]) ? 4'b1011 : 4'b1111;
										assign node53397 = (inp[15]) ? node53455 : node53398;
											assign node53398 = (inp[3]) ? node53420 : node53399;
												assign node53399 = (inp[4]) ? node53409 : node53400;
													assign node53400 = (inp[9]) ? node53406 : node53401;
														assign node53401 = (inp[12]) ? 4'b1001 : node53402;
															assign node53402 = (inp[10]) ? 4'b1001 : 4'b1101;
														assign node53406 = (inp[10]) ? 4'b1111 : 4'b1001;
													assign node53409 = (inp[9]) ? node53415 : node53410;
														assign node53410 = (inp[10]) ? 4'b1111 : node53411;
															assign node53411 = (inp[12]) ? 4'b1111 : 4'b1001;
														assign node53415 = (inp[10]) ? 4'b1011 : node53416;
															assign node53416 = (inp[2]) ? 4'b1111 : 4'b1011;
												assign node53420 = (inp[2]) ? node53434 : node53421;
													assign node53421 = (inp[12]) ? node53429 : node53422;
														assign node53422 = (inp[9]) ? node53424 : 4'b1011;
															assign node53424 = (inp[10]) ? node53426 : 4'b1111;
																assign node53426 = (inp[4]) ? 4'b1011 : 4'b1111;
														assign node53429 = (inp[4]) ? node53431 : 4'b1111;
															assign node53431 = (inp[9]) ? 4'b1011 : 4'b1111;
													assign node53434 = (inp[10]) ? node53448 : node53435;
														assign node53435 = (inp[9]) ? node53441 : node53436;
															assign node53436 = (inp[4]) ? 4'b1111 : node53437;
																assign node53437 = (inp[12]) ? 4'b1011 : 4'b1111;
															assign node53441 = (inp[4]) ? node53445 : node53442;
																assign node53442 = (inp[12]) ? 4'b1111 : 4'b1011;
																assign node53445 = (inp[12]) ? 4'b1011 : 4'b1111;
														assign node53448 = (inp[4]) ? node53452 : node53449;
															assign node53449 = (inp[9]) ? 4'b1111 : 4'b1011;
															assign node53452 = (inp[9]) ? 4'b1011 : 4'b1111;
											assign node53455 = (inp[3]) ? node53481 : node53456;
												assign node53456 = (inp[4]) ? node53468 : node53457;
													assign node53457 = (inp[9]) ? node53463 : node53458;
														assign node53458 = (inp[10]) ? 4'b1011 : node53459;
															assign node53459 = (inp[12]) ? 4'b1011 : 4'b1111;
														assign node53463 = (inp[12]) ? 4'b1101 : node53464;
															assign node53464 = (inp[10]) ? 4'b1101 : 4'b1011;
													assign node53468 = (inp[9]) ? node53476 : node53469;
														assign node53469 = (inp[2]) ? 4'b1101 : node53470;
															assign node53470 = (inp[10]) ? 4'b1101 : node53471;
																assign node53471 = (inp[12]) ? 4'b1101 : 4'b1011;
														assign node53476 = (inp[12]) ? 4'b1001 : node53477;
															assign node53477 = (inp[10]) ? 4'b1001 : 4'b1101;
												assign node53481 = (inp[9]) ? node53493 : node53482;
													assign node53482 = (inp[4]) ? node53488 : node53483;
														assign node53483 = (inp[12]) ? 4'b1001 : node53484;
															assign node53484 = (inp[10]) ? 4'b1001 : 4'b1101;
														assign node53488 = (inp[10]) ? 4'b1101 : node53489;
															assign node53489 = (inp[12]) ? 4'b1101 : 4'b1001;
													assign node53493 = (inp[4]) ? node53499 : node53494;
														assign node53494 = (inp[12]) ? 4'b1101 : node53495;
															assign node53495 = (inp[10]) ? 4'b1101 : 4'b1001;
														assign node53499 = (inp[12]) ? 4'b1001 : node53500;
															assign node53500 = (inp[10]) ? 4'b1001 : 4'b1101;
								assign node53504 = (inp[2]) ? node53814 : node53505;
									assign node53505 = (inp[14]) ? node53681 : node53506;
										assign node53506 = (inp[12]) ? node53598 : node53507;
											assign node53507 = (inp[15]) ? node53555 : node53508;
												assign node53508 = (inp[0]) ? node53526 : node53509;
													assign node53509 = (inp[3]) ? node53521 : node53510;
														assign node53510 = (inp[4]) ? node53516 : node53511;
															assign node53511 = (inp[9]) ? 4'b1011 : node53512;
																assign node53512 = (inp[10]) ? 4'b1011 : 4'b1111;
															assign node53516 = (inp[10]) ? 4'b1101 : node53517;
																assign node53517 = (inp[9]) ? 4'b1101 : 4'b1011;
														assign node53521 = (inp[4]) ? node53523 : 4'b1001;
															assign node53523 = (inp[9]) ? 4'b1001 : 4'b1101;
													assign node53526 = (inp[3]) ? node53540 : node53527;
														assign node53527 = (inp[10]) ? node53533 : node53528;
															assign node53528 = (inp[9]) ? node53530 : 4'b1001;
																assign node53530 = (inp[4]) ? 4'b1111 : 4'b1001;
															assign node53533 = (inp[9]) ? node53537 : node53534;
																assign node53534 = (inp[4]) ? 4'b1111 : 4'b1001;
																assign node53537 = (inp[4]) ? 4'b1011 : 4'b1111;
														assign node53540 = (inp[9]) ? node53548 : node53541;
															assign node53541 = (inp[10]) ? node53545 : node53542;
																assign node53542 = (inp[4]) ? 4'b1011 : 4'b1111;
																assign node53545 = (inp[4]) ? 4'b1111 : 4'b1011;
															assign node53548 = (inp[10]) ? node53552 : node53549;
																assign node53549 = (inp[4]) ? 4'b1111 : 4'b1011;
																assign node53552 = (inp[4]) ? 4'b1011 : 4'b1111;
												assign node53555 = (inp[0]) ? node53573 : node53556;
													assign node53556 = (inp[3]) ? node53566 : node53557;
														assign node53557 = (inp[9]) ? node53563 : node53558;
															assign node53558 = (inp[4]) ? 4'b1001 : node53559;
																assign node53559 = (inp[10]) ? 4'b1001 : 4'b1101;
															assign node53563 = (inp[10]) ? 4'b1011 : 4'b1111;
														assign node53566 = (inp[10]) ? node53570 : node53567;
															assign node53567 = (inp[4]) ? 4'b1011 : 4'b1111;
															assign node53570 = (inp[4]) ? 4'b1111 : 4'b1011;
													assign node53573 = (inp[3]) ? node53589 : node53574;
														assign node53574 = (inp[10]) ? node53582 : node53575;
															assign node53575 = (inp[4]) ? node53579 : node53576;
																assign node53576 = (inp[9]) ? 4'b1011 : 4'b1111;
																assign node53579 = (inp[9]) ? 4'b1101 : 4'b1011;
															assign node53582 = (inp[9]) ? node53586 : node53583;
																assign node53583 = (inp[4]) ? 4'b1101 : 4'b1011;
																assign node53586 = (inp[4]) ? 4'b1001 : 4'b1101;
														assign node53589 = (inp[10]) ? 4'b1001 : node53590;
															assign node53590 = (inp[9]) ? node53594 : node53591;
																assign node53591 = (inp[4]) ? 4'b1001 : 4'b1101;
																assign node53594 = (inp[4]) ? 4'b1101 : 4'b1001;
											assign node53598 = (inp[10]) ? node53648 : node53599;
												assign node53599 = (inp[3]) ? node53625 : node53600;
													assign node53600 = (inp[15]) ? node53614 : node53601;
														assign node53601 = (inp[0]) ? node53609 : node53602;
															assign node53602 = (inp[9]) ? node53606 : node53603;
																assign node53603 = (inp[4]) ? 4'b1101 : 4'b1011;
																assign node53606 = (inp[4]) ? 4'b1001 : 4'b1101;
															assign node53609 = (inp[4]) ? node53611 : 4'b1001;
																assign node53611 = (inp[9]) ? 4'b1011 : 4'b1111;
														assign node53614 = (inp[0]) ? node53620 : node53615;
															assign node53615 = (inp[9]) ? node53617 : 4'b1001;
																assign node53617 = (inp[4]) ? 4'b1011 : 4'b1111;
															assign node53620 = (inp[4]) ? 4'b1101 : node53621;
																assign node53621 = (inp[9]) ? 4'b1101 : 4'b1011;
													assign node53625 = (inp[0]) ? node53639 : node53626;
														assign node53626 = (inp[15]) ? node53634 : node53627;
															assign node53627 = (inp[9]) ? node53631 : node53628;
																assign node53628 = (inp[4]) ? 4'b1101 : 4'b1001;
																assign node53631 = (inp[4]) ? 4'b1001 : 4'b1101;
															assign node53634 = (inp[9]) ? node53636 : 4'b1011;
																assign node53636 = (inp[4]) ? 4'b1011 : 4'b1111;
														assign node53639 = (inp[15]) ? node53641 : 4'b1011;
															assign node53641 = (inp[4]) ? node53645 : node53642;
																assign node53642 = (inp[9]) ? 4'b1101 : 4'b1001;
																assign node53645 = (inp[9]) ? 4'b1001 : 4'b1101;
												assign node53648 = (inp[0]) ? node53664 : node53649;
													assign node53649 = (inp[15]) ? node53657 : node53650;
														assign node53650 = (inp[9]) ? node53654 : node53651;
															assign node53651 = (inp[4]) ? 4'b1101 : 4'b1001;
															assign node53654 = (inp[4]) ? 4'b1001 : 4'b1101;
														assign node53657 = (inp[3]) ? 4'b1111 : node53658;
															assign node53658 = (inp[9]) ? node53660 : 4'b1001;
																assign node53660 = (inp[4]) ? 4'b1011 : 4'b1111;
													assign node53664 = (inp[15]) ? node53674 : node53665;
														assign node53665 = (inp[4]) ? node53671 : node53666;
															assign node53666 = (inp[9]) ? 4'b1111 : node53667;
																assign node53667 = (inp[3]) ? 4'b1011 : 4'b1001;
															assign node53671 = (inp[9]) ? 4'b1011 : 4'b1111;
														assign node53674 = (inp[4]) ? node53678 : node53675;
															assign node53675 = (inp[9]) ? 4'b1101 : 4'b1011;
															assign node53678 = (inp[9]) ? 4'b1001 : 4'b1101;
										assign node53681 = (inp[15]) ? node53749 : node53682;
											assign node53682 = (inp[0]) ? node53716 : node53683;
												assign node53683 = (inp[3]) ? node53703 : node53684;
													assign node53684 = (inp[9]) ? node53692 : node53685;
														assign node53685 = (inp[4]) ? node53689 : node53686;
															assign node53686 = (inp[10]) ? 4'b1010 : 4'b1110;
															assign node53689 = (inp[10]) ? 4'b1100 : 4'b1010;
														assign node53692 = (inp[4]) ? node53698 : node53693;
															assign node53693 = (inp[10]) ? 4'b1100 : node53694;
																assign node53694 = (inp[12]) ? 4'b1100 : 4'b1010;
															assign node53698 = (inp[10]) ? 4'b1000 : node53699;
																assign node53699 = (inp[12]) ? 4'b1000 : 4'b1100;
													assign node53703 = (inp[12]) ? node53709 : node53704;
														assign node53704 = (inp[4]) ? node53706 : 4'b1000;
															assign node53706 = (inp[10]) ? 4'b1100 : 4'b1000;
														assign node53709 = (inp[4]) ? node53713 : node53710;
															assign node53710 = (inp[9]) ? 4'b1100 : 4'b1000;
															assign node53713 = (inp[9]) ? 4'b1000 : 4'b1100;
												assign node53716 = (inp[3]) ? node53730 : node53717;
													assign node53717 = (inp[9]) ? node53725 : node53718;
														assign node53718 = (inp[12]) ? 4'b1110 : node53719;
															assign node53719 = (inp[4]) ? 4'b1000 : node53720;
																assign node53720 = (inp[10]) ? 4'b1000 : 4'b1100;
														assign node53725 = (inp[4]) ? node53727 : 4'b1110;
															assign node53727 = (inp[10]) ? 4'b1010 : 4'b1110;
													assign node53730 = (inp[10]) ? node53744 : node53731;
														assign node53731 = (inp[9]) ? node53739 : node53732;
															assign node53732 = (inp[12]) ? node53736 : node53733;
																assign node53733 = (inp[4]) ? 4'b1010 : 4'b1110;
																assign node53736 = (inp[4]) ? 4'b1110 : 4'b1010;
															assign node53739 = (inp[4]) ? node53741 : 4'b1010;
																assign node53741 = (inp[12]) ? 4'b1010 : 4'b1110;
														assign node53744 = (inp[9]) ? 4'b1010 : node53745;
															assign node53745 = (inp[4]) ? 4'b1110 : 4'b1010;
											assign node53749 = (inp[0]) ? node53785 : node53750;
												assign node53750 = (inp[3]) ? node53770 : node53751;
													assign node53751 = (inp[4]) ? node53759 : node53752;
														assign node53752 = (inp[9]) ? node53754 : 4'b1000;
															assign node53754 = (inp[12]) ? 4'b1110 : node53755;
																assign node53755 = (inp[10]) ? 4'b1110 : 4'b1000;
														assign node53759 = (inp[9]) ? node53765 : node53760;
															assign node53760 = (inp[10]) ? 4'b1110 : node53761;
																assign node53761 = (inp[12]) ? 4'b1110 : 4'b1000;
															assign node53765 = (inp[10]) ? 4'b1010 : node53766;
																assign node53766 = (inp[12]) ? 4'b1010 : 4'b1110;
													assign node53770 = (inp[4]) ? node53776 : node53771;
														assign node53771 = (inp[9]) ? 4'b1110 : node53772;
															assign node53772 = (inp[12]) ? 4'b1010 : 4'b1110;
														assign node53776 = (inp[12]) ? node53782 : node53777;
															assign node53777 = (inp[10]) ? 4'b1110 : node53778;
																assign node53778 = (inp[9]) ? 4'b1110 : 4'b1010;
															assign node53782 = (inp[9]) ? 4'b1010 : 4'b1110;
												assign node53785 = (inp[3]) ? node53795 : node53786;
													assign node53786 = (inp[4]) ? 4'b1100 : node53787;
														assign node53787 = (inp[9]) ? node53789 : 4'b1010;
															assign node53789 = (inp[12]) ? 4'b1100 : node53790;
																assign node53790 = (inp[10]) ? 4'b1100 : 4'b1010;
													assign node53795 = (inp[4]) ? node53807 : node53796;
														assign node53796 = (inp[9]) ? node53802 : node53797;
															assign node53797 = (inp[10]) ? 4'b1000 : node53798;
																assign node53798 = (inp[12]) ? 4'b1000 : 4'b1100;
															assign node53802 = (inp[12]) ? 4'b1100 : node53803;
																assign node53803 = (inp[10]) ? 4'b1100 : 4'b1000;
														assign node53807 = (inp[9]) ? 4'b1000 : node53808;
															assign node53808 = (inp[10]) ? 4'b1100 : node53809;
																assign node53809 = (inp[12]) ? 4'b1100 : 4'b1000;
									assign node53814 = (inp[10]) ? node53974 : node53815;
										assign node53815 = (inp[14]) ? node53901 : node53816;
											assign node53816 = (inp[9]) ? node53862 : node53817;
												assign node53817 = (inp[4]) ? node53839 : node53818;
													assign node53818 = (inp[12]) ? node53834 : node53819;
														assign node53819 = (inp[0]) ? node53827 : node53820;
															assign node53820 = (inp[15]) ? node53824 : node53821;
																assign node53821 = (inp[3]) ? 4'b1100 : 4'b1110;
																assign node53824 = (inp[3]) ? 4'b1110 : 4'b1100;
															assign node53827 = (inp[3]) ? node53831 : node53828;
																assign node53828 = (inp[15]) ? 4'b1110 : 4'b1100;
																assign node53831 = (inp[15]) ? 4'b1100 : 4'b1110;
														assign node53834 = (inp[0]) ? 4'b1010 : node53835;
															assign node53835 = (inp[15]) ? 4'b1010 : 4'b1000;
													assign node53839 = (inp[12]) ? node53849 : node53840;
														assign node53840 = (inp[3]) ? 4'b1010 : node53841;
															assign node53841 = (inp[15]) ? node53845 : node53842;
																assign node53842 = (inp[0]) ? 4'b1000 : 4'b1010;
																assign node53845 = (inp[0]) ? 4'b1010 : 4'b1000;
														assign node53849 = (inp[3]) ? node53855 : node53850;
															assign node53850 = (inp[15]) ? 4'b1110 : node53851;
																assign node53851 = (inp[0]) ? 4'b1110 : 4'b1100;
															assign node53855 = (inp[0]) ? node53859 : node53856;
																assign node53856 = (inp[15]) ? 4'b1110 : 4'b1100;
																assign node53859 = (inp[15]) ? 4'b1100 : 4'b1110;
												assign node53862 = (inp[15]) ? node53880 : node53863;
													assign node53863 = (inp[0]) ? node53871 : node53864;
														assign node53864 = (inp[12]) ? node53868 : node53865;
															assign node53865 = (inp[3]) ? 4'b1100 : 4'b1010;
															assign node53868 = (inp[4]) ? 4'b1000 : 4'b1100;
														assign node53871 = (inp[12]) ? node53877 : node53872;
															assign node53872 = (inp[4]) ? 4'b1110 : node53873;
																assign node53873 = (inp[3]) ? 4'b1010 : 4'b1000;
															assign node53877 = (inp[4]) ? 4'b1010 : 4'b1110;
													assign node53880 = (inp[0]) ? node53888 : node53881;
														assign node53881 = (inp[4]) ? 4'b1110 : node53882;
															assign node53882 = (inp[3]) ? node53884 : 4'b1000;
																assign node53884 = (inp[12]) ? 4'b1110 : 4'b1010;
														assign node53888 = (inp[3]) ? node53894 : node53889;
															assign node53889 = (inp[12]) ? node53891 : 4'b1100;
																assign node53891 = (inp[4]) ? 4'b1000 : 4'b1100;
															assign node53894 = (inp[4]) ? node53898 : node53895;
																assign node53895 = (inp[12]) ? 4'b1100 : 4'b1000;
																assign node53898 = (inp[12]) ? 4'b1000 : 4'b1100;
											assign node53901 = (inp[9]) ? node53943 : node53902;
												assign node53902 = (inp[15]) ? node53920 : node53903;
													assign node53903 = (inp[0]) ? node53913 : node53904;
														assign node53904 = (inp[3]) ? 4'b1100 : node53905;
															assign node53905 = (inp[4]) ? node53909 : node53906;
																assign node53906 = (inp[12]) ? 4'b1010 : 4'b1110;
																assign node53909 = (inp[12]) ? 4'b1100 : 4'b1010;
														assign node53913 = (inp[3]) ? 4'b1010 : node53914;
															assign node53914 = (inp[4]) ? 4'b1110 : node53915;
																assign node53915 = (inp[12]) ? 4'b1000 : 4'b1100;
													assign node53920 = (inp[0]) ? node53928 : node53921;
														assign node53921 = (inp[3]) ? 4'b1010 : node53922;
															assign node53922 = (inp[12]) ? 4'b1000 : node53923;
																assign node53923 = (inp[4]) ? 4'b1000 : 4'b1100;
														assign node53928 = (inp[3]) ? node53936 : node53929;
															assign node53929 = (inp[4]) ? node53933 : node53930;
																assign node53930 = (inp[12]) ? 4'b1010 : 4'b1110;
																assign node53933 = (inp[12]) ? 4'b1100 : 4'b1010;
															assign node53936 = (inp[4]) ? node53940 : node53937;
																assign node53937 = (inp[12]) ? 4'b1000 : 4'b1100;
																assign node53940 = (inp[12]) ? 4'b1100 : 4'b1000;
												assign node53943 = (inp[4]) ? node53963 : node53944;
													assign node53944 = (inp[12]) ? node53952 : node53945;
														assign node53945 = (inp[0]) ? 4'b1010 : node53946;
															assign node53946 = (inp[15]) ? node53948 : 4'b1000;
																assign node53948 = (inp[3]) ? 4'b1010 : 4'b1000;
														assign node53952 = (inp[3]) ? node53958 : node53953;
															assign node53953 = (inp[0]) ? node53955 : 4'b1100;
																assign node53955 = (inp[15]) ? 4'b1100 : 4'b1110;
															assign node53958 = (inp[15]) ? node53960 : 4'b1110;
																assign node53960 = (inp[0]) ? 4'b1100 : 4'b1110;
													assign node53963 = (inp[12]) ? node53969 : node53964;
														assign node53964 = (inp[15]) ? node53966 : 4'b1100;
															assign node53966 = (inp[0]) ? 4'b1100 : 4'b1110;
														assign node53969 = (inp[15]) ? node53971 : 4'b1000;
															assign node53971 = (inp[0]) ? 4'b1000 : 4'b1010;
										assign node53974 = (inp[12]) ? node54044 : node53975;
											assign node53975 = (inp[14]) ? node54013 : node53976;
												assign node53976 = (inp[15]) ? node53996 : node53977;
													assign node53977 = (inp[0]) ? node53987 : node53978;
														assign node53978 = (inp[4]) ? node53984 : node53979;
															assign node53979 = (inp[3]) ? node53981 : 4'b1010;
																assign node53981 = (inp[9]) ? 4'b1100 : 4'b1000;
															assign node53984 = (inp[9]) ? 4'b1000 : 4'b1100;
														assign node53987 = (inp[9]) ? node53993 : node53988;
															assign node53988 = (inp[4]) ? 4'b1110 : node53989;
																assign node53989 = (inp[3]) ? 4'b1010 : 4'b1000;
															assign node53993 = (inp[4]) ? 4'b1010 : 4'b1110;
													assign node53996 = (inp[0]) ? node54004 : node53997;
														assign node53997 = (inp[3]) ? node54001 : node53998;
															assign node53998 = (inp[9]) ? 4'b1110 : 4'b1000;
															assign node54001 = (inp[9]) ? 4'b1010 : 4'b1110;
														assign node54004 = (inp[9]) ? node54010 : node54005;
															assign node54005 = (inp[4]) ? 4'b1100 : node54006;
																assign node54006 = (inp[3]) ? 4'b1000 : 4'b1010;
															assign node54010 = (inp[4]) ? 4'b1000 : 4'b1100;
												assign node54013 = (inp[15]) ? node54027 : node54014;
													assign node54014 = (inp[0]) ? node54022 : node54015;
														assign node54015 = (inp[9]) ? node54019 : node54016;
															assign node54016 = (inp[4]) ? 4'b1100 : 4'b1000;
															assign node54019 = (inp[4]) ? 4'b1000 : 4'b1100;
														assign node54022 = (inp[4]) ? node54024 : 4'b1110;
															assign node54024 = (inp[9]) ? 4'b1010 : 4'b1110;
													assign node54027 = (inp[0]) ? node54035 : node54028;
														assign node54028 = (inp[4]) ? node54032 : node54029;
															assign node54029 = (inp[9]) ? 4'b1110 : 4'b1010;
															assign node54032 = (inp[9]) ? 4'b1010 : 4'b1110;
														assign node54035 = (inp[4]) ? node54041 : node54036;
															assign node54036 = (inp[9]) ? 4'b1100 : node54037;
																assign node54037 = (inp[3]) ? 4'b1000 : 4'b1010;
															assign node54041 = (inp[9]) ? 4'b1000 : 4'b1100;
											assign node54044 = (inp[14]) ? node54078 : node54045;
												assign node54045 = (inp[0]) ? node54061 : node54046;
													assign node54046 = (inp[15]) ? node54056 : node54047;
														assign node54047 = (inp[9]) ? node54053 : node54048;
															assign node54048 = (inp[4]) ? 4'b1100 : node54049;
																assign node54049 = (inp[3]) ? 4'b1000 : 4'b1010;
															assign node54053 = (inp[4]) ? 4'b1000 : 4'b1100;
														assign node54056 = (inp[4]) ? 4'b1110 : node54057;
															assign node54057 = (inp[9]) ? 4'b1110 : 4'b1010;
													assign node54061 = (inp[15]) ? node54069 : node54062;
														assign node54062 = (inp[4]) ? node54066 : node54063;
															assign node54063 = (inp[3]) ? 4'b1010 : 4'b1000;
															assign node54066 = (inp[9]) ? 4'b1010 : 4'b1110;
														assign node54069 = (inp[9]) ? node54075 : node54070;
															assign node54070 = (inp[3]) ? node54072 : 4'b1010;
																assign node54072 = (inp[4]) ? 4'b1100 : 4'b1000;
															assign node54075 = (inp[4]) ? 4'b1000 : 4'b1100;
												assign node54078 = (inp[15]) ? node54098 : node54079;
													assign node54079 = (inp[0]) ? node54089 : node54080;
														assign node54080 = (inp[4]) ? node54086 : node54081;
															assign node54081 = (inp[9]) ? 4'b1100 : node54082;
																assign node54082 = (inp[3]) ? 4'b1000 : 4'b1010;
															assign node54086 = (inp[9]) ? 4'b1000 : 4'b1100;
														assign node54089 = (inp[3]) ? 4'b1010 : node54090;
															assign node54090 = (inp[9]) ? node54094 : node54091;
																assign node54091 = (inp[4]) ? 4'b1110 : 4'b1000;
																assign node54094 = (inp[4]) ? 4'b1010 : 4'b1110;
													assign node54098 = (inp[0]) ? node54106 : node54099;
														assign node54099 = (inp[9]) ? node54103 : node54100;
															assign node54100 = (inp[3]) ? 4'b1010 : 4'b1000;
															assign node54103 = (inp[4]) ? 4'b1010 : 4'b1110;
														assign node54106 = (inp[4]) ? node54110 : node54107;
															assign node54107 = (inp[9]) ? 4'b1100 : 4'b1010;
															assign node54110 = (inp[9]) ? 4'b1000 : 4'b1100;
					assign node54113 = (inp[8]) ? node56183 : node54114;
						assign node54114 = (inp[7]) ? node55210 : node54115;
							assign node54115 = (inp[14]) ? node54641 : node54116;
								assign node54116 = (inp[2]) ? node54410 : node54117;
									assign node54117 = (inp[3]) ? node54269 : node54118;
										assign node54118 = (inp[12]) ? node54212 : node54119;
											assign node54119 = (inp[5]) ? node54169 : node54120;
												assign node54120 = (inp[9]) ? node54144 : node54121;
													assign node54121 = (inp[10]) ? node54135 : node54122;
														assign node54122 = (inp[4]) ? node54128 : node54123;
															assign node54123 = (inp[0]) ? 4'b1101 : node54124;
																assign node54124 = (inp[15]) ? 4'b1101 : 4'b1111;
															assign node54128 = (inp[15]) ? node54132 : node54129;
																assign node54129 = (inp[0]) ? 4'b1001 : 4'b1011;
																assign node54132 = (inp[0]) ? 4'b1011 : 4'b1001;
														assign node54135 = (inp[4]) ? 4'b1101 : node54136;
															assign node54136 = (inp[15]) ? node54140 : node54137;
																assign node54137 = (inp[0]) ? 4'b1001 : 4'b1011;
																assign node54140 = (inp[0]) ? 4'b1011 : 4'b1001;
													assign node54144 = (inp[0]) ? node54154 : node54145;
														assign node54145 = (inp[15]) ? 4'b1101 : node54146;
															assign node54146 = (inp[4]) ? node54150 : node54147;
																assign node54147 = (inp[10]) ? 4'b1111 : 4'b1011;
																assign node54150 = (inp[10]) ? 4'b1011 : 4'b1111;
														assign node54154 = (inp[15]) ? node54162 : node54155;
															assign node54155 = (inp[10]) ? node54159 : node54156;
																assign node54156 = (inp[4]) ? 4'b1101 : 4'b1001;
																assign node54159 = (inp[4]) ? 4'b1001 : 4'b1101;
															assign node54162 = (inp[10]) ? node54166 : node54163;
																assign node54163 = (inp[4]) ? 4'b1111 : 4'b1011;
																assign node54166 = (inp[4]) ? 4'b1011 : 4'b1111;
												assign node54169 = (inp[9]) ? node54191 : node54170;
													assign node54170 = (inp[0]) ? node54178 : node54171;
														assign node54171 = (inp[4]) ? node54175 : node54172;
															assign node54172 = (inp[15]) ? 4'b1101 : 4'b1111;
															assign node54175 = (inp[15]) ? 4'b1001 : 4'b1101;
														assign node54178 = (inp[15]) ? node54184 : node54179;
															assign node54179 = (inp[4]) ? 4'b1111 : node54180;
																assign node54180 = (inp[10]) ? 4'b1001 : 4'b1101;
															assign node54184 = (inp[10]) ? node54188 : node54185;
																assign node54185 = (inp[4]) ? 4'b1011 : 4'b1111;
																assign node54188 = (inp[4]) ? 4'b1101 : 4'b1011;
													assign node54191 = (inp[0]) ? node54203 : node54192;
														assign node54192 = (inp[4]) ? node54200 : node54193;
															assign node54193 = (inp[10]) ? node54197 : node54194;
																assign node54194 = (inp[15]) ? 4'b1001 : 4'b1011;
																assign node54197 = (inp[15]) ? 4'b1111 : 4'b1101;
															assign node54200 = (inp[10]) ? 4'b1001 : 4'b1101;
														assign node54203 = (inp[15]) ? node54207 : node54204;
															assign node54204 = (inp[4]) ? 4'b1111 : 4'b1001;
															assign node54207 = (inp[4]) ? node54209 : 4'b1101;
																assign node54209 = (inp[10]) ? 4'b1001 : 4'b1101;
											assign node54212 = (inp[9]) ? node54240 : node54213;
												assign node54213 = (inp[4]) ? node54225 : node54214;
													assign node54214 = (inp[10]) ? node54220 : node54215;
														assign node54215 = (inp[0]) ? node54217 : 4'b1001;
															assign node54217 = (inp[15]) ? 4'b1011 : 4'b1001;
														assign node54220 = (inp[15]) ? node54222 : 4'b1011;
															assign node54222 = (inp[0]) ? 4'b1011 : 4'b1001;
													assign node54225 = (inp[15]) ? node54233 : node54226;
														assign node54226 = (inp[0]) ? node54230 : node54227;
															assign node54227 = (inp[5]) ? 4'b1101 : 4'b1111;
															assign node54230 = (inp[5]) ? 4'b1111 : 4'b1101;
														assign node54233 = (inp[0]) ? node54237 : node54234;
															assign node54234 = (inp[5]) ? 4'b1111 : 4'b1101;
															assign node54237 = (inp[5]) ? 4'b1101 : 4'b1111;
												assign node54240 = (inp[4]) ? node54256 : node54241;
													assign node54241 = (inp[5]) ? node54249 : node54242;
														assign node54242 = (inp[15]) ? node54246 : node54243;
															assign node54243 = (inp[0]) ? 4'b1101 : 4'b1111;
															assign node54246 = (inp[0]) ? 4'b1111 : 4'b1101;
														assign node54249 = (inp[15]) ? node54253 : node54250;
															assign node54250 = (inp[0]) ? 4'b1111 : 4'b1101;
															assign node54253 = (inp[0]) ? 4'b1101 : 4'b1111;
													assign node54256 = (inp[0]) ? node54264 : node54257;
														assign node54257 = (inp[15]) ? node54261 : node54258;
															assign node54258 = (inp[5]) ? 4'b1001 : 4'b1011;
															assign node54261 = (inp[5]) ? 4'b1011 : 4'b1001;
														assign node54264 = (inp[5]) ? 4'b1011 : node54265;
															assign node54265 = (inp[15]) ? 4'b1011 : 4'b1001;
										assign node54269 = (inp[15]) ? node54335 : node54270;
											assign node54270 = (inp[0]) ? node54300 : node54271;
												assign node54271 = (inp[5]) ? node54285 : node54272;
													assign node54272 = (inp[4]) ? node54282 : node54273;
														assign node54273 = (inp[9]) ? node54277 : node54274;
															assign node54274 = (inp[12]) ? 4'b1011 : 4'b1111;
															assign node54277 = (inp[12]) ? 4'b1101 : node54278;
																assign node54278 = (inp[10]) ? 4'b1101 : 4'b1011;
														assign node54282 = (inp[9]) ? 4'b1001 : 4'b1101;
													assign node54285 = (inp[10]) ? node54297 : node54286;
														assign node54286 = (inp[12]) ? node54292 : node54287;
															assign node54287 = (inp[9]) ? node54289 : 4'b1101;
																assign node54289 = (inp[4]) ? 4'b1101 : 4'b1001;
															assign node54292 = (inp[4]) ? node54294 : 4'b1001;
																assign node54294 = (inp[9]) ? 4'b1001 : 4'b1101;
														assign node54297 = (inp[12]) ? 4'b1101 : 4'b1001;
												assign node54300 = (inp[5]) ? node54314 : node54301;
													assign node54301 = (inp[10]) ? node54309 : node54302;
														assign node54302 = (inp[9]) ? 4'b1011 : node54303;
															assign node54303 = (inp[4]) ? node54305 : 4'b1001;
																assign node54305 = (inp[12]) ? 4'b1111 : 4'b1001;
														assign node54309 = (inp[4]) ? node54311 : 4'b1111;
															assign node54311 = (inp[9]) ? 4'b1011 : 4'b1111;
													assign node54314 = (inp[4]) ? node54326 : node54315;
														assign node54315 = (inp[9]) ? node54321 : node54316;
															assign node54316 = (inp[12]) ? 4'b1011 : node54317;
																assign node54317 = (inp[10]) ? 4'b1011 : 4'b1111;
															assign node54321 = (inp[12]) ? 4'b1111 : node54322;
																assign node54322 = (inp[10]) ? 4'b1111 : 4'b1011;
														assign node54326 = (inp[9]) ? node54332 : node54327;
															assign node54327 = (inp[10]) ? 4'b1111 : node54328;
																assign node54328 = (inp[12]) ? 4'b1111 : 4'b1011;
															assign node54332 = (inp[10]) ? 4'b1011 : 4'b1111;
											assign node54335 = (inp[0]) ? node54375 : node54336;
												assign node54336 = (inp[5]) ? node54352 : node54337;
													assign node54337 = (inp[9]) ? node54343 : node54338;
														assign node54338 = (inp[4]) ? node54340 : 4'b1001;
															assign node54340 = (inp[12]) ? 4'b1111 : 4'b1001;
														assign node54343 = (inp[4]) ? node54347 : node54344;
															assign node54344 = (inp[12]) ? 4'b1111 : 4'b1001;
															assign node54347 = (inp[10]) ? 4'b1011 : node54348;
																assign node54348 = (inp[12]) ? 4'b1011 : 4'b1111;
													assign node54352 = (inp[10]) ? node54364 : node54353;
														assign node54353 = (inp[4]) ? node54359 : node54354;
															assign node54354 = (inp[9]) ? node54356 : 4'b1011;
																assign node54356 = (inp[12]) ? 4'b1111 : 4'b1011;
															assign node54359 = (inp[9]) ? node54361 : 4'b1111;
																assign node54361 = (inp[12]) ? 4'b1011 : 4'b1111;
														assign node54364 = (inp[12]) ? node54370 : node54365;
															assign node54365 = (inp[4]) ? node54367 : 4'b1011;
																assign node54367 = (inp[9]) ? 4'b1011 : 4'b1111;
															assign node54370 = (inp[9]) ? node54372 : 4'b1011;
																assign node54372 = (inp[4]) ? 4'b1011 : 4'b1111;
												assign node54375 = (inp[5]) ? node54397 : node54376;
													assign node54376 = (inp[9]) ? node54386 : node54377;
														assign node54377 = (inp[4]) ? node54383 : node54378;
															assign node54378 = (inp[12]) ? 4'b1011 : node54379;
																assign node54379 = (inp[10]) ? 4'b1011 : 4'b1111;
															assign node54383 = (inp[12]) ? 4'b1101 : 4'b1011;
														assign node54386 = (inp[4]) ? node54392 : node54387;
															assign node54387 = (inp[10]) ? 4'b1101 : node54388;
																assign node54388 = (inp[12]) ? 4'b1101 : 4'b1011;
															assign node54392 = (inp[12]) ? 4'b1001 : node54393;
																assign node54393 = (inp[10]) ? 4'b1001 : 4'b1101;
													assign node54397 = (inp[10]) ? node54401 : node54398;
														assign node54398 = (inp[12]) ? 4'b1001 : 4'b1101;
														assign node54401 = (inp[12]) ? node54403 : 4'b1001;
															assign node54403 = (inp[9]) ? node54407 : node54404;
																assign node54404 = (inp[4]) ? 4'b1101 : 4'b1001;
																assign node54407 = (inp[4]) ? 4'b1001 : 4'b1101;
									assign node54410 = (inp[4]) ? node54528 : node54411;
										assign node54411 = (inp[9]) ? node54473 : node54412;
											assign node54412 = (inp[12]) ? node54450 : node54413;
												assign node54413 = (inp[10]) ? node54437 : node54414;
													assign node54414 = (inp[15]) ? node54426 : node54415;
														assign node54415 = (inp[0]) ? node54421 : node54416;
															assign node54416 = (inp[3]) ? node54418 : 4'b1110;
																assign node54418 = (inp[5]) ? 4'b1100 : 4'b1110;
															assign node54421 = (inp[3]) ? node54423 : 4'b1100;
																assign node54423 = (inp[5]) ? 4'b1110 : 4'b1100;
														assign node54426 = (inp[0]) ? node54432 : node54427;
															assign node54427 = (inp[5]) ? node54429 : 4'b1100;
																assign node54429 = (inp[3]) ? 4'b1110 : 4'b1100;
															assign node54432 = (inp[3]) ? node54434 : 4'b1110;
																assign node54434 = (inp[5]) ? 4'b1100 : 4'b1110;
													assign node54437 = (inp[15]) ? node54443 : node54438;
														assign node54438 = (inp[5]) ? 4'b1000 : node54439;
															assign node54439 = (inp[0]) ? 4'b1000 : 4'b1010;
														assign node54443 = (inp[3]) ? node54445 : 4'b1010;
															assign node54445 = (inp[0]) ? node54447 : 4'b1000;
																assign node54447 = (inp[5]) ? 4'b1000 : 4'b1010;
												assign node54450 = (inp[0]) ? node54462 : node54451;
													assign node54451 = (inp[5]) ? node54455 : node54452;
														assign node54452 = (inp[15]) ? 4'b1000 : 4'b1010;
														assign node54455 = (inp[3]) ? node54459 : node54456;
															assign node54456 = (inp[15]) ? 4'b1000 : 4'b1010;
															assign node54459 = (inp[15]) ? 4'b1010 : 4'b1000;
													assign node54462 = (inp[15]) ? node54468 : node54463;
														assign node54463 = (inp[3]) ? node54465 : 4'b1000;
															assign node54465 = (inp[5]) ? 4'b1010 : 4'b1000;
														assign node54468 = (inp[5]) ? node54470 : 4'b1010;
															assign node54470 = (inp[3]) ? 4'b1000 : 4'b1010;
											assign node54473 = (inp[12]) ? node54505 : node54474;
												assign node54474 = (inp[10]) ? node54490 : node54475;
													assign node54475 = (inp[15]) ? node54481 : node54476;
														assign node54476 = (inp[0]) ? node54478 : 4'b1010;
															assign node54478 = (inp[3]) ? 4'b1010 : 4'b1000;
														assign node54481 = (inp[5]) ? node54485 : node54482;
															assign node54482 = (inp[0]) ? 4'b1010 : 4'b1000;
															assign node54485 = (inp[3]) ? node54487 : 4'b1000;
																assign node54487 = (inp[0]) ? 4'b1000 : 4'b1010;
													assign node54490 = (inp[0]) ? node54500 : node54491;
														assign node54491 = (inp[15]) ? node54497 : node54492;
															assign node54492 = (inp[5]) ? 4'b1100 : node54493;
																assign node54493 = (inp[3]) ? 4'b1100 : 4'b1110;
															assign node54497 = (inp[5]) ? 4'b1110 : 4'b1100;
														assign node54500 = (inp[3]) ? node54502 : 4'b1110;
															assign node54502 = (inp[15]) ? 4'b1100 : 4'b1110;
												assign node54505 = (inp[0]) ? node54517 : node54506;
													assign node54506 = (inp[15]) ? node54512 : node54507;
														assign node54507 = (inp[5]) ? 4'b1100 : node54508;
															assign node54508 = (inp[3]) ? 4'b1100 : 4'b1110;
														assign node54512 = (inp[5]) ? 4'b1110 : node54513;
															assign node54513 = (inp[3]) ? 4'b1110 : 4'b1100;
													assign node54517 = (inp[15]) ? node54523 : node54518;
														assign node54518 = (inp[3]) ? 4'b1110 : node54519;
															assign node54519 = (inp[5]) ? 4'b1110 : 4'b1100;
														assign node54523 = (inp[5]) ? 4'b1100 : node54524;
															assign node54524 = (inp[3]) ? 4'b1100 : 4'b1110;
										assign node54528 = (inp[9]) ? node54580 : node54529;
											assign node54529 = (inp[12]) ? node54563 : node54530;
												assign node54530 = (inp[10]) ? node54552 : node54531;
													assign node54531 = (inp[3]) ? node54537 : node54532;
														assign node54532 = (inp[15]) ? node54534 : 4'b1010;
															assign node54534 = (inp[0]) ? 4'b1010 : 4'b1000;
														assign node54537 = (inp[5]) ? node54545 : node54538;
															assign node54538 = (inp[15]) ? node54542 : node54539;
																assign node54539 = (inp[0]) ? 4'b1000 : 4'b1010;
																assign node54542 = (inp[0]) ? 4'b1010 : 4'b1000;
															assign node54545 = (inp[15]) ? node54549 : node54546;
																assign node54546 = (inp[0]) ? 4'b1010 : 4'b1000;
																assign node54549 = (inp[0]) ? 4'b1000 : 4'b1010;
													assign node54552 = (inp[0]) ? node54556 : node54553;
														assign node54553 = (inp[15]) ? 4'b1110 : 4'b1100;
														assign node54556 = (inp[3]) ? node54560 : node54557;
															assign node54557 = (inp[15]) ? 4'b1110 : 4'b1100;
															assign node54560 = (inp[15]) ? 4'b1100 : 4'b1110;
												assign node54563 = (inp[0]) ? node54573 : node54564;
													assign node54564 = (inp[15]) ? node54568 : node54565;
														assign node54565 = (inp[10]) ? 4'b1100 : 4'b1110;
														assign node54568 = (inp[3]) ? 4'b1110 : node54569;
															assign node54569 = (inp[5]) ? 4'b1110 : 4'b1100;
													assign node54573 = (inp[15]) ? 4'b1100 : node54574;
														assign node54574 = (inp[3]) ? 4'b1110 : node54575;
															assign node54575 = (inp[5]) ? 4'b1110 : 4'b1100;
											assign node54580 = (inp[10]) ? node54612 : node54581;
												assign node54581 = (inp[12]) ? node54599 : node54582;
													assign node54582 = (inp[15]) ? node54588 : node54583;
														assign node54583 = (inp[0]) ? node54585 : 4'b1100;
															assign node54585 = (inp[3]) ? 4'b1110 : 4'b1100;
														assign node54588 = (inp[0]) ? node54594 : node54589;
															assign node54589 = (inp[5]) ? 4'b1110 : node54590;
																assign node54590 = (inp[3]) ? 4'b1110 : 4'b1100;
															assign node54594 = (inp[5]) ? 4'b1100 : node54595;
																assign node54595 = (inp[3]) ? 4'b1100 : 4'b1110;
													assign node54599 = (inp[5]) ? node54607 : node54600;
														assign node54600 = (inp[15]) ? 4'b1010 : node54601;
															assign node54601 = (inp[3]) ? node54603 : 4'b1000;
																assign node54603 = (inp[0]) ? 4'b1010 : 4'b1000;
														assign node54607 = (inp[15]) ? 4'b1000 : node54608;
															assign node54608 = (inp[0]) ? 4'b1010 : 4'b1000;
												assign node54612 = (inp[3]) ? node54634 : node54613;
													assign node54613 = (inp[5]) ? node54627 : node54614;
														assign node54614 = (inp[12]) ? node54622 : node54615;
															assign node54615 = (inp[0]) ? node54619 : node54616;
																assign node54616 = (inp[15]) ? 4'b1000 : 4'b1010;
																assign node54619 = (inp[15]) ? 4'b1010 : 4'b1000;
															assign node54622 = (inp[0]) ? 4'b1000 : node54623;
																assign node54623 = (inp[15]) ? 4'b1000 : 4'b1010;
														assign node54627 = (inp[0]) ? node54631 : node54628;
															assign node54628 = (inp[15]) ? 4'b1010 : 4'b1000;
															assign node54631 = (inp[15]) ? 4'b1000 : 4'b1010;
													assign node54634 = (inp[15]) ? node54638 : node54635;
														assign node54635 = (inp[0]) ? 4'b1010 : 4'b1000;
														assign node54638 = (inp[0]) ? 4'b1000 : 4'b1010;
								assign node54641 = (inp[2]) ? node54953 : node54642;
									assign node54642 = (inp[5]) ? node54790 : node54643;
										assign node54643 = (inp[3]) ? node54729 : node54644;
											assign node54644 = (inp[12]) ? node54692 : node54645;
												assign node54645 = (inp[4]) ? node54673 : node54646;
													assign node54646 = (inp[10]) ? node54658 : node54647;
														assign node54647 = (inp[9]) ? node54651 : node54648;
															assign node54648 = (inp[15]) ? 4'b1100 : 4'b1110;
															assign node54651 = (inp[15]) ? node54655 : node54652;
																assign node54652 = (inp[0]) ? 4'b1000 : 4'b1010;
																assign node54655 = (inp[0]) ? 4'b1010 : 4'b1000;
														assign node54658 = (inp[9]) ? node54666 : node54659;
															assign node54659 = (inp[15]) ? node54663 : node54660;
																assign node54660 = (inp[0]) ? 4'b1000 : 4'b1010;
																assign node54663 = (inp[0]) ? 4'b1010 : 4'b1000;
															assign node54666 = (inp[15]) ? node54670 : node54667;
																assign node54667 = (inp[0]) ? 4'b1100 : 4'b1110;
																assign node54670 = (inp[0]) ? 4'b1110 : 4'b1100;
													assign node54673 = (inp[9]) ? node54681 : node54674;
														assign node54674 = (inp[10]) ? node54676 : 4'b1010;
															assign node54676 = (inp[15]) ? 4'b1110 : node54677;
																assign node54677 = (inp[0]) ? 4'b1100 : 4'b1110;
														assign node54681 = (inp[10]) ? node54687 : node54682;
															assign node54682 = (inp[0]) ? 4'b1100 : node54683;
																assign node54683 = (inp[15]) ? 4'b1100 : 4'b1110;
															assign node54687 = (inp[0]) ? 4'b1010 : node54688;
																assign node54688 = (inp[15]) ? 4'b1000 : 4'b1010;
												assign node54692 = (inp[9]) ? node54708 : node54693;
													assign node54693 = (inp[4]) ? node54701 : node54694;
														assign node54694 = (inp[0]) ? node54698 : node54695;
															assign node54695 = (inp[15]) ? 4'b1000 : 4'b1010;
															assign node54698 = (inp[15]) ? 4'b1010 : 4'b1000;
														assign node54701 = (inp[0]) ? node54705 : node54702;
															assign node54702 = (inp[15]) ? 4'b1100 : 4'b1110;
															assign node54705 = (inp[15]) ? 4'b1110 : 4'b1100;
													assign node54708 = (inp[4]) ? node54716 : node54709;
														assign node54709 = (inp[15]) ? node54713 : node54710;
															assign node54710 = (inp[0]) ? 4'b1100 : 4'b1110;
															assign node54713 = (inp[0]) ? 4'b1110 : 4'b1100;
														assign node54716 = (inp[10]) ? node54722 : node54717;
															assign node54717 = (inp[15]) ? 4'b1000 : node54718;
																assign node54718 = (inp[0]) ? 4'b1000 : 4'b1010;
															assign node54722 = (inp[15]) ? node54726 : node54723;
																assign node54723 = (inp[0]) ? 4'b1000 : 4'b1010;
																assign node54726 = (inp[0]) ? 4'b1010 : 4'b1000;
											assign node54729 = (inp[15]) ? node54753 : node54730;
												assign node54730 = (inp[0]) ? node54738 : node54731;
													assign node54731 = (inp[9]) ? node54735 : node54732;
														assign node54732 = (inp[4]) ? 4'b1100 : 4'b1010;
														assign node54735 = (inp[4]) ? 4'b1000 : 4'b1100;
													assign node54738 = (inp[9]) ? node54746 : node54739;
														assign node54739 = (inp[4]) ? node54743 : node54740;
															assign node54740 = (inp[12]) ? 4'b1000 : 4'b1100;
															assign node54743 = (inp[12]) ? 4'b1110 : 4'b1000;
														assign node54746 = (inp[4]) ? node54748 : 4'b1110;
															assign node54748 = (inp[10]) ? 4'b1010 : node54749;
																assign node54749 = (inp[12]) ? 4'b1010 : 4'b1110;
												assign node54753 = (inp[0]) ? node54773 : node54754;
													assign node54754 = (inp[10]) ? node54768 : node54755;
														assign node54755 = (inp[12]) ? node54763 : node54756;
															assign node54756 = (inp[9]) ? node54760 : node54757;
																assign node54757 = (inp[4]) ? 4'b1000 : 4'b1100;
																assign node54760 = (inp[4]) ? 4'b1110 : 4'b1000;
															assign node54763 = (inp[4]) ? node54765 : 4'b1110;
																assign node54765 = (inp[9]) ? 4'b1010 : 4'b1110;
														assign node54768 = (inp[4]) ? node54770 : 4'b1110;
															assign node54770 = (inp[9]) ? 4'b1010 : 4'b1110;
													assign node54773 = (inp[9]) ? node54783 : node54774;
														assign node54774 = (inp[4]) ? node54778 : node54775;
															assign node54775 = (inp[12]) ? 4'b1010 : 4'b1110;
															assign node54778 = (inp[10]) ? 4'b1100 : node54779;
																assign node54779 = (inp[12]) ? 4'b1100 : 4'b1010;
														assign node54783 = (inp[4]) ? node54787 : node54784;
															assign node54784 = (inp[10]) ? 4'b1100 : 4'b1010;
															assign node54787 = (inp[12]) ? 4'b1000 : 4'b1100;
										assign node54790 = (inp[10]) ? node54872 : node54791;
											assign node54791 = (inp[4]) ? node54837 : node54792;
												assign node54792 = (inp[0]) ? node54808 : node54793;
													assign node54793 = (inp[15]) ? node54803 : node54794;
														assign node54794 = (inp[9]) ? node54800 : node54795;
															assign node54795 = (inp[12]) ? 4'b1010 : node54796;
																assign node54796 = (inp[3]) ? 4'b1100 : 4'b1110;
															assign node54800 = (inp[12]) ? 4'b1100 : 4'b1000;
														assign node54803 = (inp[9]) ? 4'b1110 : node54804;
															assign node54804 = (inp[3]) ? 4'b1110 : 4'b1100;
													assign node54808 = (inp[15]) ? node54824 : node54809;
														assign node54809 = (inp[3]) ? node54817 : node54810;
															assign node54810 = (inp[9]) ? node54814 : node54811;
																assign node54811 = (inp[12]) ? 4'b1000 : 4'b1100;
																assign node54814 = (inp[12]) ? 4'b1110 : 4'b1000;
															assign node54817 = (inp[9]) ? node54821 : node54818;
																assign node54818 = (inp[12]) ? 4'b1010 : 4'b1110;
																assign node54821 = (inp[12]) ? 4'b1110 : 4'b1010;
														assign node54824 = (inp[3]) ? node54832 : node54825;
															assign node54825 = (inp[9]) ? node54829 : node54826;
																assign node54826 = (inp[12]) ? 4'b1010 : 4'b1110;
																assign node54829 = (inp[12]) ? 4'b1100 : 4'b1010;
															assign node54832 = (inp[9]) ? 4'b1100 : node54833;
																assign node54833 = (inp[12]) ? 4'b1000 : 4'b1100;
												assign node54837 = (inp[12]) ? node54857 : node54838;
													assign node54838 = (inp[9]) ? node54852 : node54839;
														assign node54839 = (inp[0]) ? node54847 : node54840;
															assign node54840 = (inp[15]) ? node54844 : node54841;
																assign node54841 = (inp[3]) ? 4'b1000 : 4'b1010;
																assign node54844 = (inp[3]) ? 4'b1010 : 4'b1000;
															assign node54847 = (inp[3]) ? node54849 : 4'b1010;
																assign node54849 = (inp[15]) ? 4'b1000 : 4'b1010;
														assign node54852 = (inp[3]) ? node54854 : 4'b1100;
															assign node54854 = (inp[0]) ? 4'b1100 : 4'b1110;
													assign node54857 = (inp[9]) ? node54865 : node54858;
														assign node54858 = (inp[15]) ? node54862 : node54859;
															assign node54859 = (inp[0]) ? 4'b1110 : 4'b1100;
															assign node54862 = (inp[0]) ? 4'b1100 : 4'b1110;
														assign node54865 = (inp[3]) ? node54867 : 4'b1000;
															assign node54867 = (inp[0]) ? node54869 : 4'b1010;
																assign node54869 = (inp[15]) ? 4'b1000 : 4'b1010;
											assign node54872 = (inp[12]) ? node54916 : node54873;
												assign node54873 = (inp[4]) ? node54893 : node54874;
													assign node54874 = (inp[9]) ? node54884 : node54875;
														assign node54875 = (inp[0]) ? node54877 : 4'b1000;
															assign node54877 = (inp[3]) ? node54881 : node54878;
																assign node54878 = (inp[15]) ? 4'b1010 : 4'b1000;
																assign node54881 = (inp[15]) ? 4'b1000 : 4'b1010;
														assign node54884 = (inp[3]) ? node54888 : node54885;
															assign node54885 = (inp[15]) ? 4'b1110 : 4'b1100;
															assign node54888 = (inp[15]) ? node54890 : 4'b1110;
																assign node54890 = (inp[0]) ? 4'b1100 : 4'b1110;
													assign node54893 = (inp[9]) ? node54909 : node54894;
														assign node54894 = (inp[3]) ? node54902 : node54895;
															assign node54895 = (inp[0]) ? node54899 : node54896;
																assign node54896 = (inp[15]) ? 4'b1110 : 4'b1100;
																assign node54899 = (inp[15]) ? 4'b1100 : 4'b1110;
															assign node54902 = (inp[0]) ? node54906 : node54903;
																assign node54903 = (inp[15]) ? 4'b1110 : 4'b1100;
																assign node54906 = (inp[15]) ? 4'b1100 : 4'b1110;
														assign node54909 = (inp[15]) ? node54913 : node54910;
															assign node54910 = (inp[0]) ? 4'b1010 : 4'b1000;
															assign node54913 = (inp[0]) ? 4'b1000 : 4'b1010;
												assign node54916 = (inp[0]) ? node54938 : node54917;
													assign node54917 = (inp[15]) ? node54929 : node54918;
														assign node54918 = (inp[3]) ? node54924 : node54919;
															assign node54919 = (inp[9]) ? node54921 : 4'b1010;
																assign node54921 = (inp[4]) ? 4'b1000 : 4'b1100;
															assign node54924 = (inp[4]) ? node54926 : 4'b1100;
																assign node54926 = (inp[9]) ? 4'b1000 : 4'b1100;
														assign node54929 = (inp[3]) ? node54933 : node54930;
															assign node54930 = (inp[4]) ? 4'b1010 : 4'b1000;
															assign node54933 = (inp[4]) ? node54935 : 4'b1010;
																assign node54935 = (inp[9]) ? 4'b1010 : 4'b1110;
													assign node54938 = (inp[15]) ? node54944 : node54939;
														assign node54939 = (inp[9]) ? node54941 : 4'b1000;
															assign node54941 = (inp[4]) ? 4'b1010 : 4'b1110;
														assign node54944 = (inp[4]) ? node54950 : node54945;
															assign node54945 = (inp[9]) ? 4'b1100 : node54946;
																assign node54946 = (inp[3]) ? 4'b1000 : 4'b1010;
															assign node54950 = (inp[9]) ? 4'b1000 : 4'b1100;
									assign node54953 = (inp[12]) ? node55107 : node54954;
										assign node54954 = (inp[4]) ? node55030 : node54955;
											assign node54955 = (inp[10]) ? node54997 : node54956;
												assign node54956 = (inp[9]) ? node54976 : node54957;
													assign node54957 = (inp[3]) ? node54963 : node54958;
														assign node54958 = (inp[0]) ? node54960 : 4'b1100;
															assign node54960 = (inp[15]) ? 4'b1110 : 4'b1100;
														assign node54963 = (inp[0]) ? node54971 : node54964;
															assign node54964 = (inp[5]) ? node54968 : node54965;
																assign node54965 = (inp[15]) ? 4'b1100 : 4'b1110;
																assign node54968 = (inp[15]) ? 4'b1110 : 4'b1100;
															assign node54971 = (inp[15]) ? node54973 : 4'b1110;
																assign node54973 = (inp[5]) ? 4'b1100 : 4'b1110;
													assign node54976 = (inp[0]) ? node54986 : node54977;
														assign node54977 = (inp[15]) ? node54981 : node54978;
															assign node54978 = (inp[3]) ? 4'b1000 : 4'b1010;
															assign node54981 = (inp[5]) ? node54983 : 4'b1000;
																assign node54983 = (inp[3]) ? 4'b1010 : 4'b1000;
														assign node54986 = (inp[15]) ? node54992 : node54987;
															assign node54987 = (inp[5]) ? node54989 : 4'b1000;
																assign node54989 = (inp[3]) ? 4'b1010 : 4'b1000;
															assign node54992 = (inp[5]) ? node54994 : 4'b1010;
																assign node54994 = (inp[3]) ? 4'b1000 : 4'b1010;
												assign node54997 = (inp[9]) ? node55015 : node54998;
													assign node54998 = (inp[0]) ? node55006 : node54999;
														assign node54999 = (inp[15]) ? node55003 : node55000;
															assign node55000 = (inp[5]) ? 4'b1000 : 4'b1010;
															assign node55003 = (inp[5]) ? 4'b1010 : 4'b1000;
														assign node55006 = (inp[15]) ? node55010 : node55007;
															assign node55007 = (inp[3]) ? 4'b1010 : 4'b1000;
															assign node55010 = (inp[5]) ? node55012 : 4'b1010;
																assign node55012 = (inp[3]) ? 4'b1000 : 4'b1010;
													assign node55015 = (inp[5]) ? 4'b1110 : node55016;
														assign node55016 = (inp[15]) ? node55022 : node55017;
															assign node55017 = (inp[3]) ? node55019 : 4'b1100;
																assign node55019 = (inp[0]) ? 4'b1110 : 4'b1100;
															assign node55022 = (inp[3]) ? node55026 : node55023;
																assign node55023 = (inp[0]) ? 4'b1110 : 4'b1100;
																assign node55026 = (inp[0]) ? 4'b1100 : 4'b1110;
											assign node55030 = (inp[3]) ? node55066 : node55031;
												assign node55031 = (inp[15]) ? node55055 : node55032;
													assign node55032 = (inp[0]) ? node55042 : node55033;
														assign node55033 = (inp[10]) ? node55037 : node55034;
															assign node55034 = (inp[9]) ? 4'b1110 : 4'b1010;
															assign node55037 = (inp[9]) ? 4'b1000 : node55038;
																assign node55038 = (inp[5]) ? 4'b1100 : 4'b1110;
														assign node55042 = (inp[5]) ? node55048 : node55043;
															assign node55043 = (inp[9]) ? node55045 : 4'b1000;
																assign node55045 = (inp[10]) ? 4'b1000 : 4'b1100;
															assign node55048 = (inp[10]) ? node55052 : node55049;
																assign node55049 = (inp[9]) ? 4'b1110 : 4'b1000;
																assign node55052 = (inp[9]) ? 4'b1010 : 4'b1110;
													assign node55055 = (inp[5]) ? node55059 : node55056;
														assign node55056 = (inp[0]) ? 4'b1110 : 4'b1100;
														assign node55059 = (inp[0]) ? node55063 : node55060;
															assign node55060 = (inp[10]) ? 4'b1010 : 4'b1110;
															assign node55063 = (inp[10]) ? 4'b1100 : 4'b1010;
												assign node55066 = (inp[0]) ? node55088 : node55067;
													assign node55067 = (inp[15]) ? node55077 : node55068;
														assign node55068 = (inp[10]) ? node55074 : node55069;
															assign node55069 = (inp[5]) ? node55071 : 4'b1010;
																assign node55071 = (inp[9]) ? 4'b1100 : 4'b1000;
															assign node55074 = (inp[9]) ? 4'b1000 : 4'b1100;
														assign node55077 = (inp[5]) ? node55081 : node55078;
															assign node55078 = (inp[9]) ? 4'b1110 : 4'b1000;
															assign node55081 = (inp[9]) ? node55085 : node55082;
																assign node55082 = (inp[10]) ? 4'b1110 : 4'b1010;
																assign node55085 = (inp[10]) ? 4'b1010 : 4'b1110;
													assign node55088 = (inp[15]) ? node55094 : node55089;
														assign node55089 = (inp[9]) ? node55091 : 4'b1110;
															assign node55091 = (inp[10]) ? 4'b1010 : 4'b1110;
														assign node55094 = (inp[5]) ? node55100 : node55095;
															assign node55095 = (inp[10]) ? 4'b1100 : node55096;
																assign node55096 = (inp[9]) ? 4'b1100 : 4'b1010;
															assign node55100 = (inp[9]) ? node55104 : node55101;
																assign node55101 = (inp[10]) ? 4'b1100 : 4'b1000;
																assign node55104 = (inp[10]) ? 4'b1000 : 4'b1100;
										assign node55107 = (inp[0]) ? node55157 : node55108;
											assign node55108 = (inp[15]) ? node55132 : node55109;
												assign node55109 = (inp[3]) ? node55123 : node55110;
													assign node55110 = (inp[5]) ? node55116 : node55111;
														assign node55111 = (inp[9]) ? 4'b1010 : node55112;
															assign node55112 = (inp[4]) ? 4'b1110 : 4'b1010;
														assign node55116 = (inp[9]) ? node55120 : node55117;
															assign node55117 = (inp[4]) ? 4'b1100 : 4'b1010;
															assign node55120 = (inp[4]) ? 4'b1000 : 4'b1100;
													assign node55123 = (inp[4]) ? node55129 : node55124;
														assign node55124 = (inp[9]) ? 4'b1100 : node55125;
															assign node55125 = (inp[5]) ? 4'b1000 : 4'b1010;
														assign node55129 = (inp[9]) ? 4'b1000 : 4'b1100;
												assign node55132 = (inp[5]) ? node55148 : node55133;
													assign node55133 = (inp[3]) ? node55141 : node55134;
														assign node55134 = (inp[4]) ? node55138 : node55135;
															assign node55135 = (inp[9]) ? 4'b1100 : 4'b1000;
															assign node55138 = (inp[9]) ? 4'b1000 : 4'b1100;
														assign node55141 = (inp[9]) ? node55145 : node55142;
															assign node55142 = (inp[4]) ? 4'b1110 : 4'b1000;
															assign node55145 = (inp[4]) ? 4'b1010 : 4'b1110;
													assign node55148 = (inp[4]) ? node55154 : node55149;
														assign node55149 = (inp[9]) ? 4'b1110 : node55150;
															assign node55150 = (inp[3]) ? 4'b1010 : 4'b1000;
														assign node55154 = (inp[9]) ? 4'b1010 : 4'b1110;
											assign node55157 = (inp[15]) ? node55181 : node55158;
												assign node55158 = (inp[5]) ? node55172 : node55159;
													assign node55159 = (inp[3]) ? node55167 : node55160;
														assign node55160 = (inp[4]) ? node55164 : node55161;
															assign node55161 = (inp[9]) ? 4'b1100 : 4'b1000;
															assign node55164 = (inp[9]) ? 4'b1000 : 4'b1100;
														assign node55167 = (inp[10]) ? node55169 : 4'b1110;
															assign node55169 = (inp[9]) ? 4'b1010 : 4'b1000;
													assign node55172 = (inp[9]) ? node55178 : node55173;
														assign node55173 = (inp[4]) ? 4'b1110 : node55174;
															assign node55174 = (inp[3]) ? 4'b1010 : 4'b1000;
														assign node55178 = (inp[4]) ? 4'b1010 : 4'b1110;
												assign node55181 = (inp[3]) ? node55195 : node55182;
													assign node55182 = (inp[5]) ? node55190 : node55183;
														assign node55183 = (inp[10]) ? node55185 : 4'b1010;
															assign node55185 = (inp[4]) ? 4'b1110 : node55186;
																assign node55186 = (inp[9]) ? 4'b1110 : 4'b1010;
														assign node55190 = (inp[4]) ? node55192 : 4'b1010;
															assign node55192 = (inp[9]) ? 4'b1000 : 4'b1100;
													assign node55195 = (inp[5]) ? node55203 : node55196;
														assign node55196 = (inp[9]) ? node55200 : node55197;
															assign node55197 = (inp[4]) ? 4'b1100 : 4'b1010;
															assign node55200 = (inp[4]) ? 4'b1000 : 4'b1100;
														assign node55203 = (inp[9]) ? node55207 : node55204;
															assign node55204 = (inp[4]) ? 4'b1100 : 4'b1000;
															assign node55207 = (inp[4]) ? 4'b1000 : 4'b1100;
							assign node55210 = (inp[2]) ? node55794 : node55211;
								assign node55211 = (inp[14]) ? node55471 : node55212;
									assign node55212 = (inp[4]) ? node55354 : node55213;
										assign node55213 = (inp[9]) ? node55287 : node55214;
											assign node55214 = (inp[10]) ? node55256 : node55215;
												assign node55215 = (inp[12]) ? node55237 : node55216;
													assign node55216 = (inp[3]) ? node55232 : node55217;
														assign node55217 = (inp[5]) ? node55225 : node55218;
															assign node55218 = (inp[15]) ? node55222 : node55219;
																assign node55219 = (inp[0]) ? 4'b1100 : 4'b1110;
																assign node55222 = (inp[0]) ? 4'b1110 : 4'b1100;
															assign node55225 = (inp[0]) ? node55229 : node55226;
																assign node55226 = (inp[15]) ? 4'b1100 : 4'b1110;
																assign node55229 = (inp[15]) ? 4'b1110 : 4'b1100;
														assign node55232 = (inp[15]) ? 4'b1110 : node55233;
															assign node55233 = (inp[5]) ? 4'b1110 : 4'b1100;
													assign node55237 = (inp[3]) ? node55247 : node55238;
														assign node55238 = (inp[5]) ? 4'b1000 : node55239;
															assign node55239 = (inp[15]) ? node55243 : node55240;
																assign node55240 = (inp[0]) ? 4'b1000 : 4'b1010;
																assign node55243 = (inp[0]) ? 4'b1010 : 4'b1000;
														assign node55247 = (inp[0]) ? 4'b1010 : node55248;
															assign node55248 = (inp[5]) ? node55252 : node55249;
																assign node55249 = (inp[15]) ? 4'b1000 : 4'b1010;
																assign node55252 = (inp[15]) ? 4'b1010 : 4'b1000;
												assign node55256 = (inp[5]) ? node55274 : node55257;
													assign node55257 = (inp[12]) ? node55267 : node55258;
														assign node55258 = (inp[3]) ? node55260 : 4'b1010;
															assign node55260 = (inp[15]) ? node55264 : node55261;
																assign node55261 = (inp[0]) ? 4'b1000 : 4'b1010;
																assign node55264 = (inp[0]) ? 4'b1010 : 4'b1000;
														assign node55267 = (inp[15]) ? node55271 : node55268;
															assign node55268 = (inp[0]) ? 4'b1000 : 4'b1010;
															assign node55271 = (inp[0]) ? 4'b1010 : 4'b1000;
													assign node55274 = (inp[3]) ? node55280 : node55275;
														assign node55275 = (inp[15]) ? node55277 : 4'b1000;
															assign node55277 = (inp[0]) ? 4'b1010 : 4'b1000;
														assign node55280 = (inp[15]) ? node55284 : node55281;
															assign node55281 = (inp[0]) ? 4'b1010 : 4'b1000;
															assign node55284 = (inp[0]) ? 4'b1000 : 4'b1010;
											assign node55287 = (inp[12]) ? node55331 : node55288;
												assign node55288 = (inp[10]) ? node55314 : node55289;
													assign node55289 = (inp[3]) ? node55299 : node55290;
														assign node55290 = (inp[5]) ? node55294 : node55291;
															assign node55291 = (inp[15]) ? 4'b1000 : 4'b1010;
															assign node55294 = (inp[15]) ? 4'b1010 : node55295;
																assign node55295 = (inp[0]) ? 4'b1000 : 4'b1010;
														assign node55299 = (inp[5]) ? node55307 : node55300;
															assign node55300 = (inp[15]) ? node55304 : node55301;
																assign node55301 = (inp[0]) ? 4'b1000 : 4'b1010;
																assign node55304 = (inp[0]) ? 4'b1010 : 4'b1000;
															assign node55307 = (inp[15]) ? node55311 : node55308;
																assign node55308 = (inp[0]) ? 4'b1010 : 4'b1000;
																assign node55311 = (inp[0]) ? 4'b1000 : 4'b1010;
													assign node55314 = (inp[3]) ? node55324 : node55315;
														assign node55315 = (inp[0]) ? node55317 : 4'b1110;
															assign node55317 = (inp[15]) ? node55321 : node55318;
																assign node55318 = (inp[5]) ? 4'b1110 : 4'b1100;
																assign node55321 = (inp[5]) ? 4'b1100 : 4'b1110;
														assign node55324 = (inp[0]) ? node55328 : node55325;
															assign node55325 = (inp[15]) ? 4'b1110 : 4'b1100;
															assign node55328 = (inp[15]) ? 4'b1100 : 4'b1110;
												assign node55331 = (inp[0]) ? node55343 : node55332;
													assign node55332 = (inp[15]) ? node55338 : node55333;
														assign node55333 = (inp[3]) ? 4'b1100 : node55334;
															assign node55334 = (inp[5]) ? 4'b1100 : 4'b1110;
														assign node55338 = (inp[5]) ? 4'b1110 : node55339;
															assign node55339 = (inp[3]) ? 4'b1110 : 4'b1100;
													assign node55343 = (inp[15]) ? node55349 : node55344;
														assign node55344 = (inp[3]) ? 4'b1110 : node55345;
															assign node55345 = (inp[5]) ? 4'b1110 : 4'b1100;
														assign node55349 = (inp[5]) ? 4'b1100 : node55350;
															assign node55350 = (inp[3]) ? 4'b1100 : 4'b1110;
										assign node55354 = (inp[9]) ? node55414 : node55355;
											assign node55355 = (inp[10]) ? node55391 : node55356;
												assign node55356 = (inp[12]) ? node55376 : node55357;
													assign node55357 = (inp[5]) ? node55365 : node55358;
														assign node55358 = (inp[15]) ? node55362 : node55359;
															assign node55359 = (inp[0]) ? 4'b1000 : 4'b1010;
															assign node55362 = (inp[0]) ? 4'b1010 : 4'b1000;
														assign node55365 = (inp[3]) ? node55371 : node55366;
															assign node55366 = (inp[0]) ? node55368 : 4'b1000;
																assign node55368 = (inp[15]) ? 4'b1010 : 4'b1000;
															assign node55371 = (inp[15]) ? node55373 : 4'b1010;
																assign node55373 = (inp[0]) ? 4'b1000 : 4'b1010;
													assign node55376 = (inp[5]) ? node55386 : node55377;
														assign node55377 = (inp[3]) ? node55379 : 4'b1110;
															assign node55379 = (inp[15]) ? node55383 : node55380;
																assign node55380 = (inp[0]) ? 4'b1110 : 4'b1100;
																assign node55383 = (inp[0]) ? 4'b1100 : 4'b1110;
														assign node55386 = (inp[15]) ? 4'b1100 : node55387;
															assign node55387 = (inp[0]) ? 4'b1110 : 4'b1100;
												assign node55391 = (inp[15]) ? node55403 : node55392;
													assign node55392 = (inp[0]) ? node55398 : node55393;
														assign node55393 = (inp[3]) ? 4'b1100 : node55394;
															assign node55394 = (inp[5]) ? 4'b1100 : 4'b1110;
														assign node55398 = (inp[5]) ? 4'b1110 : node55399;
															assign node55399 = (inp[3]) ? 4'b1110 : 4'b1100;
													assign node55403 = (inp[0]) ? node55409 : node55404;
														assign node55404 = (inp[3]) ? 4'b1110 : node55405;
															assign node55405 = (inp[12]) ? 4'b1100 : 4'b1110;
														assign node55409 = (inp[3]) ? 4'b1100 : node55410;
															assign node55410 = (inp[5]) ? 4'b1100 : 4'b1110;
											assign node55414 = (inp[12]) ? node55448 : node55415;
												assign node55415 = (inp[10]) ? node55431 : node55416;
													assign node55416 = (inp[0]) ? node55422 : node55417;
														assign node55417 = (inp[3]) ? node55419 : 4'b1110;
															assign node55419 = (inp[15]) ? 4'b1110 : 4'b1100;
														assign node55422 = (inp[3]) ? node55428 : node55423;
															assign node55423 = (inp[15]) ? node55425 : 4'b1100;
																assign node55425 = (inp[5]) ? 4'b1100 : 4'b1110;
															assign node55428 = (inp[5]) ? 4'b1110 : 4'b1100;
													assign node55431 = (inp[5]) ? node55441 : node55432;
														assign node55432 = (inp[15]) ? node55434 : 4'b1000;
															assign node55434 = (inp[0]) ? node55438 : node55435;
																assign node55435 = (inp[3]) ? 4'b1010 : 4'b1000;
																assign node55438 = (inp[3]) ? 4'b1000 : 4'b1010;
														assign node55441 = (inp[15]) ? node55445 : node55442;
															assign node55442 = (inp[0]) ? 4'b1010 : 4'b1000;
															assign node55445 = (inp[0]) ? 4'b1000 : 4'b1010;
												assign node55448 = (inp[0]) ? node55460 : node55449;
													assign node55449 = (inp[15]) ? node55455 : node55450;
														assign node55450 = (inp[5]) ? 4'b1000 : node55451;
															assign node55451 = (inp[3]) ? 4'b1000 : 4'b1010;
														assign node55455 = (inp[3]) ? 4'b1010 : node55456;
															assign node55456 = (inp[5]) ? 4'b1010 : 4'b1000;
													assign node55460 = (inp[15]) ? node55466 : node55461;
														assign node55461 = (inp[5]) ? 4'b1010 : node55462;
															assign node55462 = (inp[3]) ? 4'b1010 : 4'b1000;
														assign node55466 = (inp[3]) ? 4'b1000 : node55467;
															assign node55467 = (inp[5]) ? 4'b1000 : 4'b1010;
									assign node55471 = (inp[0]) ? node55635 : node55472;
										assign node55472 = (inp[15]) ? node55558 : node55473;
											assign node55473 = (inp[3]) ? node55511 : node55474;
												assign node55474 = (inp[5]) ? node55496 : node55475;
													assign node55475 = (inp[12]) ? node55491 : node55476;
														assign node55476 = (inp[10]) ? node55484 : node55477;
															assign node55477 = (inp[9]) ? node55481 : node55478;
																assign node55478 = (inp[4]) ? 4'b0011 : 4'b0111;
																assign node55481 = (inp[4]) ? 4'b0111 : 4'b0011;
															assign node55484 = (inp[4]) ? node55488 : node55485;
																assign node55485 = (inp[9]) ? 4'b0111 : 4'b0011;
																assign node55488 = (inp[9]) ? 4'b0011 : 4'b0111;
														assign node55491 = (inp[4]) ? 4'b0011 : node55492;
															assign node55492 = (inp[9]) ? 4'b0111 : 4'b0011;
													assign node55496 = (inp[9]) ? node55506 : node55497;
														assign node55497 = (inp[4]) ? node55503 : node55498;
															assign node55498 = (inp[12]) ? 4'b0011 : node55499;
																assign node55499 = (inp[10]) ? 4'b0011 : 4'b0111;
															assign node55503 = (inp[12]) ? 4'b0101 : 4'b0011;
														assign node55506 = (inp[12]) ? 4'b0101 : node55507;
															assign node55507 = (inp[10]) ? 4'b0101 : 4'b0011;
												assign node55511 = (inp[5]) ? node55531 : node55512;
													assign node55512 = (inp[4]) ? node55522 : node55513;
														assign node55513 = (inp[9]) ? node55519 : node55514;
															assign node55514 = (inp[10]) ? 4'b0011 : node55515;
																assign node55515 = (inp[12]) ? 4'b0011 : 4'b0111;
															assign node55519 = (inp[10]) ? 4'b0101 : 4'b0011;
														assign node55522 = (inp[12]) ? node55528 : node55523;
															assign node55523 = (inp[9]) ? node55525 : 4'b0011;
																assign node55525 = (inp[10]) ? 4'b0001 : 4'b0101;
															assign node55528 = (inp[9]) ? 4'b0001 : 4'b0101;
													assign node55531 = (inp[10]) ? node55545 : node55532;
														assign node55532 = (inp[12]) ? node55538 : node55533;
															assign node55533 = (inp[4]) ? 4'b0001 : node55534;
																assign node55534 = (inp[9]) ? 4'b0001 : 4'b0101;
															assign node55538 = (inp[4]) ? node55542 : node55539;
																assign node55539 = (inp[9]) ? 4'b0101 : 4'b0001;
																assign node55542 = (inp[9]) ? 4'b0001 : 4'b0101;
														assign node55545 = (inp[12]) ? node55553 : node55546;
															assign node55546 = (inp[4]) ? node55550 : node55547;
																assign node55547 = (inp[9]) ? 4'b0101 : 4'b0001;
																assign node55550 = (inp[9]) ? 4'b0001 : 4'b0101;
															assign node55553 = (inp[9]) ? node55555 : 4'b0101;
																assign node55555 = (inp[4]) ? 4'b0001 : 4'b0101;
											assign node55558 = (inp[5]) ? node55592 : node55559;
												assign node55559 = (inp[3]) ? node55571 : node55560;
													assign node55560 = (inp[4]) ? node55564 : node55561;
														assign node55561 = (inp[9]) ? 4'b0101 : 4'b0001;
														assign node55564 = (inp[9]) ? node55566 : 4'b0101;
															assign node55566 = (inp[12]) ? 4'b0001 : node55567;
																assign node55567 = (inp[10]) ? 4'b0001 : 4'b0101;
													assign node55571 = (inp[4]) ? node55581 : node55572;
														assign node55572 = (inp[9]) ? node55578 : node55573;
															assign node55573 = (inp[12]) ? 4'b0001 : node55574;
																assign node55574 = (inp[10]) ? 4'b0001 : 4'b0101;
															assign node55578 = (inp[12]) ? 4'b0111 : 4'b0001;
														assign node55581 = (inp[9]) ? node55587 : node55582;
															assign node55582 = (inp[10]) ? 4'b0111 : node55583;
																assign node55583 = (inp[12]) ? 4'b0111 : 4'b0001;
															assign node55587 = (inp[10]) ? 4'b0011 : node55588;
																assign node55588 = (inp[12]) ? 4'b0011 : 4'b0111;
												assign node55592 = (inp[3]) ? node55612 : node55593;
													assign node55593 = (inp[4]) ? node55601 : node55594;
														assign node55594 = (inp[9]) ? node55596 : 4'b0001;
															assign node55596 = (inp[12]) ? 4'b0111 : node55597;
																assign node55597 = (inp[10]) ? 4'b0111 : 4'b0001;
														assign node55601 = (inp[9]) ? node55607 : node55602;
															assign node55602 = (inp[12]) ? 4'b0111 : node55603;
																assign node55603 = (inp[10]) ? 4'b0111 : 4'b0001;
															assign node55607 = (inp[12]) ? 4'b0011 : node55608;
																assign node55608 = (inp[10]) ? 4'b0011 : 4'b0111;
													assign node55612 = (inp[4]) ? node55624 : node55613;
														assign node55613 = (inp[9]) ? node55619 : node55614;
															assign node55614 = (inp[12]) ? 4'b0011 : node55615;
																assign node55615 = (inp[10]) ? 4'b0011 : 4'b0111;
															assign node55619 = (inp[10]) ? 4'b0111 : node55620;
																assign node55620 = (inp[12]) ? 4'b0111 : 4'b0011;
														assign node55624 = (inp[9]) ? node55630 : node55625;
															assign node55625 = (inp[12]) ? 4'b0111 : node55626;
																assign node55626 = (inp[10]) ? 4'b0111 : 4'b0011;
															assign node55630 = (inp[12]) ? 4'b0011 : node55631;
																assign node55631 = (inp[10]) ? 4'b0011 : 4'b0111;
										assign node55635 = (inp[12]) ? node55729 : node55636;
											assign node55636 = (inp[3]) ? node55678 : node55637;
												assign node55637 = (inp[15]) ? node55653 : node55638;
													assign node55638 = (inp[5]) ? node55644 : node55639;
														assign node55639 = (inp[10]) ? node55641 : 4'b0101;
															assign node55641 = (inp[4]) ? 4'b0001 : 4'b0101;
														assign node55644 = (inp[10]) ? 4'b0111 : node55645;
															assign node55645 = (inp[9]) ? node55649 : node55646;
																assign node55646 = (inp[4]) ? 4'b0001 : 4'b0101;
																assign node55649 = (inp[4]) ? 4'b0111 : 4'b0001;
													assign node55653 = (inp[5]) ? node55667 : node55654;
														assign node55654 = (inp[9]) ? node55660 : node55655;
															assign node55655 = (inp[10]) ? node55657 : 4'b0011;
																assign node55657 = (inp[4]) ? 4'b0111 : 4'b0011;
															assign node55660 = (inp[10]) ? node55664 : node55661;
																assign node55661 = (inp[4]) ? 4'b0111 : 4'b0011;
																assign node55664 = (inp[4]) ? 4'b0011 : 4'b0111;
														assign node55667 = (inp[10]) ? node55671 : node55668;
															assign node55668 = (inp[4]) ? 4'b0011 : 4'b0111;
															assign node55671 = (inp[9]) ? node55675 : node55672;
																assign node55672 = (inp[4]) ? 4'b0101 : 4'b0011;
																assign node55675 = (inp[4]) ? 4'b0001 : 4'b0101;
												assign node55678 = (inp[15]) ? node55704 : node55679;
													assign node55679 = (inp[5]) ? node55691 : node55680;
														assign node55680 = (inp[4]) ? node55686 : node55681;
															assign node55681 = (inp[9]) ? 4'b0001 : node55682;
																assign node55682 = (inp[10]) ? 4'b0001 : 4'b0101;
															assign node55686 = (inp[10]) ? 4'b0111 : node55687;
																assign node55687 = (inp[9]) ? 4'b0111 : 4'b0001;
														assign node55691 = (inp[9]) ? node55697 : node55692;
															assign node55692 = (inp[10]) ? node55694 : 4'b0111;
																assign node55694 = (inp[4]) ? 4'b0111 : 4'b0011;
															assign node55697 = (inp[10]) ? node55701 : node55698;
																assign node55698 = (inp[4]) ? 4'b0111 : 4'b0011;
																assign node55701 = (inp[4]) ? 4'b0011 : 4'b0111;
													assign node55704 = (inp[5]) ? node55716 : node55705;
														assign node55705 = (inp[10]) ? node55711 : node55706;
															assign node55706 = (inp[9]) ? node55708 : 4'b0011;
																assign node55708 = (inp[4]) ? 4'b0101 : 4'b0011;
															assign node55711 = (inp[9]) ? node55713 : 4'b0101;
																assign node55713 = (inp[4]) ? 4'b0001 : 4'b0101;
														assign node55716 = (inp[10]) ? node55722 : node55717;
															assign node55717 = (inp[4]) ? 4'b0101 : node55718;
																assign node55718 = (inp[9]) ? 4'b0001 : 4'b0101;
															assign node55722 = (inp[4]) ? node55726 : node55723;
																assign node55723 = (inp[9]) ? 4'b0101 : 4'b0001;
																assign node55726 = (inp[9]) ? 4'b0001 : 4'b0101;
											assign node55729 = (inp[10]) ? node55755 : node55730;
												assign node55730 = (inp[15]) ? node55744 : node55731;
													assign node55731 = (inp[5]) ? node55739 : node55732;
														assign node55732 = (inp[9]) ? node55736 : node55733;
															assign node55733 = (inp[4]) ? 4'b0111 : 4'b0001;
															assign node55736 = (inp[4]) ? 4'b0001 : 4'b0101;
														assign node55739 = (inp[3]) ? 4'b0011 : node55740;
															assign node55740 = (inp[4]) ? 4'b0011 : 4'b0001;
													assign node55744 = (inp[4]) ? node55752 : node55745;
														assign node55745 = (inp[9]) ? 4'b0101 : node55746;
															assign node55746 = (inp[3]) ? node55748 : 4'b0011;
																assign node55748 = (inp[5]) ? 4'b0001 : 4'b0011;
														assign node55752 = (inp[9]) ? 4'b0001 : 4'b0101;
												assign node55755 = (inp[3]) ? node55781 : node55756;
													assign node55756 = (inp[15]) ? node55770 : node55757;
														assign node55757 = (inp[5]) ? node55765 : node55758;
															assign node55758 = (inp[4]) ? node55762 : node55759;
																assign node55759 = (inp[9]) ? 4'b0101 : 4'b0001;
																assign node55762 = (inp[9]) ? 4'b0001 : 4'b0101;
															assign node55765 = (inp[9]) ? node55767 : 4'b0001;
																assign node55767 = (inp[4]) ? 4'b0011 : 4'b0111;
														assign node55770 = (inp[5]) ? node55778 : node55771;
															assign node55771 = (inp[4]) ? node55775 : node55772;
																assign node55772 = (inp[9]) ? 4'b0111 : 4'b0011;
																assign node55775 = (inp[9]) ? 4'b0011 : 4'b0111;
															assign node55778 = (inp[9]) ? 4'b0001 : 4'b0101;
													assign node55781 = (inp[15]) ? node55791 : node55782;
														assign node55782 = (inp[9]) ? node55788 : node55783;
															assign node55783 = (inp[4]) ? 4'b0111 : node55784;
																assign node55784 = (inp[5]) ? 4'b0011 : 4'b0001;
															assign node55788 = (inp[4]) ? 4'b0011 : 4'b0111;
														assign node55791 = (inp[5]) ? 4'b0001 : 4'b0011;
								assign node55794 = (inp[12]) ? node56052 : node55795;
									assign node55795 = (inp[4]) ? node55919 : node55796;
										assign node55796 = (inp[3]) ? node55848 : node55797;
											assign node55797 = (inp[0]) ? node55817 : node55798;
												assign node55798 = (inp[15]) ? node55808 : node55799;
													assign node55799 = (inp[9]) ? node55803 : node55800;
														assign node55800 = (inp[10]) ? 4'b0011 : 4'b0111;
														assign node55803 = (inp[10]) ? node55805 : 4'b0011;
															assign node55805 = (inp[14]) ? 4'b0101 : 4'b0111;
													assign node55808 = (inp[9]) ? node55812 : node55809;
														assign node55809 = (inp[10]) ? 4'b0001 : 4'b0101;
														assign node55812 = (inp[10]) ? node55814 : 4'b0001;
															assign node55814 = (inp[5]) ? 4'b0111 : 4'b0101;
												assign node55817 = (inp[15]) ? node55831 : node55818;
													assign node55818 = (inp[5]) ? node55824 : node55819;
														assign node55819 = (inp[10]) ? node55821 : 4'b0101;
															assign node55821 = (inp[9]) ? 4'b0101 : 4'b0001;
														assign node55824 = (inp[10]) ? node55828 : node55825;
															assign node55825 = (inp[9]) ? 4'b0001 : 4'b0101;
															assign node55828 = (inp[9]) ? 4'b0111 : 4'b0001;
													assign node55831 = (inp[5]) ? node55845 : node55832;
														assign node55832 = (inp[14]) ? node55838 : node55833;
															assign node55833 = (inp[10]) ? node55835 : 4'b0111;
																assign node55835 = (inp[9]) ? 4'b0111 : 4'b0011;
															assign node55838 = (inp[10]) ? node55842 : node55839;
																assign node55839 = (inp[9]) ? 4'b0011 : 4'b0111;
																assign node55842 = (inp[9]) ? 4'b0111 : 4'b0011;
														assign node55845 = (inp[10]) ? 4'b0101 : 4'b0111;
											assign node55848 = (inp[9]) ? node55882 : node55849;
												assign node55849 = (inp[10]) ? node55869 : node55850;
													assign node55850 = (inp[0]) ? node55856 : node55851;
														assign node55851 = (inp[15]) ? 4'b0101 : node55852;
															assign node55852 = (inp[5]) ? 4'b0101 : 4'b0111;
														assign node55856 = (inp[14]) ? node55864 : node55857;
															assign node55857 = (inp[15]) ? node55861 : node55858;
																assign node55858 = (inp[5]) ? 4'b0111 : 4'b0101;
																assign node55861 = (inp[5]) ? 4'b0101 : 4'b0111;
															assign node55864 = (inp[15]) ? node55866 : 4'b0101;
																assign node55866 = (inp[5]) ? 4'b0101 : 4'b0111;
													assign node55869 = (inp[15]) ? node55877 : node55870;
														assign node55870 = (inp[0]) ? node55874 : node55871;
															assign node55871 = (inp[5]) ? 4'b0001 : 4'b0011;
															assign node55874 = (inp[5]) ? 4'b0011 : 4'b0001;
														assign node55877 = (inp[0]) ? 4'b0001 : node55878;
															assign node55878 = (inp[5]) ? 4'b0011 : 4'b0001;
												assign node55882 = (inp[10]) ? node55902 : node55883;
													assign node55883 = (inp[5]) ? node55897 : node55884;
														assign node55884 = (inp[14]) ? node55890 : node55885;
															assign node55885 = (inp[0]) ? node55887 : 4'b0001;
																assign node55887 = (inp[15]) ? 4'b0011 : 4'b0001;
															assign node55890 = (inp[15]) ? node55894 : node55891;
																assign node55891 = (inp[0]) ? 4'b0001 : 4'b0011;
																assign node55894 = (inp[0]) ? 4'b0011 : 4'b0001;
														assign node55897 = (inp[0]) ? node55899 : 4'b0011;
															assign node55899 = (inp[15]) ? 4'b0001 : 4'b0011;
													assign node55902 = (inp[14]) ? node55910 : node55903;
														assign node55903 = (inp[0]) ? node55907 : node55904;
															assign node55904 = (inp[15]) ? 4'b0111 : 4'b0101;
															assign node55907 = (inp[15]) ? 4'b0101 : 4'b0111;
														assign node55910 = (inp[5]) ? node55912 : 4'b0101;
															assign node55912 = (inp[15]) ? node55916 : node55913;
																assign node55913 = (inp[0]) ? 4'b0111 : 4'b0101;
																assign node55916 = (inp[0]) ? 4'b0101 : 4'b0111;
										assign node55919 = (inp[9]) ? node55983 : node55920;
											assign node55920 = (inp[10]) ? node55958 : node55921;
												assign node55921 = (inp[3]) ? node55943 : node55922;
													assign node55922 = (inp[14]) ? node55928 : node55923;
														assign node55923 = (inp[0]) ? node55925 : 4'b0001;
															assign node55925 = (inp[15]) ? 4'b0011 : 4'b0001;
														assign node55928 = (inp[5]) ? node55936 : node55929;
															assign node55929 = (inp[15]) ? node55933 : node55930;
																assign node55930 = (inp[0]) ? 4'b0001 : 4'b0011;
																assign node55933 = (inp[0]) ? 4'b0011 : 4'b0001;
															assign node55936 = (inp[0]) ? node55940 : node55937;
																assign node55937 = (inp[15]) ? 4'b0001 : 4'b0011;
																assign node55940 = (inp[15]) ? 4'b0011 : 4'b0001;
													assign node55943 = (inp[5]) ? node55951 : node55944;
														assign node55944 = (inp[0]) ? node55948 : node55945;
															assign node55945 = (inp[15]) ? 4'b0001 : 4'b0011;
															assign node55948 = (inp[15]) ? 4'b0011 : 4'b0001;
														assign node55951 = (inp[15]) ? node55955 : node55952;
															assign node55952 = (inp[0]) ? 4'b0011 : 4'b0001;
															assign node55955 = (inp[0]) ? 4'b0001 : 4'b0011;
												assign node55958 = (inp[5]) ? node55976 : node55959;
													assign node55959 = (inp[14]) ? node55969 : node55960;
														assign node55960 = (inp[3]) ? 4'b0111 : node55961;
															assign node55961 = (inp[15]) ? node55965 : node55962;
																assign node55962 = (inp[0]) ? 4'b0101 : 4'b0111;
																assign node55965 = (inp[0]) ? 4'b0111 : 4'b0101;
														assign node55969 = (inp[3]) ? node55971 : 4'b0111;
															assign node55971 = (inp[15]) ? 4'b0111 : node55972;
																assign node55972 = (inp[0]) ? 4'b0111 : 4'b0101;
													assign node55976 = (inp[0]) ? node55980 : node55977;
														assign node55977 = (inp[15]) ? 4'b0111 : 4'b0101;
														assign node55980 = (inp[15]) ? 4'b0101 : 4'b0111;
											assign node55983 = (inp[10]) ? node56011 : node55984;
												assign node55984 = (inp[14]) ? node55996 : node55985;
													assign node55985 = (inp[3]) ? 4'b0101 : node55986;
														assign node55986 = (inp[0]) ? node55988 : 4'b0101;
															assign node55988 = (inp[15]) ? node55992 : node55989;
																assign node55989 = (inp[5]) ? 4'b0111 : 4'b0101;
																assign node55992 = (inp[5]) ? 4'b0101 : 4'b0111;
													assign node55996 = (inp[5]) ? node56004 : node55997;
														assign node55997 = (inp[3]) ? 4'b0101 : node55998;
															assign node55998 = (inp[15]) ? 4'b0111 : node55999;
																assign node55999 = (inp[0]) ? 4'b0101 : 4'b0111;
														assign node56004 = (inp[15]) ? node56008 : node56005;
															assign node56005 = (inp[0]) ? 4'b0111 : 4'b0101;
															assign node56008 = (inp[0]) ? 4'b0101 : 4'b0111;
												assign node56011 = (inp[5]) ? node56033 : node56012;
													assign node56012 = (inp[14]) ? node56024 : node56013;
														assign node56013 = (inp[15]) ? node56019 : node56014;
															assign node56014 = (inp[3]) ? node56016 : 4'b0001;
																assign node56016 = (inp[0]) ? 4'b0011 : 4'b0001;
															assign node56019 = (inp[3]) ? node56021 : 4'b0011;
																assign node56021 = (inp[0]) ? 4'b0001 : 4'b0011;
														assign node56024 = (inp[15]) ? 4'b0001 : node56025;
															assign node56025 = (inp[3]) ? node56029 : node56026;
																assign node56026 = (inp[0]) ? 4'b0001 : 4'b0011;
																assign node56029 = (inp[0]) ? 4'b0011 : 4'b0001;
													assign node56033 = (inp[14]) ? node56045 : node56034;
														assign node56034 = (inp[3]) ? node56040 : node56035;
															assign node56035 = (inp[0]) ? 4'b0001 : node56036;
																assign node56036 = (inp[15]) ? 4'b0011 : 4'b0001;
															assign node56040 = (inp[15]) ? 4'b0011 : node56041;
																assign node56041 = (inp[0]) ? 4'b0011 : 4'b0001;
														assign node56045 = (inp[0]) ? node56049 : node56046;
															assign node56046 = (inp[15]) ? 4'b0011 : 4'b0001;
															assign node56049 = (inp[15]) ? 4'b0001 : 4'b0011;
									assign node56052 = (inp[0]) ? node56104 : node56053;
										assign node56053 = (inp[15]) ? node56079 : node56054;
											assign node56054 = (inp[3]) ? node56070 : node56055;
												assign node56055 = (inp[5]) ? node56063 : node56056;
													assign node56056 = (inp[4]) ? node56060 : node56057;
														assign node56057 = (inp[9]) ? 4'b0111 : 4'b0011;
														assign node56060 = (inp[9]) ? 4'b0011 : 4'b0111;
													assign node56063 = (inp[4]) ? node56067 : node56064;
														assign node56064 = (inp[9]) ? 4'b0101 : 4'b0011;
														assign node56067 = (inp[9]) ? 4'b0001 : 4'b0101;
												assign node56070 = (inp[9]) ? node56076 : node56071;
													assign node56071 = (inp[4]) ? 4'b0101 : node56072;
														assign node56072 = (inp[5]) ? 4'b0001 : 4'b0011;
													assign node56076 = (inp[4]) ? 4'b0001 : 4'b0101;
											assign node56079 = (inp[3]) ? node56095 : node56080;
												assign node56080 = (inp[5]) ? node56088 : node56081;
													assign node56081 = (inp[4]) ? node56085 : node56082;
														assign node56082 = (inp[9]) ? 4'b0101 : 4'b0001;
														assign node56085 = (inp[9]) ? 4'b0001 : 4'b0101;
													assign node56088 = (inp[9]) ? node56092 : node56089;
														assign node56089 = (inp[4]) ? 4'b0111 : 4'b0001;
														assign node56092 = (inp[4]) ? 4'b0011 : 4'b0111;
												assign node56095 = (inp[4]) ? node56101 : node56096;
													assign node56096 = (inp[9]) ? 4'b0111 : node56097;
														assign node56097 = (inp[5]) ? 4'b0011 : 4'b0001;
													assign node56101 = (inp[9]) ? 4'b0011 : 4'b0111;
										assign node56104 = (inp[15]) ? node56144 : node56105;
											assign node56105 = (inp[5]) ? node56135 : node56106;
												assign node56106 = (inp[3]) ? node56128 : node56107;
													assign node56107 = (inp[14]) ? node56121 : node56108;
														assign node56108 = (inp[10]) ? node56116 : node56109;
															assign node56109 = (inp[4]) ? node56113 : node56110;
																assign node56110 = (inp[9]) ? 4'b0101 : 4'b0001;
																assign node56113 = (inp[9]) ? 4'b0001 : 4'b0101;
															assign node56116 = (inp[4]) ? 4'b0001 : node56117;
																assign node56117 = (inp[9]) ? 4'b0101 : 4'b0001;
														assign node56121 = (inp[10]) ? 4'b0101 : node56122;
															assign node56122 = (inp[9]) ? node56124 : 4'b0101;
																assign node56124 = (inp[4]) ? 4'b0001 : 4'b0101;
													assign node56128 = (inp[4]) ? node56132 : node56129;
														assign node56129 = (inp[9]) ? 4'b0111 : 4'b0001;
														assign node56132 = (inp[9]) ? 4'b0011 : 4'b0111;
												assign node56135 = (inp[9]) ? node56141 : node56136;
													assign node56136 = (inp[4]) ? 4'b0111 : node56137;
														assign node56137 = (inp[3]) ? 4'b0011 : 4'b0001;
													assign node56141 = (inp[4]) ? 4'b0011 : 4'b0111;
											assign node56144 = (inp[5]) ? node56168 : node56145;
												assign node56145 = (inp[3]) ? node56161 : node56146;
													assign node56146 = (inp[14]) ? node56154 : node56147;
														assign node56147 = (inp[9]) ? node56151 : node56148;
															assign node56148 = (inp[4]) ? 4'b0111 : 4'b0011;
															assign node56151 = (inp[4]) ? 4'b0011 : 4'b0111;
														assign node56154 = (inp[9]) ? node56158 : node56155;
															assign node56155 = (inp[4]) ? 4'b0111 : 4'b0011;
															assign node56158 = (inp[4]) ? 4'b0011 : 4'b0111;
													assign node56161 = (inp[4]) ? node56165 : node56162;
														assign node56162 = (inp[9]) ? 4'b0101 : 4'b0011;
														assign node56165 = (inp[9]) ? 4'b0001 : 4'b0101;
												assign node56168 = (inp[3]) ? node56176 : node56169;
													assign node56169 = (inp[4]) ? node56173 : node56170;
														assign node56170 = (inp[9]) ? 4'b0101 : 4'b0011;
														assign node56173 = (inp[9]) ? 4'b0001 : 4'b0101;
													assign node56176 = (inp[4]) ? node56180 : node56177;
														assign node56177 = (inp[9]) ? 4'b0101 : 4'b0001;
														assign node56180 = (inp[9]) ? 4'b0001 : 4'b0101;
						assign node56183 = (inp[7]) ? node57085 : node56184;
							assign node56184 = (inp[14]) ? node56726 : node56185;
								assign node56185 = (inp[2]) ? node56433 : node56186;
									assign node56186 = (inp[9]) ? node56306 : node56187;
										assign node56187 = (inp[4]) ? node56251 : node56188;
											assign node56188 = (inp[12]) ? node56228 : node56189;
												assign node56189 = (inp[10]) ? node56207 : node56190;
													assign node56190 = (inp[3]) ? node56198 : node56191;
														assign node56191 = (inp[0]) ? node56195 : node56192;
															assign node56192 = (inp[15]) ? 4'b1100 : 4'b1110;
															assign node56195 = (inp[15]) ? 4'b1110 : 4'b1100;
														assign node56198 = (inp[0]) ? node56200 : 4'b1100;
															assign node56200 = (inp[15]) ? node56204 : node56201;
																assign node56201 = (inp[5]) ? 4'b1110 : 4'b1100;
																assign node56204 = (inp[5]) ? 4'b1100 : 4'b1110;
													assign node56207 = (inp[3]) ? node56215 : node56208;
														assign node56208 = (inp[0]) ? node56212 : node56209;
															assign node56209 = (inp[15]) ? 4'b1000 : 4'b1010;
															assign node56212 = (inp[15]) ? 4'b1010 : 4'b1000;
														assign node56215 = (inp[5]) ? node56223 : node56216;
															assign node56216 = (inp[15]) ? node56220 : node56217;
																assign node56217 = (inp[0]) ? 4'b1000 : 4'b1010;
																assign node56220 = (inp[0]) ? 4'b1010 : 4'b1000;
															assign node56223 = (inp[0]) ? 4'b1010 : node56224;
																assign node56224 = (inp[15]) ? 4'b1010 : 4'b1000;
												assign node56228 = (inp[0]) ? node56240 : node56229;
													assign node56229 = (inp[15]) ? node56235 : node56230;
														assign node56230 = (inp[5]) ? node56232 : 4'b1010;
															assign node56232 = (inp[3]) ? 4'b1000 : 4'b1010;
														assign node56235 = (inp[3]) ? node56237 : 4'b1000;
															assign node56237 = (inp[5]) ? 4'b1010 : 4'b1000;
													assign node56240 = (inp[15]) ? node56246 : node56241;
														assign node56241 = (inp[3]) ? node56243 : 4'b1000;
															assign node56243 = (inp[5]) ? 4'b1010 : 4'b1000;
														assign node56246 = (inp[5]) ? node56248 : 4'b1010;
															assign node56248 = (inp[3]) ? 4'b1000 : 4'b1010;
											assign node56251 = (inp[10]) ? node56281 : node56252;
												assign node56252 = (inp[12]) ? node56266 : node56253;
													assign node56253 = (inp[5]) ? 4'b1010 : node56254;
														assign node56254 = (inp[3]) ? node56260 : node56255;
															assign node56255 = (inp[0]) ? 4'b1000 : node56256;
																assign node56256 = (inp[15]) ? 4'b1000 : 4'b1010;
															assign node56260 = (inp[0]) ? node56262 : 4'b1000;
																assign node56262 = (inp[15]) ? 4'b1010 : 4'b1000;
													assign node56266 = (inp[5]) ? node56274 : node56267;
														assign node56267 = (inp[3]) ? node56269 : 4'b1100;
															assign node56269 = (inp[15]) ? 4'b1100 : node56270;
																assign node56270 = (inp[0]) ? 4'b1110 : 4'b1100;
														assign node56274 = (inp[15]) ? node56278 : node56275;
															assign node56275 = (inp[0]) ? 4'b1110 : 4'b1100;
															assign node56278 = (inp[0]) ? 4'b1100 : 4'b1110;
												assign node56281 = (inp[3]) ? node56299 : node56282;
													assign node56282 = (inp[15]) ? node56292 : node56283;
														assign node56283 = (inp[12]) ? 4'b1110 : node56284;
															assign node56284 = (inp[5]) ? node56288 : node56285;
																assign node56285 = (inp[0]) ? 4'b1100 : 4'b1110;
																assign node56288 = (inp[0]) ? 4'b1110 : 4'b1100;
														assign node56292 = (inp[0]) ? node56296 : node56293;
															assign node56293 = (inp[5]) ? 4'b1110 : 4'b1100;
															assign node56296 = (inp[5]) ? 4'b1100 : 4'b1110;
													assign node56299 = (inp[15]) ? node56303 : node56300;
														assign node56300 = (inp[0]) ? 4'b1110 : 4'b1100;
														assign node56303 = (inp[0]) ? 4'b1100 : 4'b1110;
										assign node56306 = (inp[4]) ? node56368 : node56307;
											assign node56307 = (inp[12]) ? node56345 : node56308;
												assign node56308 = (inp[10]) ? node56326 : node56309;
													assign node56309 = (inp[15]) ? node56319 : node56310;
														assign node56310 = (inp[0]) ? node56314 : node56311;
															assign node56311 = (inp[3]) ? 4'b1000 : 4'b1010;
															assign node56314 = (inp[3]) ? node56316 : 4'b1000;
																assign node56316 = (inp[5]) ? 4'b1010 : 4'b1000;
														assign node56319 = (inp[0]) ? 4'b1010 : node56320;
															assign node56320 = (inp[5]) ? node56322 : 4'b1000;
																assign node56322 = (inp[3]) ? 4'b1010 : 4'b1000;
													assign node56326 = (inp[15]) ? node56336 : node56327;
														assign node56327 = (inp[3]) ? node56333 : node56328;
															assign node56328 = (inp[0]) ? node56330 : 4'b1110;
																assign node56330 = (inp[5]) ? 4'b1110 : 4'b1100;
															assign node56333 = (inp[0]) ? 4'b1110 : 4'b1100;
														assign node56336 = (inp[3]) ? 4'b1110 : node56337;
															assign node56337 = (inp[5]) ? node56341 : node56338;
																assign node56338 = (inp[0]) ? 4'b1110 : 4'b1100;
																assign node56341 = (inp[0]) ? 4'b1100 : 4'b1110;
												assign node56345 = (inp[15]) ? node56357 : node56346;
													assign node56346 = (inp[0]) ? node56352 : node56347;
														assign node56347 = (inp[3]) ? 4'b1100 : node56348;
															assign node56348 = (inp[5]) ? 4'b1100 : 4'b1110;
														assign node56352 = (inp[3]) ? 4'b1110 : node56353;
															assign node56353 = (inp[5]) ? 4'b1110 : 4'b1100;
													assign node56357 = (inp[10]) ? 4'b1110 : node56358;
														assign node56358 = (inp[5]) ? 4'b1110 : node56359;
															assign node56359 = (inp[3]) ? node56363 : node56360;
																assign node56360 = (inp[0]) ? 4'b1110 : 4'b1100;
																assign node56363 = (inp[0]) ? 4'b1100 : 4'b1110;
											assign node56368 = (inp[12]) ? node56410 : node56369;
												assign node56369 = (inp[10]) ? node56393 : node56370;
													assign node56370 = (inp[5]) ? node56380 : node56371;
														assign node56371 = (inp[0]) ? 4'b1110 : node56372;
															assign node56372 = (inp[15]) ? node56376 : node56373;
																assign node56373 = (inp[3]) ? 4'b1100 : 4'b1110;
																assign node56376 = (inp[3]) ? 4'b1110 : 4'b1100;
														assign node56380 = (inp[3]) ? node56386 : node56381;
															assign node56381 = (inp[15]) ? node56383 : 4'b1100;
																assign node56383 = (inp[0]) ? 4'b1100 : 4'b1110;
															assign node56386 = (inp[15]) ? node56390 : node56387;
																assign node56387 = (inp[0]) ? 4'b1110 : 4'b1100;
																assign node56390 = (inp[0]) ? 4'b1100 : 4'b1110;
													assign node56393 = (inp[0]) ? node56403 : node56394;
														assign node56394 = (inp[15]) ? node56400 : node56395;
															assign node56395 = (inp[5]) ? 4'b1000 : node56396;
																assign node56396 = (inp[3]) ? 4'b1000 : 4'b1010;
															assign node56400 = (inp[5]) ? 4'b1010 : 4'b1000;
														assign node56403 = (inp[15]) ? node56405 : 4'b1010;
															assign node56405 = (inp[3]) ? 4'b1000 : node56406;
																assign node56406 = (inp[5]) ? 4'b1000 : 4'b1010;
												assign node56410 = (inp[0]) ? node56422 : node56411;
													assign node56411 = (inp[15]) ? node56417 : node56412;
														assign node56412 = (inp[5]) ? 4'b1000 : node56413;
															assign node56413 = (inp[3]) ? 4'b1000 : 4'b1010;
														assign node56417 = (inp[3]) ? 4'b1010 : node56418;
															assign node56418 = (inp[5]) ? 4'b1010 : 4'b1000;
													assign node56422 = (inp[15]) ? node56428 : node56423;
														assign node56423 = (inp[3]) ? 4'b1010 : node56424;
															assign node56424 = (inp[5]) ? 4'b1010 : 4'b1000;
														assign node56428 = (inp[5]) ? 4'b1000 : node56429;
															assign node56429 = (inp[3]) ? 4'b1000 : 4'b1010;
									assign node56433 = (inp[5]) ? node56569 : node56434;
										assign node56434 = (inp[4]) ? node56502 : node56435;
											assign node56435 = (inp[9]) ? node56473 : node56436;
												assign node56436 = (inp[10]) ? node56458 : node56437;
													assign node56437 = (inp[12]) ? node56445 : node56438;
														assign node56438 = (inp[15]) ? node56442 : node56439;
															assign node56439 = (inp[0]) ? 4'b0101 : 4'b0111;
															assign node56442 = (inp[0]) ? 4'b0111 : 4'b0101;
														assign node56445 = (inp[3]) ? node56451 : node56446;
															assign node56446 = (inp[15]) ? node56448 : 4'b0011;
																assign node56448 = (inp[0]) ? 4'b0011 : 4'b0001;
															assign node56451 = (inp[0]) ? node56455 : node56452;
																assign node56452 = (inp[15]) ? 4'b0001 : 4'b0011;
																assign node56455 = (inp[15]) ? 4'b0011 : 4'b0001;
													assign node56458 = (inp[12]) ? node56466 : node56459;
														assign node56459 = (inp[0]) ? node56463 : node56460;
															assign node56460 = (inp[15]) ? 4'b0001 : 4'b0011;
															assign node56463 = (inp[15]) ? 4'b0011 : 4'b0001;
														assign node56466 = (inp[3]) ? 4'b0011 : node56467;
															assign node56467 = (inp[15]) ? 4'b0011 : node56468;
																assign node56468 = (inp[0]) ? 4'b0001 : 4'b0011;
												assign node56473 = (inp[12]) ? node56489 : node56474;
													assign node56474 = (inp[10]) ? node56482 : node56475;
														assign node56475 = (inp[0]) ? node56479 : node56476;
															assign node56476 = (inp[15]) ? 4'b0001 : 4'b0011;
															assign node56479 = (inp[15]) ? 4'b0011 : 4'b0001;
														assign node56482 = (inp[15]) ? node56484 : 4'b0111;
															assign node56484 = (inp[3]) ? node56486 : 4'b0101;
																assign node56486 = (inp[0]) ? 4'b0101 : 4'b0111;
													assign node56489 = (inp[15]) ? node56495 : node56490;
														assign node56490 = (inp[0]) ? node56492 : 4'b0101;
															assign node56492 = (inp[3]) ? 4'b0111 : 4'b0101;
														assign node56495 = (inp[0]) ? node56499 : node56496;
															assign node56496 = (inp[3]) ? 4'b0111 : 4'b0101;
															assign node56499 = (inp[3]) ? 4'b0101 : 4'b0111;
											assign node56502 = (inp[9]) ? node56540 : node56503;
												assign node56503 = (inp[12]) ? node56521 : node56504;
													assign node56504 = (inp[10]) ? node56512 : node56505;
														assign node56505 = (inp[0]) ? node56509 : node56506;
															assign node56506 = (inp[15]) ? 4'b0001 : 4'b0011;
															assign node56509 = (inp[15]) ? 4'b0011 : 4'b0001;
														assign node56512 = (inp[0]) ? 4'b0111 : node56513;
															assign node56513 = (inp[15]) ? node56517 : node56514;
																assign node56514 = (inp[3]) ? 4'b0101 : 4'b0111;
																assign node56517 = (inp[3]) ? 4'b0111 : 4'b0101;
													assign node56521 = (inp[0]) ? node56535 : node56522;
														assign node56522 = (inp[10]) ? node56530 : node56523;
															assign node56523 = (inp[15]) ? node56527 : node56524;
																assign node56524 = (inp[3]) ? 4'b0101 : 4'b0111;
																assign node56527 = (inp[3]) ? 4'b0111 : 4'b0101;
															assign node56530 = (inp[15]) ? node56532 : 4'b0111;
																assign node56532 = (inp[3]) ? 4'b0111 : 4'b0101;
														assign node56535 = (inp[15]) ? node56537 : 4'b0101;
															assign node56537 = (inp[3]) ? 4'b0101 : 4'b0111;
												assign node56540 = (inp[12]) ? node56558 : node56541;
													assign node56541 = (inp[10]) ? node56551 : node56542;
														assign node56542 = (inp[3]) ? node56544 : 4'b0111;
															assign node56544 = (inp[15]) ? node56548 : node56545;
																assign node56545 = (inp[0]) ? 4'b0111 : 4'b0101;
																assign node56548 = (inp[0]) ? 4'b0101 : 4'b0111;
														assign node56551 = (inp[15]) ? 4'b0001 : node56552;
															assign node56552 = (inp[0]) ? node56554 : 4'b0011;
																assign node56554 = (inp[3]) ? 4'b0011 : 4'b0001;
													assign node56558 = (inp[3]) ? 4'b0011 : node56559;
														assign node56559 = (inp[10]) ? 4'b0011 : node56560;
															assign node56560 = (inp[0]) ? node56564 : node56561;
																assign node56561 = (inp[15]) ? 4'b0001 : 4'b0011;
																assign node56564 = (inp[15]) ? 4'b0011 : 4'b0001;
										assign node56569 = (inp[3]) ? node56651 : node56570;
											assign node56570 = (inp[12]) ? node56622 : node56571;
												assign node56571 = (inp[4]) ? node56595 : node56572;
													assign node56572 = (inp[9]) ? node56582 : node56573;
														assign node56573 = (inp[10]) ? node56579 : node56574;
															assign node56574 = (inp[15]) ? 4'b0111 : node56575;
																assign node56575 = (inp[0]) ? 4'b0101 : 4'b0111;
															assign node56579 = (inp[15]) ? 4'b0001 : 4'b0011;
														assign node56582 = (inp[10]) ? node56588 : node56583;
															assign node56583 = (inp[0]) ? node56585 : 4'b0001;
																assign node56585 = (inp[15]) ? 4'b0011 : 4'b0001;
															assign node56588 = (inp[15]) ? node56592 : node56589;
																assign node56589 = (inp[0]) ? 4'b0111 : 4'b0101;
																assign node56592 = (inp[0]) ? 4'b0101 : 4'b0111;
													assign node56595 = (inp[15]) ? node56607 : node56596;
														assign node56596 = (inp[0]) ? node56604 : node56597;
															assign node56597 = (inp[9]) ? node56601 : node56598;
																assign node56598 = (inp[10]) ? 4'b0101 : 4'b0011;
																assign node56601 = (inp[10]) ? 4'b0001 : 4'b0101;
															assign node56604 = (inp[9]) ? 4'b0011 : 4'b0001;
														assign node56607 = (inp[0]) ? node56615 : node56608;
															assign node56608 = (inp[10]) ? node56612 : node56609;
																assign node56609 = (inp[9]) ? 4'b0111 : 4'b0001;
																assign node56612 = (inp[9]) ? 4'b0011 : 4'b0111;
															assign node56615 = (inp[9]) ? node56619 : node56616;
																assign node56616 = (inp[10]) ? 4'b0101 : 4'b0011;
																assign node56619 = (inp[10]) ? 4'b0001 : 4'b0101;
												assign node56622 = (inp[0]) ? node56636 : node56623;
													assign node56623 = (inp[15]) ? node56629 : node56624;
														assign node56624 = (inp[9]) ? node56626 : 4'b0011;
															assign node56626 = (inp[4]) ? 4'b0001 : 4'b0101;
														assign node56629 = (inp[9]) ? node56633 : node56630;
															assign node56630 = (inp[4]) ? 4'b0111 : 4'b0001;
															assign node56633 = (inp[4]) ? 4'b0011 : 4'b0111;
													assign node56636 = (inp[15]) ? node56644 : node56637;
														assign node56637 = (inp[9]) ? node56641 : node56638;
															assign node56638 = (inp[4]) ? 4'b0111 : 4'b0001;
															assign node56641 = (inp[4]) ? 4'b0011 : 4'b0111;
														assign node56644 = (inp[4]) ? node56648 : node56645;
															assign node56645 = (inp[9]) ? 4'b0101 : 4'b0011;
															assign node56648 = (inp[9]) ? 4'b0001 : 4'b0101;
											assign node56651 = (inp[4]) ? node56685 : node56652;
												assign node56652 = (inp[9]) ? node56670 : node56653;
													assign node56653 = (inp[12]) ? node56663 : node56654;
														assign node56654 = (inp[10]) ? node56658 : node56655;
															assign node56655 = (inp[15]) ? 4'b0111 : 4'b0101;
															assign node56658 = (inp[0]) ? 4'b0001 : node56659;
																assign node56659 = (inp[15]) ? 4'b0011 : 4'b0001;
														assign node56663 = (inp[15]) ? node56667 : node56664;
															assign node56664 = (inp[0]) ? 4'b0011 : 4'b0001;
															assign node56667 = (inp[0]) ? 4'b0001 : 4'b0011;
													assign node56670 = (inp[12]) ? node56680 : node56671;
														assign node56671 = (inp[10]) ? node56677 : node56672;
															assign node56672 = (inp[0]) ? 4'b0001 : node56673;
																assign node56673 = (inp[15]) ? 4'b0011 : 4'b0001;
															assign node56677 = (inp[15]) ? 4'b0101 : 4'b0111;
														assign node56680 = (inp[0]) ? node56682 : 4'b0101;
															assign node56682 = (inp[15]) ? 4'b0101 : 4'b0111;
												assign node56685 = (inp[9]) ? node56705 : node56686;
													assign node56686 = (inp[10]) ? node56700 : node56687;
														assign node56687 = (inp[12]) ? node56695 : node56688;
															assign node56688 = (inp[15]) ? node56692 : node56689;
																assign node56689 = (inp[0]) ? 4'b0011 : 4'b0001;
																assign node56692 = (inp[0]) ? 4'b0001 : 4'b0011;
															assign node56695 = (inp[15]) ? node56697 : 4'b0101;
																assign node56697 = (inp[0]) ? 4'b0101 : 4'b0111;
														assign node56700 = (inp[0]) ? 4'b0101 : node56701;
															assign node56701 = (inp[15]) ? 4'b0111 : 4'b0101;
													assign node56705 = (inp[12]) ? node56713 : node56706;
														assign node56706 = (inp[10]) ? 4'b0001 : node56707;
															assign node56707 = (inp[0]) ? node56709 : 4'b0101;
																assign node56709 = (inp[15]) ? 4'b0101 : 4'b0111;
														assign node56713 = (inp[10]) ? node56719 : node56714;
															assign node56714 = (inp[15]) ? 4'b0001 : node56715;
																assign node56715 = (inp[0]) ? 4'b0011 : 4'b0001;
															assign node56719 = (inp[15]) ? node56723 : node56720;
																assign node56720 = (inp[0]) ? 4'b0011 : 4'b0001;
																assign node56723 = (inp[0]) ? 4'b0001 : 4'b0011;
								assign node56726 = (inp[0]) ? node56928 : node56727;
									assign node56727 = (inp[15]) ? node56837 : node56728;
										assign node56728 = (inp[3]) ? node56790 : node56729;
											assign node56729 = (inp[5]) ? node56767 : node56730;
												assign node56730 = (inp[12]) ? node56746 : node56731;
													assign node56731 = (inp[4]) ? node56739 : node56732;
														assign node56732 = (inp[10]) ? node56736 : node56733;
															assign node56733 = (inp[9]) ? 4'b0011 : 4'b0111;
															assign node56736 = (inp[9]) ? 4'b0111 : 4'b0011;
														assign node56739 = (inp[9]) ? node56743 : node56740;
															assign node56740 = (inp[10]) ? 4'b0111 : 4'b0011;
															assign node56743 = (inp[10]) ? 4'b0011 : 4'b0111;
													assign node56746 = (inp[10]) ? node56754 : node56747;
														assign node56747 = (inp[9]) ? node56751 : node56748;
															assign node56748 = (inp[4]) ? 4'b0111 : 4'b0011;
															assign node56751 = (inp[4]) ? 4'b0011 : 4'b0111;
														assign node56754 = (inp[2]) ? node56760 : node56755;
															assign node56755 = (inp[4]) ? 4'b0111 : node56756;
																assign node56756 = (inp[9]) ? 4'b0111 : 4'b0011;
															assign node56760 = (inp[4]) ? node56764 : node56761;
																assign node56761 = (inp[9]) ? 4'b0111 : 4'b0011;
																assign node56764 = (inp[9]) ? 4'b0011 : 4'b0111;
												assign node56767 = (inp[9]) ? node56779 : node56768;
													assign node56768 = (inp[4]) ? node56774 : node56769;
														assign node56769 = (inp[12]) ? 4'b0011 : node56770;
															assign node56770 = (inp[10]) ? 4'b0011 : 4'b0111;
														assign node56774 = (inp[2]) ? node56776 : 4'b0101;
															assign node56776 = (inp[12]) ? 4'b0101 : 4'b0011;
													assign node56779 = (inp[4]) ? node56785 : node56780;
														assign node56780 = (inp[10]) ? 4'b0101 : node56781;
															assign node56781 = (inp[12]) ? 4'b0101 : 4'b0011;
														assign node56785 = (inp[2]) ? 4'b0001 : node56786;
															assign node56786 = (inp[10]) ? 4'b0001 : 4'b0101;
											assign node56790 = (inp[5]) ? node56814 : node56791;
												assign node56791 = (inp[4]) ? node56803 : node56792;
													assign node56792 = (inp[9]) ? node56798 : node56793;
														assign node56793 = (inp[10]) ? 4'b0011 : node56794;
															assign node56794 = (inp[12]) ? 4'b0011 : 4'b0111;
														assign node56798 = (inp[12]) ? 4'b0101 : node56799;
															assign node56799 = (inp[10]) ? 4'b0101 : 4'b0011;
													assign node56803 = (inp[9]) ? node56809 : node56804;
														assign node56804 = (inp[2]) ? node56806 : 4'b0101;
															assign node56806 = (inp[10]) ? 4'b0101 : 4'b0011;
														assign node56809 = (inp[10]) ? 4'b0001 : node56810;
															assign node56810 = (inp[12]) ? 4'b0001 : 4'b0101;
												assign node56814 = (inp[4]) ? node56826 : node56815;
													assign node56815 = (inp[9]) ? node56821 : node56816;
														assign node56816 = (inp[12]) ? 4'b0001 : node56817;
															assign node56817 = (inp[10]) ? 4'b0001 : 4'b0101;
														assign node56821 = (inp[12]) ? 4'b0101 : node56822;
															assign node56822 = (inp[10]) ? 4'b0101 : 4'b0001;
													assign node56826 = (inp[9]) ? node56832 : node56827;
														assign node56827 = (inp[12]) ? 4'b0101 : node56828;
															assign node56828 = (inp[10]) ? 4'b0101 : 4'b0001;
														assign node56832 = (inp[12]) ? 4'b0001 : node56833;
															assign node56833 = (inp[10]) ? 4'b0001 : 4'b0101;
										assign node56837 = (inp[3]) ? node56877 : node56838;
											assign node56838 = (inp[5]) ? node56858 : node56839;
												assign node56839 = (inp[4]) ? node56847 : node56840;
													assign node56840 = (inp[9]) ? node56842 : 4'b0001;
														assign node56842 = (inp[10]) ? 4'b0101 : node56843;
															assign node56843 = (inp[12]) ? 4'b0101 : 4'b0001;
													assign node56847 = (inp[9]) ? node56855 : node56848;
														assign node56848 = (inp[2]) ? node56850 : 4'b0101;
															assign node56850 = (inp[10]) ? 4'b0101 : node56851;
																assign node56851 = (inp[12]) ? 4'b0101 : 4'b0001;
														assign node56855 = (inp[10]) ? 4'b0001 : 4'b0101;
												assign node56858 = (inp[9]) ? node56868 : node56859;
													assign node56859 = (inp[4]) ? node56865 : node56860;
														assign node56860 = (inp[12]) ? 4'b0001 : node56861;
															assign node56861 = (inp[10]) ? 4'b0001 : 4'b0101;
														assign node56865 = (inp[12]) ? 4'b0111 : 4'b0001;
													assign node56868 = (inp[4]) ? node56874 : node56869;
														assign node56869 = (inp[10]) ? 4'b0111 : node56870;
															assign node56870 = (inp[12]) ? 4'b0111 : 4'b0001;
														assign node56874 = (inp[10]) ? 4'b0011 : 4'b0111;
											assign node56877 = (inp[5]) ? node56897 : node56878;
												assign node56878 = (inp[4]) ? node56890 : node56879;
													assign node56879 = (inp[9]) ? node56885 : node56880;
														assign node56880 = (inp[12]) ? 4'b0001 : node56881;
															assign node56881 = (inp[10]) ? 4'b0001 : 4'b0101;
														assign node56885 = (inp[12]) ? 4'b0111 : node56886;
															assign node56886 = (inp[10]) ? 4'b0111 : 4'b0001;
													assign node56890 = (inp[9]) ? node56892 : 4'b0111;
														assign node56892 = (inp[10]) ? 4'b0011 : node56893;
															assign node56893 = (inp[12]) ? 4'b0011 : 4'b0111;
												assign node56897 = (inp[10]) ? node56921 : node56898;
													assign node56898 = (inp[9]) ? node56906 : node56899;
														assign node56899 = (inp[12]) ? node56903 : node56900;
															assign node56900 = (inp[4]) ? 4'b0011 : 4'b0111;
															assign node56903 = (inp[4]) ? 4'b0111 : 4'b0011;
														assign node56906 = (inp[2]) ? node56914 : node56907;
															assign node56907 = (inp[4]) ? node56911 : node56908;
																assign node56908 = (inp[12]) ? 4'b0111 : 4'b0011;
																assign node56911 = (inp[12]) ? 4'b0011 : 4'b0111;
															assign node56914 = (inp[4]) ? node56918 : node56915;
																assign node56915 = (inp[12]) ? 4'b0111 : 4'b0011;
																assign node56918 = (inp[12]) ? 4'b0011 : 4'b0111;
													assign node56921 = (inp[9]) ? node56925 : node56922;
														assign node56922 = (inp[4]) ? 4'b0111 : 4'b0011;
														assign node56925 = (inp[4]) ? 4'b0011 : 4'b0111;
									assign node56928 = (inp[15]) ? node57004 : node56929;
										assign node56929 = (inp[5]) ? node56973 : node56930;
											assign node56930 = (inp[3]) ? node56950 : node56931;
												assign node56931 = (inp[9]) ? node56943 : node56932;
													assign node56932 = (inp[4]) ? node56938 : node56933;
														assign node56933 = (inp[12]) ? 4'b0001 : node56934;
															assign node56934 = (inp[10]) ? 4'b0001 : 4'b0101;
														assign node56938 = (inp[10]) ? 4'b0101 : node56939;
															assign node56939 = (inp[12]) ? 4'b0101 : 4'b0001;
													assign node56943 = (inp[4]) ? 4'b0001 : node56944;
														assign node56944 = (inp[10]) ? 4'b0101 : node56945;
															assign node56945 = (inp[12]) ? 4'b0101 : 4'b0001;
												assign node56950 = (inp[4]) ? node56962 : node56951;
													assign node56951 = (inp[9]) ? node56957 : node56952;
														assign node56952 = (inp[10]) ? 4'b0001 : node56953;
															assign node56953 = (inp[12]) ? 4'b0001 : 4'b0101;
														assign node56957 = (inp[12]) ? 4'b0111 : node56958;
															assign node56958 = (inp[10]) ? 4'b0111 : 4'b0001;
													assign node56962 = (inp[9]) ? node56968 : node56963;
														assign node56963 = (inp[10]) ? 4'b0111 : node56964;
															assign node56964 = (inp[12]) ? 4'b0111 : 4'b0001;
														assign node56968 = (inp[12]) ? 4'b0011 : node56969;
															assign node56969 = (inp[10]) ? 4'b0011 : 4'b0111;
											assign node56973 = (inp[3]) ? node56989 : node56974;
												assign node56974 = (inp[9]) ? node56984 : node56975;
													assign node56975 = (inp[4]) ? node56979 : node56976;
														assign node56976 = (inp[12]) ? 4'b0001 : 4'b0101;
														assign node56979 = (inp[12]) ? 4'b0111 : node56980;
															assign node56980 = (inp[10]) ? 4'b0111 : 4'b0001;
													assign node56984 = (inp[4]) ? node56986 : 4'b0111;
														assign node56986 = (inp[10]) ? 4'b0011 : 4'b0111;
												assign node56989 = (inp[9]) ? node56995 : node56990;
													assign node56990 = (inp[4]) ? node56992 : 4'b0011;
														assign node56992 = (inp[12]) ? 4'b0111 : 4'b0011;
													assign node56995 = (inp[4]) ? node57001 : node56996;
														assign node56996 = (inp[12]) ? 4'b0111 : node56997;
															assign node56997 = (inp[10]) ? 4'b0111 : 4'b0011;
														assign node57001 = (inp[10]) ? 4'b0011 : 4'b0111;
										assign node57004 = (inp[5]) ? node57048 : node57005;
											assign node57005 = (inp[3]) ? node57025 : node57006;
												assign node57006 = (inp[9]) ? node57018 : node57007;
													assign node57007 = (inp[4]) ? node57013 : node57008;
														assign node57008 = (inp[10]) ? 4'b0011 : node57009;
															assign node57009 = (inp[12]) ? 4'b0011 : 4'b0111;
														assign node57013 = (inp[12]) ? 4'b0111 : node57014;
															assign node57014 = (inp[10]) ? 4'b0111 : 4'b0011;
													assign node57018 = (inp[4]) ? node57020 : 4'b0111;
														assign node57020 = (inp[12]) ? 4'b0011 : node57021;
															assign node57021 = (inp[10]) ? 4'b0011 : 4'b0111;
												assign node57025 = (inp[9]) ? node57037 : node57026;
													assign node57026 = (inp[4]) ? node57032 : node57027;
														assign node57027 = (inp[10]) ? 4'b0011 : node57028;
															assign node57028 = (inp[12]) ? 4'b0011 : 4'b0111;
														assign node57032 = (inp[10]) ? 4'b0101 : node57033;
															assign node57033 = (inp[12]) ? 4'b0101 : 4'b0011;
													assign node57037 = (inp[4]) ? node57043 : node57038;
														assign node57038 = (inp[10]) ? 4'b0101 : node57039;
															assign node57039 = (inp[12]) ? 4'b0101 : 4'b0011;
														assign node57043 = (inp[10]) ? 4'b0001 : node57044;
															assign node57044 = (inp[12]) ? 4'b0001 : 4'b0101;
											assign node57048 = (inp[3]) ? node57068 : node57049;
												assign node57049 = (inp[4]) ? node57057 : node57050;
													assign node57050 = (inp[9]) ? node57052 : 4'b0011;
														assign node57052 = (inp[10]) ? 4'b0101 : node57053;
															assign node57053 = (inp[12]) ? 4'b0101 : 4'b0011;
													assign node57057 = (inp[9]) ? node57063 : node57058;
														assign node57058 = (inp[10]) ? 4'b0101 : node57059;
															assign node57059 = (inp[12]) ? 4'b0101 : 4'b0011;
														assign node57063 = (inp[10]) ? 4'b0001 : node57064;
															assign node57064 = (inp[12]) ? 4'b0001 : 4'b0101;
												assign node57068 = (inp[9]) ? node57078 : node57069;
													assign node57069 = (inp[4]) ? node57073 : node57070;
														assign node57070 = (inp[12]) ? 4'b0001 : 4'b0101;
														assign node57073 = (inp[12]) ? 4'b0101 : node57074;
															assign node57074 = (inp[10]) ? 4'b0101 : 4'b0001;
													assign node57078 = (inp[4]) ? 4'b0001 : node57079;
														assign node57079 = (inp[10]) ? 4'b0101 : node57080;
															assign node57080 = (inp[12]) ? 4'b0101 : 4'b0001;
							assign node57085 = (inp[2]) ? node57667 : node57086;
								assign node57086 = (inp[14]) ? node57382 : node57087;
									assign node57087 = (inp[10]) ? node57275 : node57088;
										assign node57088 = (inp[5]) ? node57178 : node57089;
											assign node57089 = (inp[9]) ? node57131 : node57090;
												assign node57090 = (inp[3]) ? node57108 : node57091;
													assign node57091 = (inp[4]) ? node57105 : node57092;
														assign node57092 = (inp[12]) ? node57100 : node57093;
															assign node57093 = (inp[15]) ? node57097 : node57094;
																assign node57094 = (inp[0]) ? 4'b0101 : 4'b0111;
																assign node57097 = (inp[0]) ? 4'b0111 : 4'b0101;
															assign node57100 = (inp[0]) ? 4'b0011 : node57101;
																assign node57101 = (inp[15]) ? 4'b0001 : 4'b0011;
														assign node57105 = (inp[12]) ? 4'b0111 : 4'b0011;
													assign node57108 = (inp[12]) ? node57120 : node57109;
														assign node57109 = (inp[4]) ? node57113 : node57110;
															assign node57110 = (inp[0]) ? 4'b0111 : 4'b0101;
															assign node57113 = (inp[0]) ? node57117 : node57114;
																assign node57114 = (inp[15]) ? 4'b0001 : 4'b0011;
																assign node57117 = (inp[15]) ? 4'b0011 : 4'b0001;
														assign node57120 = (inp[4]) ? node57124 : node57121;
															assign node57121 = (inp[15]) ? 4'b0011 : 4'b0001;
															assign node57124 = (inp[0]) ? node57128 : node57125;
																assign node57125 = (inp[15]) ? 4'b0111 : 4'b0101;
																assign node57128 = (inp[15]) ? 4'b0101 : 4'b0111;
												assign node57131 = (inp[0]) ? node57161 : node57132;
													assign node57132 = (inp[15]) ? node57148 : node57133;
														assign node57133 = (inp[3]) ? node57141 : node57134;
															assign node57134 = (inp[12]) ? node57138 : node57135;
																assign node57135 = (inp[4]) ? 4'b0111 : 4'b0011;
																assign node57138 = (inp[4]) ? 4'b0011 : 4'b0111;
															assign node57141 = (inp[4]) ? node57145 : node57142;
																assign node57142 = (inp[12]) ? 4'b0101 : 4'b0011;
																assign node57145 = (inp[12]) ? 4'b0001 : 4'b0101;
														assign node57148 = (inp[3]) ? node57154 : node57149;
															assign node57149 = (inp[4]) ? node57151 : 4'b0001;
																assign node57151 = (inp[12]) ? 4'b0001 : 4'b0101;
															assign node57154 = (inp[12]) ? node57158 : node57155;
																assign node57155 = (inp[4]) ? 4'b0111 : 4'b0001;
																assign node57158 = (inp[4]) ? 4'b0011 : 4'b0111;
													assign node57161 = (inp[15]) ? node57169 : node57162;
														assign node57162 = (inp[4]) ? node57164 : 4'b0001;
															assign node57164 = (inp[3]) ? node57166 : 4'b0001;
																assign node57166 = (inp[12]) ? 4'b0011 : 4'b0111;
														assign node57169 = (inp[3]) ? node57175 : node57170;
															assign node57170 = (inp[12]) ? node57172 : 4'b0011;
																assign node57172 = (inp[4]) ? 4'b0011 : 4'b0111;
															assign node57175 = (inp[4]) ? 4'b0001 : 4'b0011;
											assign node57178 = (inp[3]) ? node57232 : node57179;
												assign node57179 = (inp[4]) ? node57203 : node57180;
													assign node57180 = (inp[12]) ? node57194 : node57181;
														assign node57181 = (inp[9]) ? node57189 : node57182;
															assign node57182 = (inp[0]) ? node57186 : node57183;
																assign node57183 = (inp[15]) ? 4'b0101 : 4'b0111;
																assign node57186 = (inp[15]) ? 4'b0111 : 4'b0101;
															assign node57189 = (inp[0]) ? node57191 : 4'b0001;
																assign node57191 = (inp[15]) ? 4'b0011 : 4'b0001;
														assign node57194 = (inp[9]) ? node57196 : 4'b0001;
															assign node57196 = (inp[15]) ? node57200 : node57197;
																assign node57197 = (inp[0]) ? 4'b0111 : 4'b0101;
																assign node57200 = (inp[0]) ? 4'b0101 : 4'b0111;
													assign node57203 = (inp[12]) ? node57217 : node57204;
														assign node57204 = (inp[9]) ? node57212 : node57205;
															assign node57205 = (inp[15]) ? node57209 : node57206;
																assign node57206 = (inp[0]) ? 4'b0001 : 4'b0011;
																assign node57209 = (inp[0]) ? 4'b0011 : 4'b0001;
															assign node57212 = (inp[0]) ? 4'b0101 : node57213;
																assign node57213 = (inp[15]) ? 4'b0111 : 4'b0101;
														assign node57217 = (inp[9]) ? node57225 : node57218;
															assign node57218 = (inp[0]) ? node57222 : node57219;
																assign node57219 = (inp[15]) ? 4'b0111 : 4'b0101;
																assign node57222 = (inp[15]) ? 4'b0101 : 4'b0111;
															assign node57225 = (inp[15]) ? node57229 : node57226;
																assign node57226 = (inp[0]) ? 4'b0011 : 4'b0001;
																assign node57229 = (inp[0]) ? 4'b0001 : 4'b0011;
												assign node57232 = (inp[12]) ? node57250 : node57233;
													assign node57233 = (inp[4]) ? node57241 : node57234;
														assign node57234 = (inp[9]) ? node57236 : 4'b0111;
															assign node57236 = (inp[15]) ? 4'b0011 : node57237;
																assign node57237 = (inp[0]) ? 4'b0011 : 4'b0001;
														assign node57241 = (inp[9]) ? 4'b0111 : node57242;
															assign node57242 = (inp[15]) ? node57246 : node57243;
																assign node57243 = (inp[0]) ? 4'b0011 : 4'b0001;
																assign node57246 = (inp[0]) ? 4'b0001 : 4'b0011;
													assign node57250 = (inp[9]) ? node57262 : node57251;
														assign node57251 = (inp[4]) ? node57257 : node57252;
															assign node57252 = (inp[15]) ? node57254 : 4'b0001;
																assign node57254 = (inp[0]) ? 4'b0001 : 4'b0011;
															assign node57257 = (inp[15]) ? 4'b0101 : node57258;
																assign node57258 = (inp[0]) ? 4'b0111 : 4'b0101;
														assign node57262 = (inp[4]) ? node57270 : node57263;
															assign node57263 = (inp[0]) ? node57267 : node57264;
																assign node57264 = (inp[15]) ? 4'b0111 : 4'b0101;
																assign node57267 = (inp[15]) ? 4'b0101 : 4'b0111;
															assign node57270 = (inp[0]) ? 4'b0011 : node57271;
																assign node57271 = (inp[15]) ? 4'b0011 : 4'b0001;
										assign node57275 = (inp[4]) ? node57339 : node57276;
											assign node57276 = (inp[9]) ? node57306 : node57277;
												assign node57277 = (inp[0]) ? node57295 : node57278;
													assign node57278 = (inp[3]) ? node57280 : 4'b0001;
														assign node57280 = (inp[12]) ? node57288 : node57281;
															assign node57281 = (inp[5]) ? node57285 : node57282;
																assign node57282 = (inp[15]) ? 4'b0001 : 4'b0011;
																assign node57285 = (inp[15]) ? 4'b0011 : 4'b0001;
															assign node57288 = (inp[15]) ? node57292 : node57289;
																assign node57289 = (inp[5]) ? 4'b0001 : 4'b0011;
																assign node57292 = (inp[5]) ? 4'b0011 : 4'b0001;
													assign node57295 = (inp[15]) ? node57301 : node57296;
														assign node57296 = (inp[5]) ? node57298 : 4'b0001;
															assign node57298 = (inp[3]) ? 4'b0011 : 4'b0001;
														assign node57301 = (inp[5]) ? node57303 : 4'b0011;
															assign node57303 = (inp[3]) ? 4'b0001 : 4'b0011;
												assign node57306 = (inp[5]) ? node57324 : node57307;
													assign node57307 = (inp[12]) ? node57317 : node57308;
														assign node57308 = (inp[15]) ? node57310 : 4'b0101;
															assign node57310 = (inp[3]) ? node57314 : node57311;
																assign node57311 = (inp[0]) ? 4'b0111 : 4'b0101;
																assign node57314 = (inp[0]) ? 4'b0101 : 4'b0111;
														assign node57317 = (inp[3]) ? node57319 : 4'b0101;
															assign node57319 = (inp[15]) ? 4'b0101 : node57320;
																assign node57320 = (inp[0]) ? 4'b0111 : 4'b0101;
													assign node57324 = (inp[3]) ? node57332 : node57325;
														assign node57325 = (inp[15]) ? node57329 : node57326;
															assign node57326 = (inp[0]) ? 4'b0111 : 4'b0101;
															assign node57329 = (inp[0]) ? 4'b0101 : 4'b0111;
														assign node57332 = (inp[15]) ? node57336 : node57333;
															assign node57333 = (inp[0]) ? 4'b0111 : 4'b0101;
															assign node57336 = (inp[0]) ? 4'b0101 : 4'b0111;
											assign node57339 = (inp[9]) ? node57363 : node57340;
												assign node57340 = (inp[0]) ? node57352 : node57341;
													assign node57341 = (inp[15]) ? node57347 : node57342;
														assign node57342 = (inp[5]) ? 4'b0101 : node57343;
															assign node57343 = (inp[3]) ? 4'b0101 : 4'b0111;
														assign node57347 = (inp[5]) ? 4'b0111 : node57348;
															assign node57348 = (inp[3]) ? 4'b0111 : 4'b0101;
													assign node57352 = (inp[15]) ? node57358 : node57353;
														assign node57353 = (inp[5]) ? 4'b0111 : node57354;
															assign node57354 = (inp[3]) ? 4'b0111 : 4'b0101;
														assign node57358 = (inp[3]) ? 4'b0101 : node57359;
															assign node57359 = (inp[5]) ? 4'b0101 : 4'b0111;
												assign node57363 = (inp[15]) ? node57375 : node57364;
													assign node57364 = (inp[0]) ? node57370 : node57365;
														assign node57365 = (inp[5]) ? 4'b0001 : node57366;
															assign node57366 = (inp[3]) ? 4'b0001 : 4'b0011;
														assign node57370 = (inp[3]) ? 4'b0011 : node57371;
															assign node57371 = (inp[5]) ? 4'b0011 : 4'b0001;
													assign node57375 = (inp[0]) ? 4'b0001 : node57376;
														assign node57376 = (inp[5]) ? 4'b0011 : node57377;
															assign node57377 = (inp[3]) ? 4'b0011 : 4'b0001;
									assign node57382 = (inp[5]) ? node57532 : node57383;
										assign node57383 = (inp[4]) ? node57437 : node57384;
											assign node57384 = (inp[9]) ? node57410 : node57385;
												assign node57385 = (inp[12]) ? node57403 : node57386;
													assign node57386 = (inp[10]) ? node57394 : node57387;
														assign node57387 = (inp[3]) ? 4'b0100 : node57388;
															assign node57388 = (inp[15]) ? 4'b0100 : node57389;
																assign node57389 = (inp[0]) ? 4'b0100 : 4'b0110;
														assign node57394 = (inp[3]) ? 4'b0000 : node57395;
															assign node57395 = (inp[15]) ? node57399 : node57396;
																assign node57396 = (inp[0]) ? 4'b0000 : 4'b0010;
																assign node57399 = (inp[0]) ? 4'b0010 : 4'b0000;
													assign node57403 = (inp[15]) ? node57407 : node57404;
														assign node57404 = (inp[0]) ? 4'b0000 : 4'b0010;
														assign node57407 = (inp[0]) ? 4'b0010 : 4'b0000;
												assign node57410 = (inp[12]) ? node57424 : node57411;
													assign node57411 = (inp[10]) ? node57419 : node57412;
														assign node57412 = (inp[3]) ? node57414 : 4'b0000;
															assign node57414 = (inp[15]) ? 4'b0010 : node57415;
																assign node57415 = (inp[0]) ? 4'b0000 : 4'b0010;
														assign node57419 = (inp[3]) ? node57421 : 4'b0100;
															assign node57421 = (inp[15]) ? 4'b0100 : 4'b0110;
													assign node57424 = (inp[15]) ? node57432 : node57425;
														assign node57425 = (inp[3]) ? node57429 : node57426;
															assign node57426 = (inp[0]) ? 4'b0100 : 4'b0110;
															assign node57429 = (inp[0]) ? 4'b0110 : 4'b0100;
														assign node57432 = (inp[3]) ? node57434 : 4'b0110;
															assign node57434 = (inp[0]) ? 4'b0100 : 4'b0110;
											assign node57437 = (inp[9]) ? node57485 : node57438;
												assign node57438 = (inp[12]) ? node57464 : node57439;
													assign node57439 = (inp[10]) ? node57455 : node57440;
														assign node57440 = (inp[3]) ? node57448 : node57441;
															assign node57441 = (inp[15]) ? node57445 : node57442;
																assign node57442 = (inp[0]) ? 4'b0000 : 4'b0010;
																assign node57445 = (inp[0]) ? 4'b0010 : 4'b0000;
															assign node57448 = (inp[0]) ? node57452 : node57449;
																assign node57449 = (inp[15]) ? 4'b0000 : 4'b0010;
																assign node57452 = (inp[15]) ? 4'b0010 : 4'b0000;
														assign node57455 = (inp[0]) ? node57457 : 4'b0100;
															assign node57457 = (inp[15]) ? node57461 : node57458;
																assign node57458 = (inp[3]) ? 4'b0110 : 4'b0100;
																assign node57461 = (inp[3]) ? 4'b0100 : 4'b0110;
													assign node57464 = (inp[15]) ? node57470 : node57465;
														assign node57465 = (inp[10]) ? node57467 : 4'b0100;
															assign node57467 = (inp[3]) ? 4'b0100 : 4'b0110;
														assign node57470 = (inp[10]) ? node57478 : node57471;
															assign node57471 = (inp[3]) ? node57475 : node57472;
																assign node57472 = (inp[0]) ? 4'b0110 : 4'b0100;
																assign node57475 = (inp[0]) ? 4'b0100 : 4'b0110;
															assign node57478 = (inp[0]) ? node57482 : node57479;
																assign node57479 = (inp[3]) ? 4'b0110 : 4'b0100;
																assign node57482 = (inp[3]) ? 4'b0100 : 4'b0110;
												assign node57485 = (inp[12]) ? node57507 : node57486;
													assign node57486 = (inp[10]) ? node57494 : node57487;
														assign node57487 = (inp[3]) ? node57489 : 4'b0110;
															assign node57489 = (inp[15]) ? 4'b0100 : node57490;
																assign node57490 = (inp[0]) ? 4'b0110 : 4'b0100;
														assign node57494 = (inp[15]) ? node57502 : node57495;
															assign node57495 = (inp[0]) ? node57499 : node57496;
																assign node57496 = (inp[3]) ? 4'b0000 : 4'b0010;
																assign node57499 = (inp[3]) ? 4'b0010 : 4'b0000;
															assign node57502 = (inp[0]) ? 4'b0010 : node57503;
																assign node57503 = (inp[3]) ? 4'b0010 : 4'b0000;
													assign node57507 = (inp[10]) ? node57523 : node57508;
														assign node57508 = (inp[15]) ? node57516 : node57509;
															assign node57509 = (inp[3]) ? node57513 : node57510;
																assign node57510 = (inp[0]) ? 4'b0000 : 4'b0010;
																assign node57513 = (inp[0]) ? 4'b0010 : 4'b0000;
															assign node57516 = (inp[0]) ? node57520 : node57517;
																assign node57517 = (inp[3]) ? 4'b0010 : 4'b0000;
																assign node57520 = (inp[3]) ? 4'b0000 : 4'b0010;
														assign node57523 = (inp[3]) ? 4'b0000 : node57524;
															assign node57524 = (inp[15]) ? node57528 : node57525;
																assign node57525 = (inp[0]) ? 4'b0000 : 4'b0010;
																assign node57528 = (inp[0]) ? 4'b0010 : 4'b0000;
										assign node57532 = (inp[12]) ? node57612 : node57533;
											assign node57533 = (inp[4]) ? node57573 : node57534;
												assign node57534 = (inp[9]) ? node57556 : node57535;
													assign node57535 = (inp[10]) ? node57543 : node57536;
														assign node57536 = (inp[3]) ? 4'b0110 : node57537;
															assign node57537 = (inp[0]) ? node57539 : 4'b0100;
																assign node57539 = (inp[15]) ? 4'b0110 : 4'b0100;
														assign node57543 = (inp[3]) ? node57551 : node57544;
															assign node57544 = (inp[15]) ? node57548 : node57545;
																assign node57545 = (inp[0]) ? 4'b0000 : 4'b0010;
																assign node57548 = (inp[0]) ? 4'b0010 : 4'b0000;
															assign node57551 = (inp[15]) ? 4'b0000 : node57552;
																assign node57552 = (inp[0]) ? 4'b0010 : 4'b0000;
													assign node57556 = (inp[10]) ? node57566 : node57557;
														assign node57557 = (inp[3]) ? node57559 : 4'b0000;
															assign node57559 = (inp[15]) ? node57563 : node57560;
																assign node57560 = (inp[0]) ? 4'b0010 : 4'b0000;
																assign node57563 = (inp[0]) ? 4'b0000 : 4'b0010;
														assign node57566 = (inp[0]) ? node57570 : node57567;
															assign node57567 = (inp[15]) ? 4'b0110 : 4'b0100;
															assign node57570 = (inp[15]) ? 4'b0100 : 4'b0110;
												assign node57573 = (inp[0]) ? node57599 : node57574;
													assign node57574 = (inp[15]) ? node57590 : node57575;
														assign node57575 = (inp[3]) ? node57583 : node57576;
															assign node57576 = (inp[10]) ? node57580 : node57577;
																assign node57577 = (inp[9]) ? 4'b0100 : 4'b0010;
																assign node57580 = (inp[9]) ? 4'b0000 : 4'b0100;
															assign node57583 = (inp[10]) ? node57587 : node57584;
																assign node57584 = (inp[9]) ? 4'b0100 : 4'b0000;
																assign node57587 = (inp[9]) ? 4'b0000 : 4'b0100;
														assign node57590 = (inp[9]) ? node57596 : node57591;
															assign node57591 = (inp[10]) ? 4'b0110 : node57592;
																assign node57592 = (inp[3]) ? 4'b0010 : 4'b0000;
															assign node57596 = (inp[10]) ? 4'b0010 : 4'b0110;
													assign node57599 = (inp[15]) ? node57607 : node57600;
														assign node57600 = (inp[10]) ? node57604 : node57601;
															assign node57601 = (inp[9]) ? 4'b0110 : 4'b0000;
															assign node57604 = (inp[9]) ? 4'b0010 : 4'b0110;
														assign node57607 = (inp[9]) ? node57609 : 4'b0100;
															assign node57609 = (inp[10]) ? 4'b0000 : 4'b0100;
											assign node57612 = (inp[15]) ? node57636 : node57613;
												assign node57613 = (inp[0]) ? node57619 : node57614;
													assign node57614 = (inp[9]) ? 4'b0100 : node57615;
														assign node57615 = (inp[4]) ? 4'b0100 : 4'b0000;
													assign node57619 = (inp[3]) ? node57629 : node57620;
														assign node57620 = (inp[10]) ? node57622 : 4'b0110;
															assign node57622 = (inp[9]) ? node57626 : node57623;
																assign node57623 = (inp[4]) ? 4'b0110 : 4'b0000;
																assign node57626 = (inp[4]) ? 4'b0010 : 4'b0110;
														assign node57629 = (inp[9]) ? node57633 : node57630;
															assign node57630 = (inp[4]) ? 4'b0110 : 4'b0010;
															assign node57633 = (inp[4]) ? 4'b0010 : 4'b0110;
												assign node57636 = (inp[0]) ? node57652 : node57637;
													assign node57637 = (inp[3]) ? node57645 : node57638;
														assign node57638 = (inp[9]) ? node57642 : node57639;
															assign node57639 = (inp[4]) ? 4'b0110 : 4'b0000;
															assign node57642 = (inp[4]) ? 4'b0010 : 4'b0110;
														assign node57645 = (inp[9]) ? node57649 : node57646;
															assign node57646 = (inp[4]) ? 4'b0110 : 4'b0010;
															assign node57649 = (inp[4]) ? 4'b0010 : 4'b0110;
													assign node57652 = (inp[3]) ? node57660 : node57653;
														assign node57653 = (inp[9]) ? node57657 : node57654;
															assign node57654 = (inp[4]) ? 4'b0100 : 4'b0010;
															assign node57657 = (inp[4]) ? 4'b0000 : 4'b0100;
														assign node57660 = (inp[9]) ? node57664 : node57661;
															assign node57661 = (inp[4]) ? 4'b0100 : 4'b0000;
															assign node57664 = (inp[4]) ? 4'b0000 : 4'b0100;
								assign node57667 = (inp[5]) ? node57875 : node57668;
									assign node57668 = (inp[0]) ? node57776 : node57669;
										assign node57669 = (inp[15]) ? node57715 : node57670;
											assign node57670 = (inp[3]) ? node57698 : node57671;
												assign node57671 = (inp[12]) ? node57689 : node57672;
													assign node57672 = (inp[10]) ? node57680 : node57673;
														assign node57673 = (inp[4]) ? node57677 : node57674;
															assign node57674 = (inp[9]) ? 4'b0010 : 4'b0110;
															assign node57677 = (inp[9]) ? 4'b0110 : 4'b0010;
														assign node57680 = (inp[14]) ? 4'b0010 : node57681;
															assign node57681 = (inp[9]) ? node57685 : node57682;
																assign node57682 = (inp[4]) ? 4'b0110 : 4'b0010;
																assign node57685 = (inp[4]) ? 4'b0010 : 4'b0110;
													assign node57689 = (inp[10]) ? node57691 : 4'b0110;
														assign node57691 = (inp[14]) ? 4'b0110 : node57692;
															assign node57692 = (inp[9]) ? node57694 : 4'b0010;
																assign node57694 = (inp[4]) ? 4'b0010 : 4'b0110;
												assign node57698 = (inp[9]) ? node57706 : node57699;
													assign node57699 = (inp[4]) ? 4'b0100 : node57700;
														assign node57700 = (inp[10]) ? 4'b0010 : node57701;
															assign node57701 = (inp[12]) ? 4'b0010 : 4'b0110;
													assign node57706 = (inp[10]) ? node57712 : node57707;
														assign node57707 = (inp[4]) ? 4'b0100 : node57708;
															assign node57708 = (inp[12]) ? 4'b0100 : 4'b0010;
														assign node57712 = (inp[4]) ? 4'b0000 : 4'b0100;
											assign node57715 = (inp[3]) ? node57753 : node57716;
												assign node57716 = (inp[12]) ? node57746 : node57717;
													assign node57717 = (inp[4]) ? node57733 : node57718;
														assign node57718 = (inp[14]) ? node57726 : node57719;
															assign node57719 = (inp[10]) ? node57723 : node57720;
																assign node57720 = (inp[9]) ? 4'b0000 : 4'b0100;
																assign node57723 = (inp[9]) ? 4'b0100 : 4'b0000;
															assign node57726 = (inp[9]) ? node57730 : node57727;
																assign node57727 = (inp[10]) ? 4'b0000 : 4'b0100;
																assign node57730 = (inp[10]) ? 4'b0100 : 4'b0000;
														assign node57733 = (inp[14]) ? node57739 : node57734;
															assign node57734 = (inp[10]) ? node57736 : 4'b0100;
																assign node57736 = (inp[9]) ? 4'b0000 : 4'b0100;
															assign node57739 = (inp[9]) ? node57743 : node57740;
																assign node57740 = (inp[10]) ? 4'b0100 : 4'b0000;
																assign node57743 = (inp[10]) ? 4'b0000 : 4'b0100;
													assign node57746 = (inp[4]) ? node57750 : node57747;
														assign node57747 = (inp[9]) ? 4'b0100 : 4'b0000;
														assign node57750 = (inp[9]) ? 4'b0000 : 4'b0100;
												assign node57753 = (inp[4]) ? node57765 : node57754;
													assign node57754 = (inp[9]) ? node57760 : node57755;
														assign node57755 = (inp[10]) ? 4'b0000 : node57756;
															assign node57756 = (inp[12]) ? 4'b0000 : 4'b0100;
														assign node57760 = (inp[10]) ? 4'b0110 : node57761;
															assign node57761 = (inp[12]) ? 4'b0110 : 4'b0000;
													assign node57765 = (inp[9]) ? node57771 : node57766;
														assign node57766 = (inp[12]) ? 4'b0110 : node57767;
															assign node57767 = (inp[10]) ? 4'b0110 : 4'b0000;
														assign node57771 = (inp[10]) ? 4'b0010 : node57772;
															assign node57772 = (inp[14]) ? 4'b0110 : 4'b0010;
										assign node57776 = (inp[15]) ? node57832 : node57777;
											assign node57777 = (inp[3]) ? node57813 : node57778;
												assign node57778 = (inp[14]) ? node57796 : node57779;
													assign node57779 = (inp[9]) ? node57787 : node57780;
														assign node57780 = (inp[4]) ? node57784 : node57781;
															assign node57781 = (inp[12]) ? 4'b0000 : 4'b0100;
															assign node57784 = (inp[12]) ? 4'b0100 : 4'b0000;
														assign node57787 = (inp[4]) ? node57791 : node57788;
															assign node57788 = (inp[12]) ? 4'b0100 : 4'b0000;
															assign node57791 = (inp[10]) ? 4'b0000 : node57792;
																assign node57792 = (inp[12]) ? 4'b0000 : 4'b0100;
													assign node57796 = (inp[12]) ? node57808 : node57797;
														assign node57797 = (inp[10]) ? node57803 : node57798;
															assign node57798 = (inp[9]) ? 4'b0000 : node57799;
																assign node57799 = (inp[4]) ? 4'b0000 : 4'b0100;
															assign node57803 = (inp[4]) ? 4'b0100 : node57804;
																assign node57804 = (inp[9]) ? 4'b0100 : 4'b0000;
														assign node57808 = (inp[4]) ? node57810 : 4'b0100;
															assign node57810 = (inp[9]) ? 4'b0000 : 4'b0100;
												assign node57813 = (inp[9]) ? node57825 : node57814;
													assign node57814 = (inp[4]) ? node57820 : node57815;
														assign node57815 = (inp[12]) ? 4'b0000 : node57816;
															assign node57816 = (inp[10]) ? 4'b0000 : 4'b0100;
														assign node57820 = (inp[12]) ? 4'b0110 : node57821;
															assign node57821 = (inp[10]) ? 4'b0110 : 4'b0000;
													assign node57825 = (inp[4]) ? 4'b0010 : node57826;
														assign node57826 = (inp[12]) ? 4'b0110 : node57827;
															assign node57827 = (inp[10]) ? 4'b0110 : 4'b0000;
											assign node57832 = (inp[3]) ? node57852 : node57833;
												assign node57833 = (inp[4]) ? node57841 : node57834;
													assign node57834 = (inp[9]) ? node57836 : 4'b0010;
														assign node57836 = (inp[10]) ? 4'b0110 : node57837;
															assign node57837 = (inp[12]) ? 4'b0110 : 4'b0010;
													assign node57841 = (inp[9]) ? node57847 : node57842;
														assign node57842 = (inp[12]) ? 4'b0110 : node57843;
															assign node57843 = (inp[10]) ? 4'b0110 : 4'b0010;
														assign node57847 = (inp[10]) ? 4'b0010 : node57848;
															assign node57848 = (inp[12]) ? 4'b0010 : 4'b0110;
												assign node57852 = (inp[9]) ? node57864 : node57853;
													assign node57853 = (inp[4]) ? node57859 : node57854;
														assign node57854 = (inp[10]) ? 4'b0010 : node57855;
															assign node57855 = (inp[12]) ? 4'b0010 : 4'b0110;
														assign node57859 = (inp[10]) ? 4'b0100 : node57860;
															assign node57860 = (inp[12]) ? 4'b0100 : 4'b0010;
													assign node57864 = (inp[4]) ? node57870 : node57865;
														assign node57865 = (inp[10]) ? 4'b0100 : node57866;
															assign node57866 = (inp[12]) ? 4'b0100 : 4'b0010;
														assign node57870 = (inp[12]) ? 4'b0000 : node57871;
															assign node57871 = (inp[10]) ? 4'b0000 : 4'b0100;
									assign node57875 = (inp[12]) ? node58009 : node57876;
										assign node57876 = (inp[4]) ? node57944 : node57877;
											assign node57877 = (inp[0]) ? node57907 : node57878;
												assign node57878 = (inp[15]) ? node57894 : node57879;
													assign node57879 = (inp[3]) ? node57887 : node57880;
														assign node57880 = (inp[10]) ? node57884 : node57881;
															assign node57881 = (inp[9]) ? 4'b0010 : 4'b0110;
															assign node57884 = (inp[9]) ? 4'b0100 : 4'b0010;
														assign node57887 = (inp[9]) ? node57891 : node57888;
															assign node57888 = (inp[10]) ? 4'b0000 : 4'b0100;
															assign node57891 = (inp[10]) ? 4'b0100 : 4'b0000;
													assign node57894 = (inp[3]) ? node57902 : node57895;
														assign node57895 = (inp[10]) ? node57899 : node57896;
															assign node57896 = (inp[9]) ? 4'b0000 : 4'b0100;
															assign node57899 = (inp[9]) ? 4'b0110 : 4'b0000;
														assign node57902 = (inp[9]) ? 4'b0110 : node57903;
															assign node57903 = (inp[10]) ? 4'b0010 : 4'b0110;
												assign node57907 = (inp[15]) ? node57923 : node57908;
													assign node57908 = (inp[3]) ? node57916 : node57909;
														assign node57909 = (inp[9]) ? node57913 : node57910;
															assign node57910 = (inp[10]) ? 4'b0000 : 4'b0100;
															assign node57913 = (inp[10]) ? 4'b0110 : 4'b0000;
														assign node57916 = (inp[10]) ? node57920 : node57917;
															assign node57917 = (inp[9]) ? 4'b0010 : 4'b0110;
															assign node57920 = (inp[9]) ? 4'b0110 : 4'b0010;
													assign node57923 = (inp[3]) ? node57931 : node57924;
														assign node57924 = (inp[10]) ? node57928 : node57925;
															assign node57925 = (inp[9]) ? 4'b0010 : 4'b0110;
															assign node57928 = (inp[9]) ? 4'b0100 : 4'b0010;
														assign node57931 = (inp[14]) ? node57939 : node57932;
															assign node57932 = (inp[9]) ? node57936 : node57933;
																assign node57933 = (inp[10]) ? 4'b0000 : 4'b0100;
																assign node57936 = (inp[10]) ? 4'b0100 : 4'b0000;
															assign node57939 = (inp[10]) ? node57941 : 4'b0000;
																assign node57941 = (inp[9]) ? 4'b0100 : 4'b0000;
											assign node57944 = (inp[10]) ? node57984 : node57945;
												assign node57945 = (inp[9]) ? node57963 : node57946;
													assign node57946 = (inp[15]) ? node57954 : node57947;
														assign node57947 = (inp[3]) ? node57951 : node57948;
															assign node57948 = (inp[0]) ? 4'b0000 : 4'b0010;
															assign node57951 = (inp[0]) ? 4'b0010 : 4'b0000;
														assign node57954 = (inp[14]) ? node57956 : 4'b0010;
															assign node57956 = (inp[0]) ? node57960 : node57957;
																assign node57957 = (inp[3]) ? 4'b0010 : 4'b0000;
																assign node57960 = (inp[3]) ? 4'b0000 : 4'b0010;
													assign node57963 = (inp[3]) ? node57979 : node57964;
														assign node57964 = (inp[14]) ? node57972 : node57965;
															assign node57965 = (inp[0]) ? node57969 : node57966;
																assign node57966 = (inp[15]) ? 4'b0110 : 4'b0100;
																assign node57969 = (inp[15]) ? 4'b0100 : 4'b0110;
															assign node57972 = (inp[0]) ? node57976 : node57973;
																assign node57973 = (inp[15]) ? 4'b0110 : 4'b0100;
																assign node57976 = (inp[15]) ? 4'b0100 : 4'b0110;
														assign node57979 = (inp[14]) ? 4'b0110 : node57980;
															assign node57980 = (inp[0]) ? 4'b0100 : 4'b0110;
												assign node57984 = (inp[9]) ? node57992 : node57985;
													assign node57985 = (inp[0]) ? node57989 : node57986;
														assign node57986 = (inp[15]) ? 4'b0110 : 4'b0100;
														assign node57989 = (inp[15]) ? 4'b0100 : 4'b0110;
													assign node57992 = (inp[3]) ? node58000 : node57993;
														assign node57993 = (inp[15]) ? node57997 : node57994;
															assign node57994 = (inp[0]) ? 4'b0010 : 4'b0000;
															assign node57997 = (inp[0]) ? 4'b0000 : 4'b0010;
														assign node58000 = (inp[14]) ? node58006 : node58001;
															assign node58001 = (inp[15]) ? node58003 : 4'b0010;
																assign node58003 = (inp[0]) ? 4'b0000 : 4'b0010;
															assign node58006 = (inp[15]) ? 4'b0010 : 4'b0000;
										assign node58009 = (inp[15]) ? node58029 : node58010;
											assign node58010 = (inp[0]) ? node58020 : node58011;
												assign node58011 = (inp[4]) ? node58017 : node58012;
													assign node58012 = (inp[9]) ? 4'b0100 : node58013;
														assign node58013 = (inp[3]) ? 4'b0000 : 4'b0010;
													assign node58017 = (inp[9]) ? 4'b0000 : 4'b0100;
												assign node58020 = (inp[9]) ? node58026 : node58021;
													assign node58021 = (inp[4]) ? 4'b0110 : node58022;
														assign node58022 = (inp[3]) ? 4'b0010 : 4'b0000;
													assign node58026 = (inp[4]) ? 4'b0010 : 4'b0110;
											assign node58029 = (inp[0]) ? node58039 : node58030;
												assign node58030 = (inp[9]) ? node58036 : node58031;
													assign node58031 = (inp[4]) ? 4'b0110 : node58032;
														assign node58032 = (inp[3]) ? 4'b0010 : 4'b0000;
													assign node58036 = (inp[4]) ? 4'b0010 : 4'b0110;
												assign node58039 = (inp[3]) ? node58045 : node58040;
													assign node58040 = (inp[4]) ? 4'b0100 : node58041;
														assign node58041 = (inp[9]) ? 4'b0100 : 4'b0010;
													assign node58045 = (inp[9]) ? node58049 : node58046;
														assign node58046 = (inp[4]) ? 4'b0100 : 4'b0000;
														assign node58049 = (inp[4]) ? 4'b0000 : 4'b0100;
				assign node58052 = (inp[13]) ? node62116 : node58053;
					assign node58053 = (inp[8]) ? node60143 : node58054;
						assign node58054 = (inp[7]) ? node59178 : node58055;
							assign node58055 = (inp[2]) ? node58643 : node58056;
								assign node58056 = (inp[14]) ? node58356 : node58057;
									assign node58057 = (inp[3]) ? node58199 : node58058;
										assign node58058 = (inp[10]) ? node58138 : node58059;
											assign node58059 = (inp[9]) ? node58097 : node58060;
												assign node58060 = (inp[0]) ? node58078 : node58061;
													assign node58061 = (inp[15]) ? node58069 : node58062;
														assign node58062 = (inp[12]) ? node58066 : node58063;
															assign node58063 = (inp[4]) ? 4'b1011 : 4'b1111;
															assign node58066 = (inp[4]) ? 4'b1101 : 4'b1011;
														assign node58069 = (inp[4]) ? node58073 : node58070;
															assign node58070 = (inp[12]) ? 4'b1001 : 4'b1101;
															assign node58073 = (inp[12]) ? node58075 : 4'b1001;
																assign node58075 = (inp[5]) ? 4'b1111 : 4'b1101;
													assign node58078 = (inp[15]) ? node58088 : node58079;
														assign node58079 = (inp[5]) ? node58085 : node58080;
															assign node58080 = (inp[4]) ? node58082 : 4'b1001;
																assign node58082 = (inp[12]) ? 4'b1101 : 4'b1001;
															assign node58085 = (inp[4]) ? 4'b1111 : 4'b1101;
														assign node58088 = (inp[12]) ? node58092 : node58089;
															assign node58089 = (inp[4]) ? 4'b1011 : 4'b1111;
															assign node58092 = (inp[5]) ? 4'b1101 : node58093;
																assign node58093 = (inp[4]) ? 4'b1111 : 4'b1011;
												assign node58097 = (inp[5]) ? node58123 : node58098;
													assign node58098 = (inp[15]) ? node58112 : node58099;
														assign node58099 = (inp[0]) ? node58105 : node58100;
															assign node58100 = (inp[4]) ? node58102 : 4'b1111;
																assign node58102 = (inp[12]) ? 4'b1011 : 4'b1111;
															assign node58105 = (inp[4]) ? node58109 : node58106;
																assign node58106 = (inp[12]) ? 4'b1101 : 4'b1001;
																assign node58109 = (inp[12]) ? 4'b1001 : 4'b1101;
														assign node58112 = (inp[0]) ? node58116 : node58113;
															assign node58113 = (inp[12]) ? 4'b1001 : 4'b1101;
															assign node58116 = (inp[12]) ? node58120 : node58117;
																assign node58117 = (inp[4]) ? 4'b1111 : 4'b1011;
																assign node58120 = (inp[4]) ? 4'b1011 : 4'b1111;
													assign node58123 = (inp[12]) ? node58131 : node58124;
														assign node58124 = (inp[4]) ? node58126 : 4'b1011;
															assign node58126 = (inp[15]) ? 4'b1111 : node58127;
																assign node58127 = (inp[0]) ? 4'b1111 : 4'b1101;
														assign node58131 = (inp[4]) ? 4'b1011 : node58132;
															assign node58132 = (inp[0]) ? node58134 : 4'b1111;
																assign node58134 = (inp[15]) ? 4'b1101 : 4'b1111;
											assign node58138 = (inp[12]) ? node58176 : node58139;
												assign node58139 = (inp[4]) ? node58159 : node58140;
													assign node58140 = (inp[9]) ? node58146 : node58141;
														assign node58141 = (inp[15]) ? node58143 : 4'b1011;
															assign node58143 = (inp[0]) ? 4'b1011 : 4'b1001;
														assign node58146 = (inp[5]) ? node58152 : node58147;
															assign node58147 = (inp[0]) ? 4'b1111 : node58148;
																assign node58148 = (inp[15]) ? 4'b1101 : 4'b1111;
															assign node58152 = (inp[15]) ? node58156 : node58153;
																assign node58153 = (inp[0]) ? 4'b1111 : 4'b1101;
																assign node58156 = (inp[0]) ? 4'b1101 : 4'b1111;
													assign node58159 = (inp[9]) ? node58167 : node58160;
														assign node58160 = (inp[15]) ? node58162 : 4'b1101;
															assign node58162 = (inp[5]) ? node58164 : 4'b1111;
																assign node58164 = (inp[0]) ? 4'b1101 : 4'b1111;
														assign node58167 = (inp[0]) ? node58169 : 4'b1011;
															assign node58169 = (inp[15]) ? node58173 : node58170;
																assign node58170 = (inp[5]) ? 4'b1011 : 4'b1001;
																assign node58173 = (inp[5]) ? 4'b1001 : 4'b1011;
												assign node58176 = (inp[4]) ? node58188 : node58177;
													assign node58177 = (inp[9]) ? node58185 : node58178;
														assign node58178 = (inp[0]) ? node58182 : node58179;
															assign node58179 = (inp[15]) ? 4'b1001 : 4'b1011;
															assign node58182 = (inp[15]) ? 4'b1011 : 4'b1001;
														assign node58185 = (inp[15]) ? 4'b1111 : 4'b1101;
													assign node58188 = (inp[9]) ? node58190 : 4'b1111;
														assign node58190 = (inp[0]) ? 4'b1011 : node58191;
															assign node58191 = (inp[15]) ? node58195 : node58192;
																assign node58192 = (inp[5]) ? 4'b1001 : 4'b1011;
																assign node58195 = (inp[5]) ? 4'b1011 : 4'b1001;
										assign node58199 = (inp[9]) ? node58293 : node58200;
											assign node58200 = (inp[4]) ? node58244 : node58201;
												assign node58201 = (inp[12]) ? node58227 : node58202;
													assign node58202 = (inp[10]) ? node58218 : node58203;
														assign node58203 = (inp[0]) ? node58211 : node58204;
															assign node58204 = (inp[5]) ? node58208 : node58205;
																assign node58205 = (inp[15]) ? 4'b1101 : 4'b1111;
																assign node58208 = (inp[15]) ? 4'b1111 : 4'b1101;
															assign node58211 = (inp[15]) ? node58215 : node58212;
																assign node58212 = (inp[5]) ? 4'b1111 : 4'b1101;
																assign node58215 = (inp[5]) ? 4'b1101 : 4'b1111;
														assign node58218 = (inp[15]) ? 4'b1011 : node58219;
															assign node58219 = (inp[0]) ? node58223 : node58220;
																assign node58220 = (inp[5]) ? 4'b1001 : 4'b1011;
																assign node58223 = (inp[5]) ? 4'b1011 : 4'b1001;
													assign node58227 = (inp[0]) ? node58237 : node58228;
														assign node58228 = (inp[10]) ? node58234 : node58229;
															assign node58229 = (inp[5]) ? 4'b1011 : node58230;
																assign node58230 = (inp[15]) ? 4'b1001 : 4'b1011;
															assign node58234 = (inp[5]) ? 4'b1001 : 4'b1011;
														assign node58237 = (inp[10]) ? 4'b1011 : node58238;
															assign node58238 = (inp[15]) ? 4'b1011 : node58239;
																assign node58239 = (inp[5]) ? 4'b1011 : 4'b1001;
												assign node58244 = (inp[10]) ? node58270 : node58245;
													assign node58245 = (inp[12]) ? node58259 : node58246;
														assign node58246 = (inp[0]) ? node58254 : node58247;
															assign node58247 = (inp[5]) ? node58251 : node58248;
																assign node58248 = (inp[15]) ? 4'b1001 : 4'b1011;
																assign node58251 = (inp[15]) ? 4'b1011 : 4'b1001;
															assign node58254 = (inp[15]) ? node58256 : 4'b1001;
																assign node58256 = (inp[5]) ? 4'b1001 : 4'b1011;
														assign node58259 = (inp[5]) ? node58265 : node58260;
															assign node58260 = (inp[0]) ? node58262 : 4'b1101;
																assign node58262 = (inp[15]) ? 4'b1101 : 4'b1111;
															assign node58265 = (inp[15]) ? 4'b1111 : node58266;
																assign node58266 = (inp[0]) ? 4'b1111 : 4'b1101;
													assign node58270 = (inp[12]) ? node58278 : node58271;
														assign node58271 = (inp[15]) ? node58275 : node58272;
															assign node58272 = (inp[0]) ? 4'b1111 : 4'b1101;
															assign node58275 = (inp[0]) ? 4'b1101 : 4'b1111;
														assign node58278 = (inp[5]) ? node58286 : node58279;
															assign node58279 = (inp[0]) ? node58283 : node58280;
																assign node58280 = (inp[15]) ? 4'b1111 : 4'b1101;
																assign node58283 = (inp[15]) ? 4'b1101 : 4'b1111;
															assign node58286 = (inp[15]) ? node58290 : node58287;
																assign node58287 = (inp[0]) ? 4'b1111 : 4'b1101;
																assign node58290 = (inp[0]) ? 4'b1101 : 4'b1111;
											assign node58293 = (inp[4]) ? node58339 : node58294;
												assign node58294 = (inp[10]) ? node58318 : node58295;
													assign node58295 = (inp[12]) ? node58311 : node58296;
														assign node58296 = (inp[15]) ? node58304 : node58297;
															assign node58297 = (inp[5]) ? node58301 : node58298;
																assign node58298 = (inp[0]) ? 4'b1001 : 4'b1011;
																assign node58301 = (inp[0]) ? 4'b1011 : 4'b1001;
															assign node58304 = (inp[0]) ? node58308 : node58305;
																assign node58305 = (inp[5]) ? 4'b1011 : 4'b1001;
																assign node58308 = (inp[5]) ? 4'b1001 : 4'b1011;
														assign node58311 = (inp[5]) ? 4'b1101 : node58312;
															assign node58312 = (inp[0]) ? node58314 : 4'b1111;
																assign node58314 = (inp[15]) ? 4'b1101 : 4'b1111;
													assign node58318 = (inp[12]) ? node58334 : node58319;
														assign node58319 = (inp[5]) ? node58327 : node58320;
															assign node58320 = (inp[0]) ? node58324 : node58321;
																assign node58321 = (inp[15]) ? 4'b1111 : 4'b1101;
																assign node58324 = (inp[15]) ? 4'b1101 : 4'b1111;
															assign node58327 = (inp[0]) ? node58331 : node58328;
																assign node58328 = (inp[15]) ? 4'b1111 : 4'b1101;
																assign node58331 = (inp[15]) ? 4'b1101 : 4'b1111;
														assign node58334 = (inp[0]) ? 4'b1101 : node58335;
															assign node58335 = (inp[15]) ? 4'b1111 : 4'b1101;
												assign node58339 = (inp[12]) ? node58349 : node58340;
													assign node58340 = (inp[10]) ? node58342 : 4'b1111;
														assign node58342 = (inp[0]) ? node58346 : node58343;
															assign node58343 = (inp[15]) ? 4'b1011 : 4'b1001;
															assign node58346 = (inp[15]) ? 4'b1001 : 4'b1011;
													assign node58349 = (inp[0]) ? node58353 : node58350;
														assign node58350 = (inp[15]) ? 4'b1011 : 4'b1001;
														assign node58353 = (inp[15]) ? 4'b1001 : 4'b1011;
									assign node58356 = (inp[12]) ? node58524 : node58357;
										assign node58357 = (inp[4]) ? node58443 : node58358;
											assign node58358 = (inp[5]) ? node58396 : node58359;
												assign node58359 = (inp[0]) ? node58377 : node58360;
													assign node58360 = (inp[15]) ? node58368 : node58361;
														assign node58361 = (inp[10]) ? node58365 : node58362;
															assign node58362 = (inp[9]) ? 4'b1010 : 4'b1110;
															assign node58365 = (inp[9]) ? 4'b1100 : 4'b1010;
														assign node58368 = (inp[10]) ? node58372 : node58369;
															assign node58369 = (inp[9]) ? 4'b1000 : 4'b1100;
															assign node58372 = (inp[9]) ? node58374 : 4'b1000;
																assign node58374 = (inp[3]) ? 4'b1110 : 4'b1100;
													assign node58377 = (inp[15]) ? node58385 : node58378;
														assign node58378 = (inp[3]) ? 4'b1110 : node58379;
															assign node58379 = (inp[10]) ? 4'b1100 : node58380;
																assign node58380 = (inp[9]) ? 4'b1000 : 4'b1100;
														assign node58385 = (inp[3]) ? node58391 : node58386;
															assign node58386 = (inp[9]) ? 4'b1110 : node58387;
																assign node58387 = (inp[10]) ? 4'b1010 : 4'b1110;
															assign node58391 = (inp[9]) ? 4'b1010 : node58392;
																assign node58392 = (inp[10]) ? 4'b1010 : 4'b1110;
												assign node58396 = (inp[0]) ? node58420 : node58397;
													assign node58397 = (inp[3]) ? node58411 : node58398;
														assign node58398 = (inp[15]) ? node58406 : node58399;
															assign node58399 = (inp[9]) ? node58403 : node58400;
																assign node58400 = (inp[10]) ? 4'b1010 : 4'b1110;
																assign node58403 = (inp[10]) ? 4'b1100 : 4'b1010;
															assign node58406 = (inp[10]) ? node58408 : 4'b1000;
																assign node58408 = (inp[9]) ? 4'b1110 : 4'b1000;
														assign node58411 = (inp[15]) ? node58413 : 4'b1000;
															assign node58413 = (inp[10]) ? node58417 : node58414;
																assign node58414 = (inp[9]) ? 4'b1010 : 4'b1110;
																assign node58417 = (inp[9]) ? 4'b1110 : 4'b1010;
													assign node58420 = (inp[3]) ? node58434 : node58421;
														assign node58421 = (inp[15]) ? node58429 : node58422;
															assign node58422 = (inp[9]) ? node58426 : node58423;
																assign node58423 = (inp[10]) ? 4'b1000 : 4'b1100;
																assign node58426 = (inp[10]) ? 4'b1110 : 4'b1000;
															assign node58429 = (inp[10]) ? 4'b1010 : node58430;
																assign node58430 = (inp[9]) ? 4'b1010 : 4'b1110;
														assign node58434 = (inp[15]) ? node58438 : node58435;
															assign node58435 = (inp[10]) ? 4'b1110 : 4'b1010;
															assign node58438 = (inp[10]) ? node58440 : 4'b1000;
																assign node58440 = (inp[9]) ? 4'b1100 : 4'b1000;
											assign node58443 = (inp[3]) ? node58489 : node58444;
												assign node58444 = (inp[10]) ? node58466 : node58445;
													assign node58445 = (inp[9]) ? node58459 : node58446;
														assign node58446 = (inp[5]) ? node58454 : node58447;
															assign node58447 = (inp[0]) ? node58451 : node58448;
																assign node58448 = (inp[15]) ? 4'b1000 : 4'b1010;
																assign node58451 = (inp[15]) ? 4'b1010 : 4'b1000;
															assign node58454 = (inp[0]) ? 4'b1010 : node58455;
																assign node58455 = (inp[15]) ? 4'b1000 : 4'b1010;
														assign node58459 = (inp[0]) ? 4'b1100 : node58460;
															assign node58460 = (inp[5]) ? node58462 : 4'b1110;
																assign node58462 = (inp[15]) ? 4'b1110 : 4'b1100;
													assign node58466 = (inp[9]) ? node58480 : node58467;
														assign node58467 = (inp[15]) ? node58473 : node58468;
															assign node58468 = (inp[0]) ? 4'b1100 : node58469;
																assign node58469 = (inp[5]) ? 4'b1100 : 4'b1110;
															assign node58473 = (inp[5]) ? node58477 : node58474;
																assign node58474 = (inp[0]) ? 4'b1110 : 4'b1100;
																assign node58477 = (inp[0]) ? 4'b1100 : 4'b1110;
														assign node58480 = (inp[0]) ? 4'b1010 : node58481;
															assign node58481 = (inp[5]) ? node58485 : node58482;
																assign node58482 = (inp[15]) ? 4'b1000 : 4'b1010;
																assign node58485 = (inp[15]) ? 4'b1010 : 4'b1000;
												assign node58489 = (inp[9]) ? node58507 : node58490;
													assign node58490 = (inp[10]) ? node58502 : node58491;
														assign node58491 = (inp[15]) ? node58497 : node58492;
															assign node58492 = (inp[0]) ? 4'b1000 : node58493;
																assign node58493 = (inp[5]) ? 4'b1000 : 4'b1010;
															assign node58497 = (inp[5]) ? 4'b1010 : node58498;
																assign node58498 = (inp[0]) ? 4'b1010 : 4'b1000;
														assign node58502 = (inp[15]) ? node58504 : 4'b1100;
															assign node58504 = (inp[0]) ? 4'b1100 : 4'b1110;
													assign node58507 = (inp[10]) ? node58521 : node58508;
														assign node58508 = (inp[5]) ? node58514 : node58509;
															assign node58509 = (inp[0]) ? node58511 : 4'b1100;
																assign node58511 = (inp[15]) ? 4'b1100 : 4'b1110;
															assign node58514 = (inp[0]) ? node58518 : node58515;
																assign node58515 = (inp[15]) ? 4'b1110 : 4'b1100;
																assign node58518 = (inp[15]) ? 4'b1100 : 4'b1110;
														assign node58521 = (inp[15]) ? 4'b1000 : 4'b1010;
										assign node58524 = (inp[0]) ? node58596 : node58525;
											assign node58525 = (inp[10]) ? node58561 : node58526;
												assign node58526 = (inp[5]) ? node58552 : node58527;
													assign node58527 = (inp[15]) ? node58539 : node58528;
														assign node58528 = (inp[3]) ? node58534 : node58529;
															assign node58529 = (inp[4]) ? node58531 : 4'b1010;
																assign node58531 = (inp[9]) ? 4'b1010 : 4'b1110;
															assign node58534 = (inp[9]) ? node58536 : 4'b1010;
																assign node58536 = (inp[4]) ? 4'b1000 : 4'b1100;
														assign node58539 = (inp[3]) ? node58545 : node58540;
															assign node58540 = (inp[9]) ? 4'b1000 : node58541;
																assign node58541 = (inp[4]) ? 4'b1100 : 4'b1000;
															assign node58545 = (inp[4]) ? node58549 : node58546;
																assign node58546 = (inp[9]) ? 4'b1110 : 4'b1000;
																assign node58549 = (inp[9]) ? 4'b1010 : 4'b1110;
													assign node58552 = (inp[15]) ? 4'b1110 : node58553;
														assign node58553 = (inp[9]) ? 4'b1100 : node58554;
															assign node58554 = (inp[4]) ? 4'b1100 : node58555;
																assign node58555 = (inp[3]) ? 4'b1000 : 4'b1010;
												assign node58561 = (inp[9]) ? node58579 : node58562;
													assign node58562 = (inp[4]) ? node58570 : node58563;
														assign node58563 = (inp[15]) ? 4'b1000 : node58564;
															assign node58564 = (inp[5]) ? node58566 : 4'b1010;
																assign node58566 = (inp[3]) ? 4'b1000 : 4'b1010;
														assign node58570 = (inp[3]) ? 4'b1100 : node58571;
															assign node58571 = (inp[15]) ? node58575 : node58572;
																assign node58572 = (inp[5]) ? 4'b1100 : 4'b1110;
																assign node58575 = (inp[5]) ? 4'b1110 : 4'b1100;
													assign node58579 = (inp[4]) ? node58585 : node58580;
														assign node58580 = (inp[3]) ? 4'b1110 : node58581;
															assign node58581 = (inp[5]) ? 4'b1110 : 4'b1100;
														assign node58585 = (inp[15]) ? node58591 : node58586;
															assign node58586 = (inp[5]) ? 4'b1000 : node58587;
																assign node58587 = (inp[3]) ? 4'b1000 : 4'b1010;
															assign node58591 = (inp[3]) ? 4'b1010 : node58592;
																assign node58592 = (inp[5]) ? 4'b1010 : 4'b1000;
											assign node58596 = (inp[15]) ? node58618 : node58597;
												assign node58597 = (inp[3]) ? node58611 : node58598;
													assign node58598 = (inp[5]) ? node58606 : node58599;
														assign node58599 = (inp[4]) ? node58603 : node58600;
															assign node58600 = (inp[9]) ? 4'b1100 : 4'b1000;
															assign node58603 = (inp[9]) ? 4'b1000 : 4'b1100;
														assign node58606 = (inp[9]) ? node58608 : 4'b1000;
															assign node58608 = (inp[4]) ? 4'b1010 : 4'b1110;
													assign node58611 = (inp[9]) ? node58615 : node58612;
														assign node58612 = (inp[4]) ? 4'b1110 : 4'b1000;
														assign node58615 = (inp[4]) ? 4'b1010 : 4'b1110;
												assign node58618 = (inp[3]) ? node58634 : node58619;
													assign node58619 = (inp[5]) ? node58627 : node58620;
														assign node58620 = (inp[4]) ? node58624 : node58621;
															assign node58621 = (inp[9]) ? 4'b1110 : 4'b1010;
															assign node58624 = (inp[9]) ? 4'b1010 : 4'b1110;
														assign node58627 = (inp[4]) ? node58631 : node58628;
															assign node58628 = (inp[10]) ? 4'b1100 : 4'b1010;
															assign node58631 = (inp[9]) ? 4'b1000 : 4'b1100;
													assign node58634 = (inp[9]) ? node58640 : node58635;
														assign node58635 = (inp[4]) ? 4'b1100 : node58636;
															assign node58636 = (inp[5]) ? 4'b1000 : 4'b1010;
														assign node58640 = (inp[4]) ? 4'b1000 : 4'b1100;
								assign node58643 = (inp[5]) ? node58889 : node58644;
									assign node58644 = (inp[9]) ? node58756 : node58645;
										assign node58645 = (inp[4]) ? node58701 : node58646;
											assign node58646 = (inp[10]) ? node58678 : node58647;
												assign node58647 = (inp[12]) ? node58661 : node58648;
													assign node58648 = (inp[14]) ? node58654 : node58649;
														assign node58649 = (inp[0]) ? node58651 : 4'b1110;
															assign node58651 = (inp[15]) ? 4'b1110 : 4'b1100;
														assign node58654 = (inp[15]) ? node58658 : node58655;
															assign node58655 = (inp[0]) ? 4'b1100 : 4'b1110;
															assign node58658 = (inp[0]) ? 4'b1110 : 4'b1100;
													assign node58661 = (inp[3]) ? node58673 : node58662;
														assign node58662 = (inp[14]) ? node58668 : node58663;
															assign node58663 = (inp[0]) ? node58665 : 4'b1010;
																assign node58665 = (inp[15]) ? 4'b1010 : 4'b1000;
															assign node58668 = (inp[15]) ? 4'b1000 : node58669;
																assign node58669 = (inp[0]) ? 4'b1000 : 4'b1010;
														assign node58673 = (inp[0]) ? 4'b1010 : node58674;
															assign node58674 = (inp[15]) ? 4'b1000 : 4'b1010;
												assign node58678 = (inp[3]) ? node58694 : node58679;
													assign node58679 = (inp[14]) ? node58687 : node58680;
														assign node58680 = (inp[15]) ? node58684 : node58681;
															assign node58681 = (inp[0]) ? 4'b1000 : 4'b1010;
															assign node58684 = (inp[0]) ? 4'b1010 : 4'b1000;
														assign node58687 = (inp[0]) ? node58691 : node58688;
															assign node58688 = (inp[15]) ? 4'b1000 : 4'b1010;
															assign node58691 = (inp[15]) ? 4'b1010 : 4'b1000;
													assign node58694 = (inp[0]) ? node58698 : node58695;
														assign node58695 = (inp[15]) ? 4'b1000 : 4'b1010;
														assign node58698 = (inp[15]) ? 4'b1010 : 4'b1000;
											assign node58701 = (inp[12]) ? node58727 : node58702;
												assign node58702 = (inp[10]) ? node58718 : node58703;
													assign node58703 = (inp[14]) ? node58711 : node58704;
														assign node58704 = (inp[15]) ? node58708 : node58705;
															assign node58705 = (inp[0]) ? 4'b1000 : 4'b1010;
															assign node58708 = (inp[0]) ? 4'b1010 : 4'b1000;
														assign node58711 = (inp[15]) ? node58715 : node58712;
															assign node58712 = (inp[0]) ? 4'b1000 : 4'b1010;
															assign node58715 = (inp[0]) ? 4'b1010 : 4'b1000;
													assign node58718 = (inp[15]) ? 4'b1110 : node58719;
														assign node58719 = (inp[0]) ? node58723 : node58720;
															assign node58720 = (inp[3]) ? 4'b1100 : 4'b1110;
															assign node58723 = (inp[3]) ? 4'b1110 : 4'b1100;
												assign node58727 = (inp[14]) ? node58741 : node58728;
													assign node58728 = (inp[15]) ? node58730 : 4'b1110;
														assign node58730 = (inp[10]) ? node58736 : node58731;
															assign node58731 = (inp[3]) ? 4'b1110 : node58732;
																assign node58732 = (inp[0]) ? 4'b1110 : 4'b1100;
															assign node58736 = (inp[0]) ? node58738 : 4'b1110;
																assign node58738 = (inp[3]) ? 4'b1100 : 4'b1110;
													assign node58741 = (inp[15]) ? node58749 : node58742;
														assign node58742 = (inp[3]) ? node58746 : node58743;
															assign node58743 = (inp[0]) ? 4'b1100 : 4'b1110;
															assign node58746 = (inp[0]) ? 4'b1110 : 4'b1100;
														assign node58749 = (inp[0]) ? node58753 : node58750;
															assign node58750 = (inp[3]) ? 4'b1110 : 4'b1100;
															assign node58753 = (inp[3]) ? 4'b1100 : 4'b1110;
										assign node58756 = (inp[4]) ? node58828 : node58757;
											assign node58757 = (inp[10]) ? node58793 : node58758;
												assign node58758 = (inp[12]) ? node58774 : node58759;
													assign node58759 = (inp[3]) ? node58767 : node58760;
														assign node58760 = (inp[0]) ? node58764 : node58761;
															assign node58761 = (inp[15]) ? 4'b1000 : 4'b1010;
															assign node58764 = (inp[15]) ? 4'b1010 : 4'b1000;
														assign node58767 = (inp[0]) ? node58771 : node58768;
															assign node58768 = (inp[15]) ? 4'b1000 : 4'b1010;
															assign node58771 = (inp[15]) ? 4'b1010 : 4'b1000;
													assign node58774 = (inp[15]) ? node58788 : node58775;
														assign node58775 = (inp[14]) ? node58781 : node58776;
															assign node58776 = (inp[3]) ? 4'b1110 : node58777;
																assign node58777 = (inp[0]) ? 4'b1100 : 4'b1110;
															assign node58781 = (inp[0]) ? node58785 : node58782;
																assign node58782 = (inp[3]) ? 4'b1100 : 4'b1110;
																assign node58785 = (inp[3]) ? 4'b1110 : 4'b1100;
														assign node58788 = (inp[0]) ? 4'b1110 : node58789;
															assign node58789 = (inp[3]) ? 4'b1110 : 4'b1100;
												assign node58793 = (inp[14]) ? node58815 : node58794;
													assign node58794 = (inp[12]) ? node58808 : node58795;
														assign node58795 = (inp[0]) ? node58803 : node58796;
															assign node58796 = (inp[3]) ? node58800 : node58797;
																assign node58797 = (inp[15]) ? 4'b1100 : 4'b1110;
																assign node58800 = (inp[15]) ? 4'b1110 : 4'b1100;
															assign node58803 = (inp[15]) ? node58805 : 4'b1100;
																assign node58805 = (inp[3]) ? 4'b1100 : 4'b1110;
														assign node58808 = (inp[0]) ? 4'b1100 : node58809;
															assign node58809 = (inp[3]) ? node58811 : 4'b1100;
																assign node58811 = (inp[15]) ? 4'b1110 : 4'b1100;
													assign node58815 = (inp[3]) ? node58823 : node58816;
														assign node58816 = (inp[0]) ? node58820 : node58817;
															assign node58817 = (inp[15]) ? 4'b1100 : 4'b1110;
															assign node58820 = (inp[15]) ? 4'b1110 : 4'b1100;
														assign node58823 = (inp[0]) ? 4'b1110 : node58824;
															assign node58824 = (inp[15]) ? 4'b1110 : 4'b1100;
											assign node58828 = (inp[12]) ? node58856 : node58829;
												assign node58829 = (inp[10]) ? node58847 : node58830;
													assign node58830 = (inp[3]) ? node58840 : node58831;
														assign node58831 = (inp[14]) ? node58835 : node58832;
															assign node58832 = (inp[15]) ? 4'b1110 : 4'b1100;
															assign node58835 = (inp[0]) ? 4'b1100 : node58836;
																assign node58836 = (inp[15]) ? 4'b1100 : 4'b1110;
														assign node58840 = (inp[0]) ? node58844 : node58841;
															assign node58841 = (inp[15]) ? 4'b1110 : 4'b1100;
															assign node58844 = (inp[15]) ? 4'b1100 : 4'b1110;
													assign node58847 = (inp[0]) ? node58849 : 4'b1010;
														assign node58849 = (inp[3]) ? node58853 : node58850;
															assign node58850 = (inp[15]) ? 4'b1010 : 4'b1000;
															assign node58853 = (inp[15]) ? 4'b1000 : 4'b1010;
												assign node58856 = (inp[14]) ? node58876 : node58857;
													assign node58857 = (inp[3]) ? node58867 : node58858;
														assign node58858 = (inp[10]) ? node58860 : 4'b1010;
															assign node58860 = (inp[15]) ? node58864 : node58861;
																assign node58861 = (inp[0]) ? 4'b1000 : 4'b1010;
																assign node58864 = (inp[0]) ? 4'b1010 : 4'b1000;
														assign node58867 = (inp[10]) ? node58869 : 4'b1000;
															assign node58869 = (inp[15]) ? node58873 : node58870;
																assign node58870 = (inp[0]) ? 4'b1010 : 4'b1000;
																assign node58873 = (inp[0]) ? 4'b1000 : 4'b1010;
													assign node58876 = (inp[3]) ? node58884 : node58877;
														assign node58877 = (inp[0]) ? node58881 : node58878;
															assign node58878 = (inp[15]) ? 4'b1000 : 4'b1010;
															assign node58881 = (inp[15]) ? 4'b1010 : 4'b1000;
														assign node58884 = (inp[15]) ? node58886 : 4'b1010;
															assign node58886 = (inp[0]) ? 4'b1000 : 4'b1010;
									assign node58889 = (inp[14]) ? node59039 : node58890;
										assign node58890 = (inp[12]) ? node58982 : node58891;
											assign node58891 = (inp[9]) ? node58939 : node58892;
												assign node58892 = (inp[0]) ? node58920 : node58893;
													assign node58893 = (inp[15]) ? node58907 : node58894;
														assign node58894 = (inp[3]) ? node58900 : node58895;
															assign node58895 = (inp[10]) ? 4'b1100 : node58896;
																assign node58896 = (inp[4]) ? 4'b1010 : 4'b1110;
															assign node58900 = (inp[10]) ? node58904 : node58901;
																assign node58901 = (inp[4]) ? 4'b1000 : 4'b1100;
																assign node58904 = (inp[4]) ? 4'b1100 : 4'b1000;
														assign node58907 = (inp[3]) ? node58915 : node58908;
															assign node58908 = (inp[10]) ? node58912 : node58909;
																assign node58909 = (inp[4]) ? 4'b1000 : 4'b1100;
																assign node58912 = (inp[4]) ? 4'b1110 : 4'b1000;
															assign node58915 = (inp[10]) ? 4'b1110 : node58916;
																assign node58916 = (inp[4]) ? 4'b1010 : 4'b1110;
													assign node58920 = (inp[15]) ? node58930 : node58921;
														assign node58921 = (inp[3]) ? node58923 : 4'b1110;
															assign node58923 = (inp[4]) ? node58927 : node58924;
																assign node58924 = (inp[10]) ? 4'b1010 : 4'b1110;
																assign node58927 = (inp[10]) ? 4'b1110 : 4'b1010;
														assign node58930 = (inp[3]) ? node58934 : node58931;
															assign node58931 = (inp[10]) ? 4'b1010 : 4'b1110;
															assign node58934 = (inp[10]) ? 4'b1000 : node58935;
																assign node58935 = (inp[4]) ? 4'b1000 : 4'b1100;
												assign node58939 = (inp[10]) ? node58969 : node58940;
													assign node58940 = (inp[4]) ? node58954 : node58941;
														assign node58941 = (inp[3]) ? node58949 : node58942;
															assign node58942 = (inp[0]) ? node58946 : node58943;
																assign node58943 = (inp[15]) ? 4'b1000 : 4'b1010;
																assign node58946 = (inp[15]) ? 4'b1010 : 4'b1000;
															assign node58949 = (inp[0]) ? 4'b1000 : node58950;
																assign node58950 = (inp[15]) ? 4'b1010 : 4'b1000;
														assign node58954 = (inp[3]) ? node58962 : node58955;
															assign node58955 = (inp[0]) ? node58959 : node58956;
																assign node58956 = (inp[15]) ? 4'b1110 : 4'b1100;
																assign node58959 = (inp[15]) ? 4'b1100 : 4'b1110;
															assign node58962 = (inp[15]) ? node58966 : node58963;
																assign node58963 = (inp[0]) ? 4'b1110 : 4'b1100;
																assign node58966 = (inp[0]) ? 4'b1100 : 4'b1110;
													assign node58969 = (inp[4]) ? node58975 : node58970;
														assign node58970 = (inp[0]) ? 4'b1100 : node58971;
															assign node58971 = (inp[15]) ? 4'b1110 : 4'b1100;
														assign node58975 = (inp[15]) ? node58979 : node58976;
															assign node58976 = (inp[0]) ? 4'b1010 : 4'b1000;
															assign node58979 = (inp[0]) ? 4'b1000 : 4'b1010;
											assign node58982 = (inp[0]) ? node59002 : node58983;
												assign node58983 = (inp[15]) ? node58993 : node58984;
													assign node58984 = (inp[4]) ? node58990 : node58985;
														assign node58985 = (inp[9]) ? 4'b1100 : node58986;
															assign node58986 = (inp[3]) ? 4'b1000 : 4'b1010;
														assign node58990 = (inp[9]) ? 4'b1000 : 4'b1100;
													assign node58993 = (inp[9]) ? node58999 : node58994;
														assign node58994 = (inp[4]) ? 4'b1110 : node58995;
															assign node58995 = (inp[3]) ? 4'b1010 : 4'b1000;
														assign node58999 = (inp[4]) ? 4'b1010 : 4'b1110;
												assign node59002 = (inp[15]) ? node59018 : node59003;
													assign node59003 = (inp[3]) ? node59009 : node59004;
														assign node59004 = (inp[4]) ? node59006 : 4'b1000;
															assign node59006 = (inp[10]) ? 4'b1110 : 4'b1010;
														assign node59009 = (inp[10]) ? node59015 : node59010;
															assign node59010 = (inp[9]) ? 4'b1110 : node59011;
																assign node59011 = (inp[4]) ? 4'b1110 : 4'b1010;
															assign node59015 = (inp[4]) ? 4'b1010 : 4'b1110;
													assign node59018 = (inp[3]) ? node59026 : node59019;
														assign node59019 = (inp[9]) ? node59023 : node59020;
															assign node59020 = (inp[4]) ? 4'b1100 : 4'b1010;
															assign node59023 = (inp[4]) ? 4'b1000 : 4'b1100;
														assign node59026 = (inp[10]) ? node59034 : node59027;
															assign node59027 = (inp[9]) ? node59031 : node59028;
																assign node59028 = (inp[4]) ? 4'b1100 : 4'b1000;
																assign node59031 = (inp[4]) ? 4'b1000 : 4'b1100;
															assign node59034 = (inp[4]) ? node59036 : 4'b1000;
																assign node59036 = (inp[9]) ? 4'b1000 : 4'b1100;
										assign node59039 = (inp[0]) ? node59111 : node59040;
											assign node59040 = (inp[15]) ? node59082 : node59041;
												assign node59041 = (inp[3]) ? node59057 : node59042;
													assign node59042 = (inp[4]) ? node59048 : node59043;
														assign node59043 = (inp[9]) ? node59045 : 4'b1010;
															assign node59045 = (inp[12]) ? 4'b1100 : 4'b1010;
														assign node59048 = (inp[9]) ? node59054 : node59049;
															assign node59049 = (inp[12]) ? 4'b1100 : node59050;
																assign node59050 = (inp[10]) ? 4'b1100 : 4'b1010;
															assign node59054 = (inp[10]) ? 4'b1000 : 4'b1100;
													assign node59057 = (inp[12]) ? node59073 : node59058;
														assign node59058 = (inp[9]) ? node59066 : node59059;
															assign node59059 = (inp[4]) ? node59063 : node59060;
																assign node59060 = (inp[10]) ? 4'b1000 : 4'b1100;
																assign node59063 = (inp[10]) ? 4'b1100 : 4'b1000;
															assign node59066 = (inp[4]) ? node59070 : node59067;
																assign node59067 = (inp[10]) ? 4'b1100 : 4'b1000;
																assign node59070 = (inp[10]) ? 4'b1000 : 4'b1100;
														assign node59073 = (inp[10]) ? node59079 : node59074;
															assign node59074 = (inp[4]) ? 4'b1100 : node59075;
																assign node59075 = (inp[9]) ? 4'b1100 : 4'b1000;
															assign node59079 = (inp[4]) ? 4'b1000 : 4'b1100;
												assign node59082 = (inp[3]) ? node59100 : node59083;
													assign node59083 = (inp[9]) ? node59093 : node59084;
														assign node59084 = (inp[12]) ? node59090 : node59085;
															assign node59085 = (inp[10]) ? 4'b1000 : node59086;
																assign node59086 = (inp[4]) ? 4'b1000 : 4'b1100;
															assign node59090 = (inp[4]) ? 4'b1110 : 4'b1000;
														assign node59093 = (inp[4]) ? node59095 : 4'b1110;
															assign node59095 = (inp[12]) ? 4'b1010 : node59096;
																assign node59096 = (inp[10]) ? 4'b1010 : 4'b1110;
													assign node59100 = (inp[4]) ? node59102 : 4'b1110;
														assign node59102 = (inp[9]) ? node59108 : node59103;
															assign node59103 = (inp[10]) ? 4'b1110 : node59104;
																assign node59104 = (inp[12]) ? 4'b1110 : 4'b1010;
															assign node59108 = (inp[10]) ? 4'b1010 : 4'b1110;
											assign node59111 = (inp[15]) ? node59155 : node59112;
												assign node59112 = (inp[3]) ? node59132 : node59113;
													assign node59113 = (inp[4]) ? node59123 : node59114;
														assign node59114 = (inp[9]) ? node59118 : node59115;
															assign node59115 = (inp[12]) ? 4'b1000 : 4'b1100;
															assign node59118 = (inp[10]) ? 4'b1110 : node59119;
																assign node59119 = (inp[12]) ? 4'b1110 : 4'b1000;
														assign node59123 = (inp[10]) ? 4'b1110 : node59124;
															assign node59124 = (inp[9]) ? node59128 : node59125;
																assign node59125 = (inp[12]) ? 4'b1110 : 4'b1000;
																assign node59128 = (inp[12]) ? 4'b1010 : 4'b1110;
													assign node59132 = (inp[10]) ? node59148 : node59133;
														assign node59133 = (inp[4]) ? node59141 : node59134;
															assign node59134 = (inp[12]) ? node59138 : node59135;
																assign node59135 = (inp[9]) ? 4'b1010 : 4'b1110;
																assign node59138 = (inp[9]) ? 4'b1110 : 4'b1010;
															assign node59141 = (inp[12]) ? node59145 : node59142;
																assign node59142 = (inp[9]) ? 4'b1110 : 4'b1010;
																assign node59145 = (inp[9]) ? 4'b1010 : 4'b1110;
														assign node59148 = (inp[4]) ? node59152 : node59149;
															assign node59149 = (inp[9]) ? 4'b1110 : 4'b1010;
															assign node59152 = (inp[9]) ? 4'b1010 : 4'b1110;
												assign node59155 = (inp[9]) ? node59167 : node59156;
													assign node59156 = (inp[4]) ? node59162 : node59157;
														assign node59157 = (inp[12]) ? 4'b1010 : node59158;
															assign node59158 = (inp[10]) ? 4'b1010 : 4'b1110;
														assign node59162 = (inp[10]) ? 4'b1100 : node59163;
															assign node59163 = (inp[3]) ? 4'b1000 : 4'b1010;
													assign node59167 = (inp[4]) ? node59173 : node59168;
														assign node59168 = (inp[10]) ? 4'b1100 : node59169;
															assign node59169 = (inp[12]) ? 4'b1100 : 4'b1010;
														assign node59173 = (inp[12]) ? 4'b1000 : node59174;
															assign node59174 = (inp[10]) ? 4'b1000 : 4'b1100;
							assign node59178 = (inp[2]) ? node59700 : node59179;
								assign node59179 = (inp[14]) ? node59455 : node59180;
									assign node59180 = (inp[15]) ? node59306 : node59181;
										assign node59181 = (inp[0]) ? node59255 : node59182;
											assign node59182 = (inp[3]) ? node59218 : node59183;
												assign node59183 = (inp[5]) ? node59199 : node59184;
													assign node59184 = (inp[4]) ? node59194 : node59185;
														assign node59185 = (inp[12]) ? 4'b1110 : node59186;
															assign node59186 = (inp[10]) ? node59190 : node59187;
																assign node59187 = (inp[9]) ? 4'b1010 : 4'b1110;
																assign node59190 = (inp[9]) ? 4'b1110 : 4'b1010;
														assign node59194 = (inp[9]) ? 4'b1010 : node59195;
															assign node59195 = (inp[10]) ? 4'b1110 : 4'b1010;
													assign node59199 = (inp[4]) ? node59209 : node59200;
														assign node59200 = (inp[10]) ? node59206 : node59201;
															assign node59201 = (inp[9]) ? 4'b1010 : node59202;
																assign node59202 = (inp[12]) ? 4'b1010 : 4'b1110;
															assign node59206 = (inp[9]) ? 4'b1100 : 4'b1010;
														assign node59209 = (inp[9]) ? node59213 : node59210;
															assign node59210 = (inp[12]) ? 4'b1100 : 4'b1010;
															assign node59213 = (inp[10]) ? 4'b1000 : node59214;
																assign node59214 = (inp[12]) ? 4'b1000 : 4'b1100;
												assign node59218 = (inp[5]) ? node59234 : node59219;
													assign node59219 = (inp[9]) ? node59227 : node59220;
														assign node59220 = (inp[4]) ? node59224 : node59221;
															assign node59221 = (inp[10]) ? 4'b1010 : 4'b1110;
															assign node59224 = (inp[10]) ? 4'b1100 : 4'b1010;
														assign node59227 = (inp[4]) ? node59231 : node59228;
															assign node59228 = (inp[12]) ? 4'b1100 : 4'b1010;
															assign node59231 = (inp[10]) ? 4'b1000 : 4'b1100;
													assign node59234 = (inp[12]) ? node59250 : node59235;
														assign node59235 = (inp[4]) ? node59243 : node59236;
															assign node59236 = (inp[9]) ? node59240 : node59237;
																assign node59237 = (inp[10]) ? 4'b1000 : 4'b1100;
																assign node59240 = (inp[10]) ? 4'b1100 : 4'b1000;
															assign node59243 = (inp[10]) ? node59247 : node59244;
																assign node59244 = (inp[9]) ? 4'b1100 : 4'b1000;
																assign node59247 = (inp[9]) ? 4'b1000 : 4'b1100;
														assign node59250 = (inp[9]) ? node59252 : 4'b1100;
															assign node59252 = (inp[4]) ? 4'b1000 : 4'b1100;
											assign node59255 = (inp[5]) ? node59285 : node59256;
												assign node59256 = (inp[3]) ? node59274 : node59257;
													assign node59257 = (inp[12]) ? node59267 : node59258;
														assign node59258 = (inp[4]) ? node59260 : 4'b1100;
															assign node59260 = (inp[10]) ? node59264 : node59261;
																assign node59261 = (inp[9]) ? 4'b1100 : 4'b1000;
																assign node59264 = (inp[9]) ? 4'b1000 : 4'b1100;
														assign node59267 = (inp[9]) ? node59271 : node59268;
															assign node59268 = (inp[4]) ? 4'b1100 : 4'b1000;
															assign node59271 = (inp[4]) ? 4'b1000 : 4'b1100;
													assign node59274 = (inp[9]) ? node59280 : node59275;
														assign node59275 = (inp[4]) ? 4'b1110 : node59276;
															assign node59276 = (inp[10]) ? 4'b1000 : 4'b1100;
														assign node59280 = (inp[4]) ? node59282 : 4'b1110;
															assign node59282 = (inp[12]) ? 4'b1010 : 4'b1110;
												assign node59285 = (inp[4]) ? node59299 : node59286;
													assign node59286 = (inp[9]) ? node59292 : node59287;
														assign node59287 = (inp[3]) ? node59289 : 4'b1000;
															assign node59289 = (inp[12]) ? 4'b1010 : 4'b1110;
														assign node59292 = (inp[12]) ? 4'b1110 : node59293;
															assign node59293 = (inp[10]) ? 4'b1110 : node59294;
																assign node59294 = (inp[3]) ? 4'b1010 : 4'b1000;
													assign node59299 = (inp[9]) ? node59301 : 4'b1110;
														assign node59301 = (inp[12]) ? 4'b1010 : node59302;
															assign node59302 = (inp[10]) ? 4'b1010 : 4'b1110;
										assign node59306 = (inp[10]) ? node59384 : node59307;
											assign node59307 = (inp[0]) ? node59345 : node59308;
												assign node59308 = (inp[3]) ? node59332 : node59309;
													assign node59309 = (inp[5]) ? node59319 : node59310;
														assign node59310 = (inp[4]) ? 4'b1100 : node59311;
															assign node59311 = (inp[9]) ? node59315 : node59312;
																assign node59312 = (inp[12]) ? 4'b1000 : 4'b1100;
																assign node59315 = (inp[12]) ? 4'b1100 : 4'b1000;
														assign node59319 = (inp[4]) ? node59325 : node59320;
															assign node59320 = (inp[12]) ? node59322 : 4'b1000;
																assign node59322 = (inp[9]) ? 4'b1110 : 4'b1000;
															assign node59325 = (inp[12]) ? node59329 : node59326;
																assign node59326 = (inp[9]) ? 4'b1110 : 4'b1000;
																assign node59329 = (inp[9]) ? 4'b1010 : 4'b1110;
													assign node59332 = (inp[9]) ? node59338 : node59333;
														assign node59333 = (inp[5]) ? node59335 : 4'b1000;
															assign node59335 = (inp[12]) ? 4'b1110 : 4'b1010;
														assign node59338 = (inp[4]) ? node59342 : node59339;
															assign node59339 = (inp[12]) ? 4'b1110 : 4'b1010;
															assign node59342 = (inp[12]) ? 4'b1010 : 4'b1110;
												assign node59345 = (inp[5]) ? node59373 : node59346;
													assign node59346 = (inp[3]) ? node59360 : node59347;
														assign node59347 = (inp[12]) ? node59353 : node59348;
															assign node59348 = (inp[4]) ? 4'b1010 : node59349;
																assign node59349 = (inp[9]) ? 4'b1010 : 4'b1110;
															assign node59353 = (inp[9]) ? node59357 : node59354;
																assign node59354 = (inp[4]) ? 4'b1110 : 4'b1010;
																assign node59357 = (inp[4]) ? 4'b1010 : 4'b1110;
														assign node59360 = (inp[12]) ? node59366 : node59361;
															assign node59361 = (inp[4]) ? 4'b1010 : node59362;
																assign node59362 = (inp[9]) ? 4'b1010 : 4'b1110;
															assign node59366 = (inp[4]) ? node59370 : node59367;
																assign node59367 = (inp[9]) ? 4'b1100 : 4'b1010;
																assign node59370 = (inp[9]) ? 4'b1000 : 4'b1100;
													assign node59373 = (inp[4]) ? node59377 : node59374;
														assign node59374 = (inp[3]) ? 4'b1000 : 4'b1010;
														assign node59377 = (inp[12]) ? node59381 : node59378;
															assign node59378 = (inp[9]) ? 4'b1100 : 4'b1010;
															assign node59381 = (inp[9]) ? 4'b1000 : 4'b1100;
											assign node59384 = (inp[12]) ? node59418 : node59385;
												assign node59385 = (inp[9]) ? node59401 : node59386;
													assign node59386 = (inp[4]) ? node59392 : node59387;
														assign node59387 = (inp[5]) ? 4'b1000 : node59388;
															assign node59388 = (inp[0]) ? 4'b1010 : 4'b1000;
														assign node59392 = (inp[5]) ? 4'b1100 : node59393;
															assign node59393 = (inp[0]) ? node59397 : node59394;
																assign node59394 = (inp[3]) ? 4'b1110 : 4'b1100;
																assign node59397 = (inp[3]) ? 4'b1100 : 4'b1110;
													assign node59401 = (inp[4]) ? node59409 : node59402;
														assign node59402 = (inp[0]) ? node59406 : node59403;
															assign node59403 = (inp[5]) ? 4'b1110 : 4'b1100;
															assign node59406 = (inp[3]) ? 4'b1100 : 4'b1110;
														assign node59409 = (inp[5]) ? 4'b1010 : node59410;
															assign node59410 = (inp[3]) ? node59414 : node59411;
																assign node59411 = (inp[0]) ? 4'b1010 : 4'b1000;
																assign node59414 = (inp[0]) ? 4'b1000 : 4'b1010;
												assign node59418 = (inp[5]) ? node59434 : node59419;
													assign node59419 = (inp[0]) ? node59429 : node59420;
														assign node59420 = (inp[3]) ? node59422 : 4'b1100;
															assign node59422 = (inp[4]) ? node59426 : node59423;
																assign node59423 = (inp[9]) ? 4'b1110 : 4'b1000;
																assign node59426 = (inp[9]) ? 4'b1010 : 4'b1110;
														assign node59429 = (inp[4]) ? node59431 : 4'b1010;
															assign node59431 = (inp[9]) ? 4'b1010 : 4'b1110;
													assign node59434 = (inp[0]) ? node59448 : node59435;
														assign node59435 = (inp[3]) ? node59441 : node59436;
															assign node59436 = (inp[9]) ? node59438 : 4'b1000;
																assign node59438 = (inp[4]) ? 4'b1010 : 4'b1110;
															assign node59441 = (inp[4]) ? node59445 : node59442;
																assign node59442 = (inp[9]) ? 4'b1110 : 4'b1010;
																assign node59445 = (inp[9]) ? 4'b1010 : 4'b1110;
														assign node59448 = (inp[3]) ? 4'b1100 : node59449;
															assign node59449 = (inp[4]) ? 4'b1100 : node59450;
																assign node59450 = (inp[9]) ? 4'b1100 : 4'b1010;
									assign node59455 = (inp[9]) ? node59569 : node59456;
										assign node59456 = (inp[4]) ? node59520 : node59457;
											assign node59457 = (inp[10]) ? node59497 : node59458;
												assign node59458 = (inp[12]) ? node59480 : node59459;
													assign node59459 = (inp[5]) ? node59471 : node59460;
														assign node59460 = (inp[3]) ? node59466 : node59461;
															assign node59461 = (inp[0]) ? node59463 : 4'b0111;
																assign node59463 = (inp[15]) ? 4'b0111 : 4'b0101;
															assign node59466 = (inp[0]) ? 4'b0101 : node59467;
																assign node59467 = (inp[15]) ? 4'b0101 : 4'b0111;
														assign node59471 = (inp[0]) ? 4'b0111 : node59472;
															assign node59472 = (inp[3]) ? node59476 : node59473;
																assign node59473 = (inp[15]) ? 4'b0101 : 4'b0111;
																assign node59476 = (inp[15]) ? 4'b0111 : 4'b0101;
													assign node59480 = (inp[5]) ? node59488 : node59481;
														assign node59481 = (inp[0]) ? node59485 : node59482;
															assign node59482 = (inp[15]) ? 4'b0001 : 4'b0011;
															assign node59485 = (inp[15]) ? 4'b0011 : 4'b0001;
														assign node59488 = (inp[15]) ? node59490 : 4'b0001;
															assign node59490 = (inp[0]) ? node59494 : node59491;
																assign node59491 = (inp[3]) ? 4'b0011 : 4'b0001;
																assign node59494 = (inp[3]) ? 4'b0001 : 4'b0011;
												assign node59497 = (inp[0]) ? node59509 : node59498;
													assign node59498 = (inp[5]) ? node59502 : node59499;
														assign node59499 = (inp[15]) ? 4'b0001 : 4'b0011;
														assign node59502 = (inp[15]) ? node59506 : node59503;
															assign node59503 = (inp[3]) ? 4'b0001 : 4'b0011;
															assign node59506 = (inp[3]) ? 4'b0011 : 4'b0001;
													assign node59509 = (inp[15]) ? node59515 : node59510;
														assign node59510 = (inp[3]) ? node59512 : 4'b0001;
															assign node59512 = (inp[5]) ? 4'b0011 : 4'b0001;
														assign node59515 = (inp[3]) ? node59517 : 4'b0011;
															assign node59517 = (inp[5]) ? 4'b0001 : 4'b0011;
											assign node59520 = (inp[10]) ? node59552 : node59521;
												assign node59521 = (inp[12]) ? node59537 : node59522;
													assign node59522 = (inp[15]) ? node59528 : node59523;
														assign node59523 = (inp[5]) ? 4'b0001 : node59524;
															assign node59524 = (inp[0]) ? 4'b0001 : 4'b0011;
														assign node59528 = (inp[0]) ? node59532 : node59529;
															assign node59529 = (inp[5]) ? 4'b0011 : 4'b0001;
															assign node59532 = (inp[5]) ? node59534 : 4'b0011;
																assign node59534 = (inp[3]) ? 4'b0001 : 4'b0011;
													assign node59537 = (inp[0]) ? node59547 : node59538;
														assign node59538 = (inp[5]) ? 4'b0111 : node59539;
															assign node59539 = (inp[15]) ? node59543 : node59540;
																assign node59540 = (inp[3]) ? 4'b0101 : 4'b0111;
																assign node59543 = (inp[3]) ? 4'b0111 : 4'b0101;
														assign node59547 = (inp[15]) ? node59549 : 4'b0101;
															assign node59549 = (inp[5]) ? 4'b0101 : 4'b0111;
												assign node59552 = (inp[3]) ? node59562 : node59553;
													assign node59553 = (inp[0]) ? node59555 : 4'b0101;
														assign node59555 = (inp[15]) ? node59559 : node59556;
															assign node59556 = (inp[5]) ? 4'b0111 : 4'b0101;
															assign node59559 = (inp[5]) ? 4'b0101 : 4'b0111;
													assign node59562 = (inp[15]) ? node59566 : node59563;
														assign node59563 = (inp[0]) ? 4'b0111 : 4'b0101;
														assign node59566 = (inp[0]) ? 4'b0101 : 4'b0111;
										assign node59569 = (inp[4]) ? node59637 : node59570;
											assign node59570 = (inp[12]) ? node59608 : node59571;
												assign node59571 = (inp[10]) ? node59593 : node59572;
													assign node59572 = (inp[15]) ? node59582 : node59573;
														assign node59573 = (inp[3]) ? node59575 : 4'b0001;
															assign node59575 = (inp[0]) ? node59579 : node59576;
																assign node59576 = (inp[5]) ? 4'b0001 : 4'b0011;
																assign node59579 = (inp[5]) ? 4'b0011 : 4'b0001;
														assign node59582 = (inp[0]) ? node59588 : node59583;
															assign node59583 = (inp[5]) ? node59585 : 4'b0001;
																assign node59585 = (inp[3]) ? 4'b0011 : 4'b0001;
															assign node59588 = (inp[5]) ? node59590 : 4'b0011;
																assign node59590 = (inp[3]) ? 4'b0001 : 4'b0011;
													assign node59593 = (inp[15]) ? node59597 : node59594;
														assign node59594 = (inp[0]) ? 4'b0111 : 4'b0101;
														assign node59597 = (inp[0]) ? node59603 : node59598;
															assign node59598 = (inp[5]) ? 4'b0111 : node59599;
																assign node59599 = (inp[3]) ? 4'b0111 : 4'b0101;
															assign node59603 = (inp[5]) ? 4'b0101 : node59604;
																assign node59604 = (inp[3]) ? 4'b0101 : 4'b0111;
												assign node59608 = (inp[5]) ? node59622 : node59609;
													assign node59609 = (inp[0]) ? node59615 : node59610;
														assign node59610 = (inp[15]) ? node59612 : 4'b0111;
															assign node59612 = (inp[3]) ? 4'b0111 : 4'b0101;
														assign node59615 = (inp[15]) ? node59619 : node59616;
															assign node59616 = (inp[3]) ? 4'b0111 : 4'b0101;
															assign node59619 = (inp[3]) ? 4'b0101 : 4'b0111;
													assign node59622 = (inp[3]) ? node59630 : node59623;
														assign node59623 = (inp[15]) ? node59627 : node59624;
															assign node59624 = (inp[0]) ? 4'b0111 : 4'b0101;
															assign node59627 = (inp[0]) ? 4'b0101 : 4'b0111;
														assign node59630 = (inp[0]) ? node59634 : node59631;
															assign node59631 = (inp[15]) ? 4'b0111 : 4'b0101;
															assign node59634 = (inp[15]) ? 4'b0101 : 4'b0111;
											assign node59637 = (inp[12]) ? node59671 : node59638;
												assign node59638 = (inp[10]) ? node59654 : node59639;
													assign node59639 = (inp[0]) ? node59645 : node59640;
														assign node59640 = (inp[5]) ? node59642 : 4'b0101;
															assign node59642 = (inp[3]) ? 4'b0111 : 4'b0101;
														assign node59645 = (inp[15]) ? node59651 : node59646;
															assign node59646 = (inp[5]) ? 4'b0111 : node59647;
																assign node59647 = (inp[3]) ? 4'b0111 : 4'b0101;
															assign node59651 = (inp[3]) ? 4'b0101 : 4'b0111;
													assign node59654 = (inp[3]) ? node59666 : node59655;
														assign node59655 = (inp[5]) ? node59661 : node59656;
															assign node59656 = (inp[0]) ? 4'b0001 : node59657;
																assign node59657 = (inp[15]) ? 4'b0001 : 4'b0011;
															assign node59661 = (inp[15]) ? 4'b0011 : node59662;
																assign node59662 = (inp[0]) ? 4'b0011 : 4'b0001;
														assign node59666 = (inp[15]) ? node59668 : 4'b0011;
															assign node59668 = (inp[0]) ? 4'b0001 : 4'b0011;
												assign node59671 = (inp[5]) ? node59685 : node59672;
													assign node59672 = (inp[15]) ? node59678 : node59673;
														assign node59673 = (inp[0]) ? 4'b0011 : node59674;
															assign node59674 = (inp[3]) ? 4'b0001 : 4'b0011;
														assign node59678 = (inp[3]) ? node59682 : node59679;
															assign node59679 = (inp[0]) ? 4'b0011 : 4'b0001;
															assign node59682 = (inp[0]) ? 4'b0001 : 4'b0011;
													assign node59685 = (inp[3]) ? node59695 : node59686;
														assign node59686 = (inp[10]) ? node59692 : node59687;
															assign node59687 = (inp[0]) ? node59689 : 4'b0011;
																assign node59689 = (inp[15]) ? 4'b0001 : 4'b0011;
															assign node59692 = (inp[15]) ? 4'b0011 : 4'b0001;
														assign node59695 = (inp[0]) ? node59697 : 4'b0001;
															assign node59697 = (inp[15]) ? 4'b0001 : 4'b0011;
								assign node59700 = (inp[3]) ? node59948 : node59701;
									assign node59701 = (inp[4]) ? node59803 : node59702;
										assign node59702 = (inp[9]) ? node59756 : node59703;
											assign node59703 = (inp[12]) ? node59733 : node59704;
												assign node59704 = (inp[10]) ? node59720 : node59705;
													assign node59705 = (inp[14]) ? node59713 : node59706;
														assign node59706 = (inp[0]) ? node59710 : node59707;
															assign node59707 = (inp[15]) ? 4'b0101 : 4'b0111;
															assign node59710 = (inp[15]) ? 4'b0111 : 4'b0101;
														assign node59713 = (inp[0]) ? node59717 : node59714;
															assign node59714 = (inp[15]) ? 4'b0101 : 4'b0111;
															assign node59717 = (inp[15]) ? 4'b0111 : 4'b0101;
													assign node59720 = (inp[5]) ? node59726 : node59721;
														assign node59721 = (inp[0]) ? node59723 : 4'b0001;
															assign node59723 = (inp[15]) ? 4'b0011 : 4'b0001;
														assign node59726 = (inp[0]) ? node59730 : node59727;
															assign node59727 = (inp[15]) ? 4'b0001 : 4'b0011;
															assign node59730 = (inp[15]) ? 4'b0011 : 4'b0001;
												assign node59733 = (inp[14]) ? node59751 : node59734;
													assign node59734 = (inp[5]) ? node59742 : node59735;
														assign node59735 = (inp[15]) ? node59739 : node59736;
															assign node59736 = (inp[0]) ? 4'b0001 : 4'b0011;
															assign node59739 = (inp[0]) ? 4'b0011 : 4'b0001;
														assign node59742 = (inp[10]) ? 4'b0001 : node59743;
															assign node59743 = (inp[0]) ? node59747 : node59744;
																assign node59744 = (inp[15]) ? 4'b0001 : 4'b0011;
																assign node59747 = (inp[15]) ? 4'b0011 : 4'b0001;
													assign node59751 = (inp[0]) ? 4'b0011 : node59752;
														assign node59752 = (inp[15]) ? 4'b0001 : 4'b0011;
											assign node59756 = (inp[12]) ? node59782 : node59757;
												assign node59757 = (inp[10]) ? node59767 : node59758;
													assign node59758 = (inp[14]) ? 4'b0011 : node59759;
														assign node59759 = (inp[15]) ? node59763 : node59760;
															assign node59760 = (inp[0]) ? 4'b0001 : 4'b0011;
															assign node59763 = (inp[0]) ? 4'b0011 : 4'b0001;
													assign node59767 = (inp[14]) ? node59769 : 4'b0111;
														assign node59769 = (inp[5]) ? node59777 : node59770;
															assign node59770 = (inp[15]) ? node59774 : node59771;
																assign node59771 = (inp[0]) ? 4'b0101 : 4'b0111;
																assign node59774 = (inp[0]) ? 4'b0111 : 4'b0101;
															assign node59777 = (inp[0]) ? node59779 : 4'b0111;
																assign node59779 = (inp[15]) ? 4'b0101 : 4'b0111;
												assign node59782 = (inp[0]) ? node59796 : node59783;
													assign node59783 = (inp[10]) ? node59791 : node59784;
														assign node59784 = (inp[15]) ? node59788 : node59785;
															assign node59785 = (inp[5]) ? 4'b0101 : 4'b0111;
															assign node59788 = (inp[5]) ? 4'b0111 : 4'b0101;
														assign node59791 = (inp[15]) ? node59793 : 4'b0111;
															assign node59793 = (inp[14]) ? 4'b0101 : 4'b0111;
													assign node59796 = (inp[15]) ? node59800 : node59797;
														assign node59797 = (inp[5]) ? 4'b0111 : 4'b0101;
														assign node59800 = (inp[5]) ? 4'b0101 : 4'b0111;
										assign node59803 = (inp[9]) ? node59859 : node59804;
											assign node59804 = (inp[10]) ? node59828 : node59805;
												assign node59805 = (inp[12]) ? node59813 : node59806;
													assign node59806 = (inp[15]) ? node59810 : node59807;
														assign node59807 = (inp[0]) ? 4'b0001 : 4'b0011;
														assign node59810 = (inp[0]) ? 4'b0011 : 4'b0001;
													assign node59813 = (inp[5]) ? node59819 : node59814;
														assign node59814 = (inp[14]) ? node59816 : 4'b0111;
															assign node59816 = (inp[15]) ? 4'b0101 : 4'b0111;
														assign node59819 = (inp[14]) ? node59823 : node59820;
															assign node59820 = (inp[0]) ? 4'b0111 : 4'b0101;
															assign node59823 = (inp[15]) ? node59825 : 4'b0101;
																assign node59825 = (inp[0]) ? 4'b0101 : 4'b0111;
												assign node59828 = (inp[12]) ? node59846 : node59829;
													assign node59829 = (inp[15]) ? node59839 : node59830;
														assign node59830 = (inp[14]) ? 4'b0111 : node59831;
															assign node59831 = (inp[5]) ? node59835 : node59832;
																assign node59832 = (inp[0]) ? 4'b0101 : 4'b0111;
																assign node59835 = (inp[0]) ? 4'b0111 : 4'b0101;
														assign node59839 = (inp[14]) ? node59841 : 4'b0111;
															assign node59841 = (inp[5]) ? node59843 : 4'b0101;
																assign node59843 = (inp[0]) ? 4'b0101 : 4'b0111;
													assign node59846 = (inp[0]) ? node59852 : node59847;
														assign node59847 = (inp[5]) ? 4'b0101 : node59848;
															assign node59848 = (inp[14]) ? 4'b0101 : 4'b0111;
														assign node59852 = (inp[5]) ? node59856 : node59853;
															assign node59853 = (inp[15]) ? 4'b0111 : 4'b0101;
															assign node59856 = (inp[15]) ? 4'b0101 : 4'b0111;
											assign node59859 = (inp[12]) ? node59905 : node59860;
												assign node59860 = (inp[10]) ? node59890 : node59861;
													assign node59861 = (inp[14]) ? node59877 : node59862;
														assign node59862 = (inp[15]) ? node59870 : node59863;
															assign node59863 = (inp[0]) ? node59867 : node59864;
																assign node59864 = (inp[5]) ? 4'b0101 : 4'b0111;
																assign node59867 = (inp[5]) ? 4'b0111 : 4'b0101;
															assign node59870 = (inp[5]) ? node59874 : node59871;
																assign node59871 = (inp[0]) ? 4'b0111 : 4'b0101;
																assign node59874 = (inp[0]) ? 4'b0101 : 4'b0111;
														assign node59877 = (inp[5]) ? node59885 : node59878;
															assign node59878 = (inp[0]) ? node59882 : node59879;
																assign node59879 = (inp[15]) ? 4'b0101 : 4'b0111;
																assign node59882 = (inp[15]) ? 4'b0111 : 4'b0101;
															assign node59885 = (inp[15]) ? 4'b0111 : node59886;
																assign node59886 = (inp[0]) ? 4'b0111 : 4'b0101;
													assign node59890 = (inp[15]) ? node59898 : node59891;
														assign node59891 = (inp[5]) ? node59895 : node59892;
															assign node59892 = (inp[0]) ? 4'b0001 : 4'b0011;
															assign node59895 = (inp[14]) ? 4'b0001 : 4'b0011;
														assign node59898 = (inp[5]) ? node59902 : node59899;
															assign node59899 = (inp[0]) ? 4'b0011 : 4'b0001;
															assign node59902 = (inp[0]) ? 4'b0001 : 4'b0011;
												assign node59905 = (inp[10]) ? node59933 : node59906;
													assign node59906 = (inp[0]) ? node59920 : node59907;
														assign node59907 = (inp[14]) ? node59913 : node59908;
															assign node59908 = (inp[15]) ? 4'b0001 : node59909;
																assign node59909 = (inp[5]) ? 4'b0001 : 4'b0011;
															assign node59913 = (inp[5]) ? node59917 : node59914;
																assign node59914 = (inp[15]) ? 4'b0001 : 4'b0011;
																assign node59917 = (inp[15]) ? 4'b0011 : 4'b0001;
														assign node59920 = (inp[14]) ? node59926 : node59921;
															assign node59921 = (inp[15]) ? 4'b0011 : node59922;
																assign node59922 = (inp[5]) ? 4'b0011 : 4'b0001;
															assign node59926 = (inp[15]) ? node59930 : node59927;
																assign node59927 = (inp[5]) ? 4'b0011 : 4'b0001;
																assign node59930 = (inp[5]) ? 4'b0001 : 4'b0011;
													assign node59933 = (inp[0]) ? node59941 : node59934;
														assign node59934 = (inp[15]) ? node59938 : node59935;
															assign node59935 = (inp[5]) ? 4'b0001 : 4'b0011;
															assign node59938 = (inp[5]) ? 4'b0011 : 4'b0001;
														assign node59941 = (inp[15]) ? node59945 : node59942;
															assign node59942 = (inp[5]) ? 4'b0011 : 4'b0001;
															assign node59945 = (inp[5]) ? 4'b0001 : 4'b0011;
									assign node59948 = (inp[15]) ? node60054 : node59949;
										assign node59949 = (inp[0]) ? node60009 : node59950;
											assign node59950 = (inp[5]) ? node59974 : node59951;
												assign node59951 = (inp[9]) ? node59963 : node59952;
													assign node59952 = (inp[4]) ? node59958 : node59953;
														assign node59953 = (inp[10]) ? 4'b0011 : node59954;
															assign node59954 = (inp[12]) ? 4'b0011 : 4'b0111;
														assign node59958 = (inp[12]) ? 4'b0101 : node59959;
															assign node59959 = (inp[10]) ? 4'b0101 : 4'b0011;
													assign node59963 = (inp[4]) ? node59969 : node59964;
														assign node59964 = (inp[12]) ? 4'b0101 : node59965;
															assign node59965 = (inp[10]) ? 4'b0101 : 4'b0011;
														assign node59969 = (inp[10]) ? 4'b0001 : node59970;
															assign node59970 = (inp[12]) ? 4'b0001 : 4'b0101;
												assign node59974 = (inp[14]) ? node59994 : node59975;
													assign node59975 = (inp[9]) ? node59985 : node59976;
														assign node59976 = (inp[10]) ? 4'b0001 : node59977;
															assign node59977 = (inp[4]) ? node59981 : node59978;
																assign node59978 = (inp[12]) ? 4'b0001 : 4'b0101;
																assign node59981 = (inp[12]) ? 4'b0101 : 4'b0001;
														assign node59985 = (inp[4]) ? node59991 : node59986;
															assign node59986 = (inp[10]) ? 4'b0101 : node59987;
																assign node59987 = (inp[12]) ? 4'b0101 : 4'b0001;
															assign node59991 = (inp[12]) ? 4'b0001 : 4'b0101;
													assign node59994 = (inp[9]) ? node60004 : node59995;
														assign node59995 = (inp[4]) ? node59999 : node59996;
															assign node59996 = (inp[12]) ? 4'b0001 : 4'b0101;
															assign node59999 = (inp[12]) ? 4'b0101 : node60000;
																assign node60000 = (inp[10]) ? 4'b0101 : 4'b0001;
														assign node60004 = (inp[4]) ? node60006 : 4'b0101;
															assign node60006 = (inp[10]) ? 4'b0001 : 4'b0101;
											assign node60009 = (inp[5]) ? node60029 : node60010;
												assign node60010 = (inp[9]) ? node60018 : node60011;
													assign node60011 = (inp[4]) ? node60013 : 4'b0001;
														assign node60013 = (inp[10]) ? 4'b0111 : node60014;
															assign node60014 = (inp[12]) ? 4'b0111 : 4'b0001;
													assign node60018 = (inp[4]) ? node60024 : node60019;
														assign node60019 = (inp[10]) ? 4'b0111 : node60020;
															assign node60020 = (inp[12]) ? 4'b0111 : 4'b0001;
														assign node60024 = (inp[10]) ? 4'b0011 : node60025;
															assign node60025 = (inp[12]) ? 4'b0011 : 4'b0111;
												assign node60029 = (inp[12]) ? node60047 : node60030;
													assign node60030 = (inp[10]) ? node60038 : node60031;
														assign node60031 = (inp[9]) ? node60035 : node60032;
															assign node60032 = (inp[4]) ? 4'b0011 : 4'b0111;
															assign node60035 = (inp[4]) ? 4'b0111 : 4'b0011;
														assign node60038 = (inp[14]) ? node60044 : node60039;
															assign node60039 = (inp[4]) ? 4'b0111 : node60040;
																assign node60040 = (inp[9]) ? 4'b0111 : 4'b0011;
															assign node60044 = (inp[9]) ? 4'b0011 : 4'b0111;
													assign node60047 = (inp[4]) ? node60051 : node60048;
														assign node60048 = (inp[9]) ? 4'b0111 : 4'b0011;
														assign node60051 = (inp[9]) ? 4'b0011 : 4'b0111;
										assign node60054 = (inp[0]) ? node60100 : node60055;
											assign node60055 = (inp[5]) ? node60079 : node60056;
												assign node60056 = (inp[9]) ? node60068 : node60057;
													assign node60057 = (inp[4]) ? node60063 : node60058;
														assign node60058 = (inp[12]) ? 4'b0001 : node60059;
															assign node60059 = (inp[10]) ? 4'b0001 : 4'b0101;
														assign node60063 = (inp[12]) ? 4'b0111 : node60064;
															assign node60064 = (inp[10]) ? 4'b0111 : 4'b0001;
													assign node60068 = (inp[4]) ? node60074 : node60069;
														assign node60069 = (inp[10]) ? 4'b0111 : node60070;
															assign node60070 = (inp[12]) ? 4'b0111 : 4'b0001;
														assign node60074 = (inp[12]) ? 4'b0011 : node60075;
															assign node60075 = (inp[10]) ? 4'b0011 : 4'b0111;
												assign node60079 = (inp[10]) ? node60093 : node60080;
													assign node60080 = (inp[4]) ? node60088 : node60081;
														assign node60081 = (inp[9]) ? node60085 : node60082;
															assign node60082 = (inp[12]) ? 4'b0011 : 4'b0111;
															assign node60085 = (inp[12]) ? 4'b0111 : 4'b0011;
														assign node60088 = (inp[9]) ? node60090 : 4'b0111;
															assign node60090 = (inp[12]) ? 4'b0011 : 4'b0111;
													assign node60093 = (inp[9]) ? node60097 : node60094;
														assign node60094 = (inp[4]) ? 4'b0111 : 4'b0011;
														assign node60097 = (inp[4]) ? 4'b0011 : 4'b0111;
											assign node60100 = (inp[5]) ? node60122 : node60101;
												assign node60101 = (inp[9]) ? node60111 : node60102;
													assign node60102 = (inp[4]) ? node60106 : node60103;
														assign node60103 = (inp[12]) ? 4'b0011 : 4'b0111;
														assign node60106 = (inp[10]) ? 4'b0101 : node60107;
															assign node60107 = (inp[12]) ? 4'b0101 : 4'b0011;
													assign node60111 = (inp[4]) ? node60117 : node60112;
														assign node60112 = (inp[10]) ? 4'b0101 : node60113;
															assign node60113 = (inp[12]) ? 4'b0101 : 4'b0011;
														assign node60117 = (inp[10]) ? 4'b0001 : node60118;
															assign node60118 = (inp[12]) ? 4'b0001 : 4'b0101;
												assign node60122 = (inp[9]) ? node60134 : node60123;
													assign node60123 = (inp[4]) ? node60129 : node60124;
														assign node60124 = (inp[10]) ? 4'b0001 : node60125;
															assign node60125 = (inp[12]) ? 4'b0001 : 4'b0101;
														assign node60129 = (inp[12]) ? 4'b0101 : node60130;
															assign node60130 = (inp[10]) ? 4'b0101 : 4'b0001;
													assign node60134 = (inp[4]) ? node60138 : node60135;
														assign node60135 = (inp[10]) ? 4'b0101 : 4'b0001;
														assign node60138 = (inp[10]) ? 4'b0001 : node60139;
															assign node60139 = (inp[12]) ? 4'b0001 : 4'b0101;
						assign node60143 = (inp[7]) ? node61113 : node60144;
							assign node60144 = (inp[14]) ? node60690 : node60145;
								assign node60145 = (inp[2]) ? node60447 : node60146;
									assign node60146 = (inp[0]) ? node60304 : node60147;
										assign node60147 = (inp[15]) ? node60221 : node60148;
											assign node60148 = (inp[3]) ? node60184 : node60149;
												assign node60149 = (inp[5]) ? node60167 : node60150;
													assign node60150 = (inp[9]) ? node60160 : node60151;
														assign node60151 = (inp[4]) ? node60155 : node60152;
															assign node60152 = (inp[10]) ? 4'b1010 : 4'b1110;
															assign node60155 = (inp[10]) ? 4'b1110 : node60156;
																assign node60156 = (inp[12]) ? 4'b1110 : 4'b1010;
														assign node60160 = (inp[4]) ? node60162 : 4'b1110;
															assign node60162 = (inp[10]) ? 4'b1010 : node60163;
																assign node60163 = (inp[12]) ? 4'b1010 : 4'b1110;
													assign node60167 = (inp[10]) ? node60179 : node60168;
														assign node60168 = (inp[4]) ? node60174 : node60169;
															assign node60169 = (inp[9]) ? 4'b1010 : node60170;
																assign node60170 = (inp[12]) ? 4'b1010 : 4'b1110;
															assign node60174 = (inp[12]) ? 4'b1100 : node60175;
																assign node60175 = (inp[9]) ? 4'b1100 : 4'b1010;
														assign node60179 = (inp[9]) ? node60181 : 4'b1100;
															assign node60181 = (inp[4]) ? 4'b1000 : 4'b1100;
												assign node60184 = (inp[5]) ? node60204 : node60185;
													assign node60185 = (inp[9]) ? node60193 : node60186;
														assign node60186 = (inp[4]) ? 4'b1100 : node60187;
															assign node60187 = (inp[10]) ? 4'b1010 : node60188;
																assign node60188 = (inp[12]) ? 4'b1010 : 4'b1110;
														assign node60193 = (inp[4]) ? node60199 : node60194;
															assign node60194 = (inp[12]) ? 4'b1100 : node60195;
																assign node60195 = (inp[10]) ? 4'b1100 : 4'b1010;
															assign node60199 = (inp[10]) ? 4'b1000 : node60200;
																assign node60200 = (inp[12]) ? 4'b1000 : 4'b1100;
													assign node60204 = (inp[4]) ? node60212 : node60205;
														assign node60205 = (inp[9]) ? 4'b1100 : node60206;
															assign node60206 = (inp[10]) ? 4'b1000 : node60207;
																assign node60207 = (inp[12]) ? 4'b1000 : 4'b1100;
														assign node60212 = (inp[9]) ? node60216 : node60213;
															assign node60213 = (inp[10]) ? 4'b1100 : 4'b1000;
															assign node60216 = (inp[12]) ? 4'b1000 : node60217;
																assign node60217 = (inp[10]) ? 4'b1000 : 4'b1100;
											assign node60221 = (inp[3]) ? node60263 : node60222;
												assign node60222 = (inp[5]) ? node60248 : node60223;
													assign node60223 = (inp[12]) ? node60237 : node60224;
														assign node60224 = (inp[10]) ? node60230 : node60225;
															assign node60225 = (inp[4]) ? node60227 : 4'b1000;
																assign node60227 = (inp[9]) ? 4'b1100 : 4'b1000;
															assign node60230 = (inp[9]) ? node60234 : node60231;
																assign node60231 = (inp[4]) ? 4'b1100 : 4'b1000;
																assign node60234 = (inp[4]) ? 4'b1000 : 4'b1100;
														assign node60237 = (inp[10]) ? node60243 : node60238;
															assign node60238 = (inp[9]) ? node60240 : 4'b1100;
																assign node60240 = (inp[4]) ? 4'b1000 : 4'b1100;
															assign node60243 = (inp[4]) ? 4'b1100 : node60244;
																assign node60244 = (inp[9]) ? 4'b1100 : 4'b1000;
													assign node60248 = (inp[4]) ? node60258 : node60249;
														assign node60249 = (inp[9]) ? node60255 : node60250;
															assign node60250 = (inp[10]) ? 4'b1000 : node60251;
																assign node60251 = (inp[12]) ? 4'b1000 : 4'b1100;
															assign node60255 = (inp[12]) ? 4'b1110 : 4'b1000;
														assign node60258 = (inp[9]) ? node60260 : 4'b1110;
															assign node60260 = (inp[10]) ? 4'b1010 : 4'b1110;
												assign node60263 = (inp[5]) ? node60283 : node60264;
													assign node60264 = (inp[9]) ? node60272 : node60265;
														assign node60265 = (inp[4]) ? node60267 : 4'b1000;
															assign node60267 = (inp[12]) ? 4'b1110 : node60268;
																assign node60268 = (inp[10]) ? 4'b1110 : 4'b1000;
														assign node60272 = (inp[4]) ? node60278 : node60273;
															assign node60273 = (inp[10]) ? 4'b1110 : node60274;
																assign node60274 = (inp[12]) ? 4'b1110 : 4'b1000;
															assign node60278 = (inp[12]) ? 4'b1010 : node60279;
																assign node60279 = (inp[10]) ? 4'b1010 : 4'b1110;
													assign node60283 = (inp[9]) ? node60293 : node60284;
														assign node60284 = (inp[4]) ? node60288 : node60285;
															assign node60285 = (inp[10]) ? 4'b1010 : 4'b1110;
															assign node60288 = (inp[12]) ? 4'b1110 : node60289;
																assign node60289 = (inp[10]) ? 4'b1110 : 4'b1010;
														assign node60293 = (inp[4]) ? node60299 : node60294;
															assign node60294 = (inp[10]) ? 4'b1110 : node60295;
																assign node60295 = (inp[12]) ? 4'b1110 : 4'b1010;
															assign node60299 = (inp[10]) ? 4'b1010 : node60300;
																assign node60300 = (inp[12]) ? 4'b1010 : 4'b1110;
										assign node60304 = (inp[15]) ? node60378 : node60305;
											assign node60305 = (inp[5]) ? node60345 : node60306;
												assign node60306 = (inp[3]) ? node60326 : node60307;
													assign node60307 = (inp[4]) ? node60315 : node60308;
														assign node60308 = (inp[10]) ? 4'b1100 : node60309;
															assign node60309 = (inp[12]) ? 4'b1100 : node60310;
																assign node60310 = (inp[9]) ? 4'b1000 : 4'b1100;
														assign node60315 = (inp[9]) ? node60321 : node60316;
															assign node60316 = (inp[12]) ? 4'b1100 : node60317;
																assign node60317 = (inp[10]) ? 4'b1100 : 4'b1000;
															assign node60321 = (inp[10]) ? 4'b1000 : node60322;
																assign node60322 = (inp[12]) ? 4'b1000 : 4'b1100;
													assign node60326 = (inp[12]) ? node60340 : node60327;
														assign node60327 = (inp[9]) ? node60333 : node60328;
															assign node60328 = (inp[4]) ? node60330 : 4'b1000;
																assign node60330 = (inp[10]) ? 4'b1110 : 4'b1000;
															assign node60333 = (inp[4]) ? node60337 : node60334;
																assign node60334 = (inp[10]) ? 4'b1110 : 4'b1000;
																assign node60337 = (inp[10]) ? 4'b1010 : 4'b1110;
														assign node60340 = (inp[9]) ? node60342 : 4'b1110;
															assign node60342 = (inp[4]) ? 4'b1010 : 4'b1110;
												assign node60345 = (inp[3]) ? node60355 : node60346;
													assign node60346 = (inp[9]) ? node60350 : node60347;
														assign node60347 = (inp[4]) ? 4'b1110 : 4'b1000;
														assign node60350 = (inp[4]) ? node60352 : 4'b1110;
															assign node60352 = (inp[12]) ? 4'b1010 : 4'b1110;
													assign node60355 = (inp[12]) ? node60369 : node60356;
														assign node60356 = (inp[10]) ? node60362 : node60357;
															assign node60357 = (inp[4]) ? node60359 : 4'b1010;
																assign node60359 = (inp[9]) ? 4'b1110 : 4'b1010;
															assign node60362 = (inp[9]) ? node60366 : node60363;
																assign node60363 = (inp[4]) ? 4'b1110 : 4'b1010;
																assign node60366 = (inp[4]) ? 4'b1010 : 4'b1110;
														assign node60369 = (inp[10]) ? 4'b1010 : node60370;
															assign node60370 = (inp[4]) ? node60374 : node60371;
																assign node60371 = (inp[9]) ? 4'b1110 : 4'b1010;
																assign node60374 = (inp[9]) ? 4'b1010 : 4'b1110;
											assign node60378 = (inp[3]) ? node60422 : node60379;
												assign node60379 = (inp[5]) ? node60401 : node60380;
													assign node60380 = (inp[12]) ? node60394 : node60381;
														assign node60381 = (inp[10]) ? node60387 : node60382;
															assign node60382 = (inp[9]) ? 4'b1110 : node60383;
																assign node60383 = (inp[4]) ? 4'b1010 : 4'b1110;
															assign node60387 = (inp[4]) ? node60391 : node60388;
																assign node60388 = (inp[9]) ? 4'b1110 : 4'b1010;
																assign node60391 = (inp[9]) ? 4'b1010 : 4'b1110;
														assign node60394 = (inp[9]) ? node60398 : node60395;
															assign node60395 = (inp[4]) ? 4'b1110 : 4'b1010;
															assign node60398 = (inp[4]) ? 4'b1010 : 4'b1110;
													assign node60401 = (inp[9]) ? node60411 : node60402;
														assign node60402 = (inp[4]) ? node60408 : node60403;
															assign node60403 = (inp[10]) ? 4'b1010 : node60404;
																assign node60404 = (inp[12]) ? 4'b1010 : 4'b1110;
															assign node60408 = (inp[12]) ? 4'b1100 : 4'b1010;
														assign node60411 = (inp[4]) ? node60417 : node60412;
															assign node60412 = (inp[10]) ? 4'b1100 : node60413;
																assign node60413 = (inp[12]) ? 4'b1100 : 4'b1010;
															assign node60417 = (inp[10]) ? 4'b1000 : node60418;
																assign node60418 = (inp[12]) ? 4'b1000 : 4'b1100;
												assign node60422 = (inp[5]) ? node60430 : node60423;
													assign node60423 = (inp[4]) ? node60427 : node60424;
														assign node60424 = (inp[9]) ? 4'b1100 : 4'b1010;
														assign node60427 = (inp[9]) ? 4'b1000 : 4'b1100;
													assign node60430 = (inp[12]) ? node60440 : node60431;
														assign node60431 = (inp[4]) ? 4'b1000 : node60432;
															assign node60432 = (inp[9]) ? node60436 : node60433;
																assign node60433 = (inp[10]) ? 4'b1000 : 4'b1100;
																assign node60436 = (inp[10]) ? 4'b1100 : 4'b1000;
														assign node60440 = (inp[4]) ? node60444 : node60441;
															assign node60441 = (inp[9]) ? 4'b1100 : 4'b1000;
															assign node60444 = (inp[9]) ? 4'b1000 : 4'b1100;
									assign node60447 = (inp[4]) ? node60575 : node60448;
										assign node60448 = (inp[9]) ? node60512 : node60449;
											assign node60449 = (inp[10]) ? node60489 : node60450;
												assign node60450 = (inp[12]) ? node60468 : node60451;
													assign node60451 = (inp[15]) ? node60459 : node60452;
														assign node60452 = (inp[0]) ? node60454 : 4'b0111;
															assign node60454 = (inp[3]) ? node60456 : 4'b0101;
																assign node60456 = (inp[5]) ? 4'b0111 : 4'b0101;
														assign node60459 = (inp[0]) ? node60465 : node60460;
															assign node60460 = (inp[5]) ? node60462 : 4'b0101;
																assign node60462 = (inp[3]) ? 4'b0111 : 4'b0101;
															assign node60465 = (inp[3]) ? 4'b0101 : 4'b0111;
													assign node60468 = (inp[5]) ? node60480 : node60469;
														assign node60469 = (inp[3]) ? node60475 : node60470;
															assign node60470 = (inp[0]) ? 4'b0011 : node60471;
																assign node60471 = (inp[15]) ? 4'b0001 : 4'b0011;
															assign node60475 = (inp[15]) ? node60477 : 4'b0001;
																assign node60477 = (inp[0]) ? 4'b0011 : 4'b0001;
														assign node60480 = (inp[0]) ? node60482 : 4'b0011;
															assign node60482 = (inp[3]) ? node60486 : node60483;
																assign node60483 = (inp[15]) ? 4'b0011 : 4'b0001;
																assign node60486 = (inp[15]) ? 4'b0001 : 4'b0011;
												assign node60489 = (inp[15]) ? node60501 : node60490;
													assign node60490 = (inp[0]) ? node60496 : node60491;
														assign node60491 = (inp[5]) ? node60493 : 4'b0011;
															assign node60493 = (inp[3]) ? 4'b0001 : 4'b0011;
														assign node60496 = (inp[3]) ? node60498 : 4'b0001;
															assign node60498 = (inp[5]) ? 4'b0011 : 4'b0001;
													assign node60501 = (inp[0]) ? node60507 : node60502;
														assign node60502 = (inp[5]) ? node60504 : 4'b0001;
															assign node60504 = (inp[3]) ? 4'b0011 : 4'b0001;
														assign node60507 = (inp[3]) ? node60509 : 4'b0011;
															assign node60509 = (inp[5]) ? 4'b0001 : 4'b0011;
											assign node60512 = (inp[10]) ? node60552 : node60513;
												assign node60513 = (inp[12]) ? node60533 : node60514;
													assign node60514 = (inp[0]) ? node60524 : node60515;
														assign node60515 = (inp[15]) ? node60521 : node60516;
															assign node60516 = (inp[5]) ? node60518 : 4'b0011;
																assign node60518 = (inp[3]) ? 4'b0001 : 4'b0011;
															assign node60521 = (inp[3]) ? 4'b0011 : 4'b0001;
														assign node60524 = (inp[15]) ? node60530 : node60525;
															assign node60525 = (inp[5]) ? node60527 : 4'b0001;
																assign node60527 = (inp[3]) ? 4'b0011 : 4'b0001;
															assign node60530 = (inp[3]) ? 4'b0001 : 4'b0011;
													assign node60533 = (inp[0]) ? node60541 : node60534;
														assign node60534 = (inp[15]) ? 4'b0111 : node60535;
															assign node60535 = (inp[3]) ? 4'b0101 : node60536;
																assign node60536 = (inp[5]) ? 4'b0101 : 4'b0111;
														assign node60541 = (inp[15]) ? node60547 : node60542;
															assign node60542 = (inp[3]) ? 4'b0111 : node60543;
																assign node60543 = (inp[5]) ? 4'b0111 : 4'b0101;
															assign node60547 = (inp[5]) ? 4'b0101 : node60548;
																assign node60548 = (inp[3]) ? 4'b0101 : 4'b0111;
												assign node60552 = (inp[15]) ? node60564 : node60553;
													assign node60553 = (inp[0]) ? node60559 : node60554;
														assign node60554 = (inp[5]) ? 4'b0101 : node60555;
															assign node60555 = (inp[3]) ? 4'b0101 : 4'b0111;
														assign node60559 = (inp[3]) ? 4'b0111 : node60560;
															assign node60560 = (inp[5]) ? 4'b0111 : 4'b0101;
													assign node60564 = (inp[0]) ? node60570 : node60565;
														assign node60565 = (inp[5]) ? 4'b0111 : node60566;
															assign node60566 = (inp[3]) ? 4'b0111 : 4'b0101;
														assign node60570 = (inp[3]) ? 4'b0101 : node60571;
															assign node60571 = (inp[5]) ? 4'b0101 : 4'b0111;
										assign node60575 = (inp[9]) ? node60637 : node60576;
											assign node60576 = (inp[12]) ? node60600 : node60577;
												assign node60577 = (inp[10]) ? node60591 : node60578;
													assign node60578 = (inp[0]) ? node60584 : node60579;
														assign node60579 = (inp[15]) ? node60581 : 4'b0011;
															assign node60581 = (inp[3]) ? 4'b0011 : 4'b0001;
														assign node60584 = (inp[15]) ? node60586 : 4'b0001;
															assign node60586 = (inp[3]) ? node60588 : 4'b0011;
																assign node60588 = (inp[5]) ? 4'b0001 : 4'b0011;
													assign node60591 = (inp[3]) ? 4'b0101 : node60592;
														assign node60592 = (inp[5]) ? node60594 : 4'b0111;
															assign node60594 = (inp[0]) ? 4'b0101 : node60595;
																assign node60595 = (inp[15]) ? 4'b0111 : 4'b0101;
												assign node60600 = (inp[10]) ? node60616 : node60601;
													assign node60601 = (inp[5]) ? 4'b0101 : node60602;
														assign node60602 = (inp[15]) ? node60608 : node60603;
															assign node60603 = (inp[3]) ? node60605 : 4'b0101;
																assign node60605 = (inp[0]) ? 4'b0111 : 4'b0101;
															assign node60608 = (inp[3]) ? node60612 : node60609;
																assign node60609 = (inp[0]) ? 4'b0111 : 4'b0101;
																assign node60612 = (inp[0]) ? 4'b0101 : 4'b0111;
													assign node60616 = (inp[3]) ? node60632 : node60617;
														assign node60617 = (inp[15]) ? node60625 : node60618;
															assign node60618 = (inp[0]) ? node60622 : node60619;
																assign node60619 = (inp[5]) ? 4'b0101 : 4'b0111;
																assign node60622 = (inp[5]) ? 4'b0111 : 4'b0101;
															assign node60625 = (inp[0]) ? node60629 : node60626;
																assign node60626 = (inp[5]) ? 4'b0111 : 4'b0101;
																assign node60629 = (inp[5]) ? 4'b0101 : 4'b0111;
														assign node60632 = (inp[15]) ? 4'b0111 : node60633;
															assign node60633 = (inp[0]) ? 4'b0111 : 4'b0101;
											assign node60637 = (inp[12]) ? node60667 : node60638;
												assign node60638 = (inp[10]) ? node60654 : node60639;
													assign node60639 = (inp[15]) ? node60643 : node60640;
														assign node60640 = (inp[0]) ? 4'b0111 : 4'b0101;
														assign node60643 = (inp[0]) ? node60649 : node60644;
															assign node60644 = (inp[3]) ? 4'b0111 : node60645;
																assign node60645 = (inp[5]) ? 4'b0111 : 4'b0101;
															assign node60649 = (inp[5]) ? 4'b0101 : node60650;
																assign node60650 = (inp[3]) ? 4'b0101 : 4'b0111;
													assign node60654 = (inp[0]) ? node60660 : node60655;
														assign node60655 = (inp[3]) ? node60657 : 4'b0011;
															assign node60657 = (inp[15]) ? 4'b0011 : 4'b0001;
														assign node60660 = (inp[15]) ? 4'b0001 : node60661;
															assign node60661 = (inp[3]) ? 4'b0011 : node60662;
																assign node60662 = (inp[5]) ? 4'b0011 : 4'b0001;
												assign node60667 = (inp[15]) ? node60679 : node60668;
													assign node60668 = (inp[0]) ? node60674 : node60669;
														assign node60669 = (inp[3]) ? 4'b0001 : node60670;
															assign node60670 = (inp[5]) ? 4'b0001 : 4'b0011;
														assign node60674 = (inp[5]) ? 4'b0011 : node60675;
															assign node60675 = (inp[3]) ? 4'b0011 : 4'b0001;
													assign node60679 = (inp[0]) ? node60685 : node60680;
														assign node60680 = (inp[3]) ? 4'b0011 : node60681;
															assign node60681 = (inp[5]) ? 4'b0011 : 4'b0001;
														assign node60685 = (inp[5]) ? 4'b0001 : node60686;
															assign node60686 = (inp[3]) ? 4'b0001 : 4'b0011;
								assign node60690 = (inp[3]) ? node60920 : node60691;
									assign node60691 = (inp[12]) ? node60823 : node60692;
										assign node60692 = (inp[15]) ? node60756 : node60693;
											assign node60693 = (inp[0]) ? node60727 : node60694;
												assign node60694 = (inp[5]) ? node60710 : node60695;
													assign node60695 = (inp[4]) ? node60703 : node60696;
														assign node60696 = (inp[9]) ? node60700 : node60697;
															assign node60697 = (inp[10]) ? 4'b0011 : 4'b0111;
															assign node60700 = (inp[10]) ? 4'b0111 : 4'b0011;
														assign node60703 = (inp[9]) ? node60707 : node60704;
															assign node60704 = (inp[10]) ? 4'b0111 : 4'b0011;
															assign node60707 = (inp[10]) ? 4'b0011 : 4'b0111;
													assign node60710 = (inp[10]) ? node60720 : node60711;
														assign node60711 = (inp[2]) ? 4'b0011 : node60712;
															assign node60712 = (inp[4]) ? node60716 : node60713;
																assign node60713 = (inp[9]) ? 4'b0011 : 4'b0111;
																assign node60716 = (inp[9]) ? 4'b0101 : 4'b0011;
														assign node60720 = (inp[4]) ? node60724 : node60721;
															assign node60721 = (inp[9]) ? 4'b0101 : 4'b0011;
															assign node60724 = (inp[9]) ? 4'b0001 : 4'b0101;
												assign node60727 = (inp[5]) ? node60741 : node60728;
													assign node60728 = (inp[10]) ? node60736 : node60729;
														assign node60729 = (inp[9]) ? node60733 : node60730;
															assign node60730 = (inp[4]) ? 4'b0001 : 4'b0101;
															assign node60733 = (inp[4]) ? 4'b0101 : 4'b0001;
														assign node60736 = (inp[9]) ? node60738 : 4'b0101;
															assign node60738 = (inp[4]) ? 4'b0001 : 4'b0101;
													assign node60741 = (inp[10]) ? node60749 : node60742;
														assign node60742 = (inp[9]) ? node60746 : node60743;
															assign node60743 = (inp[4]) ? 4'b0001 : 4'b0101;
															assign node60746 = (inp[4]) ? 4'b0111 : 4'b0001;
														assign node60749 = (inp[9]) ? node60753 : node60750;
															assign node60750 = (inp[4]) ? 4'b0111 : 4'b0001;
															assign node60753 = (inp[4]) ? 4'b0011 : 4'b0111;
											assign node60756 = (inp[0]) ? node60794 : node60757;
												assign node60757 = (inp[5]) ? node60779 : node60758;
													assign node60758 = (inp[9]) ? node60772 : node60759;
														assign node60759 = (inp[2]) ? node60767 : node60760;
															assign node60760 = (inp[4]) ? node60764 : node60761;
																assign node60761 = (inp[10]) ? 4'b0001 : 4'b0101;
																assign node60764 = (inp[10]) ? 4'b0101 : 4'b0001;
															assign node60767 = (inp[10]) ? node60769 : 4'b0101;
																assign node60769 = (inp[4]) ? 4'b0101 : 4'b0001;
														assign node60772 = (inp[4]) ? node60776 : node60773;
															assign node60773 = (inp[10]) ? 4'b0101 : 4'b0001;
															assign node60776 = (inp[10]) ? 4'b0001 : 4'b0101;
													assign node60779 = (inp[10]) ? node60787 : node60780;
														assign node60780 = (inp[4]) ? node60784 : node60781;
															assign node60781 = (inp[9]) ? 4'b0001 : 4'b0101;
															assign node60784 = (inp[9]) ? 4'b0111 : 4'b0001;
														assign node60787 = (inp[9]) ? node60791 : node60788;
															assign node60788 = (inp[4]) ? 4'b0111 : 4'b0001;
															assign node60791 = (inp[4]) ? 4'b0011 : 4'b0111;
												assign node60794 = (inp[5]) ? node60808 : node60795;
													assign node60795 = (inp[4]) ? node60801 : node60796;
														assign node60796 = (inp[9]) ? 4'b0111 : node60797;
															assign node60797 = (inp[10]) ? 4'b0011 : 4'b0111;
														assign node60801 = (inp[9]) ? node60805 : node60802;
															assign node60802 = (inp[10]) ? 4'b0111 : 4'b0011;
															assign node60805 = (inp[10]) ? 4'b0011 : 4'b0111;
													assign node60808 = (inp[10]) ? node60816 : node60809;
														assign node60809 = (inp[4]) ? node60813 : node60810;
															assign node60810 = (inp[9]) ? 4'b0011 : 4'b0111;
															assign node60813 = (inp[9]) ? 4'b0101 : 4'b0011;
														assign node60816 = (inp[9]) ? node60820 : node60817;
															assign node60817 = (inp[2]) ? 4'b0011 : 4'b0101;
															assign node60820 = (inp[4]) ? 4'b0001 : 4'b0101;
										assign node60823 = (inp[9]) ? node60871 : node60824;
											assign node60824 = (inp[4]) ? node60832 : node60825;
												assign node60825 = (inp[0]) ? node60829 : node60826;
													assign node60826 = (inp[15]) ? 4'b0001 : 4'b0011;
													assign node60829 = (inp[15]) ? 4'b0011 : 4'b0001;
												assign node60832 = (inp[15]) ? node60848 : node60833;
													assign node60833 = (inp[2]) ? node60841 : node60834;
														assign node60834 = (inp[5]) ? node60838 : node60835;
															assign node60835 = (inp[0]) ? 4'b0101 : 4'b0111;
															assign node60838 = (inp[0]) ? 4'b0111 : 4'b0101;
														assign node60841 = (inp[0]) ? node60845 : node60842;
															assign node60842 = (inp[5]) ? 4'b0101 : 4'b0111;
															assign node60845 = (inp[5]) ? 4'b0111 : 4'b0101;
													assign node60848 = (inp[10]) ? node60864 : node60849;
														assign node60849 = (inp[2]) ? node60857 : node60850;
															assign node60850 = (inp[5]) ? node60854 : node60851;
																assign node60851 = (inp[0]) ? 4'b0111 : 4'b0101;
																assign node60854 = (inp[0]) ? 4'b0101 : 4'b0111;
															assign node60857 = (inp[0]) ? node60861 : node60858;
																assign node60858 = (inp[5]) ? 4'b0111 : 4'b0101;
																assign node60861 = (inp[5]) ? 4'b0101 : 4'b0111;
														assign node60864 = (inp[5]) ? node60868 : node60865;
															assign node60865 = (inp[0]) ? 4'b0111 : 4'b0101;
															assign node60868 = (inp[0]) ? 4'b0101 : 4'b0111;
											assign node60871 = (inp[4]) ? node60903 : node60872;
												assign node60872 = (inp[5]) ? node60896 : node60873;
													assign node60873 = (inp[10]) ? node60881 : node60874;
														assign node60874 = (inp[2]) ? 4'b0111 : node60875;
															assign node60875 = (inp[15]) ? 4'b0111 : node60876;
																assign node60876 = (inp[0]) ? 4'b0101 : 4'b0111;
														assign node60881 = (inp[2]) ? node60889 : node60882;
															assign node60882 = (inp[15]) ? node60886 : node60883;
																assign node60883 = (inp[0]) ? 4'b0101 : 4'b0111;
																assign node60886 = (inp[0]) ? 4'b0111 : 4'b0101;
															assign node60889 = (inp[0]) ? node60893 : node60890;
																assign node60890 = (inp[15]) ? 4'b0101 : 4'b0111;
																assign node60893 = (inp[15]) ? 4'b0111 : 4'b0101;
													assign node60896 = (inp[0]) ? node60900 : node60897;
														assign node60897 = (inp[15]) ? 4'b0111 : 4'b0101;
														assign node60900 = (inp[15]) ? 4'b0101 : 4'b0111;
												assign node60903 = (inp[15]) ? node60913 : node60904;
													assign node60904 = (inp[2]) ? 4'b0011 : node60905;
														assign node60905 = (inp[5]) ? node60909 : node60906;
															assign node60906 = (inp[0]) ? 4'b0001 : 4'b0011;
															assign node60909 = (inp[0]) ? 4'b0011 : 4'b0001;
													assign node60913 = (inp[0]) ? node60917 : node60914;
														assign node60914 = (inp[5]) ? 4'b0011 : 4'b0001;
														assign node60917 = (inp[5]) ? 4'b0001 : 4'b0011;
									assign node60920 = (inp[0]) ? node61012 : node60921;
										assign node60921 = (inp[15]) ? node60949 : node60922;
											assign node60922 = (inp[4]) ? node60938 : node60923;
												assign node60923 = (inp[9]) ? node60931 : node60924;
													assign node60924 = (inp[5]) ? node60926 : 4'b0011;
														assign node60926 = (inp[10]) ? 4'b0001 : node60927;
															assign node60927 = (inp[12]) ? 4'b0001 : 4'b0101;
													assign node60931 = (inp[12]) ? 4'b0101 : node60932;
														assign node60932 = (inp[10]) ? 4'b0101 : node60933;
															assign node60933 = (inp[5]) ? 4'b0001 : 4'b0011;
												assign node60938 = (inp[9]) ? node60944 : node60939;
													assign node60939 = (inp[10]) ? 4'b0101 : node60940;
														assign node60940 = (inp[12]) ? 4'b0101 : 4'b0001;
													assign node60944 = (inp[12]) ? 4'b0001 : node60945;
														assign node60945 = (inp[10]) ? 4'b0001 : 4'b0101;
											assign node60949 = (inp[5]) ? node60973 : node60950;
												assign node60950 = (inp[9]) ? node60962 : node60951;
													assign node60951 = (inp[4]) ? node60957 : node60952;
														assign node60952 = (inp[10]) ? 4'b0001 : node60953;
															assign node60953 = (inp[12]) ? 4'b0001 : 4'b0101;
														assign node60957 = (inp[10]) ? 4'b0111 : node60958;
															assign node60958 = (inp[12]) ? 4'b0111 : 4'b0001;
													assign node60962 = (inp[4]) ? node60968 : node60963;
														assign node60963 = (inp[10]) ? 4'b0111 : node60964;
															assign node60964 = (inp[12]) ? 4'b0111 : 4'b0001;
														assign node60968 = (inp[10]) ? 4'b0011 : node60969;
															assign node60969 = (inp[12]) ? 4'b0011 : 4'b0111;
												assign node60973 = (inp[2]) ? node60991 : node60974;
													assign node60974 = (inp[12]) ? node60986 : node60975;
														assign node60975 = (inp[4]) ? node60981 : node60976;
															assign node60976 = (inp[10]) ? node60978 : 4'b0111;
																assign node60978 = (inp[9]) ? 4'b0111 : 4'b0011;
															assign node60981 = (inp[9]) ? node60983 : 4'b0011;
																assign node60983 = (inp[10]) ? 4'b0011 : 4'b0111;
														assign node60986 = (inp[10]) ? 4'b0111 : node60987;
															assign node60987 = (inp[9]) ? 4'b0011 : 4'b0111;
													assign node60991 = (inp[9]) ? node61003 : node60992;
														assign node60992 = (inp[4]) ? node60998 : node60993;
															assign node60993 = (inp[12]) ? 4'b0011 : node60994;
																assign node60994 = (inp[10]) ? 4'b0011 : 4'b0111;
															assign node60998 = (inp[10]) ? 4'b0111 : node60999;
																assign node60999 = (inp[12]) ? 4'b0111 : 4'b0011;
														assign node61003 = (inp[4]) ? node61009 : node61004;
															assign node61004 = (inp[10]) ? 4'b0111 : node61005;
																assign node61005 = (inp[12]) ? 4'b0111 : 4'b0011;
															assign node61009 = (inp[12]) ? 4'b0011 : 4'b0111;
										assign node61012 = (inp[15]) ? node61074 : node61013;
											assign node61013 = (inp[5]) ? node61037 : node61014;
												assign node61014 = (inp[4]) ? node61026 : node61015;
													assign node61015 = (inp[9]) ? node61021 : node61016;
														assign node61016 = (inp[10]) ? 4'b0001 : node61017;
															assign node61017 = (inp[12]) ? 4'b0001 : 4'b0101;
														assign node61021 = (inp[10]) ? 4'b0111 : node61022;
															assign node61022 = (inp[12]) ? 4'b0111 : 4'b0001;
													assign node61026 = (inp[9]) ? node61032 : node61027;
														assign node61027 = (inp[10]) ? 4'b0111 : node61028;
															assign node61028 = (inp[12]) ? 4'b0111 : 4'b0001;
														assign node61032 = (inp[12]) ? 4'b0011 : node61033;
															assign node61033 = (inp[10]) ? 4'b0011 : 4'b0111;
												assign node61037 = (inp[2]) ? node61055 : node61038;
													assign node61038 = (inp[4]) ? node61046 : node61039;
														assign node61039 = (inp[12]) ? 4'b0011 : node61040;
															assign node61040 = (inp[9]) ? 4'b0011 : node61041;
																assign node61041 = (inp[10]) ? 4'b0011 : 4'b0111;
														assign node61046 = (inp[12]) ? node61052 : node61047;
															assign node61047 = (inp[9]) ? node61049 : 4'b0011;
																assign node61049 = (inp[10]) ? 4'b0011 : 4'b0111;
															assign node61052 = (inp[9]) ? 4'b0011 : 4'b0111;
													assign node61055 = (inp[12]) ? node61065 : node61056;
														assign node61056 = (inp[9]) ? node61058 : 4'b0111;
															assign node61058 = (inp[4]) ? node61062 : node61059;
																assign node61059 = (inp[10]) ? 4'b0111 : 4'b0011;
																assign node61062 = (inp[10]) ? 4'b0011 : 4'b0111;
														assign node61065 = (inp[10]) ? node61067 : 4'b0011;
															assign node61067 = (inp[4]) ? node61071 : node61068;
																assign node61068 = (inp[9]) ? 4'b0111 : 4'b0011;
																assign node61071 = (inp[9]) ? 4'b0011 : 4'b0111;
											assign node61074 = (inp[5]) ? node61090 : node61075;
												assign node61075 = (inp[4]) ? node61083 : node61076;
													assign node61076 = (inp[12]) ? 4'b0101 : node61077;
														assign node61077 = (inp[10]) ? node61079 : 4'b0011;
															assign node61079 = (inp[9]) ? 4'b0101 : 4'b0011;
													assign node61083 = (inp[9]) ? node61085 : 4'b0101;
														assign node61085 = (inp[12]) ? 4'b0001 : node61086;
															assign node61086 = (inp[10]) ? 4'b0001 : 4'b0101;
												assign node61090 = (inp[9]) ? node61102 : node61091;
													assign node61091 = (inp[4]) ? node61097 : node61092;
														assign node61092 = (inp[10]) ? 4'b0001 : node61093;
															assign node61093 = (inp[12]) ? 4'b0001 : 4'b0101;
														assign node61097 = (inp[12]) ? 4'b0101 : node61098;
															assign node61098 = (inp[10]) ? 4'b0101 : 4'b0001;
													assign node61102 = (inp[4]) ? node61108 : node61103;
														assign node61103 = (inp[12]) ? 4'b0101 : node61104;
															assign node61104 = (inp[10]) ? 4'b0101 : 4'b0001;
														assign node61108 = (inp[10]) ? 4'b0001 : node61109;
															assign node61109 = (inp[12]) ? 4'b0001 : 4'b0101;
							assign node61113 = (inp[2]) ? node61703 : node61114;
								assign node61114 = (inp[14]) ? node61438 : node61115;
									assign node61115 = (inp[12]) ? node61293 : node61116;
										assign node61116 = (inp[0]) ? node61200 : node61117;
											assign node61117 = (inp[4]) ? node61151 : node61118;
												assign node61118 = (inp[15]) ? node61132 : node61119;
													assign node61119 = (inp[5]) ? node61127 : node61120;
														assign node61120 = (inp[9]) ? node61124 : node61121;
															assign node61121 = (inp[10]) ? 4'b0011 : 4'b0111;
															assign node61124 = (inp[10]) ? 4'b0111 : 4'b0011;
														assign node61127 = (inp[9]) ? 4'b0101 : node61128;
															assign node61128 = (inp[10]) ? 4'b0001 : 4'b0101;
													assign node61132 = (inp[3]) ? node61142 : node61133;
														assign node61133 = (inp[5]) ? node61139 : node61134;
															assign node61134 = (inp[10]) ? node61136 : 4'b0001;
																assign node61136 = (inp[9]) ? 4'b0101 : 4'b0001;
															assign node61139 = (inp[9]) ? 4'b0001 : 4'b0101;
														assign node61142 = (inp[5]) ? node61146 : node61143;
															assign node61143 = (inp[10]) ? 4'b0111 : 4'b0101;
															assign node61146 = (inp[10]) ? 4'b0011 : node61147;
																assign node61147 = (inp[9]) ? 4'b0011 : 4'b0111;
												assign node61151 = (inp[15]) ? node61179 : node61152;
													assign node61152 = (inp[3]) ? node61166 : node61153;
														assign node61153 = (inp[5]) ? node61159 : node61154;
															assign node61154 = (inp[10]) ? 4'b0011 : node61155;
																assign node61155 = (inp[9]) ? 4'b0111 : 4'b0011;
															assign node61159 = (inp[10]) ? node61163 : node61160;
																assign node61160 = (inp[9]) ? 4'b0101 : 4'b0011;
																assign node61163 = (inp[9]) ? 4'b0001 : 4'b0101;
														assign node61166 = (inp[5]) ? node61172 : node61167;
															assign node61167 = (inp[9]) ? node61169 : 4'b0101;
																assign node61169 = (inp[10]) ? 4'b0001 : 4'b0101;
															assign node61172 = (inp[9]) ? node61176 : node61173;
																assign node61173 = (inp[10]) ? 4'b0101 : 4'b0001;
																assign node61176 = (inp[10]) ? 4'b0001 : 4'b0101;
													assign node61179 = (inp[5]) ? node61193 : node61180;
														assign node61180 = (inp[3]) ? node61188 : node61181;
															assign node61181 = (inp[9]) ? node61185 : node61182;
																assign node61182 = (inp[10]) ? 4'b0101 : 4'b0001;
																assign node61185 = (inp[10]) ? 4'b0001 : 4'b0101;
															assign node61188 = (inp[9]) ? node61190 : 4'b0001;
																assign node61190 = (inp[10]) ? 4'b0011 : 4'b0111;
														assign node61193 = (inp[3]) ? 4'b0111 : node61194;
															assign node61194 = (inp[9]) ? node61196 : 4'b0001;
																assign node61196 = (inp[10]) ? 4'b0011 : 4'b0111;
											assign node61200 = (inp[15]) ? node61242 : node61201;
												assign node61201 = (inp[3]) ? node61223 : node61202;
													assign node61202 = (inp[4]) ? node61210 : node61203;
														assign node61203 = (inp[10]) ? node61207 : node61204;
															assign node61204 = (inp[9]) ? 4'b0001 : 4'b0101;
															assign node61207 = (inp[9]) ? 4'b0101 : 4'b0001;
														assign node61210 = (inp[5]) ? node61216 : node61211;
															assign node61211 = (inp[9]) ? node61213 : 4'b0101;
																assign node61213 = (inp[10]) ? 4'b0001 : 4'b0101;
															assign node61216 = (inp[9]) ? node61220 : node61217;
																assign node61217 = (inp[10]) ? 4'b0111 : 4'b0001;
																assign node61220 = (inp[10]) ? 4'b0011 : 4'b0111;
													assign node61223 = (inp[5]) ? node61237 : node61224;
														assign node61224 = (inp[4]) ? node61230 : node61225;
															assign node61225 = (inp[10]) ? node61227 : 4'b0001;
																assign node61227 = (inp[9]) ? 4'b0111 : 4'b0001;
															assign node61230 = (inp[10]) ? node61234 : node61231;
																assign node61231 = (inp[9]) ? 4'b0111 : 4'b0001;
																assign node61234 = (inp[9]) ? 4'b0011 : 4'b0111;
														assign node61237 = (inp[10]) ? node61239 : 4'b0011;
															assign node61239 = (inp[4]) ? 4'b0011 : 4'b0111;
												assign node61242 = (inp[3]) ? node61272 : node61243;
													assign node61243 = (inp[5]) ? node61259 : node61244;
														assign node61244 = (inp[4]) ? node61252 : node61245;
															assign node61245 = (inp[9]) ? node61249 : node61246;
																assign node61246 = (inp[10]) ? 4'b0011 : 4'b0111;
																assign node61249 = (inp[10]) ? 4'b0111 : 4'b0011;
															assign node61252 = (inp[10]) ? node61256 : node61253;
																assign node61253 = (inp[9]) ? 4'b0111 : 4'b0011;
																assign node61256 = (inp[9]) ? 4'b0011 : 4'b0111;
														assign node61259 = (inp[4]) ? node61265 : node61260;
															assign node61260 = (inp[9]) ? 4'b0011 : node61261;
																assign node61261 = (inp[10]) ? 4'b0011 : 4'b0111;
															assign node61265 = (inp[9]) ? node61269 : node61266;
																assign node61266 = (inp[10]) ? 4'b0101 : 4'b0011;
																assign node61269 = (inp[10]) ? 4'b0001 : 4'b0101;
													assign node61272 = (inp[5]) ? node61286 : node61273;
														assign node61273 = (inp[10]) ? node61279 : node61274;
															assign node61274 = (inp[4]) ? node61276 : 4'b0011;
																assign node61276 = (inp[9]) ? 4'b0101 : 4'b0011;
															assign node61279 = (inp[9]) ? node61283 : node61280;
																assign node61280 = (inp[4]) ? 4'b0101 : 4'b0011;
																assign node61283 = (inp[4]) ? 4'b0001 : 4'b0101;
														assign node61286 = (inp[9]) ? node61288 : 4'b0101;
															assign node61288 = (inp[4]) ? node61290 : 4'b0001;
																assign node61290 = (inp[10]) ? 4'b0001 : 4'b0101;
										assign node61293 = (inp[10]) ? node61365 : node61294;
											assign node61294 = (inp[15]) ? node61330 : node61295;
												assign node61295 = (inp[0]) ? node61311 : node61296;
													assign node61296 = (inp[9]) ? node61308 : node61297;
														assign node61297 = (inp[4]) ? node61303 : node61298;
															assign node61298 = (inp[5]) ? node61300 : 4'b0011;
																assign node61300 = (inp[3]) ? 4'b0001 : 4'b0011;
															assign node61303 = (inp[3]) ? 4'b0101 : node61304;
																assign node61304 = (inp[5]) ? 4'b0101 : 4'b0111;
														assign node61308 = (inp[4]) ? 4'b0001 : 4'b0101;
													assign node61311 = (inp[3]) ? node61327 : node61312;
														assign node61312 = (inp[5]) ? node61320 : node61313;
															assign node61313 = (inp[9]) ? node61317 : node61314;
																assign node61314 = (inp[4]) ? 4'b0101 : 4'b0001;
																assign node61317 = (inp[4]) ? 4'b0001 : 4'b0101;
															assign node61320 = (inp[9]) ? node61324 : node61321;
																assign node61321 = (inp[4]) ? 4'b0111 : 4'b0001;
																assign node61324 = (inp[4]) ? 4'b0011 : 4'b0111;
														assign node61327 = (inp[5]) ? 4'b0011 : 4'b0111;
												assign node61330 = (inp[0]) ? node61346 : node61331;
													assign node61331 = (inp[5]) ? node61341 : node61332;
														assign node61332 = (inp[3]) ? node61334 : 4'b0001;
															assign node61334 = (inp[9]) ? node61338 : node61335;
																assign node61335 = (inp[4]) ? 4'b0111 : 4'b0001;
																assign node61338 = (inp[4]) ? 4'b0011 : 4'b0111;
														assign node61341 = (inp[4]) ? node61343 : 4'b0111;
															assign node61343 = (inp[9]) ? 4'b0011 : 4'b0111;
													assign node61346 = (inp[3]) ? node61358 : node61347;
														assign node61347 = (inp[5]) ? node61353 : node61348;
															assign node61348 = (inp[4]) ? node61350 : 4'b0111;
																assign node61350 = (inp[9]) ? 4'b0011 : 4'b0111;
															assign node61353 = (inp[9]) ? 4'b0101 : node61354;
																assign node61354 = (inp[4]) ? 4'b0101 : 4'b0011;
														assign node61358 = (inp[4]) ? node61362 : node61359;
															assign node61359 = (inp[9]) ? 4'b0101 : 4'b0001;
															assign node61362 = (inp[9]) ? 4'b0001 : 4'b0101;
											assign node61365 = (inp[15]) ? node61399 : node61366;
												assign node61366 = (inp[0]) ? node61382 : node61367;
													assign node61367 = (inp[3]) ? 4'b0101 : node61368;
														assign node61368 = (inp[5]) ? node61374 : node61369;
															assign node61369 = (inp[4]) ? 4'b0111 : node61370;
																assign node61370 = (inp[9]) ? 4'b0111 : 4'b0011;
															assign node61374 = (inp[9]) ? node61378 : node61375;
																assign node61375 = (inp[4]) ? 4'b0101 : 4'b0011;
																assign node61378 = (inp[4]) ? 4'b0001 : 4'b0101;
													assign node61382 = (inp[5]) ? node61392 : node61383;
														assign node61383 = (inp[4]) ? node61389 : node61384;
															assign node61384 = (inp[9]) ? node61386 : 4'b0001;
																assign node61386 = (inp[3]) ? 4'b0111 : 4'b0101;
															assign node61389 = (inp[9]) ? 4'b0011 : 4'b0111;
														assign node61392 = (inp[4]) ? node61396 : node61393;
															assign node61393 = (inp[9]) ? 4'b0111 : 4'b0011;
															assign node61396 = (inp[9]) ? 4'b0011 : 4'b0111;
												assign node61399 = (inp[0]) ? node61419 : node61400;
													assign node61400 = (inp[5]) ? node61410 : node61401;
														assign node61401 = (inp[4]) ? node61405 : node61402;
															assign node61402 = (inp[9]) ? 4'b0101 : 4'b0001;
															assign node61405 = (inp[9]) ? node61407 : 4'b0111;
																assign node61407 = (inp[3]) ? 4'b0011 : 4'b0001;
														assign node61410 = (inp[4]) ? node61416 : node61411;
															assign node61411 = (inp[9]) ? 4'b0111 : node61412;
																assign node61412 = (inp[3]) ? 4'b0011 : 4'b0001;
															assign node61416 = (inp[9]) ? 4'b0011 : 4'b0111;
													assign node61419 = (inp[5]) ? node61433 : node61420;
														assign node61420 = (inp[3]) ? node61426 : node61421;
															assign node61421 = (inp[4]) ? node61423 : 4'b0111;
																assign node61423 = (inp[9]) ? 4'b0011 : 4'b0111;
															assign node61426 = (inp[9]) ? node61430 : node61427;
																assign node61427 = (inp[4]) ? 4'b0101 : 4'b0011;
																assign node61430 = (inp[4]) ? 4'b0001 : 4'b0101;
														assign node61433 = (inp[9]) ? 4'b0001 : node61434;
															assign node61434 = (inp[4]) ? 4'b0101 : 4'b0001;
									assign node61438 = (inp[15]) ? node61562 : node61439;
										assign node61439 = (inp[0]) ? node61495 : node61440;
											assign node61440 = (inp[5]) ? node61472 : node61441;
												assign node61441 = (inp[3]) ? node61451 : node61442;
													assign node61442 = (inp[4]) ? node61444 : 4'b0110;
														assign node61444 = (inp[9]) ? 4'b0010 : node61445;
															assign node61445 = (inp[12]) ? 4'b0110 : node61446;
																assign node61446 = (inp[10]) ? 4'b0110 : 4'b0010;
													assign node61451 = (inp[9]) ? node61461 : node61452;
														assign node61452 = (inp[4]) ? node61456 : node61453;
															assign node61453 = (inp[10]) ? 4'b0010 : 4'b0110;
															assign node61456 = (inp[12]) ? 4'b0100 : node61457;
																assign node61457 = (inp[10]) ? 4'b0100 : 4'b0010;
														assign node61461 = (inp[4]) ? node61467 : node61462;
															assign node61462 = (inp[12]) ? 4'b0100 : node61463;
																assign node61463 = (inp[10]) ? 4'b0100 : 4'b0010;
															assign node61467 = (inp[12]) ? 4'b0000 : node61468;
																assign node61468 = (inp[10]) ? 4'b0000 : 4'b0100;
												assign node61472 = (inp[4]) ? node61484 : node61473;
													assign node61473 = (inp[9]) ? node61477 : node61474;
														assign node61474 = (inp[3]) ? 4'b0000 : 4'b0010;
														assign node61477 = (inp[10]) ? 4'b0100 : node61478;
															assign node61478 = (inp[12]) ? 4'b0100 : node61479;
																assign node61479 = (inp[3]) ? 4'b0000 : 4'b0010;
													assign node61484 = (inp[9]) ? node61490 : node61485;
														assign node61485 = (inp[10]) ? 4'b0100 : node61486;
															assign node61486 = (inp[12]) ? 4'b0100 : 4'b0000;
														assign node61490 = (inp[12]) ? 4'b0000 : node61491;
															assign node61491 = (inp[10]) ? 4'b0000 : 4'b0100;
											assign node61495 = (inp[5]) ? node61531 : node61496;
												assign node61496 = (inp[3]) ? node61512 : node61497;
													assign node61497 = (inp[9]) ? node61501 : node61498;
														assign node61498 = (inp[4]) ? 4'b0100 : 4'b0000;
														assign node61501 = (inp[4]) ? node61507 : node61502;
															assign node61502 = (inp[10]) ? 4'b0100 : node61503;
																assign node61503 = (inp[12]) ? 4'b0100 : 4'b0000;
															assign node61507 = (inp[10]) ? 4'b0000 : node61508;
																assign node61508 = (inp[12]) ? 4'b0000 : 4'b0100;
													assign node61512 = (inp[4]) ? node61522 : node61513;
														assign node61513 = (inp[9]) ? node61519 : node61514;
															assign node61514 = (inp[10]) ? 4'b0000 : node61515;
																assign node61515 = (inp[12]) ? 4'b0000 : 4'b0100;
															assign node61519 = (inp[12]) ? 4'b0110 : 4'b0000;
														assign node61522 = (inp[10]) ? node61528 : node61523;
															assign node61523 = (inp[9]) ? node61525 : 4'b0000;
																assign node61525 = (inp[12]) ? 4'b0010 : 4'b0110;
															assign node61528 = (inp[9]) ? 4'b0010 : 4'b0110;
												assign node61531 = (inp[3]) ? node61547 : node61532;
													assign node61532 = (inp[9]) ? node61540 : node61533;
														assign node61533 = (inp[4]) ? 4'b0110 : node61534;
															assign node61534 = (inp[10]) ? 4'b0000 : node61535;
																assign node61535 = (inp[12]) ? 4'b0000 : 4'b0100;
														assign node61540 = (inp[4]) ? node61542 : 4'b0110;
															assign node61542 = (inp[12]) ? 4'b0010 : node61543;
																assign node61543 = (inp[10]) ? 4'b0010 : 4'b0110;
													assign node61547 = (inp[4]) ? node61553 : node61548;
														assign node61548 = (inp[9]) ? node61550 : 4'b0010;
															assign node61550 = (inp[10]) ? 4'b0110 : 4'b0010;
														assign node61553 = (inp[9]) ? node61559 : node61554;
															assign node61554 = (inp[12]) ? 4'b0110 : node61555;
																assign node61555 = (inp[10]) ? 4'b0110 : 4'b0010;
															assign node61559 = (inp[10]) ? 4'b0010 : 4'b0110;
										assign node61562 = (inp[0]) ? node61632 : node61563;
											assign node61563 = (inp[3]) ? node61593 : node61564;
												assign node61564 = (inp[5]) ? node61580 : node61565;
													assign node61565 = (inp[4]) ? node61575 : node61566;
														assign node61566 = (inp[9]) ? node61572 : node61567;
															assign node61567 = (inp[10]) ? 4'b0000 : node61568;
																assign node61568 = (inp[12]) ? 4'b0000 : 4'b0100;
															assign node61572 = (inp[10]) ? 4'b0100 : 4'b0000;
														assign node61575 = (inp[9]) ? 4'b0000 : node61576;
															assign node61576 = (inp[12]) ? 4'b0100 : 4'b0000;
													assign node61580 = (inp[4]) ? node61586 : node61581;
														assign node61581 = (inp[12]) ? 4'b0000 : node61582;
															assign node61582 = (inp[9]) ? 4'b0000 : 4'b0100;
														assign node61586 = (inp[9]) ? node61590 : node61587;
															assign node61587 = (inp[12]) ? 4'b0110 : 4'b0000;
															assign node61590 = (inp[10]) ? 4'b0010 : 4'b0110;
												assign node61593 = (inp[5]) ? node61615 : node61594;
													assign node61594 = (inp[4]) ? node61604 : node61595;
														assign node61595 = (inp[9]) ? node61601 : node61596;
															assign node61596 = (inp[10]) ? 4'b0000 : node61597;
																assign node61597 = (inp[12]) ? 4'b0000 : 4'b0100;
															assign node61601 = (inp[12]) ? 4'b0110 : 4'b0000;
														assign node61604 = (inp[9]) ? node61610 : node61605;
															assign node61605 = (inp[12]) ? 4'b0110 : node61606;
																assign node61606 = (inp[10]) ? 4'b0110 : 4'b0000;
															assign node61610 = (inp[12]) ? 4'b0010 : node61611;
																assign node61611 = (inp[10]) ? 4'b0010 : 4'b0110;
													assign node61615 = (inp[4]) ? node61621 : node61616;
														assign node61616 = (inp[9]) ? node61618 : 4'b0010;
															assign node61618 = (inp[10]) ? 4'b0110 : 4'b0010;
														assign node61621 = (inp[9]) ? node61627 : node61622;
															assign node61622 = (inp[12]) ? 4'b0110 : node61623;
																assign node61623 = (inp[10]) ? 4'b0110 : 4'b0010;
															assign node61627 = (inp[10]) ? 4'b0010 : node61628;
																assign node61628 = (inp[12]) ? 4'b0010 : 4'b0110;
											assign node61632 = (inp[5]) ? node61670 : node61633;
												assign node61633 = (inp[3]) ? node61651 : node61634;
													assign node61634 = (inp[12]) ? node61644 : node61635;
														assign node61635 = (inp[4]) ? 4'b0010 : node61636;
															assign node61636 = (inp[10]) ? node61640 : node61637;
																assign node61637 = (inp[9]) ? 4'b0010 : 4'b0110;
																assign node61640 = (inp[9]) ? 4'b0110 : 4'b0010;
														assign node61644 = (inp[4]) ? node61648 : node61645;
															assign node61645 = (inp[9]) ? 4'b0110 : 4'b0010;
															assign node61648 = (inp[9]) ? 4'b0010 : 4'b0110;
													assign node61651 = (inp[9]) ? node61663 : node61652;
														assign node61652 = (inp[4]) ? node61658 : node61653;
															assign node61653 = (inp[10]) ? 4'b0010 : node61654;
																assign node61654 = (inp[12]) ? 4'b0010 : 4'b0110;
															assign node61658 = (inp[10]) ? 4'b0100 : node61659;
																assign node61659 = (inp[12]) ? 4'b0100 : 4'b0010;
														assign node61663 = (inp[4]) ? 4'b0000 : node61664;
															assign node61664 = (inp[10]) ? 4'b0100 : node61665;
																assign node61665 = (inp[12]) ? 4'b0100 : 4'b0010;
												assign node61670 = (inp[3]) ? node61686 : node61671;
													assign node61671 = (inp[4]) ? node61679 : node61672;
														assign node61672 = (inp[9]) ? node61676 : node61673;
															assign node61673 = (inp[12]) ? 4'b0010 : 4'b0110;
															assign node61676 = (inp[12]) ? 4'b0100 : 4'b0010;
														assign node61679 = (inp[9]) ? 4'b0000 : node61680;
															assign node61680 = (inp[12]) ? 4'b0100 : node61681;
																assign node61681 = (inp[10]) ? 4'b0100 : 4'b0010;
													assign node61686 = (inp[4]) ? node61692 : node61687;
														assign node61687 = (inp[9]) ? node61689 : 4'b0000;
															assign node61689 = (inp[12]) ? 4'b0100 : 4'b0000;
														assign node61692 = (inp[9]) ? node61698 : node61693;
															assign node61693 = (inp[12]) ? 4'b0100 : node61694;
																assign node61694 = (inp[10]) ? 4'b0100 : 4'b0000;
															assign node61698 = (inp[10]) ? 4'b0000 : node61699;
																assign node61699 = (inp[12]) ? 4'b0000 : 4'b0100;
								assign node61703 = (inp[12]) ? node61965 : node61704;
									assign node61704 = (inp[15]) ? node61840 : node61705;
										assign node61705 = (inp[0]) ? node61773 : node61706;
											assign node61706 = (inp[3]) ? node61734 : node61707;
												assign node61707 = (inp[5]) ? node61721 : node61708;
													assign node61708 = (inp[10]) ? node61716 : node61709;
														assign node61709 = (inp[4]) ? node61713 : node61710;
															assign node61710 = (inp[9]) ? 4'b0010 : 4'b0110;
															assign node61713 = (inp[9]) ? 4'b0110 : 4'b0010;
														assign node61716 = (inp[9]) ? 4'b0110 : node61717;
															assign node61717 = (inp[4]) ? 4'b0110 : 4'b0010;
													assign node61721 = (inp[9]) ? node61729 : node61722;
														assign node61722 = (inp[10]) ? node61726 : node61723;
															assign node61723 = (inp[4]) ? 4'b0010 : 4'b0110;
															assign node61726 = (inp[4]) ? 4'b0100 : 4'b0010;
														assign node61729 = (inp[4]) ? 4'b0100 : node61730;
															assign node61730 = (inp[10]) ? 4'b0100 : 4'b0010;
												assign node61734 = (inp[5]) ? node61750 : node61735;
													assign node61735 = (inp[9]) ? node61743 : node61736;
														assign node61736 = (inp[10]) ? node61740 : node61737;
															assign node61737 = (inp[4]) ? 4'b0010 : 4'b0110;
															assign node61740 = (inp[4]) ? 4'b0100 : 4'b0010;
														assign node61743 = (inp[14]) ? node61745 : 4'b0100;
															assign node61745 = (inp[4]) ? node61747 : 4'b0100;
																assign node61747 = (inp[10]) ? 4'b0000 : 4'b0100;
													assign node61750 = (inp[10]) ? node61758 : node61751;
														assign node61751 = (inp[4]) ? node61755 : node61752;
															assign node61752 = (inp[9]) ? 4'b0000 : 4'b0100;
															assign node61755 = (inp[9]) ? 4'b0100 : 4'b0000;
														assign node61758 = (inp[14]) ? node61766 : node61759;
															assign node61759 = (inp[4]) ? node61763 : node61760;
																assign node61760 = (inp[9]) ? 4'b0100 : 4'b0000;
																assign node61763 = (inp[9]) ? 4'b0000 : 4'b0100;
															assign node61766 = (inp[4]) ? node61770 : node61767;
																assign node61767 = (inp[9]) ? 4'b0100 : 4'b0000;
																assign node61770 = (inp[9]) ? 4'b0000 : 4'b0100;
											assign node61773 = (inp[5]) ? node61807 : node61774;
												assign node61774 = (inp[3]) ? node61792 : node61775;
													assign node61775 = (inp[4]) ? node61783 : node61776;
														assign node61776 = (inp[10]) ? node61780 : node61777;
															assign node61777 = (inp[9]) ? 4'b0000 : 4'b0100;
															assign node61780 = (inp[9]) ? 4'b0100 : 4'b0000;
														assign node61783 = (inp[14]) ? 4'b0100 : node61784;
															assign node61784 = (inp[10]) ? node61788 : node61785;
																assign node61785 = (inp[9]) ? 4'b0100 : 4'b0000;
																assign node61788 = (inp[9]) ? 4'b0000 : 4'b0100;
													assign node61792 = (inp[10]) ? node61800 : node61793;
														assign node61793 = (inp[4]) ? node61797 : node61794;
															assign node61794 = (inp[9]) ? 4'b0000 : 4'b0100;
															assign node61797 = (inp[9]) ? 4'b0110 : 4'b0000;
														assign node61800 = (inp[4]) ? node61804 : node61801;
															assign node61801 = (inp[9]) ? 4'b0110 : 4'b0000;
															assign node61804 = (inp[9]) ? 4'b0010 : 4'b0110;
												assign node61807 = (inp[3]) ? node61821 : node61808;
													assign node61808 = (inp[4]) ? node61814 : node61809;
														assign node61809 = (inp[9]) ? 4'b0000 : node61810;
															assign node61810 = (inp[10]) ? 4'b0000 : 4'b0100;
														assign node61814 = (inp[10]) ? node61818 : node61815;
															assign node61815 = (inp[9]) ? 4'b0110 : 4'b0000;
															assign node61818 = (inp[9]) ? 4'b0010 : 4'b0110;
													assign node61821 = (inp[14]) ? node61831 : node61822;
														assign node61822 = (inp[4]) ? 4'b0110 : node61823;
															assign node61823 = (inp[9]) ? node61827 : node61824;
																assign node61824 = (inp[10]) ? 4'b0010 : 4'b0110;
																assign node61827 = (inp[10]) ? 4'b0110 : 4'b0010;
														assign node61831 = (inp[9]) ? 4'b0010 : node61832;
															assign node61832 = (inp[4]) ? node61836 : node61833;
																assign node61833 = (inp[10]) ? 4'b0010 : 4'b0110;
																assign node61836 = (inp[10]) ? 4'b0110 : 4'b0010;
										assign node61840 = (inp[9]) ? node61908 : node61841;
											assign node61841 = (inp[0]) ? node61877 : node61842;
												assign node61842 = (inp[5]) ? node61862 : node61843;
													assign node61843 = (inp[3]) ? node61857 : node61844;
														assign node61844 = (inp[14]) ? node61850 : node61845;
															assign node61845 = (inp[10]) ? node61847 : 4'b0000;
																assign node61847 = (inp[4]) ? 4'b0100 : 4'b0000;
															assign node61850 = (inp[10]) ? node61854 : node61851;
																assign node61851 = (inp[4]) ? 4'b0000 : 4'b0100;
																assign node61854 = (inp[4]) ? 4'b0100 : 4'b0000;
														assign node61857 = (inp[10]) ? 4'b0110 : node61858;
															assign node61858 = (inp[4]) ? 4'b0000 : 4'b0100;
													assign node61862 = (inp[3]) ? node61870 : node61863;
														assign node61863 = (inp[4]) ? node61867 : node61864;
															assign node61864 = (inp[10]) ? 4'b0000 : 4'b0100;
															assign node61867 = (inp[10]) ? 4'b0110 : 4'b0000;
														assign node61870 = (inp[10]) ? node61874 : node61871;
															assign node61871 = (inp[4]) ? 4'b0010 : 4'b0110;
															assign node61874 = (inp[4]) ? 4'b0110 : 4'b0010;
												assign node61877 = (inp[5]) ? node61895 : node61878;
													assign node61878 = (inp[3]) ? node61888 : node61879;
														assign node61879 = (inp[14]) ? node61881 : 4'b0110;
															assign node61881 = (inp[4]) ? node61885 : node61882;
																assign node61882 = (inp[10]) ? 4'b0010 : 4'b0110;
																assign node61885 = (inp[10]) ? 4'b0110 : 4'b0010;
														assign node61888 = (inp[4]) ? node61892 : node61889;
															assign node61889 = (inp[10]) ? 4'b0010 : 4'b0110;
															assign node61892 = (inp[10]) ? 4'b0100 : 4'b0010;
													assign node61895 = (inp[3]) ? node61901 : node61896;
														assign node61896 = (inp[10]) ? 4'b0100 : node61897;
															assign node61897 = (inp[4]) ? 4'b0010 : 4'b0110;
														assign node61901 = (inp[10]) ? node61905 : node61902;
															assign node61902 = (inp[4]) ? 4'b0000 : 4'b0100;
															assign node61905 = (inp[4]) ? 4'b0100 : 4'b0000;
											assign node61908 = (inp[0]) ? node61934 : node61909;
												assign node61909 = (inp[3]) ? node61925 : node61910;
													assign node61910 = (inp[5]) ? node61918 : node61911;
														assign node61911 = (inp[10]) ? node61915 : node61912;
															assign node61912 = (inp[4]) ? 4'b0100 : 4'b0000;
															assign node61915 = (inp[4]) ? 4'b0000 : 4'b0100;
														assign node61918 = (inp[4]) ? node61922 : node61919;
															assign node61919 = (inp[10]) ? 4'b0110 : 4'b0000;
															assign node61922 = (inp[10]) ? 4'b0010 : 4'b0110;
													assign node61925 = (inp[4]) ? node61931 : node61926;
														assign node61926 = (inp[10]) ? 4'b0110 : node61927;
															assign node61927 = (inp[5]) ? 4'b0010 : 4'b0000;
														assign node61931 = (inp[10]) ? 4'b0010 : 4'b0110;
												assign node61934 = (inp[5]) ? node61948 : node61935;
													assign node61935 = (inp[3]) ? node61943 : node61936;
														assign node61936 = (inp[10]) ? node61940 : node61937;
															assign node61937 = (inp[4]) ? 4'b0110 : 4'b0010;
															assign node61940 = (inp[4]) ? 4'b0010 : 4'b0110;
														assign node61943 = (inp[4]) ? node61945 : 4'b0010;
															assign node61945 = (inp[10]) ? 4'b0000 : 4'b0100;
													assign node61948 = (inp[3]) ? node61956 : node61949;
														assign node61949 = (inp[4]) ? node61953 : node61950;
															assign node61950 = (inp[10]) ? 4'b0100 : 4'b0010;
															assign node61953 = (inp[10]) ? 4'b0000 : 4'b0100;
														assign node61956 = (inp[14]) ? 4'b0100 : node61957;
															assign node61957 = (inp[4]) ? node61961 : node61958;
																assign node61958 = (inp[10]) ? 4'b0100 : 4'b0000;
																assign node61961 = (inp[10]) ? 4'b0000 : 4'b0100;
									assign node61965 = (inp[15]) ? node62029 : node61966;
										assign node61966 = (inp[0]) ? node61992 : node61967;
											assign node61967 = (inp[3]) ? node61983 : node61968;
												assign node61968 = (inp[5]) ? node61976 : node61969;
													assign node61969 = (inp[9]) ? node61973 : node61970;
														assign node61970 = (inp[4]) ? 4'b0110 : 4'b0010;
														assign node61973 = (inp[4]) ? 4'b0010 : 4'b0110;
													assign node61976 = (inp[4]) ? node61980 : node61977;
														assign node61977 = (inp[9]) ? 4'b0100 : 4'b0010;
														assign node61980 = (inp[9]) ? 4'b0000 : 4'b0100;
												assign node61983 = (inp[9]) ? node61989 : node61984;
													assign node61984 = (inp[4]) ? 4'b0100 : node61985;
														assign node61985 = (inp[5]) ? 4'b0000 : 4'b0010;
													assign node61989 = (inp[4]) ? 4'b0000 : 4'b0100;
											assign node61992 = (inp[5]) ? node62020 : node61993;
												assign node61993 = (inp[3]) ? node62013 : node61994;
													assign node61994 = (inp[14]) ? node62008 : node61995;
														assign node61995 = (inp[10]) ? node62001 : node61996;
															assign node61996 = (inp[4]) ? 4'b0100 : node61997;
																assign node61997 = (inp[9]) ? 4'b0100 : 4'b0000;
															assign node62001 = (inp[9]) ? node62005 : node62002;
																assign node62002 = (inp[4]) ? 4'b0100 : 4'b0000;
																assign node62005 = (inp[4]) ? 4'b0000 : 4'b0100;
														assign node62008 = (inp[4]) ? node62010 : 4'b0000;
															assign node62010 = (inp[9]) ? 4'b0000 : 4'b0100;
													assign node62013 = (inp[9]) ? node62017 : node62014;
														assign node62014 = (inp[4]) ? 4'b0110 : 4'b0000;
														assign node62017 = (inp[4]) ? 4'b0010 : 4'b0110;
												assign node62020 = (inp[4]) ? node62026 : node62021;
													assign node62021 = (inp[9]) ? 4'b0110 : node62022;
														assign node62022 = (inp[3]) ? 4'b0010 : 4'b0000;
													assign node62026 = (inp[9]) ? 4'b0010 : 4'b0110;
										assign node62029 = (inp[0]) ? node62063 : node62030;
											assign node62030 = (inp[3]) ? node62054 : node62031;
												assign node62031 = (inp[5]) ? node62047 : node62032;
													assign node62032 = (inp[10]) ? node62040 : node62033;
														assign node62033 = (inp[4]) ? node62037 : node62034;
															assign node62034 = (inp[9]) ? 4'b0100 : 4'b0000;
															assign node62037 = (inp[9]) ? 4'b0000 : 4'b0100;
														assign node62040 = (inp[9]) ? node62044 : node62041;
															assign node62041 = (inp[4]) ? 4'b0100 : 4'b0000;
															assign node62044 = (inp[4]) ? 4'b0000 : 4'b0100;
													assign node62047 = (inp[4]) ? node62051 : node62048;
														assign node62048 = (inp[9]) ? 4'b0110 : 4'b0000;
														assign node62051 = (inp[9]) ? 4'b0010 : 4'b0110;
												assign node62054 = (inp[9]) ? node62060 : node62055;
													assign node62055 = (inp[4]) ? 4'b0110 : node62056;
														assign node62056 = (inp[5]) ? 4'b0010 : 4'b0000;
													assign node62060 = (inp[4]) ? 4'b0010 : 4'b0110;
											assign node62063 = (inp[3]) ? node62091 : node62064;
												assign node62064 = (inp[5]) ? node62084 : node62065;
													assign node62065 = (inp[14]) ? node62073 : node62066;
														assign node62066 = (inp[10]) ? node62068 : 4'b0010;
															assign node62068 = (inp[4]) ? node62070 : 4'b0010;
																assign node62070 = (inp[9]) ? 4'b0010 : 4'b0110;
														assign node62073 = (inp[10]) ? node62079 : node62074;
															assign node62074 = (inp[4]) ? 4'b0010 : node62075;
																assign node62075 = (inp[9]) ? 4'b0110 : 4'b0010;
															assign node62079 = (inp[9]) ? 4'b0110 : node62080;
																assign node62080 = (inp[4]) ? 4'b0110 : 4'b0010;
													assign node62084 = (inp[4]) ? node62088 : node62085;
														assign node62085 = (inp[9]) ? 4'b0100 : 4'b0010;
														assign node62088 = (inp[9]) ? 4'b0000 : 4'b0100;
												assign node62091 = (inp[14]) ? node62101 : node62092;
													assign node62092 = (inp[9]) ? node62098 : node62093;
														assign node62093 = (inp[4]) ? 4'b0100 : node62094;
															assign node62094 = (inp[5]) ? 4'b0000 : 4'b0010;
														assign node62098 = (inp[4]) ? 4'b0000 : 4'b0100;
													assign node62101 = (inp[5]) ? node62109 : node62102;
														assign node62102 = (inp[10]) ? 4'b0100 : node62103;
															assign node62103 = (inp[9]) ? node62105 : 4'b0100;
																assign node62105 = (inp[4]) ? 4'b0000 : 4'b0100;
														assign node62109 = (inp[10]) ? node62113 : node62110;
															assign node62110 = (inp[4]) ? 4'b0000 : 4'b0100;
															assign node62113 = (inp[4]) ? 4'b0100 : 4'b0000;
					assign node62116 = (inp[14]) ? node64786 : node62117;
						assign node62117 = (inp[15]) ? node63429 : node62118;
							assign node62118 = (inp[0]) ? node62772 : node62119;
								assign node62119 = (inp[3]) ? node62421 : node62120;
									assign node62120 = (inp[5]) ? node62282 : node62121;
										assign node62121 = (inp[4]) ? node62203 : node62122;
											assign node62122 = (inp[9]) ? node62162 : node62123;
												assign node62123 = (inp[10]) ? node62139 : node62124;
													assign node62124 = (inp[12]) ? node62132 : node62125;
														assign node62125 = (inp[7]) ? 4'b0111 : node62126;
															assign node62126 = (inp[2]) ? 4'b0110 : node62127;
																assign node62127 = (inp[8]) ? 4'b0110 : 4'b0111;
														assign node62132 = (inp[2]) ? node62134 : 4'b0010;
															assign node62134 = (inp[7]) ? node62136 : 4'b0010;
																assign node62136 = (inp[8]) ? 4'b0010 : 4'b0011;
													assign node62139 = (inp[2]) ? node62147 : node62140;
														assign node62140 = (inp[7]) ? node62144 : node62141;
															assign node62141 = (inp[8]) ? 4'b0010 : 4'b0011;
															assign node62144 = (inp[8]) ? 4'b0011 : 4'b0010;
														assign node62147 = (inp[12]) ? node62155 : node62148;
															assign node62148 = (inp[7]) ? node62152 : node62149;
																assign node62149 = (inp[8]) ? 4'b0011 : 4'b0010;
																assign node62152 = (inp[8]) ? 4'b0010 : 4'b0011;
															assign node62155 = (inp[8]) ? node62159 : node62156;
																assign node62156 = (inp[7]) ? 4'b0011 : 4'b0010;
																assign node62159 = (inp[7]) ? 4'b0010 : 4'b0011;
												assign node62162 = (inp[12]) ? node62184 : node62163;
													assign node62163 = (inp[10]) ? node62177 : node62164;
														assign node62164 = (inp[7]) ? node62172 : node62165;
															assign node62165 = (inp[8]) ? node62169 : node62166;
																assign node62166 = (inp[2]) ? 4'b0010 : 4'b0011;
																assign node62169 = (inp[2]) ? 4'b0011 : 4'b0010;
															assign node62172 = (inp[8]) ? node62174 : 4'b0011;
																assign node62174 = (inp[2]) ? 4'b0010 : 4'b0011;
														assign node62177 = (inp[2]) ? node62179 : 4'b0110;
															assign node62179 = (inp[7]) ? node62181 : 4'b0111;
																assign node62181 = (inp[8]) ? 4'b0110 : 4'b0111;
													assign node62184 = (inp[8]) ? node62190 : node62185;
														assign node62185 = (inp[7]) ? 4'b0111 : node62186;
															assign node62186 = (inp[2]) ? 4'b0110 : 4'b0111;
														assign node62190 = (inp[10]) ? node62198 : node62191;
															assign node62191 = (inp[2]) ? node62195 : node62192;
																assign node62192 = (inp[7]) ? 4'b0111 : 4'b0110;
																assign node62195 = (inp[7]) ? 4'b0110 : 4'b0111;
															assign node62198 = (inp[2]) ? 4'b0110 : node62199;
																assign node62199 = (inp[7]) ? 4'b0111 : 4'b0110;
											assign node62203 = (inp[9]) ? node62245 : node62204;
												assign node62204 = (inp[10]) ? node62228 : node62205;
													assign node62205 = (inp[12]) ? node62215 : node62206;
														assign node62206 = (inp[8]) ? node62208 : 4'b0010;
															assign node62208 = (inp[7]) ? node62212 : node62209;
																assign node62209 = (inp[2]) ? 4'b0011 : 4'b0010;
																assign node62212 = (inp[2]) ? 4'b0010 : 4'b0011;
														assign node62215 = (inp[7]) ? node62221 : node62216;
															assign node62216 = (inp[8]) ? 4'b0110 : node62217;
																assign node62217 = (inp[2]) ? 4'b0110 : 4'b0111;
															assign node62221 = (inp[8]) ? node62225 : node62222;
																assign node62222 = (inp[2]) ? 4'b0111 : 4'b0110;
																assign node62225 = (inp[2]) ? 4'b0110 : 4'b0111;
													assign node62228 = (inp[8]) ? node62240 : node62229;
														assign node62229 = (inp[12]) ? node62235 : node62230;
															assign node62230 = (inp[7]) ? 4'b0111 : node62231;
																assign node62231 = (inp[2]) ? 4'b0110 : 4'b0111;
															assign node62235 = (inp[2]) ? node62237 : 4'b0110;
																assign node62237 = (inp[7]) ? 4'b0111 : 4'b0110;
														assign node62240 = (inp[2]) ? node62242 : 4'b0111;
															assign node62242 = (inp[7]) ? 4'b0110 : 4'b0111;
												assign node62245 = (inp[12]) ? node62261 : node62246;
													assign node62246 = (inp[10]) ? node62256 : node62247;
														assign node62247 = (inp[7]) ? 4'b0110 : node62248;
															assign node62248 = (inp[8]) ? node62252 : node62249;
																assign node62249 = (inp[2]) ? 4'b0110 : 4'b0111;
																assign node62252 = (inp[2]) ? 4'b0111 : 4'b0110;
														assign node62256 = (inp[8]) ? 4'b0011 : node62257;
															assign node62257 = (inp[7]) ? 4'b0010 : 4'b0011;
													assign node62261 = (inp[10]) ? node62273 : node62262;
														assign node62262 = (inp[7]) ? node62268 : node62263;
															assign node62263 = (inp[8]) ? 4'b0010 : node62264;
																assign node62264 = (inp[2]) ? 4'b0010 : 4'b0011;
															assign node62268 = (inp[8]) ? 4'b0011 : node62269;
																assign node62269 = (inp[2]) ? 4'b0011 : 4'b0010;
														assign node62273 = (inp[8]) ? node62275 : 4'b0010;
															assign node62275 = (inp[2]) ? node62279 : node62276;
																assign node62276 = (inp[7]) ? 4'b0011 : 4'b0010;
																assign node62279 = (inp[7]) ? 4'b0010 : 4'b0011;
										assign node62282 = (inp[9]) ? node62360 : node62283;
											assign node62283 = (inp[4]) ? node62325 : node62284;
												assign node62284 = (inp[10]) ? node62300 : node62285;
													assign node62285 = (inp[12]) ? node62295 : node62286;
														assign node62286 = (inp[7]) ? 4'b0110 : node62287;
															assign node62287 = (inp[2]) ? node62291 : node62288;
																assign node62288 = (inp[8]) ? 4'b0110 : 4'b0111;
																assign node62291 = (inp[8]) ? 4'b0111 : 4'b0110;
														assign node62295 = (inp[2]) ? 4'b0010 : node62296;
															assign node62296 = (inp[7]) ? 4'b0010 : 4'b0011;
													assign node62300 = (inp[7]) ? node62316 : node62301;
														assign node62301 = (inp[12]) ? node62309 : node62302;
															assign node62302 = (inp[2]) ? node62306 : node62303;
																assign node62303 = (inp[8]) ? 4'b0010 : 4'b0011;
																assign node62306 = (inp[8]) ? 4'b0011 : 4'b0010;
															assign node62309 = (inp[2]) ? node62313 : node62310;
																assign node62310 = (inp[8]) ? 4'b0010 : 4'b0011;
																assign node62313 = (inp[8]) ? 4'b0011 : 4'b0010;
														assign node62316 = (inp[12]) ? 4'b0011 : node62317;
															assign node62317 = (inp[8]) ? node62321 : node62318;
																assign node62318 = (inp[2]) ? 4'b0011 : 4'b0010;
																assign node62321 = (inp[2]) ? 4'b0010 : 4'b0011;
												assign node62325 = (inp[12]) ? node62347 : node62326;
													assign node62326 = (inp[10]) ? node62340 : node62327;
														assign node62327 = (inp[2]) ? node62333 : node62328;
															assign node62328 = (inp[7]) ? 4'b0010 : node62329;
																assign node62329 = (inp[8]) ? 4'b0010 : 4'b0011;
															assign node62333 = (inp[7]) ? node62337 : node62334;
																assign node62334 = (inp[8]) ? 4'b0011 : 4'b0010;
																assign node62337 = (inp[8]) ? 4'b0010 : 4'b0011;
														assign node62340 = (inp[7]) ? 4'b0101 : node62341;
															assign node62341 = (inp[2]) ? node62343 : 4'b0100;
																assign node62343 = (inp[8]) ? 4'b0101 : 4'b0100;
													assign node62347 = (inp[7]) ? node62353 : node62348;
														assign node62348 = (inp[2]) ? 4'b0101 : node62349;
															assign node62349 = (inp[8]) ? 4'b0100 : 4'b0101;
														assign node62353 = (inp[8]) ? node62357 : node62354;
															assign node62354 = (inp[2]) ? 4'b0101 : 4'b0100;
															assign node62357 = (inp[2]) ? 4'b0100 : 4'b0101;
											assign node62360 = (inp[4]) ? node62392 : node62361;
												assign node62361 = (inp[12]) ? node62379 : node62362;
													assign node62362 = (inp[10]) ? node62372 : node62363;
														assign node62363 = (inp[8]) ? 4'b0011 : node62364;
															assign node62364 = (inp[7]) ? node62368 : node62365;
																assign node62365 = (inp[2]) ? 4'b0010 : 4'b0011;
																assign node62368 = (inp[2]) ? 4'b0011 : 4'b0010;
														assign node62372 = (inp[2]) ? 4'b0100 : node62373;
															assign node62373 = (inp[8]) ? 4'b0100 : node62374;
																assign node62374 = (inp[7]) ? 4'b0100 : 4'b0101;
													assign node62379 = (inp[8]) ? node62387 : node62380;
														assign node62380 = (inp[2]) ? node62384 : node62381;
															assign node62381 = (inp[7]) ? 4'b0100 : 4'b0101;
															assign node62384 = (inp[7]) ? 4'b0101 : 4'b0100;
														assign node62387 = (inp[2]) ? 4'b0101 : node62388;
															assign node62388 = (inp[7]) ? 4'b0101 : 4'b0100;
												assign node62392 = (inp[12]) ? node62406 : node62393;
													assign node62393 = (inp[10]) ? node62401 : node62394;
														assign node62394 = (inp[8]) ? node62396 : 4'b0101;
															assign node62396 = (inp[7]) ? node62398 : 4'b0100;
																assign node62398 = (inp[2]) ? 4'b0100 : 4'b0101;
														assign node62401 = (inp[7]) ? 4'b0000 : node62402;
															assign node62402 = (inp[8]) ? 4'b0000 : 4'b0001;
													assign node62406 = (inp[7]) ? node62414 : node62407;
														assign node62407 = (inp[2]) ? node62411 : node62408;
															assign node62408 = (inp[8]) ? 4'b0000 : 4'b0001;
															assign node62411 = (inp[8]) ? 4'b0001 : 4'b0000;
														assign node62414 = (inp[8]) ? node62418 : node62415;
															assign node62415 = (inp[2]) ? 4'b0001 : 4'b0000;
															assign node62418 = (inp[2]) ? 4'b0000 : 4'b0001;
									assign node62421 = (inp[5]) ? node62611 : node62422;
										assign node62422 = (inp[4]) ? node62528 : node62423;
											assign node62423 = (inp[9]) ? node62481 : node62424;
												assign node62424 = (inp[10]) ? node62452 : node62425;
													assign node62425 = (inp[12]) ? node62439 : node62426;
														assign node62426 = (inp[2]) ? node62434 : node62427;
															assign node62427 = (inp[8]) ? node62431 : node62428;
																assign node62428 = (inp[7]) ? 4'b0110 : 4'b0111;
																assign node62431 = (inp[7]) ? 4'b0111 : 4'b0110;
															assign node62434 = (inp[7]) ? node62436 : 4'b0110;
																assign node62436 = (inp[8]) ? 4'b0110 : 4'b0111;
														assign node62439 = (inp[7]) ? node62447 : node62440;
															assign node62440 = (inp[2]) ? node62444 : node62441;
																assign node62441 = (inp[8]) ? 4'b0010 : 4'b0011;
																assign node62444 = (inp[8]) ? 4'b0011 : 4'b0010;
															assign node62447 = (inp[2]) ? node62449 : 4'b0010;
																assign node62449 = (inp[8]) ? 4'b0010 : 4'b0011;
													assign node62452 = (inp[12]) ? node62468 : node62453;
														assign node62453 = (inp[2]) ? node62461 : node62454;
															assign node62454 = (inp[8]) ? node62458 : node62455;
																assign node62455 = (inp[7]) ? 4'b0010 : 4'b0011;
																assign node62458 = (inp[7]) ? 4'b0011 : 4'b0010;
															assign node62461 = (inp[8]) ? node62465 : node62462;
																assign node62462 = (inp[7]) ? 4'b0011 : 4'b0010;
																assign node62465 = (inp[7]) ? 4'b0010 : 4'b0011;
														assign node62468 = (inp[2]) ? node62476 : node62469;
															assign node62469 = (inp[8]) ? node62473 : node62470;
																assign node62470 = (inp[7]) ? 4'b0010 : 4'b0011;
																assign node62473 = (inp[7]) ? 4'b0011 : 4'b0010;
															assign node62476 = (inp[7]) ? 4'b0011 : node62477;
																assign node62477 = (inp[8]) ? 4'b0011 : 4'b0010;
												assign node62481 = (inp[10]) ? node62507 : node62482;
													assign node62482 = (inp[12]) ? node62496 : node62483;
														assign node62483 = (inp[2]) ? node62489 : node62484;
															assign node62484 = (inp[7]) ? 4'b0011 : node62485;
																assign node62485 = (inp[8]) ? 4'b0010 : 4'b0011;
															assign node62489 = (inp[7]) ? node62493 : node62490;
																assign node62490 = (inp[8]) ? 4'b0011 : 4'b0010;
																assign node62493 = (inp[8]) ? 4'b0010 : 4'b0011;
														assign node62496 = (inp[7]) ? node62502 : node62497;
															assign node62497 = (inp[8]) ? 4'b0100 : node62498;
																assign node62498 = (inp[2]) ? 4'b0100 : 4'b0101;
															assign node62502 = (inp[2]) ? 4'b0101 : node62503;
																assign node62503 = (inp[8]) ? 4'b0101 : 4'b0100;
													assign node62507 = (inp[8]) ? node62517 : node62508;
														assign node62508 = (inp[12]) ? 4'b0100 : node62509;
															assign node62509 = (inp[2]) ? node62513 : node62510;
																assign node62510 = (inp[7]) ? 4'b0100 : 4'b0101;
																assign node62513 = (inp[7]) ? 4'b0101 : 4'b0100;
														assign node62517 = (inp[12]) ? node62523 : node62518;
															assign node62518 = (inp[7]) ? node62520 : 4'b0100;
																assign node62520 = (inp[2]) ? 4'b0100 : 4'b0101;
															assign node62523 = (inp[7]) ? node62525 : 4'b0101;
																assign node62525 = (inp[2]) ? 4'b0100 : 4'b0101;
											assign node62528 = (inp[9]) ? node62574 : node62529;
												assign node62529 = (inp[10]) ? node62557 : node62530;
													assign node62530 = (inp[12]) ? node62544 : node62531;
														assign node62531 = (inp[7]) ? node62537 : node62532;
															assign node62532 = (inp[2]) ? node62534 : 4'b0011;
																assign node62534 = (inp[8]) ? 4'b0011 : 4'b0010;
															assign node62537 = (inp[8]) ? node62541 : node62538;
																assign node62538 = (inp[2]) ? 4'b0011 : 4'b0010;
																assign node62541 = (inp[2]) ? 4'b0010 : 4'b0011;
														assign node62544 = (inp[7]) ? node62552 : node62545;
															assign node62545 = (inp[2]) ? node62549 : node62546;
																assign node62546 = (inp[8]) ? 4'b0100 : 4'b0101;
																assign node62549 = (inp[8]) ? 4'b0101 : 4'b0100;
															assign node62552 = (inp[2]) ? 4'b0101 : node62553;
																assign node62553 = (inp[8]) ? 4'b0101 : 4'b0100;
													assign node62557 = (inp[7]) ? node62567 : node62558;
														assign node62558 = (inp[12]) ? 4'b0100 : node62559;
															assign node62559 = (inp[2]) ? node62563 : node62560;
																assign node62560 = (inp[8]) ? 4'b0100 : 4'b0101;
																assign node62563 = (inp[8]) ? 4'b0101 : 4'b0100;
														assign node62567 = (inp[8]) ? node62571 : node62568;
															assign node62568 = (inp[2]) ? 4'b0101 : 4'b0100;
															assign node62571 = (inp[2]) ? 4'b0100 : 4'b0101;
												assign node62574 = (inp[10]) ? node62596 : node62575;
													assign node62575 = (inp[12]) ? node62583 : node62576;
														assign node62576 = (inp[8]) ? 4'b0100 : node62577;
															assign node62577 = (inp[7]) ? 4'b0100 : node62578;
																assign node62578 = (inp[2]) ? 4'b0100 : 4'b0101;
														assign node62583 = (inp[2]) ? node62591 : node62584;
															assign node62584 = (inp[8]) ? node62588 : node62585;
																assign node62585 = (inp[7]) ? 4'b0000 : 4'b0001;
																assign node62588 = (inp[7]) ? 4'b0001 : 4'b0000;
															assign node62591 = (inp[7]) ? 4'b0000 : node62592;
																assign node62592 = (inp[8]) ? 4'b0001 : 4'b0000;
													assign node62596 = (inp[2]) ? node62604 : node62597;
														assign node62597 = (inp[7]) ? node62601 : node62598;
															assign node62598 = (inp[8]) ? 4'b0000 : 4'b0001;
															assign node62601 = (inp[8]) ? 4'b0001 : 4'b0000;
														assign node62604 = (inp[8]) ? node62608 : node62605;
															assign node62605 = (inp[7]) ? 4'b0001 : 4'b0000;
															assign node62608 = (inp[7]) ? 4'b0000 : 4'b0001;
										assign node62611 = (inp[8]) ? node62695 : node62612;
											assign node62612 = (inp[7]) ? node62656 : node62613;
												assign node62613 = (inp[2]) ? node62635 : node62614;
													assign node62614 = (inp[4]) ? node62624 : node62615;
														assign node62615 = (inp[10]) ? 4'b0001 : node62616;
															assign node62616 = (inp[9]) ? node62620 : node62617;
																assign node62617 = (inp[12]) ? 4'b0001 : 4'b0101;
																assign node62620 = (inp[12]) ? 4'b0101 : 4'b0001;
														assign node62624 = (inp[9]) ? node62630 : node62625;
															assign node62625 = (inp[12]) ? 4'b0101 : node62626;
																assign node62626 = (inp[10]) ? 4'b0101 : 4'b0001;
															assign node62630 = (inp[12]) ? 4'b0001 : node62631;
																assign node62631 = (inp[10]) ? 4'b0001 : 4'b0101;
													assign node62635 = (inp[10]) ? node62651 : node62636;
														assign node62636 = (inp[12]) ? node62644 : node62637;
															assign node62637 = (inp[9]) ? node62641 : node62638;
																assign node62638 = (inp[4]) ? 4'b0000 : 4'b0100;
																assign node62641 = (inp[4]) ? 4'b0100 : 4'b0000;
															assign node62644 = (inp[9]) ? node62648 : node62645;
																assign node62645 = (inp[4]) ? 4'b0100 : 4'b0000;
																assign node62648 = (inp[4]) ? 4'b0000 : 4'b0100;
														assign node62651 = (inp[9]) ? node62653 : 4'b0000;
															assign node62653 = (inp[4]) ? 4'b0000 : 4'b0100;
												assign node62656 = (inp[2]) ? node62678 : node62657;
													assign node62657 = (inp[10]) ? node62671 : node62658;
														assign node62658 = (inp[12]) ? node62664 : node62659;
															assign node62659 = (inp[9]) ? 4'b0000 : node62660;
																assign node62660 = (inp[4]) ? 4'b0000 : 4'b0100;
															assign node62664 = (inp[9]) ? node62668 : node62665;
																assign node62665 = (inp[4]) ? 4'b0100 : 4'b0000;
																assign node62668 = (inp[4]) ? 4'b0000 : 4'b0100;
														assign node62671 = (inp[4]) ? node62675 : node62672;
															assign node62672 = (inp[9]) ? 4'b0100 : 4'b0000;
															assign node62675 = (inp[9]) ? 4'b0000 : 4'b0100;
													assign node62678 = (inp[12]) ? node62690 : node62679;
														assign node62679 = (inp[9]) ? node62685 : node62680;
															assign node62680 = (inp[4]) ? 4'b0101 : node62681;
																assign node62681 = (inp[10]) ? 4'b0001 : 4'b0101;
															assign node62685 = (inp[10]) ? node62687 : 4'b0001;
																assign node62687 = (inp[4]) ? 4'b0001 : 4'b0101;
														assign node62690 = (inp[10]) ? node62692 : 4'b0001;
															assign node62692 = (inp[4]) ? 4'b0001 : 4'b0101;
											assign node62695 = (inp[9]) ? node62739 : node62696;
												assign node62696 = (inp[4]) ? node62712 : node62697;
													assign node62697 = (inp[10]) ? node62705 : node62698;
														assign node62698 = (inp[12]) ? node62700 : 4'b0101;
															assign node62700 = (inp[7]) ? 4'b0000 : node62701;
																assign node62701 = (inp[2]) ? 4'b0001 : 4'b0000;
														assign node62705 = (inp[7]) ? node62709 : node62706;
															assign node62706 = (inp[2]) ? 4'b0001 : 4'b0000;
															assign node62709 = (inp[2]) ? 4'b0000 : 4'b0001;
													assign node62712 = (inp[12]) ? node62726 : node62713;
														assign node62713 = (inp[10]) ? node62719 : node62714;
															assign node62714 = (inp[7]) ? 4'b0000 : node62715;
																assign node62715 = (inp[2]) ? 4'b0001 : 4'b0000;
															assign node62719 = (inp[7]) ? node62723 : node62720;
																assign node62720 = (inp[2]) ? 4'b0101 : 4'b0100;
																assign node62723 = (inp[2]) ? 4'b0100 : 4'b0101;
														assign node62726 = (inp[10]) ? node62734 : node62727;
															assign node62727 = (inp[2]) ? node62731 : node62728;
																assign node62728 = (inp[7]) ? 4'b0101 : 4'b0100;
																assign node62731 = (inp[7]) ? 4'b0100 : 4'b0101;
															assign node62734 = (inp[2]) ? node62736 : 4'b0100;
																assign node62736 = (inp[7]) ? 4'b0100 : 4'b0101;
												assign node62739 = (inp[4]) ? node62757 : node62740;
													assign node62740 = (inp[10]) ? node62750 : node62741;
														assign node62741 = (inp[12]) ? node62743 : 4'b0000;
															assign node62743 = (inp[7]) ? node62747 : node62744;
																assign node62744 = (inp[2]) ? 4'b0101 : 4'b0100;
																assign node62747 = (inp[2]) ? 4'b0100 : 4'b0101;
														assign node62750 = (inp[2]) ? node62754 : node62751;
															assign node62751 = (inp[7]) ? 4'b0101 : 4'b0100;
															assign node62754 = (inp[7]) ? 4'b0100 : 4'b0101;
													assign node62757 = (inp[10]) ? node62761 : node62758;
														assign node62758 = (inp[12]) ? 4'b0000 : 4'b0101;
														assign node62761 = (inp[12]) ? node62767 : node62762;
															assign node62762 = (inp[7]) ? 4'b0000 : node62763;
																assign node62763 = (inp[2]) ? 4'b0001 : 4'b0000;
															assign node62767 = (inp[2]) ? node62769 : 4'b0001;
																assign node62769 = (inp[7]) ? 4'b0000 : 4'b0001;
								assign node62772 = (inp[5]) ? node63106 : node62773;
									assign node62773 = (inp[3]) ? node62949 : node62774;
										assign node62774 = (inp[10]) ? node62872 : node62775;
											assign node62775 = (inp[8]) ? node62827 : node62776;
												assign node62776 = (inp[12]) ? node62798 : node62777;
													assign node62777 = (inp[9]) ? node62787 : node62778;
														assign node62778 = (inp[4]) ? node62780 : 4'b0100;
															assign node62780 = (inp[7]) ? node62784 : node62781;
																assign node62781 = (inp[2]) ? 4'b0000 : 4'b0001;
																assign node62784 = (inp[2]) ? 4'b0001 : 4'b0000;
														assign node62787 = (inp[4]) ? node62793 : node62788;
															assign node62788 = (inp[2]) ? node62790 : 4'b0000;
																assign node62790 = (inp[7]) ? 4'b0001 : 4'b0000;
															assign node62793 = (inp[2]) ? 4'b0100 : node62794;
																assign node62794 = (inp[7]) ? 4'b0100 : 4'b0101;
													assign node62798 = (inp[4]) ? node62814 : node62799;
														assign node62799 = (inp[9]) ? node62807 : node62800;
															assign node62800 = (inp[7]) ? node62804 : node62801;
																assign node62801 = (inp[2]) ? 4'b0000 : 4'b0001;
																assign node62804 = (inp[2]) ? 4'b0001 : 4'b0000;
															assign node62807 = (inp[2]) ? node62811 : node62808;
																assign node62808 = (inp[7]) ? 4'b0100 : 4'b0101;
																assign node62811 = (inp[7]) ? 4'b0101 : 4'b0100;
														assign node62814 = (inp[9]) ? node62820 : node62815;
															assign node62815 = (inp[7]) ? 4'b0101 : node62816;
																assign node62816 = (inp[2]) ? 4'b0100 : 4'b0101;
															assign node62820 = (inp[7]) ? node62824 : node62821;
																assign node62821 = (inp[2]) ? 4'b0000 : 4'b0001;
																assign node62824 = (inp[2]) ? 4'b0001 : 4'b0000;
												assign node62827 = (inp[4]) ? node62845 : node62828;
													assign node62828 = (inp[9]) ? node62836 : node62829;
														assign node62829 = (inp[12]) ? 4'b0001 : node62830;
															assign node62830 = (inp[7]) ? node62832 : 4'b0101;
																assign node62832 = (inp[2]) ? 4'b0100 : 4'b0101;
														assign node62836 = (inp[12]) ? node62842 : node62837;
															assign node62837 = (inp[7]) ? node62839 : 4'b0001;
																assign node62839 = (inp[2]) ? 4'b0000 : 4'b0001;
															assign node62842 = (inp[7]) ? 4'b0101 : 4'b0100;
													assign node62845 = (inp[2]) ? node62857 : node62846;
														assign node62846 = (inp[7]) ? node62852 : node62847;
															assign node62847 = (inp[9]) ? 4'b0000 : node62848;
																assign node62848 = (inp[12]) ? 4'b0100 : 4'b0000;
															assign node62852 = (inp[9]) ? node62854 : 4'b0001;
																assign node62854 = (inp[12]) ? 4'b0001 : 4'b0101;
														assign node62857 = (inp[7]) ? node62865 : node62858;
															assign node62858 = (inp[12]) ? node62862 : node62859;
																assign node62859 = (inp[9]) ? 4'b0101 : 4'b0001;
																assign node62862 = (inp[9]) ? 4'b0001 : 4'b0101;
															assign node62865 = (inp[12]) ? node62869 : node62866;
																assign node62866 = (inp[9]) ? 4'b0100 : 4'b0000;
																assign node62869 = (inp[9]) ? 4'b0000 : 4'b0100;
											assign node62872 = (inp[4]) ? node62918 : node62873;
												assign node62873 = (inp[9]) ? node62889 : node62874;
													assign node62874 = (inp[7]) ? node62882 : node62875;
														assign node62875 = (inp[8]) ? node62879 : node62876;
															assign node62876 = (inp[2]) ? 4'b0000 : 4'b0001;
															assign node62879 = (inp[2]) ? 4'b0001 : 4'b0000;
														assign node62882 = (inp[2]) ? node62886 : node62883;
															assign node62883 = (inp[8]) ? 4'b0001 : 4'b0000;
															assign node62886 = (inp[8]) ? 4'b0000 : 4'b0001;
													assign node62889 = (inp[8]) ? node62903 : node62890;
														assign node62890 = (inp[12]) ? node62898 : node62891;
															assign node62891 = (inp[2]) ? node62895 : node62892;
																assign node62892 = (inp[7]) ? 4'b0100 : 4'b0101;
																assign node62895 = (inp[7]) ? 4'b0101 : 4'b0100;
															assign node62898 = (inp[2]) ? node62900 : 4'b0101;
																assign node62900 = (inp[7]) ? 4'b0101 : 4'b0100;
														assign node62903 = (inp[12]) ? node62911 : node62904;
															assign node62904 = (inp[7]) ? node62908 : node62905;
																assign node62905 = (inp[2]) ? 4'b0101 : 4'b0100;
																assign node62908 = (inp[2]) ? 4'b0100 : 4'b0101;
															assign node62911 = (inp[2]) ? node62915 : node62912;
																assign node62912 = (inp[7]) ? 4'b0101 : 4'b0100;
																assign node62915 = (inp[7]) ? 4'b0100 : 4'b0101;
												assign node62918 = (inp[9]) ? node62936 : node62919;
													assign node62919 = (inp[7]) ? node62927 : node62920;
														assign node62920 = (inp[8]) ? node62924 : node62921;
															assign node62921 = (inp[2]) ? 4'b0100 : 4'b0101;
															assign node62924 = (inp[2]) ? 4'b0101 : 4'b0100;
														assign node62927 = (inp[12]) ? 4'b0101 : node62928;
															assign node62928 = (inp[2]) ? node62932 : node62929;
																assign node62929 = (inp[8]) ? 4'b0101 : 4'b0100;
																assign node62932 = (inp[8]) ? 4'b0100 : 4'b0101;
													assign node62936 = (inp[12]) ? node62938 : 4'b0001;
														assign node62938 = (inp[8]) ? node62944 : node62939;
															assign node62939 = (inp[2]) ? node62941 : 4'b0000;
																assign node62941 = (inp[7]) ? 4'b0001 : 4'b0000;
															assign node62944 = (inp[7]) ? 4'b0001 : node62945;
																assign node62945 = (inp[2]) ? 4'b0001 : 4'b0000;
										assign node62949 = (inp[9]) ? node63019 : node62950;
											assign node62950 = (inp[4]) ? node62990 : node62951;
												assign node62951 = (inp[10]) ? node62975 : node62952;
													assign node62952 = (inp[12]) ? node62964 : node62953;
														assign node62953 = (inp[7]) ? node62959 : node62954;
															assign node62954 = (inp[8]) ? node62956 : 4'b0101;
																assign node62956 = (inp[2]) ? 4'b0101 : 4'b0100;
															assign node62959 = (inp[8]) ? 4'b0100 : node62960;
																assign node62960 = (inp[2]) ? 4'b0101 : 4'b0100;
														assign node62964 = (inp[8]) ? node62970 : node62965;
															assign node62965 = (inp[2]) ? node62967 : 4'b0001;
																assign node62967 = (inp[7]) ? 4'b0001 : 4'b0000;
															assign node62970 = (inp[7]) ? 4'b0000 : node62971;
																assign node62971 = (inp[2]) ? 4'b0001 : 4'b0000;
													assign node62975 = (inp[8]) ? node62983 : node62976;
														assign node62976 = (inp[7]) ? node62980 : node62977;
															assign node62977 = (inp[2]) ? 4'b0000 : 4'b0001;
															assign node62980 = (inp[2]) ? 4'b0001 : 4'b0000;
														assign node62983 = (inp[7]) ? node62987 : node62984;
															assign node62984 = (inp[2]) ? 4'b0001 : 4'b0000;
															assign node62987 = (inp[2]) ? 4'b0000 : 4'b0001;
												assign node62990 = (inp[10]) ? node63006 : node62991;
													assign node62991 = (inp[12]) ? node63003 : node62992;
														assign node62992 = (inp[2]) ? node62998 : node62993;
															assign node62993 = (inp[8]) ? 4'b0000 : node62994;
																assign node62994 = (inp[7]) ? 4'b0000 : 4'b0001;
															assign node62998 = (inp[7]) ? 4'b0001 : node62999;
																assign node62999 = (inp[8]) ? 4'b0001 : 4'b0000;
														assign node63003 = (inp[7]) ? 4'b0111 : 4'b0110;
													assign node63006 = (inp[7]) ? node63014 : node63007;
														assign node63007 = (inp[2]) ? node63011 : node63008;
															assign node63008 = (inp[8]) ? 4'b0110 : 4'b0111;
															assign node63011 = (inp[8]) ? 4'b0111 : 4'b0110;
														assign node63014 = (inp[2]) ? node63016 : 4'b0111;
															assign node63016 = (inp[8]) ? 4'b0110 : 4'b0111;
											assign node63019 = (inp[4]) ? node63059 : node63020;
												assign node63020 = (inp[12]) ? node63040 : node63021;
													assign node63021 = (inp[10]) ? node63035 : node63022;
														assign node63022 = (inp[7]) ? node63028 : node63023;
															assign node63023 = (inp[8]) ? node63025 : 4'b0000;
																assign node63025 = (inp[2]) ? 4'b0001 : 4'b0000;
															assign node63028 = (inp[2]) ? node63032 : node63029;
																assign node63029 = (inp[8]) ? 4'b0001 : 4'b0000;
																assign node63032 = (inp[8]) ? 4'b0000 : 4'b0001;
														assign node63035 = (inp[2]) ? node63037 : 4'b0111;
															assign node63037 = (inp[8]) ? 4'b0110 : 4'b0111;
													assign node63040 = (inp[8]) ? node63054 : node63041;
														assign node63041 = (inp[10]) ? node63047 : node63042;
															assign node63042 = (inp[7]) ? 4'b0111 : node63043;
																assign node63043 = (inp[2]) ? 4'b0110 : 4'b0111;
															assign node63047 = (inp[7]) ? node63051 : node63048;
																assign node63048 = (inp[2]) ? 4'b0110 : 4'b0111;
																assign node63051 = (inp[2]) ? 4'b0111 : 4'b0110;
														assign node63054 = (inp[2]) ? 4'b0110 : node63055;
															assign node63055 = (inp[7]) ? 4'b0111 : 4'b0110;
												assign node63059 = (inp[12]) ? node63083 : node63060;
													assign node63060 = (inp[10]) ? node63070 : node63061;
														assign node63061 = (inp[8]) ? node63063 : 4'b0110;
															assign node63063 = (inp[7]) ? node63067 : node63064;
																assign node63064 = (inp[2]) ? 4'b0111 : 4'b0110;
																assign node63067 = (inp[2]) ? 4'b0110 : 4'b0111;
														assign node63070 = (inp[7]) ? node63076 : node63071;
															assign node63071 = (inp[8]) ? node63073 : 4'b0010;
																assign node63073 = (inp[2]) ? 4'b0011 : 4'b0010;
															assign node63076 = (inp[2]) ? node63080 : node63077;
																assign node63077 = (inp[8]) ? 4'b0011 : 4'b0010;
																assign node63080 = (inp[8]) ? 4'b0010 : 4'b0011;
													assign node63083 = (inp[10]) ? node63097 : node63084;
														assign node63084 = (inp[8]) ? node63090 : node63085;
															assign node63085 = (inp[2]) ? node63087 : 4'b0011;
																assign node63087 = (inp[7]) ? 4'b0011 : 4'b0010;
															assign node63090 = (inp[2]) ? node63094 : node63091;
																assign node63091 = (inp[7]) ? 4'b0011 : 4'b0010;
																assign node63094 = (inp[7]) ? 4'b0010 : 4'b0011;
														assign node63097 = (inp[7]) ? 4'b0010 : node63098;
															assign node63098 = (inp[8]) ? node63102 : node63099;
																assign node63099 = (inp[2]) ? 4'b0010 : 4'b0011;
																assign node63102 = (inp[2]) ? 4'b0011 : 4'b0010;
									assign node63106 = (inp[3]) ? node63264 : node63107;
										assign node63107 = (inp[9]) ? node63181 : node63108;
											assign node63108 = (inp[4]) ? node63152 : node63109;
												assign node63109 = (inp[12]) ? node63133 : node63110;
													assign node63110 = (inp[10]) ? node63118 : node63111;
														assign node63111 = (inp[8]) ? 4'b0100 : node63112;
															assign node63112 = (inp[7]) ? node63114 : 4'b0100;
																assign node63114 = (inp[2]) ? 4'b0101 : 4'b0100;
														assign node63118 = (inp[7]) ? node63126 : node63119;
															assign node63119 = (inp[2]) ? node63123 : node63120;
																assign node63120 = (inp[8]) ? 4'b0000 : 4'b0001;
																assign node63123 = (inp[8]) ? 4'b0001 : 4'b0000;
															assign node63126 = (inp[8]) ? node63130 : node63127;
																assign node63127 = (inp[2]) ? 4'b0001 : 4'b0000;
																assign node63130 = (inp[2]) ? 4'b0000 : 4'b0001;
													assign node63133 = (inp[10]) ? node63147 : node63134;
														assign node63134 = (inp[2]) ? node63142 : node63135;
															assign node63135 = (inp[7]) ? node63139 : node63136;
																assign node63136 = (inp[8]) ? 4'b0000 : 4'b0001;
																assign node63139 = (inp[8]) ? 4'b0001 : 4'b0000;
															assign node63142 = (inp[8]) ? 4'b0001 : node63143;
																assign node63143 = (inp[7]) ? 4'b0001 : 4'b0000;
														assign node63147 = (inp[7]) ? node63149 : 4'b0001;
															assign node63149 = (inp[8]) ? 4'b0000 : 4'b0001;
												assign node63152 = (inp[12]) ? node63168 : node63153;
													assign node63153 = (inp[10]) ? node63163 : node63154;
														assign node63154 = (inp[7]) ? node63156 : 4'b0000;
															assign node63156 = (inp[8]) ? node63160 : node63157;
																assign node63157 = (inp[2]) ? 4'b0001 : 4'b0000;
																assign node63160 = (inp[2]) ? 4'b0000 : 4'b0001;
														assign node63163 = (inp[2]) ? node63165 : 4'b0110;
															assign node63165 = (inp[8]) ? 4'b0111 : 4'b0110;
													assign node63168 = (inp[2]) ? node63176 : node63169;
														assign node63169 = (inp[8]) ? node63173 : node63170;
															assign node63170 = (inp[7]) ? 4'b0110 : 4'b0111;
															assign node63173 = (inp[7]) ? 4'b0111 : 4'b0110;
														assign node63176 = (inp[7]) ? node63178 : 4'b0110;
															assign node63178 = (inp[8]) ? 4'b0110 : 4'b0111;
											assign node63181 = (inp[4]) ? node63223 : node63182;
												assign node63182 = (inp[12]) ? node63200 : node63183;
													assign node63183 = (inp[10]) ? node63193 : node63184;
														assign node63184 = (inp[8]) ? 4'b0000 : node63185;
															assign node63185 = (inp[7]) ? node63189 : node63186;
																assign node63186 = (inp[2]) ? 4'b0000 : 4'b0001;
																assign node63189 = (inp[2]) ? 4'b0001 : 4'b0000;
														assign node63193 = (inp[7]) ? node63195 : 4'b0110;
															assign node63195 = (inp[2]) ? 4'b0110 : node63196;
																assign node63196 = (inp[8]) ? 4'b0111 : 4'b0110;
													assign node63200 = (inp[8]) ? node63216 : node63201;
														assign node63201 = (inp[10]) ? node63209 : node63202;
															assign node63202 = (inp[7]) ? node63206 : node63203;
																assign node63203 = (inp[2]) ? 4'b0110 : 4'b0111;
																assign node63206 = (inp[2]) ? 4'b0111 : 4'b0110;
															assign node63209 = (inp[2]) ? node63213 : node63210;
																assign node63210 = (inp[7]) ? 4'b0110 : 4'b0111;
																assign node63213 = (inp[7]) ? 4'b0111 : 4'b0110;
														assign node63216 = (inp[2]) ? node63220 : node63217;
															assign node63217 = (inp[7]) ? 4'b0111 : 4'b0110;
															assign node63220 = (inp[7]) ? 4'b0110 : 4'b0111;
												assign node63223 = (inp[12]) ? node63247 : node63224;
													assign node63224 = (inp[10]) ? node63238 : node63225;
														assign node63225 = (inp[7]) ? node63233 : node63226;
															assign node63226 = (inp[8]) ? node63230 : node63227;
																assign node63227 = (inp[2]) ? 4'b0110 : 4'b0111;
																assign node63230 = (inp[2]) ? 4'b0111 : 4'b0110;
															assign node63233 = (inp[8]) ? node63235 : 4'b0110;
																assign node63235 = (inp[2]) ? 4'b0110 : 4'b0111;
														assign node63238 = (inp[2]) ? 4'b0010 : node63239;
															assign node63239 = (inp[7]) ? node63243 : node63240;
																assign node63240 = (inp[8]) ? 4'b0010 : 4'b0011;
																assign node63243 = (inp[8]) ? 4'b0011 : 4'b0010;
													assign node63247 = (inp[2]) ? node63255 : node63248;
														assign node63248 = (inp[7]) ? node63252 : node63249;
															assign node63249 = (inp[8]) ? 4'b0010 : 4'b0011;
															assign node63252 = (inp[8]) ? 4'b0011 : 4'b0010;
														assign node63255 = (inp[10]) ? node63261 : node63256;
															assign node63256 = (inp[7]) ? node63258 : 4'b0010;
																assign node63258 = (inp[8]) ? 4'b0010 : 4'b0011;
															assign node63261 = (inp[7]) ? 4'b0010 : 4'b0011;
										assign node63264 = (inp[9]) ? node63348 : node63265;
											assign node63265 = (inp[4]) ? node63303 : node63266;
												assign node63266 = (inp[12]) ? node63286 : node63267;
													assign node63267 = (inp[10]) ? node63277 : node63268;
														assign node63268 = (inp[2]) ? 4'b0110 : node63269;
															assign node63269 = (inp[8]) ? node63273 : node63270;
																assign node63270 = (inp[7]) ? 4'b0110 : 4'b0111;
																assign node63273 = (inp[7]) ? 4'b0111 : 4'b0110;
														assign node63277 = (inp[8]) ? node63279 : 4'b0010;
															assign node63279 = (inp[2]) ? node63283 : node63280;
																assign node63280 = (inp[7]) ? 4'b0011 : 4'b0010;
																assign node63283 = (inp[7]) ? 4'b0010 : 4'b0011;
													assign node63286 = (inp[10]) ? node63296 : node63287;
														assign node63287 = (inp[2]) ? node63289 : 4'b0011;
															assign node63289 = (inp[7]) ? node63293 : node63290;
																assign node63290 = (inp[8]) ? 4'b0011 : 4'b0010;
																assign node63293 = (inp[8]) ? 4'b0010 : 4'b0011;
														assign node63296 = (inp[8]) ? 4'b0010 : node63297;
															assign node63297 = (inp[7]) ? node63299 : 4'b0011;
																assign node63299 = (inp[2]) ? 4'b0011 : 4'b0010;
												assign node63303 = (inp[12]) ? node63327 : node63304;
													assign node63304 = (inp[10]) ? node63314 : node63305;
														assign node63305 = (inp[7]) ? 4'b0011 : node63306;
															assign node63306 = (inp[8]) ? node63310 : node63307;
																assign node63307 = (inp[2]) ? 4'b0010 : 4'b0011;
																assign node63310 = (inp[2]) ? 4'b0011 : 4'b0010;
														assign node63314 = (inp[7]) ? node63320 : node63315;
															assign node63315 = (inp[8]) ? node63317 : 4'b0111;
																assign node63317 = (inp[2]) ? 4'b0111 : 4'b0110;
															assign node63320 = (inp[2]) ? node63324 : node63321;
																assign node63321 = (inp[8]) ? 4'b0111 : 4'b0110;
																assign node63324 = (inp[8]) ? 4'b0110 : 4'b0111;
													assign node63327 = (inp[8]) ? node63335 : node63328;
														assign node63328 = (inp[7]) ? node63332 : node63329;
															assign node63329 = (inp[2]) ? 4'b0110 : 4'b0111;
															assign node63332 = (inp[2]) ? 4'b0111 : 4'b0110;
														assign node63335 = (inp[10]) ? node63341 : node63336;
															assign node63336 = (inp[2]) ? 4'b0110 : node63337;
																assign node63337 = (inp[7]) ? 4'b0111 : 4'b0110;
															assign node63341 = (inp[7]) ? node63345 : node63342;
																assign node63342 = (inp[2]) ? 4'b0111 : 4'b0110;
																assign node63345 = (inp[2]) ? 4'b0110 : 4'b0111;
											assign node63348 = (inp[4]) ? node63392 : node63349;
												assign node63349 = (inp[12]) ? node63375 : node63350;
													assign node63350 = (inp[10]) ? node63366 : node63351;
														assign node63351 = (inp[2]) ? node63359 : node63352;
															assign node63352 = (inp[7]) ? node63356 : node63353;
																assign node63353 = (inp[8]) ? 4'b0010 : 4'b0011;
																assign node63356 = (inp[8]) ? 4'b0011 : 4'b0010;
															assign node63359 = (inp[7]) ? node63363 : node63360;
																assign node63360 = (inp[8]) ? 4'b0011 : 4'b0010;
																assign node63363 = (inp[8]) ? 4'b0010 : 4'b0011;
														assign node63366 = (inp[2]) ? 4'b0110 : node63367;
															assign node63367 = (inp[8]) ? node63371 : node63368;
																assign node63368 = (inp[7]) ? 4'b0110 : 4'b0111;
																assign node63371 = (inp[7]) ? 4'b0111 : 4'b0110;
													assign node63375 = (inp[8]) ? node63383 : node63376;
														assign node63376 = (inp[2]) ? node63380 : node63377;
															assign node63377 = (inp[7]) ? 4'b0110 : 4'b0111;
															assign node63380 = (inp[7]) ? 4'b0111 : 4'b0110;
														assign node63383 = (inp[10]) ? 4'b0110 : node63384;
															assign node63384 = (inp[7]) ? node63388 : node63385;
																assign node63385 = (inp[2]) ? 4'b0111 : 4'b0110;
																assign node63388 = (inp[2]) ? 4'b0110 : 4'b0111;
												assign node63392 = (inp[12]) ? node63408 : node63393;
													assign node63393 = (inp[10]) ? node63401 : node63394;
														assign node63394 = (inp[8]) ? node63396 : 4'b0110;
															assign node63396 = (inp[2]) ? node63398 : 4'b0111;
																assign node63398 = (inp[7]) ? 4'b0110 : 4'b0111;
														assign node63401 = (inp[2]) ? 4'b0011 : node63402;
															assign node63402 = (inp[7]) ? node63404 : 4'b0010;
																assign node63404 = (inp[8]) ? 4'b0011 : 4'b0010;
													assign node63408 = (inp[8]) ? node63422 : node63409;
														assign node63409 = (inp[10]) ? node63417 : node63410;
															assign node63410 = (inp[7]) ? node63414 : node63411;
																assign node63411 = (inp[2]) ? 4'b0010 : 4'b0011;
																assign node63414 = (inp[2]) ? 4'b0011 : 4'b0010;
															assign node63417 = (inp[7]) ? 4'b0010 : node63418;
																assign node63418 = (inp[2]) ? 4'b0010 : 4'b0011;
														assign node63422 = (inp[7]) ? node63426 : node63423;
															assign node63423 = (inp[2]) ? 4'b0011 : 4'b0010;
															assign node63426 = (inp[2]) ? 4'b0010 : 4'b0011;
							assign node63429 = (inp[0]) ? node64111 : node63430;
								assign node63430 = (inp[5]) ? node63760 : node63431;
									assign node63431 = (inp[3]) ? node63591 : node63432;
										assign node63432 = (inp[7]) ? node63522 : node63433;
											assign node63433 = (inp[12]) ? node63469 : node63434;
												assign node63434 = (inp[8]) ? node63452 : node63435;
													assign node63435 = (inp[2]) ? node63439 : node63436;
														assign node63436 = (inp[4]) ? 4'b0101 : 4'b0001;
														assign node63439 = (inp[10]) ? node63445 : node63440;
															assign node63440 = (inp[9]) ? node63442 : 4'b0100;
																assign node63442 = (inp[4]) ? 4'b0100 : 4'b0000;
															assign node63445 = (inp[9]) ? node63449 : node63446;
																assign node63446 = (inp[4]) ? 4'b0100 : 4'b0000;
																assign node63449 = (inp[4]) ? 4'b0000 : 4'b0100;
													assign node63452 = (inp[2]) ? node63460 : node63453;
														assign node63453 = (inp[4]) ? 4'b0000 : node63454;
															assign node63454 = (inp[10]) ? node63456 : 4'b0100;
																assign node63456 = (inp[9]) ? 4'b0100 : 4'b0000;
														assign node63460 = (inp[9]) ? 4'b0101 : node63461;
															assign node63461 = (inp[10]) ? node63465 : node63462;
																assign node63462 = (inp[4]) ? 4'b0001 : 4'b0101;
																assign node63465 = (inp[4]) ? 4'b0101 : 4'b0001;
												assign node63469 = (inp[10]) ? node63495 : node63470;
													assign node63470 = (inp[2]) ? node63482 : node63471;
														assign node63471 = (inp[8]) ? node63477 : node63472;
															assign node63472 = (inp[9]) ? node63474 : 4'b0001;
																assign node63474 = (inp[4]) ? 4'b0001 : 4'b0101;
															assign node63477 = (inp[4]) ? 4'b0000 : node63478;
																assign node63478 = (inp[9]) ? 4'b0100 : 4'b0000;
														assign node63482 = (inp[8]) ? node63490 : node63483;
															assign node63483 = (inp[9]) ? node63487 : node63484;
																assign node63484 = (inp[4]) ? 4'b0100 : 4'b0000;
																assign node63487 = (inp[4]) ? 4'b0000 : 4'b0100;
															assign node63490 = (inp[4]) ? node63492 : 4'b0001;
																assign node63492 = (inp[9]) ? 4'b0001 : 4'b0101;
													assign node63495 = (inp[2]) ? node63511 : node63496;
														assign node63496 = (inp[8]) ? node63504 : node63497;
															assign node63497 = (inp[4]) ? node63501 : node63498;
																assign node63498 = (inp[9]) ? 4'b0101 : 4'b0001;
																assign node63501 = (inp[9]) ? 4'b0001 : 4'b0101;
															assign node63504 = (inp[4]) ? node63508 : node63505;
																assign node63505 = (inp[9]) ? 4'b0100 : 4'b0000;
																assign node63508 = (inp[9]) ? 4'b0000 : 4'b0100;
														assign node63511 = (inp[8]) ? node63517 : node63512;
															assign node63512 = (inp[9]) ? 4'b0000 : node63513;
																assign node63513 = (inp[4]) ? 4'b0100 : 4'b0000;
															assign node63517 = (inp[4]) ? node63519 : 4'b0001;
																assign node63519 = (inp[9]) ? 4'b0001 : 4'b0101;
											assign node63522 = (inp[4]) ? node63560 : node63523;
												assign node63523 = (inp[9]) ? node63545 : node63524;
													assign node63524 = (inp[12]) ? node63536 : node63525;
														assign node63525 = (inp[10]) ? node63533 : node63526;
															assign node63526 = (inp[2]) ? node63530 : node63527;
																assign node63527 = (inp[8]) ? 4'b0101 : 4'b0100;
																assign node63530 = (inp[8]) ? 4'b0100 : 4'b0101;
															assign node63533 = (inp[8]) ? 4'b0000 : 4'b0001;
														assign node63536 = (inp[10]) ? node63540 : node63537;
															assign node63537 = (inp[2]) ? 4'b0001 : 4'b0000;
															assign node63540 = (inp[8]) ? node63542 : 4'b0000;
																assign node63542 = (inp[2]) ? 4'b0000 : 4'b0001;
													assign node63545 = (inp[8]) ? node63549 : node63546;
														assign node63546 = (inp[2]) ? 4'b0101 : 4'b0100;
														assign node63549 = (inp[2]) ? node63555 : node63550;
															assign node63550 = (inp[12]) ? 4'b0101 : node63551;
																assign node63551 = (inp[10]) ? 4'b0101 : 4'b0001;
															assign node63555 = (inp[10]) ? 4'b0100 : node63556;
																assign node63556 = (inp[12]) ? 4'b0100 : 4'b0000;
												assign node63560 = (inp[9]) ? node63578 : node63561;
													assign node63561 = (inp[10]) ? node63571 : node63562;
														assign node63562 = (inp[12]) ? 4'b0101 : node63563;
															assign node63563 = (inp[2]) ? node63567 : node63564;
																assign node63564 = (inp[8]) ? 4'b0001 : 4'b0000;
																assign node63567 = (inp[8]) ? 4'b0000 : 4'b0001;
														assign node63571 = (inp[2]) ? node63575 : node63572;
															assign node63572 = (inp[8]) ? 4'b0101 : 4'b0100;
															assign node63575 = (inp[8]) ? 4'b0100 : 4'b0101;
													assign node63578 = (inp[10]) ? node63586 : node63579;
														assign node63579 = (inp[12]) ? 4'b0000 : node63580;
															assign node63580 = (inp[2]) ? node63582 : 4'b0101;
																assign node63582 = (inp[8]) ? 4'b0100 : 4'b0101;
														assign node63586 = (inp[2]) ? 4'b0001 : node63587;
															assign node63587 = (inp[8]) ? 4'b0001 : 4'b0000;
										assign node63591 = (inp[4]) ? node63681 : node63592;
											assign node63592 = (inp[9]) ? node63636 : node63593;
												assign node63593 = (inp[10]) ? node63617 : node63594;
													assign node63594 = (inp[12]) ? node63606 : node63595;
														assign node63595 = (inp[2]) ? node63601 : node63596;
															assign node63596 = (inp[8]) ? 4'b0100 : node63597;
																assign node63597 = (inp[7]) ? 4'b0100 : 4'b0101;
															assign node63601 = (inp[8]) ? 4'b0101 : node63602;
																assign node63602 = (inp[7]) ? 4'b0101 : 4'b0100;
														assign node63606 = (inp[7]) ? node63612 : node63607;
															assign node63607 = (inp[8]) ? node63609 : 4'b0001;
																assign node63609 = (inp[2]) ? 4'b0001 : 4'b0000;
															assign node63612 = (inp[2]) ? node63614 : 4'b0000;
																assign node63614 = (inp[8]) ? 4'b0000 : 4'b0001;
													assign node63617 = (inp[2]) ? node63625 : node63618;
														assign node63618 = (inp[7]) ? node63622 : node63619;
															assign node63619 = (inp[8]) ? 4'b0000 : 4'b0001;
															assign node63622 = (inp[8]) ? 4'b0001 : 4'b0000;
														assign node63625 = (inp[12]) ? node63631 : node63626;
															assign node63626 = (inp[8]) ? node63628 : 4'b0000;
																assign node63628 = (inp[7]) ? 4'b0000 : 4'b0001;
															assign node63631 = (inp[8]) ? 4'b0000 : node63632;
																assign node63632 = (inp[7]) ? 4'b0001 : 4'b0000;
												assign node63636 = (inp[12]) ? node63664 : node63637;
													assign node63637 = (inp[10]) ? node63653 : node63638;
														assign node63638 = (inp[2]) ? node63646 : node63639;
															assign node63639 = (inp[8]) ? node63643 : node63640;
																assign node63640 = (inp[7]) ? 4'b0000 : 4'b0001;
																assign node63643 = (inp[7]) ? 4'b0001 : 4'b0000;
															assign node63646 = (inp[7]) ? node63650 : node63647;
																assign node63647 = (inp[8]) ? 4'b0001 : 4'b0000;
																assign node63650 = (inp[8]) ? 4'b0000 : 4'b0001;
														assign node63653 = (inp[8]) ? node63659 : node63654;
															assign node63654 = (inp[2]) ? node63656 : 4'b0110;
																assign node63656 = (inp[7]) ? 4'b0111 : 4'b0110;
															assign node63659 = (inp[2]) ? 4'b0111 : node63660;
																assign node63660 = (inp[7]) ? 4'b0111 : 4'b0110;
													assign node63664 = (inp[2]) ? node63674 : node63665;
														assign node63665 = (inp[10]) ? 4'b0110 : node63666;
															assign node63666 = (inp[8]) ? node63670 : node63667;
																assign node63667 = (inp[7]) ? 4'b0110 : 4'b0111;
																assign node63670 = (inp[7]) ? 4'b0111 : 4'b0110;
														assign node63674 = (inp[7]) ? node63678 : node63675;
															assign node63675 = (inp[8]) ? 4'b0111 : 4'b0110;
															assign node63678 = (inp[8]) ? 4'b0110 : 4'b0111;
											assign node63681 = (inp[9]) ? node63723 : node63682;
												assign node63682 = (inp[10]) ? node63710 : node63683;
													assign node63683 = (inp[12]) ? node63699 : node63684;
														assign node63684 = (inp[2]) ? node63692 : node63685;
															assign node63685 = (inp[7]) ? node63689 : node63686;
																assign node63686 = (inp[8]) ? 4'b0000 : 4'b0001;
																assign node63689 = (inp[8]) ? 4'b0001 : 4'b0000;
															assign node63692 = (inp[8]) ? node63696 : node63693;
																assign node63693 = (inp[7]) ? 4'b0001 : 4'b0000;
																assign node63696 = (inp[7]) ? 4'b0000 : 4'b0001;
														assign node63699 = (inp[7]) ? node63705 : node63700;
															assign node63700 = (inp[2]) ? node63702 : 4'b0110;
																assign node63702 = (inp[8]) ? 4'b0111 : 4'b0110;
															assign node63705 = (inp[2]) ? node63707 : 4'b0111;
																assign node63707 = (inp[8]) ? 4'b0110 : 4'b0111;
													assign node63710 = (inp[8]) ? node63718 : node63711;
														assign node63711 = (inp[2]) ? node63715 : node63712;
															assign node63712 = (inp[7]) ? 4'b0110 : 4'b0111;
															assign node63715 = (inp[7]) ? 4'b0111 : 4'b0110;
														assign node63718 = (inp[2]) ? 4'b0111 : node63719;
															assign node63719 = (inp[7]) ? 4'b0111 : 4'b0110;
												assign node63723 = (inp[10]) ? node63747 : node63724;
													assign node63724 = (inp[12]) ? node63738 : node63725;
														assign node63725 = (inp[7]) ? node63733 : node63726;
															assign node63726 = (inp[2]) ? node63730 : node63727;
																assign node63727 = (inp[8]) ? 4'b0110 : 4'b0111;
																assign node63730 = (inp[8]) ? 4'b0111 : 4'b0110;
															assign node63733 = (inp[8]) ? node63735 : 4'b0111;
																assign node63735 = (inp[2]) ? 4'b0110 : 4'b0111;
														assign node63738 = (inp[8]) ? node63740 : 4'b0010;
															assign node63740 = (inp[7]) ? node63744 : node63741;
																assign node63741 = (inp[2]) ? 4'b0011 : 4'b0010;
																assign node63744 = (inp[2]) ? 4'b0010 : 4'b0011;
													assign node63747 = (inp[8]) ? node63753 : node63748;
														assign node63748 = (inp[7]) ? 4'b0011 : node63749;
															assign node63749 = (inp[2]) ? 4'b0010 : 4'b0011;
														assign node63753 = (inp[2]) ? node63757 : node63754;
															assign node63754 = (inp[7]) ? 4'b0011 : 4'b0010;
															assign node63757 = (inp[7]) ? 4'b0010 : 4'b0011;
									assign node63760 = (inp[3]) ? node63922 : node63761;
										assign node63761 = (inp[9]) ? node63845 : node63762;
											assign node63762 = (inp[4]) ? node63802 : node63763;
												assign node63763 = (inp[10]) ? node63787 : node63764;
													assign node63764 = (inp[12]) ? node63774 : node63765;
														assign node63765 = (inp[2]) ? 4'b0101 : node63766;
															assign node63766 = (inp[8]) ? node63770 : node63767;
																assign node63767 = (inp[7]) ? 4'b0100 : 4'b0101;
																assign node63770 = (inp[7]) ? 4'b0101 : 4'b0100;
														assign node63774 = (inp[7]) ? node63780 : node63775;
															assign node63775 = (inp[8]) ? node63777 : 4'b0000;
																assign node63777 = (inp[2]) ? 4'b0001 : 4'b0000;
															assign node63780 = (inp[2]) ? node63784 : node63781;
																assign node63781 = (inp[8]) ? 4'b0001 : 4'b0000;
																assign node63784 = (inp[8]) ? 4'b0000 : 4'b0001;
													assign node63787 = (inp[2]) ? node63795 : node63788;
														assign node63788 = (inp[7]) ? node63792 : node63789;
															assign node63789 = (inp[8]) ? 4'b0000 : 4'b0001;
															assign node63792 = (inp[8]) ? 4'b0001 : 4'b0000;
														assign node63795 = (inp[8]) ? node63799 : node63796;
															assign node63796 = (inp[7]) ? 4'b0001 : 4'b0000;
															assign node63799 = (inp[7]) ? 4'b0000 : 4'b0001;
												assign node63802 = (inp[12]) ? node63830 : node63803;
													assign node63803 = (inp[10]) ? node63819 : node63804;
														assign node63804 = (inp[2]) ? node63812 : node63805;
															assign node63805 = (inp[8]) ? node63809 : node63806;
																assign node63806 = (inp[7]) ? 4'b0000 : 4'b0001;
																assign node63809 = (inp[7]) ? 4'b0001 : 4'b0000;
															assign node63812 = (inp[8]) ? node63816 : node63813;
																assign node63813 = (inp[7]) ? 4'b0001 : 4'b0000;
																assign node63816 = (inp[7]) ? 4'b0000 : 4'b0001;
														assign node63819 = (inp[7]) ? node63825 : node63820;
															assign node63820 = (inp[8]) ? 4'b0111 : node63821;
																assign node63821 = (inp[2]) ? 4'b0110 : 4'b0111;
															assign node63825 = (inp[2]) ? node63827 : 4'b0110;
																assign node63827 = (inp[8]) ? 4'b0110 : 4'b0111;
													assign node63830 = (inp[2]) ? node63838 : node63831;
														assign node63831 = (inp[7]) ? node63835 : node63832;
															assign node63832 = (inp[8]) ? 4'b0110 : 4'b0111;
															assign node63835 = (inp[8]) ? 4'b0111 : 4'b0110;
														assign node63838 = (inp[7]) ? node63842 : node63839;
															assign node63839 = (inp[8]) ? 4'b0111 : 4'b0110;
															assign node63842 = (inp[8]) ? 4'b0110 : 4'b0111;
											assign node63845 = (inp[4]) ? node63879 : node63846;
												assign node63846 = (inp[12]) ? node63864 : node63847;
													assign node63847 = (inp[10]) ? node63855 : node63848;
														assign node63848 = (inp[8]) ? node63850 : 4'b0000;
															assign node63850 = (inp[7]) ? node63852 : 4'b0001;
																assign node63852 = (inp[2]) ? 4'b0000 : 4'b0001;
														assign node63855 = (inp[8]) ? node63857 : 4'b0111;
															assign node63857 = (inp[7]) ? node63861 : node63858;
																assign node63858 = (inp[2]) ? 4'b0111 : 4'b0110;
																assign node63861 = (inp[2]) ? 4'b0110 : 4'b0111;
													assign node63864 = (inp[2]) ? node63872 : node63865;
														assign node63865 = (inp[8]) ? node63869 : node63866;
															assign node63866 = (inp[7]) ? 4'b0110 : 4'b0111;
															assign node63869 = (inp[7]) ? 4'b0111 : 4'b0110;
														assign node63872 = (inp[7]) ? node63876 : node63873;
															assign node63873 = (inp[8]) ? 4'b0111 : 4'b0110;
															assign node63876 = (inp[8]) ? 4'b0110 : 4'b0111;
												assign node63879 = (inp[10]) ? node63899 : node63880;
													assign node63880 = (inp[12]) ? node63892 : node63881;
														assign node63881 = (inp[7]) ? node63887 : node63882;
															assign node63882 = (inp[8]) ? 4'b0110 : node63883;
																assign node63883 = (inp[2]) ? 4'b0110 : 4'b0111;
															assign node63887 = (inp[8]) ? 4'b0111 : node63888;
																assign node63888 = (inp[2]) ? 4'b0111 : 4'b0110;
														assign node63892 = (inp[2]) ? node63894 : 4'b0011;
															assign node63894 = (inp[8]) ? 4'b0011 : node63895;
																assign node63895 = (inp[7]) ? 4'b0011 : 4'b0010;
													assign node63899 = (inp[12]) ? node63913 : node63900;
														assign node63900 = (inp[8]) ? node63908 : node63901;
															assign node63901 = (inp[7]) ? node63905 : node63902;
																assign node63902 = (inp[2]) ? 4'b0010 : 4'b0011;
																assign node63905 = (inp[2]) ? 4'b0011 : 4'b0010;
															assign node63908 = (inp[2]) ? 4'b0011 : node63909;
																assign node63909 = (inp[7]) ? 4'b0011 : 4'b0010;
														assign node63913 = (inp[2]) ? node63915 : 4'b0010;
															assign node63915 = (inp[8]) ? node63919 : node63916;
																assign node63916 = (inp[7]) ? 4'b0011 : 4'b0010;
																assign node63919 = (inp[7]) ? 4'b0010 : 4'b0011;
										assign node63922 = (inp[12]) ? node64010 : node63923;
											assign node63923 = (inp[10]) ? node63959 : node63924;
												assign node63924 = (inp[4]) ? node63940 : node63925;
													assign node63925 = (inp[9]) ? node63935 : node63926;
														assign node63926 = (inp[2]) ? 4'b0111 : node63927;
															assign node63927 = (inp[7]) ? node63931 : node63928;
																assign node63928 = (inp[8]) ? 4'b0110 : 4'b0111;
																assign node63931 = (inp[8]) ? 4'b0111 : 4'b0110;
														assign node63935 = (inp[7]) ? 4'b0011 : node63936;
															assign node63936 = (inp[2]) ? 4'b0010 : 4'b0011;
													assign node63940 = (inp[9]) ? node63948 : node63941;
														assign node63941 = (inp[2]) ? 4'b0011 : node63942;
															assign node63942 = (inp[8]) ? node63944 : 4'b0010;
																assign node63944 = (inp[7]) ? 4'b0011 : 4'b0010;
														assign node63948 = (inp[8]) ? node63954 : node63949;
															assign node63949 = (inp[2]) ? 4'b0110 : node63950;
																assign node63950 = (inp[7]) ? 4'b0110 : 4'b0111;
															assign node63954 = (inp[2]) ? node63956 : 4'b0111;
																assign node63956 = (inp[7]) ? 4'b0110 : 4'b0111;
												assign node63959 = (inp[7]) ? node63989 : node63960;
													assign node63960 = (inp[2]) ? node63976 : node63961;
														assign node63961 = (inp[8]) ? node63969 : node63962;
															assign node63962 = (inp[4]) ? node63966 : node63963;
																assign node63963 = (inp[9]) ? 4'b0111 : 4'b0011;
																assign node63966 = (inp[9]) ? 4'b0011 : 4'b0111;
															assign node63969 = (inp[4]) ? node63973 : node63970;
																assign node63970 = (inp[9]) ? 4'b0110 : 4'b0010;
																assign node63973 = (inp[9]) ? 4'b0010 : 4'b0110;
														assign node63976 = (inp[8]) ? node63984 : node63977;
															assign node63977 = (inp[4]) ? node63981 : node63978;
																assign node63978 = (inp[9]) ? 4'b0110 : 4'b0010;
																assign node63981 = (inp[9]) ? 4'b0010 : 4'b0110;
															assign node63984 = (inp[4]) ? node63986 : 4'b0111;
																assign node63986 = (inp[9]) ? 4'b0011 : 4'b0111;
													assign node63989 = (inp[8]) ? node64003 : node63990;
														assign node63990 = (inp[2]) ? node63996 : node63991;
															assign node63991 = (inp[9]) ? 4'b0110 : node63992;
																assign node63992 = (inp[4]) ? 4'b0110 : 4'b0010;
															assign node63996 = (inp[9]) ? node64000 : node63997;
																assign node63997 = (inp[4]) ? 4'b0111 : 4'b0011;
																assign node64000 = (inp[4]) ? 4'b0011 : 4'b0111;
														assign node64003 = (inp[2]) ? 4'b0010 : node64004;
															assign node64004 = (inp[4]) ? 4'b0011 : node64005;
																assign node64005 = (inp[9]) ? 4'b0111 : 4'b0011;
											assign node64010 = (inp[10]) ? node64062 : node64011;
												assign node64011 = (inp[7]) ? node64033 : node64012;
													assign node64012 = (inp[8]) ? node64020 : node64013;
														assign node64013 = (inp[2]) ? node64015 : 4'b0011;
															assign node64015 = (inp[4]) ? node64017 : 4'b0010;
																assign node64017 = (inp[9]) ? 4'b0010 : 4'b0110;
														assign node64020 = (inp[2]) ? node64028 : node64021;
															assign node64021 = (inp[9]) ? node64025 : node64022;
																assign node64022 = (inp[4]) ? 4'b0110 : 4'b0010;
																assign node64025 = (inp[4]) ? 4'b0010 : 4'b0110;
															assign node64028 = (inp[4]) ? 4'b0011 : node64029;
																assign node64029 = (inp[9]) ? 4'b0111 : 4'b0011;
													assign node64033 = (inp[2]) ? node64049 : node64034;
														assign node64034 = (inp[8]) ? node64042 : node64035;
															assign node64035 = (inp[9]) ? node64039 : node64036;
																assign node64036 = (inp[4]) ? 4'b0110 : 4'b0010;
																assign node64039 = (inp[4]) ? 4'b0010 : 4'b0110;
															assign node64042 = (inp[9]) ? node64046 : node64043;
																assign node64043 = (inp[4]) ? 4'b0111 : 4'b0011;
																assign node64046 = (inp[4]) ? 4'b0011 : 4'b0111;
														assign node64049 = (inp[8]) ? node64055 : node64050;
															assign node64050 = (inp[9]) ? 4'b0011 : node64051;
																assign node64051 = (inp[4]) ? 4'b0111 : 4'b0011;
															assign node64055 = (inp[9]) ? node64059 : node64056;
																assign node64056 = (inp[4]) ? 4'b0110 : 4'b0010;
																assign node64059 = (inp[4]) ? 4'b0010 : 4'b0110;
												assign node64062 = (inp[7]) ? node64084 : node64063;
													assign node64063 = (inp[9]) ? node64075 : node64064;
														assign node64064 = (inp[4]) ? node64068 : node64065;
															assign node64065 = (inp[2]) ? 4'b0011 : 4'b0010;
															assign node64068 = (inp[8]) ? node64072 : node64069;
																assign node64069 = (inp[2]) ? 4'b0110 : 4'b0111;
																assign node64072 = (inp[2]) ? 4'b0111 : 4'b0110;
														assign node64075 = (inp[4]) ? node64081 : node64076;
															assign node64076 = (inp[2]) ? node64078 : 4'b0111;
																assign node64078 = (inp[8]) ? 4'b0111 : 4'b0110;
															assign node64081 = (inp[2]) ? 4'b0010 : 4'b0011;
													assign node64084 = (inp[9]) ? node64100 : node64085;
														assign node64085 = (inp[4]) ? node64093 : node64086;
															assign node64086 = (inp[2]) ? node64090 : node64087;
																assign node64087 = (inp[8]) ? 4'b0011 : 4'b0010;
																assign node64090 = (inp[8]) ? 4'b0010 : 4'b0011;
															assign node64093 = (inp[2]) ? node64097 : node64094;
																assign node64094 = (inp[8]) ? 4'b0111 : 4'b0110;
																assign node64097 = (inp[8]) ? 4'b0110 : 4'b0111;
														assign node64100 = (inp[4]) ? node64106 : node64101;
															assign node64101 = (inp[2]) ? node64103 : 4'b0111;
																assign node64103 = (inp[8]) ? 4'b0110 : 4'b0111;
															assign node64106 = (inp[2]) ? 4'b0011 : node64107;
																assign node64107 = (inp[8]) ? 4'b0011 : 4'b0010;
								assign node64111 = (inp[5]) ? node64449 : node64112;
									assign node64112 = (inp[3]) ? node64286 : node64113;
										assign node64113 = (inp[4]) ? node64209 : node64114;
											assign node64114 = (inp[9]) ? node64162 : node64115;
												assign node64115 = (inp[12]) ? node64141 : node64116;
													assign node64116 = (inp[10]) ? node64128 : node64117;
														assign node64117 = (inp[8]) ? node64123 : node64118;
															assign node64118 = (inp[7]) ? node64120 : 4'b0110;
																assign node64120 = (inp[2]) ? 4'b0111 : 4'b0110;
															assign node64123 = (inp[7]) ? node64125 : 4'b0111;
																assign node64125 = (inp[2]) ? 4'b0110 : 4'b0111;
														assign node64128 = (inp[7]) ? node64134 : node64129;
															assign node64129 = (inp[8]) ? 4'b0011 : node64130;
																assign node64130 = (inp[2]) ? 4'b0010 : 4'b0011;
															assign node64134 = (inp[2]) ? node64138 : node64135;
																assign node64135 = (inp[8]) ? 4'b0011 : 4'b0010;
																assign node64138 = (inp[8]) ? 4'b0010 : 4'b0011;
													assign node64141 = (inp[8]) ? node64155 : node64142;
														assign node64142 = (inp[10]) ? node64150 : node64143;
															assign node64143 = (inp[7]) ? node64147 : node64144;
																assign node64144 = (inp[2]) ? 4'b0010 : 4'b0011;
																assign node64147 = (inp[2]) ? 4'b0011 : 4'b0010;
															assign node64150 = (inp[7]) ? node64152 : 4'b0011;
																assign node64152 = (inp[2]) ? 4'b0011 : 4'b0010;
														assign node64155 = (inp[7]) ? node64159 : node64156;
															assign node64156 = (inp[2]) ? 4'b0011 : 4'b0010;
															assign node64159 = (inp[2]) ? 4'b0010 : 4'b0011;
												assign node64162 = (inp[12]) ? node64188 : node64163;
													assign node64163 = (inp[10]) ? node64175 : node64164;
														assign node64164 = (inp[2]) ? node64170 : node64165;
															assign node64165 = (inp[8]) ? 4'b0010 : node64166;
																assign node64166 = (inp[7]) ? 4'b0010 : 4'b0011;
															assign node64170 = (inp[7]) ? node64172 : 4'b0011;
																assign node64172 = (inp[8]) ? 4'b0010 : 4'b0011;
														assign node64175 = (inp[8]) ? node64181 : node64176;
															assign node64176 = (inp[7]) ? 4'b0111 : node64177;
																assign node64177 = (inp[2]) ? 4'b0110 : 4'b0111;
															assign node64181 = (inp[2]) ? node64185 : node64182;
																assign node64182 = (inp[7]) ? 4'b0111 : 4'b0110;
																assign node64185 = (inp[7]) ? 4'b0110 : 4'b0111;
													assign node64188 = (inp[10]) ? node64204 : node64189;
														assign node64189 = (inp[2]) ? node64197 : node64190;
															assign node64190 = (inp[8]) ? node64194 : node64191;
																assign node64191 = (inp[7]) ? 4'b0110 : 4'b0111;
																assign node64194 = (inp[7]) ? 4'b0111 : 4'b0110;
															assign node64197 = (inp[8]) ? node64201 : node64198;
																assign node64198 = (inp[7]) ? 4'b0111 : 4'b0110;
																assign node64201 = (inp[7]) ? 4'b0110 : 4'b0111;
														assign node64204 = (inp[7]) ? 4'b0110 : node64205;
															assign node64205 = (inp[8]) ? 4'b0111 : 4'b0110;
											assign node64209 = (inp[9]) ? node64253 : node64210;
												assign node64210 = (inp[12]) ? node64226 : node64211;
													assign node64211 = (inp[10]) ? node64219 : node64212;
														assign node64212 = (inp[8]) ? node64214 : 4'b0011;
															assign node64214 = (inp[7]) ? node64216 : 4'b0010;
																assign node64216 = (inp[2]) ? 4'b0010 : 4'b0011;
														assign node64219 = (inp[7]) ? node64221 : 4'b0110;
															assign node64221 = (inp[8]) ? 4'b0110 : node64222;
																assign node64222 = (inp[2]) ? 4'b0111 : 4'b0110;
													assign node64226 = (inp[7]) ? node64240 : node64227;
														assign node64227 = (inp[10]) ? node64233 : node64228;
															assign node64228 = (inp[8]) ? 4'b0111 : node64229;
																assign node64229 = (inp[2]) ? 4'b0110 : 4'b0111;
															assign node64233 = (inp[8]) ? node64237 : node64234;
																assign node64234 = (inp[2]) ? 4'b0110 : 4'b0111;
																assign node64237 = (inp[2]) ? 4'b0111 : 4'b0110;
														assign node64240 = (inp[10]) ? node64248 : node64241;
															assign node64241 = (inp[2]) ? node64245 : node64242;
																assign node64242 = (inp[8]) ? 4'b0111 : 4'b0110;
																assign node64245 = (inp[8]) ? 4'b0110 : 4'b0111;
															assign node64248 = (inp[8]) ? 4'b0110 : node64249;
																assign node64249 = (inp[2]) ? 4'b0111 : 4'b0110;
												assign node64253 = (inp[10]) ? node64275 : node64254;
													assign node64254 = (inp[12]) ? node64268 : node64255;
														assign node64255 = (inp[7]) ? node64261 : node64256;
															assign node64256 = (inp[2]) ? 4'b0111 : node64257;
																assign node64257 = (inp[8]) ? 4'b0110 : 4'b0111;
															assign node64261 = (inp[2]) ? node64265 : node64262;
																assign node64262 = (inp[8]) ? 4'b0111 : 4'b0110;
																assign node64265 = (inp[8]) ? 4'b0110 : 4'b0111;
														assign node64268 = (inp[7]) ? node64270 : 4'b0011;
															assign node64270 = (inp[8]) ? node64272 : 4'b0011;
																assign node64272 = (inp[2]) ? 4'b0010 : 4'b0011;
													assign node64275 = (inp[7]) ? node64281 : node64276;
														assign node64276 = (inp[12]) ? node64278 : 4'b0011;
															assign node64278 = (inp[2]) ? 4'b0011 : 4'b0010;
														assign node64281 = (inp[12]) ? 4'b0010 : node64282;
															assign node64282 = (inp[2]) ? 4'b0011 : 4'b0010;
										assign node64286 = (inp[9]) ? node64370 : node64287;
											assign node64287 = (inp[4]) ? node64325 : node64288;
												assign node64288 = (inp[10]) ? node64312 : node64289;
													assign node64289 = (inp[12]) ? node64303 : node64290;
														assign node64290 = (inp[8]) ? node64298 : node64291;
															assign node64291 = (inp[7]) ? node64295 : node64292;
																assign node64292 = (inp[2]) ? 4'b0110 : 4'b0111;
																assign node64295 = (inp[2]) ? 4'b0111 : 4'b0110;
															assign node64298 = (inp[7]) ? 4'b0110 : node64299;
																assign node64299 = (inp[2]) ? 4'b0111 : 4'b0110;
														assign node64303 = (inp[2]) ? node64305 : 4'b0010;
															assign node64305 = (inp[8]) ? node64309 : node64306;
																assign node64306 = (inp[7]) ? 4'b0011 : 4'b0010;
																assign node64309 = (inp[7]) ? 4'b0010 : 4'b0011;
													assign node64312 = (inp[7]) ? node64320 : node64313;
														assign node64313 = (inp[2]) ? node64317 : node64314;
															assign node64314 = (inp[8]) ? 4'b0010 : 4'b0011;
															assign node64317 = (inp[8]) ? 4'b0011 : 4'b0010;
														assign node64320 = (inp[2]) ? 4'b0011 : node64321;
															assign node64321 = (inp[8]) ? 4'b0011 : 4'b0010;
												assign node64325 = (inp[10]) ? node64351 : node64326;
													assign node64326 = (inp[12]) ? node64340 : node64327;
														assign node64327 = (inp[2]) ? node64335 : node64328;
															assign node64328 = (inp[8]) ? node64332 : node64329;
																assign node64329 = (inp[7]) ? 4'b0010 : 4'b0011;
																assign node64332 = (inp[7]) ? 4'b0011 : 4'b0010;
															assign node64335 = (inp[7]) ? 4'b0011 : node64336;
																assign node64336 = (inp[8]) ? 4'b0011 : 4'b0010;
														assign node64340 = (inp[8]) ? node64346 : node64341;
															assign node64341 = (inp[2]) ? 4'b0100 : node64342;
																assign node64342 = (inp[7]) ? 4'b0100 : 4'b0101;
															assign node64346 = (inp[7]) ? 4'b0101 : node64347;
																assign node64347 = (inp[2]) ? 4'b0101 : 4'b0100;
													assign node64351 = (inp[8]) ? node64361 : node64352;
														assign node64352 = (inp[12]) ? 4'b0101 : node64353;
															assign node64353 = (inp[7]) ? node64357 : node64354;
																assign node64354 = (inp[2]) ? 4'b0100 : 4'b0101;
																assign node64357 = (inp[2]) ? 4'b0101 : 4'b0100;
														assign node64361 = (inp[12]) ? 4'b0100 : node64362;
															assign node64362 = (inp[7]) ? node64366 : node64363;
																assign node64363 = (inp[2]) ? 4'b0101 : 4'b0100;
																assign node64366 = (inp[2]) ? 4'b0100 : 4'b0101;
											assign node64370 = (inp[4]) ? node64412 : node64371;
												assign node64371 = (inp[10]) ? node64391 : node64372;
													assign node64372 = (inp[12]) ? node64380 : node64373;
														assign node64373 = (inp[2]) ? node64375 : 4'b0011;
															assign node64375 = (inp[8]) ? node64377 : 4'b0010;
																assign node64377 = (inp[7]) ? 4'b0010 : 4'b0011;
														assign node64380 = (inp[8]) ? node64386 : node64381;
															assign node64381 = (inp[2]) ? node64383 : 4'b0100;
																assign node64383 = (inp[7]) ? 4'b0101 : 4'b0100;
															assign node64386 = (inp[2]) ? node64388 : 4'b0101;
																assign node64388 = (inp[7]) ? 4'b0100 : 4'b0101;
													assign node64391 = (inp[2]) ? node64399 : node64392;
														assign node64392 = (inp[7]) ? node64396 : node64393;
															assign node64393 = (inp[8]) ? 4'b0100 : 4'b0101;
															assign node64396 = (inp[8]) ? 4'b0101 : 4'b0100;
														assign node64399 = (inp[12]) ? node64407 : node64400;
															assign node64400 = (inp[7]) ? node64404 : node64401;
																assign node64401 = (inp[8]) ? 4'b0101 : 4'b0100;
																assign node64404 = (inp[8]) ? 4'b0100 : 4'b0101;
															assign node64407 = (inp[8]) ? node64409 : 4'b0100;
																assign node64409 = (inp[7]) ? 4'b0100 : 4'b0101;
												assign node64412 = (inp[12]) ? node64432 : node64413;
													assign node64413 = (inp[10]) ? node64423 : node64414;
														assign node64414 = (inp[8]) ? node64416 : 4'b0101;
															assign node64416 = (inp[2]) ? node64420 : node64417;
																assign node64417 = (inp[7]) ? 4'b0101 : 4'b0100;
																assign node64420 = (inp[7]) ? 4'b0100 : 4'b0101;
														assign node64423 = (inp[8]) ? 4'b0000 : node64424;
															assign node64424 = (inp[2]) ? node64428 : node64425;
																assign node64425 = (inp[7]) ? 4'b0000 : 4'b0001;
																assign node64428 = (inp[7]) ? 4'b0001 : 4'b0000;
													assign node64432 = (inp[10]) ? node64442 : node64433;
														assign node64433 = (inp[2]) ? 4'b0000 : node64434;
															assign node64434 = (inp[8]) ? node64438 : node64435;
																assign node64435 = (inp[7]) ? 4'b0000 : 4'b0001;
																assign node64438 = (inp[7]) ? 4'b0001 : 4'b0000;
														assign node64442 = (inp[2]) ? node64444 : 4'b0001;
															assign node64444 = (inp[8]) ? node64446 : 4'b0001;
																assign node64446 = (inp[7]) ? 4'b0000 : 4'b0001;
									assign node64449 = (inp[3]) ? node64611 : node64450;
										assign node64450 = (inp[4]) ? node64526 : node64451;
											assign node64451 = (inp[9]) ? node64489 : node64452;
												assign node64452 = (inp[10]) ? node64468 : node64453;
													assign node64453 = (inp[12]) ? node64463 : node64454;
														assign node64454 = (inp[7]) ? node64456 : 4'b0110;
															assign node64456 = (inp[8]) ? node64460 : node64457;
																assign node64457 = (inp[2]) ? 4'b0111 : 4'b0110;
																assign node64460 = (inp[2]) ? 4'b0110 : 4'b0111;
														assign node64463 = (inp[7]) ? node64465 : 4'b0011;
															assign node64465 = (inp[2]) ? 4'b0010 : 4'b0011;
													assign node64468 = (inp[8]) ? node64482 : node64469;
														assign node64469 = (inp[12]) ? node64475 : node64470;
															assign node64470 = (inp[7]) ? 4'b0011 : node64471;
																assign node64471 = (inp[2]) ? 4'b0010 : 4'b0011;
															assign node64475 = (inp[7]) ? node64479 : node64476;
																assign node64476 = (inp[2]) ? 4'b0010 : 4'b0011;
																assign node64479 = (inp[2]) ? 4'b0011 : 4'b0010;
														assign node64482 = (inp[7]) ? node64486 : node64483;
															assign node64483 = (inp[2]) ? 4'b0011 : 4'b0010;
															assign node64486 = (inp[2]) ? 4'b0010 : 4'b0011;
												assign node64489 = (inp[10]) ? node64503 : node64490;
													assign node64490 = (inp[12]) ? node64494 : node64491;
														assign node64491 = (inp[2]) ? 4'b0010 : 4'b0011;
														assign node64494 = (inp[7]) ? node64496 : 4'b0100;
															assign node64496 = (inp[8]) ? node64500 : node64497;
																assign node64497 = (inp[2]) ? 4'b0101 : 4'b0100;
																assign node64500 = (inp[2]) ? 4'b0100 : 4'b0101;
													assign node64503 = (inp[12]) ? node64513 : node64504;
														assign node64504 = (inp[8]) ? node64506 : 4'b0100;
															assign node64506 = (inp[7]) ? node64510 : node64507;
																assign node64507 = (inp[2]) ? 4'b0101 : 4'b0100;
																assign node64510 = (inp[2]) ? 4'b0100 : 4'b0101;
														assign node64513 = (inp[7]) ? node64519 : node64514;
															assign node64514 = (inp[2]) ? node64516 : 4'b0101;
																assign node64516 = (inp[8]) ? 4'b0101 : 4'b0100;
															assign node64519 = (inp[8]) ? node64523 : node64520;
																assign node64520 = (inp[2]) ? 4'b0101 : 4'b0100;
																assign node64523 = (inp[2]) ? 4'b0100 : 4'b0101;
											assign node64526 = (inp[9]) ? node64570 : node64527;
												assign node64527 = (inp[10]) ? node64545 : node64528;
													assign node64528 = (inp[12]) ? node64532 : node64529;
														assign node64529 = (inp[7]) ? 4'b0011 : 4'b0010;
														assign node64532 = (inp[8]) ? node64540 : node64533;
															assign node64533 = (inp[2]) ? node64537 : node64534;
																assign node64534 = (inp[7]) ? 4'b0100 : 4'b0101;
																assign node64537 = (inp[7]) ? 4'b0101 : 4'b0100;
															assign node64540 = (inp[2]) ? node64542 : 4'b0101;
																assign node64542 = (inp[7]) ? 4'b0100 : 4'b0101;
													assign node64545 = (inp[7]) ? node64555 : node64546;
														assign node64546 = (inp[12]) ? 4'b0100 : node64547;
															assign node64547 = (inp[2]) ? node64551 : node64548;
																assign node64548 = (inp[8]) ? 4'b0100 : 4'b0101;
																assign node64551 = (inp[8]) ? 4'b0101 : 4'b0100;
														assign node64555 = (inp[12]) ? node64563 : node64556;
															assign node64556 = (inp[8]) ? node64560 : node64557;
																assign node64557 = (inp[2]) ? 4'b0101 : 4'b0100;
																assign node64560 = (inp[2]) ? 4'b0100 : 4'b0101;
															assign node64563 = (inp[2]) ? node64567 : node64564;
																assign node64564 = (inp[8]) ? 4'b0101 : 4'b0100;
																assign node64567 = (inp[8]) ? 4'b0100 : 4'b0101;
												assign node64570 = (inp[10]) ? node64588 : node64571;
													assign node64571 = (inp[12]) ? node64579 : node64572;
														assign node64572 = (inp[2]) ? node64574 : 4'b0100;
															assign node64574 = (inp[7]) ? node64576 : 4'b0101;
																assign node64576 = (inp[8]) ? 4'b0100 : 4'b0101;
														assign node64579 = (inp[8]) ? node64581 : 4'b0001;
															assign node64581 = (inp[7]) ? node64585 : node64582;
																assign node64582 = (inp[2]) ? 4'b0001 : 4'b0000;
																assign node64585 = (inp[2]) ? 4'b0000 : 4'b0001;
													assign node64588 = (inp[8]) ? node64604 : node64589;
														assign node64589 = (inp[12]) ? node64597 : node64590;
															assign node64590 = (inp[7]) ? node64594 : node64591;
																assign node64591 = (inp[2]) ? 4'b0000 : 4'b0001;
																assign node64594 = (inp[2]) ? 4'b0001 : 4'b0000;
															assign node64597 = (inp[7]) ? node64601 : node64598;
																assign node64598 = (inp[2]) ? 4'b0000 : 4'b0001;
																assign node64601 = (inp[2]) ? 4'b0001 : 4'b0000;
														assign node64604 = (inp[7]) ? node64608 : node64605;
															assign node64605 = (inp[2]) ? 4'b0001 : 4'b0000;
															assign node64608 = (inp[2]) ? 4'b0000 : 4'b0001;
										assign node64611 = (inp[8]) ? node64701 : node64612;
											assign node64612 = (inp[7]) ? node64660 : node64613;
												assign node64613 = (inp[2]) ? node64635 : node64614;
													assign node64614 = (inp[12]) ? node64628 : node64615;
														assign node64615 = (inp[4]) ? node64623 : node64616;
															assign node64616 = (inp[9]) ? node64620 : node64617;
																assign node64617 = (inp[10]) ? 4'b0001 : 4'b0101;
																assign node64620 = (inp[10]) ? 4'b0101 : 4'b0001;
															assign node64623 = (inp[9]) ? node64625 : 4'b0101;
																assign node64625 = (inp[10]) ? 4'b0001 : 4'b0101;
														assign node64628 = (inp[9]) ? node64632 : node64629;
															assign node64629 = (inp[4]) ? 4'b0101 : 4'b0001;
															assign node64632 = (inp[4]) ? 4'b0001 : 4'b0101;
													assign node64635 = (inp[10]) ? node64651 : node64636;
														assign node64636 = (inp[4]) ? node64644 : node64637;
															assign node64637 = (inp[9]) ? node64641 : node64638;
																assign node64638 = (inp[12]) ? 4'b0000 : 4'b0100;
																assign node64641 = (inp[12]) ? 4'b0100 : 4'b0000;
															assign node64644 = (inp[12]) ? node64648 : node64645;
																assign node64645 = (inp[9]) ? 4'b0100 : 4'b0000;
																assign node64648 = (inp[9]) ? 4'b0000 : 4'b0100;
														assign node64651 = (inp[12]) ? 4'b0000 : node64652;
															assign node64652 = (inp[4]) ? node64656 : node64653;
																assign node64653 = (inp[9]) ? 4'b0100 : 4'b0000;
																assign node64656 = (inp[9]) ? 4'b0000 : 4'b0100;
												assign node64660 = (inp[2]) ? node64684 : node64661;
													assign node64661 = (inp[4]) ? node64673 : node64662;
														assign node64662 = (inp[9]) ? node64668 : node64663;
															assign node64663 = (inp[12]) ? 4'b0000 : node64664;
																assign node64664 = (inp[10]) ? 4'b0000 : 4'b0100;
															assign node64668 = (inp[12]) ? 4'b0100 : node64669;
																assign node64669 = (inp[10]) ? 4'b0100 : 4'b0000;
														assign node64673 = (inp[9]) ? node64679 : node64674;
															assign node64674 = (inp[10]) ? 4'b0100 : node64675;
																assign node64675 = (inp[12]) ? 4'b0100 : 4'b0000;
															assign node64679 = (inp[12]) ? 4'b0000 : node64680;
																assign node64680 = (inp[10]) ? 4'b0000 : 4'b0100;
													assign node64684 = (inp[10]) ? 4'b0101 : node64685;
														assign node64685 = (inp[4]) ? node64693 : node64686;
															assign node64686 = (inp[9]) ? node64690 : node64687;
																assign node64687 = (inp[12]) ? 4'b0001 : 4'b0101;
																assign node64690 = (inp[12]) ? 4'b0101 : 4'b0001;
															assign node64693 = (inp[12]) ? node64697 : node64694;
																assign node64694 = (inp[9]) ? 4'b0101 : 4'b0001;
																assign node64697 = (inp[9]) ? 4'b0001 : 4'b0101;
											assign node64701 = (inp[2]) ? node64747 : node64702;
												assign node64702 = (inp[7]) ? node64724 : node64703;
													assign node64703 = (inp[9]) ? node64713 : node64704;
														assign node64704 = (inp[10]) ? 4'b0100 : node64705;
															assign node64705 = (inp[4]) ? node64709 : node64706;
																assign node64706 = (inp[12]) ? 4'b0000 : 4'b0100;
																assign node64709 = (inp[12]) ? 4'b0100 : 4'b0000;
														assign node64713 = (inp[4]) ? node64719 : node64714;
															assign node64714 = (inp[10]) ? 4'b0100 : node64715;
																assign node64715 = (inp[12]) ? 4'b0100 : 4'b0000;
															assign node64719 = (inp[10]) ? 4'b0000 : node64720;
																assign node64720 = (inp[12]) ? 4'b0000 : 4'b0100;
													assign node64724 = (inp[9]) ? node64736 : node64725;
														assign node64725 = (inp[4]) ? node64731 : node64726;
															assign node64726 = (inp[10]) ? 4'b0001 : node64727;
																assign node64727 = (inp[12]) ? 4'b0001 : 4'b0101;
															assign node64731 = (inp[12]) ? 4'b0101 : node64732;
																assign node64732 = (inp[10]) ? 4'b0101 : 4'b0001;
														assign node64736 = (inp[4]) ? node64742 : node64737;
															assign node64737 = (inp[12]) ? 4'b0101 : node64738;
																assign node64738 = (inp[10]) ? 4'b0101 : 4'b0001;
															assign node64742 = (inp[12]) ? 4'b0001 : node64743;
																assign node64743 = (inp[10]) ? 4'b0001 : 4'b0101;
												assign node64747 = (inp[7]) ? node64769 : node64748;
													assign node64748 = (inp[10]) ? node64762 : node64749;
														assign node64749 = (inp[9]) ? node64757 : node64750;
															assign node64750 = (inp[12]) ? node64754 : node64751;
																assign node64751 = (inp[4]) ? 4'b0001 : 4'b0101;
																assign node64754 = (inp[4]) ? 4'b0101 : 4'b0001;
															assign node64757 = (inp[4]) ? 4'b0001 : node64758;
																assign node64758 = (inp[12]) ? 4'b0101 : 4'b0001;
														assign node64762 = (inp[4]) ? node64766 : node64763;
															assign node64763 = (inp[9]) ? 4'b0101 : 4'b0001;
															assign node64766 = (inp[9]) ? 4'b0001 : 4'b0101;
													assign node64769 = (inp[10]) ? node64779 : node64770;
														assign node64770 = (inp[12]) ? node64772 : 4'b0000;
															assign node64772 = (inp[4]) ? node64776 : node64773;
																assign node64773 = (inp[9]) ? 4'b0100 : 4'b0000;
																assign node64776 = (inp[9]) ? 4'b0000 : 4'b0100;
														assign node64779 = (inp[9]) ? node64783 : node64780;
															assign node64780 = (inp[4]) ? 4'b0100 : 4'b0000;
															assign node64783 = (inp[4]) ? 4'b0000 : 4'b0100;
						assign node64786 = (inp[10]) ? node65740 : node64787;
							assign node64787 = (inp[12]) ? node65285 : node64788;
								assign node64788 = (inp[4]) ? node65006 : node64789;
									assign node64789 = (inp[9]) ? node64895 : node64790;
										assign node64790 = (inp[8]) ? node64842 : node64791;
											assign node64791 = (inp[7]) ? node64811 : node64792;
												assign node64792 = (inp[15]) ? node64804 : node64793;
													assign node64793 = (inp[0]) ? node64799 : node64794;
														assign node64794 = (inp[2]) ? 4'b0110 : node64795;
															assign node64795 = (inp[3]) ? 4'b0100 : 4'b0110;
														assign node64799 = (inp[5]) ? node64801 : 4'b0100;
															assign node64801 = (inp[3]) ? 4'b0110 : 4'b0100;
													assign node64804 = (inp[0]) ? node64806 : 4'b0100;
														assign node64806 = (inp[3]) ? node64808 : 4'b0110;
															assign node64808 = (inp[5]) ? 4'b0100 : 4'b0110;
												assign node64811 = (inp[3]) ? node64819 : node64812;
													assign node64812 = (inp[15]) ? node64816 : node64813;
														assign node64813 = (inp[0]) ? 4'b0101 : 4'b0111;
														assign node64816 = (inp[0]) ? 4'b0111 : 4'b0101;
													assign node64819 = (inp[2]) ? node64829 : node64820;
														assign node64820 = (inp[15]) ? 4'b0111 : node64821;
															assign node64821 = (inp[5]) ? node64825 : node64822;
																assign node64822 = (inp[0]) ? 4'b0101 : 4'b0111;
																assign node64825 = (inp[0]) ? 4'b0111 : 4'b0101;
														assign node64829 = (inp[0]) ? node64837 : node64830;
															assign node64830 = (inp[5]) ? node64834 : node64831;
																assign node64831 = (inp[15]) ? 4'b0101 : 4'b0111;
																assign node64834 = (inp[15]) ? 4'b0111 : 4'b0101;
															assign node64837 = (inp[15]) ? 4'b0101 : node64838;
																assign node64838 = (inp[5]) ? 4'b0111 : 4'b0101;
											assign node64842 = (inp[7]) ? node64872 : node64843;
												assign node64843 = (inp[2]) ? node64857 : node64844;
													assign node64844 = (inp[0]) ? node64852 : node64845;
														assign node64845 = (inp[3]) ? node64847 : 4'b0111;
															assign node64847 = (inp[5]) ? node64849 : 4'b0101;
																assign node64849 = (inp[15]) ? 4'b0111 : 4'b0101;
														assign node64852 = (inp[15]) ? node64854 : 4'b0101;
															assign node64854 = (inp[5]) ? 4'b0101 : 4'b0111;
													assign node64857 = (inp[0]) ? node64867 : node64858;
														assign node64858 = (inp[5]) ? node64862 : node64859;
															assign node64859 = (inp[15]) ? 4'b0101 : 4'b0111;
															assign node64862 = (inp[15]) ? 4'b0111 : node64863;
																assign node64863 = (inp[3]) ? 4'b0101 : 4'b0111;
														assign node64867 = (inp[15]) ? 4'b0111 : node64868;
															assign node64868 = (inp[3]) ? 4'b0111 : 4'b0101;
												assign node64872 = (inp[0]) ? node64884 : node64873;
													assign node64873 = (inp[15]) ? node64879 : node64874;
														assign node64874 = (inp[5]) ? node64876 : 4'b0110;
															assign node64876 = (inp[3]) ? 4'b0100 : 4'b0110;
														assign node64879 = (inp[3]) ? node64881 : 4'b0100;
															assign node64881 = (inp[5]) ? 4'b0110 : 4'b0100;
													assign node64884 = (inp[15]) ? node64890 : node64885;
														assign node64885 = (inp[3]) ? node64887 : 4'b0100;
															assign node64887 = (inp[5]) ? 4'b0110 : 4'b0100;
														assign node64890 = (inp[3]) ? node64892 : 4'b0110;
															assign node64892 = (inp[5]) ? 4'b0100 : 4'b0110;
										assign node64895 = (inp[0]) ? node64941 : node64896;
											assign node64896 = (inp[15]) ? node64918 : node64897;
												assign node64897 = (inp[5]) ? node64905 : node64898;
													assign node64898 = (inp[7]) ? node64902 : node64899;
														assign node64899 = (inp[8]) ? 4'b0011 : 4'b0010;
														assign node64902 = (inp[8]) ? 4'b0010 : 4'b0011;
													assign node64905 = (inp[3]) ? node64911 : node64906;
														assign node64906 = (inp[7]) ? 4'b0010 : node64907;
															assign node64907 = (inp[8]) ? 4'b0011 : 4'b0010;
														assign node64911 = (inp[7]) ? node64915 : node64912;
															assign node64912 = (inp[2]) ? 4'b0001 : 4'b0000;
															assign node64915 = (inp[8]) ? 4'b0000 : 4'b0001;
												assign node64918 = (inp[5]) ? node64926 : node64919;
													assign node64919 = (inp[7]) ? node64923 : node64920;
														assign node64920 = (inp[8]) ? 4'b0001 : 4'b0000;
														assign node64923 = (inp[8]) ? 4'b0000 : 4'b0001;
													assign node64926 = (inp[3]) ? node64936 : node64927;
														assign node64927 = (inp[2]) ? 4'b0000 : node64928;
															assign node64928 = (inp[7]) ? node64932 : node64929;
																assign node64929 = (inp[8]) ? 4'b0001 : 4'b0000;
																assign node64932 = (inp[8]) ? 4'b0000 : 4'b0001;
														assign node64936 = (inp[7]) ? node64938 : 4'b0010;
															assign node64938 = (inp[8]) ? 4'b0010 : 4'b0011;
											assign node64941 = (inp[15]) ? node64973 : node64942;
												assign node64942 = (inp[5]) ? node64958 : node64943;
													assign node64943 = (inp[2]) ? node64951 : node64944;
														assign node64944 = (inp[8]) ? node64948 : node64945;
															assign node64945 = (inp[7]) ? 4'b0001 : 4'b0000;
															assign node64948 = (inp[7]) ? 4'b0000 : 4'b0001;
														assign node64951 = (inp[7]) ? node64955 : node64952;
															assign node64952 = (inp[8]) ? 4'b0001 : 4'b0000;
															assign node64955 = (inp[8]) ? 4'b0000 : 4'b0001;
													assign node64958 = (inp[3]) ? node64966 : node64959;
														assign node64959 = (inp[8]) ? node64963 : node64960;
															assign node64960 = (inp[7]) ? 4'b0001 : 4'b0000;
															assign node64963 = (inp[7]) ? 4'b0000 : 4'b0001;
														assign node64966 = (inp[8]) ? node64970 : node64967;
															assign node64967 = (inp[7]) ? 4'b0011 : 4'b0010;
															assign node64970 = (inp[7]) ? 4'b0010 : 4'b0011;
												assign node64973 = (inp[3]) ? node64991 : node64974;
													assign node64974 = (inp[2]) ? node64982 : node64975;
														assign node64975 = (inp[7]) ? node64979 : node64976;
															assign node64976 = (inp[8]) ? 4'b0011 : 4'b0010;
															assign node64979 = (inp[8]) ? 4'b0010 : 4'b0011;
														assign node64982 = (inp[5]) ? node64984 : 4'b0011;
															assign node64984 = (inp[8]) ? node64988 : node64985;
																assign node64985 = (inp[7]) ? 4'b0011 : 4'b0010;
																assign node64988 = (inp[7]) ? 4'b0010 : 4'b0011;
													assign node64991 = (inp[5]) ? node64999 : node64992;
														assign node64992 = (inp[8]) ? node64996 : node64993;
															assign node64993 = (inp[7]) ? 4'b0011 : 4'b0010;
															assign node64996 = (inp[7]) ? 4'b0010 : 4'b0011;
														assign node64999 = (inp[8]) ? node65003 : node65000;
															assign node65000 = (inp[7]) ? 4'b0001 : 4'b0000;
															assign node65003 = (inp[7]) ? 4'b0000 : 4'b0001;
									assign node65006 = (inp[9]) ? node65132 : node65007;
										assign node65007 = (inp[0]) ? node65051 : node65008;
											assign node65008 = (inp[15]) ? node65034 : node65009;
												assign node65009 = (inp[3]) ? node65021 : node65010;
													assign node65010 = (inp[5]) ? node65016 : node65011;
														assign node65011 = (inp[8]) ? node65013 : 4'b0011;
															assign node65013 = (inp[7]) ? 4'b0010 : 4'b0011;
														assign node65016 = (inp[8]) ? 4'b0011 : node65017;
															assign node65017 = (inp[7]) ? 4'b0011 : 4'b0010;
													assign node65021 = (inp[5]) ? node65029 : node65022;
														assign node65022 = (inp[7]) ? node65026 : node65023;
															assign node65023 = (inp[8]) ? 4'b0011 : 4'b0010;
															assign node65026 = (inp[8]) ? 4'b0010 : 4'b0011;
														assign node65029 = (inp[7]) ? 4'b0000 : node65030;
															assign node65030 = (inp[8]) ? 4'b0001 : 4'b0000;
												assign node65034 = (inp[5]) ? node65042 : node65035;
													assign node65035 = (inp[7]) ? node65039 : node65036;
														assign node65036 = (inp[8]) ? 4'b0001 : 4'b0000;
														assign node65039 = (inp[8]) ? 4'b0000 : 4'b0001;
													assign node65042 = (inp[3]) ? node65046 : node65043;
														assign node65043 = (inp[2]) ? 4'b0001 : 4'b0000;
														assign node65046 = (inp[7]) ? 4'b0011 : node65047;
															assign node65047 = (inp[8]) ? 4'b0011 : 4'b0010;
											assign node65051 = (inp[15]) ? node65099 : node65052;
												assign node65052 = (inp[5]) ? node65078 : node65053;
													assign node65053 = (inp[3]) ? node65063 : node65054;
														assign node65054 = (inp[2]) ? node65058 : node65055;
															assign node65055 = (inp[8]) ? 4'b0001 : 4'b0000;
															assign node65058 = (inp[7]) ? node65060 : 4'b0000;
																assign node65060 = (inp[8]) ? 4'b0000 : 4'b0001;
														assign node65063 = (inp[2]) ? node65071 : node65064;
															assign node65064 = (inp[7]) ? node65068 : node65065;
																assign node65065 = (inp[8]) ? 4'b0001 : 4'b0000;
																assign node65068 = (inp[8]) ? 4'b0000 : 4'b0001;
															assign node65071 = (inp[7]) ? node65075 : node65072;
																assign node65072 = (inp[8]) ? 4'b0001 : 4'b0000;
																assign node65075 = (inp[8]) ? 4'b0000 : 4'b0001;
													assign node65078 = (inp[3]) ? node65086 : node65079;
														assign node65079 = (inp[8]) ? node65083 : node65080;
															assign node65080 = (inp[7]) ? 4'b0001 : 4'b0000;
															assign node65083 = (inp[7]) ? 4'b0000 : 4'b0001;
														assign node65086 = (inp[2]) ? node65094 : node65087;
															assign node65087 = (inp[7]) ? node65091 : node65088;
																assign node65088 = (inp[8]) ? 4'b0011 : 4'b0010;
																assign node65091 = (inp[8]) ? 4'b0010 : 4'b0011;
															assign node65094 = (inp[8]) ? 4'b0010 : node65095;
																assign node65095 = (inp[7]) ? 4'b0011 : 4'b0010;
												assign node65099 = (inp[5]) ? node65119 : node65100;
													assign node65100 = (inp[2]) ? node65106 : node65101;
														assign node65101 = (inp[8]) ? node65103 : 4'b0011;
															assign node65103 = (inp[7]) ? 4'b0010 : 4'b0011;
														assign node65106 = (inp[3]) ? node65112 : node65107;
															assign node65107 = (inp[7]) ? 4'b0010 : node65108;
																assign node65108 = (inp[8]) ? 4'b0011 : 4'b0010;
															assign node65112 = (inp[8]) ? node65116 : node65113;
																assign node65113 = (inp[7]) ? 4'b0011 : 4'b0010;
																assign node65116 = (inp[7]) ? 4'b0010 : 4'b0011;
													assign node65119 = (inp[3]) ? node65125 : node65120;
														assign node65120 = (inp[8]) ? node65122 : 4'b0010;
															assign node65122 = (inp[7]) ? 4'b0010 : 4'b0011;
														assign node65125 = (inp[8]) ? node65129 : node65126;
															assign node65126 = (inp[7]) ? 4'b0001 : 4'b0000;
															assign node65129 = (inp[7]) ? 4'b0000 : 4'b0001;
										assign node65132 = (inp[15]) ? node65220 : node65133;
											assign node65133 = (inp[0]) ? node65179 : node65134;
												assign node65134 = (inp[3]) ? node65158 : node65135;
													assign node65135 = (inp[5]) ? node65151 : node65136;
														assign node65136 = (inp[2]) ? node65144 : node65137;
															assign node65137 = (inp[8]) ? node65141 : node65138;
																assign node65138 = (inp[7]) ? 4'b0111 : 4'b0110;
																assign node65141 = (inp[7]) ? 4'b0110 : 4'b0111;
															assign node65144 = (inp[7]) ? node65148 : node65145;
																assign node65145 = (inp[8]) ? 4'b0111 : 4'b0110;
																assign node65148 = (inp[8]) ? 4'b0110 : 4'b0111;
														assign node65151 = (inp[8]) ? node65155 : node65152;
															assign node65152 = (inp[7]) ? 4'b0101 : 4'b0100;
															assign node65155 = (inp[7]) ? 4'b0100 : 4'b0101;
													assign node65158 = (inp[2]) ? node65166 : node65159;
														assign node65159 = (inp[7]) ? node65163 : node65160;
															assign node65160 = (inp[8]) ? 4'b0101 : 4'b0100;
															assign node65163 = (inp[8]) ? 4'b0100 : 4'b0101;
														assign node65166 = (inp[5]) ? node65172 : node65167;
															assign node65167 = (inp[7]) ? node65169 : 4'b0101;
																assign node65169 = (inp[8]) ? 4'b0100 : 4'b0101;
															assign node65172 = (inp[7]) ? node65176 : node65173;
																assign node65173 = (inp[8]) ? 4'b0101 : 4'b0100;
																assign node65176 = (inp[8]) ? 4'b0100 : 4'b0101;
												assign node65179 = (inp[5]) ? node65193 : node65180;
													assign node65180 = (inp[3]) ? node65188 : node65181;
														assign node65181 = (inp[7]) ? node65185 : node65182;
															assign node65182 = (inp[8]) ? 4'b0101 : 4'b0100;
															assign node65185 = (inp[8]) ? 4'b0100 : 4'b0101;
														assign node65188 = (inp[8]) ? node65190 : 4'b0110;
															assign node65190 = (inp[7]) ? 4'b0110 : 4'b0111;
													assign node65193 = (inp[2]) ? node65207 : node65194;
														assign node65194 = (inp[3]) ? node65202 : node65195;
															assign node65195 = (inp[8]) ? node65199 : node65196;
																assign node65196 = (inp[7]) ? 4'b0111 : 4'b0110;
																assign node65199 = (inp[7]) ? 4'b0110 : 4'b0111;
															assign node65202 = (inp[7]) ? node65204 : 4'b0110;
																assign node65204 = (inp[8]) ? 4'b0110 : 4'b0111;
														assign node65207 = (inp[3]) ? node65215 : node65208;
															assign node65208 = (inp[8]) ? node65212 : node65209;
																assign node65209 = (inp[7]) ? 4'b0111 : 4'b0110;
																assign node65212 = (inp[7]) ? 4'b0110 : 4'b0111;
															assign node65215 = (inp[8]) ? node65217 : 4'b0111;
																assign node65217 = (inp[7]) ? 4'b0110 : 4'b0111;
											assign node65220 = (inp[0]) ? node65254 : node65221;
												assign node65221 = (inp[3]) ? node65239 : node65222;
													assign node65222 = (inp[5]) ? node65232 : node65223;
														assign node65223 = (inp[2]) ? node65225 : 4'b0101;
															assign node65225 = (inp[8]) ? node65229 : node65226;
																assign node65226 = (inp[7]) ? 4'b0101 : 4'b0100;
																assign node65229 = (inp[7]) ? 4'b0100 : 4'b0101;
														assign node65232 = (inp[2]) ? node65234 : 4'b0110;
															assign node65234 = (inp[8]) ? node65236 : 4'b0111;
																assign node65236 = (inp[7]) ? 4'b0110 : 4'b0111;
													assign node65239 = (inp[2]) ? node65247 : node65240;
														assign node65240 = (inp[7]) ? node65244 : node65241;
															assign node65241 = (inp[8]) ? 4'b0111 : 4'b0110;
															assign node65244 = (inp[8]) ? 4'b0110 : 4'b0111;
														assign node65247 = (inp[8]) ? node65251 : node65248;
															assign node65248 = (inp[7]) ? 4'b0111 : 4'b0110;
															assign node65251 = (inp[7]) ? 4'b0110 : 4'b0111;
												assign node65254 = (inp[3]) ? node65268 : node65255;
													assign node65255 = (inp[5]) ? node65261 : node65256;
														assign node65256 = (inp[8]) ? 4'b0111 : node65257;
															assign node65257 = (inp[7]) ? 4'b0111 : 4'b0110;
														assign node65261 = (inp[7]) ? node65265 : node65262;
															assign node65262 = (inp[8]) ? 4'b0101 : 4'b0100;
															assign node65265 = (inp[8]) ? 4'b0100 : 4'b0101;
													assign node65268 = (inp[2]) ? node65276 : node65269;
														assign node65269 = (inp[7]) ? node65273 : node65270;
															assign node65270 = (inp[8]) ? 4'b0101 : 4'b0100;
															assign node65273 = (inp[8]) ? 4'b0100 : 4'b0101;
														assign node65276 = (inp[5]) ? 4'b0101 : node65277;
															assign node65277 = (inp[8]) ? node65281 : node65278;
																assign node65278 = (inp[7]) ? 4'b0101 : 4'b0100;
																assign node65281 = (inp[7]) ? 4'b0100 : 4'b0101;
								assign node65285 = (inp[7]) ? node65489 : node65286;
									assign node65286 = (inp[8]) ? node65384 : node65287;
										assign node65287 = (inp[4]) ? node65329 : node65288;
											assign node65288 = (inp[9]) ? node65308 : node65289;
												assign node65289 = (inp[15]) ? node65299 : node65290;
													assign node65290 = (inp[0]) ? node65294 : node65291;
														assign node65291 = (inp[5]) ? 4'b0000 : 4'b0010;
														assign node65294 = (inp[3]) ? node65296 : 4'b0000;
															assign node65296 = (inp[5]) ? 4'b0010 : 4'b0000;
													assign node65299 = (inp[0]) ? node65305 : node65300;
														assign node65300 = (inp[5]) ? node65302 : 4'b0000;
															assign node65302 = (inp[3]) ? 4'b0010 : 4'b0000;
														assign node65305 = (inp[3]) ? 4'b0000 : 4'b0010;
												assign node65308 = (inp[0]) ? node65320 : node65309;
													assign node65309 = (inp[15]) ? node65315 : node65310;
														assign node65310 = (inp[3]) ? 4'b0100 : node65311;
															assign node65311 = (inp[5]) ? 4'b0100 : 4'b0110;
														assign node65315 = (inp[5]) ? 4'b0110 : node65316;
															assign node65316 = (inp[3]) ? 4'b0110 : 4'b0100;
													assign node65320 = (inp[15]) ? node65326 : node65321;
														assign node65321 = (inp[3]) ? 4'b0110 : node65322;
															assign node65322 = (inp[5]) ? 4'b0110 : 4'b0100;
														assign node65326 = (inp[5]) ? 4'b0100 : 4'b0110;
											assign node65329 = (inp[9]) ? node65353 : node65330;
												assign node65330 = (inp[3]) ? node65346 : node65331;
													assign node65331 = (inp[0]) ? node65339 : node65332;
														assign node65332 = (inp[15]) ? node65336 : node65333;
															assign node65333 = (inp[5]) ? 4'b0100 : 4'b0110;
															assign node65336 = (inp[5]) ? 4'b0110 : 4'b0100;
														assign node65339 = (inp[15]) ? node65343 : node65340;
															assign node65340 = (inp[5]) ? 4'b0110 : 4'b0100;
															assign node65343 = (inp[5]) ? 4'b0100 : 4'b0110;
													assign node65346 = (inp[0]) ? node65350 : node65347;
														assign node65347 = (inp[15]) ? 4'b0110 : 4'b0100;
														assign node65350 = (inp[15]) ? 4'b0100 : 4'b0110;
												assign node65353 = (inp[3]) ? node65371 : node65354;
													assign node65354 = (inp[0]) ? node65362 : node65355;
														assign node65355 = (inp[5]) ? node65359 : node65356;
															assign node65356 = (inp[15]) ? 4'b0000 : 4'b0010;
															assign node65359 = (inp[15]) ? 4'b0010 : 4'b0000;
														assign node65362 = (inp[2]) ? 4'b0010 : node65363;
															assign node65363 = (inp[15]) ? node65367 : node65364;
																assign node65364 = (inp[5]) ? 4'b0010 : 4'b0000;
																assign node65367 = (inp[5]) ? 4'b0000 : 4'b0010;
													assign node65371 = (inp[5]) ? node65377 : node65372;
														assign node65372 = (inp[15]) ? 4'b0000 : node65373;
															assign node65373 = (inp[0]) ? 4'b0010 : 4'b0000;
														assign node65377 = (inp[0]) ? node65381 : node65378;
															assign node65378 = (inp[15]) ? 4'b0010 : 4'b0000;
															assign node65381 = (inp[15]) ? 4'b0000 : 4'b0010;
										assign node65384 = (inp[3]) ? node65444 : node65385;
											assign node65385 = (inp[9]) ? node65407 : node65386;
												assign node65386 = (inp[4]) ? node65394 : node65387;
													assign node65387 = (inp[0]) ? node65391 : node65388;
														assign node65388 = (inp[15]) ? 4'b0001 : 4'b0011;
														assign node65391 = (inp[15]) ? 4'b0011 : 4'b0001;
													assign node65394 = (inp[5]) ? node65402 : node65395;
														assign node65395 = (inp[15]) ? node65399 : node65396;
															assign node65396 = (inp[0]) ? 4'b0101 : 4'b0111;
															assign node65399 = (inp[0]) ? 4'b0111 : 4'b0101;
														assign node65402 = (inp[15]) ? 4'b0101 : node65403;
															assign node65403 = (inp[0]) ? 4'b0111 : 4'b0101;
												assign node65407 = (inp[4]) ? node65429 : node65408;
													assign node65408 = (inp[0]) ? node65416 : node65409;
														assign node65409 = (inp[15]) ? node65413 : node65410;
															assign node65410 = (inp[5]) ? 4'b0101 : 4'b0111;
															assign node65413 = (inp[5]) ? 4'b0111 : 4'b0101;
														assign node65416 = (inp[2]) ? node65424 : node65417;
															assign node65417 = (inp[15]) ? node65421 : node65418;
																assign node65418 = (inp[5]) ? 4'b0111 : 4'b0101;
																assign node65421 = (inp[5]) ? 4'b0101 : 4'b0111;
															assign node65424 = (inp[15]) ? 4'b0101 : node65425;
																assign node65425 = (inp[5]) ? 4'b0111 : 4'b0101;
													assign node65429 = (inp[5]) ? node65437 : node65430;
														assign node65430 = (inp[15]) ? node65434 : node65431;
															assign node65431 = (inp[0]) ? 4'b0001 : 4'b0011;
															assign node65434 = (inp[0]) ? 4'b0011 : 4'b0001;
														assign node65437 = (inp[0]) ? node65441 : node65438;
															assign node65438 = (inp[15]) ? 4'b0011 : 4'b0001;
															assign node65441 = (inp[15]) ? 4'b0001 : 4'b0011;
											assign node65444 = (inp[0]) ? node65458 : node65445;
												assign node65445 = (inp[15]) ? node65453 : node65446;
													assign node65446 = (inp[9]) ? node65450 : node65447;
														assign node65447 = (inp[4]) ? 4'b0101 : 4'b0011;
														assign node65450 = (inp[4]) ? 4'b0001 : 4'b0101;
													assign node65453 = (inp[9]) ? node65455 : 4'b0111;
														assign node65455 = (inp[4]) ? 4'b0011 : 4'b0111;
												assign node65458 = (inp[15]) ? node65482 : node65459;
													assign node65459 = (inp[2]) ? node65475 : node65460;
														assign node65460 = (inp[5]) ? node65468 : node65461;
															assign node65461 = (inp[4]) ? node65465 : node65462;
																assign node65462 = (inp[9]) ? 4'b0111 : 4'b0001;
																assign node65465 = (inp[9]) ? 4'b0011 : 4'b0111;
															assign node65468 = (inp[9]) ? node65472 : node65469;
																assign node65469 = (inp[4]) ? 4'b0111 : 4'b0011;
																assign node65472 = (inp[4]) ? 4'b0011 : 4'b0111;
														assign node65475 = (inp[4]) ? node65479 : node65476;
															assign node65476 = (inp[9]) ? 4'b0111 : 4'b0011;
															assign node65479 = (inp[9]) ? 4'b0011 : 4'b0111;
													assign node65482 = (inp[9]) ? 4'b0101 : node65483;
														assign node65483 = (inp[4]) ? 4'b0101 : node65484;
															assign node65484 = (inp[2]) ? 4'b0001 : 4'b0011;
									assign node65489 = (inp[8]) ? node65613 : node65490;
										assign node65490 = (inp[15]) ? node65562 : node65491;
											assign node65491 = (inp[0]) ? node65533 : node65492;
												assign node65492 = (inp[5]) ? node65512 : node65493;
													assign node65493 = (inp[3]) ? node65505 : node65494;
														assign node65494 = (inp[2]) ? node65500 : node65495;
															assign node65495 = (inp[9]) ? 4'b0111 : node65496;
																assign node65496 = (inp[4]) ? 4'b0111 : 4'b0011;
															assign node65500 = (inp[4]) ? node65502 : 4'b0111;
																assign node65502 = (inp[9]) ? 4'b0011 : 4'b0111;
														assign node65505 = (inp[4]) ? node65509 : node65506;
															assign node65506 = (inp[9]) ? 4'b0101 : 4'b0011;
															assign node65509 = (inp[9]) ? 4'b0001 : 4'b0101;
													assign node65512 = (inp[2]) ? node65518 : node65513;
														assign node65513 = (inp[9]) ? 4'b0101 : node65514;
															assign node65514 = (inp[4]) ? 4'b0101 : 4'b0001;
														assign node65518 = (inp[3]) ? node65526 : node65519;
															assign node65519 = (inp[9]) ? node65523 : node65520;
																assign node65520 = (inp[4]) ? 4'b0101 : 4'b0011;
																assign node65523 = (inp[4]) ? 4'b0001 : 4'b0101;
															assign node65526 = (inp[9]) ? node65530 : node65527;
																assign node65527 = (inp[4]) ? 4'b0101 : 4'b0001;
																assign node65530 = (inp[4]) ? 4'b0001 : 4'b0101;
												assign node65533 = (inp[5]) ? node65555 : node65534;
													assign node65534 = (inp[3]) ? node65548 : node65535;
														assign node65535 = (inp[2]) ? node65543 : node65536;
															assign node65536 = (inp[9]) ? node65540 : node65537;
																assign node65537 = (inp[4]) ? 4'b0101 : 4'b0001;
																assign node65540 = (inp[4]) ? 4'b0001 : 4'b0101;
															assign node65543 = (inp[4]) ? 4'b0001 : node65544;
																assign node65544 = (inp[9]) ? 4'b0101 : 4'b0001;
														assign node65548 = (inp[9]) ? node65552 : node65549;
															assign node65549 = (inp[4]) ? 4'b0111 : 4'b0001;
															assign node65552 = (inp[4]) ? 4'b0011 : 4'b0111;
													assign node65555 = (inp[4]) ? node65559 : node65556;
														assign node65556 = (inp[9]) ? 4'b0111 : 4'b0001;
														assign node65559 = (inp[9]) ? 4'b0011 : 4'b0111;
											assign node65562 = (inp[0]) ? node65588 : node65563;
												assign node65563 = (inp[3]) ? node65579 : node65564;
													assign node65564 = (inp[5]) ? node65572 : node65565;
														assign node65565 = (inp[9]) ? node65569 : node65566;
															assign node65566 = (inp[4]) ? 4'b0101 : 4'b0001;
															assign node65569 = (inp[4]) ? 4'b0001 : 4'b0101;
														assign node65572 = (inp[4]) ? node65576 : node65573;
															assign node65573 = (inp[9]) ? 4'b0111 : 4'b0001;
															assign node65576 = (inp[9]) ? 4'b0011 : 4'b0111;
													assign node65579 = (inp[9]) ? node65585 : node65580;
														assign node65580 = (inp[4]) ? 4'b0111 : node65581;
															assign node65581 = (inp[5]) ? 4'b0011 : 4'b0001;
														assign node65585 = (inp[4]) ? 4'b0011 : 4'b0111;
												assign node65588 = (inp[5]) ? node65604 : node65589;
													assign node65589 = (inp[3]) ? node65597 : node65590;
														assign node65590 = (inp[9]) ? node65594 : node65591;
															assign node65591 = (inp[4]) ? 4'b0111 : 4'b0011;
															assign node65594 = (inp[4]) ? 4'b0011 : 4'b0111;
														assign node65597 = (inp[9]) ? node65601 : node65598;
															assign node65598 = (inp[4]) ? 4'b0101 : 4'b0011;
															assign node65601 = (inp[2]) ? 4'b0101 : 4'b0001;
													assign node65604 = (inp[9]) ? node65610 : node65605;
														assign node65605 = (inp[4]) ? 4'b0101 : node65606;
															assign node65606 = (inp[3]) ? 4'b0001 : 4'b0011;
														assign node65610 = (inp[4]) ? 4'b0001 : 4'b0101;
										assign node65613 = (inp[5]) ? node65673 : node65614;
											assign node65614 = (inp[15]) ? node65648 : node65615;
												assign node65615 = (inp[0]) ? node65633 : node65616;
													assign node65616 = (inp[3]) ? node65626 : node65617;
														assign node65617 = (inp[2]) ? 4'b0110 : node65618;
															assign node65618 = (inp[4]) ? node65622 : node65619;
																assign node65619 = (inp[9]) ? 4'b0110 : 4'b0010;
																assign node65622 = (inp[9]) ? 4'b0010 : 4'b0110;
														assign node65626 = (inp[9]) ? node65630 : node65627;
															assign node65627 = (inp[4]) ? 4'b0100 : 4'b0010;
															assign node65630 = (inp[4]) ? 4'b0000 : 4'b0100;
													assign node65633 = (inp[3]) ? node65641 : node65634;
														assign node65634 = (inp[9]) ? node65638 : node65635;
															assign node65635 = (inp[4]) ? 4'b0100 : 4'b0000;
															assign node65638 = (inp[4]) ? 4'b0000 : 4'b0100;
														assign node65641 = (inp[2]) ? node65643 : 4'b0110;
															assign node65643 = (inp[9]) ? node65645 : 4'b0000;
																assign node65645 = (inp[4]) ? 4'b0010 : 4'b0110;
												assign node65648 = (inp[9]) ? node65658 : node65649;
													assign node65649 = (inp[4]) ? node65651 : 4'b0010;
														assign node65651 = (inp[3]) ? node65655 : node65652;
															assign node65652 = (inp[0]) ? 4'b0110 : 4'b0100;
															assign node65655 = (inp[0]) ? 4'b0100 : 4'b0110;
													assign node65658 = (inp[4]) ? node65666 : node65659;
														assign node65659 = (inp[0]) ? node65663 : node65660;
															assign node65660 = (inp[3]) ? 4'b0110 : 4'b0100;
															assign node65663 = (inp[3]) ? 4'b0100 : 4'b0110;
														assign node65666 = (inp[0]) ? node65670 : node65667;
															assign node65667 = (inp[3]) ? 4'b0010 : 4'b0000;
															assign node65670 = (inp[3]) ? 4'b0000 : 4'b0010;
											assign node65673 = (inp[9]) ? node65715 : node65674;
												assign node65674 = (inp[4]) ? node65702 : node65675;
													assign node65675 = (inp[3]) ? node65689 : node65676;
														assign node65676 = (inp[2]) ? node65682 : node65677;
															assign node65677 = (inp[0]) ? 4'b0010 : node65678;
																assign node65678 = (inp[15]) ? 4'b0000 : 4'b0010;
															assign node65682 = (inp[0]) ? node65686 : node65683;
																assign node65683 = (inp[15]) ? 4'b0000 : 4'b0010;
																assign node65686 = (inp[15]) ? 4'b0010 : 4'b0000;
														assign node65689 = (inp[2]) ? node65695 : node65690;
															assign node65690 = (inp[15]) ? node65692 : 4'b0000;
																assign node65692 = (inp[0]) ? 4'b0000 : 4'b0010;
															assign node65695 = (inp[15]) ? node65699 : node65696;
																assign node65696 = (inp[0]) ? 4'b0010 : 4'b0000;
																assign node65699 = (inp[0]) ? 4'b0000 : 4'b0010;
													assign node65702 = (inp[2]) ? node65710 : node65703;
														assign node65703 = (inp[0]) ? node65707 : node65704;
															assign node65704 = (inp[15]) ? 4'b0110 : 4'b0100;
															assign node65707 = (inp[3]) ? 4'b0110 : 4'b0100;
														assign node65710 = (inp[15]) ? node65712 : 4'b0100;
															assign node65712 = (inp[0]) ? 4'b0100 : 4'b0110;
												assign node65715 = (inp[4]) ? node65723 : node65716;
													assign node65716 = (inp[15]) ? node65720 : node65717;
														assign node65717 = (inp[0]) ? 4'b0110 : 4'b0100;
														assign node65720 = (inp[0]) ? 4'b0100 : 4'b0110;
													assign node65723 = (inp[3]) ? node65735 : node65724;
														assign node65724 = (inp[2]) ? node65730 : node65725;
															assign node65725 = (inp[0]) ? node65727 : 4'b0000;
																assign node65727 = (inp[15]) ? 4'b0000 : 4'b0010;
															assign node65730 = (inp[0]) ? 4'b0010 : node65731;
																assign node65731 = (inp[15]) ? 4'b0010 : 4'b0000;
														assign node65735 = (inp[0]) ? 4'b0000 : node65736;
															assign node65736 = (inp[15]) ? 4'b0010 : 4'b0000;
							assign node65740 = (inp[5]) ? node66108 : node65741;
								assign node65741 = (inp[8]) ? node65945 : node65742;
									assign node65742 = (inp[7]) ? node65828 : node65743;
										assign node65743 = (inp[0]) ? node65797 : node65744;
											assign node65744 = (inp[15]) ? node65766 : node65745;
												assign node65745 = (inp[3]) ? node65759 : node65746;
													assign node65746 = (inp[2]) ? node65754 : node65747;
														assign node65747 = (inp[4]) ? node65751 : node65748;
															assign node65748 = (inp[9]) ? 4'b0110 : 4'b0010;
															assign node65751 = (inp[12]) ? 4'b0010 : 4'b0110;
														assign node65754 = (inp[9]) ? 4'b0010 : node65755;
															assign node65755 = (inp[4]) ? 4'b0110 : 4'b0010;
													assign node65759 = (inp[4]) ? node65763 : node65760;
														assign node65760 = (inp[9]) ? 4'b0100 : 4'b0010;
														assign node65763 = (inp[9]) ? 4'b0000 : 4'b0100;
												assign node65766 = (inp[3]) ? node65790 : node65767;
													assign node65767 = (inp[12]) ? node65781 : node65768;
														assign node65768 = (inp[2]) ? node65776 : node65769;
															assign node65769 = (inp[4]) ? node65773 : node65770;
																assign node65770 = (inp[9]) ? 4'b0100 : 4'b0000;
																assign node65773 = (inp[9]) ? 4'b0000 : 4'b0100;
															assign node65776 = (inp[9]) ? node65778 : 4'b0000;
																assign node65778 = (inp[4]) ? 4'b0000 : 4'b0100;
														assign node65781 = (inp[2]) ? 4'b0100 : node65782;
															assign node65782 = (inp[4]) ? node65786 : node65783;
																assign node65783 = (inp[9]) ? 4'b0100 : 4'b0000;
																assign node65786 = (inp[9]) ? 4'b0000 : 4'b0100;
													assign node65790 = (inp[9]) ? node65794 : node65791;
														assign node65791 = (inp[4]) ? 4'b0110 : 4'b0000;
														assign node65794 = (inp[4]) ? 4'b0010 : 4'b0110;
											assign node65797 = (inp[15]) ? node65813 : node65798;
												assign node65798 = (inp[3]) ? node65806 : node65799;
													assign node65799 = (inp[4]) ? node65803 : node65800;
														assign node65800 = (inp[9]) ? 4'b0100 : 4'b0000;
														assign node65803 = (inp[9]) ? 4'b0000 : 4'b0100;
													assign node65806 = (inp[4]) ? node65810 : node65807;
														assign node65807 = (inp[9]) ? 4'b0110 : 4'b0000;
														assign node65810 = (inp[9]) ? 4'b0010 : 4'b0110;
												assign node65813 = (inp[3]) ? node65821 : node65814;
													assign node65814 = (inp[4]) ? node65818 : node65815;
														assign node65815 = (inp[9]) ? 4'b0110 : 4'b0010;
														assign node65818 = (inp[9]) ? 4'b0010 : 4'b0110;
													assign node65821 = (inp[9]) ? node65825 : node65822;
														assign node65822 = (inp[4]) ? 4'b0100 : 4'b0010;
														assign node65825 = (inp[4]) ? 4'b0000 : 4'b0100;
										assign node65828 = (inp[9]) ? node65890 : node65829;
											assign node65829 = (inp[4]) ? node65855 : node65830;
												assign node65830 = (inp[12]) ? node65848 : node65831;
													assign node65831 = (inp[2]) ? node65839 : node65832;
														assign node65832 = (inp[0]) ? node65836 : node65833;
															assign node65833 = (inp[15]) ? 4'b0001 : 4'b0011;
															assign node65836 = (inp[15]) ? 4'b0011 : 4'b0001;
														assign node65839 = (inp[3]) ? node65843 : node65840;
															assign node65840 = (inp[15]) ? 4'b0011 : 4'b0001;
															assign node65843 = (inp[0]) ? 4'b0011 : node65844;
																assign node65844 = (inp[15]) ? 4'b0001 : 4'b0011;
													assign node65848 = (inp[0]) ? node65852 : node65849;
														assign node65849 = (inp[15]) ? 4'b0001 : 4'b0011;
														assign node65852 = (inp[15]) ? 4'b0011 : 4'b0001;
												assign node65855 = (inp[3]) ? node65877 : node65856;
													assign node65856 = (inp[2]) ? node65870 : node65857;
														assign node65857 = (inp[12]) ? node65863 : node65858;
															assign node65858 = (inp[15]) ? 4'b0111 : node65859;
																assign node65859 = (inp[0]) ? 4'b0101 : 4'b0111;
															assign node65863 = (inp[0]) ? node65867 : node65864;
																assign node65864 = (inp[15]) ? 4'b0101 : 4'b0111;
																assign node65867 = (inp[15]) ? 4'b0111 : 4'b0101;
														assign node65870 = (inp[15]) ? node65874 : node65871;
															assign node65871 = (inp[0]) ? 4'b0101 : 4'b0111;
															assign node65874 = (inp[0]) ? 4'b0111 : 4'b0101;
													assign node65877 = (inp[2]) ? node65885 : node65878;
														assign node65878 = (inp[0]) ? node65882 : node65879;
															assign node65879 = (inp[15]) ? 4'b0111 : 4'b0101;
															assign node65882 = (inp[15]) ? 4'b0101 : 4'b0111;
														assign node65885 = (inp[15]) ? node65887 : 4'b0101;
															assign node65887 = (inp[0]) ? 4'b0101 : 4'b0111;
											assign node65890 = (inp[4]) ? node65920 : node65891;
												assign node65891 = (inp[12]) ? node65905 : node65892;
													assign node65892 = (inp[3]) ? node65898 : node65893;
														assign node65893 = (inp[2]) ? node65895 : 4'b0101;
															assign node65895 = (inp[15]) ? 4'b0101 : 4'b0111;
														assign node65898 = (inp[0]) ? node65902 : node65899;
															assign node65899 = (inp[15]) ? 4'b0111 : 4'b0101;
															assign node65902 = (inp[15]) ? 4'b0101 : 4'b0111;
													assign node65905 = (inp[0]) ? node65913 : node65906;
														assign node65906 = (inp[15]) ? node65910 : node65907;
															assign node65907 = (inp[3]) ? 4'b0101 : 4'b0111;
															assign node65910 = (inp[3]) ? 4'b0111 : 4'b0101;
														assign node65913 = (inp[15]) ? node65917 : node65914;
															assign node65914 = (inp[3]) ? 4'b0111 : 4'b0101;
															assign node65917 = (inp[3]) ? 4'b0101 : 4'b0111;
												assign node65920 = (inp[15]) ? node65936 : node65921;
													assign node65921 = (inp[2]) ? node65929 : node65922;
														assign node65922 = (inp[0]) ? node65926 : node65923;
															assign node65923 = (inp[3]) ? 4'b0001 : 4'b0011;
															assign node65926 = (inp[3]) ? 4'b0011 : 4'b0001;
														assign node65929 = (inp[3]) ? node65933 : node65930;
															assign node65930 = (inp[0]) ? 4'b0001 : 4'b0011;
															assign node65933 = (inp[0]) ? 4'b0011 : 4'b0001;
													assign node65936 = (inp[12]) ? node65938 : 4'b0011;
														assign node65938 = (inp[3]) ? node65942 : node65939;
															assign node65939 = (inp[0]) ? 4'b0011 : 4'b0001;
															assign node65942 = (inp[0]) ? 4'b0001 : 4'b0011;
									assign node65945 = (inp[7]) ? node66029 : node65946;
										assign node65946 = (inp[9]) ? node65984 : node65947;
											assign node65947 = (inp[4]) ? node65955 : node65948;
												assign node65948 = (inp[0]) ? node65952 : node65949;
													assign node65949 = (inp[15]) ? 4'b0001 : 4'b0011;
													assign node65952 = (inp[15]) ? 4'b0011 : 4'b0001;
												assign node65955 = (inp[2]) ? node65969 : node65956;
													assign node65956 = (inp[3]) ? node65962 : node65957;
														assign node65957 = (inp[0]) ? 4'b0101 : node65958;
															assign node65958 = (inp[15]) ? 4'b0101 : 4'b0111;
														assign node65962 = (inp[0]) ? node65966 : node65963;
															assign node65963 = (inp[15]) ? 4'b0111 : 4'b0101;
															assign node65966 = (inp[15]) ? 4'b0101 : 4'b0111;
													assign node65969 = (inp[3]) ? node65977 : node65970;
														assign node65970 = (inp[0]) ? node65974 : node65971;
															assign node65971 = (inp[15]) ? 4'b0101 : 4'b0111;
															assign node65974 = (inp[15]) ? 4'b0111 : 4'b0101;
														assign node65977 = (inp[0]) ? node65981 : node65978;
															assign node65978 = (inp[15]) ? 4'b0111 : 4'b0101;
															assign node65981 = (inp[15]) ? 4'b0101 : 4'b0111;
											assign node65984 = (inp[4]) ? node66014 : node65985;
												assign node65985 = (inp[15]) ? node66001 : node65986;
													assign node65986 = (inp[12]) ? node65994 : node65987;
														assign node65987 = (inp[3]) ? node65991 : node65988;
															assign node65988 = (inp[0]) ? 4'b0101 : 4'b0111;
															assign node65991 = (inp[0]) ? 4'b0111 : 4'b0101;
														assign node65994 = (inp[0]) ? node65998 : node65995;
															assign node65995 = (inp[3]) ? 4'b0101 : 4'b0111;
															assign node65998 = (inp[3]) ? 4'b0111 : 4'b0101;
													assign node66001 = (inp[2]) ? node66009 : node66002;
														assign node66002 = (inp[3]) ? node66006 : node66003;
															assign node66003 = (inp[0]) ? 4'b0111 : 4'b0101;
															assign node66006 = (inp[0]) ? 4'b0101 : 4'b0111;
														assign node66009 = (inp[0]) ? 4'b0101 : node66010;
															assign node66010 = (inp[3]) ? 4'b0111 : 4'b0101;
												assign node66014 = (inp[15]) ? node66022 : node66015;
													assign node66015 = (inp[0]) ? node66019 : node66016;
														assign node66016 = (inp[3]) ? 4'b0001 : 4'b0011;
														assign node66019 = (inp[3]) ? 4'b0011 : 4'b0001;
													assign node66022 = (inp[0]) ? node66026 : node66023;
														assign node66023 = (inp[3]) ? 4'b0011 : 4'b0001;
														assign node66026 = (inp[3]) ? 4'b0001 : 4'b0011;
										assign node66029 = (inp[0]) ? node66069 : node66030;
											assign node66030 = (inp[15]) ? node66054 : node66031;
												assign node66031 = (inp[3]) ? node66047 : node66032;
													assign node66032 = (inp[2]) ? node66040 : node66033;
														assign node66033 = (inp[9]) ? node66037 : node66034;
															assign node66034 = (inp[4]) ? 4'b0110 : 4'b0010;
															assign node66037 = (inp[4]) ? 4'b0010 : 4'b0110;
														assign node66040 = (inp[9]) ? node66044 : node66041;
															assign node66041 = (inp[4]) ? 4'b0110 : 4'b0010;
															assign node66044 = (inp[4]) ? 4'b0010 : 4'b0110;
													assign node66047 = (inp[4]) ? node66051 : node66048;
														assign node66048 = (inp[9]) ? 4'b0100 : 4'b0010;
														assign node66051 = (inp[9]) ? 4'b0000 : 4'b0100;
												assign node66054 = (inp[3]) ? node66062 : node66055;
													assign node66055 = (inp[4]) ? node66059 : node66056;
														assign node66056 = (inp[9]) ? 4'b0100 : 4'b0000;
														assign node66059 = (inp[9]) ? 4'b0000 : 4'b0100;
													assign node66062 = (inp[9]) ? node66066 : node66063;
														assign node66063 = (inp[4]) ? 4'b0110 : 4'b0000;
														assign node66066 = (inp[4]) ? 4'b0010 : 4'b0110;
											assign node66069 = (inp[15]) ? node66087 : node66070;
												assign node66070 = (inp[3]) ? node66080 : node66071;
													assign node66071 = (inp[2]) ? 4'b0000 : node66072;
														assign node66072 = (inp[9]) ? node66076 : node66073;
															assign node66073 = (inp[4]) ? 4'b0100 : 4'b0000;
															assign node66076 = (inp[4]) ? 4'b0000 : 4'b0100;
													assign node66080 = (inp[9]) ? node66084 : node66081;
														assign node66081 = (inp[4]) ? 4'b0110 : 4'b0000;
														assign node66084 = (inp[4]) ? 4'b0010 : 4'b0110;
												assign node66087 = (inp[3]) ? node66101 : node66088;
													assign node66088 = (inp[12]) ? node66096 : node66089;
														assign node66089 = (inp[9]) ? node66093 : node66090;
															assign node66090 = (inp[4]) ? 4'b0110 : 4'b0010;
															assign node66093 = (inp[4]) ? 4'b0010 : 4'b0110;
														assign node66096 = (inp[4]) ? 4'b0110 : node66097;
															assign node66097 = (inp[9]) ? 4'b0110 : 4'b0010;
													assign node66101 = (inp[4]) ? node66105 : node66102;
														assign node66102 = (inp[9]) ? 4'b0100 : 4'b0010;
														assign node66105 = (inp[9]) ? 4'b0000 : 4'b0100;
								assign node66108 = (inp[7]) ? node66308 : node66109;
									assign node66109 = (inp[8]) ? node66253 : node66110;
										assign node66110 = (inp[2]) ? node66164 : node66111;
											assign node66111 = (inp[0]) ? node66141 : node66112;
												assign node66112 = (inp[15]) ? node66132 : node66113;
													assign node66113 = (inp[12]) ? node66119 : node66114;
														assign node66114 = (inp[9]) ? node66116 : 4'b0100;
															assign node66116 = (inp[4]) ? 4'b0000 : 4'b0100;
														assign node66119 = (inp[3]) ? node66127 : node66120;
															assign node66120 = (inp[9]) ? node66124 : node66121;
																assign node66121 = (inp[4]) ? 4'b0100 : 4'b0010;
																assign node66124 = (inp[4]) ? 4'b0000 : 4'b0100;
															assign node66127 = (inp[4]) ? 4'b0100 : node66128;
																assign node66128 = (inp[9]) ? 4'b0100 : 4'b0000;
													assign node66132 = (inp[4]) ? node66138 : node66133;
														assign node66133 = (inp[9]) ? 4'b0110 : node66134;
															assign node66134 = (inp[3]) ? 4'b0010 : 4'b0000;
														assign node66138 = (inp[9]) ? 4'b0010 : 4'b0110;
												assign node66141 = (inp[15]) ? node66155 : node66142;
													assign node66142 = (inp[3]) ? node66150 : node66143;
														assign node66143 = (inp[4]) ? node66147 : node66144;
															assign node66144 = (inp[9]) ? 4'b0110 : 4'b0000;
															assign node66147 = (inp[9]) ? 4'b0010 : 4'b0110;
														assign node66150 = (inp[4]) ? 4'b0010 : node66151;
															assign node66151 = (inp[12]) ? 4'b0010 : 4'b0110;
													assign node66155 = (inp[4]) ? node66161 : node66156;
														assign node66156 = (inp[9]) ? 4'b0100 : node66157;
															assign node66157 = (inp[3]) ? 4'b0000 : 4'b0010;
														assign node66161 = (inp[9]) ? 4'b0000 : 4'b0100;
											assign node66164 = (inp[12]) ? node66206 : node66165;
												assign node66165 = (inp[3]) ? node66185 : node66166;
													assign node66166 = (inp[15]) ? node66180 : node66167;
														assign node66167 = (inp[0]) ? node66173 : node66168;
															assign node66168 = (inp[9]) ? node66170 : 4'b0010;
																assign node66170 = (inp[4]) ? 4'b0000 : 4'b0100;
															assign node66173 = (inp[9]) ? node66177 : node66174;
																assign node66174 = (inp[4]) ? 4'b0110 : 4'b0000;
																assign node66177 = (inp[4]) ? 4'b0010 : 4'b0110;
														assign node66180 = (inp[4]) ? node66182 : 4'b0010;
															assign node66182 = (inp[9]) ? 4'b0010 : 4'b0110;
													assign node66185 = (inp[9]) ? node66195 : node66186;
														assign node66186 = (inp[4]) ? 4'b0100 : node66187;
															assign node66187 = (inp[15]) ? node66191 : node66188;
																assign node66188 = (inp[0]) ? 4'b0010 : 4'b0000;
																assign node66191 = (inp[0]) ? 4'b0000 : 4'b0010;
														assign node66195 = (inp[4]) ? node66201 : node66196;
															assign node66196 = (inp[15]) ? node66198 : 4'b0110;
																assign node66198 = (inp[0]) ? 4'b0100 : 4'b0110;
															assign node66201 = (inp[15]) ? 4'b0010 : node66202;
																assign node66202 = (inp[0]) ? 4'b0010 : 4'b0000;
												assign node66206 = (inp[9]) ? node66236 : node66207;
													assign node66207 = (inp[4]) ? node66223 : node66208;
														assign node66208 = (inp[15]) ? node66216 : node66209;
															assign node66209 = (inp[0]) ? node66213 : node66210;
																assign node66210 = (inp[3]) ? 4'b0000 : 4'b0010;
																assign node66213 = (inp[3]) ? 4'b0010 : 4'b0000;
															assign node66216 = (inp[0]) ? node66220 : node66217;
																assign node66217 = (inp[3]) ? 4'b0010 : 4'b0000;
																assign node66220 = (inp[3]) ? 4'b0000 : 4'b0010;
														assign node66223 = (inp[3]) ? node66229 : node66224;
															assign node66224 = (inp[15]) ? node66226 : 4'b0110;
																assign node66226 = (inp[0]) ? 4'b0100 : 4'b0110;
															assign node66229 = (inp[15]) ? node66233 : node66230;
																assign node66230 = (inp[0]) ? 4'b0110 : 4'b0100;
																assign node66233 = (inp[0]) ? 4'b0100 : 4'b0110;
													assign node66236 = (inp[4]) ? node66248 : node66237;
														assign node66237 = (inp[3]) ? node66243 : node66238;
															assign node66238 = (inp[15]) ? 4'b0100 : node66239;
																assign node66239 = (inp[0]) ? 4'b0110 : 4'b0100;
															assign node66243 = (inp[0]) ? 4'b0110 : node66244;
																assign node66244 = (inp[15]) ? 4'b0110 : 4'b0100;
														assign node66248 = (inp[15]) ? node66250 : 4'b0000;
															assign node66250 = (inp[0]) ? 4'b0000 : 4'b0010;
										assign node66253 = (inp[15]) ? node66273 : node66254;
											assign node66254 = (inp[0]) ? node66264 : node66255;
												assign node66255 = (inp[4]) ? node66261 : node66256;
													assign node66256 = (inp[9]) ? 4'b0101 : node66257;
														assign node66257 = (inp[3]) ? 4'b0001 : 4'b0011;
													assign node66261 = (inp[9]) ? 4'b0001 : 4'b0101;
												assign node66264 = (inp[4]) ? node66270 : node66265;
													assign node66265 = (inp[9]) ? 4'b0111 : node66266;
														assign node66266 = (inp[3]) ? 4'b0011 : 4'b0001;
													assign node66270 = (inp[9]) ? 4'b0011 : 4'b0111;
											assign node66273 = (inp[0]) ? node66283 : node66274;
												assign node66274 = (inp[9]) ? node66280 : node66275;
													assign node66275 = (inp[4]) ? 4'b0111 : node66276;
														assign node66276 = (inp[3]) ? 4'b0011 : 4'b0001;
													assign node66280 = (inp[4]) ? 4'b0011 : 4'b0111;
												assign node66283 = (inp[2]) ? node66297 : node66284;
													assign node66284 = (inp[3]) ? node66290 : node66285;
														assign node66285 = (inp[9]) ? node66287 : 4'b0011;
															assign node66287 = (inp[4]) ? 4'b0001 : 4'b0101;
														assign node66290 = (inp[4]) ? node66294 : node66291;
															assign node66291 = (inp[9]) ? 4'b0101 : 4'b0001;
															assign node66294 = (inp[9]) ? 4'b0001 : 4'b0101;
													assign node66297 = (inp[3]) ? node66303 : node66298;
														assign node66298 = (inp[4]) ? node66300 : 4'b0101;
															assign node66300 = (inp[9]) ? 4'b0001 : 4'b0101;
														assign node66303 = (inp[9]) ? 4'b0101 : node66304;
															assign node66304 = (inp[4]) ? 4'b0101 : 4'b0001;
									assign node66308 = (inp[8]) ? node66378 : node66309;
										assign node66309 = (inp[0]) ? node66343 : node66310;
											assign node66310 = (inp[15]) ? node66334 : node66311;
												assign node66311 = (inp[3]) ? node66319 : node66312;
													assign node66312 = (inp[9]) ? node66316 : node66313;
														assign node66313 = (inp[4]) ? 4'b0101 : 4'b0011;
														assign node66316 = (inp[4]) ? 4'b0001 : 4'b0101;
													assign node66319 = (inp[12]) ? node66327 : node66320;
														assign node66320 = (inp[4]) ? node66324 : node66321;
															assign node66321 = (inp[9]) ? 4'b0101 : 4'b0001;
															assign node66324 = (inp[9]) ? 4'b0001 : 4'b0101;
														assign node66327 = (inp[2]) ? node66329 : 4'b0001;
															assign node66329 = (inp[9]) ? 4'b0001 : node66330;
																assign node66330 = (inp[4]) ? 4'b0101 : 4'b0001;
												assign node66334 = (inp[9]) ? node66340 : node66335;
													assign node66335 = (inp[4]) ? 4'b0111 : node66336;
														assign node66336 = (inp[3]) ? 4'b0011 : 4'b0001;
													assign node66340 = (inp[4]) ? 4'b0011 : 4'b0111;
											assign node66343 = (inp[15]) ? node66369 : node66344;
												assign node66344 = (inp[3]) ? node66352 : node66345;
													assign node66345 = (inp[9]) ? node66349 : node66346;
														assign node66346 = (inp[4]) ? 4'b0111 : 4'b0001;
														assign node66349 = (inp[4]) ? 4'b0011 : 4'b0111;
													assign node66352 = (inp[12]) ? node66360 : node66353;
														assign node66353 = (inp[4]) ? node66357 : node66354;
															assign node66354 = (inp[9]) ? 4'b0111 : 4'b0011;
															assign node66357 = (inp[9]) ? 4'b0011 : 4'b0111;
														assign node66360 = (inp[2]) ? node66362 : 4'b0111;
															assign node66362 = (inp[9]) ? node66366 : node66363;
																assign node66363 = (inp[4]) ? 4'b0111 : 4'b0011;
																assign node66366 = (inp[4]) ? 4'b0011 : 4'b0111;
												assign node66369 = (inp[9]) ? node66375 : node66370;
													assign node66370 = (inp[4]) ? 4'b0101 : node66371;
														assign node66371 = (inp[3]) ? 4'b0001 : 4'b0011;
													assign node66375 = (inp[4]) ? 4'b0001 : 4'b0101;
										assign node66378 = (inp[4]) ? node66448 : node66379;
											assign node66379 = (inp[9]) ? node66427 : node66380;
												assign node66380 = (inp[12]) ? node66412 : node66381;
													assign node66381 = (inp[2]) ? node66397 : node66382;
														assign node66382 = (inp[0]) ? node66390 : node66383;
															assign node66383 = (inp[15]) ? node66387 : node66384;
																assign node66384 = (inp[3]) ? 4'b0000 : 4'b0010;
																assign node66387 = (inp[3]) ? 4'b0010 : 4'b0000;
															assign node66390 = (inp[15]) ? node66394 : node66391;
																assign node66391 = (inp[3]) ? 4'b0010 : 4'b0000;
																assign node66394 = (inp[3]) ? 4'b0000 : 4'b0010;
														assign node66397 = (inp[3]) ? node66405 : node66398;
															assign node66398 = (inp[15]) ? node66402 : node66399;
																assign node66399 = (inp[0]) ? 4'b0000 : 4'b0010;
																assign node66402 = (inp[0]) ? 4'b0010 : 4'b0000;
															assign node66405 = (inp[0]) ? node66409 : node66406;
																assign node66406 = (inp[15]) ? 4'b0010 : 4'b0000;
																assign node66409 = (inp[15]) ? 4'b0000 : 4'b0010;
													assign node66412 = (inp[15]) ? node66420 : node66413;
														assign node66413 = (inp[2]) ? 4'b0000 : node66414;
															assign node66414 = (inp[0]) ? node66416 : 4'b0000;
																assign node66416 = (inp[3]) ? 4'b0010 : 4'b0000;
														assign node66420 = (inp[3]) ? node66424 : node66421;
															assign node66421 = (inp[0]) ? 4'b0010 : 4'b0000;
															assign node66424 = (inp[0]) ? 4'b0000 : 4'b0010;
												assign node66427 = (inp[2]) ? node66433 : node66428;
													assign node66428 = (inp[0]) ? 4'b0110 : node66429;
														assign node66429 = (inp[15]) ? 4'b0110 : 4'b0100;
													assign node66433 = (inp[12]) ? node66441 : node66434;
														assign node66434 = (inp[3]) ? 4'b0100 : node66435;
															assign node66435 = (inp[0]) ? 4'b0100 : node66436;
																assign node66436 = (inp[15]) ? 4'b0110 : 4'b0100;
														assign node66441 = (inp[0]) ? node66445 : node66442;
															assign node66442 = (inp[15]) ? 4'b0110 : 4'b0100;
															assign node66445 = (inp[15]) ? 4'b0100 : 4'b0110;
											assign node66448 = (inp[9]) ? node66480 : node66449;
												assign node66449 = (inp[3]) ? node66473 : node66450;
													assign node66450 = (inp[12]) ? node66466 : node66451;
														assign node66451 = (inp[2]) ? node66459 : node66452;
															assign node66452 = (inp[15]) ? node66456 : node66453;
																assign node66453 = (inp[0]) ? 4'b0110 : 4'b0100;
																assign node66456 = (inp[0]) ? 4'b0100 : 4'b0110;
															assign node66459 = (inp[0]) ? node66463 : node66460;
																assign node66460 = (inp[15]) ? 4'b0110 : 4'b0100;
																assign node66463 = (inp[15]) ? 4'b0100 : 4'b0110;
														assign node66466 = (inp[0]) ? node66470 : node66467;
															assign node66467 = (inp[15]) ? 4'b0110 : 4'b0100;
															assign node66470 = (inp[15]) ? 4'b0100 : 4'b0110;
													assign node66473 = (inp[15]) ? node66477 : node66474;
														assign node66474 = (inp[0]) ? 4'b0110 : 4'b0100;
														assign node66477 = (inp[0]) ? 4'b0100 : 4'b0110;
												assign node66480 = (inp[12]) ? node66488 : node66481;
													assign node66481 = (inp[0]) ? node66485 : node66482;
														assign node66482 = (inp[15]) ? 4'b0010 : 4'b0000;
														assign node66485 = (inp[15]) ? 4'b0000 : 4'b0010;
													assign node66488 = (inp[15]) ? node66492 : node66489;
														assign node66489 = (inp[0]) ? 4'b0010 : 4'b0000;
														assign node66492 = (inp[0]) ? 4'b0000 : 4'b0010;

endmodule