module dtc_split25_bm39 (
	input  wire [14-1:0] inp,
	output wire [14-1:0] outp
);

	wire [14-1:0] node1;
	wire [14-1:0] node3;
	wire [14-1:0] node4;
	wire [14-1:0] node5;
	wire [14-1:0] node6;
	wire [14-1:0] node7;
	wire [14-1:0] node8;
	wire [14-1:0] node9;
	wire [14-1:0] node10;
	wire [14-1:0] node11;
	wire [14-1:0] node12;
	wire [14-1:0] node17;
	wire [14-1:0] node18;
	wire [14-1:0] node19;
	wire [14-1:0] node21;
	wire [14-1:0] node24;
	wire [14-1:0] node25;
	wire [14-1:0] node29;
	wire [14-1:0] node30;
	wire [14-1:0] node33;
	wire [14-1:0] node36;
	wire [14-1:0] node37;
	wire [14-1:0] node38;
	wire [14-1:0] node39;
	wire [14-1:0] node40;
	wire [14-1:0] node44;
	wire [14-1:0] node47;
	wire [14-1:0] node50;
	wire [14-1:0] node51;
	wire [14-1:0] node52;
	wire [14-1:0] node53;
	wire [14-1:0] node57;
	wire [14-1:0] node59;
	wire [14-1:0] node62;
	wire [14-1:0] node65;
	wire [14-1:0] node66;
	wire [14-1:0] node67;
	wire [14-1:0] node68;
	wire [14-1:0] node70;
	wire [14-1:0] node72;
	wire [14-1:0] node75;
	wire [14-1:0] node76;
	wire [14-1:0] node79;
	wire [14-1:0] node82;
	wire [14-1:0] node83;
	wire [14-1:0] node84;
	wire [14-1:0] node87;
	wire [14-1:0] node90;
	wire [14-1:0] node91;
	wire [14-1:0] node94;
	wire [14-1:0] node97;
	wire [14-1:0] node98;
	wire [14-1:0] node99;
	wire [14-1:0] node104;
	wire [14-1:0] node105;
	wire [14-1:0] node106;
	wire [14-1:0] node107;
	wire [14-1:0] node108;
	wire [14-1:0] node111;
	wire [14-1:0] node112;
	wire [14-1:0] node116;
	wire [14-1:0] node117;
	wire [14-1:0] node118;
	wire [14-1:0] node120;
	wire [14-1:0] node123;
	wire [14-1:0] node126;
	wire [14-1:0] node127;
	wire [14-1:0] node130;
	wire [14-1:0] node131;
	wire [14-1:0] node134;
	wire [14-1:0] node137;
	wire [14-1:0] node138;
	wire [14-1:0] node139;
	wire [14-1:0] node141;
	wire [14-1:0] node144;
	wire [14-1:0] node146;
	wire [14-1:0] node147;
	wire [14-1:0] node151;
	wire [14-1:0] node152;
	wire [14-1:0] node153;
	wire [14-1:0] node156;
	wire [14-1:0] node158;
	wire [14-1:0] node161;
	wire [14-1:0] node162;
	wire [14-1:0] node165;
	wire [14-1:0] node168;
	wire [14-1:0] node169;
	wire [14-1:0] node170;
	wire [14-1:0] node171;
	wire [14-1:0] node173;
	wire [14-1:0] node176;
	wire [14-1:0] node177;
	wire [14-1:0] node179;
	wire [14-1:0] node183;
	wire [14-1:0] node184;
	wire [14-1:0] node185;
	wire [14-1:0] node189;
	wire [14-1:0] node190;
	wire [14-1:0] node193;
	wire [14-1:0] node195;
	wire [14-1:0] node199;
	wire [14-1:0] node200;
	wire [14-1:0] node201;
	wire [14-1:0] node202;
	wire [14-1:0] node203;
	wire [14-1:0] node204;
	wire [14-1:0] node206;
	wire [14-1:0] node208;
	wire [14-1:0] node211;
	wire [14-1:0] node212;
	wire [14-1:0] node215;
	wire [14-1:0] node218;
	wire [14-1:0] node219;
	wire [14-1:0] node220;
	wire [14-1:0] node223;
	wire [14-1:0] node226;
	wire [14-1:0] node229;
	wire [14-1:0] node230;
	wire [14-1:0] node231;
	wire [14-1:0] node234;
	wire [14-1:0] node235;
	wire [14-1:0] node237;
	wire [14-1:0] node240;
	wire [14-1:0] node241;
	wire [14-1:0] node246;
	wire [14-1:0] node247;
	wire [14-1:0] node249;
	wire [14-1:0] node250;
	wire [14-1:0] node251;
	wire [14-1:0] node252;
	wire [14-1:0] node256;
	wire [14-1:0] node257;
	wire [14-1:0] node260;
	wire [14-1:0] node263;
	wire [14-1:0] node264;
	wire [14-1:0] node269;
	wire [14-1:0] node271;
	wire [14-1:0] node272;
	wire [14-1:0] node273;
	wire [14-1:0] node274;
	wire [14-1:0] node277;
	wire [14-1:0] node278;
	wire [14-1:0] node282;
	wire [14-1:0] node283;
	wire [14-1:0] node286;
	wire [14-1:0] node290;
	wire [14-1:0] node291;
	wire [14-1:0] node292;
	wire [14-1:0] node293;
	wire [14-1:0] node294;
	wire [14-1:0] node295;
	wire [14-1:0] node297;
	wire [14-1:0] node298;
	wire [14-1:0] node300;
	wire [14-1:0] node303;
	wire [14-1:0] node306;
	wire [14-1:0] node307;
	wire [14-1:0] node308;
	wire [14-1:0] node309;
	wire [14-1:0] node313;
	wire [14-1:0] node316;
	wire [14-1:0] node317;
	wire [14-1:0] node318;
	wire [14-1:0] node323;
	wire [14-1:0] node324;
	wire [14-1:0] node325;
	wire [14-1:0] node327;
	wire [14-1:0] node330;
	wire [14-1:0] node332;
	wire [14-1:0] node335;
	wire [14-1:0] node336;
	wire [14-1:0] node337;
	wire [14-1:0] node340;
	wire [14-1:0] node341;
	wire [14-1:0] node345;
	wire [14-1:0] node346;
	wire [14-1:0] node347;
	wire [14-1:0] node351;
	wire [14-1:0] node354;
	wire [14-1:0] node355;
	wire [14-1:0] node356;
	wire [14-1:0] node357;
	wire [14-1:0] node359;
	wire [14-1:0] node362;
	wire [14-1:0] node363;
	wire [14-1:0] node368;
	wire [14-1:0] node370;
	wire [14-1:0] node371;
	wire [14-1:0] node372;
	wire [14-1:0] node375;
	wire [14-1:0] node379;
	wire [14-1:0] node381;
	wire [14-1:0] node382;
	wire [14-1:0] node383;
	wire [14-1:0] node384;
	wire [14-1:0] node385;
	wire [14-1:0] node392;
	wire [14-1:0] node393;
	wire [14-1:0] node394;
	wire [14-1:0] node396;
	wire [14-1:0] node397;
	wire [14-1:0] node398;
	wire [14-1:0] node399;
	wire [14-1:0] node403;
	wire [14-1:0] node404;
	wire [14-1:0] node405;
	wire [14-1:0] node409;
	wire [14-1:0] node412;
	wire [14-1:0] node417;
	wire [14-1:0] node418;
	wire [14-1:0] node419;
	wire [14-1:0] node420;
	wire [14-1:0] node421;
	wire [14-1:0] node422;
	wire [14-1:0] node423;
	wire [14-1:0] node424;
	wire [14-1:0] node427;
	wire [14-1:0] node430;
	wire [14-1:0] node431;
	wire [14-1:0] node432;
	wire [14-1:0] node433;
	wire [14-1:0] node439;
	wire [14-1:0] node440;
	wire [14-1:0] node441;
	wire [14-1:0] node442;
	wire [14-1:0] node444;
	wire [14-1:0] node447;
	wire [14-1:0] node448;
	wire [14-1:0] node451;
	wire [14-1:0] node454;
	wire [14-1:0] node457;
	wire [14-1:0] node458;
	wire [14-1:0] node459;
	wire [14-1:0] node462;
	wire [14-1:0] node465;
	wire [14-1:0] node468;
	wire [14-1:0] node469;
	wire [14-1:0] node470;
	wire [14-1:0] node471;
	wire [14-1:0] node474;
	wire [14-1:0] node475;
	wire [14-1:0] node478;
	wire [14-1:0] node481;
	wire [14-1:0] node482;
	wire [14-1:0] node484;
	wire [14-1:0] node489;
	wire [14-1:0] node490;
	wire [14-1:0] node491;
	wire [14-1:0] node492;
	wire [14-1:0] node493;
	wire [14-1:0] node496;
	wire [14-1:0] node497;
	wire [14-1:0] node500;
	wire [14-1:0] node501;
	wire [14-1:0] node505;
	wire [14-1:0] node506;
	wire [14-1:0] node507;
	wire [14-1:0] node512;
	wire [14-1:0] node513;
	wire [14-1:0] node514;
	wire [14-1:0] node517;
	wire [14-1:0] node518;
	wire [14-1:0] node524;
	wire [14-1:0] node525;
	wire [14-1:0] node526;
	wire [14-1:0] node527;
	wire [14-1:0] node528;
	wire [14-1:0] node529;
	wire [14-1:0] node531;
	wire [14-1:0] node533;
	wire [14-1:0] node536;
	wire [14-1:0] node537;
	wire [14-1:0] node541;
	wire [14-1:0] node542;
	wire [14-1:0] node544;
	wire [14-1:0] node548;
	wire [14-1:0] node549;
	wire [14-1:0] node550;
	wire [14-1:0] node552;
	wire [14-1:0] node555;
	wire [14-1:0] node559;
	wire [14-1:0] node561;
	wire [14-1:0] node562;
	wire [14-1:0] node564;
	wire [14-1:0] node567;
	wire [14-1:0] node568;
	wire [14-1:0] node569;
	wire [14-1:0] node572;
	wire [14-1:0] node576;
	wire [14-1:0] node577;
	wire [14-1:0] node579;
	wire [14-1:0] node580;
	wire [14-1:0] node581;
	wire [14-1:0] node582;
	wire [14-1:0] node583;
	wire [14-1:0] node586;
	wire [14-1:0] node590;
	wire [14-1:0] node592;
	wire [14-1:0] node594;
	wire [14-1:0] node597;
	wire [14-1:0] node598;
	wire [14-1:0] node604;
	wire [14-1:0] node605;
	wire [14-1:0] node606;
	wire [14-1:0] node607;
	wire [14-1:0] node608;
	wire [14-1:0] node609;
	wire [14-1:0] node610;
	wire [14-1:0] node611;
	wire [14-1:0] node612;
	wire [14-1:0] node613;
	wire [14-1:0] node614;
	wire [14-1:0] node618;
	wire [14-1:0] node619;
	wire [14-1:0] node624;
	wire [14-1:0] node625;
	wire [14-1:0] node626;
	wire [14-1:0] node629;
	wire [14-1:0] node630;
	wire [14-1:0] node634;
	wire [14-1:0] node636;
	wire [14-1:0] node637;
	wire [14-1:0] node640;
	wire [14-1:0] node643;
	wire [14-1:0] node644;
	wire [14-1:0] node645;
	wire [14-1:0] node646;
	wire [14-1:0] node647;
	wire [14-1:0] node651;
	wire [14-1:0] node652;
	wire [14-1:0] node656;
	wire [14-1:0] node657;
	wire [14-1:0] node658;
	wire [14-1:0] node663;
	wire [14-1:0] node664;
	wire [14-1:0] node665;
	wire [14-1:0] node667;
	wire [14-1:0] node670;
	wire [14-1:0] node671;
	wire [14-1:0] node674;
	wire [14-1:0] node677;
	wire [14-1:0] node678;
	wire [14-1:0] node680;
	wire [14-1:0] node683;
	wire [14-1:0] node686;
	wire [14-1:0] node687;
	wire [14-1:0] node688;
	wire [14-1:0] node689;
	wire [14-1:0] node690;
	wire [14-1:0] node694;
	wire [14-1:0] node696;
	wire [14-1:0] node697;
	wire [14-1:0] node700;
	wire [14-1:0] node703;
	wire [14-1:0] node704;
	wire [14-1:0] node705;
	wire [14-1:0] node706;
	wire [14-1:0] node709;
	wire [14-1:0] node712;
	wire [14-1:0] node713;
	wire [14-1:0] node714;
	wire [14-1:0] node719;
	wire [14-1:0] node721;
	wire [14-1:0] node722;
	wire [14-1:0] node726;
	wire [14-1:0] node727;
	wire [14-1:0] node728;
	wire [14-1:0] node729;
	wire [14-1:0] node730;
	wire [14-1:0] node733;
	wire [14-1:0] node734;
	wire [14-1:0] node738;
	wire [14-1:0] node740;
	wire [14-1:0] node743;
	wire [14-1:0] node744;
	wire [14-1:0] node746;
	wire [14-1:0] node749;
	wire [14-1:0] node750;
	wire [14-1:0] node753;
	wire [14-1:0] node756;
	wire [14-1:0] node757;
	wire [14-1:0] node758;
	wire [14-1:0] node759;
	wire [14-1:0] node762;
	wire [14-1:0] node764;
	wire [14-1:0] node767;
	wire [14-1:0] node768;
	wire [14-1:0] node772;
	wire [14-1:0] node774;
	wire [14-1:0] node775;
	wire [14-1:0] node776;
	wire [14-1:0] node781;
	wire [14-1:0] node782;
	wire [14-1:0] node783;
	wire [14-1:0] node784;
	wire [14-1:0] node785;
	wire [14-1:0] node786;
	wire [14-1:0] node788;
	wire [14-1:0] node791;
	wire [14-1:0] node792;
	wire [14-1:0] node794;
	wire [14-1:0] node795;
	wire [14-1:0] node800;
	wire [14-1:0] node802;
	wire [14-1:0] node804;
	wire [14-1:0] node807;
	wire [14-1:0] node808;
	wire [14-1:0] node809;
	wire [14-1:0] node812;
	wire [14-1:0] node813;
	wire [14-1:0] node814;
	wire [14-1:0] node818;
	wire [14-1:0] node821;
	wire [14-1:0] node823;
	wire [14-1:0] node824;
	wire [14-1:0] node826;
	wire [14-1:0] node829;
	wire [14-1:0] node832;
	wire [14-1:0] node833;
	wire [14-1:0] node834;
	wire [14-1:0] node835;
	wire [14-1:0] node836;
	wire [14-1:0] node839;
	wire [14-1:0] node841;
	wire [14-1:0] node844;
	wire [14-1:0] node845;
	wire [14-1:0] node847;
	wire [14-1:0] node852;
	wire [14-1:0] node853;
	wire [14-1:0] node855;
	wire [14-1:0] node857;
	wire [14-1:0] node860;
	wire [14-1:0] node861;
	wire [14-1:0] node863;
	wire [14-1:0] node866;
	wire [14-1:0] node869;
	wire [14-1:0] node870;
	wire [14-1:0] node871;
	wire [14-1:0] node872;
	wire [14-1:0] node874;
	wire [14-1:0] node876;
	wire [14-1:0] node879;
	wire [14-1:0] node880;
	wire [14-1:0] node881;
	wire [14-1:0] node884;
	wire [14-1:0] node886;
	wire [14-1:0] node892;
	wire [14-1:0] node893;
	wire [14-1:0] node894;
	wire [14-1:0] node895;
	wire [14-1:0] node896;
	wire [14-1:0] node897;
	wire [14-1:0] node899;
	wire [14-1:0] node900;
	wire [14-1:0] node902;
	wire [14-1:0] node906;
	wire [14-1:0] node907;
	wire [14-1:0] node908;
	wire [14-1:0] node911;
	wire [14-1:0] node914;
	wire [14-1:0] node915;
	wire [14-1:0] node916;
	wire [14-1:0] node920;
	wire [14-1:0] node922;
	wire [14-1:0] node925;
	wire [14-1:0] node926;
	wire [14-1:0] node927;
	wire [14-1:0] node928;
	wire [14-1:0] node932;
	wire [14-1:0] node933;
	wire [14-1:0] node935;
	wire [14-1:0] node938;
	wire [14-1:0] node942;
	wire [14-1:0] node943;
	wire [14-1:0] node944;
	wire [14-1:0] node945;
	wire [14-1:0] node946;
	wire [14-1:0] node948;
	wire [14-1:0] node951;
	wire [14-1:0] node953;
	wire [14-1:0] node956;
	wire [14-1:0] node959;
	wire [14-1:0] node962;
	wire [14-1:0] node963;
	wire [14-1:0] node965;
	wire [14-1:0] node966;
	wire [14-1:0] node971;
	wire [14-1:0] node972;
	wire [14-1:0] node973;
	wire [14-1:0] node974;
	wire [14-1:0] node975;
	wire [14-1:0] node977;
	wire [14-1:0] node980;
	wire [14-1:0] node983;
	wire [14-1:0] node984;
	wire [14-1:0] node985;
	wire [14-1:0] node988;
	wire [14-1:0] node991;
	wire [14-1:0] node993;
	wire [14-1:0] node996;
	wire [14-1:0] node997;
	wire [14-1:0] node999;
	wire [14-1:0] node1002;
	wire [14-1:0] node1003;
	wire [14-1:0] node1004;
	wire [14-1:0] node1008;
	wire [14-1:0] node1009;
	wire [14-1:0] node1012;
	wire [14-1:0] node1015;
	wire [14-1:0] node1016;
	wire [14-1:0] node1017;
	wire [14-1:0] node1018;
	wire [14-1:0] node1021;
	wire [14-1:0] node1023;
	wire [14-1:0] node1026;
	wire [14-1:0] node1027;
	wire [14-1:0] node1032;
	wire [14-1:0] node1033;
	wire [14-1:0] node1034;
	wire [14-1:0] node1035;
	wire [14-1:0] node1036;
	wire [14-1:0] node1037;
	wire [14-1:0] node1040;
	wire [14-1:0] node1042;
	wire [14-1:0] node1044;
	wire [14-1:0] node1047;
	wire [14-1:0] node1048;
	wire [14-1:0] node1049;
	wire [14-1:0] node1053;
	wire [14-1:0] node1054;
	wire [14-1:0] node1056;
	wire [14-1:0] node1059;
	wire [14-1:0] node1061;
	wire [14-1:0] node1064;
	wire [14-1:0] node1065;
	wire [14-1:0] node1066;
	wire [14-1:0] node1067;
	wire [14-1:0] node1072;
	wire [14-1:0] node1074;
	wire [14-1:0] node1075;
	wire [14-1:0] node1076;
	wire [14-1:0] node1083;
	wire [14-1:0] node1084;
	wire [14-1:0] node1085;
	wire [14-1:0] node1086;
	wire [14-1:0] node1087;
	wire [14-1:0] node1088;
	wire [14-1:0] node1089;
	wire [14-1:0] node1090;
	wire [14-1:0] node1091;
	wire [14-1:0] node1093;
	wire [14-1:0] node1096;
	wire [14-1:0] node1099;
	wire [14-1:0] node1100;
	wire [14-1:0] node1101;
	wire [14-1:0] node1104;
	wire [14-1:0] node1107;
	wire [14-1:0] node1109;
	wire [14-1:0] node1112;
	wire [14-1:0] node1113;
	wire [14-1:0] node1114;
	wire [14-1:0] node1116;
	wire [14-1:0] node1119;
	wire [14-1:0] node1122;
	wire [14-1:0] node1123;
	wire [14-1:0] node1125;
	wire [14-1:0] node1128;
	wire [14-1:0] node1129;
	wire [14-1:0] node1133;
	wire [14-1:0] node1134;
	wire [14-1:0] node1135;
	wire [14-1:0] node1137;
	wire [14-1:0] node1140;
	wire [14-1:0] node1142;
	wire [14-1:0] node1145;
	wire [14-1:0] node1146;
	wire [14-1:0] node1150;
	wire [14-1:0] node1151;
	wire [14-1:0] node1152;
	wire [14-1:0] node1153;
	wire [14-1:0] node1155;
	wire [14-1:0] node1158;
	wire [14-1:0] node1159;
	wire [14-1:0] node1162;
	wire [14-1:0] node1163;
	wire [14-1:0] node1167;
	wire [14-1:0] node1168;
	wire [14-1:0] node1169;
	wire [14-1:0] node1171;
	wire [14-1:0] node1177;
	wire [14-1:0] node1178;
	wire [14-1:0] node1179;
	wire [14-1:0] node1180;
	wire [14-1:0] node1182;
	wire [14-1:0] node1183;
	wire [14-1:0] node1187;
	wire [14-1:0] node1188;
	wire [14-1:0] node1190;
	wire [14-1:0] node1193;
	wire [14-1:0] node1195;
	wire [14-1:0] node1198;
	wire [14-1:0] node1199;
	wire [14-1:0] node1200;
	wire [14-1:0] node1203;
	wire [14-1:0] node1207;
	wire [14-1:0] node1208;
	wire [14-1:0] node1209;
	wire [14-1:0] node1210;
	wire [14-1:0] node1213;
	wire [14-1:0] node1215;
	wire [14-1:0] node1218;
	wire [14-1:0] node1219;
	wire [14-1:0] node1220;
	wire [14-1:0] node1223;
	wire [14-1:0] node1226;
	wire [14-1:0] node1228;
	wire [14-1:0] node1231;
	wire [14-1:0] node1232;
	wire [14-1:0] node1233;
	wire [14-1:0] node1235;
	wire [14-1:0] node1238;
	wire [14-1:0] node1239;
	wire [14-1:0] node1244;
	wire [14-1:0] node1245;
	wire [14-1:0] node1246;
	wire [14-1:0] node1247;
	wire [14-1:0] node1248;
	wire [14-1:0] node1249;
	wire [14-1:0] node1250;
	wire [14-1:0] node1253;
	wire [14-1:0] node1254;
	wire [14-1:0] node1257;
	wire [14-1:0] node1260;
	wire [14-1:0] node1261;
	wire [14-1:0] node1265;
	wire [14-1:0] node1266;
	wire [14-1:0] node1267;
	wire [14-1:0] node1270;
	wire [14-1:0] node1273;
	wire [14-1:0] node1274;
	wire [14-1:0] node1277;
	wire [14-1:0] node1278;
	wire [14-1:0] node1281;
	wire [14-1:0] node1284;
	wire [14-1:0] node1285;
	wire [14-1:0] node1286;
	wire [14-1:0] node1287;
	wire [14-1:0] node1290;
	wire [14-1:0] node1293;
	wire [14-1:0] node1294;
	wire [14-1:0] node1297;
	wire [14-1:0] node1300;
	wire [14-1:0] node1301;
	wire [14-1:0] node1305;
	wire [14-1:0] node1306;
	wire [14-1:0] node1308;
	wire [14-1:0] node1309;
	wire [14-1:0] node1310;
	wire [14-1:0] node1311;
	wire [14-1:0] node1315;
	wire [14-1:0] node1318;
	wire [14-1:0] node1319;
	wire [14-1:0] node1321;
	wire [14-1:0] node1326;
	wire [14-1:0] node1327;
	wire [14-1:0] node1328;
	wire [14-1:0] node1329;
	wire [14-1:0] node1331;
	wire [14-1:0] node1337;
	wire [14-1:0] node1338;
	wire [14-1:0] node1339;
	wire [14-1:0] node1340;
	wire [14-1:0] node1341;
	wire [14-1:0] node1342;
	wire [14-1:0] node1343;
	wire [14-1:0] node1345;
	wire [14-1:0] node1351;
	wire [14-1:0] node1352;
	wire [14-1:0] node1353;
	wire [14-1:0] node1354;
	wire [14-1:0] node1355;
	wire [14-1:0] node1359;
	wire [14-1:0] node1360;
	wire [14-1:0] node1362;
	wire [14-1:0] node1366;
	wire [14-1:0] node1367;
	wire [14-1:0] node1368;
	wire [14-1:0] node1371;
	wire [14-1:0] node1374;
	wire [14-1:0] node1375;
	wire [14-1:0] node1376;
	wire [14-1:0] node1381;
	wire [14-1:0] node1382;
	wire [14-1:0] node1383;
	wire [14-1:0] node1384;
	wire [14-1:0] node1387;
	wire [14-1:0] node1388;
	wire [14-1:0] node1392;
	wire [14-1:0] node1396;
	wire [14-1:0] node1398;
	wire [14-1:0] node1399;
	wire [14-1:0] node1400;
	wire [14-1:0] node1401;
	wire [14-1:0] node1405;
	wire [14-1:0] node1407;
	wire [14-1:0] node1408;
	wire [14-1:0] node1414;
	wire [14-1:0] node1415;
	wire [14-1:0] node1416;
	wire [14-1:0] node1417;
	wire [14-1:0] node1418;
	wire [14-1:0] node1419;
	wire [14-1:0] node1420;
	wire [14-1:0] node1421;
	wire [14-1:0] node1423;
	wire [14-1:0] node1425;
	wire [14-1:0] node1426;
	wire [14-1:0] node1430;
	wire [14-1:0] node1431;
	wire [14-1:0] node1432;
	wire [14-1:0] node1433;
	wire [14-1:0] node1435;
	wire [14-1:0] node1439;
	wire [14-1:0] node1442;
	wire [14-1:0] node1443;
	wire [14-1:0] node1447;
	wire [14-1:0] node1448;
	wire [14-1:0] node1449;
	wire [14-1:0] node1450;
	wire [14-1:0] node1453;
	wire [14-1:0] node1456;
	wire [14-1:0] node1458;
	wire [14-1:0] node1461;
	wire [14-1:0] node1462;
	wire [14-1:0] node1463;
	wire [14-1:0] node1468;
	wire [14-1:0] node1469;
	wire [14-1:0] node1470;
	wire [14-1:0] node1472;
	wire [14-1:0] node1473;
	wire [14-1:0] node1477;
	wire [14-1:0] node1478;
	wire [14-1:0] node1479;
	wire [14-1:0] node1484;
	wire [14-1:0] node1485;
	wire [14-1:0] node1486;
	wire [14-1:0] node1487;
	wire [14-1:0] node1491;
	wire [14-1:0] node1493;
	wire [14-1:0] node1496;
	wire [14-1:0] node1499;
	wire [14-1:0] node1500;
	wire [14-1:0] node1501;
	wire [14-1:0] node1502;
	wire [14-1:0] node1503;
	wire [14-1:0] node1504;
	wire [14-1:0] node1507;
	wire [14-1:0] node1511;
	wire [14-1:0] node1512;
	wire [14-1:0] node1515;
	wire [14-1:0] node1516;
	wire [14-1:0] node1519;
	wire [14-1:0] node1522;
	wire [14-1:0] node1523;
	wire [14-1:0] node1524;
	wire [14-1:0] node1529;
	wire [14-1:0] node1530;
	wire [14-1:0] node1531;
	wire [14-1:0] node1532;
	wire [14-1:0] node1533;
	wire [14-1:0] node1538;
	wire [14-1:0] node1540;
	wire [14-1:0] node1544;
	wire [14-1:0] node1545;
	wire [14-1:0] node1546;
	wire [14-1:0] node1547;
	wire [14-1:0] node1548;
	wire [14-1:0] node1549;
	wire [14-1:0] node1550;
	wire [14-1:0] node1553;
	wire [14-1:0] node1554;
	wire [14-1:0] node1558;
	wire [14-1:0] node1559;
	wire [14-1:0] node1562;
	wire [14-1:0] node1564;
	wire [14-1:0] node1567;
	wire [14-1:0] node1568;
	wire [14-1:0] node1572;
	wire [14-1:0] node1573;
	wire [14-1:0] node1574;
	wire [14-1:0] node1575;
	wire [14-1:0] node1576;
	wire [14-1:0] node1580;
	wire [14-1:0] node1584;
	wire [14-1:0] node1585;
	wire [14-1:0] node1586;
	wire [14-1:0] node1591;
	wire [14-1:0] node1592;
	wire [14-1:0] node1594;
	wire [14-1:0] node1595;
	wire [14-1:0] node1599;
	wire [14-1:0] node1600;
	wire [14-1:0] node1601;
	wire [14-1:0] node1602;
	wire [14-1:0] node1606;
	wire [14-1:0] node1611;
	wire [14-1:0] node1612;
	wire [14-1:0] node1613;
	wire [14-1:0] node1614;
	wire [14-1:0] node1615;
	wire [14-1:0] node1616;
	wire [14-1:0] node1617;
	wire [14-1:0] node1618;
	wire [14-1:0] node1620;
	wire [14-1:0] node1623;
	wire [14-1:0] node1624;
	wire [14-1:0] node1628;
	wire [14-1:0] node1629;
	wire [14-1:0] node1631;
	wire [14-1:0] node1632;
	wire [14-1:0] node1636;
	wire [14-1:0] node1639;
	wire [14-1:0] node1640;
	wire [14-1:0] node1641;
	wire [14-1:0] node1645;
	wire [14-1:0] node1646;
	wire [14-1:0] node1647;
	wire [14-1:0] node1652;
	wire [14-1:0] node1653;
	wire [14-1:0] node1654;
	wire [14-1:0] node1655;
	wire [14-1:0] node1658;
	wire [14-1:0] node1660;
	wire [14-1:0] node1663;
	wire [14-1:0] node1667;
	wire [14-1:0] node1669;
	wire [14-1:0] node1670;
	wire [14-1:0] node1671;
	wire [14-1:0] node1674;
	wire [14-1:0] node1677;
	wire [14-1:0] node1678;
	wire [14-1:0] node1680;
	wire [14-1:0] node1684;
	wire [14-1:0] node1685;
	wire [14-1:0] node1687;
	wire [14-1:0] node1688;
	wire [14-1:0] node1689;
	wire [14-1:0] node1692;
	wire [14-1:0] node1695;
	wire [14-1:0] node1696;
	wire [14-1:0] node1698;
	wire [14-1:0] node1699;
	wire [14-1:0] node1705;
	wire [14-1:0] node1706;
	wire [14-1:0] node1707;
	wire [14-1:0] node1708;
	wire [14-1:0] node1709;
	wire [14-1:0] node1711;
	wire [14-1:0] node1713;
	wire [14-1:0] node1715;
	wire [14-1:0] node1718;
	wire [14-1:0] node1719;
	wire [14-1:0] node1726;
	wire [14-1:0] node1728;
	wire [14-1:0] node1729;
	wire [14-1:0] node1730;
	wire [14-1:0] node1731;
	wire [14-1:0] node1732;
	wire [14-1:0] node1733;
	wire [14-1:0] node1734;
	wire [14-1:0] node1736;
	wire [14-1:0] node1739;
	wire [14-1:0] node1741;
	wire [14-1:0] node1744;
	wire [14-1:0] node1745;
	wire [14-1:0] node1748;
	wire [14-1:0] node1750;
	wire [14-1:0] node1753;
	wire [14-1:0] node1754;
	wire [14-1:0] node1755;
	wire [14-1:0] node1758;
	wire [14-1:0] node1762;
	wire [14-1:0] node1763;
	wire [14-1:0] node1764;
	wire [14-1:0] node1765;
	wire [14-1:0] node1771;
	wire [14-1:0] node1773;
	wire [14-1:0] node1774;
	wire [14-1:0] node1775;
	wire [14-1:0] node1776;
	wire [14-1:0] node1778;
	wire [14-1:0] node1781;
	wire [14-1:0] node1782;
	wire [14-1:0] node1788;
	wire [14-1:0] node1790;
	wire [14-1:0] node1792;
	wire [14-1:0] node1794;
	wire [14-1:0] node1796;
	wire [14-1:0] node1798;

	assign outp = (inp[8]) ? node604 : node1;
		assign node1 = (inp[13]) ? node3 : 14'b00000000000000;
			assign node3 = (inp[5]) ? node417 : node4;
				assign node4 = (inp[3]) ? node290 : node5;
					assign node5 = (inp[2]) ? node199 : node6;
						assign node6 = (inp[10]) ? node104 : node7;
							assign node7 = (inp[4]) ? node65 : node8;
								assign node8 = (inp[7]) ? node36 : node9;
									assign node9 = (inp[12]) ? node17 : node10;
										assign node10 = (inp[6]) ? 14'b00000000000001 : node11;
											assign node11 = (inp[1]) ? 14'b00000000000001 : node12;
												assign node12 = (inp[0]) ? 14'b00000000000001 : 14'b10000000001000;
										assign node17 = (inp[6]) ? node29 : node18;
											assign node18 = (inp[1]) ? node24 : node19;
												assign node19 = (inp[9]) ? node21 : 14'b00000000000001;
													assign node21 = (inp[11]) ? 14'b01000010010100 : 14'b01000000000100;
												assign node24 = (inp[0]) ? 14'b00000000000001 : node25;
													assign node25 = (inp[11]) ? 14'b01010010100100 : 14'b01010010000100;
											assign node29 = (inp[0]) ? node33 : node30;
												assign node30 = (inp[9]) ? 14'b01010000010100 : 14'b01010000110100;
												assign node33 = (inp[9]) ? 14'b01000000010100 : 14'b01000000110100;
									assign node36 = (inp[12]) ? node50 : node37;
										assign node37 = (inp[0]) ? node47 : node38;
											assign node38 = (inp[11]) ? node44 : node39;
												assign node39 = (inp[6]) ? 14'b00010000110010 : node40;
													assign node40 = (inp[9]) ? 14'b00010010000010 : 14'b00010010100010;
												assign node44 = (inp[9]) ? 14'b00010000000010 : 14'b00000000000001;
											assign node47 = (inp[9]) ? 14'b00000010010010 : 14'b00000010110010;
										assign node50 = (inp[1]) ? node62 : node51;
											assign node51 = (inp[6]) ? node57 : node52;
												assign node52 = (inp[0]) ? 14'b00000010110000 : node53;
													assign node53 = (inp[9]) ? 14'b00000000000000 : 14'b00000000000001;
												assign node57 = (inp[9]) ? node59 : 14'b00010000110000;
													assign node59 = (inp[0]) ? 14'b00000000010000 : 14'b00010000010000;
											assign node62 = (inp[9]) ? 14'b00010010000000 : 14'b00000000000001;
								assign node65 = (inp[0]) ? node97 : node66;
									assign node66 = (inp[6]) ? node82 : node67;
										assign node67 = (inp[1]) ? node75 : node68;
											assign node68 = (inp[9]) ? node70 : 14'b00000000000001;
												assign node70 = (inp[12]) ? node72 : 14'b00100000000110;
													assign node72 = (inp[7]) ? 14'b00100000000100 : 14'b00100100000100;
											assign node75 = (inp[7]) ? node79 : node76;
												assign node76 = (inp[11]) ? 14'b00110110100110 : 14'b00110110100100;
												assign node79 = (inp[9]) ? 14'b00110010000100 : 14'b00110010100100;
										assign node82 = (inp[9]) ? node90 : node83;
											assign node83 = (inp[12]) ? node87 : node84;
												assign node84 = (inp[7]) ? 14'b00110000110110 : 14'b00110100110110;
												assign node87 = (inp[1]) ? 14'b00110100100100 : 14'b00110100110100;
											assign node90 = (inp[7]) ? node94 : node91;
												assign node91 = (inp[12]) ? 14'b00110100010100 : 14'b00110100010110;
												assign node94 = (inp[1]) ? 14'b00110000000100 : 14'b00110000010100;
									assign node97 = (inp[1]) ? 14'b00000000000001 : node98;
										assign node98 = (inp[12]) ? 14'b00100100010100 : node99;
											assign node99 = (inp[7]) ? 14'b00100010010110 : 14'b00100110110110;
							assign node104 = (inp[1]) ? node168 : node105;
								assign node105 = (inp[12]) ? node137 : node106;
									assign node106 = (inp[6]) ? node116 : node107;
										assign node107 = (inp[9]) ? node111 : node108;
											assign node108 = (inp[7]) ? 14'b01100010110010 : 14'b00100110110010;
											assign node111 = (inp[4]) ? 14'b00100010010010 : node112;
												assign node112 = (inp[7]) ? 14'b01100010010010 : 14'b01100110010010;
										assign node116 = (inp[4]) ? node126 : node117;
											assign node117 = (inp[9]) ? node123 : node118;
												assign node118 = (inp[11]) ? node120 : 14'b01110000110010;
													assign node120 = (inp[0]) ? 14'b01100100110010 : 14'b01110100110010;
												assign node123 = (inp[0]) ? 14'b01100100010010 : 14'b01110100010010;
											assign node126 = (inp[0]) ? node130 : node127;
												assign node127 = (inp[9]) ? 14'b00110100010010 : 14'b00110100110010;
												assign node130 = (inp[7]) ? node134 : node131;
													assign node131 = (inp[9]) ? 14'b00100100010010 : 14'b00100100110010;
													assign node134 = (inp[9]) ? 14'b00100000010010 : 14'b00100000110010;
									assign node137 = (inp[0]) ? node151 : node138;
										assign node138 = (inp[6]) ? node144 : node139;
											assign node139 = (inp[9]) ? node141 : 14'b00000000000001;
												assign node141 = (inp[7]) ? 14'b01100000000000 : 14'b01100100000000;
											assign node144 = (inp[4]) ? node146 : 14'b01110000110000;
												assign node146 = (inp[7]) ? 14'b00110000010000 : node147;
													assign node147 = (inp[9]) ? 14'b00110100010000 : 14'b00110100110000;
										assign node151 = (inp[7]) ? node161 : node152;
											assign node152 = (inp[4]) ? node156 : node153;
												assign node153 = (inp[6]) ? 14'b01100100010000 : 14'b01100110010000;
												assign node156 = (inp[9]) ? node158 : 14'b00100110110000;
													assign node158 = (inp[6]) ? 14'b00100100010000 : 14'b00100110010000;
											assign node161 = (inp[6]) ? node165 : node162;
												assign node162 = (inp[9]) ? 14'b01100010010000 : 14'b01100010110000;
												assign node165 = (inp[9]) ? 14'b01100000010000 : 14'b01100000110000;
								assign node168 = (inp[0]) ? 14'b00000000000001 : node169;
									assign node169 = (inp[7]) ? node183 : node170;
										assign node170 = (inp[6]) ? node176 : node171;
											assign node171 = (inp[4]) ? node173 : 14'b01110110000000;
												assign node173 = (inp[9]) ? 14'b00110110000010 : 14'b00110110100000;
											assign node176 = (inp[4]) ? 14'b00110100100000 : node177;
												assign node177 = (inp[12]) ? node179 : 14'b01110100100010;
													assign node179 = (inp[9]) ? 14'b01110100000000 : 14'b01110100100000;
										assign node183 = (inp[9]) ? node189 : node184;
											assign node184 = (inp[6]) ? 14'b00110000100000 : node185;
												assign node185 = (inp[12]) ? 14'b01110010100000 : 14'b01110010100010;
											assign node189 = (inp[12]) ? node193 : node190;
												assign node190 = (inp[11]) ? 14'b01110000000010 : 14'b00110000000010;
												assign node193 = (inp[6]) ? node195 : 14'b00110010000000;
													assign node195 = (inp[4]) ? 14'b00110000000000 : 14'b01110000000000;
						assign node199 = (inp[10]) ? node269 : node200;
							assign node200 = (inp[4]) ? node246 : node201;
								assign node201 = (inp[0]) ? node229 : node202;
									assign node202 = (inp[9]) ? node218 : node203;
										assign node203 = (inp[12]) ? node211 : node204;
											assign node204 = (inp[7]) ? node206 : 14'b01110100100110;
												assign node206 = (inp[6]) ? node208 : 14'b01110010100110;
													assign node208 = (inp[1]) ? 14'b01110000100110 : 14'b01110000110110;
											assign node211 = (inp[1]) ? node215 : node212;
												assign node212 = (inp[7]) ? 14'b01110000110100 : 14'b01110100110100;
												assign node215 = (inp[7]) ? 14'b01110000100100 : 14'b01110100100100;
										assign node218 = (inp[12]) ? node226 : node219;
											assign node219 = (inp[1]) ? node223 : node220;
												assign node220 = (inp[7]) ? 14'b01110000010110 : 14'b01110100010110;
												assign node223 = (inp[7]) ? 14'b01110000000110 : 14'b01110100000110;
											assign node226 = (inp[1]) ? 14'b01110010000100 : 14'b01100000000100;
									assign node229 = (inp[1]) ? 14'b00000000000001 : node230;
										assign node230 = (inp[12]) ? node234 : node231;
											assign node231 = (inp[9]) ? 14'b01100110010110 : 14'b01100110110110;
											assign node234 = (inp[7]) ? node240 : node235;
												assign node235 = (inp[6]) ? node237 : 14'b01100110010100;
													assign node237 = (inp[11]) ? 14'b01100100110100 : 14'b01100100010100;
												assign node240 = (inp[11]) ? 14'b01100000010100 : node241;
													assign node241 = (inp[9]) ? 14'b01100010010100 : 14'b01100010110100;
								assign node246 = (inp[7]) ? 14'b00000000000001 : node247;
									assign node247 = (inp[12]) ? node249 : 14'b00000000000001;
										assign node249 = (inp[1]) ? node263 : node250;
											assign node250 = (inp[6]) ? node256 : node251;
												assign node251 = (inp[0]) ? 14'b00000110110100 : node252;
													assign node252 = (inp[9]) ? 14'b00000100000100 : 14'b00000000000001;
												assign node256 = (inp[9]) ? node260 : node257;
													assign node257 = (inp[0]) ? 14'b00000100110100 : 14'b00010100110100;
													assign node260 = (inp[11]) ? 14'b00000100010100 : 14'b00010100010100;
											assign node263 = (inp[0]) ? 14'b00000000000001 : node264;
												assign node264 = (inp[6]) ? 14'b00010100000100 : 14'b00010110000100;
							assign node269 = (inp[4]) ? node271 : 14'b00000000000001;
								assign node271 = (inp[7]) ? 14'b00000000000001 : node272;
									assign node272 = (inp[1]) ? node282 : node273;
										assign node273 = (inp[6]) ? node277 : node274;
											assign node274 = (inp[9]) ? 14'b00000100000000 : 14'b00000000000001;
											assign node277 = (inp[12]) ? 14'b00010100110000 : node278;
												assign node278 = (inp[0]) ? 14'b00000100010010 : 14'b00010100010010;
										assign node282 = (inp[12]) ? node286 : node283;
											assign node283 = (inp[6]) ? 14'b00010100100010 : 14'b00010110100010;
											assign node286 = (inp[9]) ? 14'b00010100000000 : 14'b00010110100000;
					assign node290 = (inp[0]) ? node392 : node291;
						assign node291 = (inp[6]) ? node379 : node292;
							assign node292 = (inp[2]) ? node354 : node293;
								assign node293 = (inp[1]) ? node323 : node294;
									assign node294 = (inp[4]) ? node306 : node295;
										assign node295 = (inp[10]) ? node297 : 14'b00010010010000;
											assign node297 = (inp[7]) ? node303 : node298;
												assign node298 = (inp[12]) ? node300 : 14'b01110110010010;
													assign node300 = (inp[11]) ? 14'b01110110110000 : 14'b01110110010000;
												assign node303 = (inp[12]) ? 14'b01110010110000 : 14'b01110010110010;
										assign node306 = (inp[9]) ? node316 : node307;
											assign node307 = (inp[7]) ? node313 : node308;
												assign node308 = (inp[12]) ? 14'b00110110110100 : node309;
													assign node309 = (inp[10]) ? 14'b00110110110010 : 14'b00110110110110;
												assign node313 = (inp[10]) ? 14'b00110010110010 : 14'b00110010110110;
											assign node316 = (inp[10]) ? 14'b00110110010010 : node317;
												assign node317 = (inp[7]) ? 14'b00110010010110 : node318;
													assign node318 = (inp[11]) ? 14'b00110110010100 : 14'b00110110010110;
									assign node323 = (inp[10]) ? node335 : node324;
										assign node324 = (inp[4]) ? node330 : node325;
											assign node325 = (inp[12]) ? node327 : 14'b00000000000001;
												assign node327 = (inp[7]) ? 14'b00000010000000 : 14'b01000010100100;
											assign node330 = (inp[12]) ? node332 : 14'b00100110100110;
												assign node332 = (inp[11]) ? 14'b00100010000100 : 14'b00100010100100;
										assign node335 = (inp[7]) ? node345 : node336;
											assign node336 = (inp[12]) ? node340 : node337;
												assign node337 = (inp[11]) ? 14'b00100110000010 : 14'b01100110000010;
												assign node340 = (inp[4]) ? 14'b00100110000000 : node341;
													assign node341 = (inp[9]) ? 14'b01100110000000 : 14'b01100110100000;
											assign node345 = (inp[12]) ? node351 : node346;
												assign node346 = (inp[9]) ? 14'b00100010000010 : node347;
													assign node347 = (inp[11]) ? 14'b00100010100010 : 14'b01100010100010;
												assign node351 = (inp[11]) ? 14'b00100010100000 : 14'b00100010000000;
								assign node354 = (inp[10]) ? node368 : node355;
									assign node355 = (inp[4]) ? 14'b00000000000001 : node356;
										assign node356 = (inp[1]) ? node362 : node357;
											assign node357 = (inp[7]) ? node359 : 14'b01110110110100;
												assign node359 = (inp[11]) ? 14'b01110010010110 : 14'b01110010010100;
											assign node362 = (inp[9]) ? 14'b01100110000100 : node363;
												assign node363 = (inp[7]) ? 14'b01100010100100 : 14'b01100110100100;
									assign node368 = (inp[4]) ? node370 : 14'b00000000000001;
										assign node370 = (inp[7]) ? 14'b00000000000001 : node371;
											assign node371 = (inp[1]) ? node375 : node372;
												assign node372 = (inp[11]) ? 14'b00010110110010 : 14'b00010110110000;
												assign node375 = (inp[12]) ? 14'b00000110000000 : 14'b00000110100010;
							assign node379 = (inp[2]) ? node381 : 14'b00000000000001;
								assign node381 = (inp[11]) ? 14'b00000000000001 : node382;
									assign node382 = (inp[12]) ? 14'b00000000000001 : node383;
										assign node383 = (inp[4]) ? 14'b10000001001010 : node384;
											assign node384 = (inp[1]) ? 14'b00000000000001 : node385;
												assign node385 = (inp[7]) ? 14'b00000000000001 : 14'b10000001001000;
						assign node392 = (inp[9]) ? 14'b00000000000001 : node393;
							assign node393 = (inp[1]) ? 14'b00000000000001 : node394;
								assign node394 = (inp[6]) ? node396 : 14'b00000000000001;
									assign node396 = (inp[10]) ? node412 : node397;
										assign node397 = (inp[12]) ? node403 : node398;
											assign node398 = (inp[4]) ? 14'b00100100100110 : node399;
												assign node399 = (inp[7]) ? 14'b00000000100010 : 14'b00000000000001;
											assign node403 = (inp[2]) ? node409 : node404;
												assign node404 = (inp[4]) ? 14'b00100000100100 : node405;
													assign node405 = (inp[7]) ? 14'b00000000100000 : 14'b01000000100100;
												assign node409 = (inp[11]) ? 14'b01100000100100 : 14'b01100100100100;
										assign node412 = (inp[4]) ? 14'b00100000100000 : 14'b00000000000001;
				assign node417 = (inp[10]) ? 14'b00000000000001 : node418;
					assign node418 = (inp[12]) ? node524 : node419;
						assign node419 = (inp[0]) ? node489 : node420;
							assign node420 = (inp[7]) ? node468 : node421;
								assign node421 = (inp[1]) ? node439 : node422;
									assign node422 = (inp[3]) ? node430 : node423;
										assign node423 = (inp[9]) ? node427 : node424;
											assign node424 = (inp[6]) ? 14'b01010100110010 : 14'b00000000000001;
											assign node427 = (inp[4]) ? 14'b01000000000010 : 14'b01000100000010;
										assign node430 = (inp[6]) ? 14'b00000000000001 : node431;
											assign node431 = (inp[4]) ? 14'b01010010010010 : node432;
												assign node432 = (inp[2]) ? 14'b01010110110010 : node433;
													assign node433 = (inp[9]) ? 14'b01010110010110 : 14'b01010110110110;
									assign node439 = (inp[2]) ? node457 : node440;
										assign node440 = (inp[3]) ? node454 : node441;
											assign node441 = (inp[9]) ? node447 : node442;
												assign node442 = (inp[6]) ? node444 : 14'b00010110100110;
													assign node444 = (inp[4]) ? 14'b00010100100110 : 14'b01010100100110;
												assign node447 = (inp[4]) ? node451 : node448;
													assign node448 = (inp[6]) ? 14'b01010100000110 : 14'b01010110000110;
													assign node451 = (inp[11]) ? 14'b00010110000110 : 14'b00010100000110;
											assign node454 = (inp[4]) ? 14'b00000000000001 : 14'b01000110000110;
										assign node457 = (inp[9]) ? node465 : node458;
											assign node458 = (inp[3]) ? node462 : node459;
												assign node459 = (inp[4]) ? 14'b01010000100010 : 14'b01010100100010;
												assign node462 = (inp[11]) ? 14'b01000010100010 : 14'b01000110100010;
											assign node465 = (inp[6]) ? 14'b01010100000010 : 14'b01010110000010;
								assign node468 = (inp[2]) ? 14'b00000000000001 : node469;
									assign node469 = (inp[3]) ? node481 : node470;
										assign node470 = (inp[6]) ? node474 : node471;
											assign node471 = (inp[4]) ? 14'b00010010100110 : 14'b00000000000001;
											assign node474 = (inp[4]) ? node478 : node475;
												assign node475 = (inp[1]) ? 14'b01010000100110 : 14'b01010000110110;
												assign node478 = (inp[11]) ? 14'b00010000100110 : 14'b00010000000110;
										assign node481 = (inp[6]) ? 14'b00000000000001 : node482;
											assign node482 = (inp[1]) ? node484 : 14'b00010010110110;
												assign node484 = (inp[4]) ? 14'b00000010000110 : 14'b01000010100110;
							assign node489 = (inp[1]) ? 14'b00000000000001 : node490;
								assign node490 = (inp[3]) ? node512 : node491;
									assign node491 = (inp[7]) ? node505 : node492;
										assign node492 = (inp[2]) ? node496 : node493;
											assign node493 = (inp[9]) ? 14'b00000100010110 : 14'b00000110110110;
											assign node496 = (inp[4]) ? node500 : node497;
												assign node497 = (inp[6]) ? 14'b01000100010010 : 14'b01000110010010;
												assign node500 = (inp[9]) ? 14'b01000010010010 : node501;
													assign node501 = (inp[6]) ? 14'b01000000110010 : 14'b01000010110010;
										assign node505 = (inp[2]) ? 14'b00000000000001 : node506;
											assign node506 = (inp[11]) ? 14'b01000000010110 : node507;
												assign node507 = (inp[9]) ? 14'b00000010010110 : 14'b00000010110110;
									assign node512 = (inp[9]) ? 14'b00000000000001 : node513;
										assign node513 = (inp[7]) ? node517 : node514;
											assign node514 = (inp[4]) ? 14'b01000000100010 : 14'b01000100100010;
											assign node517 = (inp[2]) ? 14'b00000000000001 : node518;
												assign node518 = (inp[4]) ? 14'b00000000100110 : 14'b01000000100110;
						assign node524 = (inp[4]) ? node576 : node525;
							assign node525 = (inp[7]) ? node559 : node526;
								assign node526 = (inp[0]) ? node548 : node527;
									assign node527 = (inp[6]) ? node541 : node528;
										assign node528 = (inp[2]) ? node536 : node529;
											assign node529 = (inp[9]) ? node531 : 14'b01010110110100;
												assign node531 = (inp[1]) ? node533 : 14'b01000100000100;
													assign node533 = (inp[3]) ? 14'b01000110000100 : 14'b01010110000100;
											assign node536 = (inp[9]) ? 14'b01010110010000 : node537;
												assign node537 = (inp[3]) ? 14'b01000110100000 : 14'b01010110100000;
										assign node541 = (inp[3]) ? 14'b00000000000001 : node542;
											assign node542 = (inp[2]) ? node544 : 14'b01010100110100;
												assign node544 = (inp[1]) ? 14'b01010100000000 : 14'b01010100010000;
									assign node548 = (inp[1]) ? 14'b00000000000001 : node549;
										assign node549 = (inp[3]) ? node555 : node550;
											assign node550 = (inp[6]) ? node552 : 14'b01000110010100;
												assign node552 = (inp[9]) ? 14'b01000100010100 : 14'b01000100110100;
											assign node555 = (inp[6]) ? 14'b01000100100000 : 14'b00000000000001;
								assign node559 = (inp[2]) ? node561 : 14'b00000000000001;
									assign node561 = (inp[1]) ? node567 : node562;
										assign node562 = (inp[3]) ? node564 : 14'b01000010110000;
											assign node564 = (inp[9]) ? 14'b01010010010000 : 14'b01010010110000;
										assign node567 = (inp[0]) ? 14'b00000000000001 : node568;
											assign node568 = (inp[11]) ? node572 : node569;
												assign node569 = (inp[6]) ? 14'b01010000000000 : 14'b01010010000000;
												assign node572 = (inp[6]) ? 14'b00000000000001 : 14'b01000010000000;
							assign node576 = (inp[2]) ? 14'b00000000000001 : node577;
								assign node577 = (inp[7]) ? node579 : 14'b00000000000001;
									assign node579 = (inp[1]) ? node597 : node580;
										assign node580 = (inp[6]) ? node590 : node581;
											assign node581 = (inp[3]) ? 14'b00010010110100 : node582;
												assign node582 = (inp[0]) ? node586 : node583;
													assign node583 = (inp[11]) ? 14'b00000000000100 : 14'b00000000000001;
													assign node586 = (inp[9]) ? 14'b00000010010100 : 14'b00000010110100;
											assign node590 = (inp[3]) ? node592 : 14'b00010000110100;
												assign node592 = (inp[11]) ? node594 : 14'b00000000000001;
													assign node594 = (inp[0]) ? 14'b00000000100100 : 14'b00000000000001;
										assign node597 = (inp[0]) ? 14'b00000000000001 : node598;
											assign node598 = (inp[11]) ? 14'b00000010000100 : 14'b00000000000001;
		assign node604 = (inp[0]) ? node1414 : node605;
			assign node605 = (inp[2]) ? node1083 : node606;
				assign node606 = (inp[12]) ? node892 : node607;
					assign node607 = (inp[3]) ? node781 : node608;
						assign node608 = (inp[6]) ? node686 : node609;
							assign node609 = (inp[1]) ? node643 : node610;
								assign node610 = (inp[9]) ? node624 : node611;
									assign node611 = (inp[13]) ? 14'b00000000000001 : node612;
										assign node612 = (inp[5]) ? node618 : node613;
											assign node613 = (inp[4]) ? 14'b00000000000001 : node614;
												assign node614 = (inp[10]) ? 14'b00000000000001 : 14'b10000000001000;
											assign node618 = (inp[11]) ? 14'b00000000000001 : node619;
												assign node619 = (inp[4]) ? 14'b01100110110000 : 14'b00100110110010;
									assign node624 = (inp[13]) ? node634 : node625;
										assign node625 = (inp[10]) ? node629 : node626;
											assign node626 = (inp[4]) ? 14'b01101110010110 : 14'b01100110010100;
											assign node629 = (inp[11]) ? 14'b00000000000001 : node630;
												assign node630 = (inp[5]) ? 14'b01100100000000 : 14'b01101100000000;
										assign node634 = (inp[7]) ? node636 : 14'b00100100000000;
											assign node636 = (inp[4]) ? node640 : node637;
												assign node637 = (inp[5]) ? 14'b01100000000000 : 14'b00000000000000;
												assign node640 = (inp[5]) ? 14'b00100000000000 : 14'b00100000000100;
								assign node643 = (inp[13]) ? node663 : node644;
									assign node644 = (inp[10]) ? node656 : node645;
										assign node645 = (inp[11]) ? node651 : node646;
											assign node646 = (inp[4]) ? 14'b01101010010110 : node647;
												assign node647 = (inp[5]) ? 14'b00100000000010 : 14'b00000000000001;
											assign node651 = (inp[7]) ? 14'b01100010010100 : node652;
												assign node652 = (inp[9]) ? 14'b01101000000100 : 14'b01111010000100;
										assign node656 = (inp[11]) ? 14'b00000000000001 : node657;
											assign node657 = (inp[7]) ? 14'b01101010110000 : node658;
												assign node658 = (inp[9]) ? 14'b01100000000000 : 14'b01110010000010;
									assign node663 = (inp[4]) ? node677 : node664;
										assign node664 = (inp[5]) ? node670 : node665;
											assign node665 = (inp[7]) ? node667 : 14'b00000000000001;
												assign node667 = (inp[9]) ? 14'b00010010000000 : 14'b00010010100000;
											assign node670 = (inp[9]) ? node674 : node671;
												assign node671 = (inp[7]) ? 14'b01110010100000 : 14'b01110110100000;
												assign node674 = (inp[7]) ? 14'b01110010000000 : 14'b01110110000000;
										assign node677 = (inp[7]) ? node683 : node678;
											assign node678 = (inp[5]) ? node680 : 14'b00110110100100;
												assign node680 = (inp[9]) ? 14'b00110110000000 : 14'b00110110100000;
											assign node683 = (inp[9]) ? 14'b00110010000100 : 14'b00110010100100;
							assign node686 = (inp[5]) ? node726 : node687;
								assign node687 = (inp[4]) ? node703 : node688;
									assign node688 = (inp[7]) ? node694 : node689;
										assign node689 = (inp[13]) ? 14'b00000000000001 : node690;
											assign node690 = (inp[1]) ? 14'b00000000000001 : 14'b01111100010100;
										assign node694 = (inp[13]) ? node696 : 14'b00000000000001;
											assign node696 = (inp[9]) ? node700 : node697;
												assign node697 = (inp[1]) ? 14'b00010000100000 : 14'b00010000110000;
												assign node700 = (inp[1]) ? 14'b00010000000000 : 14'b00010000010000;
									assign node703 = (inp[11]) ? node719 : node704;
										assign node704 = (inp[13]) ? node712 : node705;
											assign node705 = (inp[10]) ? node709 : node706;
												assign node706 = (inp[1]) ? 14'b01101000110110 : 14'b01101100110110;
												assign node709 = (inp[9]) ? 14'b01111100010000 : 14'b01111100110000;
											assign node712 = (inp[1]) ? 14'b00110100000100 : node713;
												assign node713 = (inp[9]) ? 14'b00110000010100 : node714;
													assign node714 = (inp[10]) ? 14'b00110000110100 : 14'b00110100110100;
										assign node719 = (inp[13]) ? node721 : 14'b00000000000001;
											assign node721 = (inp[7]) ? 14'b00110000000100 : node722;
												assign node722 = (inp[1]) ? 14'b00110100100100 : 14'b00110100010100;
								assign node726 = (inp[9]) ? node756 : node727;
									assign node727 = (inp[7]) ? node743 : node728;
										assign node728 = (inp[1]) ? node738 : node729;
											assign node729 = (inp[10]) ? node733 : node730;
												assign node730 = (inp[4]) ? 14'b00110100110000 : 14'b01110100110000;
												assign node733 = (inp[13]) ? 14'b01110100110000 : node734;
													assign node734 = (inp[4]) ? 14'b01110100110000 : 14'b01110100110010;
											assign node738 = (inp[13]) ? node740 : 14'b01110000110000;
												assign node740 = (inp[4]) ? 14'b00110100100000 : 14'b01110100100000;
										assign node743 = (inp[13]) ? node749 : node744;
											assign node744 = (inp[1]) ? node746 : 14'b01100100110110;
												assign node746 = (inp[4]) ? 14'b01100000110000 : 14'b00100000110010;
											assign node749 = (inp[1]) ? node753 : node750;
												assign node750 = (inp[4]) ? 14'b00110000110000 : 14'b01110000110000;
												assign node753 = (inp[4]) ? 14'b00110000100000 : 14'b01110000100000;
									assign node756 = (inp[11]) ? node772 : node757;
										assign node757 = (inp[10]) ? node767 : node758;
											assign node758 = (inp[4]) ? node762 : node759;
												assign node759 = (inp[1]) ? 14'b00110000010010 : 14'b00110100010010;
												assign node762 = (inp[1]) ? node764 : 14'b01100100010110;
													assign node764 = (inp[7]) ? 14'b01100000010110 : 14'b01110000010110;
											assign node767 = (inp[1]) ? 14'b00110100000000 : node768;
												assign node768 = (inp[7]) ? 14'b01100100010000 : 14'b01110100010000;
										assign node772 = (inp[13]) ? node774 : 14'b00000000000001;
											assign node774 = (inp[4]) ? 14'b00110000000000 : node775;
												assign node775 = (inp[7]) ? 14'b01110000010000 : node776;
													assign node776 = (inp[10]) ? 14'b01110100000000 : 14'b01110100010000;
						assign node781 = (inp[6]) ? node869 : node782;
							assign node782 = (inp[9]) ? node832 : node783;
								assign node783 = (inp[5]) ? node807 : node784;
									assign node784 = (inp[4]) ? node800 : node785;
										assign node785 = (inp[1]) ? node791 : node786;
											assign node786 = (inp[7]) ? node788 : 14'b00000000000001;
												assign node788 = (inp[13]) ? 14'b00010010110000 : 14'b00000000000001;
											assign node791 = (inp[11]) ? 14'b01111010110100 : node792;
												assign node792 = (inp[10]) ? node794 : 14'b00000010100000;
													assign node794 = (inp[13]) ? 14'b00000000000001 : node795;
														assign node795 = (inp[7]) ? 14'b00000000000001 : 14'b01111010110010;
										assign node800 = (inp[13]) ? node802 : 14'b00000000000001;
											assign node802 = (inp[1]) ? node804 : 14'b00110110110100;
												assign node804 = (inp[7]) ? 14'b00100010100100 : 14'b00100110100100;
									assign node807 = (inp[11]) ? node821 : node808;
										assign node808 = (inp[10]) ? node812 : node809;
											assign node809 = (inp[7]) ? 14'b00110010110000 : 14'b01110010110110;
											assign node812 = (inp[13]) ? node818 : node813;
												assign node813 = (inp[4]) ? 14'b01110110110000 : node814;
													assign node814 = (inp[1]) ? 14'b01110010110010 : 14'b01110110110010;
												assign node818 = (inp[1]) ? 14'b01100110100000 : 14'b01110110110000;
										assign node821 = (inp[13]) ? node823 : 14'b00000000000001;
											assign node823 = (inp[1]) ? node829 : node824;
												assign node824 = (inp[4]) ? node826 : 14'b01110010110000;
													assign node826 = (inp[7]) ? 14'b00110010110000 : 14'b00110110110000;
												assign node829 = (inp[4]) ? 14'b00100010100000 : 14'b01100110100000;
								assign node832 = (inp[13]) ? node852 : node833;
									assign node833 = (inp[7]) ? 14'b00000000000001 : node834;
										assign node834 = (inp[11]) ? node844 : node835;
											assign node835 = (inp[10]) ? node839 : node836;
												assign node836 = (inp[5]) ? 14'b01110110010110 : 14'b01111110010110;
												assign node839 = (inp[4]) ? node841 : 14'b01110110010010;
													assign node841 = (inp[5]) ? 14'b01110010010000 : 14'b01111110010000;
											assign node844 = (inp[4]) ? 14'b00000000000001 : node845;
												assign node845 = (inp[5]) ? node847 : 14'b00000000000001;
													assign node847 = (inp[1]) ? 14'b01110010010100 : 14'b01110110010100;
									assign node852 = (inp[4]) ? node860 : node853;
										assign node853 = (inp[7]) ? node855 : 14'b00000000000001;
											assign node855 = (inp[11]) ? node857 : 14'b00000010000000;
												assign node857 = (inp[5]) ? 14'b01110010010000 : 14'b00010010010000;
										assign node860 = (inp[1]) ? node866 : node861;
											assign node861 = (inp[7]) ? node863 : 14'b00110110010100;
												assign node863 = (inp[10]) ? 14'b00110010010100 : 14'b00110010010000;
											assign node866 = (inp[5]) ? 14'b00100010000000 : 14'b00100010000100;
							assign node869 = (inp[13]) ? 14'b00000000000001 : node870;
								assign node870 = (inp[9]) ? 14'b00000000000001 : node871;
									assign node871 = (inp[7]) ? node879 : node872;
										assign node872 = (inp[1]) ? node874 : 14'b00000000000001;
											assign node874 = (inp[11]) ? node876 : 14'b00000000000001;
												assign node876 = (inp[5]) ? 14'b01110000100100 : 14'b01111000100100;
										assign node879 = (inp[11]) ? 14'b00000000000001 : node880;
											assign node880 = (inp[5]) ? node884 : node881;
												assign node881 = (inp[10]) ? 14'b01101000100000 : 14'b00000000000001;
												assign node884 = (inp[10]) ? node886 : 14'b01100100100110;
													assign node886 = (inp[1]) ? 14'b01100000100010 : 14'b01100100100010;
					assign node892 = (inp[5]) ? node1032 : node893;
						assign node893 = (inp[13]) ? node971 : node894;
							assign node894 = (inp[3]) ? node942 : node895;
								assign node895 = (inp[10]) ? node925 : node896;
									assign node896 = (inp[11]) ? node906 : node897;
										assign node897 = (inp[6]) ? node899 : 14'b00000000000001;
											assign node899 = (inp[4]) ? 14'b00000000000001 : node900;
												assign node900 = (inp[9]) ? node902 : 14'b01001000110110;
													assign node902 = (inp[1]) ? 14'b01011000010110 : 14'b01011100010110;
										assign node906 = (inp[9]) ? node914 : node907;
											assign node907 = (inp[1]) ? node911 : node908;
												assign node908 = (inp[4]) ? 14'b01011100110000 : 14'b01001100110100;
												assign node911 = (inp[6]) ? 14'b01001000110000 : 14'b01001010110000;
											assign node914 = (inp[4]) ? node920 : node915;
												assign node915 = (inp[6]) ? 14'b01001000010100 : node916;
													assign node916 = (inp[1]) ? 14'b01001000000100 : 14'b01001100000100;
												assign node920 = (inp[6]) ? node922 : 14'b01001000000000;
													assign node922 = (inp[1]) ? 14'b01001000010000 : 14'b01001100010000;
									assign node925 = (inp[11]) ? 14'b00000000000001 : node926;
										assign node926 = (inp[4]) ? node932 : node927;
											assign node927 = (inp[7]) ? 14'b01001010110010 : node928;
												assign node928 = (inp[9]) ? 14'b01011100010010 : 14'b01011100110010;
											assign node932 = (inp[7]) ? node938 : node933;
												assign node933 = (inp[9]) ? node935 : 14'b00111000110000;
													assign node935 = (inp[1]) ? 14'b00111000010000 : 14'b00111100010000;
												assign node938 = (inp[6]) ? 14'b00101100010000 : 14'b00101110110000;
								assign node942 = (inp[7]) ? node962 : node943;
									assign node943 = (inp[6]) ? node959 : node944;
										assign node944 = (inp[11]) ? node956 : node945;
											assign node945 = (inp[4]) ? node951 : node946;
												assign node946 = (inp[1]) ? node948 : 14'b01011110110110;
													assign node948 = (inp[9]) ? 14'b01011010010010 : 14'b01011010110010;
												assign node951 = (inp[10]) ? node953 : 14'b00000000000001;
													assign node953 = (inp[1]) ? 14'b00111010110000 : 14'b00111110110000;
											assign node956 = (inp[10]) ? 14'b00000000000001 : 14'b01011010110000;
										assign node959 = (inp[1]) ? 14'b01011000100100 : 14'b00000000000001;
									assign node962 = (inp[1]) ? 14'b00000000000001 : node963;
										assign node963 = (inp[6]) ? node965 : 14'b00000000000001;
											assign node965 = (inp[9]) ? 14'b00000000000001 : node966;
												assign node966 = (inp[10]) ? 14'b01001100100010 : 14'b01001100100110;
							assign node971 = (inp[6]) ? node1015 : node972;
								assign node972 = (inp[7]) ? node996 : node973;
									assign node973 = (inp[3]) ? node983 : node974;
										assign node974 = (inp[1]) ? node980 : node975;
											assign node975 = (inp[9]) ? node977 : 14'b00000000000001;
												assign node977 = (inp[4]) ? 14'b00000100000100 : 14'b01000100000100;
											assign node980 = (inp[4]) ? 14'b00010110100100 : 14'b01010110000100;
										assign node983 = (inp[1]) ? node991 : node984;
											assign node984 = (inp[4]) ? node988 : node985;
												assign node985 = (inp[10]) ? 14'b01010110110100 : 14'b01010110010100;
												assign node988 = (inp[11]) ? 14'b00010110010100 : 14'b00010110110100;
											assign node991 = (inp[9]) ? node993 : 14'b01000110100100;
												assign node993 = (inp[4]) ? 14'b00000110000100 : 14'b01000110000100;
									assign node996 = (inp[1]) ? node1002 : node997;
										assign node997 = (inp[3]) ? node999 : 14'b00000000000001;
											assign node999 = (inp[4]) ? 14'b00010010110100 : 14'b01010010010100;
										assign node1002 = (inp[4]) ? node1008 : node1003;
											assign node1003 = (inp[3]) ? 14'b01000010100100 : node1004;
												assign node1004 = (inp[9]) ? 14'b01010010000100 : 14'b01010010100100;
											assign node1008 = (inp[9]) ? node1012 : node1009;
												assign node1009 = (inp[3]) ? 14'b00000010100100 : 14'b00010010100100;
												assign node1012 = (inp[3]) ? 14'b00000010000100 : 14'b00010010000100;
								assign node1015 = (inp[3]) ? 14'b00000000000001 : node1016;
									assign node1016 = (inp[9]) ? node1026 : node1017;
										assign node1017 = (inp[1]) ? node1021 : node1018;
											assign node1018 = (inp[10]) ? 14'b01010100110100 : 14'b00010100110100;
											assign node1021 = (inp[4]) ? node1023 : 14'b01010000100100;
												assign node1023 = (inp[7]) ? 14'b00010000100100 : 14'b00010100100100;
										assign node1026 = (inp[1]) ? 14'b01010100000100 : node1027;
											assign node1027 = (inp[4]) ? 14'b00010000010100 : 14'b01010000010100;
						assign node1032 = (inp[10]) ? 14'b00000000000001 : node1033;
							assign node1033 = (inp[13]) ? 14'b00000000000001 : node1034;
								assign node1034 = (inp[3]) ? node1064 : node1035;
									assign node1035 = (inp[6]) ? node1047 : node1036;
										assign node1036 = (inp[7]) ? node1040 : node1037;
											assign node1037 = (inp[9]) ? 14'b01000100000110 : 14'b00000000000001;
											assign node1040 = (inp[9]) ? node1042 : 14'b01000110110010;
												assign node1042 = (inp[11]) ? node1044 : 14'b01000010010010;
													assign node1044 = (inp[1]) ? 14'b01000010010000 : 14'b01000110010000;
										assign node1047 = (inp[9]) ? node1053 : node1048;
											assign node1048 = (inp[11]) ? 14'b01010000110000 : node1049;
												assign node1049 = (inp[7]) ? 14'b01000000110110 : 14'b01010000110110;
											assign node1053 = (inp[11]) ? node1059 : node1054;
												assign node1054 = (inp[7]) ? node1056 : 14'b01010100010110;
													assign node1056 = (inp[4]) ? 14'b01000100010010 : 14'b01000100010110;
												assign node1059 = (inp[7]) ? node1061 : 14'b01010100010100;
													assign node1061 = (inp[1]) ? 14'b01000000010100 : 14'b01000100010100;
									assign node1064 = (inp[7]) ? node1072 : node1065;
										assign node1065 = (inp[6]) ? 14'b00000000000001 : node1066;
											assign node1066 = (inp[1]) ? 14'b01010010010110 : node1067;
												assign node1067 = (inp[4]) ? 14'b01010110110000 : 14'b01010110110100;
										assign node1072 = (inp[6]) ? node1074 : 14'b00000000000001;
											assign node1074 = (inp[9]) ? 14'b00000000000001 : node1075;
												assign node1075 = (inp[4]) ? 14'b01000100100010 : node1076;
													assign node1076 = (inp[11]) ? 14'b01000000100100 : 14'b01000000100110;
				assign node1083 = (inp[4]) ? node1337 : node1084;
					assign node1084 = (inp[5]) ? node1244 : node1085;
						assign node1085 = (inp[13]) ? node1177 : node1086;
							assign node1086 = (inp[11]) ? node1150 : node1087;
								assign node1087 = (inp[3]) ? node1133 : node1088;
									assign node1088 = (inp[12]) ? node1112 : node1089;
										assign node1089 = (inp[10]) ? node1099 : node1090;
											assign node1090 = (inp[6]) ? node1096 : node1091;
												assign node1091 = (inp[1]) ? node1093 : 14'b00000000000001;
													assign node1093 = (inp[7]) ? 14'b00001010110000 : 14'b00011010000000;
												assign node1096 = (inp[7]) ? 14'b00001100010000 : 14'b00011100010000;
											assign node1099 = (inp[1]) ? node1107 : node1100;
												assign node1100 = (inp[7]) ? node1104 : node1101;
													assign node1101 = (inp[6]) ? 14'b00111100010010 : 14'b00101100000010;
													assign node1104 = (inp[9]) ? 14'b00101110010010 : 14'b00101110110010;
												assign node1107 = (inp[9]) ? node1109 : 14'b00111000110010;
													assign node1109 = (inp[7]) ? 14'b00101000010010 : 14'b00101000000010;
										assign node1112 = (inp[1]) ? node1122 : node1113;
											assign node1113 = (inp[7]) ? node1119 : node1114;
												assign node1114 = (inp[6]) ? node1116 : 14'b00001100000110;
													assign node1116 = (inp[10]) ? 14'b00011100010010 : 14'b00011100010110;
												assign node1119 = (inp[6]) ? 14'b00001100110110 : 14'b00001110010110;
											assign node1122 = (inp[6]) ? node1128 : node1123;
												assign node1123 = (inp[7]) ? node1125 : 14'b00011010000110;
													assign node1125 = (inp[9]) ? 14'b00001010010010 : 14'b00001010110110;
												assign node1128 = (inp[10]) ? 14'b00001000110010 : node1129;
													assign node1129 = (inp[7]) ? 14'b00001000110110 : 14'b00011000110110;
									assign node1133 = (inp[9]) ? node1145 : node1134;
										assign node1134 = (inp[1]) ? node1140 : node1135;
											assign node1135 = (inp[10]) ? node1137 : 14'b00000000000001;
												assign node1137 = (inp[12]) ? 14'b00000000000001 : 14'b00111110110010;
											assign node1140 = (inp[12]) ? node1142 : 14'b00101000100010;
												assign node1142 = (inp[6]) ? 14'b00011000100110 : 14'b00011010110110;
										assign node1145 = (inp[7]) ? 14'b00000000000001 : node1146;
											assign node1146 = (inp[12]) ? 14'b00011110010010 : 14'b00000000000001;
								assign node1150 = (inp[10]) ? 14'b00000000000001 : node1151;
									assign node1151 = (inp[3]) ? node1167 : node1152;
										assign node1152 = (inp[7]) ? node1158 : node1153;
											assign node1153 = (inp[6]) ? node1155 : 14'b00000000000001;
												assign node1155 = (inp[1]) ? 14'b00011000110100 : 14'b00011100110100;
											assign node1158 = (inp[12]) ? node1162 : node1159;
												assign node1159 = (inp[9]) ? 14'b00101000010100 : 14'b00101000110100;
												assign node1162 = (inp[6]) ? 14'b00001000010100 : node1163;
													assign node1163 = (inp[9]) ? 14'b00001010010100 : 14'b00001010110100;
										assign node1167 = (inp[7]) ? 14'b00000000000001 : node1168;
											assign node1168 = (inp[6]) ? 14'b00000000000001 : node1169;
												assign node1169 = (inp[1]) ? node1171 : 14'b00111110010100;
													assign node1171 = (inp[12]) ? 14'b00011010010100 : 14'b00111010010100;
							assign node1177 = (inp[12]) ? node1207 : node1178;
								assign node1178 = (inp[3]) ? node1198 : node1179;
									assign node1179 = (inp[6]) ? node1187 : node1180;
										assign node1180 = (inp[9]) ? node1182 : 14'b00000000000001;
											assign node1182 = (inp[1]) ? 14'b01110110000100 : node1183;
												assign node1183 = (inp[7]) ? 14'b01100000000100 : 14'b01100100000100;
										assign node1187 = (inp[1]) ? node1193 : node1188;
											assign node1188 = (inp[9]) ? node1190 : 14'b01110000110100;
												assign node1190 = (inp[7]) ? 14'b01110000010100 : 14'b01110100010100;
											assign node1193 = (inp[7]) ? node1195 : 14'b01110100100100;
												assign node1195 = (inp[10]) ? 14'b01110000100100 : 14'b01110000000100;
									assign node1198 = (inp[6]) ? 14'b00000000000001 : node1199;
										assign node1199 = (inp[1]) ? node1203 : node1200;
											assign node1200 = (inp[7]) ? 14'b01110010010100 : 14'b01110110010100;
											assign node1203 = (inp[7]) ? 14'b01100010000100 : 14'b01100110100100;
								assign node1207 = (inp[6]) ? node1231 : node1208;
									assign node1208 = (inp[3]) ? node1218 : node1209;
										assign node1209 = (inp[1]) ? node1213 : node1210;
											assign node1210 = (inp[9]) ? 14'b01000100000000 : 14'b00000000000001;
											assign node1213 = (inp[10]) ? node1215 : 14'b01010010000000;
												assign node1215 = (inp[7]) ? 14'b01010010100000 : 14'b01010110100000;
										assign node1218 = (inp[1]) ? node1226 : node1219;
											assign node1219 = (inp[9]) ? node1223 : node1220;
												assign node1220 = (inp[11]) ? 14'b01010110110000 : 14'b01010010110000;
												assign node1223 = (inp[7]) ? 14'b01010010010000 : 14'b01010110010000;
											assign node1226 = (inp[7]) ? node1228 : 14'b01000110000000;
												assign node1228 = (inp[10]) ? 14'b01000010100000 : 14'b01000010000000;
									assign node1231 = (inp[3]) ? 14'b00000000000001 : node1232;
										assign node1232 = (inp[9]) ? node1238 : node1233;
											assign node1233 = (inp[7]) ? node1235 : 14'b01010100100000;
												assign node1235 = (inp[10]) ? 14'b01010000100000 : 14'b01010000110000;
											assign node1238 = (inp[1]) ? 14'b01010000000000 : node1239;
												assign node1239 = (inp[7]) ? 14'b01010000010000 : 14'b01010100010000;
						assign node1244 = (inp[13]) ? node1326 : node1245;
							assign node1245 = (inp[10]) ? node1305 : node1246;
								assign node1246 = (inp[7]) ? node1284 : node1247;
									assign node1247 = (inp[6]) ? node1265 : node1248;
										assign node1248 = (inp[3]) ? node1260 : node1249;
											assign node1249 = (inp[1]) ? node1253 : node1250;
												assign node1250 = (inp[9]) ? 14'b00000100000100 : 14'b00000000000001;
												assign node1253 = (inp[9]) ? node1257 : node1254;
													assign node1254 = (inp[11]) ? 14'b00110010000100 : 14'b00010010000110;
													assign node1257 = (inp[12]) ? 14'b00000000000100 : 14'b00000000000000;
											assign node1260 = (inp[11]) ? 14'b00010010010100 : node1261;
												assign node1261 = (inp[1]) ? 14'b00010010010000 : 14'b00010110010000;
										assign node1265 = (inp[12]) ? node1273 : node1266;
											assign node1266 = (inp[9]) ? node1270 : node1267;
												assign node1267 = (inp[11]) ? 14'b00110000100100 : 14'b00010000100000;
												assign node1270 = (inp[11]) ? 14'b00000000000001 : 14'b00010000010000;
											assign node1273 = (inp[1]) ? node1277 : node1274;
												assign node1274 = (inp[9]) ? 14'b00010100010110 : 14'b00010100110110;
												assign node1277 = (inp[3]) ? node1281 : node1278;
													assign node1278 = (inp[11]) ? 14'b00010000110100 : 14'b00010000110110;
													assign node1281 = (inp[11]) ? 14'b00010000100100 : 14'b00010000100110;
									assign node1284 = (inp[3]) ? node1300 : node1285;
										assign node1285 = (inp[11]) ? node1293 : node1286;
											assign node1286 = (inp[9]) ? node1290 : node1287;
												assign node1287 = (inp[6]) ? 14'b00000000110000 : 14'b00000010110000;
												assign node1290 = (inp[6]) ? 14'b00000100010000 : 14'b00000110010000;
											assign node1293 = (inp[1]) ? node1297 : node1294;
												assign node1294 = (inp[6]) ? 14'b00100100010100 : 14'b00100110010100;
												assign node1297 = (inp[9]) ? 14'b00100000010100 : 14'b00100000110100;
										assign node1300 = (inp[9]) ? 14'b00000000000001 : node1301;
											assign node1301 = (inp[6]) ? 14'b00000100100000 : 14'b00000000000001;
								assign node1305 = (inp[11]) ? 14'b00000000000001 : node1306;
									assign node1306 = (inp[12]) ? node1308 : 14'b00000000000001;
										assign node1308 = (inp[6]) ? node1318 : node1309;
											assign node1309 = (inp[1]) ? node1315 : node1310;
												assign node1310 = (inp[9]) ? 14'b00010110010010 : node1311;
													assign node1311 = (inp[7]) ? 14'b00000110110010 : 14'b00010110110010;
												assign node1315 = (inp[7]) ? 14'b00000010010010 : 14'b00010010000010;
											assign node1318 = (inp[9]) ? 14'b00000000000001 : node1319;
												assign node1319 = (inp[1]) ? node1321 : 14'b00000100110010;
													assign node1321 = (inp[3]) ? 14'b00010000100010 : 14'b00010000110010;
							assign node1326 = (inp[9]) ? 14'b00000000000001 : node1327;
								assign node1327 = (inp[3]) ? 14'b00000000000001 : node1328;
									assign node1328 = (inp[6]) ? 14'b00000000000001 : node1329;
										assign node1329 = (inp[7]) ? node1331 : 14'b00000000000001;
											assign node1331 = (inp[12]) ? 14'b10001000001000 : 14'b00000000000001;
					assign node1337 = (inp[12]) ? 14'b00000000000001 : node1338;
						assign node1338 = (inp[11]) ? node1396 : node1339;
							assign node1339 = (inp[5]) ? node1351 : node1340;
								assign node1340 = (inp[13]) ? 14'b00000000000001 : node1341;
									assign node1341 = (inp[3]) ? 14'b00000000000001 : node1342;
										assign node1342 = (inp[10]) ? 14'b00000000000001 : node1343;
											assign node1343 = (inp[6]) ? node1345 : 14'b00000000000001;
												assign node1345 = (inp[1]) ? 14'b00101000110110 : 14'b00101100110110;
								assign node1351 = (inp[13]) ? node1381 : node1352;
									assign node1352 = (inp[1]) ? node1366 : node1353;
										assign node1353 = (inp[3]) ? node1359 : node1354;
											assign node1354 = (inp[10]) ? 14'b00000000000001 : node1355;
												assign node1355 = (inp[7]) ? 14'b00100100110110 : 14'b00110100110110;
											assign node1359 = (inp[9]) ? 14'b00000000000001 : node1360;
												assign node1360 = (inp[7]) ? node1362 : 14'b00000000000001;
													assign node1362 = (inp[6]) ? 14'b00100100100000 : 14'b00000000000001;
										assign node1366 = (inp[10]) ? node1374 : node1367;
											assign node1367 = (inp[6]) ? node1371 : node1368;
												assign node1368 = (inp[7]) ? 14'b00100010110110 : 14'b00110010110110;
												assign node1371 = (inp[9]) ? 14'b00100000010110 : 14'b00100000100110;
											assign node1374 = (inp[6]) ? 14'b00000000000001 : node1375;
												assign node1375 = (inp[3]) ? 14'b00110010110000 : node1376;
													assign node1376 = (inp[9]) ? 14'b00100010010000 : 14'b00110010000000;
									assign node1381 = (inp[7]) ? 14'b00000000000001 : node1382;
										assign node1382 = (inp[6]) ? node1392 : node1383;
											assign node1383 = (inp[10]) ? node1387 : node1384;
												assign node1384 = (inp[9]) ? 14'b00010110010000 : 14'b00010110110000;
												assign node1387 = (inp[3]) ? 14'b00000110000000 : node1388;
													assign node1388 = (inp[9]) ? 14'b00010110000000 : 14'b00010110100000;
											assign node1392 = (inp[3]) ? 14'b00000000000001 : 14'b00010100110000;
							assign node1396 = (inp[13]) ? node1398 : 14'b00000000000001;
								assign node1398 = (inp[9]) ? 14'b00000000000001 : node1399;
									assign node1399 = (inp[7]) ? node1405 : node1400;
										assign node1400 = (inp[3]) ? 14'b00010110110000 : node1401;
											assign node1401 = (inp[6]) ? 14'b00010100100000 : 14'b00000000000001;
										assign node1405 = (inp[6]) ? node1407 : 14'b00000000000001;
											assign node1407 = (inp[10]) ? 14'b00000000000001 : node1408;
												assign node1408 = (inp[3]) ? 14'b10000000000000 : 14'b00000000000001;
			assign node1414 = (inp[7]) ? node1726 : node1415;
				assign node1415 = (inp[1]) ? node1611 : node1416;
					assign node1416 = (inp[3]) ? node1544 : node1417;
						assign node1417 = (inp[2]) ? node1499 : node1418;
							assign node1418 = (inp[13]) ? node1468 : node1419;
								assign node1419 = (inp[6]) ? node1447 : node1420;
									assign node1420 = (inp[9]) ? node1430 : node1421;
										assign node1421 = (inp[5]) ? node1423 : 14'b01011110100010;
											assign node1423 = (inp[4]) ? node1425 : 14'b01010110100100;
												assign node1425 = (inp[12]) ? 14'b01010110100010 : node1426;
													assign node1426 = (inp[10]) ? 14'b01110110100000 : 14'b01110110100110;
										assign node1430 = (inp[10]) ? node1442 : node1431;
											assign node1431 = (inp[12]) ? node1439 : node1432;
												assign node1432 = (inp[4]) ? 14'b01111110000110 : node1433;
													assign node1433 = (inp[5]) ? node1435 : 14'b00000000000001;
														assign node1435 = (inp[11]) ? 14'b01110110000100 : 14'b00110110000010;
												assign node1439 = (inp[5]) ? 14'b01010110000010 : 14'b01011110000110;
											assign node1442 = (inp[12]) ? 14'b00000000000001 : node1443;
												assign node1443 = (inp[5]) ? 14'b01110110000000 : 14'b00000000000001;
									assign node1447 = (inp[11]) ? node1461 : node1448;
										assign node1448 = (inp[4]) ? node1456 : node1449;
											assign node1449 = (inp[12]) ? node1453 : node1450;
												assign node1450 = (inp[5]) ? 14'b00110100100010 : 14'b00000000000001;
												assign node1453 = (inp[5]) ? 14'b00000000000001 : 14'b01011100000110;
											assign node1456 = (inp[10]) ? node1458 : 14'b01110100100110;
												assign node1458 = (inp[12]) ? 14'b00111100000000 : 14'b01110100000000;
										assign node1461 = (inp[10]) ? 14'b00000000000001 : node1462;
											assign node1462 = (inp[9]) ? 14'b01110100000100 : node1463;
												assign node1463 = (inp[12]) ? 14'b01010100100000 : 14'b00000000000001;
								assign node1468 = (inp[4]) ? node1484 : node1469;
									assign node1469 = (inp[5]) ? node1477 : node1470;
										assign node1470 = (inp[12]) ? node1472 : 14'b00000000000001;
											assign node1472 = (inp[9]) ? 14'b01000110010100 : node1473;
												assign node1473 = (inp[11]) ? 14'b01000110110100 : 14'b01000100110100;
										assign node1477 = (inp[12]) ? 14'b00000000000001 : node1478;
											assign node1478 = (inp[9]) ? 14'b01100100010000 : node1479;
												assign node1479 = (inp[6]) ? 14'b01100100110000 : 14'b01100110110000;
									assign node1484 = (inp[5]) ? node1496 : node1485;
										assign node1485 = (inp[12]) ? node1491 : node1486;
											assign node1486 = (inp[6]) ? 14'b00100100010100 : node1487;
												assign node1487 = (inp[9]) ? 14'b00100110010100 : 14'b00100110110100;
											assign node1491 = (inp[6]) ? node1493 : 14'b00000110010100;
												assign node1493 = (inp[9]) ? 14'b00000100010100 : 14'b00000100110100;
										assign node1496 = (inp[9]) ? 14'b00100100010000 : 14'b00100100110000;
							assign node1499 = (inp[4]) ? node1529 : node1500;
								assign node1500 = (inp[5]) ? node1522 : node1501;
									assign node1501 = (inp[13]) ? node1511 : node1502;
										assign node1502 = (inp[10]) ? 14'b00000000000001 : node1503;
											assign node1503 = (inp[9]) ? node1507 : node1504;
												assign node1504 = (inp[11]) ? 14'b00111110100100 : 14'b00011110100000;
												assign node1507 = (inp[6]) ? 14'b00111100000100 : 14'b00011110000100;
										assign node1511 = (inp[12]) ? node1515 : node1512;
											assign node1512 = (inp[6]) ? 14'b01100100010100 : 14'b01100110010100;
											assign node1515 = (inp[6]) ? node1519 : node1516;
												assign node1516 = (inp[9]) ? 14'b01000110010000 : 14'b01000110110000;
												assign node1519 = (inp[9]) ? 14'b01000100010000 : 14'b01000100110000;
									assign node1522 = (inp[13]) ? 14'b00000000000001 : node1523;
										assign node1523 = (inp[10]) ? 14'b00000000000001 : node1524;
											assign node1524 = (inp[9]) ? 14'b00010100000000 : 14'b00010100100110;
								assign node1529 = (inp[12]) ? 14'b00000000000001 : node1530;
									assign node1530 = (inp[11]) ? node1538 : node1531;
										assign node1531 = (inp[13]) ? 14'b00000000000001 : node1532;
											assign node1532 = (inp[10]) ? 14'b00110110100000 : node1533;
												assign node1533 = (inp[5]) ? 14'b00110100000110 : 14'b00111100100110;
										assign node1538 = (inp[5]) ? node1540 : 14'b00000000000001;
											assign node1540 = (inp[9]) ? 14'b00000110010000 : 14'b00000000000001;
						assign node1544 = (inp[9]) ? 14'b00000000000001 : node1545;
							assign node1545 = (inp[13]) ? node1591 : node1546;
								assign node1546 = (inp[4]) ? node1572 : node1547;
									assign node1547 = (inp[10]) ? node1567 : node1548;
										assign node1548 = (inp[6]) ? node1558 : node1549;
											assign node1549 = (inp[12]) ? node1553 : node1550;
												assign node1550 = (inp[2]) ? 14'b00100110100100 : 14'b01100110100100;
												assign node1553 = (inp[5]) ? 14'b00000110100110 : node1554;
													assign node1554 = (inp[11]) ? 14'b00001110100100 : 14'b00001110100110;
											assign node1558 = (inp[2]) ? node1562 : node1559;
												assign node1559 = (inp[5]) ? 14'b01000110000100 : 14'b01001110000100;
												assign node1562 = (inp[11]) ? node1564 : 14'b00001110000000;
													assign node1564 = (inp[12]) ? 14'b00001110000100 : 14'b00101110000100;
										assign node1567 = (inp[11]) ? 14'b00000000000001 : node1568;
											assign node1568 = (inp[5]) ? 14'b01100110000010 : 14'b01101110000010;
									assign node1572 = (inp[2]) ? node1584 : node1573;
										assign node1573 = (inp[11]) ? 14'b00000000000001 : node1574;
											assign node1574 = (inp[12]) ? node1580 : node1575;
												assign node1575 = (inp[10]) ? 14'b01100110000000 : node1576;
													assign node1576 = (inp[5]) ? 14'b01100110000110 : 14'b01101110000110;
												assign node1580 = (inp[5]) ? 14'b01000110100010 : 14'b00000000000001;
										assign node1584 = (inp[11]) ? 14'b00000000000001 : node1585;
											assign node1585 = (inp[12]) ? 14'b00000000000001 : node1586;
												assign node1586 = (inp[10]) ? 14'b00000000000001 : 14'b00101110000110;
								assign node1591 = (inp[6]) ? node1599 : node1592;
									assign node1592 = (inp[2]) ? node1594 : 14'b00000000000001;
										assign node1594 = (inp[11]) ? 14'b00000000000001 : node1595;
											assign node1595 = (inp[10]) ? 14'b10000001000000 : 14'b00000000000001;
									assign node1599 = (inp[12]) ? 14'b00000000000001 : node1600;
										assign node1600 = (inp[4]) ? node1606 : node1601;
											assign node1601 = (inp[2]) ? 14'b00000000000001 : node1602;
												assign node1602 = (inp[5]) ? 14'b01100100100000 : 14'b00000000000001;
											assign node1606 = (inp[5]) ? 14'b00100100100000 : 14'b00100100100100;
					assign node1611 = (inp[13]) ? node1705 : node1612;
						assign node1612 = (inp[6]) ? node1684 : node1613;
							assign node1613 = (inp[9]) ? node1667 : node1614;
								assign node1614 = (inp[11]) ? node1652 : node1615;
									assign node1615 = (inp[4]) ? node1639 : node1616;
										assign node1616 = (inp[12]) ? node1628 : node1617;
											assign node1617 = (inp[5]) ? node1623 : node1618;
												assign node1618 = (inp[2]) ? node1620 : 14'b00000000000001;
													assign node1620 = (inp[10]) ? 14'b00101010100010 : 14'b00001010100000;
												assign node1623 = (inp[2]) ? 14'b00000010100000 : node1624;
													assign node1624 = (inp[3]) ? 14'b00100010100010 : 14'b00110010100010;
											assign node1628 = (inp[10]) ? node1636 : node1629;
												assign node1629 = (inp[2]) ? node1631 : 14'b01010010100110;
													assign node1631 = (inp[5]) ? 14'b00000010100110 : node1632;
														assign node1632 = (inp[3]) ? 14'b00001010100110 : 14'b00011010100110;
												assign node1636 = (inp[2]) ? 14'b00011010100010 : 14'b01001010100010;
										assign node1639 = (inp[12]) ? node1645 : node1640;
											assign node1640 = (inp[2]) ? 14'b00111010100110 : node1641;
												assign node1641 = (inp[3]) ? 14'b01101010100000 : 14'b01110010100000;
											assign node1645 = (inp[2]) ? 14'b00000000000001 : node1646;
												assign node1646 = (inp[3]) ? 14'b00000000000001 : node1647;
													assign node1647 = (inp[10]) ? 14'b00111010100000 : 14'b01010010100010;
									assign node1652 = (inp[10]) ? 14'b00000000000001 : node1653;
										assign node1653 = (inp[3]) ? node1663 : node1654;
											assign node1654 = (inp[12]) ? node1658 : node1655;
												assign node1655 = (inp[5]) ? 14'b01110010100100 : 14'b01111010100100;
												assign node1658 = (inp[4]) ? node1660 : 14'b01011010100100;
													assign node1660 = (inp[5]) ? 14'b01010010100000 : 14'b01011010100000;
											assign node1663 = (inp[12]) ? 14'b00000010100100 : 14'b00000000000001;
								assign node1667 = (inp[3]) ? node1669 : 14'b00000000000001;
									assign node1669 = (inp[5]) ? node1677 : node1670;
										assign node1670 = (inp[4]) ? node1674 : node1671;
											assign node1671 = (inp[11]) ? 14'b01101010000100 : 14'b00101010000010;
											assign node1674 = (inp[10]) ? 14'b00101010000000 : 14'b00000000000001;
										assign node1677 = (inp[10]) ? 14'b00000000000001 : node1678;
											assign node1678 = (inp[12]) ? node1680 : 14'b00000000000001;
												assign node1680 = (inp[11]) ? 14'b01000010000100 : 14'b01000010000010;
							assign node1684 = (inp[3]) ? 14'b00000000000001 : node1685;
								assign node1685 = (inp[9]) ? node1687 : 14'b00000000000001;
									assign node1687 = (inp[10]) ? node1695 : node1688;
										assign node1688 = (inp[12]) ? node1692 : node1689;
											assign node1689 = (inp[11]) ? 14'b00111000000100 : 14'b01111000000110;
											assign node1692 = (inp[4]) ? 14'b00000000000001 : 14'b00011000000100;
										assign node1695 = (inp[11]) ? 14'b00000000000001 : node1696;
											assign node1696 = (inp[12]) ? node1698 : 14'b01111000000010;
												assign node1698 = (inp[4]) ? 14'b00000000000001 : node1699;
													assign node1699 = (inp[2]) ? 14'b00010000000010 : 14'b00000000000001;
						assign node1705 = (inp[3]) ? 14'b00000000000001 : node1706;
							assign node1706 = (inp[6]) ? 14'b00000000000001 : node1707;
								assign node1707 = (inp[9]) ? 14'b00000000000001 : node1708;
									assign node1708 = (inp[4]) ? node1718 : node1709;
										assign node1709 = (inp[5]) ? node1711 : 14'b00000000000001;
											assign node1711 = (inp[10]) ? node1713 : 14'b10000000001010;
												assign node1713 = (inp[12]) ? node1715 : 14'b00000000000001;
													assign node1715 = (inp[2]) ? 14'b00000000000001 : 14'b10001001001000;
										assign node1718 = (inp[5]) ? 14'b00000000000001 : node1719;
											assign node1719 = (inp[12]) ? 14'b00000000000001 : 14'b10000001000010;
				assign node1726 = (inp[13]) ? node1728 : 14'b00000000000001;
					assign node1728 = (inp[1]) ? node1788 : node1729;
						assign node1729 = (inp[3]) ? node1771 : node1730;
							assign node1730 = (inp[5]) ? node1762 : node1731;
								assign node1731 = (inp[4]) ? node1753 : node1732;
									assign node1732 = (inp[6]) ? node1744 : node1733;
										assign node1733 = (inp[9]) ? node1739 : node1734;
											assign node1734 = (inp[10]) ? node1736 : 14'b00000010110000;
												assign node1736 = (inp[12]) ? 14'b01000010110100 : 14'b01100010110100;
											assign node1739 = (inp[12]) ? node1741 : 14'b01100010010100;
												assign node1741 = (inp[2]) ? 14'b01000010010000 : 14'b01000010010100;
										assign node1744 = (inp[9]) ? node1748 : node1745;
											assign node1745 = (inp[2]) ? 14'b01000000110000 : 14'b01000000110100;
											assign node1748 = (inp[12]) ? node1750 : 14'b00000000010000;
												assign node1750 = (inp[2]) ? 14'b01000000010000 : 14'b01000000010100;
									assign node1753 = (inp[2]) ? 14'b00000000000001 : node1754;
										assign node1754 = (inp[9]) ? node1758 : node1755;
											assign node1755 = (inp[6]) ? 14'b00000000110100 : 14'b00000010110100;
											assign node1758 = (inp[6]) ? 14'b00100000010100 : 14'b00000010010100;
								assign node1762 = (inp[12]) ? 14'b00000000000001 : node1763;
									assign node1763 = (inp[2]) ? 14'b00000000000001 : node1764;
										assign node1764 = (inp[9]) ? 14'b01100010010000 : node1765;
											assign node1765 = (inp[4]) ? 14'b00100010110000 : 14'b01100010110000;
							assign node1771 = (inp[6]) ? node1773 : 14'b00000000000001;
								assign node1773 = (inp[5]) ? 14'b00000000000001 : node1774;
									assign node1774 = (inp[9]) ? 14'b00000000000001 : node1775;
										assign node1775 = (inp[2]) ? node1781 : node1776;
											assign node1776 = (inp[4]) ? node1778 : 14'b00000000100000;
												assign node1778 = (inp[12]) ? 14'b00000000100100 : 14'b00100000100100;
											assign node1781 = (inp[4]) ? 14'b00000000000001 : node1782;
												assign node1782 = (inp[10]) ? 14'b01100000100100 : 14'b01000000100000;
						assign node1788 = (inp[12]) ? node1790 : 14'b00000000000001;
							assign node1790 = (inp[3]) ? node1792 : 14'b00000000000001;
								assign node1792 = (inp[5]) ? node1794 : 14'b00000000000001;
									assign node1794 = (inp[2]) ? node1796 : 14'b00000000000001;
										assign node1796 = (inp[9]) ? node1798 : 14'b00000000000001;
											assign node1798 = (inp[6]) ? 14'b10001001000000 : 14'b10001000000000;

endmodule