module dtc_split66_bm40 (
	input  wire [16-1:0] inp,
	output wire [40-1:0] outp
);

	wire [40-1:0] node1;
	wire [40-1:0] node2;
	wire [40-1:0] node5;
	wire [40-1:0] node6;
	wire [40-1:0] node8;
	wire [40-1:0] node9;
	wire [40-1:0] node11;
	wire [40-1:0] node12;
	wire [40-1:0] node17;
	wire [40-1:0] node18;
	wire [40-1:0] node19;
	wire [40-1:0] node20;
	wire [40-1:0] node21;
	wire [40-1:0] node24;
	wire [40-1:0] node27;
	wire [40-1:0] node28;
	wire [40-1:0] node31;
	wire [40-1:0] node33;
	wire [40-1:0] node34;
	wire [40-1:0] node36;
	wire [40-1:0] node39;
	wire [40-1:0] node40;
	wire [40-1:0] node43;
	wire [40-1:0] node46;
	wire [40-1:0] node47;
	wire [40-1:0] node49;
	wire [40-1:0] node50;
	wire [40-1:0] node51;
	wire [40-1:0] node53;
	wire [40-1:0] node55;
	wire [40-1:0] node57;
	wire [40-1:0] node58;
	wire [40-1:0] node61;
	wire [40-1:0] node64;
	wire [40-1:0] node65;
	wire [40-1:0] node67;
	wire [40-1:0] node69;
	wire [40-1:0] node71;
	wire [40-1:0] node74;
	wire [40-1:0] node75;
	wire [40-1:0] node77;
	wire [40-1:0] node79;
	wire [40-1:0] node83;
	wire [40-1:0] node85;
	wire [40-1:0] node87;
	wire [40-1:0] node89;
	wire [40-1:0] node90;
	wire [40-1:0] node92;
	wire [40-1:0] node95;
	wire [40-1:0] node96;
	wire [40-1:0] node99;
	wire [40-1:0] node102;
	wire [40-1:0] node103;
	wire [40-1:0] node106;
	wire [40-1:0] node107;
	wire [40-1:0] node109;
	wire [40-1:0] node111;
	wire [40-1:0] node113;
	wire [40-1:0] node115;
	wire [40-1:0] node117;
	wire [40-1:0] node120;
	wire [40-1:0] node121;
	wire [40-1:0] node123;
	wire [40-1:0] node125;
	wire [40-1:0] node126;
	wire [40-1:0] node128;
	wire [40-1:0] node131;
	wire [40-1:0] node132;
	wire [40-1:0] node135;
	wire [40-1:0] node138;
	wire [40-1:0] node139;
	wire [40-1:0] node141;
	wire [40-1:0] node143;
	wire [40-1:0] node145;
	wire [40-1:0] node148;
	wire [40-1:0] node151;
	wire [40-1:0] node152;
	wire [40-1:0] node154;
	wire [40-1:0] node156;
	wire [40-1:0] node157;
	wire [40-1:0] node158;
	wire [40-1:0] node160;
	wire [40-1:0] node162;
	wire [40-1:0] node163;
	wire [40-1:0] node164;
	wire [40-1:0] node168;
	wire [40-1:0] node169;
	wire [40-1:0] node172;
	wire [40-1:0] node175;
	wire [40-1:0] node176;
	wire [40-1:0] node178;
	wire [40-1:0] node180;
	wire [40-1:0] node182;
	wire [40-1:0] node185;
	wire [40-1:0] node186;
	wire [40-1:0] node188;
	wire [40-1:0] node190;
	wire [40-1:0] node195;
	wire [40-1:0] node196;
	wire [40-1:0] node198;
	wire [40-1:0] node200;
	wire [40-1:0] node201;
	wire [40-1:0] node203;
	wire [40-1:0] node206;
	wire [40-1:0] node207;
	wire [40-1:0] node210;
	wire [40-1:0] node213;
	wire [40-1:0] node214;
	wire [40-1:0] node217;
	wire [40-1:0] node218;
	wire [40-1:0] node220;
	wire [40-1:0] node222;
	wire [40-1:0] node224;
	wire [40-1:0] node226;
	wire [40-1:0] node228;
	wire [40-1:0] node231;
	wire [40-1:0] node232;
	wire [40-1:0] node234;
	wire [40-1:0] node236;
	wire [40-1:0] node237;
	wire [40-1:0] node238;
	wire [40-1:0] node242;
	wire [40-1:0] node243;
	wire [40-1:0] node246;
	wire [40-1:0] node249;
	wire [40-1:0] node250;
	wire [40-1:0] node252;
	wire [40-1:0] node254;
	wire [40-1:0] node255;
	wire [40-1:0] node258;
	wire [40-1:0] node261;
	wire [40-1:0] node264;
	wire [40-1:0] node265;
	wire [40-1:0] node266;
	wire [40-1:0] node269;
	wire [40-1:0] node270;
	wire [40-1:0] node271;
	wire [40-1:0] node272;
	wire [40-1:0] node273;
	wire [40-1:0] node276;
	wire [40-1:0] node279;
	wire [40-1:0] node280;
	wire [40-1:0] node283;
	wire [40-1:0] node286;
	wire [40-1:0] node287;
	wire [40-1:0] node288;
	wire [40-1:0] node291;
	wire [40-1:0] node294;
	wire [40-1:0] node295;
	wire [40-1:0] node298;
	wire [40-1:0] node301;
	wire [40-1:0] node302;
	wire [40-1:0] node303;
	wire [40-1:0] node304;
	wire [40-1:0] node307;
	wire [40-1:0] node310;
	wire [40-1:0] node311;
	wire [40-1:0] node314;
	wire [40-1:0] node317;
	wire [40-1:0] node318;
	wire [40-1:0] node319;
	wire [40-1:0] node322;
	wire [40-1:0] node325;
	wire [40-1:0] node326;
	wire [40-1:0] node329;
	wire [40-1:0] node332;
	wire [40-1:0] node333;
	wire [40-1:0] node336;
	wire [40-1:0] node338;
	wire [40-1:0] node339;
	wire [40-1:0] node340;
	wire [40-1:0] node341;
	wire [40-1:0] node342;
	wire [40-1:0] node343;
	wire [40-1:0] node344;
	wire [40-1:0] node345;
	wire [40-1:0] node346;
	wire [40-1:0] node347;
	wire [40-1:0] node350;
	wire [40-1:0] node353;
	wire [40-1:0] node354;
	wire [40-1:0] node357;
	wire [40-1:0] node360;
	wire [40-1:0] node361;
	wire [40-1:0] node362;
	wire [40-1:0] node365;
	wire [40-1:0] node368;
	wire [40-1:0] node369;
	wire [40-1:0] node372;
	wire [40-1:0] node375;
	wire [40-1:0] node376;
	wire [40-1:0] node377;
	wire [40-1:0] node378;
	wire [40-1:0] node381;
	wire [40-1:0] node384;
	wire [40-1:0] node385;
	wire [40-1:0] node388;
	wire [40-1:0] node391;
	wire [40-1:0] node392;
	wire [40-1:0] node393;
	wire [40-1:0] node396;
	wire [40-1:0] node399;
	wire [40-1:0] node400;
	wire [40-1:0] node403;
	wire [40-1:0] node406;
	wire [40-1:0] node407;
	wire [40-1:0] node408;
	wire [40-1:0] node409;
	wire [40-1:0] node410;
	wire [40-1:0] node413;
	wire [40-1:0] node416;
	wire [40-1:0] node417;
	wire [40-1:0] node420;
	wire [40-1:0] node423;
	wire [40-1:0] node424;
	wire [40-1:0] node425;
	wire [40-1:0] node428;
	wire [40-1:0] node431;
	wire [40-1:0] node432;
	wire [40-1:0] node435;
	wire [40-1:0] node438;
	wire [40-1:0] node439;
	wire [40-1:0] node440;
	wire [40-1:0] node441;
	wire [40-1:0] node444;
	wire [40-1:0] node447;
	wire [40-1:0] node448;
	wire [40-1:0] node451;
	wire [40-1:0] node454;
	wire [40-1:0] node455;
	wire [40-1:0] node456;
	wire [40-1:0] node459;
	wire [40-1:0] node462;
	wire [40-1:0] node463;
	wire [40-1:0] node466;
	wire [40-1:0] node469;
	wire [40-1:0] node470;
	wire [40-1:0] node471;
	wire [40-1:0] node472;
	wire [40-1:0] node473;
	wire [40-1:0] node474;
	wire [40-1:0] node477;
	wire [40-1:0] node480;
	wire [40-1:0] node481;
	wire [40-1:0] node484;
	wire [40-1:0] node487;
	wire [40-1:0] node488;
	wire [40-1:0] node489;
	wire [40-1:0] node492;
	wire [40-1:0] node495;
	wire [40-1:0] node496;
	wire [40-1:0] node499;
	wire [40-1:0] node502;
	wire [40-1:0] node503;
	wire [40-1:0] node504;
	wire [40-1:0] node505;
	wire [40-1:0] node508;
	wire [40-1:0] node511;
	wire [40-1:0] node512;
	wire [40-1:0] node515;
	wire [40-1:0] node518;
	wire [40-1:0] node519;
	wire [40-1:0] node520;
	wire [40-1:0] node523;
	wire [40-1:0] node526;
	wire [40-1:0] node527;
	wire [40-1:0] node530;
	wire [40-1:0] node533;
	wire [40-1:0] node534;
	wire [40-1:0] node535;
	wire [40-1:0] node536;
	wire [40-1:0] node537;
	wire [40-1:0] node540;
	wire [40-1:0] node543;
	wire [40-1:0] node544;
	wire [40-1:0] node547;
	wire [40-1:0] node550;
	wire [40-1:0] node551;
	wire [40-1:0] node552;
	wire [40-1:0] node555;
	wire [40-1:0] node558;
	wire [40-1:0] node559;
	wire [40-1:0] node562;
	wire [40-1:0] node565;
	wire [40-1:0] node566;
	wire [40-1:0] node567;
	wire [40-1:0] node568;
	wire [40-1:0] node571;
	wire [40-1:0] node574;
	wire [40-1:0] node575;
	wire [40-1:0] node578;
	wire [40-1:0] node581;
	wire [40-1:0] node582;
	wire [40-1:0] node583;
	wire [40-1:0] node586;
	wire [40-1:0] node589;
	wire [40-1:0] node590;
	wire [40-1:0] node593;
	wire [40-1:0] node596;
	wire [40-1:0] node597;
	wire [40-1:0] node598;
	wire [40-1:0] node599;
	wire [40-1:0] node601;
	wire [40-1:0] node602;
	wire [40-1:0] node603;
	wire [40-1:0] node606;
	wire [40-1:0] node612;
	wire [40-1:0] node613;
	wire [40-1:0] node614;
	wire [40-1:0] node615;
	wire [40-1:0] node616;
	wire [40-1:0] node617;
	wire [40-1:0] node620;
	wire [40-1:0] node623;
	wire [40-1:0] node624;
	wire [40-1:0] node627;
	wire [40-1:0] node630;
	wire [40-1:0] node631;
	wire [40-1:0] node632;
	wire [40-1:0] node635;
	wire [40-1:0] node638;
	wire [40-1:0] node639;
	wire [40-1:0] node642;
	wire [40-1:0] node645;
	wire [40-1:0] node646;
	wire [40-1:0] node647;
	wire [40-1:0] node648;
	wire [40-1:0] node651;
	wire [40-1:0] node654;
	wire [40-1:0] node655;
	wire [40-1:0] node658;
	wire [40-1:0] node661;
	wire [40-1:0] node662;
	wire [40-1:0] node663;
	wire [40-1:0] node666;
	wire [40-1:0] node669;
	wire [40-1:0] node670;
	wire [40-1:0] node673;
	wire [40-1:0] node676;
	wire [40-1:0] node677;
	wire [40-1:0] node678;
	wire [40-1:0] node679;
	wire [40-1:0] node680;
	wire [40-1:0] node683;
	wire [40-1:0] node686;
	wire [40-1:0] node687;
	wire [40-1:0] node690;
	wire [40-1:0] node693;
	wire [40-1:0] node694;
	wire [40-1:0] node695;
	wire [40-1:0] node698;
	wire [40-1:0] node701;
	wire [40-1:0] node702;
	wire [40-1:0] node705;
	wire [40-1:0] node708;
	wire [40-1:0] node709;
	wire [40-1:0] node710;
	wire [40-1:0] node711;
	wire [40-1:0] node714;
	wire [40-1:0] node717;
	wire [40-1:0] node718;
	wire [40-1:0] node721;
	wire [40-1:0] node724;
	wire [40-1:0] node725;
	wire [40-1:0] node726;
	wire [40-1:0] node729;
	wire [40-1:0] node732;
	wire [40-1:0] node733;
	wire [40-1:0] node736;
	wire [40-1:0] node739;
	wire [40-1:0] node740;
	wire [40-1:0] node741;
	wire [40-1:0] node742;
	wire [40-1:0] node743;
	wire [40-1:0] node745;
	wire [40-1:0] node746;
	wire [40-1:0] node747;
	wire [40-1:0] node751;
	wire [40-1:0] node752;
	wire [40-1:0] node755;
	wire [40-1:0] node758;
	wire [40-1:0] node759;
	wire [40-1:0] node760;
	wire [40-1:0] node761;
	wire [40-1:0] node764;
	wire [40-1:0] node769;
	wire [40-1:0] node770;
	wire [40-1:0] node771;
	wire [40-1:0] node773;
	wire [40-1:0] node774;
	wire [40-1:0] node778;
	wire [40-1:0] node779;
	wire [40-1:0] node781;
	wire [40-1:0] node787;
	wire [40-1:0] node788;
	wire [40-1:0] node789;
	wire [40-1:0] node791;
	wire [40-1:0] node793;
	wire [40-1:0] node795;
	wire [40-1:0] node796;
	wire [40-1:0] node799;
	wire [40-1:0] node803;
	wire [40-1:0] node804;
	wire [40-1:0] node805;
	wire [40-1:0] node806;
	wire [40-1:0] node807;
	wire [40-1:0] node808;
	wire [40-1:0] node811;
	wire [40-1:0] node814;
	wire [40-1:0] node815;
	wire [40-1:0] node818;
	wire [40-1:0] node821;
	wire [40-1:0] node822;
	wire [40-1:0] node823;
	wire [40-1:0] node826;
	wire [40-1:0] node829;
	wire [40-1:0] node830;
	wire [40-1:0] node833;
	wire [40-1:0] node836;
	wire [40-1:0] node837;
	wire [40-1:0] node838;
	wire [40-1:0] node839;
	wire [40-1:0] node842;
	wire [40-1:0] node845;
	wire [40-1:0] node846;
	wire [40-1:0] node849;
	wire [40-1:0] node852;
	wire [40-1:0] node853;
	wire [40-1:0] node854;
	wire [40-1:0] node857;
	wire [40-1:0] node860;
	wire [40-1:0] node861;
	wire [40-1:0] node864;
	wire [40-1:0] node867;
	wire [40-1:0] node868;
	wire [40-1:0] node869;
	wire [40-1:0] node870;
	wire [40-1:0] node871;
	wire [40-1:0] node874;
	wire [40-1:0] node877;
	wire [40-1:0] node878;
	wire [40-1:0] node881;
	wire [40-1:0] node884;
	wire [40-1:0] node885;
	wire [40-1:0] node886;
	wire [40-1:0] node889;
	wire [40-1:0] node892;
	wire [40-1:0] node893;
	wire [40-1:0] node896;
	wire [40-1:0] node899;
	wire [40-1:0] node900;
	wire [40-1:0] node901;
	wire [40-1:0] node902;
	wire [40-1:0] node905;
	wire [40-1:0] node908;
	wire [40-1:0] node909;
	wire [40-1:0] node912;
	wire [40-1:0] node915;
	wire [40-1:0] node916;
	wire [40-1:0] node917;
	wire [40-1:0] node920;
	wire [40-1:0] node923;
	wire [40-1:0] node924;
	wire [40-1:0] node927;
	wire [40-1:0] node930;
	wire [40-1:0] node931;
	wire [40-1:0] node932;
	wire [40-1:0] node934;
	wire [40-1:0] node935;
	wire [40-1:0] node936;
	wire [40-1:0] node938;
	wire [40-1:0] node941;
	wire [40-1:0] node942;
	wire [40-1:0] node946;
	wire [40-1:0] node947;
	wire [40-1:0] node949;
	wire [40-1:0] node952;
	wire [40-1:0] node953;
	wire [40-1:0] node957;
	wire [40-1:0] node958;
	wire [40-1:0] node959;
	wire [40-1:0] node961;
	wire [40-1:0] node963;
	wire [40-1:0] node965;
	wire [40-1:0] node966;
	wire [40-1:0] node969;
	wire [40-1:0] node972;
	wire [40-1:0] node973;
	wire [40-1:0] node975;
	wire [40-1:0] node977;
	wire [40-1:0] node978;
	wire [40-1:0] node981;
	wire [40-1:0] node984;
	wire [40-1:0] node985;
	wire [40-1:0] node987;
	wire [40-1:0] node988;
	wire [40-1:0] node991;
	wire [40-1:0] node994;
	wire [40-1:0] node995;
	wire [40-1:0] node996;
	wire [40-1:0] node999;
	wire [40-1:0] node1004;
	wire [40-1:0] node1005;
	wire [40-1:0] node1006;
	wire [40-1:0] node1008;
	wire [40-1:0] node1009;
	wire [40-1:0] node1010;
	wire [40-1:0] node1011;
	wire [40-1:0] node1012;
	wire [40-1:0] node1015;
	wire [40-1:0] node1018;
	wire [40-1:0] node1019;
	wire [40-1:0] node1022;
	wire [40-1:0] node1025;
	wire [40-1:0] node1026;
	wire [40-1:0] node1027;
	wire [40-1:0] node1030;
	wire [40-1:0] node1033;
	wire [40-1:0] node1034;
	wire [40-1:0] node1037;
	wire [40-1:0] node1040;
	wire [40-1:0] node1041;
	wire [40-1:0] node1042;
	wire [40-1:0] node1043;
	wire [40-1:0] node1046;
	wire [40-1:0] node1049;
	wire [40-1:0] node1050;
	wire [40-1:0] node1053;
	wire [40-1:0] node1056;
	wire [40-1:0] node1057;
	wire [40-1:0] node1058;
	wire [40-1:0] node1061;
	wire [40-1:0] node1064;
	wire [40-1:0] node1065;
	wire [40-1:0] node1068;
	wire [40-1:0] node1071;
	wire [40-1:0] node1072;
	wire [40-1:0] node1073;
	wire [40-1:0] node1074;
	wire [40-1:0] node1075;
	wire [40-1:0] node1076;
	wire [40-1:0] node1079;
	wire [40-1:0] node1082;
	wire [40-1:0] node1083;
	wire [40-1:0] node1086;
	wire [40-1:0] node1089;
	wire [40-1:0] node1090;
	wire [40-1:0] node1091;
	wire [40-1:0] node1094;
	wire [40-1:0] node1097;
	wire [40-1:0] node1098;
	wire [40-1:0] node1101;
	wire [40-1:0] node1104;
	wire [40-1:0] node1105;
	wire [40-1:0] node1106;
	wire [40-1:0] node1107;
	wire [40-1:0] node1110;
	wire [40-1:0] node1113;
	wire [40-1:0] node1114;
	wire [40-1:0] node1117;
	wire [40-1:0] node1120;
	wire [40-1:0] node1121;
	wire [40-1:0] node1122;
	wire [40-1:0] node1125;
	wire [40-1:0] node1128;
	wire [40-1:0] node1129;
	wire [40-1:0] node1132;
	wire [40-1:0] node1136;
	wire [40-1:0] node1137;
	wire [40-1:0] node1138;
	wire [40-1:0] node1140;
	wire [40-1:0] node1141;
	wire [40-1:0] node1142;
	wire [40-1:0] node1143;
	wire [40-1:0] node1146;
	wire [40-1:0] node1149;
	wire [40-1:0] node1150;
	wire [40-1:0] node1153;
	wire [40-1:0] node1156;
	wire [40-1:0] node1157;
	wire [40-1:0] node1158;
	wire [40-1:0] node1161;
	wire [40-1:0] node1164;
	wire [40-1:0] node1165;
	wire [40-1:0] node1168;
	wire [40-1:0] node1171;
	wire [40-1:0] node1172;
	wire [40-1:0] node1173;
	wire [40-1:0] node1174;
	wire [40-1:0] node1175;
	wire [40-1:0] node1178;
	wire [40-1:0] node1181;
	wire [40-1:0] node1182;
	wire [40-1:0] node1185;
	wire [40-1:0] node1188;
	wire [40-1:0] node1189;
	wire [40-1:0] node1190;
	wire [40-1:0] node1193;
	wire [40-1:0] node1196;
	wire [40-1:0] node1197;
	wire [40-1:0] node1200;
	wire [40-1:0] node1204;
	wire [40-1:0] node1205;
	wire [40-1:0] node1206;
	wire [40-1:0] node1208;
	wire [40-1:0] node1209;
	wire [40-1:0] node1210;
	wire [40-1:0] node1213;
	wire [40-1:0] node1216;
	wire [40-1:0] node1217;
	wire [40-1:0] node1220;
	wire [40-1:0] node1223;
	wire [40-1:0] node1224;
	wire [40-1:0] node1225;
	wire [40-1:0] node1226;
	wire [40-1:0] node1229;
	wire [40-1:0] node1232;
	wire [40-1:0] node1233;
	wire [40-1:0] node1236;
	wire [40-1:0] node1240;
	wire [40-1:0] node1241;
	wire [40-1:0] node1243;
	wire [40-1:0] node1244;
	wire [40-1:0] node1245;
	wire [40-1:0] node1248;
	wire [40-1:0] node1251;
	wire [40-1:0] node1252;
	wire [40-1:0] node1255;
	wire [40-1:0] node1258;
	wire [40-1:0] node1259;
	wire [40-1:0] node1260;
	wire [40-1:0] node1261;
	wire [40-1:0] node1264;
	wire [40-1:0] node1267;
	wire [40-1:0] node1268;
	wire [40-1:0] node1271;

	assign outp = (inp[9]) ? node264 : node1;
		assign node1 = (inp[4]) ? node5 : node2;
			assign node2 = (inp[1]) ? 40'b0000000001000000000000000000000000000000 : 40'b0000000000000000000000000000000000000000;
			assign node5 = (inp[1]) ? node17 : node6;
				assign node6 = (inp[7]) ? node8 : 40'b0000000000000000000000000000000000000000;
					assign node8 = (inp[11]) ? 40'b0000000000000000000000000000000000000000 : node9;
						assign node9 = (inp[8]) ? node11 : 40'b0000000000000000000000000000000000000000;
							assign node11 = (inp[3]) ? 40'b0000000000000000000000000000000000000000 : node12;
								assign node12 = (inp[14]) ? 40'b0000000000000000000000000000000000000000 : 40'b0000000000000000100000000000000000000000;
				assign node17 = (inp[7]) ? node151 : node18;
					assign node18 = (inp[8]) ? node46 : node19;
						assign node19 = (inp[14]) ? node27 : node20;
							assign node20 = (inp[3]) ? node24 : node21;
								assign node21 = (inp[11]) ? 40'b0000000000000010000001000000000000000000 : 40'b0000000000000010000000000100000000000000;
								assign node24 = (inp[11]) ? 40'b0000000000000001010000000100000000000000 : 40'b0000000000100010000000000000000000000000;
							assign node27 = (inp[11]) ? node31 : node28;
								assign node28 = (inp[3]) ? 40'b0000000000100000000000000000000010000000 : 40'b0000000000000000000000000100000010000000;
								assign node31 = (inp[3]) ? node33 : 40'b0000000000000000000001000000000010000000;
									assign node33 = (inp[13]) ? node39 : node34;
										assign node34 = (inp[0]) ? node36 : 40'b0000000000000000000000000000000000000000;
											assign node36 = (inp[10]) ? 40'b0000000000000000010000010000000010000000 : 40'b0000000000000000000000000000000000000000;
										assign node39 = (inp[10]) ? node43 : node40;
											assign node40 = (inp[0]) ? 40'b0000000000000010010000010000000000000000 : 40'b0000000000000000000000000000000000000000;
											assign node43 = (inp[0]) ? 40'b0000000000000000000000000000000000000000 : 40'b0000000000000010010000010000000010000000;
						assign node46 = (inp[14]) ? node102 : node47;
							assign node47 = (inp[0]) ? node49 : 40'b0000000000000000000000000000000000000000;
								assign node49 = (inp[11]) ? node83 : node50;
									assign node50 = (inp[3]) ? node64 : node51;
										assign node51 = (inp[12]) ? node53 : 40'b0000000000000000000000000000000000000000;
											assign node53 = (inp[15]) ? node55 : 40'b0000000000000000000000000000000000000000;
												assign node55 = (inp[2]) ? node57 : 40'b0000000000000000000000000000000000000000;
													assign node57 = (inp[6]) ? node61 : node58;
														assign node58 = (inp[5]) ? 40'b0000000000000000000000000000000000000000 : 40'b0000000000000000000000000000000000000000;
														assign node61 = (inp[5]) ? 40'b0000000000000000000000000000000000000000 : 40'b0000000000000000010000100000000000000010;
										assign node64 = (inp[13]) ? node74 : node65;
											assign node65 = (inp[12]) ? node67 : 40'b0000000000000000000000000000000000000000;
												assign node67 = (inp[15]) ? node69 : 40'b0000000000000000000000000000000000000000;
													assign node69 = (inp[2]) ? node71 : 40'b0000000000000000000000000000000000000000;
														assign node71 = (inp[10]) ? 40'b0000000000000000000000000000000000000000 : 40'b0000000000000001010000000000000000000000;
											assign node74 = (inp[10]) ? 40'b0000000000000000000000000000001000000000 : node75;
												assign node75 = (inp[5]) ? node77 : 40'b0000000000000000000000000000000000000000;
													assign node77 = (inp[12]) ? node79 : 40'b0000000000000000000000000000000000000000;
														assign node79 = (inp[15]) ? 40'b0000000000000000000000000000000000000000 : 40'b0000000000000000000000000000000000000000;
									assign node83 = (inp[3]) ? node85 : 40'b0000000000000000000000000000000000000000;
										assign node85 = (inp[12]) ? node87 : 40'b0000000000000000000000000000000000000000;
											assign node87 = (inp[15]) ? node89 : 40'b0000000000000000000000000000000000000000;
												assign node89 = (inp[6]) ? node95 : node90;
													assign node90 = (inp[5]) ? node92 : 40'b0000000000000000000000000000000000000000;
														assign node92 = (inp[2]) ? 40'b0000000000000000000000000000000000000000 : 40'b0000000000000000000000000000000000000000;
													assign node95 = (inp[10]) ? node99 : node96;
														assign node96 = (inp[2]) ? 40'b0000000000000000000000000000000000000000 : 40'b0000000010000000010000000000010000000000;
														assign node99 = (inp[13]) ? 40'b0000000000000000000000000000000000000000 : 40'b0000000000000000000000000000000000000000;
							assign node102 = (inp[3]) ? node106 : node103;
								assign node103 = (inp[11]) ? 40'b0000000000001000010000100100000001000000 : 40'b0000000000000000010100100100000001000000;
								assign node106 = (inp[0]) ? node120 : node107;
									assign node107 = (inp[12]) ? node109 : 40'b0000000000000000000000000000000000000000;
										assign node109 = (inp[5]) ? node111 : 40'b0000000000000000000000000000000000000000;
											assign node111 = (inp[6]) ? node113 : 40'b0000000000000000000000000000000000000000;
												assign node113 = (inp[2]) ? node115 : 40'b0000000000000000000000000000000000000000;
													assign node115 = (inp[15]) ? node117 : 40'b0000000000000000000000000000000000000000;
														assign node117 = (inp[11]) ? 40'b0000000000001000000000000000000001000000 : 40'b0000000000000000000100000000000001000000;
									assign node120 = (inp[10]) ? node138 : node121;
										assign node121 = (inp[15]) ? node123 : 40'b0000000000000000000000000000000000000000;
											assign node123 = (inp[12]) ? node125 : 40'b0000000000000000000000000000000000000000;
												assign node125 = (inp[2]) ? node131 : node126;
													assign node126 = (inp[6]) ? node128 : 40'b0000000000000000000000000000000000000000;
														assign node128 = (inp[5]) ? 40'b0000000010001010010000100000000001000000 : 40'b0000000000000000000000000000000000000000;
													assign node131 = (inp[13]) ? node135 : node132;
														assign node132 = (inp[6]) ? 40'b0000000000000000000000000000000000000000 : 40'b0000000000000001010000000000001001000000;
														assign node135 = (inp[11]) ? 40'b0000000000000000000000000000000000000000 : 40'b0000000000000000000000000000000000000000;
										assign node138 = (inp[13]) ? node148 : node139;
											assign node139 = (inp[6]) ? node141 : 40'b0000000000000000000000000000000000000000;
												assign node141 = (inp[15]) ? node143 : 40'b0000000000000000000000000000000000000000;
													assign node143 = (inp[12]) ? node145 : 40'b0000000000000000000000000000000000000000;
														assign node145 = (inp[5]) ? 40'b0000000010000000010000100000000011000000 : 40'b0000000000000000000000000000000000000000;
											assign node148 = (inp[11]) ? 40'b0000000010001000000000000000000001000010 : 40'b0000000000000000000100000000001001000010;
					assign node151 = (inp[14]) ? node195 : node152;
						assign node152 = (inp[8]) ? node154 : 40'b0000000000000000000000000000000000000000;
							assign node154 = (inp[0]) ? node156 : 40'b0000000000000000000000000000000000000000;
								assign node156 = (inp[11]) ? 40'b0000000000000000000000000000000000000000 : node157;
									assign node157 = (inp[3]) ? node175 : node158;
										assign node158 = (inp[15]) ? node160 : 40'b0000000000000000000000000000000000000000;
											assign node160 = (inp[12]) ? node162 : 40'b0000000000000000000000000000000000000000;
												assign node162 = (inp[2]) ? node168 : node163;
													assign node163 = (inp[10]) ? 40'b0000000000000000000000000000000000000000 : node164;
														assign node164 = (inp[5]) ? 40'b0000000000000000000000000000000000000000 : 40'b0000000000000000000000000000000000000000;
													assign node168 = (inp[6]) ? node172 : node169;
														assign node169 = (inp[5]) ? 40'b0000000000000000000000000000000000000000 : 40'b0000000000000000000000000000000000000000;
														assign node172 = (inp[5]) ? 40'b0000000000000000000000000000000000000000 : 40'b0000000000000000000000100000000100000010;
										assign node175 = (inp[10]) ? node185 : node176;
											assign node176 = (inp[15]) ? node178 : 40'b0000000000000000000000000000000000000000;
												assign node178 = (inp[12]) ? node180 : 40'b0000000000000000000000000000000000000000;
													assign node180 = (inp[2]) ? node182 : 40'b0000000000000000000000000000000000000000;
														assign node182 = (inp[5]) ? 40'b0000000000000010000000100000001100000000 : 40'b0000000000000000000000000000000000000000;
											assign node185 = (inp[13]) ? 40'b0000000000000000000000010000000100000000 : node186;
												assign node186 = (inp[12]) ? node188 : 40'b0000000000000000000000000000000000000000;
													assign node188 = (inp[2]) ? node190 : 40'b0000000000000000000000000000000000000000;
														assign node190 = (inp[15]) ? 40'b0000000000000000000000100000000110000000 : 40'b0000000000000000000000000000000000000000;
						assign node195 = (inp[8]) ? node213 : node196;
							assign node196 = (inp[11]) ? node198 : 40'b0000000000000000000000000000000000000000;
								assign node198 = (inp[3]) ? node200 : 40'b0000000000000000000000000000000000000000;
									assign node200 = (inp[13]) ? node206 : node201;
										assign node201 = (inp[0]) ? node203 : 40'b0000000000000000000000000000000000000000;
											assign node203 = (inp[10]) ? 40'b0000000000000000000000010000000110000000 : 40'b0000000000000000000000000000000000000000;
										assign node206 = (inp[0]) ? node210 : node207;
											assign node207 = (inp[10]) ? 40'b0000000000000010000000010000000110000000 : 40'b0000000000000000000000000000000000000000;
											assign node210 = (inp[10]) ? 40'b0000000000000000000000000000000000000000 : 40'b0000000000000010000000010000000100000000;
							assign node213 = (inp[3]) ? node217 : node214;
								assign node214 = (inp[11]) ? 40'b0100000000000000000000100100000100000001 : 40'b0100000000000000000000101100000100000000;
								assign node217 = (inp[0]) ? node231 : node218;
									assign node218 = (inp[12]) ? node220 : 40'b0000000000000000000000000000000000000000;
										assign node220 = (inp[5]) ? node222 : 40'b0000000000000000000000000000000000000000;
											assign node222 = (inp[2]) ? node224 : 40'b0000000000000000000000000000000000000000;
												assign node224 = (inp[6]) ? node226 : 40'b0000000000000000000000000000000000000000;
													assign node226 = (inp[15]) ? node228 : 40'b0000000000000000000000000000000000000000;
														assign node228 = (inp[11]) ? 40'b0100000000000000000000000000000000000001 : 40'b0100000000000000000000001000000000000000;
									assign node231 = (inp[10]) ? node249 : node232;
										assign node232 = (inp[15]) ? node234 : 40'b0000000000000000000000000000000000000000;
											assign node234 = (inp[12]) ? node236 : 40'b0000000000000000000000000000000000000000;
												assign node236 = (inp[13]) ? node242 : node237;
													assign node237 = (inp[11]) ? 40'b0000000000000000000000000000000000000000 : node238;
														assign node238 = (inp[2]) ? 40'b0100000000000001000000001000000100000010 : 40'b0000000000000000000000000000000000000000;
													assign node242 = (inp[2]) ? node246 : node243;
														assign node243 = (inp[5]) ? 40'b0100000010000010000000100000000100000000 : 40'b0000000000000000000000000000000000000000;
														assign node246 = (inp[11]) ? 40'b0100000000000010000000100000000100000001 : 40'b0000000000000000000000000000000000000000;
										assign node249 = (inp[13]) ? node261 : node250;
											assign node250 = (inp[12]) ? node252 : 40'b0000000000000000000000000000000000000000;
												assign node252 = (inp[15]) ? node254 : 40'b0000000000000000000000000000000000000000;
													assign node254 = (inp[2]) ? node258 : node255;
														assign node255 = (inp[5]) ? 40'b0100000010000000000000100000000110000000 : 40'b0000000000000000000000000000000000000000;
														assign node258 = (inp[5]) ? 40'b0000000000000000000000000000000000000000 : 40'b0100000000000000000000100000000110000010;
											assign node261 = (inp[11]) ? 40'b0100000000000000000000010000000100000001 : 40'b0100000000000000000000011000000100000000;
		assign node264 = (inp[1]) ? node332 : node265;
			assign node265 = (inp[8]) ? node269 : node266;
				assign node266 = (inp[4]) ? 40'b0000000001000000000000000000000000000100 : 40'b0000000000000000000000000000000000000100;
				assign node269 = (inp[7]) ? node301 : node270;
					assign node270 = (inp[3]) ? node286 : node271;
						assign node271 = (inp[14]) ? node279 : node272;
							assign node272 = (inp[11]) ? node276 : node273;
								assign node273 = (inp[4]) ? 40'b0000000001000010010100100000001001000100 : 40'b0000000000000010010100100000001001000100;
								assign node276 = (inp[4]) ? 40'b0000000001000010010100100000000001000110 : 40'b0000000000000010010100100000000001000110;
							assign node279 = (inp[11]) ? node283 : node280;
								assign node280 = (inp[4]) ? 40'b0000000001001010010000100000001001000100 : 40'b0000000000001010010000100000001001000100;
								assign node283 = (inp[4]) ? 40'b0000000001001010010000100000000001000110 : 40'b0000000000001010010000100000000001000110;
						assign node286 = (inp[11]) ? node294 : node287;
							assign node287 = (inp[14]) ? node291 : node288;
								assign node288 = (inp[4]) ? 40'b0000000001000000010100100000001011000100 : 40'b0000000000000000010100100000001011000100;
								assign node291 = (inp[4]) ? 40'b0000000001001000010000100000001011000100 : 40'b0000000000001000010000100000001011000100;
							assign node294 = (inp[14]) ? node298 : node295;
								assign node295 = (inp[4]) ? 40'b0000000001000000010100100000000011000110 : 40'b0000000000000000010100100000000011000110;
								assign node298 = (inp[4]) ? 40'b0000000001001000010000100000000011000110 : 40'b0000000000001000010000100000000011000110;
					assign node301 = (inp[11]) ? node317 : node302;
						assign node302 = (inp[3]) ? node310 : node303;
							assign node303 = (inp[14]) ? node307 : node304;
								assign node304 = (inp[4]) ? 40'b0100000001000010000000101000001100000100 : 40'b0100000000000010000000101000001100000100;
								assign node307 = (inp[4]) ? 40'b0100000001000010000000100000001100000101 : 40'b0100000000000010000000100000001100000101;
							assign node310 = (inp[14]) ? node314 : node311;
								assign node311 = (inp[4]) ? 40'b0100000001000000000000101000001110000100 : 40'b0100000000000000000000101000001110000100;
								assign node314 = (inp[4]) ? 40'b0100000001000000000000100000001110000101 : 40'b0100000000000000000000100000001110000101;
						assign node317 = (inp[3]) ? node325 : node318;
							assign node318 = (inp[14]) ? node322 : node319;
								assign node319 = (inp[4]) ? 40'b0100000001000010000000101000000100000110 : 40'b0100000000000010000000101000000100000110;
								assign node322 = (inp[4]) ? 40'b0100000001000010000000100000000100000111 : 40'b0100000000000010000000100000000100000111;
							assign node325 = (inp[14]) ? node329 : node326;
								assign node326 = (inp[4]) ? 40'b0100000001000000000000101000000110000110 : 40'b0100000000000000000000101000000110000110;
								assign node329 = (inp[4]) ? 40'b0100000001000000000000100000000110000111 : 40'b0100000000000000000000100000000110000111;
			assign node332 = (inp[4]) ? node336 : node333;
				assign node333 = (inp[8]) ? 40'b0000000001000000000000000000000000000000 : 40'b0000100001000000000000000000000000000000;
				assign node336 = (inp[8]) ? node338 : 40'b0000100000000000000000000000000000000000;
					assign node338 = (inp[7]) ? node930 : node339;
						assign node339 = (inp[3]) ? node739 : node340;
							assign node340 = (inp[14]) ? node596 : node341;
								assign node341 = (inp[0]) ? node469 : node342;
									assign node342 = (inp[15]) ? node406 : node343;
										assign node343 = (inp[13]) ? node375 : node344;
											assign node344 = (inp[11]) ? node360 : node345;
												assign node345 = (inp[10]) ? node353 : node346;
													assign node346 = (inp[5]) ? node350 : node347;
														assign node347 = (inp[6]) ? 40'b0001000000011101010010000010101000010000 : 40'b1001000000010101010010000000101000010000;
														assign node350 = (inp[6]) ? 40'b0001000000010101010010000001101000010000 : 40'b0001000000010101010110000010101000010000;
													assign node353 = (inp[5]) ? node357 : node354;
														assign node354 = (inp[6]) ? 40'b0001000000011001010010000010101000010000 : 40'b1001000000010001010010000000101000010000;
														assign node357 = (inp[6]) ? 40'b0001000000010001010010000001101000010000 : 40'b0001000000010001010110000010101000010000;
												assign node360 = (inp[10]) ? node368 : node361;
													assign node361 = (inp[12]) ? node365 : node362;
														assign node362 = (inp[2]) ? 40'b0001000000010101010110000010101000000000 : 40'b1001000000010101010010000000101000000000;
														assign node365 = (inp[2]) ? 40'b0001000000010101010010000011101000000000 : 40'b0001000000011101010010000010101000000000;
													assign node368 = (inp[6]) ? node372 : node369;
														assign node369 = (inp[12]) ? 40'b0001000000010001010110000010101000000000 : 40'b1001000000010001010110000010101000000000;
														assign node372 = (inp[5]) ? 40'b0001000000010001010010000001101000000000 : 40'b0001000000011001010110000010101000000000;
											assign node375 = (inp[10]) ? node391 : node376;
												assign node376 = (inp[11]) ? node384 : node377;
													assign node377 = (inp[5]) ? node381 : node378;
														assign node378 = (inp[6]) ? 40'b0001000000011101010010000010001000010000 : 40'b1001000000010101010010000000001000010000;
														assign node381 = (inp[6]) ? 40'b0001000000010101010010000001001000010000 : 40'b0001000000010101010110000010001000010000;
													assign node384 = (inp[2]) ? node388 : node385;
														assign node385 = (inp[12]) ? 40'b0001000000011101010010000010001000000000 : 40'b1001000000010101010110000010001000000000;
														assign node388 = (inp[12]) ? 40'b0001000000010101010010000001001000000000 : 40'b0001000000011101010110000010001000000000;
												assign node391 = (inp[11]) ? node399 : node392;
													assign node392 = (inp[5]) ? node396 : node393;
														assign node393 = (inp[6]) ? 40'b0001000000011001010010000010001000010000 : 40'b1001000000010001010010000000001000010000;
														assign node396 = (inp[12]) ? 40'b0001000000010001010010000011001000010000 : 40'b0001000000010001010110000010001000010000;
													assign node399 = (inp[5]) ? node403 : node400;
														assign node400 = (inp[6]) ? 40'b0001000000011001010010000010001000000000 : 40'b1001000000010001010010000000001000000000;
														assign node403 = (inp[6]) ? 40'b0001000000010001010010000001001000000000 : 40'b0001000000010001010110000010001000000000;
										assign node406 = (inp[11]) ? node438 : node407;
											assign node407 = (inp[13]) ? node423 : node408;
												assign node408 = (inp[10]) ? node416 : node409;
													assign node409 = (inp[6]) ? node413 : node410;
														assign node410 = (inp[5]) ? 40'b0001000000000101010110000010101000010000 : 40'b1001000000000101010010000000101000010000;
														assign node413 = (inp[5]) ? 40'b0001000000000101010010000001101000010000 : 40'b0001000000001101010010000010101000010000;
													assign node416 = (inp[12]) ? node420 : node417;
														assign node417 = (inp[2]) ? 40'b0001000000000001010110000010101000010000 : 40'b1001000000000001010010000000101000010000;
														assign node420 = (inp[2]) ? 40'b0001000000000001010010000001101000010000 : 40'b0001000000001001010010000010101000010000;
												assign node423 = (inp[10]) ? node431 : node424;
													assign node424 = (inp[12]) ? node428 : node425;
														assign node425 = (inp[2]) ? 40'b0001000000000101010110000010001000010000 : 40'b1001000000000101010010000000001000010000;
														assign node428 = (inp[6]) ? 40'b0001000000001101010010000011001000010000 : 40'b0001000000000101010010000001001000010000;
													assign node431 = (inp[5]) ? node435 : node432;
														assign node432 = (inp[2]) ? 40'b0001000000000001010110000010001000010000 : 40'b1001000000000001010010000000001000010000;
														assign node435 = (inp[6]) ? 40'b0001000000000001010010000001001000010000 : 40'b0001000000000001010110000010001000010000;
											assign node438 = (inp[10]) ? node454 : node439;
												assign node439 = (inp[13]) ? node447 : node440;
													assign node440 = (inp[6]) ? node444 : node441;
														assign node441 = (inp[5]) ? 40'b0001000000000101010110000010101000000000 : 40'b1001000000000101010010000000101000000000;
														assign node444 = (inp[12]) ? 40'b0001000000001101010010000011101000000000 : 40'b0001000000000101010110000010101000000000;
													assign node447 = (inp[6]) ? node451 : node448;
														assign node448 = (inp[5]) ? 40'b0001000000000101010110000010001000000000 : 40'b1001000000000101010010000000001000000000;
														assign node451 = (inp[5]) ? 40'b0001000000000101010010000001001000000000 : 40'b0001000000001101010010000010001000000000;
												assign node454 = (inp[13]) ? node462 : node455;
													assign node455 = (inp[12]) ? node459 : node456;
														assign node456 = (inp[2]) ? 40'b0001000000000001010110000010101000000000 : 40'b1001000000000001010010000000101000000000;
														assign node459 = (inp[2]) ? 40'b0001000000000001010110000011101000000000 : 40'b0001000000001001010010000010101000000000;
													assign node462 = (inp[2]) ? node466 : node463;
														assign node463 = (inp[5]) ? 40'b0001000000001001010110000010001000000000 : 40'b1001000000001001010010000010001000000000;
														assign node466 = (inp[12]) ? 40'b0001000000000001010010000001001000000000 : 40'b0001000000000001010110000010001000000000;
									assign node469 = (inp[15]) ? node533 : node470;
										assign node470 = (inp[13]) ? node502 : node471;
											assign node471 = (inp[10]) ? node487 : node472;
												assign node472 = (inp[11]) ? node480 : node473;
													assign node473 = (inp[6]) ? node477 : node474;
														assign node474 = (inp[5]) ? 40'b0000000000010101010110000010101000010000 : 40'b1000000000010101010010000010101000010000;
														assign node477 = (inp[12]) ? 40'b0000000000011101010010000011101000010000 : 40'b0000000000010101010110000011101000010000;
													assign node480 = (inp[2]) ? node484 : node481;
														assign node481 = (inp[12]) ? 40'b0000000000011101010010000010101000000000 : 40'b1000000000010101010010000000101000000000;
														assign node484 = (inp[12]) ? 40'b0000000000010101010010000001101000000000 : 40'b0000000000010101010110000010101000000000;
												assign node487 = (inp[11]) ? node495 : node488;
													assign node488 = (inp[5]) ? node492 : node489;
														assign node489 = (inp[6]) ? 40'b0000000000011001010010000010101000010000 : 40'b1000000000010001010010000001101000010000;
														assign node492 = (inp[2]) ? 40'b0000000000010001010110000011101000010000 : 40'b0000000000010001010110000010101000010000;
													assign node495 = (inp[5]) ? node499 : node496;
														assign node496 = (inp[6]) ? 40'b0000000000011001010010000010101000000000 : 40'b1000000000010001010010000010101000000000;
														assign node499 = (inp[2]) ? 40'b0000000000010001010110000011101000000000 : 40'b0000000000011001010010000010101000000000;
											assign node502 = (inp[11]) ? node518 : node503;
												assign node503 = (inp[10]) ? node511 : node504;
													assign node504 = (inp[12]) ? node508 : node505;
														assign node505 = (inp[2]) ? 40'b0000000000010101010110000010001000010000 : 40'b1000000000010101010010000000001000010000;
														assign node508 = (inp[2]) ? 40'b0000000000010101010010000001001000010000 : 40'b0000000000011101010010000010001000010000;
													assign node511 = (inp[6]) ? node515 : node512;
														assign node512 = (inp[5]) ? 40'b0000000000010001010110000010001000010000 : 40'b1000000000010001010010000010001000010000;
														assign node515 = (inp[5]) ? 40'b0000000000010001010010000001001000010000 : 40'b0000000000011001010110000010001000010000;
												assign node518 = (inp[10]) ? node526 : node519;
													assign node519 = (inp[6]) ? node523 : node520;
														assign node520 = (inp[12]) ? 40'b0000000000010101010010000001001000000000 : 40'b1000000000010101010110000010001000000000;
														assign node523 = (inp[5]) ? 40'b0000000000010101010010000001001000000000 : 40'b0000000000011101010010000010001000000000;
													assign node526 = (inp[12]) ? node530 : node527;
														assign node527 = (inp[6]) ? 40'b1000000000011001010010000010001000000000 : 40'b1000000000010001010110000010001000000000;
														assign node530 = (inp[2]) ? 40'b0000000000010001010010000001001000000000 : 40'b0000000000011001010010000010001000000000;
										assign node533 = (inp[13]) ? node565 : node534;
											assign node534 = (inp[11]) ? node550 : node535;
												assign node535 = (inp[10]) ? node543 : node536;
													assign node536 = (inp[6]) ? node540 : node537;
														assign node537 = (inp[5]) ? 40'b0000000000000101010110000010101000010000 : 40'b1000000000000101010010000000101000010000;
														assign node540 = (inp[2]) ? 40'b0000000000000101010010000001101000010000 : 40'b0000000000000101010010000001101000010000;
													assign node543 = (inp[2]) ? node547 : node544;
														assign node544 = (inp[12]) ? 40'b0000000000001001010010000010101000010000 : 40'b1000000000000001010010000000101000010000;
														assign node547 = (inp[6]) ? 40'b0000000000000001010110000011101000010000 : 40'b0000000000000001010110000010101000010000;
												assign node550 = (inp[10]) ? node558 : node551;
													assign node551 = (inp[6]) ? node555 : node552;
														assign node552 = (inp[12]) ? 40'b0000000000000101010010000001101000000000 : 40'b1000000000000101010110000010101000000000;
														assign node555 = (inp[12]) ? 40'b0000000000001101010010000011101000000000 : 40'b0000000000000101010010000001101000000000;
													assign node558 = (inp[5]) ? node562 : node559;
														assign node559 = (inp[6]) ? 40'b0000000000001001010110000010101000000000 : 40'b1000000000000001010010000000101000000000;
														assign node562 = (inp[6]) ? 40'b0000000000000001010010000001101000000000 : 40'b0000000000000001010110000010101000000000;
											assign node565 = (inp[10]) ? node581 : node566;
												assign node566 = (inp[11]) ? node574 : node567;
													assign node567 = (inp[6]) ? node571 : node568;
														assign node568 = (inp[2]) ? 40'b0000000000000101010110000010001000010000 : 40'b0000000000001101010110000010001000010000;
														assign node571 = (inp[12]) ? 40'b0000000000001101010010000011001000010000 : 40'b0000000000000101010010000001001000010000;
													assign node574 = (inp[5]) ? node578 : node575;
														assign node575 = (inp[6]) ? 40'b0000000000001101010010000010001000000000 : 40'b1000000000000101010010000000001000000000;
														assign node578 = (inp[2]) ? 40'b0000000000000101010110000011001000000000 : 40'b1000000000000101010110000010001000000000;
												assign node581 = (inp[11]) ? node589 : node582;
													assign node582 = (inp[5]) ? node586 : node583;
														assign node583 = (inp[2]) ? 40'b1000000000000001010010000000001000010000 : 40'b1000000000001001010010000010001000010000;
														assign node586 = (inp[6]) ? 40'b0000000000000001010010000011001000010000 : 40'b0000000000000001010110000010001000010000;
													assign node589 = (inp[2]) ? node593 : node590;
														assign node590 = (inp[12]) ? 40'b0000000000001001010010000010001000000000 : 40'b1000000000000001010010000000001000000000;
														assign node593 = (inp[12]) ? 40'b0000000000000001010010000011001000000000 : 40'b0000000000001001010110000010001000000000;
								assign node596 = (inp[11]) ? node612 : node597;
									assign node597 = (inp[5]) ? 40'b0000000000000000000000000000000000000000 : node598;
										assign node598 = (inp[6]) ? 40'b0000000000000000000000000000000000000000 : node599;
											assign node599 = (inp[2]) ? node601 : 40'b0000000000000000000000000000000000000000;
												assign node601 = (inp[12]) ? 40'b0000000000000000000000000000000000000000 : node602;
													assign node602 = (inp[15]) ? node606 : node603;
														assign node603 = (inp[10]) ? 40'b0000000000000000000000000000000000000000 : 40'b1000000000010100001000000000000000000000;
														assign node606 = (inp[13]) ? 40'b0000000000000000000000000000000000000000 : 40'b0000000000000000000000000000000000000000;
									assign node612 = (inp[13]) ? node676 : node613;
										assign node613 = (inp[15]) ? node645 : node614;
											assign node614 = (inp[10]) ? node630 : node615;
												assign node615 = (inp[0]) ? node623 : node616;
													assign node616 = (inp[2]) ? node620 : node617;
														assign node617 = (inp[5]) ? 40'b0001010000011100000000000010100000000000 : 40'b1001010000011100000000000010100000000000;
														assign node620 = (inp[12]) ? 40'b0001010000010100000000000001100000000000 : 40'b0001010000010100000100000010100000000000;
													assign node623 = (inp[6]) ? node627 : node624;
														assign node624 = (inp[5]) ? 40'b0000010000010100000100000010100000000000 : 40'b1000010000010100000000000000100000000000;
														assign node627 = (inp[2]) ? 40'b0000010000010100000000000001100000000000 : 40'b0000010000011100000000000010100000000000;
												assign node630 = (inp[0]) ? node638 : node631;
													assign node631 = (inp[6]) ? node635 : node632;
														assign node632 = (inp[5]) ? 40'b0001010000010000000100000010100000000000 : 40'b1001010000010000000000000000100000000000;
														assign node635 = (inp[5]) ? 40'b0001010000010000000000000011100000000000 : 40'b0001010000011000000000000010100000000000;
													assign node638 = (inp[12]) ? node642 : node639;
														assign node639 = (inp[2]) ? 40'b0000010000010000000100000010100000000000 : 40'b1000010000010000000000000000100000000000;
														assign node642 = (inp[6]) ? 40'b0000010000011000000000000011100000000000 : 40'b1000010000011000000000000010100000000000;
											assign node645 = (inp[0]) ? node661 : node646;
												assign node646 = (inp[10]) ? node654 : node647;
													assign node647 = (inp[5]) ? node651 : node648;
														assign node648 = (inp[6]) ? 40'b0001010000001100000000000010100000000000 : 40'b1001010000000100000000000010100000000000;
														assign node651 = (inp[2]) ? 40'b0001010000000100000100000011100000000000 : 40'b1001010000000100000000000001100000000000;
													assign node654 = (inp[6]) ? node658 : node655;
														assign node655 = (inp[5]) ? 40'b0001010000000000000100000010100000000000 : 40'b1001010000000000000000000000100000000000;
														assign node658 = (inp[12]) ? 40'b0001010000001000000000000011100000000000 : 40'b0001010000000000000100000010100000000000;
												assign node661 = (inp[10]) ? node669 : node662;
													assign node662 = (inp[12]) ? node666 : node663;
														assign node663 = (inp[6]) ? 40'b0000010000000100000100000011100000000000 : 40'b1000010000000100000100000010100000000000;
														assign node666 = (inp[6]) ? 40'b0000010000001100000000000011100000000000 : 40'b0000010000001100000000000010100000000000;
													assign node669 = (inp[2]) ? node673 : node670;
														assign node670 = (inp[5]) ? 40'b0000010000001000000000000011100000000000 : 40'b1000010000001000000000000010100000000000;
														assign node673 = (inp[12]) ? 40'b0000010000000000000000000001100000000000 : 40'b0000010000000000000100000010100000000000;
										assign node676 = (inp[15]) ? node708 : node677;
											assign node677 = (inp[10]) ? node693 : node678;
												assign node678 = (inp[0]) ? node686 : node679;
													assign node679 = (inp[2]) ? node683 : node680;
														assign node680 = (inp[5]) ? 40'b0001010000010100000100000010000000000000 : 40'b1001010000011100000000000010000000000000;
														assign node683 = (inp[12]) ? 40'b0001010000010100000000000001000000000000 : 40'b0001010000010100000100000010000000000000;
													assign node686 = (inp[12]) ? node690 : node687;
														assign node687 = (inp[2]) ? 40'b0000010000010100000100000010000000000000 : 40'b1000010000010100000000000000000000000000;
														assign node690 = (inp[2]) ? 40'b0000010000010100000000000001000000000000 : 40'b0000010000011100000000000010000000000000;
												assign node693 = (inp[0]) ? node701 : node694;
													assign node694 = (inp[2]) ? node698 : node695;
														assign node695 = (inp[12]) ? 40'b0001010000011000000000000010000000000000 : 40'b1001010000010000000000000000000000000000;
														assign node698 = (inp[5]) ? 40'b0001010000010000000100000011000000000000 : 40'b0001010000011000000000000011000000000000;
													assign node701 = (inp[6]) ? node705 : node702;
														assign node702 = (inp[12]) ? 40'b0000010000010000000100000011000000000000 : 40'b1000010000010000000100000010000000000000;
														assign node705 = (inp[12]) ? 40'b0000010000011000000000000011000000000000 : 40'b0000010000010000000100000010000000000000;
											assign node708 = (inp[10]) ? node724 : node709;
												assign node709 = (inp[0]) ? node717 : node710;
													assign node710 = (inp[5]) ? node714 : node711;
														assign node711 = (inp[6]) ? 40'b0001010000001100000000000010000000000000 : 40'b1001010000000100000000000000000000000000;
														assign node714 = (inp[6]) ? 40'b0001010000000100000000000011000000000000 : 40'b0001010000000100000100000010000000000000;
													assign node717 = (inp[5]) ? node721 : node718;
														assign node718 = (inp[6]) ? 40'b0000010000001100000000000010000000000000 : 40'b1000010000000100000000000000000000000000;
														assign node721 = (inp[6]) ? 40'b0000010000000100000000000001000000000000 : 40'b0000010000000100000100000010000000000000;
												assign node724 = (inp[0]) ? node732 : node725;
													assign node725 = (inp[12]) ? node729 : node726;
														assign node726 = (inp[2]) ? 40'b0001010000000000000100000010000000000000 : 40'b1001010000000000000000000010000000000000;
														assign node729 = (inp[5]) ? 40'b0001010000000000000000000011000000000000 : 40'b1001010000000000000000000001000000000000;
													assign node732 = (inp[2]) ? node736 : node733;
														assign node733 = (inp[5]) ? 40'b1000010000000000000100000010000000000000 : 40'b1000010000001000000000000010000000000000;
														assign node736 = (inp[12]) ? 40'b0000010000000000000000000001000000000000 : 40'b0000010000000000000100000010000000000000;
							assign node739 = (inp[11]) ? node787 : node740;
								assign node740 = (inp[14]) ? 40'b0000000000000000000000000000000000000000 : node741;
									assign node741 = (inp[6]) ? node769 : node742;
										assign node742 = (inp[13]) ? node758 : node743;
											assign node743 = (inp[15]) ? node745 : 40'b0000000000000000000000000000000000000000;
												assign node745 = (inp[5]) ? node751 : node746;
													assign node746 = (inp[12]) ? 40'b0000000000000000000000000000000000000000 : node747;
														assign node747 = (inp[2]) ? 40'b1000000000000000000100000010100000100000 : 40'b0000000000000000000000000000000000000000;
													assign node751 = (inp[2]) ? node755 : node752;
														assign node752 = (inp[0]) ? 40'b0000000000000100000100000010100000100000 : 40'b0000000000000000000000000000000000000000;
														assign node755 = (inp[12]) ? 40'b0000000000000000000100000011100000100000 : 40'b0000000000000000000100000010100000100000;
											assign node758 = (inp[5]) ? 40'b0000000000000000000000000000000000000000 : node759;
												assign node759 = (inp[15]) ? 40'b0000000000000000000000000000000000000000 : node760;
													assign node760 = (inp[0]) ? node764 : node761;
														assign node761 = (inp[10]) ? 40'b1001000000010000000000000000000000100000 : 40'b0000000000000000000000000000000000000000;
														assign node764 = (inp[10]) ? 40'b0000000000000000000000000000000000000000 : 40'b1000000000010100000000000000000000100000;
										assign node769 = (inp[12]) ? 40'b0000000000000000000000000000000000000000 : node770;
											assign node770 = (inp[15]) ? node778 : node771;
												assign node771 = (inp[13]) ? node773 : 40'b0000000000000000000000000000000000000000;
													assign node773 = (inp[2]) ? 40'b0000000000000000000000000000000000000000 : node774;
														assign node774 = (inp[5]) ? 40'b0000000000000000000000000000000000000000 : 40'b1000000000011000000000000010000000100000;
												assign node778 = (inp[13]) ? 40'b0000000000000000000000000000000000000000 : node779;
													assign node779 = (inp[0]) ? node781 : 40'b0000000000000000000000000000000000000000;
														assign node781 = (inp[10]) ? 40'b0000000000000000000000000000000000000000 : 40'b0000000000000100000100000010100000100000;
								assign node787 = (inp[14]) ? node803 : node788;
									assign node788 = (inp[6]) ? 40'b0000000000000000000000000000000000000000 : node789;
										assign node789 = (inp[5]) ? node791 : 40'b0000000000000000000000000000000000000000;
											assign node791 = (inp[2]) ? node793 : 40'b0000000000000000000000000000000000000000;
												assign node793 = (inp[12]) ? node795 : 40'b0000000000000000000000000000000000000000;
													assign node795 = (inp[10]) ? node799 : node796;
														assign node796 = (inp[0]) ? 40'b0000000000000100001100000010000000010000 : 40'b0000000000000000000000000000000000000000;
														assign node799 = (inp[0]) ? 40'b0000000000000000000000000000000000000000 : 40'b0001000000000000001000000000100000010000;
									assign node803 = (inp[13]) ? node867 : node804;
										assign node804 = (inp[0]) ? node836 : node805;
											assign node805 = (inp[10]) ? node821 : node806;
												assign node806 = (inp[15]) ? node814 : node807;
													assign node807 = (inp[2]) ? node811 : node808;
														assign node808 = (inp[12]) ? 40'b0011000000011100000000000010100000000000 : 40'b1011000000010100000000000000100000000000;
														assign node811 = (inp[12]) ? 40'b0011000000010100000000000001100000000000 : 40'b0011000000010100000100000010100000000000;
													assign node814 = (inp[12]) ? node818 : node815;
														assign node815 = (inp[2]) ? 40'b0011000000000100000100000010100000000000 : 40'b1011000000000100000000000000100000000000;
														assign node818 = (inp[2]) ? 40'b0011000000000100000000000001100000000000 : 40'b0011000000001100000000000010100000000000;
												assign node821 = (inp[15]) ? node829 : node822;
													assign node822 = (inp[6]) ? node826 : node823;
														assign node823 = (inp[12]) ? 40'b1011000000010000000000000011100000000000 : 40'b1011000000010000000100000010100000000000;
														assign node826 = (inp[5]) ? 40'b0011000000010000000000000001100000000000 : 40'b0011000000011000000000000010100000000000;
													assign node829 = (inp[2]) ? node833 : node830;
														assign node830 = (inp[12]) ? 40'b0011000000001000000000000010100000000000 : 40'b1011000000000000000000000000100000000000;
														assign node833 = (inp[12]) ? 40'b0011000000000000000000000001100000000000 : 40'b0011000000000000000100000010100000000000;
											assign node836 = (inp[10]) ? node852 : node837;
												assign node837 = (inp[15]) ? node845 : node838;
													assign node838 = (inp[12]) ? node842 : node839;
														assign node839 = (inp[2]) ? 40'b0010000000010100000100000010100000000000 : 40'b1010000000010100000000000000100000000000;
														assign node842 = (inp[6]) ? 40'b0010000000011100000000000011100000000000 : 40'b1010000000010100000000000000100000000000;
													assign node845 = (inp[6]) ? node849 : node846;
														assign node846 = (inp[5]) ? 40'b0010000000000100000100000010100000000000 : 40'b1010000000000100000000000000100000000000;
														assign node849 = (inp[5]) ? 40'b0010000000000100000100000011100000000000 : 40'b0010000000001100000000000010100000000000;
												assign node852 = (inp[15]) ? node860 : node853;
													assign node853 = (inp[2]) ? node857 : node854;
														assign node854 = (inp[12]) ? 40'b0010000000011000000000000010100000000000 : 40'b1010000000010000000000000000100000000000;
														assign node857 = (inp[12]) ? 40'b0010000000010000000000000001100000000000 : 40'b0010000000010000000100000010100000000000;
													assign node860 = (inp[2]) ? node864 : node861;
														assign node861 = (inp[12]) ? 40'b0010000000001000000000000010100000000000 : 40'b1010000000000000000000000000100000000000;
														assign node864 = (inp[5]) ? 40'b0010000000000000000100000011100000000000 : 40'b1010000000000000000100000010100000000000;
										assign node867 = (inp[10]) ? node899 : node868;
											assign node868 = (inp[0]) ? node884 : node869;
												assign node869 = (inp[15]) ? node877 : node870;
													assign node870 = (inp[5]) ? node874 : node871;
														assign node871 = (inp[2]) ? 40'b0011000000011100000100000010000000000000 : 40'b1011000000011100000000000010000000000000;
														assign node874 = (inp[6]) ? 40'b0011000000010100000000000001000000000000 : 40'b0011000000010100000100000010000000000000;
													assign node877 = (inp[12]) ? node881 : node878;
														assign node878 = (inp[5]) ? 40'b0011000000000100000100000010000000000000 : 40'b0011000000001100000100000010000000000000;
														assign node881 = (inp[2]) ? 40'b0011000000000100000000000001000000000000 : 40'b0011000000001100000000000010000000000000;
												assign node884 = (inp[5]) ? node892 : node885;
													assign node885 = (inp[6]) ? node889 : node886;
														assign node886 = (inp[2]) ? 40'b1010000000010100000100000010000000000000 : 40'b1010000000001100000000000010000000000000;
														assign node889 = (inp[15]) ? 40'b0010000000001100000000000010000000000000 : 40'b0010000000011100000000000010000000000000;
													assign node892 = (inp[6]) ? node896 : node893;
														assign node893 = (inp[12]) ? 40'b0010000000000100000100000011000000000000 : 40'b0010000000010100000100000010000000000000;
														assign node896 = (inp[12]) ? 40'b0010000000010100000000000001000000000000 : 40'b0010000000010100000100000011000000000000;
											assign node899 = (inp[15]) ? node915 : node900;
												assign node900 = (inp[5]) ? node908 : node901;
													assign node901 = (inp[6]) ? node905 : node902;
														assign node902 = (inp[2]) ? 40'b1010000000010000000100000010000000000000 : 40'b1011000000010000000000000000000000000000;
														assign node905 = (inp[0]) ? 40'b0010000000011000000000000010000000000000 : 40'b0011000000011000000000000010000000000000;
													assign node908 = (inp[0]) ? node912 : node909;
														assign node909 = (inp[2]) ? 40'b0011000000010000000100000011000000000000 : 40'b0011000000010000000000000001000000000000;
														assign node912 = (inp[6]) ? 40'b0010000000010000000000000001000000000000 : 40'b0010000000010000000100000010000000000000;
												assign node915 = (inp[0]) ? node923 : node916;
													assign node916 = (inp[12]) ? node920 : node917;
														assign node917 = (inp[5]) ? 40'b0011000000000000000100000010000000000000 : 40'b0011000000000000000100000010000000000000;
														assign node920 = (inp[2]) ? 40'b0011000000000000000000000001000000000000 : 40'b0011000000001000000000000010000000000000;
													assign node923 = (inp[2]) ? node927 : node924;
														assign node924 = (inp[12]) ? 40'b0010000000001000000000000010000000000000 : 40'b1010000000000000000000000001000000000000;
														assign node927 = (inp[12]) ? 40'b0010000000000000000000000001000000000000 : 40'b0010000000000000000100000010000000000000;
						assign node930 = (inp[3]) ? node1004 : node931;
							assign node931 = (inp[14]) ? node957 : node932;
								assign node932 = (inp[11]) ? node934 : 40'b0000000000000000000000000000000000000000;
									assign node934 = (inp[15]) ? node946 : node935;
										assign node935 = (inp[0]) ? node941 : node936;
											assign node936 = (inp[10]) ? node938 : 40'b0000000000000000000000000000000000000000;
												assign node938 = (inp[13]) ? 40'b1001001000010000000000000000000000001000 : 40'b1001001000010000000000000000100000001000;
											assign node941 = (inp[10]) ? 40'b0000000000000000000000000000000000000000 : node942;
												assign node942 = (inp[13]) ? 40'b1000001000010100000000000000000000001000 : 40'b1000001000010100000000000000100000001000;
										assign node946 = (inp[10]) ? node952 : node947;
											assign node947 = (inp[0]) ? node949 : 40'b0000000000000000000000000000000000000000;
												assign node949 = (inp[13]) ? 40'b0000001000000100000100000010000000001000 : 40'b0000001000000100000100000010100000001000;
											assign node952 = (inp[0]) ? 40'b0000000000000000000000000000000000000000 : node953;
												assign node953 = (inp[13]) ? 40'b0001001000000000000100000010000000001000 : 40'b0001001000000000000100000010100000001000;
								assign node957 = (inp[11]) ? 40'b0000000000000000000000000000000000000000 : node958;
									assign node958 = (inp[15]) ? node972 : node959;
										assign node959 = (inp[13]) ? node961 : 40'b0000000000000000000000000000000000000000;
											assign node961 = (inp[10]) ? node963 : 40'b0000000000000000000000000000000000000000;
												assign node963 = (inp[0]) ? node965 : 40'b0000000000000000000000000000000000000000;
													assign node965 = (inp[6]) ? node969 : node966;
														assign node966 = (inp[5]) ? 40'b0000001100010000000100000010000000000000 : 40'b1000001100010000000000000000000000000000;
														assign node969 = (inp[5]) ? 40'b0000001100010000000000000001000000000000 : 40'b0000001100011000000000000010000000000000;
										assign node972 = (inp[0]) ? node984 : node973;
											assign node973 = (inp[13]) ? node975 : 40'b0000000000000000000000000000000000000000;
												assign node975 = (inp[10]) ? node977 : 40'b0000000000000000000000000000000000000000;
													assign node977 = (inp[5]) ? node981 : node978;
														assign node978 = (inp[2]) ? 40'b0001001100001000000000000011000000000000 : 40'b1001001100001000000000000010000000000000;
														assign node981 = (inp[6]) ? 40'b0001001100000000000000000001000000000000 : 40'b0001001100000000000100000010000000000000;
											assign node984 = (inp[13]) ? node994 : node985;
												assign node985 = (inp[10]) ? node987 : 40'b0000000000000000000000000000000000000000;
													assign node987 = (inp[5]) ? node991 : node988;
														assign node988 = (inp[12]) ? 40'b1000001100001000000000000011100000000000 : 40'b1000001100001000000100000010100000000000;
														assign node991 = (inp[12]) ? 40'b0000001100001000000100000011100000000000 : 40'b1000001100000000000100000011100000000000;
												assign node994 = (inp[10]) ? 40'b0000000000000000000000000000000000000000 : node995;
													assign node995 = (inp[5]) ? node999 : node996;
														assign node996 = (inp[6]) ? 40'b0000001100001100000000000010000000000000 : 40'b1000001100000100000000000010000000000000;
														assign node999 = (inp[6]) ? 40'b0000001100000100000000000001000000000000 : 40'b0000001100000100000100000010000000000000;
							assign node1004 = (inp[13]) ? node1136 : node1005;
								assign node1005 = (inp[14]) ? node1071 : node1006;
									assign node1006 = (inp[11]) ? node1008 : 40'b0000000000000000000000000000000000000000;
										assign node1008 = (inp[0]) ? node1040 : node1009;
											assign node1009 = (inp[15]) ? node1025 : node1010;
												assign node1010 = (inp[10]) ? node1018 : node1011;
													assign node1011 = (inp[5]) ? node1015 : node1012;
														assign node1012 = (inp[6]) ? 40'b0001001000011100000000000010100000001000 : 40'b1001001000010100000000000000100000001000;
														assign node1015 = (inp[12]) ? 40'b0001001000011100000100000011100000001000 : 40'b1001001000010100000100000011100000001000;
													assign node1018 = (inp[6]) ? node1022 : node1019;
														assign node1019 = (inp[5]) ? 40'b0001001000010000000100000010100000001000 : 40'b1001001000010000000000000000100000001000;
														assign node1022 = (inp[5]) ? 40'b0001001000010000000000000001100000001000 : 40'b0001001000011000000000000010100000001000;
												assign node1025 = (inp[10]) ? node1033 : node1026;
													assign node1026 = (inp[12]) ? node1030 : node1027;
														assign node1027 = (inp[2]) ? 40'b0001001000000100000100000010100000001000 : 40'b1001001000000100000000000010100000001000;
														assign node1030 = (inp[6]) ? 40'b0001001000001100000000000011100000001000 : 40'b0001001000000100000100000010100000001000;
													assign node1033 = (inp[2]) ? node1037 : node1034;
														assign node1034 = (inp[5]) ? 40'b0001001000000000000000000001100000001000 : 40'b1001001000001000000000000010100000001000;
														assign node1037 = (inp[12]) ? 40'b0001001000000000000000000001100000001000 : 40'b0001001000000000000100000010100000001000;
											assign node1040 = (inp[15]) ? node1056 : node1041;
												assign node1041 = (inp[10]) ? node1049 : node1042;
													assign node1042 = (inp[5]) ? node1046 : node1043;
														assign node1043 = (inp[6]) ? 40'b0000001000011100000000000010100000001000 : 40'b1000001000010100000000000010100000001000;
														assign node1046 = (inp[6]) ? 40'b0000001000010100000000000001100000001000 : 40'b0000001000010100000100000010100000001000;
													assign node1049 = (inp[5]) ? node1053 : node1050;
														assign node1050 = (inp[2]) ? 40'b0000001000010000000100000010100000001000 : 40'b1000001000011000000000000010100000001000;
														assign node1053 = (inp[6]) ? 40'b0000001000010000000000000001100000001000 : 40'b0000001000010000000100000010100000001000;
												assign node1056 = (inp[10]) ? node1064 : node1057;
													assign node1057 = (inp[2]) ? node1061 : node1058;
														assign node1058 = (inp[12]) ? 40'b0000001000001100000000000010100000001000 : 40'b1000001000000100000000000000100000001000;
														assign node1061 = (inp[5]) ? 40'b0000001000000100000100000011100000001000 : 40'b1000001000000100000000000000100000001000;
													assign node1064 = (inp[5]) ? node1068 : node1065;
														assign node1065 = (inp[6]) ? 40'b0000001000001000000100000010100000001000 : 40'b1000001000000000000000000010100000001000;
														assign node1068 = (inp[6]) ? 40'b0000001000000000000000000001100000001000 : 40'b0000001000000000000100000010100000001000;
									assign node1071 = (inp[11]) ? 40'b0000000000000000000000000000000000000000 : node1072;
										assign node1072 = (inp[10]) ? node1104 : node1073;
											assign node1073 = (inp[0]) ? node1089 : node1074;
												assign node1074 = (inp[15]) ? node1082 : node1075;
													assign node1075 = (inp[2]) ? node1079 : node1076;
														assign node1076 = (inp[12]) ? 40'b0001001000011100000000000010100000000000 : 40'b1001001000010100000000000000100000000000;
														assign node1079 = (inp[12]) ? 40'b0001001000010100000000000011100000000000 : 40'b0001001000010100000100000010100000000000;
													assign node1082 = (inp[5]) ? node1086 : node1083;
														assign node1083 = (inp[6]) ? 40'b0001001000001100000000000010100000000000 : 40'b1001001000000100000000000000100000000000;
														assign node1086 = (inp[6]) ? 40'b0001001000000100000000000001100000000000 : 40'b0001001000000100000100000010100000000000;
												assign node1089 = (inp[15]) ? node1097 : node1090;
													assign node1090 = (inp[2]) ? node1094 : node1091;
														assign node1091 = (inp[6]) ? 40'b0000001000011100000000000011100000000000 : 40'b0000001000011100000000000010100000000000;
														assign node1094 = (inp[12]) ? 40'b0000001000010100000000000001100000000000 : 40'b0000001000010100000100000010100000000000;
													assign node1097 = (inp[12]) ? node1101 : node1098;
														assign node1098 = (inp[6]) ? 40'b0000001000001100000100000010100000000000 : 40'b1000001000000100000100000010100000000000;
														assign node1101 = (inp[2]) ? 40'b0000001000000100000000000011100000000000 : 40'b0000001000001100000000000010100000000000;
											assign node1104 = (inp[15]) ? node1120 : node1105;
												assign node1105 = (inp[0]) ? node1113 : node1106;
													assign node1106 = (inp[5]) ? node1110 : node1107;
														assign node1107 = (inp[2]) ? 40'b0001001000011000000100000010100000000000 : 40'b1001001000011000000000000010100000000000;
														assign node1110 = (inp[2]) ? 40'b0001001000010000000000000001100000000000 : 40'b0001001000011000000000000011100000000000;
													assign node1113 = (inp[5]) ? node1117 : node1114;
														assign node1114 = (inp[6]) ? 40'b0000001000011000000000000010100000000000 : 40'b1000001000010000000000000010100000000000;
														assign node1117 = (inp[6]) ? 40'b0000001000010000000000000001100000000000 : 40'b0000001000010000000100000010100000000000;
												assign node1120 = (inp[0]) ? node1128 : node1121;
													assign node1121 = (inp[12]) ? node1125 : node1122;
														assign node1122 = (inp[2]) ? 40'b0001001000000000000100000010100000000000 : 40'b1001001000000000000000000000100000000000;
														assign node1125 = (inp[2]) ? 40'b0001001000000000000000000001100000000000 : 40'b0001001000001000000000000010100000000000;
													assign node1128 = (inp[6]) ? node1132 : node1129;
														assign node1129 = (inp[12]) ? 40'b0000001000001000000000000010100000000000 : 40'b1000001000000000000100000010100000000000;
														assign node1132 = (inp[5]) ? 40'b0000001000000000000000000001100000000000 : 40'b0000001000001000000000000010100000000000;
								assign node1136 = (inp[0]) ? node1204 : node1137;
									assign node1137 = (inp[11]) ? node1171 : node1138;
										assign node1138 = (inp[14]) ? node1140 : 40'b0000000000000000000000000000000000000000;
											assign node1140 = (inp[15]) ? node1156 : node1141;
												assign node1141 = (inp[10]) ? node1149 : node1142;
													assign node1142 = (inp[6]) ? node1146 : node1143;
														assign node1143 = (inp[5]) ? 40'b0001001000010100000100000010000000000000 : 40'b1001001000010100000000000010000000000000;
														assign node1146 = (inp[12]) ? 40'b0001001000011100000000000011000000000000 : 40'b0001001000011100000000000010000000000000;
													assign node1149 = (inp[5]) ? node1153 : node1150;
														assign node1150 = (inp[12]) ? 40'b1001001000010000000000000001000000000000 : 40'b1001001000010000000000000010000000000000;
														assign node1153 = (inp[2]) ? 40'b0001001000010000000100000011000000000000 : 40'b1001001000010000000100000010000000000000;
												assign node1156 = (inp[10]) ? node1164 : node1157;
													assign node1157 = (inp[12]) ? node1161 : node1158;
														assign node1158 = (inp[6]) ? 40'b0001001000000100000000000001000000000000 : 40'b1001001000000100000100000010000000000000;
														assign node1161 = (inp[2]) ? 40'b0001001000000100000000000001000000000000 : 40'b0001001000001100000000000010000000000000;
													assign node1164 = (inp[2]) ? node1168 : node1165;
														assign node1165 = (inp[12]) ? 40'b0001001000001000000000000010000000000000 : 40'b1001001000000000000000000010000000000000;
														assign node1168 = (inp[12]) ? 40'b0001001000000000000000000001000000000000 : 40'b0001001000000000000100000010000000000000;
										assign node1171 = (inp[14]) ? 40'b0000000000000000000000000000000000000000 : node1172;
											assign node1172 = (inp[15]) ? node1188 : node1173;
												assign node1173 = (inp[10]) ? node1181 : node1174;
													assign node1174 = (inp[6]) ? node1178 : node1175;
														assign node1175 = (inp[5]) ? 40'b0001001000010100000100000010000000001000 : 40'b1001001000010100000000000001000000001000;
														assign node1178 = (inp[5]) ? 40'b0001001000010100000000000001000000001000 : 40'b0001001000011100000000000010000000001000;
													assign node1181 = (inp[6]) ? node1185 : node1182;
														assign node1182 = (inp[5]) ? 40'b0001001000010000000100000010000000001000 : 40'b1001001000010000000000000000000000001000;
														assign node1185 = (inp[12]) ? 40'b0001001000011000000000000011000000001000 : 40'b1001001000010000000000000000000000001000;
												assign node1188 = (inp[2]) ? node1196 : node1189;
													assign node1189 = (inp[10]) ? node1193 : node1190;
														assign node1190 = (inp[5]) ? 40'b0001001000001100000000000010000000001000 : 40'b1001001000001100000000000010000000001000;
														assign node1193 = (inp[5]) ? 40'b0001001000000000000100000010000000001000 : 40'b1001001000001000000000000010000000001000;
													assign node1196 = (inp[12]) ? node1200 : node1197;
														assign node1197 = (inp[10]) ? 40'b0001001000000000000100000010000000001000 : 40'b0001001000000100000100000010000000001000;
														assign node1200 = (inp[10]) ? 40'b0001001000000000000000000011000000001000 : 40'b0001001000000100000000000001000000001000;
									assign node1204 = (inp[15]) ? node1240 : node1205;
										assign node1205 = (inp[14]) ? node1223 : node1206;
											assign node1206 = (inp[11]) ? node1208 : 40'b0000000000000000000000000000000000000000;
												assign node1208 = (inp[10]) ? node1216 : node1209;
													assign node1209 = (inp[6]) ? node1213 : node1210;
														assign node1210 = (inp[5]) ? 40'b0000001000010100000100000010000000001000 : 40'b1000001000010100000000000010000000001000;
														assign node1213 = (inp[12]) ? 40'b0000001000011100000000000011000000001000 : 40'b0000001000011100000000000010000000001000;
													assign node1216 = (inp[6]) ? node1220 : node1217;
														assign node1217 = (inp[2]) ? 40'b1000001000010000000000000001000000001000 : 40'b1000001000011000000100000010000000001000;
														assign node1220 = (inp[5]) ? 40'b0000001000010000000000000001000000001000 : 40'b0000001000011000000000000010000000001000;
											assign node1223 = (inp[11]) ? 40'b0000000000000000000000000000000000000000 : node1224;
												assign node1224 = (inp[10]) ? node1232 : node1225;
													assign node1225 = (inp[12]) ? node1229 : node1226;
														assign node1226 = (inp[2]) ? 40'b0000001000010100000100000010000000000000 : 40'b1000001000010100000000000000000000000000;
														assign node1229 = (inp[6]) ? 40'b0000001000011100000000000011000000000000 : 40'b0000001000010100000100000010000000000000;
													assign node1232 = (inp[5]) ? node1236 : node1233;
														assign node1233 = (inp[6]) ? 40'b0000001000011000000100000010000000000000 : 40'b1000001000010000000000000000000000000000;
														assign node1236 = (inp[6]) ? 40'b0000001000010000000000000001000000000000 : 40'b0000001000010000000100000010000000000000;
										assign node1240 = (inp[14]) ? node1258 : node1241;
											assign node1241 = (inp[11]) ? node1243 : 40'b0000000000000000000000000000000000000000;
												assign node1243 = (inp[10]) ? node1251 : node1244;
													assign node1244 = (inp[5]) ? node1248 : node1245;
														assign node1245 = (inp[6]) ? 40'b0000001000001100000000000010000000001000 : 40'b1000001000000100000000000000000000001000;
														assign node1248 = (inp[12]) ? 40'b0000001000000100000000000011000000001000 : 40'b1000001000000100000000000001000000001000;
													assign node1251 = (inp[12]) ? node1255 : node1252;
														assign node1252 = (inp[2]) ? 40'b0000001000000000000100000010000000001000 : 40'b1000001000000000000000000010000000001000;
														assign node1255 = (inp[2]) ? 40'b0000001000000000000000000011000000001000 : 40'b0000001000001000000000000010000000001000;
											assign node1258 = (inp[11]) ? 40'b0000000000000000000000000000000000000000 : node1259;
												assign node1259 = (inp[10]) ? node1267 : node1260;
													assign node1260 = (inp[2]) ? node1264 : node1261;
														assign node1261 = (inp[6]) ? 40'b1000001000000100000000000001000000000000 : 40'b1000001000000100000100000010000000000000;
														assign node1264 = (inp[5]) ? 40'b0000001000000100000100000011000000000000 : 40'b0000001000001100000000000011000000000000;
													assign node1267 = (inp[5]) ? node1271 : node1268;
														assign node1268 = (inp[6]) ? 40'b0000001000001000000000000010000000000000 : 40'b1000001000000000000000000010000000000000;
														assign node1271 = (inp[6]) ? 40'b0000001000000000000000000001000000000000 : 40'b0000001000000000000100000010000000000000;

endmodule