module dtc_split75_bm60 (
	input  wire [12-1:0] inp,
	output wire [3-1:0] outp
);

	wire [3-1:0] node1;
	wire [3-1:0] node2;
	wire [3-1:0] node3;
	wire [3-1:0] node5;
	wire [3-1:0] node7;
	wire [3-1:0] node8;
	wire [3-1:0] node10;
	wire [3-1:0] node12;
	wire [3-1:0] node14;
	wire [3-1:0] node17;
	wire [3-1:0] node18;
	wire [3-1:0] node20;
	wire [3-1:0] node22;
	wire [3-1:0] node26;
	wire [3-1:0] node28;
	wire [3-1:0] node30;
	wire [3-1:0] node31;
	wire [3-1:0] node33;
	wire [3-1:0] node37;
	wire [3-1:0] node38;
	wire [3-1:0] node39;
	wire [3-1:0] node40;
	wire [3-1:0] node42;
	wire [3-1:0] node44;
	wire [3-1:0] node47;
	wire [3-1:0] node48;
	wire [3-1:0] node49;
	wire [3-1:0] node51;
	wire [3-1:0] node53;
	wire [3-1:0] node58;
	wire [3-1:0] node59;
	wire [3-1:0] node62;
	wire [3-1:0] node65;
	wire [3-1:0] node66;
	wire [3-1:0] node68;
	wire [3-1:0] node69;
	wire [3-1:0] node71;
	wire [3-1:0] node72;
	wire [3-1:0] node74;
	wire [3-1:0] node78;
	wire [3-1:0] node80;
	wire [3-1:0] node82;
	wire [3-1:0] node84;
	wire [3-1:0] node87;
	wire [3-1:0] node89;
	wire [3-1:0] node90;
	wire [3-1:0] node92;
	wire [3-1:0] node96;
	wire [3-1:0] node97;
	wire [3-1:0] node98;
	wire [3-1:0] node99;
	wire [3-1:0] node101;
	wire [3-1:0] node102;
	wire [3-1:0] node104;
	wire [3-1:0] node106;
	wire [3-1:0] node108;
	wire [3-1:0] node112;
	wire [3-1:0] node113;
	wire [3-1:0] node114;
	wire [3-1:0] node115;
	wire [3-1:0] node117;
	wire [3-1:0] node119;
	wire [3-1:0] node125;
	wire [3-1:0] node126;
	wire [3-1:0] node127;
	wire [3-1:0] node129;
	wire [3-1:0] node131;
	wire [3-1:0] node135;
	wire [3-1:0] node137;
	wire [3-1:0] node138;
	wire [3-1:0] node140;
	wire [3-1:0] node142;
	wire [3-1:0] node144;
	wire [3-1:0] node148;
	wire [3-1:0] node149;
	wire [3-1:0] node150;
	wire [3-1:0] node152;
	wire [3-1:0] node153;
	wire [3-1:0] node155;
	wire [3-1:0] node157;
	wire [3-1:0] node159;
	wire [3-1:0] node162;
	wire [3-1:0] node163;
	wire [3-1:0] node165;
	wire [3-1:0] node167;
	wire [3-1:0] node171;
	wire [3-1:0] node173;
	wire [3-1:0] node174;
	wire [3-1:0] node176;
	wire [3-1:0] node180;
	wire [3-1:0] node181;
	wire [3-1:0] node182;
	wire [3-1:0] node183;
	wire [3-1:0] node184;
	wire [3-1:0] node186;
	wire [3-1:0] node188;
	wire [3-1:0] node192;
	wire [3-1:0] node194;
	wire [3-1:0] node196;
	wire [3-1:0] node198;
	wire [3-1:0] node201;
	wire [3-1:0] node203;
	wire [3-1:0] node205;
	wire [3-1:0] node208;
	wire [3-1:0] node209;
	wire [3-1:0] node210;
	wire [3-1:0] node212;
	wire [3-1:0] node214;
	wire [3-1:0] node216;
	wire [3-1:0] node219;
	wire [3-1:0] node220;
	wire [3-1:0] node222;
	wire [3-1:0] node224;
	wire [3-1:0] node228;
	wire [3-1:0] node229;
	wire [3-1:0] node231;
	wire [3-1:0] node234;
	wire [3-1:0] node235;
	wire [3-1:0] node237;
	wire [3-1:0] node239;
	wire [3-1:0] node242;
	wire [3-1:0] node244;
	wire [3-1:0] node246;

	assign outp = (inp[2]) ? node96 : node1;
		assign node1 = (inp[4]) ? node37 : node2;
			assign node2 = (inp[10]) ? node26 : node3;
				assign node3 = (inp[5]) ? node5 : 3'b111;
					assign node5 = (inp[9]) ? node7 : 3'b111;
						assign node7 = (inp[7]) ? node17 : node8;
							assign node8 = (inp[8]) ? node10 : 3'b111;
								assign node10 = (inp[11]) ? node12 : 3'b111;
									assign node12 = (inp[6]) ? node14 : 3'b111;
										assign node14 = (inp[3]) ? 3'b110 : 3'b111;
							assign node17 = (inp[3]) ? 3'b110 : node18;
								assign node18 = (inp[6]) ? node20 : 3'b111;
									assign node20 = (inp[11]) ? node22 : 3'b111;
										assign node22 = (inp[8]) ? 3'b110 : 3'b111;
				assign node26 = (inp[5]) ? node28 : 3'b110;
					assign node28 = (inp[9]) ? node30 : 3'b110;
						assign node30 = (inp[3]) ? 3'b011 : node31;
							assign node31 = (inp[8]) ? node33 : 3'b110;
								assign node33 = (inp[7]) ? 3'b111 : 3'b110;
			assign node37 = (inp[3]) ? node65 : node38;
				assign node38 = (inp[5]) ? node58 : node39;
					assign node39 = (inp[10]) ? node47 : node40;
						assign node40 = (inp[7]) ? node42 : 3'b110;
							assign node42 = (inp[8]) ? node44 : 3'b110;
								assign node44 = (inp[9]) ? 3'b111 : 3'b110;
						assign node47 = (inp[7]) ? 3'b110 : node48;
							assign node48 = (inp[9]) ? 3'b110 : node49;
								assign node49 = (inp[8]) ? node51 : 3'b111;
									assign node51 = (inp[6]) ? node53 : 3'b111;
										assign node53 = (inp[11]) ? 3'b110 : 3'b111;
					assign node58 = (inp[9]) ? node62 : node59;
						assign node59 = (inp[10]) ? 3'b110 : 3'b111;
						assign node62 = (inp[10]) ? 3'b011 : 3'b111;
				assign node65 = (inp[5]) ? node87 : node66;
					assign node66 = (inp[9]) ? node68 : 3'b011;
						assign node68 = (inp[7]) ? node78 : node69;
							assign node69 = (inp[11]) ? node71 : 3'b011;
								assign node71 = (inp[10]) ? 3'b011 : node72;
									assign node72 = (inp[8]) ? node74 : 3'b011;
										assign node74 = (inp[6]) ? 3'b010 : 3'b011;
							assign node78 = (inp[10]) ? node80 : 3'b010;
								assign node80 = (inp[6]) ? node82 : 3'b011;
									assign node82 = (inp[8]) ? node84 : 3'b011;
										assign node84 = (inp[11]) ? 3'b010 : 3'b011;
					assign node87 = (inp[9]) ? node89 : 3'b010;
						assign node89 = (inp[10]) ? 3'b010 : node90;
							assign node90 = (inp[7]) ? node92 : 3'b010;
								assign node92 = (inp[8]) ? 3'b011 : 3'b010;
		assign node96 = (inp[4]) ? node148 : node97;
			assign node97 = (inp[10]) ? node125 : node98;
				assign node98 = (inp[5]) ? node112 : node99;
					assign node99 = (inp[3]) ? node101 : 3'b011;
						assign node101 = (inp[9]) ? 3'b010 : node102;
							assign node102 = (inp[7]) ? node104 : 3'b011;
								assign node104 = (inp[8]) ? node106 : 3'b011;
									assign node106 = (inp[6]) ? node108 : 3'b011;
										assign node108 = (inp[11]) ? 3'b010 : 3'b011;
					assign node112 = (inp[7]) ? 3'b010 : node113;
						assign node113 = (inp[3]) ? 3'b010 : node114;
							assign node114 = (inp[9]) ? 3'b010 : node115;
								assign node115 = (inp[6]) ? node117 : 3'b011;
									assign node117 = (inp[11]) ? node119 : 3'b011;
										assign node119 = (inp[8]) ? 3'b010 : 3'b011;
				assign node125 = (inp[3]) ? node135 : node126;
					assign node126 = (inp[5]) ? 3'b011 : node127;
						assign node127 = (inp[9]) ? node129 : 3'b010;
							assign node129 = (inp[7]) ? node131 : 3'b010;
								assign node131 = (inp[8]) ? 3'b011 : 3'b010;
					assign node135 = (inp[5]) ? node137 : 3'b111;
						assign node137 = (inp[9]) ? 3'b110 : node138;
							assign node138 = (inp[11]) ? node140 : 3'b111;
								assign node140 = (inp[7]) ? node142 : 3'b111;
									assign node142 = (inp[8]) ? node144 : 3'b111;
										assign node144 = (inp[6]) ? 3'b110 : 3'b111;
			assign node148 = (inp[3]) ? node180 : node149;
				assign node149 = (inp[5]) ? node171 : node150;
					assign node150 = (inp[9]) ? node152 : 3'b101;
						assign node152 = (inp[7]) ? node162 : node153;
							assign node153 = (inp[8]) ? node155 : 3'b101;
								assign node155 = (inp[10]) ? node157 : 3'b101;
									assign node157 = (inp[11]) ? node159 : 3'b101;
										assign node159 = (inp[6]) ? 3'b100 : 3'b101;
							assign node162 = (inp[10]) ? 3'b100 : node163;
								assign node163 = (inp[8]) ? node165 : 3'b101;
									assign node165 = (inp[6]) ? node167 : 3'b101;
										assign node167 = (inp[11]) ? 3'b100 : 3'b101;
					assign node171 = (inp[9]) ? node173 : 3'b100;
						assign node173 = (inp[10]) ? 3'b001 : node174;
							assign node174 = (inp[8]) ? node176 : 3'b100;
								assign node176 = (inp[7]) ? 3'b101 : 3'b100;
				assign node180 = (inp[10]) ? node208 : node181;
					assign node181 = (inp[9]) ? node201 : node182;
						assign node182 = (inp[5]) ? node192 : node183;
							assign node183 = (inp[7]) ? 3'b000 : node184;
								assign node184 = (inp[11]) ? node186 : 3'b001;
									assign node186 = (inp[8]) ? node188 : 3'b001;
										assign node188 = (inp[6]) ? 3'b000 : 3'b001;
							assign node192 = (inp[7]) ? node194 : 3'b001;
								assign node194 = (inp[8]) ? node196 : 3'b001;
									assign node196 = (inp[11]) ? node198 : 3'b001;
										assign node198 = (inp[6]) ? 3'b000 : 3'b001;
						assign node201 = (inp[8]) ? node203 : 3'b000;
							assign node203 = (inp[7]) ? node205 : 3'b000;
								assign node205 = (inp[5]) ? 3'b000 : 3'b001;
					assign node208 = (inp[9]) ? node228 : node209;
						assign node209 = (inp[7]) ? node219 : node210;
							assign node210 = (inp[8]) ? node212 : 3'b101;
								assign node212 = (inp[6]) ? node214 : 3'b101;
									assign node214 = (inp[5]) ? node216 : 3'b101;
										assign node216 = (inp[11]) ? 3'b100 : 3'b101;
							assign node219 = (inp[5]) ? 3'b100 : node220;
								assign node220 = (inp[6]) ? node222 : 3'b101;
									assign node222 = (inp[8]) ? node224 : 3'b101;
										assign node224 = (inp[11]) ? 3'b100 : 3'b101;
						assign node228 = (inp[5]) ? node234 : node229;
							assign node229 = (inp[8]) ? node231 : 3'b100;
								assign node231 = (inp[7]) ? 3'b101 : 3'b100;
							assign node234 = (inp[7]) ? node242 : node235;
								assign node235 = (inp[6]) ? node237 : 3'b001;
									assign node237 = (inp[11]) ? node239 : 3'b001;
										assign node239 = (inp[8]) ? 3'b000 : 3'b001;
								assign node242 = (inp[8]) ? node244 : 3'b000;
									assign node244 = (inp[11]) ? node246 : 3'b001;
										assign node246 = (inp[6]) ? 3'b000 : 3'b001;

endmodule