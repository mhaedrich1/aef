module dtc_split25_bm60 (
	input  wire [12-1:0] inp,
	output wire [3-1:0] outp
);

	wire [3-1:0] node1;
	wire [3-1:0] node2;
	wire [3-1:0] node3;
	wire [3-1:0] node5;
	wire [3-1:0] node7;
	wire [3-1:0] node9;
	wire [3-1:0] node10;
	wire [3-1:0] node12;
	wire [3-1:0] node13;
	wire [3-1:0] node17;
	wire [3-1:0] node18;
	wire [3-1:0] node19;
	wire [3-1:0] node24;
	wire [3-1:0] node26;
	wire [3-1:0] node28;
	wire [3-1:0] node29;
	wire [3-1:0] node33;
	wire [3-1:0] node34;
	wire [3-1:0] node35;
	wire [3-1:0] node36;
	wire [3-1:0] node37;
	wire [3-1:0] node38;
	wire [3-1:0] node43;
	wire [3-1:0] node44;
	wire [3-1:0] node46;
	wire [3-1:0] node47;
	wire [3-1:0] node51;
	wire [3-1:0] node52;
	wire [3-1:0] node56;
	wire [3-1:0] node57;
	wire [3-1:0] node60;
	wire [3-1:0] node63;
	wire [3-1:0] node64;
	wire [3-1:0] node65;
	wire [3-1:0] node67;
	wire [3-1:0] node68;
	wire [3-1:0] node70;
	wire [3-1:0] node75;
	wire [3-1:0] node77;
	wire [3-1:0] node78;
	wire [3-1:0] node80;
	wire [3-1:0] node84;
	wire [3-1:0] node85;
	wire [3-1:0] node86;
	wire [3-1:0] node87;
	wire [3-1:0] node89;
	wire [3-1:0] node90;
	wire [3-1:0] node92;
	wire [3-1:0] node94;
	wire [3-1:0] node96;
	wire [3-1:0] node100;
	wire [3-1:0] node101;
	wire [3-1:0] node102;
	wire [3-1:0] node107;
	wire [3-1:0] node108;
	wire [3-1:0] node109;
	wire [3-1:0] node111;
	wire [3-1:0] node113;
	wire [3-1:0] node117;
	wire [3-1:0] node119;
	wire [3-1:0] node122;
	wire [3-1:0] node123;
	wire [3-1:0] node124;
	wire [3-1:0] node125;
	wire [3-1:0] node126;
	wire [3-1:0] node128;
	wire [3-1:0] node130;
	wire [3-1:0] node134;
	wire [3-1:0] node136;
	wire [3-1:0] node137;
	wire [3-1:0] node141;
	wire [3-1:0] node142;
	wire [3-1:0] node144;
	wire [3-1:0] node146;
	wire [3-1:0] node149;
	wire [3-1:0] node152;
	wire [3-1:0] node153;
	wire [3-1:0] node154;
	wire [3-1:0] node156;
	wire [3-1:0] node158;
	wire [3-1:0] node160;
	wire [3-1:0] node163;
	wire [3-1:0] node165;
	wire [3-1:0] node167;
	wire [3-1:0] node170;
	wire [3-1:0] node171;
	wire [3-1:0] node172;
	wire [3-1:0] node174;
	wire [3-1:0] node176;
	wire [3-1:0] node179;
	wire [3-1:0] node180;
	wire [3-1:0] node184;
	wire [3-1:0] node185;
	wire [3-1:0] node187;
	wire [3-1:0] node190;
	wire [3-1:0] node192;
	wire [3-1:0] node194;

	assign outp = (inp[2]) ? node84 : node1;
		assign node1 = (inp[4]) ? node33 : node2;
			assign node2 = (inp[10]) ? node24 : node3;
				assign node3 = (inp[11]) ? node5 : 3'b111;
					assign node5 = (inp[5]) ? node7 : 3'b111;
						assign node7 = (inp[9]) ? node9 : 3'b111;
							assign node9 = (inp[7]) ? node17 : node10;
								assign node10 = (inp[6]) ? node12 : 3'b111;
									assign node12 = (inp[0]) ? 3'b111 : node13;
										assign node13 = (inp[8]) ? 3'b110 : 3'b111;
								assign node17 = (inp[3]) ? 3'b110 : node18;
									assign node18 = (inp[1]) ? 3'b111 : node19;
										assign node19 = (inp[6]) ? 3'b110 : 3'b111;
				assign node24 = (inp[5]) ? node26 : 3'b110;
					assign node26 = (inp[9]) ? node28 : 3'b110;
						assign node28 = (inp[3]) ? 3'b011 : node29;
							assign node29 = (inp[8]) ? 3'b111 : 3'b110;
			assign node33 = (inp[3]) ? node63 : node34;
				assign node34 = (inp[5]) ? node56 : node35;
					assign node35 = (inp[8]) ? node43 : node36;
						assign node36 = (inp[7]) ? 3'b110 : node37;
							assign node37 = (inp[9]) ? 3'b110 : node38;
								assign node38 = (inp[10]) ? 3'b111 : 3'b110;
						assign node43 = (inp[9]) ? node51 : node44;
							assign node44 = (inp[10]) ? node46 : 3'b110;
								assign node46 = (inp[7]) ? 3'b110 : node47;
									assign node47 = (inp[11]) ? 3'b110 : 3'b111;
							assign node51 = (inp[10]) ? 3'b110 : node52;
								assign node52 = (inp[7]) ? 3'b111 : 3'b110;
					assign node56 = (inp[9]) ? node60 : node57;
						assign node57 = (inp[10]) ? 3'b110 : 3'b111;
						assign node60 = (inp[10]) ? 3'b011 : 3'b111;
				assign node63 = (inp[5]) ? node75 : node64;
					assign node64 = (inp[10]) ? 3'b011 : node65;
						assign node65 = (inp[9]) ? node67 : 3'b011;
							assign node67 = (inp[7]) ? 3'b010 : node68;
								assign node68 = (inp[11]) ? node70 : 3'b011;
									assign node70 = (inp[8]) ? 3'b010 : 3'b011;
					assign node75 = (inp[8]) ? node77 : 3'b010;
						assign node77 = (inp[10]) ? 3'b010 : node78;
							assign node78 = (inp[9]) ? node80 : 3'b010;
								assign node80 = (inp[7]) ? 3'b011 : 3'b010;
		assign node84 = (inp[4]) ? node122 : node85;
			assign node85 = (inp[10]) ? node107 : node86;
				assign node86 = (inp[5]) ? node100 : node87;
					assign node87 = (inp[3]) ? node89 : 3'b011;
						assign node89 = (inp[9]) ? 3'b010 : node90;
							assign node90 = (inp[7]) ? node92 : 3'b011;
								assign node92 = (inp[6]) ? node94 : 3'b011;
									assign node94 = (inp[11]) ? node96 : 3'b011;
										assign node96 = (inp[8]) ? 3'b010 : 3'b011;
					assign node100 = (inp[3]) ? 3'b010 : node101;
						assign node101 = (inp[9]) ? 3'b010 : node102;
							assign node102 = (inp[7]) ? 3'b010 : 3'b011;
				assign node107 = (inp[3]) ? node117 : node108;
					assign node108 = (inp[5]) ? 3'b011 : node109;
						assign node109 = (inp[7]) ? node111 : 3'b010;
							assign node111 = (inp[9]) ? node113 : 3'b010;
								assign node113 = (inp[8]) ? 3'b011 : 3'b010;
					assign node117 = (inp[9]) ? node119 : 3'b111;
						assign node119 = (inp[5]) ? 3'b110 : 3'b111;
			assign node122 = (inp[3]) ? node152 : node123;
				assign node123 = (inp[5]) ? node141 : node124;
					assign node124 = (inp[10]) ? node134 : node125;
						assign node125 = (inp[0]) ? 3'b101 : node126;
							assign node126 = (inp[7]) ? node128 : 3'b101;
								assign node128 = (inp[9]) ? node130 : 3'b101;
									assign node130 = (inp[6]) ? 3'b100 : 3'b101;
						assign node134 = (inp[9]) ? node136 : 3'b101;
							assign node136 = (inp[7]) ? 3'b100 : node137;
								assign node137 = (inp[6]) ? 3'b100 : 3'b101;
					assign node141 = (inp[10]) ? node149 : node142;
						assign node142 = (inp[7]) ? node144 : 3'b100;
							assign node144 = (inp[8]) ? node146 : 3'b100;
								assign node146 = (inp[9]) ? 3'b101 : 3'b100;
						assign node149 = (inp[9]) ? 3'b001 : 3'b100;
				assign node152 = (inp[10]) ? node170 : node153;
					assign node153 = (inp[9]) ? node163 : node154;
						assign node154 = (inp[7]) ? node156 : 3'b001;
							assign node156 = (inp[5]) ? node158 : 3'b000;
								assign node158 = (inp[11]) ? node160 : 3'b001;
									assign node160 = (inp[8]) ? 3'b000 : 3'b001;
						assign node163 = (inp[8]) ? node165 : 3'b000;
							assign node165 = (inp[7]) ? node167 : 3'b000;
								assign node167 = (inp[5]) ? 3'b000 : 3'b001;
					assign node170 = (inp[9]) ? node184 : node171;
						assign node171 = (inp[7]) ? node179 : node172;
							assign node172 = (inp[8]) ? node174 : 3'b101;
								assign node174 = (inp[5]) ? node176 : 3'b101;
									assign node176 = (inp[6]) ? 3'b100 : 3'b101;
							assign node179 = (inp[5]) ? 3'b100 : node180;
								assign node180 = (inp[6]) ? 3'b100 : 3'b101;
						assign node184 = (inp[5]) ? node190 : node185;
							assign node185 = (inp[8]) ? node187 : 3'b100;
								assign node187 = (inp[7]) ? 3'b101 : 3'b100;
							assign node190 = (inp[7]) ? node192 : 3'b001;
								assign node192 = (inp[8]) ? node194 : 3'b000;
									assign node194 = (inp[6]) ? 3'b000 : 3'b001;

endmodule