module dtc_split125_bm96 (
	input  wire [12-1:0] inp,
	output wire [3-1:0] outp
);

	wire [3-1:0] node1;
	wire [3-1:0] node2;
	wire [3-1:0] node4;
	wire [3-1:0] node5;
	wire [3-1:0] node7;
	wire [3-1:0] node9;
	wire [3-1:0] node14;
	wire [3-1:0] node16;
	wire [3-1:0] node17;
	wire [3-1:0] node18;
	wire [3-1:0] node19;
	wire [3-1:0] node21;
	wire [3-1:0] node22;
	wire [3-1:0] node27;
	wire [3-1:0] node28;
	wire [3-1:0] node29;
	wire [3-1:0] node30;
	wire [3-1:0] node31;
	wire [3-1:0] node34;
	wire [3-1:0] node37;
	wire [3-1:0] node38;
	wire [3-1:0] node43;
	wire [3-1:0] node44;
	wire [3-1:0] node46;
	wire [3-1:0] node49;
	wire [3-1:0] node50;
	wire [3-1:0] node51;
	wire [3-1:0] node55;
	wire [3-1:0] node56;
	wire [3-1:0] node60;
	wire [3-1:0] node61;
	wire [3-1:0] node62;
	wire [3-1:0] node63;
	wire [3-1:0] node64;
	wire [3-1:0] node65;
	wire [3-1:0] node70;
	wire [3-1:0] node71;
	wire [3-1:0] node74;
	wire [3-1:0] node77;
	wire [3-1:0] node78;
	wire [3-1:0] node81;
	wire [3-1:0] node83;
	wire [3-1:0] node86;
	wire [3-1:0] node87;
	wire [3-1:0] node88;
	wire [3-1:0] node89;
	wire [3-1:0] node93;
	wire [3-1:0] node95;
	wire [3-1:0] node96;
	wire [3-1:0] node100;
	wire [3-1:0] node101;
	wire [3-1:0] node104;
	wire [3-1:0] node105;
	wire [3-1:0] node107;

	assign outp = (inp[7]) ? node14 : node1;
		assign node1 = (inp[10]) ? 3'b000 : node2;
			assign node2 = (inp[2]) ? node4 : 3'b000;
				assign node4 = (inp[11]) ? 3'b000 : node5;
					assign node5 = (inp[4]) ? node7 : 3'b000;
						assign node7 = (inp[3]) ? node9 : 3'b000;
							assign node9 = (inp[8]) ? 3'b100 : 3'b000;
		assign node14 = (inp[6]) ? node16 : 3'b000;
			assign node16 = (inp[3]) ? node60 : node17;
				assign node17 = (inp[4]) ? node27 : node18;
					assign node18 = (inp[1]) ? 3'b011 : node19;
						assign node19 = (inp[9]) ? node21 : 3'b011;
							assign node21 = (inp[10]) ? 3'b101 : node22;
								assign node22 = (inp[5]) ? 3'b011 : 3'b111;
					assign node27 = (inp[0]) ? node43 : node28;
						assign node28 = (inp[1]) ? 3'b010 : node29;
							assign node29 = (inp[11]) ? node37 : node30;
								assign node30 = (inp[5]) ? node34 : node31;
									assign node31 = (inp[10]) ? 3'b001 : 3'b010;
									assign node34 = (inp[2]) ? 3'b001 : 3'b000;
								assign node37 = (inp[5]) ? 3'b010 : node38;
									assign node38 = (inp[9]) ? 3'b001 : 3'b010;
						assign node43 = (inp[9]) ? node49 : node44;
							assign node44 = (inp[2]) ? node46 : 3'b001;
								assign node46 = (inp[10]) ? 3'b010 : 3'b001;
							assign node49 = (inp[2]) ? node55 : node50;
								assign node50 = (inp[10]) ? 3'b010 : node51;
									assign node51 = (inp[11]) ? 3'b101 : 3'b110;
								assign node55 = (inp[10]) ? 3'b001 : node56;
									assign node56 = (inp[8]) ? 3'b101 : 3'b001;
				assign node60 = (inp[1]) ? node86 : node61;
					assign node61 = (inp[0]) ? node77 : node62;
						assign node62 = (inp[5]) ? node70 : node63;
							assign node63 = (inp[4]) ? 3'b110 : node64;
								assign node64 = (inp[11]) ? 3'b111 : node65;
									assign node65 = (inp[2]) ? 3'b110 : 3'b111;
							assign node70 = (inp[9]) ? node74 : node71;
								assign node71 = (inp[10]) ? 3'b001 : 3'b011;
								assign node74 = (inp[4]) ? 3'b010 : 3'b011;
						assign node77 = (inp[11]) ? node81 : node78;
							assign node78 = (inp[4]) ? 3'b110 : 3'b111;
							assign node81 = (inp[9]) ? node83 : 3'b110;
								assign node83 = (inp[4]) ? 3'b100 : 3'b110;
					assign node86 = (inp[4]) ? node100 : node87;
						assign node87 = (inp[11]) ? node93 : node88;
							assign node88 = (inp[0]) ? 3'b101 : node89;
								assign node89 = (inp[9]) ? 3'b101 : 3'b100;
							assign node93 = (inp[9]) ? node95 : 3'b100;
								assign node95 = (inp[0]) ? 3'b100 : node96;
									assign node96 = (inp[5]) ? 3'b100 : 3'b101;
						assign node100 = (inp[0]) ? node104 : node101;
							assign node101 = (inp[9]) ? 3'b010 : 3'b001;
							assign node104 = (inp[9]) ? 3'b000 : node105;
								assign node105 = (inp[8]) ? node107 : 3'b100;
									assign node107 = (inp[10]) ? 3'b010 : 3'b110;

endmodule