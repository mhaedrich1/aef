module dtc_split25_bm45 (
	input  wire [16-1:0] inp,
	output wire [46-1:0] outp
);

	wire [46-1:0] node1;
	wire [46-1:0] node2;
	wire [46-1:0] node4;
	wire [46-1:0] node6;
	wire [46-1:0] node8;
	wire [46-1:0] node10;
	wire [46-1:0] node12;
	wire [46-1:0] node14;
	wire [46-1:0] node15;
	wire [46-1:0] node16;
	wire [46-1:0] node18;
	wire [46-1:0] node19;
	wire [46-1:0] node24;
	wire [46-1:0] node26;
	wire [46-1:0] node27;
	wire [46-1:0] node29;
	wire [46-1:0] node31;
	wire [46-1:0] node35;
	wire [46-1:0] node37;
	wire [46-1:0] node38;
	wire [46-1:0] node39;
	wire [46-1:0] node40;
	wire [46-1:0] node41;
	wire [46-1:0] node45;
	wire [46-1:0] node47;
	wire [46-1:0] node49;
	wire [46-1:0] node50;
	wire [46-1:0] node52;
	wire [46-1:0] node53;
	wire [46-1:0] node55;
	wire [46-1:0] node56;
	wire [46-1:0] node58;
	wire [46-1:0] node64;
	wire [46-1:0] node65;
	wire [46-1:0] node66;
	wire [46-1:0] node70;
	wire [46-1:0] node71;
	wire [46-1:0] node74;
	wire [46-1:0] node77;
	wire [46-1:0] node78;
	wire [46-1:0] node79;
	wire [46-1:0] node80;
	wire [46-1:0] node83;
	wire [46-1:0] node85;
	wire [46-1:0] node87;
	wire [46-1:0] node89;
	wire [46-1:0] node90;
	wire [46-1:0] node93;
	wire [46-1:0] node94;
	wire [46-1:0] node95;
	wire [46-1:0] node99;
	wire [46-1:0] node100;
	wire [46-1:0] node101;
	wire [46-1:0] node106;
	wire [46-1:0] node107;
	wire [46-1:0] node109;
	wire [46-1:0] node110;
	wire [46-1:0] node112;
	wire [46-1:0] node113;
	wire [46-1:0] node115;
	wire [46-1:0] node120;
	wire [46-1:0] node122;
	wire [46-1:0] node124;
	wire [46-1:0] node126;
	wire [46-1:0] node127;
	wire [46-1:0] node129;
	wire [46-1:0] node131;
	wire [46-1:0] node133;
	wire [46-1:0] node137;
	wire [46-1:0] node139;
	wire [46-1:0] node140;
	wire [46-1:0] node142;
	wire [46-1:0] node144;
	wire [46-1:0] node146;
	wire [46-1:0] node148;
	wire [46-1:0] node149;
	wire [46-1:0] node151;
	wire [46-1:0] node155;
	wire [46-1:0] node157;
	wire [46-1:0] node159;
	wire [46-1:0] node160;
	wire [46-1:0] node161;
	wire [46-1:0] node162;
	wire [46-1:0] node164;
	wire [46-1:0] node166;
	wire [46-1:0] node170;
	wire [46-1:0] node171;
	wire [46-1:0] node172;
	wire [46-1:0] node173;
	wire [46-1:0] node178;
	wire [46-1:0] node179;
	wire [46-1:0] node180;
	wire [46-1:0] node183;
	wire [46-1:0] node187;
	wire [46-1:0] node188;
	wire [46-1:0] node189;
	wire [46-1:0] node194;
	wire [46-1:0] node195;
	wire [46-1:0] node196;
	wire [46-1:0] node199;
	wire [46-1:0] node200;
	wire [46-1:0] node201;
	wire [46-1:0] node202;
	wire [46-1:0] node203;
	wire [46-1:0] node206;
	wire [46-1:0] node209;
	wire [46-1:0] node210;
	wire [46-1:0] node213;
	wire [46-1:0] node216;
	wire [46-1:0] node217;
	wire [46-1:0] node218;
	wire [46-1:0] node221;
	wire [46-1:0] node224;
	wire [46-1:0] node225;
	wire [46-1:0] node228;
	wire [46-1:0] node231;
	wire [46-1:0] node232;
	wire [46-1:0] node233;
	wire [46-1:0] node234;
	wire [46-1:0] node237;
	wire [46-1:0] node240;
	wire [46-1:0] node241;
	wire [46-1:0] node244;
	wire [46-1:0] node247;
	wire [46-1:0] node248;
	wire [46-1:0] node249;
	wire [46-1:0] node252;
	wire [46-1:0] node255;
	wire [46-1:0] node256;
	wire [46-1:0] node259;
	wire [46-1:0] node262;
	wire [46-1:0] node263;
	wire [46-1:0] node266;
	wire [46-1:0] node268;
	wire [46-1:0] node269;
	wire [46-1:0] node270;
	wire [46-1:0] node271;
	wire [46-1:0] node272;
	wire [46-1:0] node273;
	wire [46-1:0] node274;
	wire [46-1:0] node275;
	wire [46-1:0] node276;
	wire [46-1:0] node277;
	wire [46-1:0] node280;
	wire [46-1:0] node283;
	wire [46-1:0] node284;
	wire [46-1:0] node288;
	wire [46-1:0] node289;
	wire [46-1:0] node290;
	wire [46-1:0] node293;
	wire [46-1:0] node296;
	wire [46-1:0] node297;
	wire [46-1:0] node299;
	wire [46-1:0] node302;
	wire [46-1:0] node305;
	wire [46-1:0] node306;
	wire [46-1:0] node307;
	wire [46-1:0] node308;
	wire [46-1:0] node311;
	wire [46-1:0] node314;
	wire [46-1:0] node317;
	wire [46-1:0] node318;
	wire [46-1:0] node321;
	wire [46-1:0] node322;
	wire [46-1:0] node324;
	wire [46-1:0] node328;
	wire [46-1:0] node329;
	wire [46-1:0] node330;
	wire [46-1:0] node331;
	wire [46-1:0] node333;
	wire [46-1:0] node334;
	wire [46-1:0] node338;
	wire [46-1:0] node339;
	wire [46-1:0] node341;
	wire [46-1:0] node344;
	wire [46-1:0] node346;
	wire [46-1:0] node349;
	wire [46-1:0] node350;
	wire [46-1:0] node352;
	wire [46-1:0] node356;
	wire [46-1:0] node357;
	wire [46-1:0] node358;
	wire [46-1:0] node359;
	wire [46-1:0] node361;
	wire [46-1:0] node364;
	wire [46-1:0] node367;
	wire [46-1:0] node370;
	wire [46-1:0] node371;
	wire [46-1:0] node373;
	wire [46-1:0] node374;
	wire [46-1:0] node377;
	wire [46-1:0] node381;
	wire [46-1:0] node382;
	wire [46-1:0] node383;
	wire [46-1:0] node384;
	wire [46-1:0] node385;
	wire [46-1:0] node386;
	wire [46-1:0] node387;
	wire [46-1:0] node391;
	wire [46-1:0] node393;
	wire [46-1:0] node396;
	wire [46-1:0] node397;
	wire [46-1:0] node398;
	wire [46-1:0] node402;
	wire [46-1:0] node403;
	wire [46-1:0] node407;
	wire [46-1:0] node408;
	wire [46-1:0] node409;
	wire [46-1:0] node413;
	wire [46-1:0] node415;
	wire [46-1:0] node418;
	wire [46-1:0] node419;
	wire [46-1:0] node420;
	wire [46-1:0] node421;
	wire [46-1:0] node426;
	wire [46-1:0] node427;
	wire [46-1:0] node428;
	wire [46-1:0] node429;
	wire [46-1:0] node433;
	wire [46-1:0] node434;
	wire [46-1:0] node438;
	wire [46-1:0] node439;
	wire [46-1:0] node442;
	wire [46-1:0] node445;
	wire [46-1:0] node446;
	wire [46-1:0] node447;
	wire [46-1:0] node448;
	wire [46-1:0] node449;
	wire [46-1:0] node450;
	wire [46-1:0] node454;
	wire [46-1:0] node455;
	wire [46-1:0] node458;
	wire [46-1:0] node461;
	wire [46-1:0] node463;
	wire [46-1:0] node466;
	wire [46-1:0] node467;
	wire [46-1:0] node469;
	wire [46-1:0] node472;
	wire [46-1:0] node475;
	wire [46-1:0] node476;
	wire [46-1:0] node477;
	wire [46-1:0] node478;
	wire [46-1:0] node480;
	wire [46-1:0] node483;
	wire [46-1:0] node486;
	wire [46-1:0] node487;
	wire [46-1:0] node490;
	wire [46-1:0] node493;
	wire [46-1:0] node494;
	wire [46-1:0] node495;
	wire [46-1:0] node498;
	wire [46-1:0] node501;
	wire [46-1:0] node502;
	wire [46-1:0] node503;
	wire [46-1:0] node507;
	wire [46-1:0] node510;
	wire [46-1:0] node511;
	wire [46-1:0] node513;
	wire [46-1:0] node515;
	wire [46-1:0] node516;
	wire [46-1:0] node518;
	wire [46-1:0] node519;
	wire [46-1:0] node523;
	wire [46-1:0] node524;
	wire [46-1:0] node526;
	wire [46-1:0] node529;
	wire [46-1:0] node530;
	wire [46-1:0] node533;
	wire [46-1:0] node536;
	wire [46-1:0] node537;
	wire [46-1:0] node538;
	wire [46-1:0] node539;
	wire [46-1:0] node540;
	wire [46-1:0] node541;
	wire [46-1:0] node542;
	wire [46-1:0] node546;
	wire [46-1:0] node549;
	wire [46-1:0] node550;
	wire [46-1:0] node552;
	wire [46-1:0] node555;
	wire [46-1:0] node558;
	wire [46-1:0] node559;
	wire [46-1:0] node560;
	wire [46-1:0] node563;
	wire [46-1:0] node566;
	wire [46-1:0] node569;
	wire [46-1:0] node570;
	wire [46-1:0] node571;
	wire [46-1:0] node572;
	wire [46-1:0] node575;
	wire [46-1:0] node578;
	wire [46-1:0] node579;
	wire [46-1:0] node583;
	wire [46-1:0] node584;
	wire [46-1:0] node585;
	wire [46-1:0] node588;
	wire [46-1:0] node591;
	wire [46-1:0] node592;
	wire [46-1:0] node595;
	wire [46-1:0] node596;
	wire [46-1:0] node600;
	wire [46-1:0] node601;
	wire [46-1:0] node602;
	wire [46-1:0] node603;
	wire [46-1:0] node604;
	wire [46-1:0] node608;
	wire [46-1:0] node609;
	wire [46-1:0] node610;
	wire [46-1:0] node613;
	wire [46-1:0] node616;
	wire [46-1:0] node619;
	wire [46-1:0] node620;
	wire [46-1:0] node621;
	wire [46-1:0] node625;
	wire [46-1:0] node626;
	wire [46-1:0] node627;
	wire [46-1:0] node631;
	wire [46-1:0] node633;
	wire [46-1:0] node636;
	wire [46-1:0] node637;
	wire [46-1:0] node638;
	wire [46-1:0] node641;
	wire [46-1:0] node642;
	wire [46-1:0] node645;
	wire [46-1:0] node646;
	wire [46-1:0] node650;
	wire [46-1:0] node651;
	wire [46-1:0] node652;
	wire [46-1:0] node654;
	wire [46-1:0] node658;
	wire [46-1:0] node661;
	wire [46-1:0] node662;
	wire [46-1:0] node663;
	wire [46-1:0] node664;
	wire [46-1:0] node666;
	wire [46-1:0] node667;
	wire [46-1:0] node668;
	wire [46-1:0] node669;
	wire [46-1:0] node671;
	wire [46-1:0] node675;
	wire [46-1:0] node677;
	wire [46-1:0] node680;
	wire [46-1:0] node682;
	wire [46-1:0] node683;
	wire [46-1:0] node687;
	wire [46-1:0] node688;
	wire [46-1:0] node689;
	wire [46-1:0] node692;
	wire [46-1:0] node693;
	wire [46-1:0] node696;
	wire [46-1:0] node701;
	wire [46-1:0] node702;
	wire [46-1:0] node703;
	wire [46-1:0] node704;
	wire [46-1:0] node705;
	wire [46-1:0] node706;
	wire [46-1:0] node708;
	wire [46-1:0] node711;
	wire [46-1:0] node713;
	wire [46-1:0] node716;
	wire [46-1:0] node717;
	wire [46-1:0] node720;
	wire [46-1:0] node721;
	wire [46-1:0] node724;
	wire [46-1:0] node727;
	wire [46-1:0] node728;
	wire [46-1:0] node729;
	wire [46-1:0] node731;
	wire [46-1:0] node734;
	wire [46-1:0] node736;
	wire [46-1:0] node737;
	wire [46-1:0] node741;
	wire [46-1:0] node742;
	wire [46-1:0] node744;
	wire [46-1:0] node747;
	wire [46-1:0] node748;
	wire [46-1:0] node749;
	wire [46-1:0] node752;
	wire [46-1:0] node755;
	wire [46-1:0] node758;
	wire [46-1:0] node759;
	wire [46-1:0] node760;
	wire [46-1:0] node761;
	wire [46-1:0] node763;
	wire [46-1:0] node766;
	wire [46-1:0] node767;
	wire [46-1:0] node768;
	wire [46-1:0] node771;
	wire [46-1:0] node774;
	wire [46-1:0] node775;
	wire [46-1:0] node779;
	wire [46-1:0] node782;
	wire [46-1:0] node783;
	wire [46-1:0] node784;
	wire [46-1:0] node786;
	wire [46-1:0] node789;
	wire [46-1:0] node791;
	wire [46-1:0] node794;
	wire [46-1:0] node797;
	wire [46-1:0] node798;
	wire [46-1:0] node799;
	wire [46-1:0] node800;
	wire [46-1:0] node801;
	wire [46-1:0] node804;
	wire [46-1:0] node805;
	wire [46-1:0] node806;
	wire [46-1:0] node810;
	wire [46-1:0] node812;
	wire [46-1:0] node815;
	wire [46-1:0] node816;
	wire [46-1:0] node818;
	wire [46-1:0] node819;
	wire [46-1:0] node824;
	wire [46-1:0] node825;
	wire [46-1:0] node826;
	wire [46-1:0] node827;
	wire [46-1:0] node830;
	wire [46-1:0] node833;
	wire [46-1:0] node834;
	wire [46-1:0] node838;
	wire [46-1:0] node839;
	wire [46-1:0] node842;
	wire [46-1:0] node843;
	wire [46-1:0] node845;
	wire [46-1:0] node848;
	wire [46-1:0] node850;
	wire [46-1:0] node853;
	wire [46-1:0] node854;
	wire [46-1:0] node855;
	wire [46-1:0] node856;
	wire [46-1:0] node857;
	wire [46-1:0] node859;
	wire [46-1:0] node862;
	wire [46-1:0] node865;
	wire [46-1:0] node866;
	wire [46-1:0] node867;
	wire [46-1:0] node872;
	wire [46-1:0] node873;
	wire [46-1:0] node874;
	wire [46-1:0] node877;
	wire [46-1:0] node880;
	wire [46-1:0] node881;
	wire [46-1:0] node884;
	wire [46-1:0] node887;
	wire [46-1:0] node888;
	wire [46-1:0] node889;
	wire [46-1:0] node891;
	wire [46-1:0] node893;
	wire [46-1:0] node896;
	wire [46-1:0] node897;
	wire [46-1:0] node898;
	wire [46-1:0] node903;
	wire [46-1:0] node906;
	wire [46-1:0] node907;
	wire [46-1:0] node908;
	wire [46-1:0] node909;
	wire [46-1:0] node911;
	wire [46-1:0] node913;
	wire [46-1:0] node915;
	wire [46-1:0] node917;
	wire [46-1:0] node919;
	wire [46-1:0] node922;
	wire [46-1:0] node923;
	wire [46-1:0] node925;
	wire [46-1:0] node927;
	wire [46-1:0] node929;
	wire [46-1:0] node930;
	wire [46-1:0] node933;
	wire [46-1:0] node935;
	wire [46-1:0] node938;
	wire [46-1:0] node939;
	wire [46-1:0] node940;
	wire [46-1:0] node941;
	wire [46-1:0] node944;
	wire [46-1:0] node945;
	wire [46-1:0] node948;
	wire [46-1:0] node951;
	wire [46-1:0] node952;
	wire [46-1:0] node953;
	wire [46-1:0] node956;
	wire [46-1:0] node958;
	wire [46-1:0] node961;
	wire [46-1:0] node962;
	wire [46-1:0] node964;
	wire [46-1:0] node968;
	wire [46-1:0] node969;
	wire [46-1:0] node971;
	wire [46-1:0] node972;
	wire [46-1:0] node976;
	wire [46-1:0] node977;
	wire [46-1:0] node978;
	wire [46-1:0] node980;
	wire [46-1:0] node983;
	wire [46-1:0] node987;
	wire [46-1:0] node988;
	wire [46-1:0] node989;
	wire [46-1:0] node990;
	wire [46-1:0] node991;
	wire [46-1:0] node992;
	wire [46-1:0] node993;
	wire [46-1:0] node996;
	wire [46-1:0] node998;
	wire [46-1:0] node1001;
	wire [46-1:0] node1003;
	wire [46-1:0] node1006;
	wire [46-1:0] node1007;
	wire [46-1:0] node1008;
	wire [46-1:0] node1011;
	wire [46-1:0] node1014;
	wire [46-1:0] node1016;
	wire [46-1:0] node1018;
	wire [46-1:0] node1021;
	wire [46-1:0] node1022;
	wire [46-1:0] node1024;
	wire [46-1:0] node1027;
	wire [46-1:0] node1028;
	wire [46-1:0] node1031;
	wire [46-1:0] node1032;
	wire [46-1:0] node1034;
	wire [46-1:0] node1037;
	wire [46-1:0] node1040;
	wire [46-1:0] node1041;
	wire [46-1:0] node1042;
	wire [46-1:0] node1043;
	wire [46-1:0] node1044;
	wire [46-1:0] node1045;
	wire [46-1:0] node1049;
	wire [46-1:0] node1050;
	wire [46-1:0] node1054;
	wire [46-1:0] node1055;
	wire [46-1:0] node1059;
	wire [46-1:0] node1060;
	wire [46-1:0] node1063;
	wire [46-1:0] node1064;
	wire [46-1:0] node1067;
	wire [46-1:0] node1070;
	wire [46-1:0] node1071;
	wire [46-1:0] node1072;
	wire [46-1:0] node1074;
	wire [46-1:0] node1077;
	wire [46-1:0] node1078;
	wire [46-1:0] node1081;
	wire [46-1:0] node1082;
	wire [46-1:0] node1085;
	wire [46-1:0] node1088;
	wire [46-1:0] node1089;
	wire [46-1:0] node1090;
	wire [46-1:0] node1091;
	wire [46-1:0] node1095;
	wire [46-1:0] node1098;
	wire [46-1:0] node1099;
	wire [46-1:0] node1102;
	wire [46-1:0] node1105;
	wire [46-1:0] node1106;
	wire [46-1:0] node1107;
	wire [46-1:0] node1108;
	wire [46-1:0] node1109;
	wire [46-1:0] node1110;
	wire [46-1:0] node1112;
	wire [46-1:0] node1116;
	wire [46-1:0] node1119;
	wire [46-1:0] node1120;
	wire [46-1:0] node1121;
	wire [46-1:0] node1124;
	wire [46-1:0] node1128;
	wire [46-1:0] node1129;
	wire [46-1:0] node1130;
	wire [46-1:0] node1131;
	wire [46-1:0] node1134;
	wire [46-1:0] node1137;
	wire [46-1:0] node1138;
	wire [46-1:0] node1139;
	wire [46-1:0] node1143;
	wire [46-1:0] node1146;
	wire [46-1:0] node1147;
	wire [46-1:0] node1149;
	wire [46-1:0] node1152;
	wire [46-1:0] node1153;
	wire [46-1:0] node1156;
	wire [46-1:0] node1157;
	wire [46-1:0] node1161;
	wire [46-1:0] node1162;
	wire [46-1:0] node1163;
	wire [46-1:0] node1164;
	wire [46-1:0] node1166;
	wire [46-1:0] node1170;
	wire [46-1:0] node1171;
	wire [46-1:0] node1172;
	wire [46-1:0] node1175;
	wire [46-1:0] node1177;
	wire [46-1:0] node1180;
	wire [46-1:0] node1181;
	wire [46-1:0] node1185;
	wire [46-1:0] node1186;
	wire [46-1:0] node1187;
	wire [46-1:0] node1188;
	wire [46-1:0] node1191;
	wire [46-1:0] node1194;
	wire [46-1:0] node1195;
	wire [46-1:0] node1199;
	wire [46-1:0] node1200;
	wire [46-1:0] node1201;
	wire [46-1:0] node1202;
	wire [46-1:0] node1206;
	wire [46-1:0] node1209;
	wire [46-1:0] node1210;
	wire [46-1:0] node1213;
	wire [46-1:0] node1215;
	wire [46-1:0] node1218;
	wire [46-1:0] node1219;
	wire [46-1:0] node1220;
	wire [46-1:0] node1221;
	wire [46-1:0] node1223;
	wire [46-1:0] node1224;
	wire [46-1:0] node1227;
	wire [46-1:0] node1230;
	wire [46-1:0] node1231;
	wire [46-1:0] node1232;
	wire [46-1:0] node1235;
	wire [46-1:0] node1239;
	wire [46-1:0] node1240;
	wire [46-1:0] node1242;
	wire [46-1:0] node1243;
	wire [46-1:0] node1246;
	wire [46-1:0] node1249;
	wire [46-1:0] node1250;
	wire [46-1:0] node1251;
	wire [46-1:0] node1254;
	wire [46-1:0] node1258;
	wire [46-1:0] node1259;
	wire [46-1:0] node1260;
	wire [46-1:0] node1262;
	wire [46-1:0] node1263;
	wire [46-1:0] node1266;
	wire [46-1:0] node1269;
	wire [46-1:0] node1270;
	wire [46-1:0] node1271;
	wire [46-1:0] node1274;

	assign outp = (inp[1]) ? node194 : node1;
		assign node1 = (inp[15]) ? node35 : node2;
			assign node2 = (inp[7]) ? node4 : 46'b0000000000000000000000000000000000000000000000;
				assign node4 = (inp[8]) ? node6 : 46'b0000000000000000000000000000000000000000000000;
					assign node6 = (inp[3]) ? node8 : 46'b0000000000000000000000000000000000000000000000;
						assign node8 = (inp[6]) ? node10 : 46'b0000000000000000000000000000000000000000000000;
							assign node10 = (inp[12]) ? node12 : 46'b0000000000000000000000000000000000000000000000;
								assign node12 = (inp[5]) ? node14 : 46'b0000000000000000000000000000000000000000000000;
									assign node14 = (inp[4]) ? node24 : node15;
										assign node15 = (inp[9]) ? 46'b0000000000000000000000000000000000000000000000 : node16;
											assign node16 = (inp[13]) ? node18 : 46'b0000000000000000000000000000000000000000000000;
												assign node18 = (inp[11]) ? 46'b0000000000000000000000000000000000000000000000 : node19;
													assign node19 = (inp[0]) ? 46'b0000000000000000000000000000000000000000000000 : 46'b0000000000000000000000000000000000000100000000;
										assign node24 = (inp[14]) ? node26 : 46'b0000000000000000000000000000000000000000000000;
											assign node26 = (inp[11]) ? 46'b0000000000000000000000000000000000000000000000 : node27;
												assign node27 = (inp[13]) ? node29 : 46'b0000000000000000000000000000000000000000000000;
													assign node29 = (inp[10]) ? node31 : 46'b0000000000000000000000000000000000000000000000;
														assign node31 = (inp[0]) ? 46'b0000000001000000000000000000001000000000000000 : 46'b0000000000000000000000000000000000000000000000;
			assign node35 = (inp[3]) ? node37 : 46'b0000000000000000000000000000001000000000000000;
				assign node37 = (inp[9]) ? node77 : node38;
					assign node38 = (inp[11]) ? node64 : node39;
						assign node39 = (inp[13]) ? node45 : node40;
							assign node40 = (inp[2]) ? 46'b0000000000000000000000000000000000000000000000 : node41;
								assign node41 = (inp[0]) ? 46'b0000000000001000000000000010000000000000000000 : 46'b0000001000001000000000000000000000000000000000;
							assign node45 = (inp[14]) ? node47 : 46'b0000000000000000000000000000000000000000000000;
								assign node47 = (inp[8]) ? node49 : 46'b0000000000000000000000000000000000000000000000;
									assign node49 = (inp[7]) ? 46'b0000000000000000000000000000000000000000000000 : node50;
										assign node50 = (inp[5]) ? node52 : 46'b0000000000000000000000000000000000000000000000;
											assign node52 = (inp[0]) ? 46'b0000000000000000000000000000000000000000000000 : node53;
												assign node53 = (inp[12]) ? node55 : 46'b0000000000000000000000000000000000000000000000;
													assign node55 = (inp[2]) ? 46'b0000010000000000010000010000000001000010000000 : node56;
														assign node56 = (inp[6]) ? node58 : 46'b0000000000000000000000000000000000000000000000;
															assign node58 = (inp[10]) ? 46'b0000000000000000000000000000000000000000000000 : 46'b0000010000000000010100000000000100000000010000;
						assign node64 = (inp[13]) ? node70 : node65;
							assign node65 = (inp[2]) ? 46'b0000000000000000000000000000000000000000000000 : node66;
								assign node66 = (inp[0]) ? 46'b0000010000000000000000000010000000000000000000 : 46'b0000011000000000000000000000000000000000000000;
							assign node70 = (inp[2]) ? node74 : node71;
								assign node71 = (inp[0]) ? 46'b0000001000000000011000000100000000000000010000 : 46'b0000001000000000010000000100000000000000010010;
								assign node74 = (inp[0]) ? 46'b0000001000000000010010000000010000000010000000 : 46'b0000001000000000010010100000000000000010000000;
					assign node77 = (inp[2]) ? node137 : node78;
						assign node78 = (inp[0]) ? node106 : node79;
							assign node79 = (inp[13]) ? node83 : node80;
								assign node80 = (inp[11]) ? 46'b0000010100000000000000000000000000000000000000 : 46'b0000000100001000000000000000000000000000000000;
								assign node83 = (inp[5]) ? node85 : 46'b0000000000000000000000000000000000000000000000;
									assign node85 = (inp[14]) ? node87 : 46'b0000000000000000000000000000000000000000000000;
										assign node87 = (inp[4]) ? node89 : 46'b0000000000000000000000000000000000000000000000;
											assign node89 = (inp[6]) ? node93 : node90;
												assign node90 = (inp[11]) ? 46'b0000000000000000000000000100000000000000000010 : 46'b0000000000000000000000000000000000000000000000;
												assign node93 = (inp[8]) ? node99 : node94;
													assign node94 = (inp[7]) ? 46'b0000000000011000010000000100000000000000010010 : node95;
														assign node95 = (inp[11]) ? 46'b0000000000000000000000000000000000000000000000 : 46'b0000010000010000010000000000000000000000010000;
													assign node99 = (inp[10]) ? 46'b0000000000000000000000000000000000000000000000 : node100;
														assign node100 = (inp[7]) ? 46'b0000000000001000010000000000000100000000010000 : node101;
															assign node101 = (inp[11]) ? 46'b0010000000000000000000000100000100000000010010 : 46'b0010000000000000000000000000000100000000010000;
							assign node106 = (inp[11]) ? node120 : node107;
								assign node107 = (inp[13]) ? node109 : 46'b0010001000000000000000000000000000000000010000;
									assign node109 = (inp[7]) ? 46'b0000000000000000000000000000000000000000000000 : node110;
										assign node110 = (inp[14]) ? node112 : 46'b0000000000000000000000000000000000000000000000;
											assign node112 = (inp[8]) ? 46'b0000000000000000000000000000000000000000000000 : node113;
												assign node113 = (inp[10]) ? node115 : 46'b0000000000000000000000000000000000000000000000;
													assign node115 = (inp[4]) ? 46'b0010000000010000000000000000000000000000010100 : 46'b0000000000000000000000000000000000000000000000;
								assign node120 = (inp[8]) ? node122 : 46'b0000000000000000000000000000000000000000000000;
									assign node122 = (inp[13]) ? node124 : 46'b0000000000000000000000000000000000000000000000;
										assign node124 = (inp[5]) ? node126 : 46'b0000000000000000000000000000000000000000000000;
											assign node126 = (inp[6]) ? 46'b0000000000000000000000000000000000000000000000 : node127;
												assign node127 = (inp[10]) ? node129 : 46'b0000000000000000000000000000000000000000000000;
													assign node129 = (inp[14]) ? node131 : 46'b0000000000000000000000000000000000000000000000;
														assign node131 = (inp[7]) ? node133 : 46'b0000000000000000001000000100000001000000000000;
															assign node133 = (inp[12]) ? 46'b0000000000000000000000000000000000000000000000 : 46'b0000000000000000001000000100000000000000000000;
						assign node137 = (inp[13]) ? node139 : 46'b0000000000000000000000000000000000000000000000;
							assign node139 = (inp[6]) ? node155 : node140;
								assign node140 = (inp[0]) ? node142 : 46'b0000000000000000000000000000000000000000000000;
									assign node142 = (inp[10]) ? node144 : 46'b0000000000000000000000000000000000000000000000;
										assign node144 = (inp[5]) ? node146 : 46'b0000000000000000000000000000000000000000000000;
											assign node146 = (inp[8]) ? node148 : 46'b0000000000000000000000000000000000000000000000;
												assign node148 = (inp[12]) ? 46'b0000000000000000000000000000000000000000000000 : node149;
													assign node149 = (inp[11]) ? node151 : 46'b0000000000000000000000000000000000000000000000;
														assign node151 = (inp[7]) ? 46'b0000000000000000000010000000010000000000000000 : 46'b0000000000000000000000000000000000000000000000;
								assign node155 = (inp[14]) ? node157 : 46'b0000000000000000000000000000000000000000000000;
									assign node157 = (inp[5]) ? node159 : 46'b0000000000000000000000000000000000000000000000;
										assign node159 = (inp[0]) ? node187 : node160;
											assign node160 = (inp[11]) ? node170 : node161;
												assign node161 = (inp[8]) ? 46'b0000000000000000000000000000000000000000000000 : node162;
													assign node162 = (inp[7]) ? node164 : 46'b0000010000010000010000000000000000000010000000;
														assign node164 = (inp[4]) ? node166 : 46'b0000000000000000000000000000000000000000000000;
															assign node166 = (inp[10]) ? 46'b0000000000011000010000000000000000000010000000 : 46'b0000000000000000000000000000000000000000000000;
												assign node170 = (inp[10]) ? node178 : node171;
													assign node171 = (inp[7]) ? 46'b0000000000000000000000000000000000000000000000 : node172;
														assign node172 = (inp[12]) ? 46'b0000010000000000010010100000000100000010000000 : node173;
															assign node173 = (inp[8]) ? 46'b0000000000000000000000000000000000000000000000 : 46'b0000000000000000000000000000000000000000000000;
													assign node178 = (inp[12]) ? 46'b0000000000000000000000000000000000000000000000 : node179;
														assign node179 = (inp[7]) ? node183 : node180;
															assign node180 = (inp[4]) ? 46'b0010000000010000000010100000000000000010000000 : 46'b0010000000000000000010110000000000000010000000;
															assign node183 = (inp[8]) ? 46'b0000000000001000010010110000000000000010000000 : 46'b0000000000011000010010100000000000000010000000;
											assign node187 = (inp[10]) ? 46'b0000000000000000000000000000000000000000000000 : node188;
												assign node188 = (inp[7]) ? 46'b0000000000000000000000000000000000000000000000 : node189;
													assign node189 = (inp[11]) ? 46'b0000010000000000010010000000010100000010000000 : 46'b0000000000000000000000000000000000000000000000;
		assign node194 = (inp[15]) ? node262 : node195;
			assign node195 = (inp[13]) ? node199 : node196;
				assign node196 = (inp[3]) ? 46'b0000100000000000000000000000001000000000000000 : 46'b0000100000000000000000000000000000000000000000;
				assign node199 = (inp[2]) ? node231 : node200;
					assign node200 = (inp[11]) ? node216 : node201;
						assign node201 = (inp[0]) ? node209 : node202;
							assign node202 = (inp[9]) ? node206 : node203;
								assign node203 = (inp[3]) ? 46'b0000100000001000010000010100001000000000010010 : 46'b0000100000001000010000010100000000000000010010;
								assign node206 = (inp[3]) ? 46'b0000110000000000010000010100001000000000010010 : 46'b0000110000000000010000010100000000000000010010;
							assign node209 = (inp[9]) ? node213 : node210;
								assign node210 = (inp[3]) ? 46'b0000100000001000010000000100001100000000010010 : 46'b0000100000001000010000000100000100000000010010;
								assign node213 = (inp[3]) ? 46'b0000110000000000010000000100001100000000010010 : 46'b0000110000000000010000000100000100000000010010;
						assign node216 = (inp[9]) ? node224 : node217;
							assign node217 = (inp[0]) ? node221 : node218;
								assign node218 = (inp[3]) ? 46'b0000100000001000011000010100001000000000010000 : 46'b0000100000001000011000010100000000000000010000;
								assign node221 = (inp[3]) ? 46'b0000100000001000011000000100001100000000010000 : 46'b0000100000001000011000000100000100000000010000;
							assign node224 = (inp[0]) ? node228 : node225;
								assign node225 = (inp[3]) ? 46'b0000110000000000011000010100001000000000010000 : 46'b0000110000000000011000010100000000000000010000;
								assign node228 = (inp[3]) ? 46'b0000110000000000011000000100001100000000010000 : 46'b0000110000000000011000000100000100000000010000;
					assign node231 = (inp[0]) ? node247 : node232;
						assign node232 = (inp[11]) ? node240 : node233;
							assign node233 = (inp[9]) ? node237 : node234;
								assign node234 = (inp[3]) ? 46'b0000100000001000010010110000001000000010000000 : 46'b0000100000001000010010110000000000000010000000;
								assign node237 = (inp[3]) ? 46'b0000110000000000010010110000001000000010000000 : 46'b0000110000000000010010110000000000000010000000;
							assign node240 = (inp[9]) ? node244 : node241;
								assign node241 = (inp[3]) ? 46'b0000100000001000010010010000011000000010000000 : 46'b0000100000001000010010010000010000000010000000;
								assign node244 = (inp[3]) ? 46'b0000110000000000010010010000011000000010000000 : 46'b0000110000000000010010010000010000000010000000;
						assign node247 = (inp[11]) ? node255 : node248;
							assign node248 = (inp[9]) ? node252 : node249;
								assign node249 = (inp[3]) ? 46'b0000100000001000010010100000001100000010000000 : 46'b0000100000001000010010100000000100000010000000;
								assign node252 = (inp[3]) ? 46'b0000110000000000010010100000001100000010000000 : 46'b0000110000000000010010100000000100000010000000;
							assign node255 = (inp[9]) ? node259 : node256;
								assign node256 = (inp[3]) ? 46'b0000100000001000010010000000011100000010000000 : 46'b0000100000001000010010000000010100000010000000;
								assign node259 = (inp[3]) ? 46'b0000110000000000010010000000011100000010000000 : 46'b0000110000000000010010000000010100000010000000;
			assign node262 = (inp[13]) ? node266 : node263;
				assign node263 = (inp[3]) ? 46'b0000000000000000000000000000000000000000001000 : 46'b0000000000000000000000000000001000000000001000;
				assign node266 = (inp[3]) ? node268 : 46'b0000000000000000000000000000001000000000000000;
					assign node268 = (inp[2]) ? node906 : node269;
						assign node269 = (inp[9]) ? node661 : node270;
							assign node270 = (inp[11]) ? node510 : node271;
								assign node271 = (inp[12]) ? node381 : node272;
									assign node272 = (inp[0]) ? node328 : node273;
										assign node273 = (inp[6]) ? node305 : node274;
											assign node274 = (inp[7]) ? node288 : node275;
												assign node275 = (inp[5]) ? node283 : node276;
													assign node276 = (inp[8]) ? node280 : node277;
														assign node277 = (inp[10]) ? 46'b0011000000000000001000010001100010110001010010 : 46'b0011000000000100001000010001100010110001010000;
														assign node280 = (inp[14]) ? 46'b0011000000000010001000010001100010110001010000 : 46'b0011000000000000001000010001100010110001010010;
													assign node283 = (inp[8]) ? 46'b0010000000000000000000010001100010110001010010 : node284;
														assign node284 = (inp[14]) ? 46'b0010000000000010001000010001100010110001010000 : 46'b0010000000000100001000010001100010110001010000;
												assign node288 = (inp[4]) ? node296 : node289;
													assign node289 = (inp[10]) ? node293 : node290;
														assign node290 = (inp[14]) ? 46'b0011000000000100001000010001000010110001010000 : 46'b0011000000000100000000010000000010110001010000;
														assign node293 = (inp[5]) ? 46'b0010000000000100000000010001000010110001010010 : 46'b0011000000000100000000010001000010110001010010;
													assign node296 = (inp[14]) ? node302 : node297;
														assign node297 = (inp[8]) ? node299 : 46'b0011000000000100001000010001000010110001010000;
															assign node299 = (inp[10]) ? 46'b0011000000000010000000010001000010110001010010 : 46'b0011000000000000001000010001000010110001010010;
														assign node302 = (inp[5]) ? 46'b0010000000000010001000010001000010110001010000 : 46'b0011000000000010001000010001000010110001010000;
											assign node305 = (inp[7]) ? node317 : node306;
												assign node306 = (inp[5]) ? node314 : node307;
													assign node307 = (inp[4]) ? node311 : node308;
														assign node308 = (inp[10]) ? 46'b0011000000000000001000010001100010010001010010 : 46'b0011000000000100000000010001100010010001010010;
														assign node311 = (inp[14]) ? 46'b0011000000000010001000010001100010010001010000 : 46'b0011000000000000001000010001100010010001010010;
													assign node314 = (inp[8]) ? 46'b0010000000000010000000010001100010010001010010 : 46'b0010000000000100000000010001100010010001010010;
												assign node317 = (inp[5]) ? node321 : node318;
													assign node318 = (inp[14]) ? 46'b0011000000000000001000010001000010010001010010 : 46'b0011000000000100000000010001000010010001010010;
													assign node321 = (inp[10]) ? 46'b0010000000000000000000010001000010010001010010 : node322;
														assign node322 = (inp[4]) ? node324 : 46'b0010000000000100001000010001000010010001010000;
															assign node324 = (inp[14]) ? 46'b0010000000000000001000010001000010010001010000 : 46'b0010000000000100001000010001000010010001010000;
										assign node328 = (inp[6]) ? node356 : node329;
											assign node329 = (inp[7]) ? node349 : node330;
												assign node330 = (inp[8]) ? node338 : node331;
													assign node331 = (inp[5]) ? node333 : 46'b0011000000000100001000010001100010110000010000;
														assign node333 = (inp[4]) ? 46'b0010000000000110000000010000100010110000010000 : node334;
															assign node334 = (inp[10]) ? 46'b0010000000000100000000010001100010110000010010 : 46'b0010000000000100000000010000100010110000010000;
													assign node338 = (inp[14]) ? node344 : node339;
														assign node339 = (inp[4]) ? node341 : 46'b0011000000000000000000010001100010110000010010;
															assign node341 = (inp[5]) ? 46'b0010000000000000001000010001100010110000010010 : 46'b0011000000000000001000010001100010110000010010;
														assign node344 = (inp[4]) ? node346 : 46'b0010000000000010000000010001100010110000010010;
															assign node346 = (inp[10]) ? 46'b0010000000000010000000010000100010110000010000 : 46'b0010000000000010001000010001100010110000010000;
												assign node349 = (inp[8]) ? 46'b0010000000000010001000010001000010110000010000 : node350;
													assign node350 = (inp[4]) ? node352 : 46'b0010000000000100001000010001000010110000010000;
														assign node352 = (inp[14]) ? 46'b0010000000000000001000010001000010110000010000 : 46'b0010000000000100001000010001000010110000010000;
											assign node356 = (inp[7]) ? node370 : node357;
												assign node357 = (inp[5]) ? node367 : node358;
													assign node358 = (inp[8]) ? node364 : node359;
														assign node359 = (inp[4]) ? node361 : 46'b0011000000000100001000010001100010010000010000;
															assign node361 = (inp[14]) ? 46'b0011000000000000001000010001100010010000010000 : 46'b0011000000000100001000010001100010010000010000;
														assign node364 = (inp[4]) ? 46'b0011000000000010001000010001100010010000010000 : 46'b0011000000000110000000010000100010010000010000;
													assign node367 = (inp[10]) ? 46'b0010000000000100000000010001100010010000010010 : 46'b0010000000000100001000010001100010010000010000;
												assign node370 = (inp[5]) ? 46'b0010000000000000001000010001000010010000010010 : node371;
													assign node371 = (inp[10]) ? node373 : 46'b0011000000000110000000010000000010010000010000;
														assign node373 = (inp[4]) ? node377 : node374;
															assign node374 = (inp[8]) ? 46'b0011000000000010000000010001000010010000010010 : 46'b0011000000000000000000010001000010010000010010;
															assign node377 = (inp[14]) ? 46'b0011000000000010001000010001000010010000010000 : 46'b0011000000000110000000010000000010010000010000;
									assign node381 = (inp[0]) ? node445 : node382;
										assign node382 = (inp[7]) ? node418 : node383;
											assign node383 = (inp[5]) ? node407 : node384;
												assign node384 = (inp[10]) ? node396 : node385;
													assign node385 = (inp[4]) ? node391 : node386;
														assign node386 = (inp[8]) ? 46'b0011000000000110000000010000100000110001010000 : node387;
															assign node387 = (inp[14]) ? 46'b0011000000000100001000010001100000110001010000 : 46'b0011000000000100000000010000100000110001010000;
														assign node391 = (inp[14]) ? node393 : 46'b0011000000000100001000010001100000110001010000;
															assign node393 = (inp[8]) ? 46'b0011000000000010001000010001100000110001010000 : 46'b0011000000000000001000010001100000110001010000;
													assign node396 = (inp[8]) ? node402 : node397;
														assign node397 = (inp[14]) ? 46'b0011000000000010001000010001100000110001010000 : node398;
															assign node398 = (inp[6]) ? 46'b0011000000000110000000010000100000010001010000 : 46'b0011000000000110000000010000100000110001010000;
														assign node402 = (inp[14]) ? 46'b0011000000000010000000010000100000110001010000 : node403;
															assign node403 = (inp[4]) ? 46'b0011000000000010000000010001100000110001010010 : 46'b0011000000000000000000010001100000110001010010;
												assign node407 = (inp[10]) ? node413 : node408;
													assign node408 = (inp[8]) ? 46'b0010000000000000001000010001100000010001010010 : node409;
														assign node409 = (inp[4]) ? 46'b0010000000000100001000010001100000010001010000 : 46'b0010000000000100001000010001100000110001010000;
													assign node413 = (inp[14]) ? node415 : 46'b0010000000000100000000010001100000110001010010;
														assign node415 = (inp[8]) ? 46'b0010000000000010000000010001100000110001010010 : 46'b0010000000000010001000010001100000110001010000;
											assign node418 = (inp[8]) ? node426 : node419;
												assign node419 = (inp[14]) ? 46'b0010000000000100001000010001000000110001010000 : node420;
													assign node420 = (inp[4]) ? 46'b0010000000000110000000010000000000110001010000 : node421;
														assign node421 = (inp[6]) ? 46'b0010000000000100000000010000000000010001010000 : 46'b0010000000000100000000010000000000110001010000;
												assign node426 = (inp[6]) ? node438 : node427;
													assign node427 = (inp[4]) ? node433 : node428;
														assign node428 = (inp[10]) ? 46'b0010000000000010000000010001000000110001010010 : node429;
															assign node429 = (inp[5]) ? 46'b0010000000000110000000010000000000110001010000 : 46'b0011000000000110000000010000000000110001010000;
														assign node433 = (inp[14]) ? 46'b0010000000000010001000010001000000110001010000 : node434;
															assign node434 = (inp[10]) ? 46'b0010000000000010000000010001000000110001010010 : 46'b0011000000000000001000010001000000110001010010;
													assign node438 = (inp[10]) ? node442 : node439;
														assign node439 = (inp[5]) ? 46'b0010000000000010001000010001000000010001010000 : 46'b0011000000000010001000010001000000010001010000;
														assign node442 = (inp[4]) ? 46'b0011000000000010000000010000000000010001010000 : 46'b0011000000000010000000010001000000010001010010;
										assign node445 = (inp[6]) ? node475 : node446;
											assign node446 = (inp[7]) ? node466 : node447;
												assign node447 = (inp[5]) ? node461 : node448;
													assign node448 = (inp[14]) ? node454 : node449;
														assign node449 = (inp[8]) ? 46'b0011000000000100000000010001100000110000010010 : node450;
															assign node450 = (inp[4]) ? 46'b0011000000000110000000010000100000110000010000 : 46'b0011000000000100000000010000100000110000010000;
														assign node454 = (inp[8]) ? node458 : node455;
															assign node455 = (inp[10]) ? 46'b0011000000000000001000010001100000110000010010 : 46'b0011000000000000001000010001100000110000010000;
															assign node458 = (inp[4]) ? 46'b0011000000000010001000010001100000110000010000 : 46'b0011000000000010000000010000100000110000010000;
													assign node461 = (inp[14]) ? node463 : 46'b0010000000000100000000010001100000110000010010;
														assign node463 = (inp[8]) ? 46'b0010000000000110000000010000100000110000010000 : 46'b0010000000000100001000010001100000110000010000;
												assign node466 = (inp[4]) ? node472 : node467;
													assign node467 = (inp[14]) ? node469 : 46'b0010000000000100000000010001000000110000010010;
														assign node469 = (inp[5]) ? 46'b0010000000000010000000010001000000110000010010 : 46'b0011000000000010000000010001000000110000010010;
													assign node472 = (inp[8]) ? 46'b0010000000000010000000010000000000110000010000 : 46'b0010000000000010001000010001000000110000010000;
											assign node475 = (inp[5]) ? node493 : node476;
												assign node476 = (inp[7]) ? node486 : node477;
													assign node477 = (inp[10]) ? node483 : node478;
														assign node478 = (inp[14]) ? node480 : 46'b0011000000000000001000010001100000010000010010;
															assign node480 = (inp[4]) ? 46'b0011000000000000001000010001100000010000010000 : 46'b0011000000000100001000010001100000010000010000;
														assign node483 = (inp[4]) ? 46'b0011000000000010000000010001100000010000010010 : 46'b0011000000000100000000010001100000010000010010;
													assign node486 = (inp[4]) ? node490 : node487;
														assign node487 = (inp[8]) ? 46'b0011000000000000000000010001000000010000010010 : 46'b0011000000000000001000010001000000010000010010;
														assign node490 = (inp[10]) ? 46'b0011000000000110000000010000000000010000010000 : 46'b0011000000000010001000010001000000010000010000;
												assign node493 = (inp[4]) ? node501 : node494;
													assign node494 = (inp[7]) ? node498 : node495;
														assign node495 = (inp[14]) ? 46'b0010000000000010000000010001100000010000010010 : 46'b0010000000000000000000010001100000010000010010;
														assign node498 = (inp[14]) ? 46'b0010000000000000001000010001000000010000010010 : 46'b0010000000000100000000010001000000010000010010;
													assign node501 = (inp[7]) ? node507 : node502;
														assign node502 = (inp[10]) ? 46'b0010000000000010000000010000100000010000010000 : node503;
															assign node503 = (inp[14]) ? 46'b0010000000000010001000010001100000010000010000 : 46'b0010000000000100001000010001100000010000010000;
														assign node507 = (inp[14]) ? 46'b0010000000000010001000010001000000010000010000 : 46'b0010000000000010000000010001000000010000010010;
								assign node510 = (inp[0]) ? node536 : node511;
									assign node511 = (inp[7]) ? node513 : 46'b0000000000000000000000000000000000000000000000;
										assign node513 = (inp[5]) ? node515 : 46'b0000000000000000000000000000000000000000000000;
											assign node515 = (inp[4]) ? node523 : node516;
												assign node516 = (inp[10]) ? node518 : 46'b0000000000000000000000000000000000000000000000;
													assign node518 = (inp[12]) ? 46'b0000000000000100000001000001000000100000000010 : node519;
														assign node519 = (inp[6]) ? 46'b0000000000000000000001000001000010000000000010 : 46'b0000000000000000000000000000000000000000000000;
												assign node523 = (inp[14]) ? node529 : node524;
													assign node524 = (inp[10]) ? node526 : 46'b0000000000000000000000000000000000000000000000;
														assign node526 = (inp[6]) ? 46'b0000000000000110000001000000000010000000000000 : 46'b0000000000000000000000000000000000000000000000;
													assign node529 = (inp[10]) ? node533 : node530;
														assign node530 = (inp[8]) ? 46'b0000000000000010001001000001000000100000000000 : 46'b0000000000000000001001000001000000100000000000;
														assign node533 = (inp[6]) ? 46'b0000000000000000000000000000000000000000000000 : 46'b0000000000000010000001000000000000100000000000;
									assign node536 = (inp[12]) ? node600 : node537;
										assign node537 = (inp[6]) ? node569 : node538;
											assign node538 = (inp[7]) ? node558 : node539;
												assign node539 = (inp[14]) ? node549 : node540;
													assign node540 = (inp[8]) ? node546 : node541;
														assign node541 = (inp[5]) ? 46'b0100000000000100000000000001100010100000000010 : node542;
															assign node542 = (inp[10]) ? 46'b0101000000000110000000000000100010100000000000 : 46'b0101000000000100000000000000100010100000000000;
														assign node546 = (inp[10]) ? 46'b0101000000000010000000000001100010100000000010 : 46'b0101000000000000001000000001100010100000000010;
													assign node549 = (inp[10]) ? node555 : node550;
														assign node550 = (inp[8]) ? node552 : 46'b0100000000000000001000000001100010100000000000;
															assign node552 = (inp[5]) ? 46'b0100000000000010001000000001100010100000000000 : 46'b0101000000000010001000000001100010100000000000;
														assign node555 = (inp[5]) ? 46'b0100000000000010000000000000100010100000000000 : 46'b0101000000000010000000000000100010100000000000;
												assign node558 = (inp[4]) ? node566 : node559;
													assign node559 = (inp[5]) ? node563 : node560;
														assign node560 = (inp[14]) ? 46'b0101000000000000001000000001000010100000000010 : 46'b0101000000000100000000000001000010100000000010;
														assign node563 = (inp[14]) ? 46'b0100000000000010000000000001000010100000000010 : 46'b0100000000000000000000000001000010100000000010;
													assign node566 = (inp[5]) ? 46'b0100000000000010000000000000000010100000000000 : 46'b0101000000000010000000000000000010100000000000;
											assign node569 = (inp[10]) ? node583 : node570;
												assign node570 = (inp[5]) ? node578 : node571;
													assign node571 = (inp[7]) ? node575 : node572;
														assign node572 = (inp[8]) ? 46'b0101000000000100000000000001100010000000000010 : 46'b0101000000000100000000000000100010000000000000;
														assign node575 = (inp[8]) ? 46'b0101000000000110000000000000000010000000000000 : 46'b0101000000000100000000000000000010000000000000;
													assign node578 = (inp[8]) ? 46'b0100000000000100000000000001100010000000000010 : node579;
														assign node579 = (inp[7]) ? 46'b0100000000000100001000000001000010000000000000 : 46'b0100000000000100001000000001100010000000000000;
												assign node583 = (inp[4]) ? node591 : node584;
													assign node584 = (inp[14]) ? node588 : node585;
														assign node585 = (inp[8]) ? 46'b0101000000000000000000000001100010000000000010 : 46'b0101000000000100000000000001100010000000000010;
														assign node588 = (inp[7]) ? 46'b0101000000000010000000000001000010000000000010 : 46'b0101000000000010000000000001100010000000000010;
													assign node591 = (inp[8]) ? node595 : node592;
														assign node592 = (inp[5]) ? 46'b0100000000000010001000000001100010000000000000 : 46'b0101000000000010001000000001100010000000000000;
														assign node595 = (inp[14]) ? 46'b0100000000000010000000000000100010000000000000 : node596;
															assign node596 = (inp[7]) ? 46'b0100000000000010000000000001000010000000000010 : 46'b0100000000000010000000000001100010000000000010;
										assign node600 = (inp[5]) ? node636 : node601;
											assign node601 = (inp[7]) ? node619 : node602;
												assign node602 = (inp[6]) ? node608 : node603;
													assign node603 = (inp[8]) ? 46'b0101000000000010000000000001100000100000000010 : node604;
														assign node604 = (inp[10]) ? 46'b0101000000000010001000000001100000100000000000 : 46'b0101000000000000001000000001100000100000000000;
													assign node608 = (inp[4]) ? node616 : node609;
														assign node609 = (inp[10]) ? node613 : node610;
															assign node610 = (inp[14]) ? 46'b0101000000000110000000000000100000000000000000 : 46'b0101000000000100000000000000100000000000000000;
															assign node613 = (inp[14]) ? 46'b0101000000000000001000000001100000000000000010 : 46'b0101000000000100000000000001100000000000000010;
														assign node616 = (inp[10]) ? 46'b0101000000000010000000000001100000000000000010 : 46'b0101000000000010001000000001100000000000000000;
												assign node619 = (inp[6]) ? node625 : node620;
													assign node620 = (inp[10]) ? 46'b0101000000000100000000000001000000100000000010 : node621;
														assign node621 = (inp[14]) ? 46'b0101000000000110000000000000000000100000000000 : 46'b0101000000000100000000000000000000100000000000;
													assign node625 = (inp[10]) ? node631 : node626;
														assign node626 = (inp[8]) ? 46'b0101000000000000001000000001000000000000000010 : node627;
															assign node627 = (inp[14]) ? 46'b0101000000000100001000000001000000000000000000 : 46'b0101000000000100000000000000000000000000000000;
														assign node631 = (inp[8]) ? node633 : 46'b0101000000000000001000000001000000000000000010;
															assign node633 = (inp[14]) ? 46'b0101000000000010000000000001000000000000000010 : 46'b0101000000000000000000000001000000000000000010;
											assign node636 = (inp[6]) ? node650 : node637;
												assign node637 = (inp[7]) ? node641 : node638;
													assign node638 = (inp[8]) ? 46'b0100000000000110000000000000100000100000000000 : 46'b0100000000000100001000000001100000100000000000;
													assign node641 = (inp[14]) ? node645 : node642;
														assign node642 = (inp[8]) ? 46'b0100000000000100000000000001000000100000000010 : 46'b0100000000000100000000000000000000100000000000;
														assign node645 = (inp[8]) ? 46'b0100000000000010000000000001000000100000000010 : node646;
															assign node646 = (inp[4]) ? 46'b0100000000000000001000000001000000100000000000 : 46'b0100000000000000001000000001000000100000000010;
												assign node650 = (inp[10]) ? node658 : node651;
													assign node651 = (inp[8]) ? 46'b0100000000000010001000000001000000000000000000 : node652;
														assign node652 = (inp[7]) ? node654 : 46'b0100000000000000001000000001100000000000000000;
															assign node654 = (inp[14]) ? 46'b0100000000000100001000000001000000000000000000 : 46'b0100000000000100000000000000000000000000000000;
													assign node658 = (inp[7]) ? 46'b0100000000000100000000000001000000000000000010 : 46'b0100000000000100000000000001100000000000000010;
							assign node661 = (inp[11]) ? node701 : node662;
								assign node662 = (inp[0]) ? 46'b0000000000000000000000000000000000000000000000 : node663;
									assign node663 = (inp[7]) ? node687 : node664;
										assign node664 = (inp[5]) ? node666 : 46'b0000000000000000000000000000000000000000000000;
											assign node666 = (inp[4]) ? node680 : node667;
												assign node667 = (inp[14]) ? node675 : node668;
													assign node668 = (inp[12]) ? 46'b0000000000000000000000001001100000100000000010 : node669;
														assign node669 = (inp[10]) ? node671 : 46'b0000000000000100000000001001100010100000000010;
															assign node671 = (inp[8]) ? 46'b0000000000000000000000001001100010100000000010 : 46'b0000000000000100000000001001100010100000000010;
													assign node675 = (inp[10]) ? node677 : 46'b0000000000000000000000000000000000000000000000;
														assign node677 = (inp[12]) ? 46'b0000000000000000001000001001100000000000000010 : 46'b0000000000000000001000001001100010000000000010;
												assign node680 = (inp[8]) ? node682 : 46'b0000000000000000000000000000000000000000000000;
													assign node682 = (inp[14]) ? 46'b0000000000000000000000000000000000000000000000 : node683;
														assign node683 = (inp[12]) ? 46'b0000000000000010000000001001100000000000000010 : 46'b0000000000000000001000001001100010100000000010;
										assign node687 = (inp[5]) ? 46'b0000000000000000000000000000000000000000000000 : node688;
											assign node688 = (inp[6]) ? node692 : node689;
												assign node689 = (inp[10]) ? 46'b0000000000000000000000000000000000000000000000 : 46'b0001000000000100000000001000000000100000000000;
												assign node692 = (inp[14]) ? node696 : node693;
													assign node693 = (inp[10]) ? 46'b0001000000000110000000001000000010000000000000 : 46'b0001000000000100000000001000000000000000000000;
													assign node696 = (inp[12]) ? 46'b0001000000000100001000001001000000000000000000 : 46'b0001000000000100001000001001000010000000000000;
								assign node701 = (inp[0]) ? node797 : node702;
									assign node702 = (inp[7]) ? node758 : node703;
										assign node703 = (inp[6]) ? node727 : node704;
											assign node704 = (inp[12]) ? node716 : node705;
												assign node705 = (inp[8]) ? node711 : node706;
													assign node706 = (inp[4]) ? node708 : 46'b1001000000000100001000000001100010100000000000;
														assign node708 = (inp[14]) ? 46'b1000000000000000001000000001100010100000000000 : 46'b1000000000000100001000000001100010100000000000;
													assign node711 = (inp[10]) ? node713 : 46'b1001000000000110000000000000100010100000000000;
														assign node713 = (inp[5]) ? 46'b1000000000000000000000000001100010100000000010 : 46'b1001000000000010000000000001100010100000000010;
												assign node716 = (inp[4]) ? node720 : node717;
													assign node717 = (inp[8]) ? 46'b1001000000000000000000000001100000100000000010 : 46'b1000000000000000001000000001100000100000000010;
													assign node720 = (inp[8]) ? node724 : node721;
														assign node721 = (inp[14]) ? 46'b1001000000000000001000000001100000100000000000 : 46'b1001000000000100001000000001100000100000000000;
														assign node724 = (inp[14]) ? 46'b1001000000000010001000000001100000100000000000 : 46'b1001000000000000001000000001100000100000000010;
											assign node727 = (inp[5]) ? node741 : node728;
												assign node728 = (inp[14]) ? node734 : node729;
													assign node729 = (inp[12]) ? node731 : 46'b1001000000000100000000000001100010000000000010;
														assign node731 = (inp[10]) ? 46'b1001000000000000000000000001100000000000000010 : 46'b1001000000000000001000000001100000000000000010;
													assign node734 = (inp[8]) ? node736 : 46'b1001000000000100001000000001100010000000000000;
														assign node736 = (inp[12]) ? 46'b1001000000000110000000000000100000000000000000 : node737;
															assign node737 = (inp[4]) ? 46'b1001000000000010000000000000100010000000000000 : 46'b1001000000000110000000000000100010000000000000;
												assign node741 = (inp[12]) ? node747 : node742;
													assign node742 = (inp[14]) ? node744 : 46'b1000000000000100000000000001100010000000000010;
														assign node744 = (inp[4]) ? 46'b1000000000000010001000000001100010000000000000 : 46'b1000000000000100001000000001100010000000000000;
													assign node747 = (inp[10]) ? node755 : node748;
														assign node748 = (inp[4]) ? node752 : node749;
															assign node749 = (inp[14]) ? 46'b1000000000000100001000000001100000000000000000 : 46'b1000000000000100000000000000100000000000000000;
															assign node752 = (inp[14]) ? 46'b1000000000000000001000000001100000000000000000 : 46'b1000000000000100001000000001100000000000000000;
														assign node755 = (inp[14]) ? 46'b1000000000000010000000000000100000000000000000 : 46'b1000000000000110000000000000100000000000000000;
										assign node758 = (inp[12]) ? node782 : node759;
											assign node759 = (inp[4]) ? node779 : node760;
												assign node760 = (inp[5]) ? node766 : node761;
													assign node761 = (inp[14]) ? node763 : 46'b1001000000000100000000000001000010100000000010;
														assign node763 = (inp[6]) ? 46'b1001000000000100001000000001000010000000000000 : 46'b1001000000000100001000000001000010100000000000;
													assign node766 = (inp[10]) ? node774 : node767;
														assign node767 = (inp[8]) ? node771 : node768;
															assign node768 = (inp[6]) ? 46'b1000000000000100000000000000000010000000000000 : 46'b1000000000000100000000000000000010100000000000;
															assign node771 = (inp[6]) ? 46'b1000000000000100000000000001000010000000000010 : 46'b1000000000000100000000000001000010100000000010;
														assign node774 = (inp[8]) ? 46'b1000000000000000000000000001000010000000000010 : node775;
															assign node775 = (inp[14]) ? 46'b1000000000000000001000000001000010100000000010 : 46'b1000000000000100000000000001000010100000000010;
												assign node779 = (inp[8]) ? 46'b1001000000000010000000000000000010100000000000 : 46'b1001000000000110000000000000000010100000000000;
											assign node782 = (inp[5]) ? node794 : node783;
												assign node783 = (inp[6]) ? node789 : node784;
													assign node784 = (inp[8]) ? node786 : 46'b1001000000000000001000000001000000100000000010;
														assign node786 = (inp[4]) ? 46'b1001000000000000001000000001000000100000000010 : 46'b1001000000000010000000000001000000100000000010;
													assign node789 = (inp[14]) ? node791 : 46'b1001000000000100000000000001000000000000000010;
														assign node791 = (inp[4]) ? 46'b1001000000000010001000000001000000000000000000 : 46'b1001000000000100001000000001000000000000000000;
												assign node794 = (inp[10]) ? 46'b1000000000000110000000000000000000100000000000 : 46'b1000000000000100001000000001000000100000000000;
									assign node797 = (inp[5]) ? node853 : node798;
										assign node798 = (inp[12]) ? node824 : node799;
											assign node799 = (inp[4]) ? node815 : node800;
												assign node800 = (inp[10]) ? node804 : node801;
													assign node801 = (inp[14]) ? 46'b0001000000000100001000000001000010001000000000 : 46'b0001000000000100000000000000000010001000000000;
													assign node804 = (inp[14]) ? node810 : node805;
														assign node805 = (inp[8]) ? 46'b0001000000000000000000000001000010001000000010 : node806;
															assign node806 = (inp[7]) ? 46'b0001000000000100000000000001000010001000000010 : 46'b0001000000000100000000000001100010001000000010;
														assign node810 = (inp[6]) ? node812 : 46'b0001000000000000001000000001000010101000000010;
															assign node812 = (inp[7]) ? 46'b0001000000000000001000000001000010001000000010 : 46'b0001000000000000001000000001100010001000000010;
												assign node815 = (inp[7]) ? 46'b0001000000000010000000000001000010001000000010 : node816;
													assign node816 = (inp[10]) ? node818 : 46'b0001000000000000001000000001100010101000000000;
														assign node818 = (inp[8]) ? 46'b0001000000000010000000000000100010101000000000 : node819;
															assign node819 = (inp[6]) ? 46'b0001000000000110000000000000100010001000000000 : 46'b0001000000000110000000000000100010101000000000;
											assign node824 = (inp[6]) ? node838 : node825;
												assign node825 = (inp[10]) ? node833 : node826;
													assign node826 = (inp[4]) ? node830 : node827;
														assign node827 = (inp[14]) ? 46'b0001000000000100001000000001000000101000000000 : 46'b0001000000000100000000000000000000101000000000;
														assign node830 = (inp[8]) ? 46'b0001000000000010001000000001000000101000000000 : 46'b0001000000000000001000000001100000101000000000;
													assign node833 = (inp[7]) ? 46'b0001000000000000000000000001000000101000000010 : node834;
														assign node834 = (inp[4]) ? 46'b0001000000000010000000000001100000101000000010 : 46'b0001000000000000000000000001100000101000000010;
												assign node838 = (inp[14]) ? node842 : node839;
													assign node839 = (inp[10]) ? 46'b0001000000000110000000000000100000001000000000 : 46'b0001000000000100000000000000100000001000000000;
													assign node842 = (inp[4]) ? node848 : node843;
														assign node843 = (inp[10]) ? node845 : 46'b0001000000000110000000000000000000001000000000;
															assign node845 = (inp[8]) ? 46'b0001000000000010000000000001000000001000000010 : 46'b0001000000000000001000000001000000001000000010;
														assign node848 = (inp[7]) ? node850 : 46'b0001000000000010001000000001100000001000000000;
															assign node850 = (inp[8]) ? 46'b0001000000000010000000000000000000001000000000 : 46'b0001000000000010001000000001000000001000000000;
										assign node853 = (inp[10]) ? node887 : node854;
											assign node854 = (inp[4]) ? node872 : node855;
												assign node855 = (inp[12]) ? node865 : node856;
													assign node856 = (inp[8]) ? node862 : node857;
														assign node857 = (inp[7]) ? node859 : 46'b0000000000000100001000000001100010001000000000;
															assign node859 = (inp[6]) ? 46'b0000000000000100001000000001000010001000000000 : 46'b0000000000000100001000000001000010101000000000;
														assign node862 = (inp[7]) ? 46'b0000000000000110000000000000000010101000000000 : 46'b0000000000000110000000000000100010001000000000;
													assign node865 = (inp[14]) ? 46'b0000000000000100001000000001100000001000000000 : node866;
														assign node866 = (inp[8]) ? 46'b0000000000000100000000000001100000001000000010 : node867;
															assign node867 = (inp[7]) ? 46'b0000000000000100000000000000000000001000000000 : 46'b0000000000000100000000000000100000001000000000;
												assign node872 = (inp[12]) ? node880 : node873;
													assign node873 = (inp[14]) ? node877 : node874;
														assign node874 = (inp[6]) ? 46'b0000000000000100001000000001100010001000000000 : 46'b0000000000000100001000000001100010101000000000;
														assign node877 = (inp[6]) ? 46'b0000000000000000001000000001100010001000000000 : 46'b0000000000000000001000000001100010101000000000;
													assign node880 = (inp[8]) ? node884 : node881;
														assign node881 = (inp[14]) ? 46'b0000000000000000001000000001100000101000000000 : 46'b0000000000000100001000000001100000101000000000;
														assign node884 = (inp[6]) ? 46'b0000000000000000001000000001100000001000000010 : 46'b0000000000000000001000000001100000101000000010;
											assign node887 = (inp[7]) ? node903 : node888;
												assign node888 = (inp[12]) ? node896 : node889;
													assign node889 = (inp[8]) ? node891 : 46'b0000000000000000001000000001100010001000000010;
														assign node891 = (inp[14]) ? node893 : 46'b0000000000000000000000000001100010101000000010;
															assign node893 = (inp[6]) ? 46'b0000000000000010000000000001100010001000000010 : 46'b0000000000000010000000000001100010101000000010;
													assign node896 = (inp[4]) ? 46'b0000000000000010000000000000100000101000000000 : node897;
														assign node897 = (inp[14]) ? 46'b0000000000000010000000000001100000101000000010 : node898;
															assign node898 = (inp[8]) ? 46'b0000000000000000000000000001100000101000000010 : 46'b0000000000000100000000000001100000101000000010;
												assign node903 = (inp[6]) ? 46'b0000000000000000001000000001000000001000000010 : 46'b0000000000000000001000000001000000101000000010;
						assign node906 = (inp[11]) ? node1218 : node907;
							assign node907 = (inp[9]) ? node987 : node908;
								assign node908 = (inp[5]) ? node922 : node909;
									assign node909 = (inp[0]) ? node911 : 46'b0000000000000000000000000000000000000000000000;
										assign node911 = (inp[12]) ? node913 : 46'b0000000000000000000000000000000000000000000000;
											assign node913 = (inp[7]) ? node915 : 46'b0000000000000000000000000000000000000000000000;
												assign node915 = (inp[6]) ? node917 : 46'b0000000000000000000000000000000000000000000000;
													assign node917 = (inp[14]) ? node919 : 46'b0001000000000101000000000001000000000000100010;
														assign node919 = (inp[4]) ? 46'b0001000000000011001000000001000000000000100000 : 46'b0001000000000001001000000001000000000000100010;
									assign node922 = (inp[7]) ? node938 : node923;
										assign node923 = (inp[0]) ? node925 : 46'b0000000000000000000000000000000000000000000000;
											assign node925 = (inp[12]) ? node927 : 46'b0000000000000000000000000000000000000000000000;
												assign node927 = (inp[6]) ? node929 : 46'b0000000000000000000000000000000000000000000000;
													assign node929 = (inp[8]) ? node933 : node930;
														assign node930 = (inp[14]) ? 46'b0000000000000101001000000001100000000000100000 : 46'b0000000000000101000000000000100000000000100000;
														assign node933 = (inp[10]) ? node935 : 46'b0000000000000001001000000001100000000000100010;
															assign node935 = (inp[4]) ? 46'b0000000000000011000000000001100000000000100010 : 46'b0000000000000001000000000001100000000000100010;
										assign node938 = (inp[0]) ? node968 : node939;
											assign node939 = (inp[10]) ? node951 : node940;
												assign node940 = (inp[6]) ? node944 : node941;
													assign node941 = (inp[12]) ? 46'b0000000000100100001001000001000000100000000000 : 46'b0000000000100100001001000001000010100000000000;
													assign node944 = (inp[4]) ? node948 : node945;
														assign node945 = (inp[8]) ? 46'b0000000000100100000001000001000000000000000010 : 46'b0000000000100100000001000000000000000000000000;
														assign node948 = (inp[12]) ? 46'b0000000000100100001001000001000000000000000000 : 46'b0000000000100100001001000001000010000000000000;
												assign node951 = (inp[12]) ? node961 : node952;
													assign node952 = (inp[8]) ? node956 : node953;
														assign node953 = (inp[4]) ? 46'b0000000000100010001001000001000010100000000000 : 46'b0000000000100000001001000001000010000000000010;
														assign node956 = (inp[6]) ? node958 : 46'b0000000000100010000001000001000010100000000010;
															assign node958 = (inp[4]) ? 46'b0000000000100010000001000000000010000000000000 : 46'b0000000000100010000001000001000010000000000010;
													assign node961 = (inp[6]) ? 46'b0000000000100010000001000001000000000000000010 : node962;
														assign node962 = (inp[8]) ? node964 : 46'b0000000000100100000001000001000000100000000010;
															assign node964 = (inp[4]) ? 46'b0000000000100010000001000001000000100000000010 : 46'b0000000000100000000001000001000000100000000010;
											assign node968 = (inp[6]) ? node976 : node969;
												assign node969 = (inp[12]) ? node971 : 46'b0000000000000000000000000000000000000000000000;
													assign node971 = (inp[8]) ? 46'b0000000000000001001000000001000000100000100010 : node972;
														assign node972 = (inp[14]) ? 46'b0000000000000101001000000001000000100000100000 : 46'b0000000000000101000000000000000000100000100000;
												assign node976 = (inp[12]) ? 46'b0000000000000000000000000000000000000000000000 : node977;
													assign node977 = (inp[14]) ? node983 : node978;
														assign node978 = (inp[10]) ? node980 : 46'b0000000000000101000000000001000010000000100010;
															assign node980 = (inp[8]) ? 46'b0000000000000001000000000001000010000000100010 : 46'b0000000000000101000000000001000010000000100010;
														assign node983 = (inp[4]) ? 46'b0000000000000011001000000001000010000000100000 : 46'b0000000000000001001000000001000010000000100010;
								assign node987 = (inp[0]) ? node1105 : node988;
									assign node988 = (inp[12]) ? node1040 : node989;
										assign node989 = (inp[7]) ? node1021 : node990;
											assign node990 = (inp[6]) ? node1006 : node991;
												assign node991 = (inp[8]) ? node1001 : node992;
													assign node992 = (inp[4]) ? node996 : node993;
														assign node993 = (inp[10]) ? 46'b0000000000100000001000000001100010100000100010 : 46'b0000000000100100001000000001100010100000100000;
														assign node996 = (inp[10]) ? node998 : 46'b0001000000100100001000000001100010100000100000;
															assign node998 = (inp[5]) ? 46'b0000000000100110000000000000100010100000100000 : 46'b0001000000100110000000000000100010100000100000;
													assign node1001 = (inp[4]) ? node1003 : 46'b0001000000100010000000000001100010100000100010;
														assign node1003 = (inp[5]) ? 46'b0000000000100000001000000001100010100000100010 : 46'b0001000000100000001000000001100010100000100010;
												assign node1006 = (inp[5]) ? node1014 : node1007;
													assign node1007 = (inp[14]) ? node1011 : node1008;
														assign node1008 = (inp[10]) ? 46'b0001000000100000000000000001100010000000100010 : 46'b0001000000100100000000000000100010000000100000;
														assign node1011 = (inp[10]) ? 46'b0001000000100000001000000001100010000000100010 : 46'b0001000000100010001000000001100010000000100000;
													assign node1014 = (inp[10]) ? node1016 : 46'b0000000000100000001000000001100010000000100000;
														assign node1016 = (inp[4]) ? node1018 : 46'b0000000000100010000000000001100010000000100010;
															assign node1018 = (inp[8]) ? 46'b0000000000100010000000000000100010000000100000 : 46'b0000000000100110000000000000100010000000100000;
											assign node1021 = (inp[5]) ? node1027 : node1022;
												assign node1022 = (inp[8]) ? node1024 : 46'b0001000000100100000000000000000010100000100000;
													assign node1024 = (inp[14]) ? 46'b0001000000100010000000000000000010000000100000 : 46'b0001000000100000001000000001000010000000100010;
												assign node1027 = (inp[6]) ? node1031 : node1028;
													assign node1028 = (inp[8]) ? 46'b0000000000100000000000000001000010100000100010 : 46'b0000000000100000001000000001000010100000100010;
													assign node1031 = (inp[4]) ? node1037 : node1032;
														assign node1032 = (inp[10]) ? node1034 : 46'b0000000000100110000000000000000010000000100000;
															assign node1034 = (inp[14]) ? 46'b0000000000100000001000000001000010000000100010 : 46'b0000000000100100000000000001000010000000100010;
														assign node1037 = (inp[8]) ? 46'b0000000000100000001000000001000010000000100010 : 46'b0000000000100000001000000001000010000000100000;
										assign node1040 = (inp[7]) ? node1070 : node1041;
											assign node1041 = (inp[5]) ? node1059 : node1042;
												assign node1042 = (inp[6]) ? node1054 : node1043;
													assign node1043 = (inp[10]) ? node1049 : node1044;
														assign node1044 = (inp[14]) ? 46'b0001000000100110000000000000100000100000100000 : node1045;
															assign node1045 = (inp[8]) ? 46'b0001000000100100000000000001100000100000100010 : 46'b0001000000100100000000000000100000100000100000;
														assign node1049 = (inp[4]) ? 46'b0001000000100110000000000000100000100000100000 : node1050;
															assign node1050 = (inp[8]) ? 46'b0001000000100010000000000001100000100000100010 : 46'b0001000000100000001000000001100000100000100010;
													assign node1054 = (inp[14]) ? 46'b0001000000100010000000000000100000000000100000 : node1055;
														assign node1055 = (inp[4]) ? 46'b0001000000100000001000000001100000000000100010 : 46'b0001000000100100000000000001100000000000100010;
												assign node1059 = (inp[14]) ? node1063 : node1060;
													assign node1060 = (inp[4]) ? 46'b0000000000100010000000000001100000100000100010 : 46'b0000000000100000000000000001100000100000100010;
													assign node1063 = (inp[8]) ? node1067 : node1064;
														assign node1064 = (inp[6]) ? 46'b0000000000100100001000000001100000000000100000 : 46'b0000000000100100001000000001100000100000100000;
														assign node1067 = (inp[6]) ? 46'b0000000000100110000000000000100000000000100000 : 46'b0000000000100110000000000000100000100000100000;
											assign node1070 = (inp[5]) ? node1088 : node1071;
												assign node1071 = (inp[4]) ? node1077 : node1072;
													assign node1072 = (inp[10]) ? node1074 : 46'b0001000000100100000000000001000000000000100010;
														assign node1074 = (inp[6]) ? 46'b0001000000100000001000000001000000000000100010 : 46'b0001000000100000001000000001000000100000100010;
													assign node1077 = (inp[10]) ? node1081 : node1078;
														assign node1078 = (inp[8]) ? 46'b0001000000100000001000000001000000100000100010 : 46'b0001000000100100001000000001000000100000100000;
														assign node1081 = (inp[6]) ? node1085 : node1082;
															assign node1082 = (inp[8]) ? 46'b0001000000100010000000000000000000100000100000 : 46'b0001000000100110000000000000000000100000100000;
															assign node1085 = (inp[8]) ? 46'b0001000000100010000000000000000000000000100000 : 46'b0001000000100010001000000001000000000000100000;
												assign node1088 = (inp[10]) ? node1098 : node1089;
													assign node1089 = (inp[4]) ? node1095 : node1090;
														assign node1090 = (inp[6]) ? 46'b0000000000100100000000000001000000000000100010 : node1091;
															assign node1091 = (inp[14]) ? 46'b0000000000100110000000000000000000100000100000 : 46'b0000000000100100000000000000000000100000100000;
														assign node1095 = (inp[8]) ? 46'b0000000000100000001000000001000000100000100010 : 46'b0000000000100100001000000001000000100000100000;
													assign node1098 = (inp[4]) ? node1102 : node1099;
														assign node1099 = (inp[14]) ? 46'b0000000000100000001000000001000000100000100010 : 46'b0000000000100000000000000001000000100000100010;
														assign node1102 = (inp[6]) ? 46'b0000000000100010000000000001000000000000100010 : 46'b0000000000100010000000000001000000100000100010;
									assign node1105 = (inp[5]) ? node1161 : node1106;
										assign node1106 = (inp[6]) ? node1128 : node1107;
											assign node1107 = (inp[10]) ? node1119 : node1108;
												assign node1108 = (inp[8]) ? node1116 : node1109;
													assign node1109 = (inp[12]) ? 46'b0001000000000100001000000001000000100000100000 : node1110;
														assign node1110 = (inp[4]) ? node1112 : 46'b0001000000000100001000000001000010100000100000;
															assign node1112 = (inp[14]) ? 46'b0001000000000000001000000001000010100000100000 : 46'b0001000000000100001000000001000010100000100000;
													assign node1116 = (inp[14]) ? 46'b0001000000000110000000000000000010100000100000 : 46'b0001000000000100000000000001000010100000100010;
												assign node1119 = (inp[4]) ? 46'b0001000000000010001000000001100000100000100000 : node1120;
													assign node1120 = (inp[12]) ? node1124 : node1121;
														assign node1121 = (inp[7]) ? 46'b0001000000000000001000000001000010100000100010 : 46'b0001000000000000001000000001100010100000100010;
														assign node1124 = (inp[7]) ? 46'b0001000000000000001000000001000000100000100010 : 46'b0001000000000000001000000001100000100000100010;
											assign node1128 = (inp[8]) ? node1146 : node1129;
												assign node1129 = (inp[7]) ? node1137 : node1130;
													assign node1130 = (inp[10]) ? node1134 : node1131;
														assign node1131 = (inp[14]) ? 46'b0001000000000000001000000001100010000000100000 : 46'b0001000000000100000000000000100010000000100000;
														assign node1134 = (inp[12]) ? 46'b0001000000000100000000000001100000000000100010 : 46'b0001000000000100000000000001100010000000100010;
													assign node1137 = (inp[14]) ? node1143 : node1138;
														assign node1138 = (inp[10]) ? 46'b0001000000000110000000000000000010000000100000 : node1139;
															assign node1139 = (inp[4]) ? 46'b0001000000000100001000000001000010000000100000 : 46'b0001000000000100000000000000000000000000100000;
														assign node1143 = (inp[12]) ? 46'b0001000000000100001000000001000000000000100000 : 46'b0001000000000100001000000001000010000000100000;
												assign node1146 = (inp[14]) ? node1152 : node1147;
													assign node1147 = (inp[7]) ? node1149 : 46'b0001000000000010000000000001100010000000100010;
														assign node1149 = (inp[10]) ? 46'b0001000000000000000000000001000000000000100010 : 46'b0001000000000000001000000001000010000000100010;
													assign node1152 = (inp[12]) ? node1156 : node1153;
														assign node1153 = (inp[10]) ? 46'b0001000000000010000000000000000010000000100000 : 46'b0001000000000110000000000000000010000000100000;
														assign node1156 = (inp[7]) ? 46'b0001000000000010000000000001000000000000100010 : node1157;
															assign node1157 = (inp[10]) ? 46'b0001000000000010000000000000100000000000100000 : 46'b0001000000000010001000000001100000000000100000;
										assign node1161 = (inp[6]) ? node1185 : node1162;
											assign node1162 = (inp[7]) ? node1170 : node1163;
												assign node1163 = (inp[12]) ? 46'b0000000000000100001000000001100000100000100000 : node1164;
													assign node1164 = (inp[8]) ? node1166 : 46'b0000000000000100000000000001100010100000100010;
														assign node1166 = (inp[4]) ? 46'b0000000000000010000000000001100010100000100010 : 46'b0000000000000000000000000001100010100000100010;
												assign node1170 = (inp[12]) ? node1180 : node1171;
													assign node1171 = (inp[10]) ? node1175 : node1172;
														assign node1172 = (inp[8]) ? 46'b0000000000000110000000000000000010100000100000 : 46'b0000000000000100000000000000000010100000100000;
														assign node1175 = (inp[8]) ? node1177 : 46'b0000000000000110000000000000000010100000100000;
															assign node1177 = (inp[4]) ? 46'b0000000000000010000000000000000010100000100000 : 46'b0000000000000010000000000001000010100000100010;
													assign node1180 = (inp[10]) ? 46'b0000000000000010000000000001000000100000100010 : node1181;
														assign node1181 = (inp[4]) ? 46'b0000000000000010001000000001000000100000100000 : 46'b0000000000000110000000000000000000100000100000;
											assign node1185 = (inp[12]) ? node1199 : node1186;
												assign node1186 = (inp[7]) ? node1194 : node1187;
													assign node1187 = (inp[14]) ? node1191 : node1188;
														assign node1188 = (inp[10]) ? 46'b0000000000000110000000000000100010000000100000 : 46'b0000000000000100001000000001100010000000100000;
														assign node1191 = (inp[8]) ? 46'b0000000000000010000000000001100010000000100010 : 46'b0000000000000000001000000001100010000000100010;
													assign node1194 = (inp[14]) ? 46'b0000000000000010001000000001000010000000100000 : node1195;
														assign node1195 = (inp[4]) ? 46'b0000000000000000001000000001000010000000100010 : 46'b0000000000000000000000000001000010000000100010;
												assign node1199 = (inp[4]) ? node1209 : node1200;
													assign node1200 = (inp[10]) ? node1206 : node1201;
														assign node1201 = (inp[8]) ? 46'b0000000000000110000000000000000000000000100000 : node1202;
															assign node1202 = (inp[14]) ? 46'b0000000000000100001000000001000000000000100000 : 46'b0000000000000100000000000000000000000000100000;
														assign node1206 = (inp[7]) ? 46'b0000000000000100000000000001000000000000100010 : 46'b0000000000000100000000000001100000000000100010;
													assign node1209 = (inp[7]) ? node1213 : node1210;
														assign node1210 = (inp[8]) ? 46'b0000000000000000001000000001100000000000100010 : 46'b0000000000000100001000000001100000000000100000;
														assign node1213 = (inp[14]) ? node1215 : 46'b0000000000000000001000000001000000000000100010;
															assign node1215 = (inp[10]) ? 46'b0000000000000010001000000001000000000000100000 : 46'b0000000000000000001000000001000000000000100000;
							assign node1218 = (inp[9]) ? node1258 : node1219;
								assign node1219 = (inp[0]) ? node1239 : node1220;
									assign node1220 = (inp[6]) ? node1230 : node1221;
										assign node1221 = (inp[12]) ? node1223 : 46'b0000000000000000000000000000000000000000000000;
											assign node1223 = (inp[7]) ? node1227 : node1224;
												assign node1224 = (inp[5]) ? 46'b0000000000100000001000000001100000100000100000 : 46'b0001000000100000001000000001100000100000100000;
												assign node1227 = (inp[5]) ? 46'b0000000000100000001000000001000000100000100000 : 46'b0001000000100000001000000001000000100000100000;
										assign node1230 = (inp[12]) ? 46'b0000000000000000000000000000000000000000000000 : node1231;
											assign node1231 = (inp[5]) ? node1235 : node1232;
												assign node1232 = (inp[7]) ? 46'b0001000000100010000000000000000010000000100000 : 46'b0001000000100010000000000000100010000000100000;
												assign node1235 = (inp[7]) ? 46'b0000000000100010000000000000000010000000100000 : 46'b0000000000100010000000000000100010000000100000;
									assign node1239 = (inp[7]) ? node1249 : node1240;
										assign node1240 = (inp[5]) ? node1242 : 46'b0000000000000000000000000000000000000000000000;
											assign node1242 = (inp[6]) ? node1246 : node1243;
												assign node1243 = (inp[12]) ? 46'b0000000010000000000000000001100000100000000010 : 46'b0000000010000000000000000001100010100000000010;
												assign node1246 = (inp[12]) ? 46'b0000000010000000000000000001100000000000000010 : 46'b0000000010000000000000000001100010000000000010;
										assign node1249 = (inp[5]) ? 46'b0000000000000000000000000000000000000000000000 : node1250;
											assign node1250 = (inp[6]) ? node1254 : node1251;
												assign node1251 = (inp[12]) ? 46'b0001000010000100000000000000000000100000000000 : 46'b0001000010000100000000000000000010100000000000;
												assign node1254 = (inp[12]) ? 46'b0001000010000100000000000000000000000000000000 : 46'b0001000010000100000000000000000010000000000000;
								assign node1258 = (inp[0]) ? 46'b0000000000000000000000000000000000000000000000 : node1259;
									assign node1259 = (inp[7]) ? node1269 : node1260;
										assign node1260 = (inp[5]) ? node1262 : 46'b0000000000000000000000000000000000000000000000;
											assign node1262 = (inp[12]) ? node1266 : node1263;
												assign node1263 = (inp[6]) ? 46'b0000000010000000000000000001100010000001000010 : 46'b0000000010000000000000000001100010100001000010;
												assign node1266 = (inp[6]) ? 46'b0000000010000000000000000001100000000001000010 : 46'b0000000010000000000000000001100000100001000010;
										assign node1269 = (inp[5]) ? 46'b0000000000000000000000000000000000000000000000 : node1270;
											assign node1270 = (inp[12]) ? node1274 : node1271;
												assign node1271 = (inp[6]) ? 46'b0001000010000100000000000000000010000001000000 : 46'b0001000010000100000000000000000010100001000000;
												assign node1274 = (inp[6]) ? 46'b0001000010000100000000000000000000000001000000 : 46'b0001000010000100000000000000000000100001000000;

endmodule