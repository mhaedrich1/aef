module dtc_split875_bm66 (
	input  wire [16-1:0] inp,
	output wire [4-1:0] outp
);

	wire [4-1:0] node1;
	wire [4-1:0] node2;
	wire [4-1:0] node3;
	wire [4-1:0] node4;
	wire [4-1:0] node6;
	wire [4-1:0] node7;
	wire [4-1:0] node9;
	wire [4-1:0] node11;
	wire [4-1:0] node13;
	wire [4-1:0] node14;
	wire [4-1:0] node16;
	wire [4-1:0] node18;
	wire [4-1:0] node20;
	wire [4-1:0] node23;
	wire [4-1:0] node24;
	wire [4-1:0] node26;
	wire [4-1:0] node28;
	wire [4-1:0] node32;
	wire [4-1:0] node33;
	wire [4-1:0] node34;
	wire [4-1:0] node36;
	wire [4-1:0] node37;
	wire [4-1:0] node39;
	wire [4-1:0] node41;
	wire [4-1:0] node43;
	wire [4-1:0] node47;
	wire [4-1:0] node48;
	wire [4-1:0] node49;
	wire [4-1:0] node50;
	wire [4-1:0] node52;
	wire [4-1:0] node54;
	wire [4-1:0] node61;
	wire [4-1:0] node62;
	wire [4-1:0] node64;
	wire [4-1:0] node66;
	wire [4-1:0] node68;
	wire [4-1:0] node70;
	wire [4-1:0] node73;
	wire [4-1:0] node74;
	wire [4-1:0] node76;
	wire [4-1:0] node78;
	wire [4-1:0] node80;
	wire [4-1:0] node81;
	wire [4-1:0] node83;
	wire [4-1:0] node87;
	wire [4-1:0] node88;
	wire [4-1:0] node89;
	wire [4-1:0] node90;
	wire [4-1:0] node92;
	wire [4-1:0] node94;
	wire [4-1:0] node100;
	wire [4-1:0] node101;
	wire [4-1:0] node102;
	wire [4-1:0] node104;
	wire [4-1:0] node106;
	wire [4-1:0] node107;
	wire [4-1:0] node109;
	wire [4-1:0] node110;
	wire [4-1:0] node112;
	wire [4-1:0] node114;
	wire [4-1:0] node116;
	wire [4-1:0] node120;
	wire [4-1:0] node121;
	wire [4-1:0] node122;
	wire [4-1:0] node123;
	wire [4-1:0] node125;
	wire [4-1:0] node127;
	wire [4-1:0] node133;
	wire [4-1:0] node134;
	wire [4-1:0] node135;
	wire [4-1:0] node137;
	wire [4-1:0] node138;
	wire [4-1:0] node140;
	wire [4-1:0] node142;
	wire [4-1:0] node144;
	wire [4-1:0] node146;
	wire [4-1:0] node150;
	wire [4-1:0] node151;
	wire [4-1:0] node152;
	wire [4-1:0] node154;
	wire [4-1:0] node155;
	wire [4-1:0] node157;
	wire [4-1:0] node159;
	wire [4-1:0] node166;
	wire [4-1:0] node167;
	wire [4-1:0] node169;
	wire [4-1:0] node171;
	wire [4-1:0] node172;
	wire [4-1:0] node173;
	wire [4-1:0] node175;
	wire [4-1:0] node177;
	wire [4-1:0] node182;
	wire [4-1:0] node183;
	wire [4-1:0] node184;
	wire [4-1:0] node185;
	wire [4-1:0] node187;
	wire [4-1:0] node189;
	wire [4-1:0] node191;
	wire [4-1:0] node196;
	wire [4-1:0] node198;
	wire [4-1:0] node200;
	wire [4-1:0] node201;
	wire [4-1:0] node203;
	wire [4-1:0] node205;
	wire [4-1:0] node207;
	wire [4-1:0] node209;
	wire [4-1:0] node213;
	wire [4-1:0] node214;
	wire [4-1:0] node215;
	wire [4-1:0] node216;
	wire [4-1:0] node217;
	wire [4-1:0] node218;
	wire [4-1:0] node220;
	wire [4-1:0] node221;
	wire [4-1:0] node222;
	wire [4-1:0] node224;
	wire [4-1:0] node226;
	wire [4-1:0] node228;
	wire [4-1:0] node233;
	wire [4-1:0] node234;
	wire [4-1:0] node235;
	wire [4-1:0] node237;
	wire [4-1:0] node239;
	wire [4-1:0] node244;
	wire [4-1:0] node245;
	wire [4-1:0] node247;
	wire [4-1:0] node249;
	wire [4-1:0] node252;
	wire [4-1:0] node253;
	wire [4-1:0] node254;
	wire [4-1:0] node256;
	wire [4-1:0] node257;
	wire [4-1:0] node259;
	wire [4-1:0] node261;
	wire [4-1:0] node267;
	wire [4-1:0] node268;
	wire [4-1:0] node270;
	wire [4-1:0] node272;
	wire [4-1:0] node274;
	wire [4-1:0] node276;
	wire [4-1:0] node278;
	wire [4-1:0] node281;
	wire [4-1:0] node282;
	wire [4-1:0] node286;
	wire [4-1:0] node287;
	wire [4-1:0] node288;
	wire [4-1:0] node289;
	wire [4-1:0] node291;
	wire [4-1:0] node293;
	wire [4-1:0] node294;
	wire [4-1:0] node296;
	wire [4-1:0] node298;
	wire [4-1:0] node300;
	wire [4-1:0] node305;
	wire [4-1:0] node306;
	wire [4-1:0] node308;
	wire [4-1:0] node309;
	wire [4-1:0] node311;
	wire [4-1:0] node313;
	wire [4-1:0] node315;
	wire [4-1:0] node317;
	wire [4-1:0] node322;
	wire [4-1:0] node323;
	wire [4-1:0] node324;
	wire [4-1:0] node325;
	wire [4-1:0] node326;
	wire [4-1:0] node328;
	wire [4-1:0] node330;
	wire [4-1:0] node335;
	wire [4-1:0] node337;
	wire [4-1:0] node338;
	wire [4-1:0] node339;
	wire [4-1:0] node340;
	wire [4-1:0] node342;
	wire [4-1:0] node344;
	wire [4-1:0] node350;
	wire [4-1:0] node352;
	wire [4-1:0] node353;
	wire [4-1:0] node354;
	wire [4-1:0] node356;
	wire [4-1:0] node358;
	wire [4-1:0] node360;
	wire [4-1:0] node362;
	wire [4-1:0] node367;
	wire [4-1:0] node368;
	wire [4-1:0] node369;
	wire [4-1:0] node370;
	wire [4-1:0] node371;
	wire [4-1:0] node372;
	wire [4-1:0] node374;
	wire [4-1:0] node376;
	wire [4-1:0] node378;
	wire [4-1:0] node382;
	wire [4-1:0] node384;
	wire [4-1:0] node385;
	wire [4-1:0] node387;
	wire [4-1:0] node388;
	wire [4-1:0] node390;
	wire [4-1:0] node392;
	wire [4-1:0] node397;
	wire [4-1:0] node398;
	wire [4-1:0] node400;
	wire [4-1:0] node401;
	wire [4-1:0] node402;
	wire [4-1:0] node404;
	wire [4-1:0] node406;
	wire [4-1:0] node408;
	wire [4-1:0] node413;
	wire [4-1:0] node415;
	wire [4-1:0] node416;
	wire [4-1:0] node418;
	wire [4-1:0] node420;
	wire [4-1:0] node424;
	wire [4-1:0] node425;
	wire [4-1:0] node426;
	wire [4-1:0] node428;
	wire [4-1:0] node430;
	wire [4-1:0] node433;
	wire [4-1:0] node435;
	wire [4-1:0] node437;
	wire [4-1:0] node438;
	wire [4-1:0] node439;
	wire [4-1:0] node441;
	wire [4-1:0] node443;
	wire [4-1:0] node448;
	wire [4-1:0] node450;
	wire [4-1:0] node452;
	wire [4-1:0] node454;
	wire [4-1:0] node457;
	wire [4-1:0] node458;
	wire [4-1:0] node459;
	wire [4-1:0] node460;
	wire [4-1:0] node461;
	wire [4-1:0] node462;
	wire [4-1:0] node463;
	wire [4-1:0] node464;
	wire [4-1:0] node466;
	wire [4-1:0] node468;
	wire [4-1:0] node474;
	wire [4-1:0] node476;
	wire [4-1:0] node477;
	wire [4-1:0] node479;
	wire [4-1:0] node481;
	wire [4-1:0] node483;
	wire [4-1:0] node488;
	wire [4-1:0] node490;
	wire [4-1:0] node492;
	wire [4-1:0] node494;
	wire [4-1:0] node495;
	wire [4-1:0] node496;
	wire [4-1:0] node498;
	wire [4-1:0] node500;
	wire [4-1:0] node504;
	wire [4-1:0] node506;
	wire [4-1:0] node508;
	wire [4-1:0] node510;
	wire [4-1:0] node513;
	wire [4-1:0] node514;
	wire [4-1:0] node515;
	wire [4-1:0] node516;
	wire [4-1:0] node517;
	wire [4-1:0] node519;
	wire [4-1:0] node521;
	wire [4-1:0] node526;
	wire [4-1:0] node529;
	wire [4-1:0] node531;
	wire [4-1:0] node533;
	wire [4-1:0] node534;
	wire [4-1:0] node536;
	wire [4-1:0] node538;
	wire [4-1:0] node542;
	wire [4-1:0] node543;
	wire [4-1:0] node544;
	wire [4-1:0] node545;
	wire [4-1:0] node546;
	wire [4-1:0] node547;
	wire [4-1:0] node548;
	wire [4-1:0] node550;
	wire [4-1:0] node552;
	wire [4-1:0] node553;
	wire [4-1:0] node554;
	wire [4-1:0] node556;
	wire [4-1:0] node558;
	wire [4-1:0] node564;
	wire [4-1:0] node565;
	wire [4-1:0] node567;
	wire [4-1:0] node569;
	wire [4-1:0] node570;
	wire [4-1:0] node572;
	wire [4-1:0] node576;
	wire [4-1:0] node578;
	wire [4-1:0] node580;
	wire [4-1:0] node583;
	wire [4-1:0] node584;
	wire [4-1:0] node586;
	wire [4-1:0] node587;
	wire [4-1:0] node588;
	wire [4-1:0] node590;
	wire [4-1:0] node591;
	wire [4-1:0] node593;
	wire [4-1:0] node595;
	wire [4-1:0] node601;
	wire [4-1:0] node603;
	wire [4-1:0] node604;
	wire [4-1:0] node606;
	wire [4-1:0] node608;
	wire [4-1:0] node609;
	wire [4-1:0] node611;
	wire [4-1:0] node613;
	wire [4-1:0] node618;
	wire [4-1:0] node619;
	wire [4-1:0] node620;
	wire [4-1:0] node621;
	wire [4-1:0] node623;
	wire [4-1:0] node625;
	wire [4-1:0] node628;
	wire [4-1:0] node630;
	wire [4-1:0] node632;
	wire [4-1:0] node634;
	wire [4-1:0] node636;
	wire [4-1:0] node640;
	wire [4-1:0] node641;
	wire [4-1:0] node642;
	wire [4-1:0] node644;
	wire [4-1:0] node646;
	wire [4-1:0] node648;
	wire [4-1:0] node650;
	wire [4-1:0] node652;
	wire [4-1:0] node654;
	wire [4-1:0] node657;
	wire [4-1:0] node658;
	wire [4-1:0] node659;
	wire [4-1:0] node660;
	wire [4-1:0] node661;
	wire [4-1:0] node663;
	wire [4-1:0] node665;
	wire [4-1:0] node673;
	wire [4-1:0] node674;
	wire [4-1:0] node675;
	wire [4-1:0] node676;
	wire [4-1:0] node677;
	wire [4-1:0] node678;
	wire [4-1:0] node679;
	wire [4-1:0] node683;
	wire [4-1:0] node685;
	wire [4-1:0] node687;
	wire [4-1:0] node689;
	wire [4-1:0] node691;
	wire [4-1:0] node693;
	wire [4-1:0] node696;
	wire [4-1:0] node697;
	wire [4-1:0] node698;
	wire [4-1:0] node699;
	wire [4-1:0] node701;
	wire [4-1:0] node706;
	wire [4-1:0] node708;
	wire [4-1:0] node711;
	wire [4-1:0] node713;
	wire [4-1:0] node716;
	wire [4-1:0] node717;
	wire [4-1:0] node719;
	wire [4-1:0] node720;
	wire [4-1:0] node721;
	wire [4-1:0] node722;
	wire [4-1:0] node724;
	wire [4-1:0] node726;
	wire [4-1:0] node728;
	wire [4-1:0] node734;
	wire [4-1:0] node735;
	wire [4-1:0] node737;
	wire [4-1:0] node738;
	wire [4-1:0] node740;
	wire [4-1:0] node742;
	wire [4-1:0] node747;
	wire [4-1:0] node748;
	wire [4-1:0] node749;
	wire [4-1:0] node751;
	wire [4-1:0] node752;
	wire [4-1:0] node754;
	wire [4-1:0] node756;
	wire [4-1:0] node758;
	wire [4-1:0] node760;
	wire [4-1:0] node762;
	wire [4-1:0] node766;
	wire [4-1:0] node767;
	wire [4-1:0] node769;
	wire [4-1:0] node771;
	wire [4-1:0] node773;
	wire [4-1:0] node775;
	wire [4-1:0] node779;
	wire [4-1:0] node780;
	wire [4-1:0] node781;
	wire [4-1:0] node782;
	wire [4-1:0] node784;
	wire [4-1:0] node786;
	wire [4-1:0] node787;
	wire [4-1:0] node789;
	wire [4-1:0] node791;
	wire [4-1:0] node796;
	wire [4-1:0] node798;
	wire [4-1:0] node800;
	wire [4-1:0] node803;
	wire [4-1:0] node805;
	wire [4-1:0] node806;
	wire [4-1:0] node808;
	wire [4-1:0] node809;
	wire [4-1:0] node810;
	wire [4-1:0] node812;
	wire [4-1:0] node814;
	wire [4-1:0] node820;
	wire [4-1:0] node821;
	wire [4-1:0] node822;
	wire [4-1:0] node823;
	wire [4-1:0] node824;
	wire [4-1:0] node826;
	wire [4-1:0] node828;
	wire [4-1:0] node830;
	wire [4-1:0] node831;
	wire [4-1:0] node833;
	wire [4-1:0] node835;
	wire [4-1:0] node837;
	wire [4-1:0] node840;
	wire [4-1:0] node841;
	wire [4-1:0] node843;
	wire [4-1:0] node845;
	wire [4-1:0] node849;
	wire [4-1:0] node850;
	wire [4-1:0] node851;
	wire [4-1:0] node853;
	wire [4-1:0] node854;
	wire [4-1:0] node856;
	wire [4-1:0] node858;
	wire [4-1:0] node860;
	wire [4-1:0] node864;
	wire [4-1:0] node865;
	wire [4-1:0] node866;
	wire [4-1:0] node867;
	wire [4-1:0] node869;
	wire [4-1:0] node871;
	wire [4-1:0] node877;
	wire [4-1:0] node879;
	wire [4-1:0] node881;
	wire [4-1:0] node884;
	wire [4-1:0] node885;
	wire [4-1:0] node887;
	wire [4-1:0] node889;
	wire [4-1:0] node891;
	wire [4-1:0] node892;
	wire [4-1:0] node894;
	wire [4-1:0] node898;
	wire [4-1:0] node899;
	wire [4-1:0] node900;
	wire [4-1:0] node901;
	wire [4-1:0] node903;
	wire [4-1:0] node905;
	wire [4-1:0] node910;
	wire [4-1:0] node912;
	wire [4-1:0] node913;
	wire [4-1:0] node915;
	wire [4-1:0] node916;
	wire [4-1:0] node918;
	wire [4-1:0] node920;
	wire [4-1:0] node925;
	wire [4-1:0] node926;
	wire [4-1:0] node927;
	wire [4-1:0] node928;
	wire [4-1:0] node930;
	wire [4-1:0] node932;
	wire [4-1:0] node934;
	wire [4-1:0] node936;
	wire [4-1:0] node939;
	wire [4-1:0] node941;
	wire [4-1:0] node942;
	wire [4-1:0] node943;
	wire [4-1:0] node944;
	wire [4-1:0] node946;
	wire [4-1:0] node948;
	wire [4-1:0] node954;
	wire [4-1:0] node955;
	wire [4-1:0] node956;
	wire [4-1:0] node958;
	wire [4-1:0] node960;
	wire [4-1:0] node962;
	wire [4-1:0] node964;
	wire [4-1:0] node966;
	wire [4-1:0] node970;
	wire [4-1:0] node971;
	wire [4-1:0] node972;
	wire [4-1:0] node974;
	wire [4-1:0] node976;
	wire [4-1:0] node981;
	wire [4-1:0] node982;
	wire [4-1:0] node983;
	wire [4-1:0] node985;
	wire [4-1:0] node986;
	wire [4-1:0] node987;
	wire [4-1:0] node989;
	wire [4-1:0] node991;
	wire [4-1:0] node993;
	wire [4-1:0] node998;
	wire [4-1:0] node1001;
	wire [4-1:0] node1002;
	wire [4-1:0] node1004;
	wire [4-1:0] node1006;
	wire [4-1:0] node1008;
	wire [4-1:0] node1010;
	wire [4-1:0] node1013;
	wire [4-1:0] node1014;
	wire [4-1:0] node1015;
	wire [4-1:0] node1017;
	wire [4-1:0] node1019;
	wire [4-1:0] node1021;
	wire [4-1:0] node1023;
	wire [4-1:0] node1028;
	wire [4-1:0] node1029;
	wire [4-1:0] node1030;
	wire [4-1:0] node1031;
	wire [4-1:0] node1032;
	wire [4-1:0] node1033;
	wire [4-1:0] node1034;
	wire [4-1:0] node1036;
	wire [4-1:0] node1038;
	wire [4-1:0] node1040;
	wire [4-1:0] node1042;
	wire [4-1:0] node1045;
	wire [4-1:0] node1046;
	wire [4-1:0] node1047;
	wire [4-1:0] node1049;
	wire [4-1:0] node1051;
	wire [4-1:0] node1057;
	wire [4-1:0] node1058;
	wire [4-1:0] node1060;
	wire [4-1:0] node1062;
	wire [4-1:0] node1064;
	wire [4-1:0] node1067;
	wire [4-1:0] node1068;
	wire [4-1:0] node1071;
	wire [4-1:0] node1074;
	wire [4-1:0] node1075;
	wire [4-1:0] node1077;
	wire [4-1:0] node1078;
	wire [4-1:0] node1079;
	wire [4-1:0] node1080;
	wire [4-1:0] node1082;
	wire [4-1:0] node1084;
	wire [4-1:0] node1090;
	wire [4-1:0] node1091;
	wire [4-1:0] node1093;
	wire [4-1:0] node1094;
	wire [4-1:0] node1095;
	wire [4-1:0] node1097;
	wire [4-1:0] node1099;
	wire [4-1:0] node1104;
	wire [4-1:0] node1106;
	wire [4-1:0] node1109;
	wire [4-1:0] node1110;
	wire [4-1:0] node1111;
	wire [4-1:0] node1112;
	wire [4-1:0] node1113;
	wire [4-1:0] node1115;
	wire [4-1:0] node1117;
	wire [4-1:0] node1122;
	wire [4-1:0] node1124;
	wire [4-1:0] node1126;
	wire [4-1:0] node1127;
	wire [4-1:0] node1128;
	wire [4-1:0] node1130;
	wire [4-1:0] node1132;
	wire [4-1:0] node1136;
	wire [4-1:0] node1138;
	wire [4-1:0] node1140;
	wire [4-1:0] node1142;
	wire [4-1:0] node1145;
	wire [4-1:0] node1146;
	wire [4-1:0] node1147;
	wire [4-1:0] node1149;
	wire [4-1:0] node1150;
	wire [4-1:0] node1152;
	wire [4-1:0] node1154;
	wire [4-1:0] node1156;
	wire [4-1:0] node1161;
	wire [4-1:0] node1162;
	wire [4-1:0] node1164;
	wire [4-1:0] node1166;
	wire [4-1:0] node1168;
	wire [4-1:0] node1172;
	wire [4-1:0] node1173;
	wire [4-1:0] node1174;
	wire [4-1:0] node1175;
	wire [4-1:0] node1177;
	wire [4-1:0] node1179;
	wire [4-1:0] node1180;
	wire [4-1:0] node1182;
	wire [4-1:0] node1184;
	wire [4-1:0] node1186;
	wire [4-1:0] node1189;
	wire [4-1:0] node1190;
	wire [4-1:0] node1192;
	wire [4-1:0] node1194;
	wire [4-1:0] node1198;
	wire [4-1:0] node1200;
	wire [4-1:0] node1202;
	wire [4-1:0] node1203;
	wire [4-1:0] node1205;
	wire [4-1:0] node1209;
	wire [4-1:0] node1210;
	wire [4-1:0] node1211;
	wire [4-1:0] node1212;
	wire [4-1:0] node1214;
	wire [4-1:0] node1215;
	wire [4-1:0] node1219;
	wire [4-1:0] node1220;
	wire [4-1:0] node1221;
	wire [4-1:0] node1222;
	wire [4-1:0] node1223;
	wire [4-1:0] node1224;
	wire [4-1:0] node1226;
	wire [4-1:0] node1229;
	wire [4-1:0] node1230;
	wire [4-1:0] node1234;
	wire [4-1:0] node1235;
	wire [4-1:0] node1237;
	wire [4-1:0] node1240;
	wire [4-1:0] node1243;
	wire [4-1:0] node1244;
	wire [4-1:0] node1245;
	wire [4-1:0] node1249;
	wire [4-1:0] node1251;
	wire [4-1:0] node1254;
	wire [4-1:0] node1255;
	wire [4-1:0] node1257;
	wire [4-1:0] node1260;
	wire [4-1:0] node1261;
	wire [4-1:0] node1265;
	wire [4-1:0] node1266;
	wire [4-1:0] node1268;
	wire [4-1:0] node1269;
	wire [4-1:0] node1273;
	wire [4-1:0] node1275;
	wire [4-1:0] node1278;
	wire [4-1:0] node1279;
	wire [4-1:0] node1282;
	wire [4-1:0] node1285;
	wire [4-1:0] node1286;
	wire [4-1:0] node1288;
	wire [4-1:0] node1289;
	wire [4-1:0] node1290;
	wire [4-1:0] node1292;
	wire [4-1:0] node1294;
	wire [4-1:0] node1298;
	wire [4-1:0] node1300;
	wire [4-1:0] node1302;
	wire [4-1:0] node1304;
	wire [4-1:0] node1307;
	wire [4-1:0] node1309;
	wire [4-1:0] node1311;
	wire [4-1:0] node1312;
	wire [4-1:0] node1316;
	wire [4-1:0] node1317;
	wire [4-1:0] node1318;
	wire [4-1:0] node1319;
	wire [4-1:0] node1321;
	wire [4-1:0] node1322;
	wire [4-1:0] node1324;
	wire [4-1:0] node1326;
	wire [4-1:0] node1328;
	wire [4-1:0] node1332;
	wire [4-1:0] node1333;
	wire [4-1:0] node1334;
	wire [4-1:0] node1335;
	wire [4-1:0] node1337;
	wire [4-1:0] node1339;
	wire [4-1:0] node1345;
	wire [4-1:0] node1346;
	wire [4-1:0] node1347;
	wire [4-1:0] node1349;
	wire [4-1:0] node1351;
	wire [4-1:0] node1355;
	wire [4-1:0] node1357;
	wire [4-1:0] node1358;
	wire [4-1:0] node1360;
	wire [4-1:0] node1362;
	wire [4-1:0] node1364;
	wire [4-1:0] node1368;
	wire [4-1:0] node1369;
	wire [4-1:0] node1370;
	wire [4-1:0] node1372;
	wire [4-1:0] node1373;
	wire [4-1:0] node1375;
	wire [4-1:0] node1377;
	wire [4-1:0] node1379;
	wire [4-1:0] node1382;
	wire [4-1:0] node1383;
	wire [4-1:0] node1385;
	wire [4-1:0] node1387;
	wire [4-1:0] node1391;
	wire [4-1:0] node1393;
	wire [4-1:0] node1394;
	wire [4-1:0] node1396;
	wire [4-1:0] node1400;
	wire [4-1:0] node1401;
	wire [4-1:0] node1402;
	wire [4-1:0] node1403;
	wire [4-1:0] node1404;
	wire [4-1:0] node1406;
	wire [4-1:0] node1408;
	wire [4-1:0] node1412;
	wire [4-1:0] node1414;
	wire [4-1:0] node1416;
	wire [4-1:0] node1418;
	wire [4-1:0] node1421;
	wire [4-1:0] node1423;
	wire [4-1:0] node1425;
	wire [4-1:0] node1428;
	wire [4-1:0] node1429;
	wire [4-1:0] node1430;
	wire [4-1:0] node1432;
	wire [4-1:0] node1434;
	wire [4-1:0] node1436;
	wire [4-1:0] node1439;
	wire [4-1:0] node1440;
	wire [4-1:0] node1442;
	wire [4-1:0] node1444;
	wire [4-1:0] node1448;
	wire [4-1:0] node1449;
	wire [4-1:0] node1451;
	wire [4-1:0] node1454;
	wire [4-1:0] node1455;
	wire [4-1:0] node1457;
	wire [4-1:0] node1459;
	wire [4-1:0] node1462;
	wire [4-1:0] node1464;
	wire [4-1:0] node1466;

	assign outp = (inp[10]) ? node542 : node1;
		assign node1 = (inp[5]) ? node213 : node2;
			assign node2 = (inp[4]) ? node100 : node3;
				assign node3 = (inp[14]) ? node61 : node4;
					assign node4 = (inp[13]) ? node6 : 4'b1111;
						assign node6 = (inp[12]) ? node32 : node7;
							assign node7 = (inp[9]) ? node9 : 4'b1111;
								assign node9 = (inp[8]) ? node11 : 4'b1111;
									assign node11 = (inp[2]) ? node13 : 4'b1111;
										assign node13 = (inp[6]) ? node23 : node14;
											assign node14 = (inp[11]) ? node16 : 4'b1111;
												assign node16 = (inp[7]) ? node18 : 4'b1111;
													assign node18 = (inp[1]) ? node20 : 4'b1111;
														assign node20 = (inp[15]) ? 4'b1101 : 4'b1111;
											assign node23 = (inp[7]) ? 4'b1101 : node24;
												assign node24 = (inp[11]) ? node26 : 4'b1111;
													assign node26 = (inp[1]) ? node28 : 4'b1111;
														assign node28 = (inp[15]) ? 4'b1101 : 4'b1111;
							assign node32 = (inp[2]) ? 4'b1101 : node33;
								assign node33 = (inp[6]) ? node47 : node34;
									assign node34 = (inp[9]) ? node36 : 4'b1111;
										assign node36 = (inp[8]) ? 4'b1101 : node37;
											assign node37 = (inp[1]) ? node39 : 4'b1111;
												assign node39 = (inp[15]) ? node41 : 4'b1111;
													assign node41 = (inp[7]) ? node43 : 4'b1111;
														assign node43 = (inp[11]) ? 4'b1101 : 4'b1111;
									assign node47 = (inp[9]) ? 4'b1101 : node48;
										assign node48 = (inp[7]) ? 4'b1101 : node49;
											assign node49 = (inp[8]) ? 4'b1101 : node50;
												assign node50 = (inp[11]) ? node52 : 4'b1111;
													assign node52 = (inp[15]) ? node54 : 4'b1111;
														assign node54 = (inp[1]) ? 4'b1101 : 4'b1111;
					assign node61 = (inp[13]) ? node73 : node62;
						assign node62 = (inp[6]) ? node64 : 4'b1101;
							assign node64 = (inp[12]) ? node66 : 4'b1101;
								assign node66 = (inp[8]) ? node68 : 4'b1101;
									assign node68 = (inp[9]) ? node70 : 4'b1101;
										assign node70 = (inp[2]) ? 4'b1011 : 4'b1101;
						assign node73 = (inp[12]) ? node87 : node74;
							assign node74 = (inp[2]) ? node76 : 4'b1101;
								assign node76 = (inp[8]) ? node78 : 4'b1101;
									assign node78 = (inp[9]) ? node80 : 4'b1101;
										assign node80 = (inp[6]) ? 4'b1011 : node81;
											assign node81 = (inp[15]) ? node83 : 4'b1101;
												assign node83 = (inp[7]) ? 4'b1111 : 4'b1101;
							assign node87 = (inp[6]) ? 4'b1011 : node88;
								assign node88 = (inp[9]) ? 4'b1111 : node89;
									assign node89 = (inp[2]) ? 4'b1111 : node90;
										assign node90 = (inp[15]) ? node92 : 4'b1101;
											assign node92 = (inp[7]) ? node94 : 4'b1101;
												assign node94 = (inp[8]) ? 4'b1111 : 4'b1101;
				assign node100 = (inp[14]) ? node166 : node101;
					assign node101 = (inp[12]) ? node133 : node102;
						assign node102 = (inp[13]) ? node104 : 4'b1011;
							assign node104 = (inp[2]) ? node106 : 4'b1011;
								assign node106 = (inp[9]) ? node120 : node107;
									assign node107 = (inp[6]) ? node109 : 4'b1011;
										assign node109 = (inp[8]) ? 4'b1001 : node110;
											assign node110 = (inp[11]) ? node112 : 4'b1011;
												assign node112 = (inp[7]) ? node114 : 4'b1011;
													assign node114 = (inp[1]) ? node116 : 4'b1011;
														assign node116 = (inp[15]) ? 4'b1001 : 4'b1011;
									assign node120 = (inp[7]) ? 4'b1001 : node121;
										assign node121 = (inp[6]) ? 4'b1001 : node122;
											assign node122 = (inp[8]) ? 4'b1001 : node123;
												assign node123 = (inp[11]) ? node125 : 4'b1011;
													assign node125 = (inp[1]) ? node127 : 4'b1011;
														assign node127 = (inp[15]) ? 4'b1001 : 4'b1011;
						assign node133 = (inp[13]) ? 4'b1001 : node134;
							assign node134 = (inp[2]) ? node150 : node135;
								assign node135 = (inp[6]) ? node137 : 4'b1011;
									assign node137 = (inp[9]) ? 4'b1001 : node138;
										assign node138 = (inp[15]) ? node140 : 4'b1011;
											assign node140 = (inp[1]) ? node142 : 4'b1011;
												assign node142 = (inp[8]) ? node144 : 4'b1011;
													assign node144 = (inp[11]) ? node146 : 4'b1011;
														assign node146 = (inp[7]) ? 4'b1001 : 4'b1011;
								assign node150 = (inp[9]) ? 4'b1001 : node151;
									assign node151 = (inp[6]) ? 4'b1001 : node152;
										assign node152 = (inp[8]) ? node154 : 4'b1011;
											assign node154 = (inp[7]) ? 4'b1001 : node155;
												assign node155 = (inp[11]) ? node157 : 4'b1011;
													assign node157 = (inp[15]) ? node159 : 4'b1011;
														assign node159 = (inp[1]) ? 4'b1001 : 4'b1011;
					assign node166 = (inp[12]) ? node182 : node167;
						assign node167 = (inp[13]) ? node169 : 4'b1001;
							assign node169 = (inp[2]) ? node171 : 4'b1001;
								assign node171 = (inp[6]) ? 4'b1111 : node172;
									assign node172 = (inp[9]) ? 4'b1011 : node173;
										assign node173 = (inp[8]) ? node175 : 4'b1001;
											assign node175 = (inp[7]) ? node177 : 4'b1001;
												assign node177 = (inp[15]) ? 4'b1011 : 4'b1001;
						assign node182 = (inp[6]) ? node196 : node183;
							assign node183 = (inp[13]) ? 4'b1011 : node184;
								assign node184 = (inp[2]) ? 4'b1011 : node185;
									assign node185 = (inp[8]) ? node187 : 4'b1001;
										assign node187 = (inp[15]) ? node189 : 4'b1001;
											assign node189 = (inp[9]) ? node191 : 4'b1001;
												assign node191 = (inp[7]) ? 4'b1011 : 4'b1001;
							assign node196 = (inp[13]) ? node198 : 4'b1110;
								assign node198 = (inp[2]) ? node200 : 4'b1110;
									assign node200 = (inp[9]) ? 4'b1100 : node201;
										assign node201 = (inp[11]) ? node203 : 4'b1110;
											assign node203 = (inp[7]) ? node205 : 4'b1110;
												assign node205 = (inp[8]) ? node207 : 4'b1110;
													assign node207 = (inp[1]) ? node209 : 4'b1110;
														assign node209 = (inp[15]) ? 4'b1100 : 4'b1110;
			assign node213 = (inp[12]) ? node367 : node214;
				assign node214 = (inp[6]) ? node286 : node215;
					assign node215 = (inp[13]) ? node267 : node216;
						assign node216 = (inp[4]) ? node244 : node217;
							assign node217 = (inp[2]) ? node233 : node218;
								assign node218 = (inp[14]) ? node220 : 4'b1001;
									assign node220 = (inp[9]) ? 4'b1001 : node221;
										assign node221 = (inp[8]) ? 4'b1001 : node222;
											assign node222 = (inp[7]) ? node224 : 4'b1011;
												assign node224 = (inp[11]) ? node226 : 4'b1011;
													assign node226 = (inp[15]) ? node228 : 4'b1011;
														assign node228 = (inp[1]) ? 4'b1001 : 4'b1011;
								assign node233 = (inp[14]) ? 4'b1001 : node234;
									assign node234 = (inp[9]) ? 4'b1011 : node235;
										assign node235 = (inp[15]) ? node237 : 4'b1001;
											assign node237 = (inp[7]) ? node239 : 4'b1001;
												assign node239 = (inp[8]) ? 4'b1011 : 4'b1001;
							assign node244 = (inp[14]) ? node252 : node245;
								assign node245 = (inp[9]) ? node247 : 4'b1101;
									assign node247 = (inp[8]) ? node249 : 4'b1101;
										assign node249 = (inp[2]) ? 4'b1011 : 4'b1101;
								assign node252 = (inp[9]) ? 4'b1001 : node253;
									assign node253 = (inp[2]) ? 4'b1001 : node254;
										assign node254 = (inp[8]) ? node256 : 4'b1011;
											assign node256 = (inp[7]) ? 4'b1001 : node257;
												assign node257 = (inp[15]) ? node259 : 4'b1011;
													assign node259 = (inp[11]) ? node261 : 4'b1011;
														assign node261 = (inp[1]) ? 4'b1001 : 4'b1011;
						assign node267 = (inp[2]) ? node281 : node268;
							assign node268 = (inp[14]) ? node270 : 4'b1011;
								assign node270 = (inp[9]) ? node272 : 4'b1001;
									assign node272 = (inp[15]) ? node274 : 4'b1001;
										assign node274 = (inp[4]) ? node276 : 4'b1001;
											assign node276 = (inp[7]) ? node278 : 4'b1001;
												assign node278 = (inp[8]) ? 4'b1011 : 4'b1001;
							assign node281 = (inp[4]) ? 4'b1011 : node282;
								assign node282 = (inp[14]) ? 4'b1111 : 4'b1011;
					assign node286 = (inp[14]) ? node322 : node287;
						assign node287 = (inp[4]) ? node305 : node288;
							assign node288 = (inp[13]) ? 4'b1101 : node289;
								assign node289 = (inp[9]) ? node291 : 4'b1111;
									assign node291 = (inp[2]) ? node293 : 4'b1111;
										assign node293 = (inp[8]) ? 4'b1101 : node294;
											assign node294 = (inp[15]) ? node296 : 4'b1111;
												assign node296 = (inp[7]) ? node298 : 4'b1111;
													assign node298 = (inp[11]) ? node300 : 4'b1111;
														assign node300 = (inp[1]) ? 4'b1101 : 4'b1111;
							assign node305 = (inp[13]) ? 4'b1001 : node306;
								assign node306 = (inp[2]) ? node308 : 4'b1011;
									assign node308 = (inp[9]) ? 4'b1001 : node309;
										assign node309 = (inp[11]) ? node311 : 4'b1011;
											assign node311 = (inp[8]) ? node313 : 4'b1011;
												assign node313 = (inp[7]) ? node315 : 4'b1011;
													assign node315 = (inp[1]) ? node317 : 4'b1011;
														assign node317 = (inp[15]) ? 4'b1001 : 4'b1011;
						assign node322 = (inp[4]) ? node350 : node323;
							assign node323 = (inp[13]) ? node335 : node324;
								assign node324 = (inp[2]) ? 4'b1111 : node325;
									assign node325 = (inp[9]) ? 4'b1111 : node326;
										assign node326 = (inp[7]) ? node328 : 4'b1101;
											assign node328 = (inp[15]) ? node330 : 4'b1101;
												assign node330 = (inp[8]) ? 4'b1111 : 4'b1101;
								assign node335 = (inp[2]) ? node337 : 4'b1111;
									assign node337 = (inp[8]) ? 4'b1101 : node338;
										assign node338 = (inp[9]) ? 4'b1101 : node339;
											assign node339 = (inp[7]) ? 4'b1101 : node340;
												assign node340 = (inp[1]) ? node342 : 4'b1111;
													assign node342 = (inp[11]) ? node344 : 4'b1111;
														assign node344 = (inp[15]) ? 4'b1101 : 4'b1111;
							assign node350 = (inp[13]) ? node352 : 4'b1110;
								assign node352 = (inp[9]) ? 4'b1100 : node353;
									assign node353 = (inp[2]) ? 4'b1100 : node354;
										assign node354 = (inp[11]) ? node356 : 4'b1110;
											assign node356 = (inp[1]) ? node358 : 4'b1110;
												assign node358 = (inp[8]) ? node360 : 4'b1110;
													assign node360 = (inp[7]) ? node362 : 4'b1110;
														assign node362 = (inp[15]) ? 4'b1100 : 4'b1110;
				assign node367 = (inp[6]) ? node457 : node368;
					assign node368 = (inp[14]) ? node424 : node369;
						assign node369 = (inp[4]) ? node397 : node370;
							assign node370 = (inp[2]) ? node382 : node371;
								assign node371 = (inp[13]) ? 4'b1110 : node372;
									assign node372 = (inp[15]) ? node374 : 4'b1100;
										assign node374 = (inp[8]) ? node376 : 4'b1100;
											assign node376 = (inp[7]) ? node378 : 4'b1100;
												assign node378 = (inp[9]) ? 4'b1110 : 4'b1100;
								assign node382 = (inp[13]) ? node384 : 4'b1110;
									assign node384 = (inp[9]) ? 4'b1100 : node385;
										assign node385 = (inp[8]) ? node387 : 4'b1110;
											assign node387 = (inp[7]) ? 4'b1100 : node388;
												assign node388 = (inp[11]) ? node390 : 4'b1110;
													assign node390 = (inp[15]) ? node392 : 4'b1110;
														assign node392 = (inp[1]) ? 4'b1100 : 4'b1110;
							assign node397 = (inp[13]) ? node413 : node398;
								assign node398 = (inp[2]) ? node400 : 4'b1110;
									assign node400 = (inp[9]) ? 4'b1100 : node401;
										assign node401 = (inp[8]) ? 4'b1100 : node402;
											assign node402 = (inp[7]) ? node404 : 4'b1110;
												assign node404 = (inp[1]) ? node406 : 4'b1110;
													assign node406 = (inp[15]) ? node408 : 4'b1110;
														assign node408 = (inp[11]) ? 4'b1100 : 4'b1110;
								assign node413 = (inp[2]) ? node415 : 4'b1100;
									assign node415 = (inp[9]) ? 4'b1110 : node416;
										assign node416 = (inp[7]) ? node418 : 4'b1100;
											assign node418 = (inp[8]) ? node420 : 4'b1100;
												assign node420 = (inp[15]) ? 4'b1110 : 4'b1100;
						assign node424 = (inp[13]) ? node448 : node425;
							assign node425 = (inp[4]) ? node433 : node426;
								assign node426 = (inp[9]) ? node428 : 4'b1100;
									assign node428 = (inp[2]) ? node430 : 4'b1100;
										assign node430 = (inp[8]) ? 4'b1010 : 4'b1100;
								assign node433 = (inp[9]) ? node435 : 4'b1110;
									assign node435 = (inp[2]) ? node437 : 4'b1110;
										assign node437 = (inp[8]) ? 4'b1100 : node438;
											assign node438 = (inp[7]) ? 4'b1100 : node439;
												assign node439 = (inp[15]) ? node441 : 4'b1110;
													assign node441 = (inp[1]) ? node443 : 4'b1110;
														assign node443 = (inp[11]) ? 4'b1100 : 4'b1110;
							assign node448 = (inp[4]) ? node450 : 4'b1010;
								assign node450 = (inp[8]) ? node452 : 4'b1100;
									assign node452 = (inp[2]) ? node454 : 4'b1100;
										assign node454 = (inp[9]) ? 4'b1010 : 4'b1100;
					assign node457 = (inp[13]) ? node513 : node458;
						assign node458 = (inp[4]) ? node488 : node459;
							assign node459 = (inp[2]) ? 4'b1000 : node460;
								assign node460 = (inp[14]) ? node474 : node461;
									assign node461 = (inp[8]) ? 4'b1000 : node462;
										assign node462 = (inp[9]) ? 4'b1000 : node463;
											assign node463 = (inp[7]) ? 4'b1000 : node464;
												assign node464 = (inp[11]) ? node466 : 4'b1010;
													assign node466 = (inp[15]) ? node468 : 4'b1010;
														assign node468 = (inp[1]) ? 4'b1000 : 4'b1010;
									assign node474 = (inp[9]) ? node476 : 4'b1010;
										assign node476 = (inp[8]) ? 4'b1000 : node477;
											assign node477 = (inp[15]) ? node479 : 4'b1010;
												assign node479 = (inp[11]) ? node481 : 4'b1010;
													assign node481 = (inp[1]) ? node483 : 4'b1010;
														assign node483 = (inp[7]) ? 4'b1000 : 4'b1010;
							assign node488 = (inp[8]) ? node490 : 4'b1010;
								assign node490 = (inp[2]) ? node492 : 4'b1010;
									assign node492 = (inp[9]) ? node494 : 4'b1010;
										assign node494 = (inp[7]) ? node504 : node495;
											assign node495 = (inp[14]) ? 4'b1010 : node496;
												assign node496 = (inp[15]) ? node498 : 4'b1010;
													assign node498 = (inp[11]) ? node500 : 4'b1010;
														assign node500 = (inp[1]) ? 4'b1000 : 4'b1010;
											assign node504 = (inp[14]) ? node506 : 4'b1000;
												assign node506 = (inp[11]) ? node508 : 4'b1010;
													assign node508 = (inp[1]) ? node510 : 4'b1010;
														assign node510 = (inp[15]) ? 4'b1000 : 4'b1010;
						assign node513 = (inp[4]) ? node529 : node514;
							assign node514 = (inp[2]) ? node526 : node515;
								assign node515 = (inp[14]) ? 4'b1000 : node516;
									assign node516 = (inp[9]) ? 4'b1010 : node517;
										assign node517 = (inp[8]) ? node519 : 4'b1000;
											assign node519 = (inp[15]) ? node521 : 4'b1000;
												assign node521 = (inp[7]) ? 4'b1010 : 4'b1000;
								assign node526 = (inp[14]) ? 4'b1110 : 4'b1010;
							assign node529 = (inp[15]) ? node531 : 4'b1000;
								assign node531 = (inp[7]) ? node533 : 4'b1000;
									assign node533 = (inp[14]) ? 4'b1000 : node534;
										assign node534 = (inp[2]) ? node536 : 4'b1000;
											assign node536 = (inp[9]) ? node538 : 4'b1000;
												assign node538 = (inp[8]) ? 4'b1010 : 4'b1000;
		assign node542 = (inp[5]) ? node820 : node543;
			assign node543 = (inp[4]) ? node673 : node544;
				assign node544 = (inp[6]) ? node618 : node545;
					assign node545 = (inp[14]) ? node583 : node546;
						assign node546 = (inp[13]) ? node564 : node547;
							assign node547 = (inp[2]) ? 4'b1100 : node548;
								assign node548 = (inp[12]) ? node550 : 4'b1100;
									assign node550 = (inp[9]) ? node552 : 4'b1110;
										assign node552 = (inp[7]) ? 4'b1100 : node553;
											assign node553 = (inp[8]) ? 4'b1100 : node554;
												assign node554 = (inp[1]) ? node556 : 4'b1110;
													assign node556 = (inp[15]) ? node558 : 4'b1110;
														assign node558 = (inp[11]) ? 4'b1100 : 4'b1110;
							assign node564 = (inp[2]) ? node576 : node565;
								assign node565 = (inp[8]) ? node567 : 4'b1100;
									assign node567 = (inp[15]) ? node569 : 4'b1100;
										assign node569 = (inp[12]) ? 4'b1100 : node570;
											assign node570 = (inp[9]) ? node572 : 4'b1100;
												assign node572 = (inp[7]) ? 4'b1110 : 4'b1100;
								assign node576 = (inp[12]) ? node578 : 4'b1110;
									assign node578 = (inp[8]) ? node580 : 4'b1100;
										assign node580 = (inp[9]) ? 4'b1010 : 4'b1100;
						assign node583 = (inp[12]) ? node601 : node584;
							assign node584 = (inp[13]) ? node586 : 4'b1110;
								assign node586 = (inp[2]) ? 4'b1100 : node587;
									assign node587 = (inp[9]) ? 4'b1100 : node588;
										assign node588 = (inp[8]) ? node590 : 4'b1110;
											assign node590 = (inp[7]) ? 4'b1100 : node591;
												assign node591 = (inp[1]) ? node593 : 4'b1110;
													assign node593 = (inp[15]) ? node595 : 4'b1110;
														assign node595 = (inp[11]) ? 4'b1100 : 4'b1110;
							assign node601 = (inp[13]) ? node603 : 4'b1010;
								assign node603 = (inp[2]) ? 4'b1000 : node604;
									assign node604 = (inp[8]) ? node606 : 4'b1010;
										assign node606 = (inp[9]) ? node608 : 4'b1010;
											assign node608 = (inp[7]) ? 4'b1000 : node609;
												assign node609 = (inp[11]) ? node611 : 4'b1010;
													assign node611 = (inp[1]) ? node613 : 4'b1010;
														assign node613 = (inp[15]) ? 4'b1000 : 4'b1010;
					assign node618 = (inp[14]) ? node640 : node619;
						assign node619 = (inp[13]) ? 4'b1010 : node620;
							assign node620 = (inp[12]) ? node628 : node621;
								assign node621 = (inp[8]) ? node623 : 4'b1100;
									assign node623 = (inp[2]) ? node625 : 4'b1100;
										assign node625 = (inp[9]) ? 4'b1010 : 4'b1100;
								assign node628 = (inp[7]) ? node630 : 4'b1000;
									assign node630 = (inp[15]) ? node632 : 4'b1000;
										assign node632 = (inp[9]) ? node634 : 4'b1000;
											assign node634 = (inp[2]) ? node636 : 4'b1000;
												assign node636 = (inp[8]) ? 4'b1010 : 4'b1000;
						assign node640 = (inp[13]) ? 4'b1000 : node641;
							assign node641 = (inp[2]) ? node657 : node642;
								assign node642 = (inp[9]) ? node644 : 4'b1010;
									assign node644 = (inp[15]) ? node646 : 4'b1010;
										assign node646 = (inp[8]) ? node648 : 4'b1010;
											assign node648 = (inp[11]) ? node650 : 4'b1010;
												assign node650 = (inp[12]) ? node652 : 4'b1010;
													assign node652 = (inp[7]) ? node654 : 4'b1010;
														assign node654 = (inp[1]) ? 4'b1000 : 4'b1010;
								assign node657 = (inp[7]) ? 4'b1000 : node658;
									assign node658 = (inp[8]) ? 4'b1000 : node659;
										assign node659 = (inp[9]) ? 4'b1000 : node660;
											assign node660 = (inp[12]) ? 4'b1000 : node661;
												assign node661 = (inp[1]) ? node663 : 4'b1010;
													assign node663 = (inp[15]) ? node665 : 4'b1010;
														assign node665 = (inp[11]) ? 4'b1000 : 4'b1010;
				assign node673 = (inp[12]) ? node747 : node674;
					assign node674 = (inp[6]) ? node716 : node675;
						assign node675 = (inp[14]) ? node711 : node676;
							assign node676 = (inp[8]) ? node696 : node677;
								assign node677 = (inp[13]) ? node683 : node678;
									assign node678 = (inp[9]) ? 4'b1010 : node679;
										assign node679 = (inp[2]) ? 4'b1010 : 4'b1000;
									assign node683 = (inp[11]) ? node685 : 4'b1010;
										assign node685 = (inp[9]) ? node687 : 4'b1010;
											assign node687 = (inp[15]) ? node689 : 4'b1010;
												assign node689 = (inp[7]) ? node691 : 4'b1010;
													assign node691 = (inp[2]) ? node693 : 4'b1010;
														assign node693 = (inp[1]) ? 4'b1000 : 4'b1010;
								assign node696 = (inp[13]) ? node706 : node697;
									assign node697 = (inp[9]) ? 4'b1010 : node698;
										assign node698 = (inp[2]) ? 4'b1010 : node699;
											assign node699 = (inp[7]) ? node701 : 4'b1000;
												assign node701 = (inp[15]) ? 4'b1010 : 4'b1000;
									assign node706 = (inp[9]) ? node708 : 4'b1010;
										assign node708 = (inp[2]) ? 4'b1000 : 4'b1010;
							assign node711 = (inp[13]) ? node713 : 4'b1000;
								assign node713 = (inp[2]) ? 4'b1110 : 4'b1000;
						assign node716 = (inp[14]) ? node734 : node717;
							assign node717 = (inp[13]) ? node719 : 4'b1110;
								assign node719 = (inp[9]) ? 4'b1100 : node720;
									assign node720 = (inp[2]) ? 4'b1100 : node721;
										assign node721 = (inp[8]) ? 4'b1100 : node722;
											assign node722 = (inp[11]) ? node724 : 4'b1110;
												assign node724 = (inp[7]) ? node726 : 4'b1110;
													assign node726 = (inp[1]) ? node728 : 4'b1110;
														assign node728 = (inp[15]) ? 4'b1100 : 4'b1110;
							assign node734 = (inp[13]) ? 4'b1110 : node735;
								assign node735 = (inp[2]) ? node737 : 4'b1100;
									assign node737 = (inp[9]) ? 4'b1110 : node738;
										assign node738 = (inp[15]) ? node740 : 4'b1100;
											assign node740 = (inp[8]) ? node742 : 4'b1100;
												assign node742 = (inp[7]) ? 4'b1110 : 4'b1100;
					assign node747 = (inp[6]) ? node779 : node748;
						assign node748 = (inp[14]) ? node766 : node749;
							assign node749 = (inp[13]) ? node751 : 4'b1111;
								assign node751 = (inp[2]) ? 4'b1101 : node752;
									assign node752 = (inp[9]) ? node754 : 4'b1111;
										assign node754 = (inp[15]) ? node756 : 4'b1111;
											assign node756 = (inp[1]) ? node758 : 4'b1111;
												assign node758 = (inp[11]) ? node760 : 4'b1111;
													assign node760 = (inp[8]) ? node762 : 4'b1111;
														assign node762 = (inp[7]) ? 4'b1101 : 4'b1111;
							assign node766 = (inp[13]) ? 4'b1111 : node767;
								assign node767 = (inp[7]) ? node769 : 4'b1101;
									assign node769 = (inp[15]) ? node771 : 4'b1101;
										assign node771 = (inp[8]) ? node773 : 4'b1101;
											assign node773 = (inp[9]) ? node775 : 4'b1101;
												assign node775 = (inp[2]) ? 4'b1111 : 4'b1101;
						assign node779 = (inp[14]) ? node803 : node780;
							assign node780 = (inp[2]) ? node796 : node781;
								assign node781 = (inp[13]) ? 4'b1101 : node782;
									assign node782 = (inp[8]) ? node784 : 4'b1111;
										assign node784 = (inp[9]) ? node786 : 4'b1111;
											assign node786 = (inp[7]) ? 4'b1101 : node787;
												assign node787 = (inp[15]) ? node789 : 4'b1111;
													assign node789 = (inp[1]) ? node791 : 4'b1111;
														assign node791 = (inp[11]) ? 4'b1101 : 4'b1111;
								assign node796 = (inp[8]) ? node798 : 4'b1101;
									assign node798 = (inp[13]) ? node800 : 4'b1101;
										assign node800 = (inp[9]) ? 4'b1011 : 4'b1101;
							assign node803 = (inp[13]) ? node805 : 4'b1011;
								assign node805 = (inp[2]) ? 4'b1001 : node806;
									assign node806 = (inp[9]) ? node808 : 4'b1011;
										assign node808 = (inp[7]) ? 4'b1001 : node809;
											assign node809 = (inp[8]) ? 4'b1001 : node810;
												assign node810 = (inp[15]) ? node812 : 4'b1011;
													assign node812 = (inp[1]) ? node814 : 4'b1011;
														assign node814 = (inp[11]) ? 4'b1001 : 4'b1011;
			assign node820 = (inp[12]) ? node1028 : node821;
				assign node821 = (inp[6]) ? node925 : node822;
					assign node822 = (inp[13]) ? node884 : node823;
						assign node823 = (inp[4]) ? node849 : node824;
							assign node824 = (inp[2]) ? node826 : 4'b0111;
								assign node826 = (inp[9]) ? node828 : 4'b0111;
									assign node828 = (inp[8]) ? node830 : 4'b0111;
										assign node830 = (inp[14]) ? node840 : node831;
											assign node831 = (inp[7]) ? node833 : 4'b0111;
												assign node833 = (inp[15]) ? node835 : 4'b0111;
													assign node835 = (inp[1]) ? node837 : 4'b0111;
														assign node837 = (inp[11]) ? 4'b0101 : 4'b0111;
											assign node840 = (inp[7]) ? 4'b0101 : node841;
												assign node841 = (inp[15]) ? node843 : 4'b0111;
													assign node843 = (inp[11]) ? node845 : 4'b0111;
														assign node845 = (inp[1]) ? 4'b0101 : 4'b0111;
							assign node849 = (inp[2]) ? node877 : node850;
								assign node850 = (inp[14]) ? node864 : node851;
									assign node851 = (inp[9]) ? node853 : 4'b0111;
										assign node853 = (inp[8]) ? 4'b0101 : node854;
											assign node854 = (inp[15]) ? node856 : 4'b0111;
												assign node856 = (inp[1]) ? node858 : 4'b0111;
													assign node858 = (inp[11]) ? node860 : 4'b0111;
														assign node860 = (inp[7]) ? 4'b0101 : 4'b0111;
									assign node864 = (inp[9]) ? 4'b0101 : node865;
										assign node865 = (inp[7]) ? 4'b0101 : node866;
											assign node866 = (inp[8]) ? 4'b0101 : node867;
												assign node867 = (inp[1]) ? node869 : 4'b0111;
													assign node869 = (inp[11]) ? node871 : 4'b0111;
														assign node871 = (inp[15]) ? 4'b0101 : 4'b0111;
								assign node877 = (inp[9]) ? node879 : 4'b0101;
									assign node879 = (inp[8]) ? node881 : 4'b0101;
										assign node881 = (inp[14]) ? 4'b0011 : 4'b0101;
						assign node884 = (inp[4]) ? node898 : node885;
							assign node885 = (inp[8]) ? node887 : 4'b0101;
								assign node887 = (inp[2]) ? node889 : 4'b0101;
									assign node889 = (inp[9]) ? node891 : 4'b0101;
										assign node891 = (inp[14]) ? 4'b0011 : node892;
											assign node892 = (inp[15]) ? node894 : 4'b0101;
												assign node894 = (inp[7]) ? 4'b0111 : 4'b0101;
							assign node898 = (inp[14]) ? node910 : node899;
								assign node899 = (inp[9]) ? 4'b0111 : node900;
									assign node900 = (inp[2]) ? 4'b0111 : node901;
										assign node901 = (inp[7]) ? node903 : 4'b0101;
											assign node903 = (inp[15]) ? node905 : 4'b0101;
												assign node905 = (inp[8]) ? 4'b0111 : 4'b0101;
								assign node910 = (inp[2]) ? node912 : 4'b0011;
									assign node912 = (inp[9]) ? 4'b0001 : node913;
										assign node913 = (inp[8]) ? node915 : 4'b0011;
											assign node915 = (inp[7]) ? 4'b0001 : node916;
												assign node916 = (inp[11]) ? node918 : 4'b0011;
													assign node918 = (inp[15]) ? node920 : 4'b0011;
														assign node920 = (inp[1]) ? 4'b0001 : 4'b0011;
					assign node925 = (inp[14]) ? node981 : node926;
						assign node926 = (inp[13]) ? node954 : node927;
							assign node927 = (inp[2]) ? node939 : node928;
								assign node928 = (inp[4]) ? node930 : 4'b0011;
									assign node930 = (inp[8]) ? node932 : 4'b0001;
										assign node932 = (inp[7]) ? node934 : 4'b0001;
											assign node934 = (inp[9]) ? node936 : 4'b0001;
												assign node936 = (inp[15]) ? 4'b0011 : 4'b0001;
								assign node939 = (inp[9]) ? node941 : 4'b0011;
									assign node941 = (inp[4]) ? 4'b0011 : node942;
										assign node942 = (inp[8]) ? 4'b0001 : node943;
											assign node943 = (inp[7]) ? 4'b0001 : node944;
												assign node944 = (inp[11]) ? node946 : 4'b0011;
													assign node946 = (inp[1]) ? node948 : 4'b0011;
														assign node948 = (inp[15]) ? 4'b0001 : 4'b0011;
							assign node954 = (inp[2]) ? node970 : node955;
								assign node955 = (inp[9]) ? 4'b0001 : node956;
									assign node956 = (inp[4]) ? node958 : 4'b0001;
										assign node958 = (inp[1]) ? node960 : 4'b0011;
											assign node960 = (inp[11]) ? node962 : 4'b0011;
												assign node962 = (inp[15]) ? node964 : 4'b0011;
													assign node964 = (inp[8]) ? node966 : 4'b0011;
														assign node966 = (inp[7]) ? 4'b0001 : 4'b0011;
								assign node970 = (inp[4]) ? 4'b0001 : node971;
									assign node971 = (inp[9]) ? 4'b0011 : node972;
										assign node972 = (inp[15]) ? node974 : 4'b0001;
											assign node974 = (inp[8]) ? node976 : 4'b0001;
												assign node976 = (inp[7]) ? 4'b0011 : 4'b0001;
						assign node981 = (inp[4]) ? node1001 : node982;
							assign node982 = (inp[13]) ? node998 : node983;
								assign node983 = (inp[2]) ? node985 : 4'b0011;
									assign node985 = (inp[9]) ? 4'b0001 : node986;
										assign node986 = (inp[8]) ? 4'b0001 : node987;
											assign node987 = (inp[1]) ? node989 : 4'b0011;
												assign node989 = (inp[7]) ? node991 : 4'b0011;
													assign node991 = (inp[11]) ? node993 : 4'b0011;
														assign node993 = (inp[15]) ? 4'b0001 : 4'b0011;
								assign node998 = (inp[2]) ? 4'b0111 : 4'b0001;
							assign node1001 = (inp[2]) ? node1013 : node1002;
								assign node1002 = (inp[13]) ? node1004 : 4'b0110;
									assign node1004 = (inp[9]) ? node1006 : 4'b0100;
										assign node1006 = (inp[8]) ? node1008 : 4'b0100;
											assign node1008 = (inp[15]) ? node1010 : 4'b0100;
												assign node1010 = (inp[7]) ? 4'b0110 : 4'b0100;
								assign node1013 = (inp[13]) ? 4'b0110 : node1014;
									assign node1014 = (inp[9]) ? 4'b0100 : node1015;
										assign node1015 = (inp[15]) ? node1017 : 4'b0110;
											assign node1017 = (inp[11]) ? node1019 : 4'b0110;
												assign node1019 = (inp[8]) ? node1021 : 4'b0110;
													assign node1021 = (inp[1]) ? node1023 : 4'b0110;
														assign node1023 = (inp[7]) ? 4'b0100 : 4'b0110;
				assign node1028 = (inp[4]) ? node1172 : node1029;
					assign node1029 = (inp[14]) ? node1109 : node1030;
						assign node1030 = (inp[13]) ? node1074 : node1031;
							assign node1031 = (inp[2]) ? node1057 : node1032;
								assign node1032 = (inp[9]) ? 4'b0100 : node1033;
									assign node1033 = (inp[8]) ? node1045 : node1034;
										assign node1034 = (inp[1]) ? node1036 : 4'b0110;
											assign node1036 = (inp[6]) ? node1038 : 4'b0110;
												assign node1038 = (inp[15]) ? node1040 : 4'b0110;
													assign node1040 = (inp[11]) ? node1042 : 4'b0110;
														assign node1042 = (inp[7]) ? 4'b0100 : 4'b0110;
										assign node1045 = (inp[7]) ? 4'b0100 : node1046;
											assign node1046 = (inp[6]) ? 4'b0100 : node1047;
												assign node1047 = (inp[1]) ? node1049 : 4'b0110;
													assign node1049 = (inp[15]) ? node1051 : 4'b0110;
														assign node1051 = (inp[11]) ? 4'b0100 : 4'b0110;
								assign node1057 = (inp[9]) ? node1067 : node1058;
									assign node1058 = (inp[7]) ? node1060 : 4'b0100;
										assign node1060 = (inp[15]) ? node1062 : 4'b0100;
											assign node1062 = (inp[8]) ? node1064 : 4'b0100;
												assign node1064 = (inp[6]) ? 4'b0110 : 4'b0100;
									assign node1067 = (inp[8]) ? node1071 : node1068;
										assign node1068 = (inp[6]) ? 4'b0110 : 4'b0100;
										assign node1071 = (inp[6]) ? 4'b0110 : 4'b0010;
							assign node1074 = (inp[6]) ? node1090 : node1075;
								assign node1075 = (inp[2]) ? node1077 : 4'b0010;
									assign node1077 = (inp[7]) ? 4'b0000 : node1078;
										assign node1078 = (inp[9]) ? 4'b0000 : node1079;
											assign node1079 = (inp[8]) ? 4'b0000 : node1080;
												assign node1080 = (inp[11]) ? node1082 : 4'b0010;
													assign node1082 = (inp[15]) ? node1084 : 4'b0010;
														assign node1084 = (inp[1]) ? 4'b0000 : 4'b0010;
								assign node1090 = (inp[2]) ? node1104 : node1091;
									assign node1091 = (inp[9]) ? node1093 : 4'b0110;
										assign node1093 = (inp[7]) ? 4'b0100 : node1094;
											assign node1094 = (inp[8]) ? 4'b0100 : node1095;
												assign node1095 = (inp[1]) ? node1097 : 4'b0110;
													assign node1097 = (inp[11]) ? node1099 : 4'b0110;
														assign node1099 = (inp[15]) ? 4'b0100 : 4'b0110;
									assign node1104 = (inp[8]) ? node1106 : 4'b0100;
										assign node1106 = (inp[9]) ? 4'b0010 : 4'b0100;
						assign node1109 = (inp[2]) ? node1145 : node1110;
							assign node1110 = (inp[6]) ? node1122 : node1111;
								assign node1111 = (inp[13]) ? 4'b0000 : node1112;
									assign node1112 = (inp[9]) ? 4'b0010 : node1113;
										assign node1113 = (inp[15]) ? node1115 : 4'b0000;
											assign node1115 = (inp[8]) ? node1117 : 4'b0000;
												assign node1117 = (inp[7]) ? 4'b0010 : 4'b0000;
								assign node1122 = (inp[9]) ? node1124 : 4'b0010;
									assign node1124 = (inp[8]) ? node1126 : 4'b0010;
										assign node1126 = (inp[13]) ? node1136 : node1127;
											assign node1127 = (inp[7]) ? 4'b0000 : node1128;
												assign node1128 = (inp[1]) ? node1130 : 4'b0010;
													assign node1130 = (inp[11]) ? node1132 : 4'b0010;
														assign node1132 = (inp[15]) ? 4'b0000 : 4'b0010;
											assign node1136 = (inp[15]) ? node1138 : 4'b0010;
												assign node1138 = (inp[1]) ? node1140 : 4'b0010;
													assign node1140 = (inp[7]) ? node1142 : 4'b0010;
														assign node1142 = (inp[11]) ? 4'b0000 : 4'b0010;
							assign node1145 = (inp[6]) ? node1161 : node1146;
								assign node1146 = (inp[13]) ? 4'b0110 : node1147;
									assign node1147 = (inp[9]) ? node1149 : 4'b0010;
										assign node1149 = (inp[8]) ? 4'b0000 : node1150;
											assign node1150 = (inp[7]) ? node1152 : 4'b0010;
												assign node1152 = (inp[11]) ? node1154 : 4'b0010;
													assign node1154 = (inp[15]) ? node1156 : 4'b0010;
														assign node1156 = (inp[1]) ? 4'b0000 : 4'b0010;
								assign node1161 = (inp[13]) ? 4'b0000 : node1162;
									assign node1162 = (inp[9]) ? node1164 : 4'b0000;
										assign node1164 = (inp[15]) ? node1166 : 4'b0000;
											assign node1166 = (inp[7]) ? node1168 : 4'b0000;
												assign node1168 = (inp[8]) ? 4'b0010 : 4'b0000;
					assign node1172 = (inp[14]) ? node1316 : node1173;
						assign node1173 = (inp[6]) ? node1209 : node1174;
							assign node1174 = (inp[2]) ? node1198 : node1175;
								assign node1175 = (inp[9]) ? node1177 : 4'b0111;
									assign node1177 = (inp[8]) ? node1179 : 4'b0111;
										assign node1179 = (inp[7]) ? node1189 : node1180;
											assign node1180 = (inp[15]) ? node1182 : 4'b0111;
												assign node1182 = (inp[1]) ? node1184 : 4'b0111;
													assign node1184 = (inp[13]) ? node1186 : 4'b0111;
														assign node1186 = (inp[11]) ? 4'b0101 : 4'b0111;
											assign node1189 = (inp[13]) ? 4'b0101 : node1190;
												assign node1190 = (inp[1]) ? node1192 : 4'b0111;
													assign node1192 = (inp[15]) ? node1194 : 4'b0111;
														assign node1194 = (inp[11]) ? 4'b0101 : 4'b0111;
								assign node1198 = (inp[9]) ? node1200 : 4'b0101;
									assign node1200 = (inp[8]) ? node1202 : 4'b0101;
										assign node1202 = (inp[13]) ? 4'b0011 : node1203;
											assign node1203 = (inp[7]) ? node1205 : 4'b0101;
												assign node1205 = (inp[15]) ? 4'b0111 : 4'b0101;
							assign node1209 = (inp[13]) ? node1285 : node1210;
								assign node1210 = (inp[9]) ? node1278 : node1211;
									assign node1211 = (inp[15]) ? node1219 : node1212;
										assign node1212 = (inp[2]) ? node1214 : 4'b0101;
											assign node1214 = (inp[8]) ? 4'b0101 : node1215;
												assign node1215 = (inp[7]) ? 4'b0101 : 4'b0111;
										assign node1219 = (inp[11]) ? node1265 : node1220;
											assign node1220 = (inp[3]) ? node1254 : node1221;
												assign node1221 = (inp[1]) ? node1243 : node1222;
													assign node1222 = (inp[0]) ? node1234 : node1223;
														assign node1223 = (inp[8]) ? node1229 : node1224;
															assign node1224 = (inp[2]) ? node1226 : 4'b0101;
																assign node1226 = (inp[7]) ? 4'b0101 : 4'b0111;
															assign node1229 = (inp[2]) ? 4'b0101 : node1230;
																assign node1230 = (inp[7]) ? 4'b0111 : 4'b0101;
														assign node1234 = (inp[7]) ? node1240 : node1235;
															assign node1235 = (inp[2]) ? node1237 : 4'b0101;
																assign node1237 = (inp[8]) ? 4'b0101 : 4'b0111;
															assign node1240 = (inp[8]) ? 4'b0111 : 4'b0101;
													assign node1243 = (inp[7]) ? node1249 : node1244;
														assign node1244 = (inp[8]) ? 4'b0101 : node1245;
															assign node1245 = (inp[2]) ? 4'b0111 : 4'b0101;
														assign node1249 = (inp[8]) ? node1251 : 4'b0101;
															assign node1251 = (inp[2]) ? 4'b0101 : 4'b0111;
												assign node1254 = (inp[2]) ? node1260 : node1255;
													assign node1255 = (inp[7]) ? node1257 : 4'b0101;
														assign node1257 = (inp[8]) ? 4'b0111 : 4'b0101;
													assign node1260 = (inp[7]) ? 4'b0101 : node1261;
														assign node1261 = (inp[8]) ? 4'b0101 : 4'b0111;
											assign node1265 = (inp[7]) ? node1273 : node1266;
												assign node1266 = (inp[2]) ? node1268 : 4'b0101;
													assign node1268 = (inp[1]) ? 4'b0101 : node1269;
														assign node1269 = (inp[8]) ? 4'b0101 : 4'b0111;
												assign node1273 = (inp[8]) ? node1275 : 4'b0101;
													assign node1275 = (inp[2]) ? 4'b0101 : 4'b0111;
									assign node1278 = (inp[8]) ? node1282 : node1279;
										assign node1279 = (inp[2]) ? 4'b0101 : 4'b0111;
										assign node1282 = (inp[2]) ? 4'b0011 : 4'b0111;
								assign node1285 = (inp[9]) ? node1307 : node1286;
									assign node1286 = (inp[8]) ? node1288 : 4'b0011;
										assign node1288 = (inp[2]) ? node1298 : node1289;
											assign node1289 = (inp[7]) ? 4'b0001 : node1290;
												assign node1290 = (inp[15]) ? node1292 : 4'b0011;
													assign node1292 = (inp[1]) ? node1294 : 4'b0011;
														assign node1294 = (inp[11]) ? 4'b0001 : 4'b0011;
											assign node1298 = (inp[15]) ? node1300 : 4'b0011;
												assign node1300 = (inp[1]) ? node1302 : 4'b0011;
													assign node1302 = (inp[7]) ? node1304 : 4'b0011;
														assign node1304 = (inp[11]) ? 4'b0001 : 4'b0011;
									assign node1307 = (inp[7]) ? node1309 : 4'b0001;
										assign node1309 = (inp[8]) ? node1311 : 4'b0001;
											assign node1311 = (inp[2]) ? 4'b0001 : node1312;
												assign node1312 = (inp[15]) ? 4'b0011 : 4'b0001;
						assign node1316 = (inp[6]) ? node1368 : node1317;
							assign node1317 = (inp[2]) ? node1345 : node1318;
								assign node1318 = (inp[9]) ? node1332 : node1319;
									assign node1319 = (inp[13]) ? node1321 : 4'b0011;
										assign node1321 = (inp[8]) ? 4'b0001 : node1322;
											assign node1322 = (inp[11]) ? node1324 : 4'b0011;
												assign node1324 = (inp[15]) ? node1326 : 4'b0011;
													assign node1326 = (inp[7]) ? node1328 : 4'b0011;
														assign node1328 = (inp[1]) ? 4'b0001 : 4'b0011;
									assign node1332 = (inp[13]) ? 4'b0001 : node1333;
										assign node1333 = (inp[8]) ? 4'b0001 : node1334;
											assign node1334 = (inp[7]) ? 4'b0001 : node1335;
												assign node1335 = (inp[1]) ? node1337 : 4'b0011;
													assign node1337 = (inp[15]) ? node1339 : 4'b0011;
														assign node1339 = (inp[11]) ? 4'b0001 : 4'b0011;
								assign node1345 = (inp[13]) ? node1355 : node1346;
									assign node1346 = (inp[9]) ? 4'b0011 : node1347;
										assign node1347 = (inp[8]) ? node1349 : 4'b0001;
											assign node1349 = (inp[15]) ? node1351 : 4'b0001;
												assign node1351 = (inp[7]) ? 4'b0011 : 4'b0001;
									assign node1355 = (inp[9]) ? node1357 : 4'b0111;
										assign node1357 = (inp[8]) ? 4'b0101 : node1358;
											assign node1358 = (inp[1]) ? node1360 : 4'b0111;
												assign node1360 = (inp[15]) ? node1362 : 4'b0111;
													assign node1362 = (inp[11]) ? node1364 : 4'b0111;
														assign node1364 = (inp[7]) ? 4'b0101 : 4'b0111;
							assign node1368 = (inp[13]) ? node1400 : node1369;
								assign node1369 = (inp[9]) ? node1391 : node1370;
									assign node1370 = (inp[8]) ? node1372 : 4'b0110;
										assign node1372 = (inp[2]) ? node1382 : node1373;
											assign node1373 = (inp[7]) ? node1375 : 4'b0110;
												assign node1375 = (inp[1]) ? node1377 : 4'b0110;
													assign node1377 = (inp[15]) ? node1379 : 4'b0110;
														assign node1379 = (inp[11]) ? 4'b0100 : 4'b0110;
											assign node1382 = (inp[7]) ? 4'b0100 : node1383;
												assign node1383 = (inp[15]) ? node1385 : 4'b0110;
													assign node1385 = (inp[1]) ? node1387 : 4'b0110;
														assign node1387 = (inp[11]) ? 4'b0100 : 4'b0110;
									assign node1391 = (inp[8]) ? node1393 : 4'b0100;
										assign node1393 = (inp[2]) ? 4'b0010 : node1394;
											assign node1394 = (inp[15]) ? node1396 : 4'b0100;
												assign node1396 = (inp[7]) ? 4'b0110 : 4'b0100;
								assign node1400 = (inp[2]) ? node1428 : node1401;
									assign node1401 = (inp[8]) ? node1421 : node1402;
										assign node1402 = (inp[9]) ? node1412 : node1403;
											assign node1403 = (inp[7]) ? 4'b0000 : node1404;
												assign node1404 = (inp[15]) ? node1406 : 4'b0010;
													assign node1406 = (inp[1]) ? node1408 : 4'b0010;
														assign node1408 = (inp[11]) ? 4'b0000 : 4'b0010;
											assign node1412 = (inp[11]) ? node1414 : 4'b0010;
												assign node1414 = (inp[15]) ? node1416 : 4'b0010;
													assign node1416 = (inp[1]) ? node1418 : 4'b0010;
														assign node1418 = (inp[7]) ? 4'b0000 : 4'b0010;
										assign node1421 = (inp[7]) ? node1423 : 4'b0000;
											assign node1423 = (inp[15]) ? node1425 : 4'b0000;
												assign node1425 = (inp[9]) ? 4'b0000 : 4'b0010;
									assign node1428 = (inp[8]) ? node1448 : node1429;
										assign node1429 = (inp[9]) ? node1439 : node1430;
											assign node1430 = (inp[7]) ? node1432 : 4'b0110;
												assign node1432 = (inp[15]) ? node1434 : 4'b0110;
													assign node1434 = (inp[11]) ? node1436 : 4'b0110;
														assign node1436 = (inp[1]) ? 4'b0100 : 4'b0110;
											assign node1439 = (inp[7]) ? 4'b0100 : node1440;
												assign node1440 = (inp[11]) ? node1442 : 4'b0110;
													assign node1442 = (inp[1]) ? node1444 : 4'b0110;
														assign node1444 = (inp[15]) ? 4'b0100 : 4'b0110;
										assign node1448 = (inp[9]) ? node1454 : node1449;
											assign node1449 = (inp[7]) ? node1451 : 4'b0100;
												assign node1451 = (inp[15]) ? 4'b0110 : 4'b0100;
											assign node1454 = (inp[7]) ? node1462 : node1455;
												assign node1455 = (inp[1]) ? node1457 : 4'b0010;
													assign node1457 = (inp[15]) ? node1459 : 4'b0010;
														assign node1459 = (inp[11]) ? 4'b0000 : 4'b0010;
												assign node1462 = (inp[15]) ? node1464 : 4'b0000;
													assign node1464 = (inp[1]) ? node1466 : 4'b0010;
														assign node1466 = (inp[11]) ? 4'b0000 : 4'b0010;

endmodule