module dtc_split75_bm66 (
	input  wire [16-1:0] inp,
	output wire [4-1:0] outp
);

	wire [4-1:0] node1;
	wire [4-1:0] node2;
	wire [4-1:0] node3;
	wire [4-1:0] node4;
	wire [4-1:0] node6;
	wire [4-1:0] node7;
	wire [4-1:0] node9;
	wire [4-1:0] node11;
	wire [4-1:0] node13;
	wire [4-1:0] node14;
	wire [4-1:0] node16;
	wire [4-1:0] node18;
	wire [4-1:0] node20;
	wire [4-1:0] node23;
	wire [4-1:0] node24;
	wire [4-1:0] node26;
	wire [4-1:0] node28;
	wire [4-1:0] node32;
	wire [4-1:0] node33;
	wire [4-1:0] node34;
	wire [4-1:0] node36;
	wire [4-1:0] node37;
	wire [4-1:0] node39;
	wire [4-1:0] node41;
	wire [4-1:0] node43;
	wire [4-1:0] node47;
	wire [4-1:0] node48;
	wire [4-1:0] node49;
	wire [4-1:0] node50;
	wire [4-1:0] node52;
	wire [4-1:0] node54;
	wire [4-1:0] node61;
	wire [4-1:0] node62;
	wire [4-1:0] node64;
	wire [4-1:0] node66;
	wire [4-1:0] node68;
	wire [4-1:0] node70;
	wire [4-1:0] node73;
	wire [4-1:0] node74;
	wire [4-1:0] node76;
	wire [4-1:0] node78;
	wire [4-1:0] node80;
	wire [4-1:0] node81;
	wire [4-1:0] node83;
	wire [4-1:0] node87;
	wire [4-1:0] node88;
	wire [4-1:0] node89;
	wire [4-1:0] node90;
	wire [4-1:0] node92;
	wire [4-1:0] node94;
	wire [4-1:0] node100;
	wire [4-1:0] node101;
	wire [4-1:0] node102;
	wire [4-1:0] node103;
	wire [4-1:0] node105;
	wire [4-1:0] node107;
	wire [4-1:0] node109;
	wire [4-1:0] node110;
	wire [4-1:0] node111;
	wire [4-1:0] node113;
	wire [4-1:0] node115;
	wire [4-1:0] node120;
	wire [4-1:0] node121;
	wire [4-1:0] node123;
	wire [4-1:0] node124;
	wire [4-1:0] node126;
	wire [4-1:0] node127;
	wire [4-1:0] node129;
	wire [4-1:0] node131;
	wire [4-1:0] node137;
	wire [4-1:0] node138;
	wire [4-1:0] node140;
	wire [4-1:0] node142;
	wire [4-1:0] node143;
	wire [4-1:0] node145;
	wire [4-1:0] node147;
	wire [4-1:0] node151;
	wire [4-1:0] node152;
	wire [4-1:0] node153;
	wire [4-1:0] node155;
	wire [4-1:0] node157;
	wire [4-1:0] node159;
	wire [4-1:0] node164;
	wire [4-1:0] node165;
	wire [4-1:0] node166;
	wire [4-1:0] node168;
	wire [4-1:0] node170;
	wire [4-1:0] node171;
	wire [4-1:0] node172;
	wire [4-1:0] node174;
	wire [4-1:0] node176;
	wire [4-1:0] node178;
	wire [4-1:0] node183;
	wire [4-1:0] node184;
	wire [4-1:0] node185;
	wire [4-1:0] node186;
	wire [4-1:0] node188;
	wire [4-1:0] node190;
	wire [4-1:0] node192;
	wire [4-1:0] node194;
	wire [4-1:0] node200;
	wire [4-1:0] node201;
	wire [4-1:0] node203;
	wire [4-1:0] node206;
	wire [4-1:0] node208;
	wire [4-1:0] node210;
	wire [4-1:0] node211;
	wire [4-1:0] node213;
	wire [4-1:0] node215;
	wire [4-1:0] node217;
	wire [4-1:0] node219;
	wire [4-1:0] node223;
	wire [4-1:0] node224;
	wire [4-1:0] node225;
	wire [4-1:0] node226;
	wire [4-1:0] node227;
	wire [4-1:0] node228;
	wire [4-1:0] node230;
	wire [4-1:0] node231;
	wire [4-1:0] node233;
	wire [4-1:0] node235;
	wire [4-1:0] node239;
	wire [4-1:0] node240;
	wire [4-1:0] node241;
	wire [4-1:0] node242;
	wire [4-1:0] node244;
	wire [4-1:0] node246;
	wire [4-1:0] node248;
	wire [4-1:0] node254;
	wire [4-1:0] node255;
	wire [4-1:0] node257;
	wire [4-1:0] node259;
	wire [4-1:0] node262;
	wire [4-1:0] node263;
	wire [4-1:0] node264;
	wire [4-1:0] node266;
	wire [4-1:0] node267;
	wire [4-1:0] node269;
	wire [4-1:0] node271;
	wire [4-1:0] node277;
	wire [4-1:0] node278;
	wire [4-1:0] node280;
	wire [4-1:0] node282;
	wire [4-1:0] node284;
	wire [4-1:0] node286;
	wire [4-1:0] node288;
	wire [4-1:0] node291;
	wire [4-1:0] node292;
	wire [4-1:0] node296;
	wire [4-1:0] node297;
	wire [4-1:0] node298;
	wire [4-1:0] node299;
	wire [4-1:0] node301;
	wire [4-1:0] node303;
	wire [4-1:0] node304;
	wire [4-1:0] node306;
	wire [4-1:0] node308;
	wire [4-1:0] node310;
	wire [4-1:0] node315;
	wire [4-1:0] node316;
	wire [4-1:0] node318;
	wire [4-1:0] node319;
	wire [4-1:0] node321;
	wire [4-1:0] node323;
	wire [4-1:0] node325;
	wire [4-1:0] node327;
	wire [4-1:0] node332;
	wire [4-1:0] node333;
	wire [4-1:0] node334;
	wire [4-1:0] node335;
	wire [4-1:0] node336;
	wire [4-1:0] node338;
	wire [4-1:0] node340;
	wire [4-1:0] node345;
	wire [4-1:0] node347;
	wire [4-1:0] node348;
	wire [4-1:0] node349;
	wire [4-1:0] node350;
	wire [4-1:0] node352;
	wire [4-1:0] node354;
	wire [4-1:0] node360;
	wire [4-1:0] node362;
	wire [4-1:0] node363;
	wire [4-1:0] node364;
	wire [4-1:0] node366;
	wire [4-1:0] node368;
	wire [4-1:0] node370;
	wire [4-1:0] node375;
	wire [4-1:0] node376;
	wire [4-1:0] node377;
	wire [4-1:0] node378;
	wire [4-1:0] node379;
	wire [4-1:0] node380;
	wire [4-1:0] node383;
	wire [4-1:0] node385;
	wire [4-1:0] node387;
	wire [4-1:0] node388;
	wire [4-1:0] node390;
	wire [4-1:0] node392;
	wire [4-1:0] node396;
	wire [4-1:0] node397;
	wire [4-1:0] node398;
	wire [4-1:0] node400;
	wire [4-1:0] node402;
	wire [4-1:0] node406;
	wire [4-1:0] node409;
	wire [4-1:0] node410;
	wire [4-1:0] node412;
	wire [4-1:0] node413;
	wire [4-1:0] node414;
	wire [4-1:0] node416;
	wire [4-1:0] node418;
	wire [4-1:0] node420;
	wire [4-1:0] node425;
	wire [4-1:0] node427;
	wire [4-1:0] node428;
	wire [4-1:0] node430;
	wire [4-1:0] node432;
	wire [4-1:0] node436;
	wire [4-1:0] node437;
	wire [4-1:0] node438;
	wire [4-1:0] node440;
	wire [4-1:0] node442;
	wire [4-1:0] node445;
	wire [4-1:0] node447;
	wire [4-1:0] node449;
	wire [4-1:0] node450;
	wire [4-1:0] node451;
	wire [4-1:0] node453;
	wire [4-1:0] node455;
	wire [4-1:0] node460;
	wire [4-1:0] node462;
	wire [4-1:0] node464;
	wire [4-1:0] node466;
	wire [4-1:0] node469;
	wire [4-1:0] node470;
	wire [4-1:0] node471;
	wire [4-1:0] node472;
	wire [4-1:0] node473;
	wire [4-1:0] node474;
	wire [4-1:0] node475;
	wire [4-1:0] node476;
	wire [4-1:0] node478;
	wire [4-1:0] node480;
	wire [4-1:0] node486;
	wire [4-1:0] node488;
	wire [4-1:0] node489;
	wire [4-1:0] node491;
	wire [4-1:0] node492;
	wire [4-1:0] node493;
	wire [4-1:0] node495;
	wire [4-1:0] node502;
	wire [4-1:0] node504;
	wire [4-1:0] node506;
	wire [4-1:0] node508;
	wire [4-1:0] node509;
	wire [4-1:0] node510;
	wire [4-1:0] node512;
	wire [4-1:0] node514;
	wire [4-1:0] node518;
	wire [4-1:0] node520;
	wire [4-1:0] node522;
	wire [4-1:0] node524;
	wire [4-1:0] node527;
	wire [4-1:0] node528;
	wire [4-1:0] node529;
	wire [4-1:0] node530;
	wire [4-1:0] node531;
	wire [4-1:0] node533;
	wire [4-1:0] node535;
	wire [4-1:0] node540;
	wire [4-1:0] node543;
	wire [4-1:0] node545;
	wire [4-1:0] node547;
	wire [4-1:0] node549;
	wire [4-1:0] node551;
	wire [4-1:0] node552;
	wire [4-1:0] node556;
	wire [4-1:0] node557;
	wire [4-1:0] node558;
	wire [4-1:0] node559;
	wire [4-1:0] node560;
	wire [4-1:0] node561;
	wire [4-1:0] node562;
	wire [4-1:0] node564;
	wire [4-1:0] node566;
	wire [4-1:0] node567;
	wire [4-1:0] node568;
	wire [4-1:0] node570;
	wire [4-1:0] node572;
	wire [4-1:0] node578;
	wire [4-1:0] node579;
	wire [4-1:0] node581;
	wire [4-1:0] node583;
	wire [4-1:0] node585;
	wire [4-1:0] node586;
	wire [4-1:0] node590;
	wire [4-1:0] node592;
	wire [4-1:0] node594;
	wire [4-1:0] node597;
	wire [4-1:0] node598;
	wire [4-1:0] node600;
	wire [4-1:0] node601;
	wire [4-1:0] node602;
	wire [4-1:0] node604;
	wire [4-1:0] node605;
	wire [4-1:0] node607;
	wire [4-1:0] node609;
	wire [4-1:0] node615;
	wire [4-1:0] node617;
	wire [4-1:0] node618;
	wire [4-1:0] node620;
	wire [4-1:0] node622;
	wire [4-1:0] node623;
	wire [4-1:0] node625;
	wire [4-1:0] node627;
	wire [4-1:0] node632;
	wire [4-1:0] node633;
	wire [4-1:0] node634;
	wire [4-1:0] node635;
	wire [4-1:0] node637;
	wire [4-1:0] node639;
	wire [4-1:0] node642;
	wire [4-1:0] node644;
	wire [4-1:0] node646;
	wire [4-1:0] node648;
	wire [4-1:0] node650;
	wire [4-1:0] node654;
	wire [4-1:0] node655;
	wire [4-1:0] node656;
	wire [4-1:0] node658;
	wire [4-1:0] node660;
	wire [4-1:0] node662;
	wire [4-1:0] node664;
	wire [4-1:0] node666;
	wire [4-1:0] node668;
	wire [4-1:0] node671;
	wire [4-1:0] node672;
	wire [4-1:0] node673;
	wire [4-1:0] node674;
	wire [4-1:0] node675;
	wire [4-1:0] node677;
	wire [4-1:0] node679;
	wire [4-1:0] node687;
	wire [4-1:0] node688;
	wire [4-1:0] node689;
	wire [4-1:0] node690;
	wire [4-1:0] node691;
	wire [4-1:0] node692;
	wire [4-1:0] node693;
	wire [4-1:0] node697;
	wire [4-1:0] node699;
	wire [4-1:0] node701;
	wire [4-1:0] node703;
	wire [4-1:0] node705;
	wire [4-1:0] node707;
	wire [4-1:0] node710;
	wire [4-1:0] node711;
	wire [4-1:0] node712;
	wire [4-1:0] node713;
	wire [4-1:0] node714;
	wire [4-1:0] node715;
	wire [4-1:0] node719;
	wire [4-1:0] node721;
	wire [4-1:0] node724;
	wire [4-1:0] node725;
	wire [4-1:0] node726;
	wire [4-1:0] node727;
	wire [4-1:0] node731;
	wire [4-1:0] node733;
	wire [4-1:0] node736;
	wire [4-1:0] node737;
	wire [4-1:0] node738;
	wire [4-1:0] node742;
	wire [4-1:0] node744;
	wire [4-1:0] node747;
	wire [4-1:0] node748;
	wire [4-1:0] node749;
	wire [4-1:0] node750;
	wire [4-1:0] node754;
	wire [4-1:0] node756;
	wire [4-1:0] node759;
	wire [4-1:0] node760;
	wire [4-1:0] node761;
	wire [4-1:0] node762;
	wire [4-1:0] node766;
	wire [4-1:0] node768;
	wire [4-1:0] node771;
	wire [4-1:0] node772;
	wire [4-1:0] node773;
	wire [4-1:0] node777;
	wire [4-1:0] node779;
	wire [4-1:0] node782;
	wire [4-1:0] node783;
	wire [4-1:0] node784;
	wire [4-1:0] node785;
	wire [4-1:0] node786;
	wire [4-1:0] node790;
	wire [4-1:0] node792;
	wire [4-1:0] node795;
	wire [4-1:0] node796;
	wire [4-1:0] node797;
	wire [4-1:0] node798;
	wire [4-1:0] node799;
	wire [4-1:0] node803;
	wire [4-1:0] node806;
	wire [4-1:0] node807;
	wire [4-1:0] node808;
	wire [4-1:0] node812;
	wire [4-1:0] node815;
	wire [4-1:0] node816;
	wire [4-1:0] node817;
	wire [4-1:0] node821;
	wire [4-1:0] node823;
	wire [4-1:0] node826;
	wire [4-1:0] node828;
	wire [4-1:0] node830;
	wire [4-1:0] node833;
	wire [4-1:0] node835;
	wire [4-1:0] node838;
	wire [4-1:0] node839;
	wire [4-1:0] node841;
	wire [4-1:0] node843;
	wire [4-1:0] node844;
	wire [4-1:0] node846;
	wire [4-1:0] node848;
	wire [4-1:0] node852;
	wire [4-1:0] node853;
	wire [4-1:0] node854;
	wire [4-1:0] node855;
	wire [4-1:0] node856;
	wire [4-1:0] node858;
	wire [4-1:0] node860;
	wire [4-1:0] node862;
	wire [4-1:0] node869;
	wire [4-1:0] node870;
	wire [4-1:0] node871;
	wire [4-1:0] node873;
	wire [4-1:0] node874;
	wire [4-1:0] node876;
	wire [4-1:0] node878;
	wire [4-1:0] node880;
	wire [4-1:0] node882;
	wire [4-1:0] node884;
	wire [4-1:0] node888;
	wire [4-1:0] node889;
	wire [4-1:0] node891;
	wire [4-1:0] node893;
	wire [4-1:0] node895;
	wire [4-1:0] node897;
	wire [4-1:0] node901;
	wire [4-1:0] node902;
	wire [4-1:0] node903;
	wire [4-1:0] node904;
	wire [4-1:0] node906;
	wire [4-1:0] node908;
	wire [4-1:0] node909;
	wire [4-1:0] node911;
	wire [4-1:0] node913;
	wire [4-1:0] node918;
	wire [4-1:0] node920;
	wire [4-1:0] node922;
	wire [4-1:0] node925;
	wire [4-1:0] node927;
	wire [4-1:0] node928;
	wire [4-1:0] node930;
	wire [4-1:0] node931;
	wire [4-1:0] node932;
	wire [4-1:0] node934;
	wire [4-1:0] node936;
	wire [4-1:0] node942;
	wire [4-1:0] node943;
	wire [4-1:0] node944;
	wire [4-1:0] node945;
	wire [4-1:0] node946;
	wire [4-1:0] node948;
	wire [4-1:0] node950;
	wire [4-1:0] node952;
	wire [4-1:0] node953;
	wire [4-1:0] node955;
	wire [4-1:0] node957;
	wire [4-1:0] node959;
	wire [4-1:0] node962;
	wire [4-1:0] node963;
	wire [4-1:0] node965;
	wire [4-1:0] node967;
	wire [4-1:0] node971;
	wire [4-1:0] node972;
	wire [4-1:0] node973;
	wire [4-1:0] node975;
	wire [4-1:0] node976;
	wire [4-1:0] node978;
	wire [4-1:0] node980;
	wire [4-1:0] node982;
	wire [4-1:0] node986;
	wire [4-1:0] node987;
	wire [4-1:0] node988;
	wire [4-1:0] node989;
	wire [4-1:0] node991;
	wire [4-1:0] node993;
	wire [4-1:0] node999;
	wire [4-1:0] node1001;
	wire [4-1:0] node1003;
	wire [4-1:0] node1006;
	wire [4-1:0] node1007;
	wire [4-1:0] node1009;
	wire [4-1:0] node1011;
	wire [4-1:0] node1013;
	wire [4-1:0] node1014;
	wire [4-1:0] node1016;
	wire [4-1:0] node1020;
	wire [4-1:0] node1021;
	wire [4-1:0] node1022;
	wire [4-1:0] node1023;
	wire [4-1:0] node1025;
	wire [4-1:0] node1027;
	wire [4-1:0] node1032;
	wire [4-1:0] node1034;
	wire [4-1:0] node1035;
	wire [4-1:0] node1037;
	wire [4-1:0] node1038;
	wire [4-1:0] node1040;
	wire [4-1:0] node1042;
	wire [4-1:0] node1047;
	wire [4-1:0] node1048;
	wire [4-1:0] node1049;
	wire [4-1:0] node1050;
	wire [4-1:0] node1052;
	wire [4-1:0] node1054;
	wire [4-1:0] node1055;
	wire [4-1:0] node1056;
	wire [4-1:0] node1058;
	wire [4-1:0] node1060;
	wire [4-1:0] node1065;
	wire [4-1:0] node1066;
	wire [4-1:0] node1068;
	wire [4-1:0] node1070;
	wire [4-1:0] node1072;
	wire [4-1:0] node1076;
	wire [4-1:0] node1077;
	wire [4-1:0] node1079;
	wire [4-1:0] node1080;
	wire [4-1:0] node1082;
	wire [4-1:0] node1084;
	wire [4-1:0] node1088;
	wire [4-1:0] node1089;
	wire [4-1:0] node1090;
	wire [4-1:0] node1092;
	wire [4-1:0] node1094;
	wire [4-1:0] node1096;
	wire [4-1:0] node1098;
	wire [4-1:0] node1103;
	wire [4-1:0] node1104;
	wire [4-1:0] node1105;
	wire [4-1:0] node1108;
	wire [4-1:0] node1109;
	wire [4-1:0] node1110;
	wire [4-1:0] node1111;
	wire [4-1:0] node1113;
	wire [4-1:0] node1115;
	wire [4-1:0] node1117;
	wire [4-1:0] node1123;
	wire [4-1:0] node1124;
	wire [4-1:0] node1126;
	wire [4-1:0] node1128;
	wire [4-1:0] node1130;
	wire [4-1:0] node1132;
	wire [4-1:0] node1135;
	wire [4-1:0] node1136;
	wire [4-1:0] node1137;
	wire [4-1:0] node1139;
	wire [4-1:0] node1141;
	wire [4-1:0] node1143;
	wire [4-1:0] node1145;
	wire [4-1:0] node1150;
	wire [4-1:0] node1151;
	wire [4-1:0] node1152;
	wire [4-1:0] node1153;
	wire [4-1:0] node1154;
	wire [4-1:0] node1155;
	wire [4-1:0] node1156;
	wire [4-1:0] node1158;
	wire [4-1:0] node1160;
	wire [4-1:0] node1162;
	wire [4-1:0] node1164;
	wire [4-1:0] node1167;
	wire [4-1:0] node1168;
	wire [4-1:0] node1169;
	wire [4-1:0] node1171;
	wire [4-1:0] node1173;
	wire [4-1:0] node1179;
	wire [4-1:0] node1180;
	wire [4-1:0] node1182;
	wire [4-1:0] node1184;
	wire [4-1:0] node1186;
	wire [4-1:0] node1189;
	wire [4-1:0] node1190;
	wire [4-1:0] node1193;
	wire [4-1:0] node1196;
	wire [4-1:0] node1197;
	wire [4-1:0] node1199;
	wire [4-1:0] node1200;
	wire [4-1:0] node1201;
	wire [4-1:0] node1202;
	wire [4-1:0] node1204;
	wire [4-1:0] node1206;
	wire [4-1:0] node1212;
	wire [4-1:0] node1213;
	wire [4-1:0] node1215;
	wire [4-1:0] node1216;
	wire [4-1:0] node1217;
	wire [4-1:0] node1219;
	wire [4-1:0] node1221;
	wire [4-1:0] node1226;
	wire [4-1:0] node1228;
	wire [4-1:0] node1231;
	wire [4-1:0] node1232;
	wire [4-1:0] node1233;
	wire [4-1:0] node1234;
	wire [4-1:0] node1235;
	wire [4-1:0] node1237;
	wire [4-1:0] node1239;
	wire [4-1:0] node1244;
	wire [4-1:0] node1246;
	wire [4-1:0] node1248;
	wire [4-1:0] node1249;
	wire [4-1:0] node1250;
	wire [4-1:0] node1252;
	wire [4-1:0] node1254;
	wire [4-1:0] node1258;
	wire [4-1:0] node1260;
	wire [4-1:0] node1262;
	wire [4-1:0] node1264;
	wire [4-1:0] node1267;
	wire [4-1:0] node1268;
	wire [4-1:0] node1269;
	wire [4-1:0] node1271;
	wire [4-1:0] node1272;
	wire [4-1:0] node1274;
	wire [4-1:0] node1276;
	wire [4-1:0] node1278;
	wire [4-1:0] node1283;
	wire [4-1:0] node1284;
	wire [4-1:0] node1286;
	wire [4-1:0] node1288;
	wire [4-1:0] node1290;
	wire [4-1:0] node1294;
	wire [4-1:0] node1295;
	wire [4-1:0] node1296;
	wire [4-1:0] node1297;
	wire [4-1:0] node1298;
	wire [4-1:0] node1300;
	wire [4-1:0] node1302;
	wire [4-1:0] node1304;
	wire [4-1:0] node1307;
	wire [4-1:0] node1309;
	wire [4-1:0] node1311;
	wire [4-1:0] node1313;
	wire [4-1:0] node1315;
	wire [4-1:0] node1317;
	wire [4-1:0] node1320;
	wire [4-1:0] node1321;
	wire [4-1:0] node1323;
	wire [4-1:0] node1325;
	wire [4-1:0] node1327;
	wire [4-1:0] node1330;
	wire [4-1:0] node1331;
	wire [4-1:0] node1332;
	wire [4-1:0] node1333;
	wire [4-1:0] node1335;
	wire [4-1:0] node1337;
	wire [4-1:0] node1342;
	wire [4-1:0] node1345;
	wire [4-1:0] node1346;
	wire [4-1:0] node1347;
	wire [4-1:0] node1349;
	wire [4-1:0] node1351;
	wire [4-1:0] node1352;
	wire [4-1:0] node1354;
	wire [4-1:0] node1356;
	wire [4-1:0] node1360;
	wire [4-1:0] node1362;
	wire [4-1:0] node1365;
	wire [4-1:0] node1366;
	wire [4-1:0] node1368;
	wire [4-1:0] node1369;
	wire [4-1:0] node1371;
	wire [4-1:0] node1372;
	wire [4-1:0] node1374;
	wire [4-1:0] node1378;
	wire [4-1:0] node1380;
	wire [4-1:0] node1382;
	wire [4-1:0] node1384;
	wire [4-1:0] node1387;
	wire [4-1:0] node1389;
	wire [4-1:0] node1390;
	wire [4-1:0] node1392;
	wire [4-1:0] node1396;
	wire [4-1:0] node1397;
	wire [4-1:0] node1398;
	wire [4-1:0] node1399;
	wire [4-1:0] node1401;
	wire [4-1:0] node1402;
	wire [4-1:0] node1404;
	wire [4-1:0] node1406;
	wire [4-1:0] node1408;
	wire [4-1:0] node1412;
	wire [4-1:0] node1413;
	wire [4-1:0] node1414;
	wire [4-1:0] node1415;
	wire [4-1:0] node1417;
	wire [4-1:0] node1419;
	wire [4-1:0] node1425;
	wire [4-1:0] node1426;
	wire [4-1:0] node1427;
	wire [4-1:0] node1429;
	wire [4-1:0] node1431;
	wire [4-1:0] node1435;
	wire [4-1:0] node1437;
	wire [4-1:0] node1438;
	wire [4-1:0] node1440;
	wire [4-1:0] node1442;
	wire [4-1:0] node1444;
	wire [4-1:0] node1448;
	wire [4-1:0] node1449;
	wire [4-1:0] node1450;
	wire [4-1:0] node1452;
	wire [4-1:0] node1453;
	wire [4-1:0] node1455;
	wire [4-1:0] node1457;
	wire [4-1:0] node1459;
	wire [4-1:0] node1462;
	wire [4-1:0] node1463;
	wire [4-1:0] node1465;
	wire [4-1:0] node1467;
	wire [4-1:0] node1471;
	wire [4-1:0] node1473;
	wire [4-1:0] node1474;
	wire [4-1:0] node1476;
	wire [4-1:0] node1480;
	wire [4-1:0] node1481;
	wire [4-1:0] node1482;
	wire [4-1:0] node1483;
	wire [4-1:0] node1485;
	wire [4-1:0] node1487;
	wire [4-1:0] node1488;
	wire [4-1:0] node1492;
	wire [4-1:0] node1494;
	wire [4-1:0] node1496;
	wire [4-1:0] node1498;
	wire [4-1:0] node1501;
	wire [4-1:0] node1502;
	wire [4-1:0] node1504;
	wire [4-1:0] node1508;
	wire [4-1:0] node1509;
	wire [4-1:0] node1510;
	wire [4-1:0] node1512;
	wire [4-1:0] node1514;
	wire [4-1:0] node1516;
	wire [4-1:0] node1519;
	wire [4-1:0] node1520;
	wire [4-1:0] node1522;
	wire [4-1:0] node1524;
	wire [4-1:0] node1528;
	wire [4-1:0] node1529;
	wire [4-1:0] node1531;
	wire [4-1:0] node1534;
	wire [4-1:0] node1535;
	wire [4-1:0] node1537;
	wire [4-1:0] node1539;
	wire [4-1:0] node1542;
	wire [4-1:0] node1544;
	wire [4-1:0] node1546;

	assign outp = (inp[10]) ? node556 : node1;
		assign node1 = (inp[5]) ? node223 : node2;
			assign node2 = (inp[4]) ? node100 : node3;
				assign node3 = (inp[14]) ? node61 : node4;
					assign node4 = (inp[13]) ? node6 : 4'b1111;
						assign node6 = (inp[12]) ? node32 : node7;
							assign node7 = (inp[2]) ? node9 : 4'b1111;
								assign node9 = (inp[9]) ? node11 : 4'b1111;
									assign node11 = (inp[8]) ? node13 : 4'b1111;
										assign node13 = (inp[7]) ? node23 : node14;
											assign node14 = (inp[1]) ? node16 : 4'b1111;
												assign node16 = (inp[15]) ? node18 : 4'b1111;
													assign node18 = (inp[11]) ? node20 : 4'b1111;
														assign node20 = (inp[6]) ? 4'b1101 : 4'b1111;
											assign node23 = (inp[6]) ? 4'b1101 : node24;
												assign node24 = (inp[15]) ? node26 : 4'b1111;
													assign node26 = (inp[11]) ? node28 : 4'b1111;
														assign node28 = (inp[1]) ? 4'b1101 : 4'b1111;
							assign node32 = (inp[2]) ? 4'b1101 : node33;
								assign node33 = (inp[6]) ? node47 : node34;
									assign node34 = (inp[9]) ? node36 : 4'b1111;
										assign node36 = (inp[8]) ? 4'b1101 : node37;
											assign node37 = (inp[7]) ? node39 : 4'b1111;
												assign node39 = (inp[11]) ? node41 : 4'b1111;
													assign node41 = (inp[15]) ? node43 : 4'b1111;
														assign node43 = (inp[1]) ? 4'b1101 : 4'b1111;
									assign node47 = (inp[9]) ? 4'b1101 : node48;
										assign node48 = (inp[7]) ? 4'b1101 : node49;
											assign node49 = (inp[8]) ? 4'b1101 : node50;
												assign node50 = (inp[1]) ? node52 : 4'b1111;
													assign node52 = (inp[15]) ? node54 : 4'b1111;
														assign node54 = (inp[11]) ? 4'b1101 : 4'b1111;
					assign node61 = (inp[13]) ? node73 : node62;
						assign node62 = (inp[12]) ? node64 : 4'b1101;
							assign node64 = (inp[9]) ? node66 : 4'b1101;
								assign node66 = (inp[2]) ? node68 : 4'b1101;
									assign node68 = (inp[8]) ? node70 : 4'b1101;
										assign node70 = (inp[6]) ? 4'b1011 : 4'b1101;
						assign node73 = (inp[12]) ? node87 : node74;
							assign node74 = (inp[8]) ? node76 : 4'b1101;
								assign node76 = (inp[2]) ? node78 : 4'b1101;
									assign node78 = (inp[9]) ? node80 : 4'b1101;
										assign node80 = (inp[6]) ? 4'b1011 : node81;
											assign node81 = (inp[15]) ? node83 : 4'b1101;
												assign node83 = (inp[7]) ? 4'b1111 : 4'b1101;
							assign node87 = (inp[6]) ? 4'b1011 : node88;
								assign node88 = (inp[9]) ? 4'b1111 : node89;
									assign node89 = (inp[2]) ? 4'b1111 : node90;
										assign node90 = (inp[8]) ? node92 : 4'b1101;
											assign node92 = (inp[15]) ? node94 : 4'b1101;
												assign node94 = (inp[7]) ? 4'b1111 : 4'b1101;
				assign node100 = (inp[6]) ? node164 : node101;
					assign node101 = (inp[14]) ? node137 : node102;
						assign node102 = (inp[12]) ? node120 : node103;
							assign node103 = (inp[2]) ? node105 : 4'b1011;
								assign node105 = (inp[13]) ? node107 : 4'b1011;
									assign node107 = (inp[9]) ? node109 : 4'b1011;
										assign node109 = (inp[8]) ? 4'b1001 : node110;
											assign node110 = (inp[7]) ? 4'b1001 : node111;
												assign node111 = (inp[11]) ? node113 : 4'b1011;
													assign node113 = (inp[1]) ? node115 : 4'b1011;
														assign node115 = (inp[15]) ? 4'b1001 : 4'b1011;
							assign node120 = (inp[13]) ? 4'b1001 : node121;
								assign node121 = (inp[2]) ? node123 : 4'b1011;
									assign node123 = (inp[9]) ? 4'b1001 : node124;
										assign node124 = (inp[8]) ? node126 : 4'b1011;
											assign node126 = (inp[7]) ? 4'b1001 : node127;
												assign node127 = (inp[1]) ? node129 : 4'b1011;
													assign node129 = (inp[11]) ? node131 : 4'b1011;
														assign node131 = (inp[15]) ? 4'b1001 : 4'b1011;
						assign node137 = (inp[12]) ? node151 : node138;
							assign node138 = (inp[2]) ? node140 : 4'b1001;
								assign node140 = (inp[13]) ? node142 : 4'b1001;
									assign node142 = (inp[9]) ? 4'b1011 : node143;
										assign node143 = (inp[7]) ? node145 : 4'b1001;
											assign node145 = (inp[15]) ? node147 : 4'b1001;
												assign node147 = (inp[8]) ? 4'b1011 : 4'b1001;
							assign node151 = (inp[13]) ? 4'b1011 : node152;
								assign node152 = (inp[2]) ? 4'b1011 : node153;
									assign node153 = (inp[7]) ? node155 : 4'b1001;
										assign node155 = (inp[8]) ? node157 : 4'b1001;
											assign node157 = (inp[9]) ? node159 : 4'b1001;
												assign node159 = (inp[15]) ? 4'b1011 : 4'b1001;
					assign node164 = (inp[14]) ? node200 : node165;
						assign node165 = (inp[12]) ? node183 : node166;
							assign node166 = (inp[2]) ? node168 : 4'b1011;
								assign node168 = (inp[13]) ? node170 : 4'b1011;
									assign node170 = (inp[9]) ? 4'b1001 : node171;
										assign node171 = (inp[8]) ? 4'b1001 : node172;
											assign node172 = (inp[7]) ? node174 : 4'b1011;
												assign node174 = (inp[1]) ? node176 : 4'b1011;
													assign node176 = (inp[15]) ? node178 : 4'b1011;
														assign node178 = (inp[11]) ? 4'b1001 : 4'b1011;
							assign node183 = (inp[2]) ? 4'b1001 : node184;
								assign node184 = (inp[13]) ? 4'b1001 : node185;
									assign node185 = (inp[9]) ? 4'b1001 : node186;
										assign node186 = (inp[7]) ? node188 : 4'b1011;
											assign node188 = (inp[15]) ? node190 : 4'b1011;
												assign node190 = (inp[11]) ? node192 : 4'b1011;
													assign node192 = (inp[1]) ? node194 : 4'b1011;
														assign node194 = (inp[8]) ? 4'b1001 : 4'b1011;
						assign node200 = (inp[12]) ? node206 : node201;
							assign node201 = (inp[2]) ? node203 : 4'b1001;
								assign node203 = (inp[13]) ? 4'b1111 : 4'b1001;
							assign node206 = (inp[2]) ? node208 : 4'b1110;
								assign node208 = (inp[13]) ? node210 : 4'b1110;
									assign node210 = (inp[9]) ? 4'b1100 : node211;
										assign node211 = (inp[1]) ? node213 : 4'b1110;
											assign node213 = (inp[8]) ? node215 : 4'b1110;
												assign node215 = (inp[15]) ? node217 : 4'b1110;
													assign node217 = (inp[11]) ? node219 : 4'b1110;
														assign node219 = (inp[7]) ? 4'b1100 : 4'b1110;
			assign node223 = (inp[12]) ? node375 : node224;
				assign node224 = (inp[6]) ? node296 : node225;
					assign node225 = (inp[13]) ? node277 : node226;
						assign node226 = (inp[4]) ? node254 : node227;
							assign node227 = (inp[14]) ? node239 : node228;
								assign node228 = (inp[2]) ? node230 : 4'b1001;
									assign node230 = (inp[9]) ? 4'b1011 : node231;
										assign node231 = (inp[8]) ? node233 : 4'b1001;
											assign node233 = (inp[7]) ? node235 : 4'b1001;
												assign node235 = (inp[15]) ? 4'b1011 : 4'b1001;
								assign node239 = (inp[8]) ? 4'b1001 : node240;
									assign node240 = (inp[9]) ? 4'b1001 : node241;
										assign node241 = (inp[2]) ? 4'b1001 : node242;
											assign node242 = (inp[15]) ? node244 : 4'b1011;
												assign node244 = (inp[1]) ? node246 : 4'b1011;
													assign node246 = (inp[11]) ? node248 : 4'b1011;
														assign node248 = (inp[7]) ? 4'b1001 : 4'b1011;
							assign node254 = (inp[14]) ? node262 : node255;
								assign node255 = (inp[2]) ? node257 : 4'b1101;
									assign node257 = (inp[9]) ? node259 : 4'b1101;
										assign node259 = (inp[8]) ? 4'b1011 : 4'b1101;
								assign node262 = (inp[9]) ? 4'b1001 : node263;
									assign node263 = (inp[2]) ? 4'b1001 : node264;
										assign node264 = (inp[8]) ? node266 : 4'b1011;
											assign node266 = (inp[7]) ? 4'b1001 : node267;
												assign node267 = (inp[1]) ? node269 : 4'b1011;
													assign node269 = (inp[15]) ? node271 : 4'b1011;
														assign node271 = (inp[11]) ? 4'b1001 : 4'b1011;
						assign node277 = (inp[2]) ? node291 : node278;
							assign node278 = (inp[14]) ? node280 : 4'b1011;
								assign node280 = (inp[9]) ? node282 : 4'b1001;
									assign node282 = (inp[8]) ? node284 : 4'b1001;
										assign node284 = (inp[4]) ? node286 : 4'b1001;
											assign node286 = (inp[15]) ? node288 : 4'b1001;
												assign node288 = (inp[7]) ? 4'b1011 : 4'b1001;
							assign node291 = (inp[4]) ? 4'b1011 : node292;
								assign node292 = (inp[14]) ? 4'b1111 : 4'b1011;
					assign node296 = (inp[14]) ? node332 : node297;
						assign node297 = (inp[4]) ? node315 : node298;
							assign node298 = (inp[13]) ? 4'b1101 : node299;
								assign node299 = (inp[2]) ? node301 : 4'b1111;
									assign node301 = (inp[9]) ? node303 : 4'b1111;
										assign node303 = (inp[8]) ? 4'b1101 : node304;
											assign node304 = (inp[7]) ? node306 : 4'b1111;
												assign node306 = (inp[15]) ? node308 : 4'b1111;
													assign node308 = (inp[11]) ? node310 : 4'b1111;
														assign node310 = (inp[1]) ? 4'b1101 : 4'b1111;
							assign node315 = (inp[13]) ? 4'b1001 : node316;
								assign node316 = (inp[2]) ? node318 : 4'b1011;
									assign node318 = (inp[9]) ? 4'b1001 : node319;
										assign node319 = (inp[7]) ? node321 : 4'b1011;
											assign node321 = (inp[15]) ? node323 : 4'b1011;
												assign node323 = (inp[1]) ? node325 : 4'b1011;
													assign node325 = (inp[11]) ? node327 : 4'b1011;
														assign node327 = (inp[8]) ? 4'b1001 : 4'b1011;
						assign node332 = (inp[4]) ? node360 : node333;
							assign node333 = (inp[2]) ? node345 : node334;
								assign node334 = (inp[13]) ? 4'b1111 : node335;
									assign node335 = (inp[9]) ? 4'b1111 : node336;
										assign node336 = (inp[8]) ? node338 : 4'b1101;
											assign node338 = (inp[7]) ? node340 : 4'b1101;
												assign node340 = (inp[15]) ? 4'b1111 : 4'b1101;
								assign node345 = (inp[13]) ? node347 : 4'b1111;
									assign node347 = (inp[7]) ? 4'b1101 : node348;
										assign node348 = (inp[9]) ? 4'b1101 : node349;
											assign node349 = (inp[8]) ? 4'b1101 : node350;
												assign node350 = (inp[1]) ? node352 : 4'b1111;
													assign node352 = (inp[11]) ? node354 : 4'b1111;
														assign node354 = (inp[15]) ? 4'b1101 : 4'b1111;
							assign node360 = (inp[13]) ? node362 : 4'b1110;
								assign node362 = (inp[2]) ? 4'b1100 : node363;
									assign node363 = (inp[9]) ? 4'b1100 : node364;
										assign node364 = (inp[1]) ? node366 : 4'b1110;
											assign node366 = (inp[8]) ? node368 : 4'b1110;
												assign node368 = (inp[11]) ? node370 : 4'b1110;
													assign node370 = (inp[7]) ? 4'b1100 : 4'b1110;
				assign node375 = (inp[6]) ? node469 : node376;
					assign node376 = (inp[14]) ? node436 : node377;
						assign node377 = (inp[4]) ? node409 : node378;
							assign node378 = (inp[9]) ? node396 : node379;
								assign node379 = (inp[2]) ? node383 : node380;
									assign node380 = (inp[13]) ? 4'b1110 : 4'b1100;
									assign node383 = (inp[8]) ? node385 : 4'b1110;
										assign node385 = (inp[13]) ? node387 : 4'b1110;
											assign node387 = (inp[7]) ? 4'b1100 : node388;
												assign node388 = (inp[11]) ? node390 : 4'b1110;
													assign node390 = (inp[15]) ? node392 : 4'b1110;
														assign node392 = (inp[1]) ? 4'b1100 : 4'b1110;
								assign node396 = (inp[13]) ? node406 : node397;
									assign node397 = (inp[2]) ? 4'b1110 : node398;
										assign node398 = (inp[7]) ? node400 : 4'b1100;
											assign node400 = (inp[15]) ? node402 : 4'b1100;
												assign node402 = (inp[8]) ? 4'b1110 : 4'b1100;
									assign node406 = (inp[2]) ? 4'b1100 : 4'b1110;
							assign node409 = (inp[13]) ? node425 : node410;
								assign node410 = (inp[2]) ? node412 : 4'b1110;
									assign node412 = (inp[9]) ? 4'b1100 : node413;
										assign node413 = (inp[8]) ? 4'b1100 : node414;
											assign node414 = (inp[7]) ? node416 : 4'b1110;
												assign node416 = (inp[11]) ? node418 : 4'b1110;
													assign node418 = (inp[1]) ? node420 : 4'b1110;
														assign node420 = (inp[15]) ? 4'b1100 : 4'b1110;
								assign node425 = (inp[2]) ? node427 : 4'b1100;
									assign node427 = (inp[9]) ? 4'b1110 : node428;
										assign node428 = (inp[8]) ? node430 : 4'b1100;
											assign node430 = (inp[15]) ? node432 : 4'b1100;
												assign node432 = (inp[7]) ? 4'b1110 : 4'b1100;
						assign node436 = (inp[13]) ? node460 : node437;
							assign node437 = (inp[4]) ? node445 : node438;
								assign node438 = (inp[8]) ? node440 : 4'b1100;
									assign node440 = (inp[2]) ? node442 : 4'b1100;
										assign node442 = (inp[9]) ? 4'b1010 : 4'b1100;
								assign node445 = (inp[9]) ? node447 : 4'b1110;
									assign node447 = (inp[2]) ? node449 : 4'b1110;
										assign node449 = (inp[8]) ? 4'b1100 : node450;
											assign node450 = (inp[7]) ? 4'b1100 : node451;
												assign node451 = (inp[11]) ? node453 : 4'b1110;
													assign node453 = (inp[1]) ? node455 : 4'b1110;
														assign node455 = (inp[15]) ? 4'b1100 : 4'b1110;
							assign node460 = (inp[4]) ? node462 : 4'b1010;
								assign node462 = (inp[8]) ? node464 : 4'b1100;
									assign node464 = (inp[9]) ? node466 : 4'b1100;
										assign node466 = (inp[2]) ? 4'b1010 : 4'b1100;
					assign node469 = (inp[13]) ? node527 : node470;
						assign node470 = (inp[4]) ? node502 : node471;
							assign node471 = (inp[2]) ? 4'b1000 : node472;
								assign node472 = (inp[14]) ? node486 : node473;
									assign node473 = (inp[8]) ? 4'b1000 : node474;
										assign node474 = (inp[9]) ? 4'b1000 : node475;
											assign node475 = (inp[7]) ? 4'b1000 : node476;
												assign node476 = (inp[15]) ? node478 : 4'b1010;
													assign node478 = (inp[11]) ? node480 : 4'b1010;
														assign node480 = (inp[1]) ? 4'b1000 : 4'b1010;
									assign node486 = (inp[9]) ? node488 : 4'b1010;
										assign node488 = (inp[8]) ? 4'b1000 : node489;
											assign node489 = (inp[11]) ? node491 : 4'b1010;
												assign node491 = (inp[0]) ? 4'b1010 : node492;
													assign node492 = (inp[3]) ? 4'b1010 : node493;
														assign node493 = (inp[1]) ? node495 : 4'b1010;
															assign node495 = (inp[7]) ? 4'b1000 : 4'b1010;
							assign node502 = (inp[8]) ? node504 : 4'b1010;
								assign node504 = (inp[2]) ? node506 : 4'b1010;
									assign node506 = (inp[9]) ? node508 : 4'b1010;
										assign node508 = (inp[14]) ? node518 : node509;
											assign node509 = (inp[7]) ? 4'b1000 : node510;
												assign node510 = (inp[15]) ? node512 : 4'b1010;
													assign node512 = (inp[11]) ? node514 : 4'b1010;
														assign node514 = (inp[1]) ? 4'b1000 : 4'b1010;
											assign node518 = (inp[15]) ? node520 : 4'b1010;
												assign node520 = (inp[7]) ? node522 : 4'b1010;
													assign node522 = (inp[11]) ? node524 : 4'b1010;
														assign node524 = (inp[1]) ? 4'b1000 : 4'b1010;
						assign node527 = (inp[4]) ? node543 : node528;
							assign node528 = (inp[2]) ? node540 : node529;
								assign node529 = (inp[14]) ? 4'b1000 : node530;
									assign node530 = (inp[9]) ? 4'b1010 : node531;
										assign node531 = (inp[15]) ? node533 : 4'b1000;
											assign node533 = (inp[7]) ? node535 : 4'b1000;
												assign node535 = (inp[8]) ? 4'b1010 : 4'b1000;
								assign node540 = (inp[14]) ? 4'b1110 : 4'b1010;
							assign node543 = (inp[8]) ? node545 : 4'b1000;
								assign node545 = (inp[7]) ? node547 : 4'b1000;
									assign node547 = (inp[15]) ? node549 : 4'b1000;
										assign node549 = (inp[9]) ? node551 : 4'b1000;
											assign node551 = (inp[14]) ? 4'b1000 : node552;
												assign node552 = (inp[2]) ? 4'b1010 : 4'b1000;
		assign node556 = (inp[5]) ? node942 : node557;
			assign node557 = (inp[4]) ? node687 : node558;
				assign node558 = (inp[6]) ? node632 : node559;
					assign node559 = (inp[14]) ? node597 : node560;
						assign node560 = (inp[13]) ? node578 : node561;
							assign node561 = (inp[2]) ? 4'b1100 : node562;
								assign node562 = (inp[12]) ? node564 : 4'b1100;
									assign node564 = (inp[9]) ? node566 : 4'b1110;
										assign node566 = (inp[8]) ? 4'b1100 : node567;
											assign node567 = (inp[7]) ? 4'b1100 : node568;
												assign node568 = (inp[11]) ? node570 : 4'b1110;
													assign node570 = (inp[15]) ? node572 : 4'b1110;
														assign node572 = (inp[1]) ? 4'b1100 : 4'b1110;
							assign node578 = (inp[2]) ? node590 : node579;
								assign node579 = (inp[15]) ? node581 : 4'b1100;
									assign node581 = (inp[8]) ? node583 : 4'b1100;
										assign node583 = (inp[7]) ? node585 : 4'b1100;
											assign node585 = (inp[12]) ? 4'b1100 : node586;
												assign node586 = (inp[9]) ? 4'b1110 : 4'b1100;
								assign node590 = (inp[12]) ? node592 : 4'b1110;
									assign node592 = (inp[9]) ? node594 : 4'b1100;
										assign node594 = (inp[8]) ? 4'b1010 : 4'b1100;
						assign node597 = (inp[12]) ? node615 : node598;
							assign node598 = (inp[13]) ? node600 : 4'b1110;
								assign node600 = (inp[9]) ? 4'b1100 : node601;
									assign node601 = (inp[2]) ? 4'b1100 : node602;
										assign node602 = (inp[8]) ? node604 : 4'b1110;
											assign node604 = (inp[7]) ? 4'b1100 : node605;
												assign node605 = (inp[11]) ? node607 : 4'b1110;
													assign node607 = (inp[15]) ? node609 : 4'b1110;
														assign node609 = (inp[1]) ? 4'b1100 : 4'b1110;
							assign node615 = (inp[13]) ? node617 : 4'b1010;
								assign node617 = (inp[2]) ? 4'b1000 : node618;
									assign node618 = (inp[9]) ? node620 : 4'b1010;
										assign node620 = (inp[8]) ? node622 : 4'b1010;
											assign node622 = (inp[7]) ? 4'b1000 : node623;
												assign node623 = (inp[15]) ? node625 : 4'b1010;
													assign node625 = (inp[1]) ? node627 : 4'b1010;
														assign node627 = (inp[11]) ? 4'b1000 : 4'b1010;
					assign node632 = (inp[14]) ? node654 : node633;
						assign node633 = (inp[13]) ? 4'b1010 : node634;
							assign node634 = (inp[12]) ? node642 : node635;
								assign node635 = (inp[9]) ? node637 : 4'b1100;
									assign node637 = (inp[8]) ? node639 : 4'b1100;
										assign node639 = (inp[2]) ? 4'b1010 : 4'b1100;
								assign node642 = (inp[9]) ? node644 : 4'b1000;
									assign node644 = (inp[8]) ? node646 : 4'b1000;
										assign node646 = (inp[2]) ? node648 : 4'b1000;
											assign node648 = (inp[15]) ? node650 : 4'b1000;
												assign node650 = (inp[7]) ? 4'b1010 : 4'b1000;
						assign node654 = (inp[13]) ? 4'b1000 : node655;
							assign node655 = (inp[2]) ? node671 : node656;
								assign node656 = (inp[11]) ? node658 : 4'b1010;
									assign node658 = (inp[9]) ? node660 : 4'b1010;
										assign node660 = (inp[15]) ? node662 : 4'b1010;
											assign node662 = (inp[8]) ? node664 : 4'b1010;
												assign node664 = (inp[12]) ? node666 : 4'b1010;
													assign node666 = (inp[7]) ? node668 : 4'b1010;
														assign node668 = (inp[1]) ? 4'b1000 : 4'b1010;
								assign node671 = (inp[9]) ? 4'b1000 : node672;
									assign node672 = (inp[7]) ? 4'b1000 : node673;
										assign node673 = (inp[12]) ? 4'b1000 : node674;
											assign node674 = (inp[8]) ? 4'b1000 : node675;
												assign node675 = (inp[15]) ? node677 : 4'b1010;
													assign node677 = (inp[11]) ? node679 : 4'b1010;
														assign node679 = (inp[1]) ? 4'b1000 : 4'b1010;
				assign node687 = (inp[12]) ? node869 : node688;
					assign node688 = (inp[6]) ? node838 : node689;
						assign node689 = (inp[14]) ? node833 : node690;
							assign node690 = (inp[8]) ? node710 : node691;
								assign node691 = (inp[9]) ? node697 : node692;
									assign node692 = (inp[2]) ? 4'b1010 : node693;
										assign node693 = (inp[13]) ? 4'b1010 : 4'b1000;
									assign node697 = (inp[2]) ? node699 : 4'b1010;
										assign node699 = (inp[15]) ? node701 : 4'b1010;
											assign node701 = (inp[1]) ? node703 : 4'b1010;
												assign node703 = (inp[7]) ? node705 : 4'b1010;
													assign node705 = (inp[11]) ? node707 : 4'b1010;
														assign node707 = (inp[13]) ? 4'b1000 : 4'b1010;
								assign node710 = (inp[7]) ? node782 : node711;
									assign node711 = (inp[1]) ? node747 : node712;
										assign node712 = (inp[0]) ? node724 : node713;
											assign node713 = (inp[2]) ? node719 : node714;
												assign node714 = (inp[13]) ? 4'b1010 : node715;
													assign node715 = (inp[9]) ? 4'b1010 : 4'b1000;
												assign node719 = (inp[13]) ? node721 : 4'b1010;
													assign node721 = (inp[9]) ? 4'b1000 : 4'b1010;
											assign node724 = (inp[11]) ? node736 : node725;
												assign node725 = (inp[2]) ? node731 : node726;
													assign node726 = (inp[9]) ? 4'b1010 : node727;
														assign node727 = (inp[13]) ? 4'b1010 : 4'b1000;
													assign node731 = (inp[9]) ? node733 : 4'b1010;
														assign node733 = (inp[13]) ? 4'b1000 : 4'b1010;
												assign node736 = (inp[2]) ? node742 : node737;
													assign node737 = (inp[9]) ? 4'b1010 : node738;
														assign node738 = (inp[13]) ? 4'b1010 : 4'b1000;
													assign node742 = (inp[9]) ? node744 : 4'b1010;
														assign node744 = (inp[13]) ? 4'b1000 : 4'b1010;
										assign node747 = (inp[0]) ? node759 : node748;
											assign node748 = (inp[2]) ? node754 : node749;
												assign node749 = (inp[9]) ? 4'b1010 : node750;
													assign node750 = (inp[13]) ? 4'b1010 : 4'b1000;
												assign node754 = (inp[9]) ? node756 : 4'b1010;
													assign node756 = (inp[13]) ? 4'b1000 : 4'b1010;
											assign node759 = (inp[3]) ? node771 : node760;
												assign node760 = (inp[9]) ? node766 : node761;
													assign node761 = (inp[2]) ? 4'b1010 : node762;
														assign node762 = (inp[13]) ? 4'b1010 : 4'b1000;
													assign node766 = (inp[2]) ? node768 : 4'b1010;
														assign node768 = (inp[13]) ? 4'b1000 : 4'b1010;
												assign node771 = (inp[2]) ? node777 : node772;
													assign node772 = (inp[9]) ? 4'b1010 : node773;
														assign node773 = (inp[13]) ? 4'b1010 : 4'b1000;
													assign node777 = (inp[9]) ? node779 : 4'b1010;
														assign node779 = (inp[13]) ? 4'b1000 : 4'b1010;
									assign node782 = (inp[15]) ? node826 : node783;
										assign node783 = (inp[3]) ? node795 : node784;
											assign node784 = (inp[9]) ? node790 : node785;
												assign node785 = (inp[2]) ? 4'b1010 : node786;
													assign node786 = (inp[13]) ? 4'b1010 : 4'b1000;
												assign node790 = (inp[2]) ? node792 : 4'b1010;
													assign node792 = (inp[13]) ? 4'b1000 : 4'b1010;
											assign node795 = (inp[1]) ? node815 : node796;
												assign node796 = (inp[0]) ? node806 : node797;
													assign node797 = (inp[13]) ? node803 : node798;
														assign node798 = (inp[2]) ? 4'b1010 : node799;
															assign node799 = (inp[9]) ? 4'b1010 : 4'b1000;
														assign node803 = (inp[9]) ? 4'b1000 : 4'b1010;
													assign node806 = (inp[2]) ? node812 : node807;
														assign node807 = (inp[9]) ? 4'b1010 : node808;
															assign node808 = (inp[13]) ? 4'b1010 : 4'b1000;
														assign node812 = (inp[9]) ? 4'b1000 : 4'b1010;
												assign node815 = (inp[2]) ? node821 : node816;
													assign node816 = (inp[13]) ? 4'b1010 : node817;
														assign node817 = (inp[9]) ? 4'b1010 : 4'b1000;
													assign node821 = (inp[13]) ? node823 : 4'b1010;
														assign node823 = (inp[9]) ? 4'b1000 : 4'b1010;
										assign node826 = (inp[13]) ? node828 : 4'b1010;
											assign node828 = (inp[2]) ? node830 : 4'b1010;
												assign node830 = (inp[9]) ? 4'b1000 : 4'b1010;
							assign node833 = (inp[13]) ? node835 : 4'b1000;
								assign node835 = (inp[2]) ? 4'b1110 : 4'b1000;
						assign node838 = (inp[13]) ? node852 : node839;
							assign node839 = (inp[14]) ? node841 : 4'b1110;
								assign node841 = (inp[2]) ? node843 : 4'b1100;
									assign node843 = (inp[9]) ? 4'b1110 : node844;
										assign node844 = (inp[8]) ? node846 : 4'b1100;
											assign node846 = (inp[15]) ? node848 : 4'b1100;
												assign node848 = (inp[7]) ? 4'b1110 : 4'b1100;
							assign node852 = (inp[14]) ? 4'b1110 : node853;
								assign node853 = (inp[8]) ? 4'b1100 : node854;
									assign node854 = (inp[2]) ? 4'b1100 : node855;
										assign node855 = (inp[9]) ? 4'b1100 : node856;
											assign node856 = (inp[1]) ? node858 : 4'b1110;
												assign node858 = (inp[15]) ? node860 : 4'b1110;
													assign node860 = (inp[7]) ? node862 : 4'b1110;
														assign node862 = (inp[11]) ? 4'b1100 : 4'b1110;
					assign node869 = (inp[6]) ? node901 : node870;
						assign node870 = (inp[14]) ? node888 : node871;
							assign node871 = (inp[13]) ? node873 : 4'b1111;
								assign node873 = (inp[2]) ? 4'b1101 : node874;
									assign node874 = (inp[9]) ? node876 : 4'b1111;
										assign node876 = (inp[1]) ? node878 : 4'b1111;
											assign node878 = (inp[11]) ? node880 : 4'b1111;
												assign node880 = (inp[7]) ? node882 : 4'b1111;
													assign node882 = (inp[8]) ? node884 : 4'b1111;
														assign node884 = (inp[15]) ? 4'b1101 : 4'b1111;
							assign node888 = (inp[13]) ? 4'b1111 : node889;
								assign node889 = (inp[2]) ? node891 : 4'b1101;
									assign node891 = (inp[7]) ? node893 : 4'b1101;
										assign node893 = (inp[8]) ? node895 : 4'b1101;
											assign node895 = (inp[9]) ? node897 : 4'b1101;
												assign node897 = (inp[15]) ? 4'b1111 : 4'b1101;
						assign node901 = (inp[14]) ? node925 : node902;
							assign node902 = (inp[13]) ? node918 : node903;
								assign node903 = (inp[2]) ? 4'b1101 : node904;
									assign node904 = (inp[9]) ? node906 : 4'b1111;
										assign node906 = (inp[8]) ? node908 : 4'b1111;
											assign node908 = (inp[7]) ? 4'b1101 : node909;
												assign node909 = (inp[1]) ? node911 : 4'b1111;
													assign node911 = (inp[15]) ? node913 : 4'b1111;
														assign node913 = (inp[11]) ? 4'b1101 : 4'b1111;
								assign node918 = (inp[2]) ? node920 : 4'b1101;
									assign node920 = (inp[9]) ? node922 : 4'b1101;
										assign node922 = (inp[8]) ? 4'b1011 : 4'b1101;
							assign node925 = (inp[13]) ? node927 : 4'b1011;
								assign node927 = (inp[2]) ? 4'b1001 : node928;
									assign node928 = (inp[9]) ? node930 : 4'b1011;
										assign node930 = (inp[8]) ? 4'b1001 : node931;
											assign node931 = (inp[7]) ? 4'b1001 : node932;
												assign node932 = (inp[15]) ? node934 : 4'b1011;
													assign node934 = (inp[1]) ? node936 : 4'b1011;
														assign node936 = (inp[11]) ? 4'b1001 : 4'b1011;
			assign node942 = (inp[12]) ? node1150 : node943;
				assign node943 = (inp[6]) ? node1047 : node944;
					assign node944 = (inp[13]) ? node1006 : node945;
						assign node945 = (inp[4]) ? node971 : node946;
							assign node946 = (inp[8]) ? node948 : 4'b0111;
								assign node948 = (inp[9]) ? node950 : 4'b0111;
									assign node950 = (inp[2]) ? node952 : 4'b0111;
										assign node952 = (inp[14]) ? node962 : node953;
											assign node953 = (inp[15]) ? node955 : 4'b0111;
												assign node955 = (inp[1]) ? node957 : 4'b0111;
													assign node957 = (inp[11]) ? node959 : 4'b0111;
														assign node959 = (inp[7]) ? 4'b0101 : 4'b0111;
											assign node962 = (inp[7]) ? 4'b0101 : node963;
												assign node963 = (inp[15]) ? node965 : 4'b0111;
													assign node965 = (inp[1]) ? node967 : 4'b0111;
														assign node967 = (inp[11]) ? 4'b0101 : 4'b0111;
							assign node971 = (inp[2]) ? node999 : node972;
								assign node972 = (inp[14]) ? node986 : node973;
									assign node973 = (inp[9]) ? node975 : 4'b0111;
										assign node975 = (inp[8]) ? 4'b0101 : node976;
											assign node976 = (inp[11]) ? node978 : 4'b0111;
												assign node978 = (inp[7]) ? node980 : 4'b0111;
													assign node980 = (inp[1]) ? node982 : 4'b0111;
														assign node982 = (inp[15]) ? 4'b0101 : 4'b0111;
									assign node986 = (inp[7]) ? 4'b0101 : node987;
										assign node987 = (inp[8]) ? 4'b0101 : node988;
											assign node988 = (inp[9]) ? 4'b0101 : node989;
												assign node989 = (inp[11]) ? node991 : 4'b0111;
													assign node991 = (inp[15]) ? node993 : 4'b0111;
														assign node993 = (inp[1]) ? 4'b0101 : 4'b0111;
								assign node999 = (inp[8]) ? node1001 : 4'b0101;
									assign node1001 = (inp[9]) ? node1003 : 4'b0101;
										assign node1003 = (inp[14]) ? 4'b0011 : 4'b0101;
						assign node1006 = (inp[4]) ? node1020 : node1007;
							assign node1007 = (inp[8]) ? node1009 : 4'b0101;
								assign node1009 = (inp[9]) ? node1011 : 4'b0101;
									assign node1011 = (inp[2]) ? node1013 : 4'b0101;
										assign node1013 = (inp[14]) ? 4'b0011 : node1014;
											assign node1014 = (inp[15]) ? node1016 : 4'b0101;
												assign node1016 = (inp[7]) ? 4'b0111 : 4'b0101;
							assign node1020 = (inp[14]) ? node1032 : node1021;
								assign node1021 = (inp[2]) ? 4'b0111 : node1022;
									assign node1022 = (inp[9]) ? 4'b0111 : node1023;
										assign node1023 = (inp[8]) ? node1025 : 4'b0101;
											assign node1025 = (inp[15]) ? node1027 : 4'b0101;
												assign node1027 = (inp[7]) ? 4'b0111 : 4'b0101;
								assign node1032 = (inp[2]) ? node1034 : 4'b0011;
									assign node1034 = (inp[9]) ? 4'b0001 : node1035;
										assign node1035 = (inp[8]) ? node1037 : 4'b0011;
											assign node1037 = (inp[7]) ? 4'b0001 : node1038;
												assign node1038 = (inp[15]) ? node1040 : 4'b0011;
													assign node1040 = (inp[1]) ? node1042 : 4'b0011;
														assign node1042 = (inp[11]) ? 4'b0001 : 4'b0011;
					assign node1047 = (inp[14]) ? node1103 : node1048;
						assign node1048 = (inp[13]) ? node1076 : node1049;
							assign node1049 = (inp[4]) ? node1065 : node1050;
								assign node1050 = (inp[2]) ? node1052 : 4'b0011;
									assign node1052 = (inp[9]) ? node1054 : 4'b0011;
										assign node1054 = (inp[8]) ? 4'b0001 : node1055;
											assign node1055 = (inp[7]) ? 4'b0001 : node1056;
												assign node1056 = (inp[11]) ? node1058 : 4'b0011;
													assign node1058 = (inp[1]) ? node1060 : 4'b0011;
														assign node1060 = (inp[15]) ? 4'b0001 : 4'b0011;
								assign node1065 = (inp[2]) ? 4'b0011 : node1066;
									assign node1066 = (inp[8]) ? node1068 : 4'b0001;
										assign node1068 = (inp[7]) ? node1070 : 4'b0001;
											assign node1070 = (inp[15]) ? node1072 : 4'b0001;
												assign node1072 = (inp[9]) ? 4'b0011 : 4'b0001;
							assign node1076 = (inp[4]) ? node1088 : node1077;
								assign node1077 = (inp[2]) ? node1079 : 4'b0001;
									assign node1079 = (inp[9]) ? 4'b0011 : node1080;
										assign node1080 = (inp[15]) ? node1082 : 4'b0001;
											assign node1082 = (inp[7]) ? node1084 : 4'b0001;
												assign node1084 = (inp[8]) ? 4'b0011 : 4'b0001;
								assign node1088 = (inp[9]) ? 4'b0001 : node1089;
									assign node1089 = (inp[2]) ? 4'b0001 : node1090;
										assign node1090 = (inp[11]) ? node1092 : 4'b0011;
											assign node1092 = (inp[1]) ? node1094 : 4'b0011;
												assign node1094 = (inp[15]) ? node1096 : 4'b0011;
													assign node1096 = (inp[7]) ? node1098 : 4'b0011;
														assign node1098 = (inp[8]) ? 4'b0001 : 4'b0011;
						assign node1103 = (inp[4]) ? node1123 : node1104;
							assign node1104 = (inp[2]) ? node1108 : node1105;
								assign node1105 = (inp[13]) ? 4'b0001 : 4'b0011;
								assign node1108 = (inp[13]) ? 4'b0111 : node1109;
									assign node1109 = (inp[9]) ? 4'b0001 : node1110;
										assign node1110 = (inp[8]) ? 4'b0001 : node1111;
											assign node1111 = (inp[11]) ? node1113 : 4'b0011;
												assign node1113 = (inp[15]) ? node1115 : 4'b0011;
													assign node1115 = (inp[7]) ? node1117 : 4'b0011;
														assign node1117 = (inp[1]) ? 4'b0001 : 4'b0011;
							assign node1123 = (inp[2]) ? node1135 : node1124;
								assign node1124 = (inp[13]) ? node1126 : 4'b0110;
									assign node1126 = (inp[8]) ? node1128 : 4'b0100;
										assign node1128 = (inp[9]) ? node1130 : 4'b0100;
											assign node1130 = (inp[15]) ? node1132 : 4'b0100;
												assign node1132 = (inp[7]) ? 4'b0110 : 4'b0100;
								assign node1135 = (inp[13]) ? 4'b0110 : node1136;
									assign node1136 = (inp[9]) ? 4'b0100 : node1137;
										assign node1137 = (inp[7]) ? node1139 : 4'b0110;
											assign node1139 = (inp[15]) ? node1141 : 4'b0110;
												assign node1141 = (inp[1]) ? node1143 : 4'b0110;
													assign node1143 = (inp[8]) ? node1145 : 4'b0110;
														assign node1145 = (inp[11]) ? 4'b0100 : 4'b0110;
				assign node1150 = (inp[4]) ? node1294 : node1151;
					assign node1151 = (inp[14]) ? node1231 : node1152;
						assign node1152 = (inp[13]) ? node1196 : node1153;
							assign node1153 = (inp[2]) ? node1179 : node1154;
								assign node1154 = (inp[9]) ? 4'b0100 : node1155;
									assign node1155 = (inp[8]) ? node1167 : node1156;
										assign node1156 = (inp[15]) ? node1158 : 4'b0110;
											assign node1158 = (inp[7]) ? node1160 : 4'b0110;
												assign node1160 = (inp[6]) ? node1162 : 4'b0110;
													assign node1162 = (inp[11]) ? node1164 : 4'b0110;
														assign node1164 = (inp[1]) ? 4'b0100 : 4'b0110;
										assign node1167 = (inp[6]) ? 4'b0100 : node1168;
											assign node1168 = (inp[7]) ? 4'b0100 : node1169;
												assign node1169 = (inp[1]) ? node1171 : 4'b0110;
													assign node1171 = (inp[15]) ? node1173 : 4'b0110;
														assign node1173 = (inp[11]) ? 4'b0100 : 4'b0110;
								assign node1179 = (inp[9]) ? node1189 : node1180;
									assign node1180 = (inp[6]) ? node1182 : 4'b0100;
										assign node1182 = (inp[8]) ? node1184 : 4'b0100;
											assign node1184 = (inp[15]) ? node1186 : 4'b0100;
												assign node1186 = (inp[7]) ? 4'b0110 : 4'b0100;
									assign node1189 = (inp[8]) ? node1193 : node1190;
										assign node1190 = (inp[6]) ? 4'b0110 : 4'b0100;
										assign node1193 = (inp[6]) ? 4'b0110 : 4'b0010;
							assign node1196 = (inp[6]) ? node1212 : node1197;
								assign node1197 = (inp[2]) ? node1199 : 4'b0010;
									assign node1199 = (inp[9]) ? 4'b0000 : node1200;
										assign node1200 = (inp[8]) ? 4'b0000 : node1201;
											assign node1201 = (inp[7]) ? 4'b0000 : node1202;
												assign node1202 = (inp[11]) ? node1204 : 4'b0010;
													assign node1204 = (inp[15]) ? node1206 : 4'b0010;
														assign node1206 = (inp[1]) ? 4'b0000 : 4'b0010;
								assign node1212 = (inp[2]) ? node1226 : node1213;
									assign node1213 = (inp[9]) ? node1215 : 4'b0110;
										assign node1215 = (inp[8]) ? 4'b0100 : node1216;
											assign node1216 = (inp[7]) ? 4'b0100 : node1217;
												assign node1217 = (inp[1]) ? node1219 : 4'b0110;
													assign node1219 = (inp[15]) ? node1221 : 4'b0110;
														assign node1221 = (inp[11]) ? 4'b0100 : 4'b0110;
									assign node1226 = (inp[8]) ? node1228 : 4'b0100;
										assign node1228 = (inp[9]) ? 4'b0010 : 4'b0100;
						assign node1231 = (inp[2]) ? node1267 : node1232;
							assign node1232 = (inp[6]) ? node1244 : node1233;
								assign node1233 = (inp[13]) ? 4'b0000 : node1234;
									assign node1234 = (inp[9]) ? 4'b0010 : node1235;
										assign node1235 = (inp[7]) ? node1237 : 4'b0000;
											assign node1237 = (inp[8]) ? node1239 : 4'b0000;
												assign node1239 = (inp[15]) ? 4'b0010 : 4'b0000;
								assign node1244 = (inp[8]) ? node1246 : 4'b0010;
									assign node1246 = (inp[9]) ? node1248 : 4'b0010;
										assign node1248 = (inp[7]) ? node1258 : node1249;
											assign node1249 = (inp[13]) ? 4'b0010 : node1250;
												assign node1250 = (inp[1]) ? node1252 : 4'b0010;
													assign node1252 = (inp[11]) ? node1254 : 4'b0010;
														assign node1254 = (inp[0]) ? 4'b0000 : 4'b0010;
											assign node1258 = (inp[13]) ? node1260 : 4'b0000;
												assign node1260 = (inp[15]) ? node1262 : 4'b0010;
													assign node1262 = (inp[1]) ? node1264 : 4'b0010;
														assign node1264 = (inp[11]) ? 4'b0000 : 4'b0010;
							assign node1267 = (inp[6]) ? node1283 : node1268;
								assign node1268 = (inp[13]) ? 4'b0110 : node1269;
									assign node1269 = (inp[9]) ? node1271 : 4'b0010;
										assign node1271 = (inp[8]) ? 4'b0000 : node1272;
											assign node1272 = (inp[15]) ? node1274 : 4'b0010;
												assign node1274 = (inp[11]) ? node1276 : 4'b0010;
													assign node1276 = (inp[7]) ? node1278 : 4'b0010;
														assign node1278 = (inp[1]) ? 4'b0000 : 4'b0010;
								assign node1283 = (inp[13]) ? 4'b0000 : node1284;
									assign node1284 = (inp[15]) ? node1286 : 4'b0000;
										assign node1286 = (inp[8]) ? node1288 : 4'b0000;
											assign node1288 = (inp[7]) ? node1290 : 4'b0000;
												assign node1290 = (inp[9]) ? 4'b0010 : 4'b0000;
					assign node1294 = (inp[14]) ? node1396 : node1295;
						assign node1295 = (inp[13]) ? node1345 : node1296;
							assign node1296 = (inp[2]) ? node1320 : node1297;
								assign node1297 = (inp[9]) ? node1307 : node1298;
									assign node1298 = (inp[6]) ? node1300 : 4'b0111;
										assign node1300 = (inp[7]) ? node1302 : 4'b0101;
											assign node1302 = (inp[8]) ? node1304 : 4'b0101;
												assign node1304 = (inp[15]) ? 4'b0111 : 4'b0101;
									assign node1307 = (inp[11]) ? node1309 : 4'b0111;
										assign node1309 = (inp[7]) ? node1311 : 4'b0111;
											assign node1311 = (inp[1]) ? node1313 : 4'b0111;
												assign node1313 = (inp[15]) ? node1315 : 4'b0111;
													assign node1315 = (inp[8]) ? node1317 : 4'b0111;
														assign node1317 = (inp[6]) ? 4'b0111 : 4'b0101;
								assign node1320 = (inp[6]) ? node1330 : node1321;
									assign node1321 = (inp[15]) ? node1323 : 4'b0101;
										assign node1323 = (inp[7]) ? node1325 : 4'b0101;
											assign node1325 = (inp[8]) ? node1327 : 4'b0101;
												assign node1327 = (inp[9]) ? 4'b0111 : 4'b0101;
									assign node1330 = (inp[9]) ? node1342 : node1331;
										assign node1331 = (inp[8]) ? 4'b0101 : node1332;
											assign node1332 = (inp[7]) ? 4'b0101 : node1333;
												assign node1333 = (inp[15]) ? node1335 : 4'b0111;
													assign node1335 = (inp[1]) ? node1337 : 4'b0111;
														assign node1337 = (inp[11]) ? 4'b0101 : 4'b0111;
										assign node1342 = (inp[8]) ? 4'b0011 : 4'b0101;
							assign node1345 = (inp[6]) ? node1365 : node1346;
								assign node1346 = (inp[2]) ? node1360 : node1347;
									assign node1347 = (inp[9]) ? node1349 : 4'b0111;
										assign node1349 = (inp[8]) ? node1351 : 4'b0111;
											assign node1351 = (inp[7]) ? 4'b0101 : node1352;
												assign node1352 = (inp[1]) ? node1354 : 4'b0111;
													assign node1354 = (inp[15]) ? node1356 : 4'b0111;
														assign node1356 = (inp[11]) ? 4'b0101 : 4'b0111;
									assign node1360 = (inp[8]) ? node1362 : 4'b0101;
										assign node1362 = (inp[9]) ? 4'b0011 : 4'b0101;
								assign node1365 = (inp[9]) ? node1387 : node1366;
									assign node1366 = (inp[8]) ? node1368 : 4'b0011;
										assign node1368 = (inp[7]) ? node1378 : node1369;
											assign node1369 = (inp[11]) ? node1371 : 4'b0011;
												assign node1371 = (inp[2]) ? 4'b0011 : node1372;
													assign node1372 = (inp[15]) ? node1374 : 4'b0011;
														assign node1374 = (inp[1]) ? 4'b0001 : 4'b0011;
											assign node1378 = (inp[2]) ? node1380 : 4'b0001;
												assign node1380 = (inp[1]) ? node1382 : 4'b0011;
													assign node1382 = (inp[11]) ? node1384 : 4'b0011;
														assign node1384 = (inp[15]) ? 4'b0001 : 4'b0011;
									assign node1387 = (inp[8]) ? node1389 : 4'b0001;
										assign node1389 = (inp[2]) ? 4'b0001 : node1390;
											assign node1390 = (inp[15]) ? node1392 : 4'b0001;
												assign node1392 = (inp[7]) ? 4'b0011 : 4'b0001;
						assign node1396 = (inp[6]) ? node1448 : node1397;
							assign node1397 = (inp[2]) ? node1425 : node1398;
								assign node1398 = (inp[9]) ? node1412 : node1399;
									assign node1399 = (inp[13]) ? node1401 : 4'b0011;
										assign node1401 = (inp[8]) ? 4'b0001 : node1402;
											assign node1402 = (inp[1]) ? node1404 : 4'b0011;
												assign node1404 = (inp[11]) ? node1406 : 4'b0011;
													assign node1406 = (inp[15]) ? node1408 : 4'b0011;
														assign node1408 = (inp[7]) ? 4'b0001 : 4'b0011;
									assign node1412 = (inp[13]) ? 4'b0001 : node1413;
										assign node1413 = (inp[7]) ? 4'b0001 : node1414;
											assign node1414 = (inp[8]) ? 4'b0001 : node1415;
												assign node1415 = (inp[11]) ? node1417 : 4'b0011;
													assign node1417 = (inp[15]) ? node1419 : 4'b0011;
														assign node1419 = (inp[1]) ? 4'b0001 : 4'b0011;
								assign node1425 = (inp[13]) ? node1435 : node1426;
									assign node1426 = (inp[9]) ? 4'b0011 : node1427;
										assign node1427 = (inp[15]) ? node1429 : 4'b0001;
											assign node1429 = (inp[8]) ? node1431 : 4'b0001;
												assign node1431 = (inp[7]) ? 4'b0011 : 4'b0001;
									assign node1435 = (inp[9]) ? node1437 : 4'b0111;
										assign node1437 = (inp[8]) ? 4'b0101 : node1438;
											assign node1438 = (inp[7]) ? node1440 : 4'b0111;
												assign node1440 = (inp[15]) ? node1442 : 4'b0111;
													assign node1442 = (inp[11]) ? node1444 : 4'b0111;
														assign node1444 = (inp[1]) ? 4'b0101 : 4'b0111;
							assign node1448 = (inp[13]) ? node1480 : node1449;
								assign node1449 = (inp[9]) ? node1471 : node1450;
									assign node1450 = (inp[8]) ? node1452 : 4'b0110;
										assign node1452 = (inp[2]) ? node1462 : node1453;
											assign node1453 = (inp[7]) ? node1455 : 4'b0110;
												assign node1455 = (inp[15]) ? node1457 : 4'b0110;
													assign node1457 = (inp[11]) ? node1459 : 4'b0110;
														assign node1459 = (inp[1]) ? 4'b0100 : 4'b0110;
											assign node1462 = (inp[7]) ? 4'b0100 : node1463;
												assign node1463 = (inp[11]) ? node1465 : 4'b0110;
													assign node1465 = (inp[15]) ? node1467 : 4'b0110;
														assign node1467 = (inp[1]) ? 4'b0100 : 4'b0110;
									assign node1471 = (inp[8]) ? node1473 : 4'b0100;
										assign node1473 = (inp[2]) ? 4'b0010 : node1474;
											assign node1474 = (inp[7]) ? node1476 : 4'b0100;
												assign node1476 = (inp[15]) ? 4'b0110 : 4'b0100;
								assign node1480 = (inp[2]) ? node1508 : node1481;
									assign node1481 = (inp[8]) ? node1501 : node1482;
										assign node1482 = (inp[7]) ? node1492 : node1483;
											assign node1483 = (inp[15]) ? node1485 : 4'b0010;
												assign node1485 = (inp[1]) ? node1487 : 4'b0010;
													assign node1487 = (inp[9]) ? 4'b0010 : node1488;
														assign node1488 = (inp[11]) ? 4'b0000 : 4'b0010;
											assign node1492 = (inp[9]) ? node1494 : 4'b0000;
												assign node1494 = (inp[11]) ? node1496 : 4'b0010;
													assign node1496 = (inp[1]) ? node1498 : 4'b0010;
														assign node1498 = (inp[15]) ? 4'b0000 : 4'b0010;
										assign node1501 = (inp[9]) ? 4'b0000 : node1502;
											assign node1502 = (inp[7]) ? node1504 : 4'b0000;
												assign node1504 = (inp[15]) ? 4'b0010 : 4'b0000;
									assign node1508 = (inp[8]) ? node1528 : node1509;
										assign node1509 = (inp[9]) ? node1519 : node1510;
											assign node1510 = (inp[1]) ? node1512 : 4'b0110;
												assign node1512 = (inp[11]) ? node1514 : 4'b0110;
													assign node1514 = (inp[15]) ? node1516 : 4'b0110;
														assign node1516 = (inp[7]) ? 4'b0100 : 4'b0110;
											assign node1519 = (inp[7]) ? 4'b0100 : node1520;
												assign node1520 = (inp[11]) ? node1522 : 4'b0110;
													assign node1522 = (inp[15]) ? node1524 : 4'b0110;
														assign node1524 = (inp[1]) ? 4'b0100 : 4'b0110;
										assign node1528 = (inp[9]) ? node1534 : node1529;
											assign node1529 = (inp[15]) ? node1531 : 4'b0100;
												assign node1531 = (inp[7]) ? 4'b0110 : 4'b0100;
											assign node1534 = (inp[7]) ? node1542 : node1535;
												assign node1535 = (inp[15]) ? node1537 : 4'b0010;
													assign node1537 = (inp[1]) ? node1539 : 4'b0010;
														assign node1539 = (inp[11]) ? 4'b0000 : 4'b0010;
												assign node1542 = (inp[15]) ? node1544 : 4'b0000;
													assign node1544 = (inp[11]) ? node1546 : 4'b0010;
														assign node1546 = (inp[1]) ? 4'b0000 : 4'b0010;

endmodule