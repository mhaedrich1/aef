module dtc_split125_bm21 (
	input  wire [10-1:0] inp,
	output wire [10-1:0] outp
);

	wire [10-1:0] node1;
	wire [10-1:0] node2;
	wire [10-1:0] node3;
	wire [10-1:0] node4;
	wire [10-1:0] node5;
	wire [10-1:0] node6;
	wire [10-1:0] node7;
	wire [10-1:0] node11;
	wire [10-1:0] node12;
	wire [10-1:0] node16;
	wire [10-1:0] node17;
	wire [10-1:0] node20;
	wire [10-1:0] node23;
	wire [10-1:0] node25;
	wire [10-1:0] node28;
	wire [10-1:0] node30;
	wire [10-1:0] node31;
	wire [10-1:0] node34;
	wire [10-1:0] node35;
	wire [10-1:0] node39;
	wire [10-1:0] node40;
	wire [10-1:0] node41;
	wire [10-1:0] node42;
	wire [10-1:0] node43;
	wire [10-1:0] node44;
	wire [10-1:0] node50;
	wire [10-1:0] node52;
	wire [10-1:0] node53;
	wire [10-1:0] node55;
	wire [10-1:0] node59;
	wire [10-1:0] node60;
	wire [10-1:0] node61;
	wire [10-1:0] node62;
	wire [10-1:0] node64;
	wire [10-1:0] node67;
	wire [10-1:0] node70;
	wire [10-1:0] node71;
	wire [10-1:0] node73;
	wire [10-1:0] node76;
	wire [10-1:0] node79;
	wire [10-1:0] node80;
	wire [10-1:0] node82;
	wire [10-1:0] node84;
	wire [10-1:0] node87;
	wire [10-1:0] node89;
	wire [10-1:0] node92;
	wire [10-1:0] node93;
	wire [10-1:0] node94;
	wire [10-1:0] node95;
	wire [10-1:0] node97;
	wire [10-1:0] node98;
	wire [10-1:0] node102;
	wire [10-1:0] node103;
	wire [10-1:0] node104;
	wire [10-1:0] node106;
	wire [10-1:0] node110;
	wire [10-1:0] node112;
	wire [10-1:0] node113;
	wire [10-1:0] node117;
	wire [10-1:0] node118;
	wire [10-1:0] node119;
	wire [10-1:0] node122;
	wire [10-1:0] node124;
	wire [10-1:0] node127;
	wire [10-1:0] node129;
	wire [10-1:0] node130;
	wire [10-1:0] node134;
	wire [10-1:0] node135;
	wire [10-1:0] node136;
	wire [10-1:0] node137;
	wire [10-1:0] node139;
	wire [10-1:0] node140;
	wire [10-1:0] node143;
	wire [10-1:0] node147;
	wire [10-1:0] node148;
	wire [10-1:0] node151;
	wire [10-1:0] node154;
	wire [10-1:0] node155;
	wire [10-1:0] node156;
	wire [10-1:0] node159;
	wire [10-1:0] node160;
	wire [10-1:0] node162;
	wire [10-1:0] node166;
	wire [10-1:0] node167;
	wire [10-1:0] node170;
	wire [10-1:0] node172;
	wire [10-1:0] node173;

	assign outp = (inp[6]) ? node92 : node1;
		assign node1 = (inp[5]) ? node39 : node2;
			assign node2 = (inp[8]) ? node28 : node3;
				assign node3 = (inp[3]) ? node23 : node4;
					assign node4 = (inp[7]) ? node16 : node5;
						assign node5 = (inp[1]) ? node11 : node6;
							assign node6 = (inp[9]) ? 10'b0011111111 : node7;
								assign node7 = (inp[0]) ? 10'b0011111111 : 10'b0111111111;
							assign node11 = (inp[2]) ? 10'b0001111111 : node12;
								assign node12 = (inp[0]) ? 10'b0001111111 : 10'b0011111111;
						assign node16 = (inp[1]) ? node20 : node17;
							assign node17 = (inp[9]) ? 10'b0001111111 : 10'b0011111111;
							assign node20 = (inp[0]) ? 10'b0000111111 : 10'b0001111111;
					assign node23 = (inp[0]) ? node25 : 10'b0001111111;
						assign node25 = (inp[7]) ? 10'b0000111111 : 10'b0000011111;
				assign node28 = (inp[7]) ? node30 : 10'b0000111111;
					assign node30 = (inp[4]) ? node34 : node31;
						assign node31 = (inp[2]) ? 10'b0000111111 : 10'b0001111111;
						assign node34 = (inp[3]) ? 10'b0000011111 : node35;
							assign node35 = (inp[2]) ? 10'b0000011111 : 10'b0000111111;
			assign node39 = (inp[3]) ? node59 : node40;
				assign node40 = (inp[8]) ? node50 : node41;
					assign node41 = (inp[4]) ? 10'b0000111111 : node42;
						assign node42 = (inp[7]) ? 10'b0000111111 : node43;
							assign node43 = (inp[2]) ? 10'b0001111111 : node44;
								assign node44 = (inp[0]) ? 10'b0001111111 : 10'b0011111111;
					assign node50 = (inp[1]) ? node52 : 10'b0000111111;
						assign node52 = (inp[2]) ? 10'b0000001111 : node53;
							assign node53 = (inp[7]) ? node55 : 10'b0000111111;
								assign node55 = (inp[0]) ? 10'b0000001111 : 10'b0000011111;
				assign node59 = (inp[7]) ? node79 : node60;
					assign node60 = (inp[9]) ? node70 : node61;
						assign node61 = (inp[8]) ? node67 : node62;
							assign node62 = (inp[2]) ? node64 : 10'b0000111111;
								assign node64 = (inp[0]) ? 10'b0000011111 : 10'b0000111111;
							assign node67 = (inp[1]) ? 10'b0000001111 : 10'b0000011111;
						assign node70 = (inp[0]) ? node76 : node71;
							assign node71 = (inp[4]) ? node73 : 10'b0000011111;
								assign node73 = (inp[2]) ? 10'b0000001111 : 10'b0000011111;
							assign node76 = (inp[8]) ? 10'b0000000111 : 10'b0000001111;
					assign node79 = (inp[2]) ? node87 : node80;
						assign node80 = (inp[8]) ? node82 : 10'b0000111111;
							assign node82 = (inp[1]) ? node84 : 10'b0000001111;
								assign node84 = (inp[4]) ? 10'b0000000111 : 10'b0000001111;
						assign node87 = (inp[9]) ? node89 : 10'b0000000111;
							assign node89 = (inp[8]) ? 10'b0000000001 : 10'b0000000011;
		assign node92 = (inp[9]) ? node134 : node93;
			assign node93 = (inp[3]) ? node117 : node94;
				assign node94 = (inp[5]) ? node102 : node95;
					assign node95 = (inp[7]) ? node97 : 10'b0000111111;
						assign node97 = (inp[0]) ? 10'b0000001111 : node98;
							assign node98 = (inp[4]) ? 10'b0000011111 : 10'b0000111111;
					assign node102 = (inp[4]) ? node110 : node103;
						assign node103 = (inp[8]) ? 10'b0000011111 : node104;
							assign node104 = (inp[0]) ? node106 : 10'b0000111111;
								assign node106 = (inp[2]) ? 10'b0000011111 : 10'b0000111111;
						assign node110 = (inp[2]) ? node112 : 10'b0000011111;
							assign node112 = (inp[1]) ? 10'b0000001111 : node113;
								assign node113 = (inp[8]) ? 10'b0000001111 : 10'b0000011111;
				assign node117 = (inp[1]) ? node127 : node118;
					assign node118 = (inp[7]) ? node122 : node119;
						assign node119 = (inp[2]) ? 10'b0000011111 : 10'b0001111111;
						assign node122 = (inp[4]) ? node124 : 10'b0000011111;
							assign node124 = (inp[8]) ? 10'b0000011111 : 10'b0000001111;
					assign node127 = (inp[4]) ? node129 : 10'b0000011111;
						assign node129 = (inp[5]) ? 10'b0000000111 : node130;
							assign node130 = (inp[8]) ? 10'b0000011111 : 10'b0000001111;
			assign node134 = (inp[0]) ? node154 : node135;
				assign node135 = (inp[5]) ? node147 : node136;
					assign node136 = (inp[1]) ? 10'b0000011111 : node137;
						assign node137 = (inp[4]) ? node139 : 10'b0000111111;
							assign node139 = (inp[3]) ? node143 : node140;
								assign node140 = (inp[8]) ? 10'b0000011111 : 10'b0000111111;
								assign node143 = (inp[8]) ? 10'b0000001111 : 10'b0000011111;
					assign node147 = (inp[2]) ? node151 : node148;
						assign node148 = (inp[7]) ? 10'b0000001111 : 10'b0000011111;
						assign node151 = (inp[1]) ? 10'b0000000001 : 10'b0000000111;
				assign node154 = (inp[5]) ? node166 : node155;
					assign node155 = (inp[2]) ? node159 : node156;
						assign node156 = (inp[7]) ? 10'b0000001111 : 10'b0000011111;
						assign node159 = (inp[3]) ? 10'b0000000011 : node160;
							assign node160 = (inp[4]) ? node162 : 10'b0000001111;
								assign node162 = (inp[7]) ? 10'b0000000111 : 10'b0000001111;
					assign node166 = (inp[4]) ? node170 : node167;
						assign node167 = (inp[1]) ? 10'b0000000111 : 10'b0000011111;
						assign node170 = (inp[1]) ? node172 : 10'b0000000111;
							assign node172 = (inp[8]) ? 10'b0000000001 : node173;
								assign node173 = (inp[7]) ? 10'b0000000011 : 10'b0000000111;

endmodule