module dtc_split33_bm57 (
	input  wire [12-1:0] inp,
	output wire [3-1:0] outp
);

	wire [3-1:0] node1;
	wire [3-1:0] node2;
	wire [3-1:0] node3;
	wire [3-1:0] node4;
	wire [3-1:0] node5;
	wire [3-1:0] node6;
	wire [3-1:0] node7;
	wire [3-1:0] node8;
	wire [3-1:0] node9;
	wire [3-1:0] node12;
	wire [3-1:0] node13;
	wire [3-1:0] node16;
	wire [3-1:0] node18;
	wire [3-1:0] node21;
	wire [3-1:0] node23;
	wire [3-1:0] node26;
	wire [3-1:0] node27;
	wire [3-1:0] node30;
	wire [3-1:0] node32;
	wire [3-1:0] node33;
	wire [3-1:0] node36;
	wire [3-1:0] node39;
	wire [3-1:0] node40;
	wire [3-1:0] node41;
	wire [3-1:0] node42;
	wire [3-1:0] node45;
	wire [3-1:0] node48;
	wire [3-1:0] node49;
	wire [3-1:0] node52;
	wire [3-1:0] node54;
	wire [3-1:0] node57;
	wire [3-1:0] node58;
	wire [3-1:0] node59;
	wire [3-1:0] node63;
	wire [3-1:0] node64;
	wire [3-1:0] node67;
	wire [3-1:0] node69;
	wire [3-1:0] node72;
	wire [3-1:0] node73;
	wire [3-1:0] node74;
	wire [3-1:0] node76;
	wire [3-1:0] node77;
	wire [3-1:0] node80;
	wire [3-1:0] node83;
	wire [3-1:0] node84;
	wire [3-1:0] node85;
	wire [3-1:0] node88;
	wire [3-1:0] node89;
	wire [3-1:0] node92;
	wire [3-1:0] node95;
	wire [3-1:0] node96;
	wire [3-1:0] node97;
	wire [3-1:0] node100;
	wire [3-1:0] node104;
	wire [3-1:0] node105;
	wire [3-1:0] node106;
	wire [3-1:0] node108;
	wire [3-1:0] node109;
	wire [3-1:0] node112;
	wire [3-1:0] node115;
	wire [3-1:0] node116;
	wire [3-1:0] node119;
	wire [3-1:0] node120;
	wire [3-1:0] node124;
	wire [3-1:0] node125;
	wire [3-1:0] node126;
	wire [3-1:0] node129;
	wire [3-1:0] node130;
	wire [3-1:0] node132;
	wire [3-1:0] node136;
	wire [3-1:0] node137;
	wire [3-1:0] node141;
	wire [3-1:0] node142;
	wire [3-1:0] node143;
	wire [3-1:0] node144;
	wire [3-1:0] node146;
	wire [3-1:0] node148;
	wire [3-1:0] node151;
	wire [3-1:0] node153;
	wire [3-1:0] node155;
	wire [3-1:0] node158;
	wire [3-1:0] node159;
	wire [3-1:0] node160;
	wire [3-1:0] node161;
	wire [3-1:0] node162;
	wire [3-1:0] node166;
	wire [3-1:0] node168;
	wire [3-1:0] node169;
	wire [3-1:0] node172;
	wire [3-1:0] node176;
	wire [3-1:0] node178;
	wire [3-1:0] node179;
	wire [3-1:0] node182;
	wire [3-1:0] node185;
	wire [3-1:0] node186;
	wire [3-1:0] node187;
	wire [3-1:0] node188;
	wire [3-1:0] node190;
	wire [3-1:0] node192;
	wire [3-1:0] node195;
	wire [3-1:0] node197;
	wire [3-1:0] node198;
	wire [3-1:0] node202;
	wire [3-1:0] node203;
	wire [3-1:0] node205;
	wire [3-1:0] node207;
	wire [3-1:0] node210;
	wire [3-1:0] node211;
	wire [3-1:0] node215;
	wire [3-1:0] node216;
	wire [3-1:0] node219;
	wire [3-1:0] node220;
	wire [3-1:0] node223;
	wire [3-1:0] node224;
	wire [3-1:0] node228;
	wire [3-1:0] node229;
	wire [3-1:0] node230;
	wire [3-1:0] node231;
	wire [3-1:0] node232;
	wire [3-1:0] node233;
	wire [3-1:0] node237;
	wire [3-1:0] node238;
	wire [3-1:0] node239;
	wire [3-1:0] node240;
	wire [3-1:0] node244;
	wire [3-1:0] node248;
	wire [3-1:0] node249;
	wire [3-1:0] node250;
	wire [3-1:0] node251;
	wire [3-1:0] node252;
	wire [3-1:0] node257;
	wire [3-1:0] node259;
	wire [3-1:0] node262;
	wire [3-1:0] node263;
	wire [3-1:0] node264;
	wire [3-1:0] node265;
	wire [3-1:0] node269;
	wire [3-1:0] node270;
	wire [3-1:0] node272;
	wire [3-1:0] node276;
	wire [3-1:0] node278;
	wire [3-1:0] node281;
	wire [3-1:0] node282;
	wire [3-1:0] node283;
	wire [3-1:0] node284;
	wire [3-1:0] node285;
	wire [3-1:0] node288;
	wire [3-1:0] node291;
	wire [3-1:0] node292;
	wire [3-1:0] node295;
	wire [3-1:0] node298;
	wire [3-1:0] node299;
	wire [3-1:0] node300;
	wire [3-1:0] node303;
	wire [3-1:0] node304;
	wire [3-1:0] node309;
	wire [3-1:0] node310;
	wire [3-1:0] node311;
	wire [3-1:0] node313;
	wire [3-1:0] node314;
	wire [3-1:0] node315;
	wire [3-1:0] node320;
	wire [3-1:0] node323;
	wire [3-1:0] node324;
	wire [3-1:0] node326;
	wire [3-1:0] node329;
	wire [3-1:0] node330;
	wire [3-1:0] node334;
	wire [3-1:0] node335;
	wire [3-1:0] node336;
	wire [3-1:0] node337;
	wire [3-1:0] node338;
	wire [3-1:0] node339;
	wire [3-1:0] node342;
	wire [3-1:0] node343;
	wire [3-1:0] node344;
	wire [3-1:0] node348;
	wire [3-1:0] node351;
	wire [3-1:0] node352;
	wire [3-1:0] node353;
	wire [3-1:0] node355;
	wire [3-1:0] node359;
	wire [3-1:0] node362;
	wire [3-1:0] node363;
	wire [3-1:0] node365;
	wire [3-1:0] node366;
	wire [3-1:0] node368;
	wire [3-1:0] node372;
	wire [3-1:0] node374;
	wire [3-1:0] node377;
	wire [3-1:0] node378;
	wire [3-1:0] node379;
	wire [3-1:0] node381;
	wire [3-1:0] node384;
	wire [3-1:0] node385;
	wire [3-1:0] node389;
	wire [3-1:0] node390;
	wire [3-1:0] node391;
	wire [3-1:0] node393;
	wire [3-1:0] node396;
	wire [3-1:0] node399;
	wire [3-1:0] node401;
	wire [3-1:0] node402;
	wire [3-1:0] node406;
	wire [3-1:0] node407;
	wire [3-1:0] node408;
	wire [3-1:0] node409;
	wire [3-1:0] node410;
	wire [3-1:0] node414;
	wire [3-1:0] node415;
	wire [3-1:0] node417;
	wire [3-1:0] node420;
	wire [3-1:0] node422;
	wire [3-1:0] node425;
	wire [3-1:0] node426;
	wire [3-1:0] node427;
	wire [3-1:0] node431;
	wire [3-1:0] node434;
	wire [3-1:0] node435;
	wire [3-1:0] node436;
	wire [3-1:0] node437;
	wire [3-1:0] node439;
	wire [3-1:0] node443;
	wire [3-1:0] node446;
	wire [3-1:0] node447;
	wire [3-1:0] node448;
	wire [3-1:0] node450;
	wire [3-1:0] node452;
	wire [3-1:0] node457;
	wire [3-1:0] node458;
	wire [3-1:0] node459;
	wire [3-1:0] node460;
	wire [3-1:0] node461;
	wire [3-1:0] node462;
	wire [3-1:0] node463;
	wire [3-1:0] node467;
	wire [3-1:0] node468;
	wire [3-1:0] node469;
	wire [3-1:0] node470;
	wire [3-1:0] node475;
	wire [3-1:0] node476;
	wire [3-1:0] node477;
	wire [3-1:0] node480;
	wire [3-1:0] node483;
	wire [3-1:0] node484;
	wire [3-1:0] node488;
	wire [3-1:0] node489;
	wire [3-1:0] node490;
	wire [3-1:0] node491;
	wire [3-1:0] node493;
	wire [3-1:0] node497;
	wire [3-1:0] node499;
	wire [3-1:0] node500;
	wire [3-1:0] node503;
	wire [3-1:0] node506;
	wire [3-1:0] node507;
	wire [3-1:0] node508;
	wire [3-1:0] node509;
	wire [3-1:0] node514;
	wire [3-1:0] node515;
	wire [3-1:0] node517;
	wire [3-1:0] node521;
	wire [3-1:0] node522;
	wire [3-1:0] node523;
	wire [3-1:0] node525;
	wire [3-1:0] node526;
	wire [3-1:0] node528;
	wire [3-1:0] node529;
	wire [3-1:0] node533;
	wire [3-1:0] node535;
	wire [3-1:0] node538;
	wire [3-1:0] node540;
	wire [3-1:0] node541;
	wire [3-1:0] node543;
	wire [3-1:0] node547;
	wire [3-1:0] node548;
	wire [3-1:0] node549;
	wire [3-1:0] node550;
	wire [3-1:0] node552;
	wire [3-1:0] node553;
	wire [3-1:0] node559;
	wire [3-1:0] node560;
	wire [3-1:0] node561;
	wire [3-1:0] node565;
	wire [3-1:0] node567;
	wire [3-1:0] node570;
	wire [3-1:0] node571;
	wire [3-1:0] node572;
	wire [3-1:0] node573;
	wire [3-1:0] node574;
	wire [3-1:0] node577;
	wire [3-1:0] node578;
	wire [3-1:0] node581;
	wire [3-1:0] node584;
	wire [3-1:0] node585;
	wire [3-1:0] node588;
	wire [3-1:0] node589;
	wire [3-1:0] node592;
	wire [3-1:0] node595;
	wire [3-1:0] node596;
	wire [3-1:0] node597;
	wire [3-1:0] node599;
	wire [3-1:0] node602;
	wire [3-1:0] node605;
	wire [3-1:0] node606;
	wire [3-1:0] node608;
	wire [3-1:0] node611;
	wire [3-1:0] node614;
	wire [3-1:0] node615;
	wire [3-1:0] node616;
	wire [3-1:0] node617;
	wire [3-1:0] node619;
	wire [3-1:0] node622;
	wire [3-1:0] node623;
	wire [3-1:0] node624;
	wire [3-1:0] node628;
	wire [3-1:0] node631;
	wire [3-1:0] node633;
	wire [3-1:0] node634;
	wire [3-1:0] node637;
	wire [3-1:0] node640;
	wire [3-1:0] node641;
	wire [3-1:0] node642;
	wire [3-1:0] node645;
	wire [3-1:0] node646;
	wire [3-1:0] node649;
	wire [3-1:0] node652;
	wire [3-1:0] node653;
	wire [3-1:0] node654;
	wire [3-1:0] node657;
	wire [3-1:0] node660;
	wire [3-1:0] node662;
	wire [3-1:0] node664;
	wire [3-1:0] node667;
	wire [3-1:0] node668;
	wire [3-1:0] node669;
	wire [3-1:0] node670;
	wire [3-1:0] node671;
	wire [3-1:0] node672;
	wire [3-1:0] node673;
	wire [3-1:0] node675;
	wire [3-1:0] node678;
	wire [3-1:0] node679;
	wire [3-1:0] node683;
	wire [3-1:0] node684;
	wire [3-1:0] node685;
	wire [3-1:0] node689;
	wire [3-1:0] node692;
	wire [3-1:0] node693;
	wire [3-1:0] node695;
	wire [3-1:0] node697;
	wire [3-1:0] node698;
	wire [3-1:0] node701;
	wire [3-1:0] node704;
	wire [3-1:0] node707;
	wire [3-1:0] node708;
	wire [3-1:0] node709;
	wire [3-1:0] node710;
	wire [3-1:0] node712;
	wire [3-1:0] node715;
	wire [3-1:0] node717;
	wire [3-1:0] node721;
	wire [3-1:0] node723;
	wire [3-1:0] node724;
	wire [3-1:0] node725;
	wire [3-1:0] node726;
	wire [3-1:0] node732;
	wire [3-1:0] node733;
	wire [3-1:0] node734;
	wire [3-1:0] node735;
	wire [3-1:0] node736;
	wire [3-1:0] node741;
	wire [3-1:0] node742;
	wire [3-1:0] node746;
	wire [3-1:0] node747;
	wire [3-1:0] node748;
	wire [3-1:0] node752;
	wire [3-1:0] node753;
	wire [3-1:0] node757;
	wire [3-1:0] node758;
	wire [3-1:0] node759;
	wire [3-1:0] node760;
	wire [3-1:0] node761;
	wire [3-1:0] node764;
	wire [3-1:0] node765;
	wire [3-1:0] node766;
	wire [3-1:0] node767;
	wire [3-1:0] node773;
	wire [3-1:0] node774;
	wire [3-1:0] node777;
	wire [3-1:0] node780;
	wire [3-1:0] node781;
	wire [3-1:0] node782;
	wire [3-1:0] node784;
	wire [3-1:0] node785;
	wire [3-1:0] node788;
	wire [3-1:0] node791;
	wire [3-1:0] node794;
	wire [3-1:0] node795;
	wire [3-1:0] node797;
	wire [3-1:0] node799;
	wire [3-1:0] node802;
	wire [3-1:0] node803;
	wire [3-1:0] node807;
	wire [3-1:0] node808;
	wire [3-1:0] node809;
	wire [3-1:0] node810;
	wire [3-1:0] node812;
	wire [3-1:0] node815;
	wire [3-1:0] node816;
	wire [3-1:0] node819;
	wire [3-1:0] node823;
	wire [3-1:0] node824;
	wire [3-1:0] node826;
	wire [3-1:0] node827;
	wire [3-1:0] node830;
	wire [3-1:0] node834;
	wire [3-1:0] node835;
	wire [3-1:0] node836;
	wire [3-1:0] node837;
	wire [3-1:0] node838;
	wire [3-1:0] node839;
	wire [3-1:0] node840;
	wire [3-1:0] node842;
	wire [3-1:0] node843;
	wire [3-1:0] node844;
	wire [3-1:0] node847;
	wire [3-1:0] node851;
	wire [3-1:0] node852;
	wire [3-1:0] node853;
	wire [3-1:0] node858;
	wire [3-1:0] node859;
	wire [3-1:0] node861;
	wire [3-1:0] node862;
	wire [3-1:0] node865;
	wire [3-1:0] node866;
	wire [3-1:0] node870;
	wire [3-1:0] node871;
	wire [3-1:0] node874;
	wire [3-1:0] node876;
	wire [3-1:0] node879;
	wire [3-1:0] node880;
	wire [3-1:0] node881;
	wire [3-1:0] node882;
	wire [3-1:0] node883;
	wire [3-1:0] node886;
	wire [3-1:0] node890;
	wire [3-1:0] node891;
	wire [3-1:0] node893;
	wire [3-1:0] node894;
	wire [3-1:0] node896;
	wire [3-1:0] node900;
	wire [3-1:0] node902;
	wire [3-1:0] node905;
	wire [3-1:0] node906;
	wire [3-1:0] node907;
	wire [3-1:0] node911;
	wire [3-1:0] node912;
	wire [3-1:0] node914;
	wire [3-1:0] node915;
	wire [3-1:0] node920;
	wire [3-1:0] node921;
	wire [3-1:0] node922;
	wire [3-1:0] node923;
	wire [3-1:0] node924;
	wire [3-1:0] node925;
	wire [3-1:0] node927;
	wire [3-1:0] node930;
	wire [3-1:0] node931;
	wire [3-1:0] node934;
	wire [3-1:0] node936;
	wire [3-1:0] node940;
	wire [3-1:0] node941;
	wire [3-1:0] node942;
	wire [3-1:0] node947;
	wire [3-1:0] node948;
	wire [3-1:0] node949;
	wire [3-1:0] node951;
	wire [3-1:0] node954;
	wire [3-1:0] node955;
	wire [3-1:0] node960;
	wire [3-1:0] node961;
	wire [3-1:0] node962;
	wire [3-1:0] node963;
	wire [3-1:0] node967;
	wire [3-1:0] node968;
	wire [3-1:0] node969;
	wire [3-1:0] node971;
	wire [3-1:0] node976;
	wire [3-1:0] node977;
	wire [3-1:0] node978;
	wire [3-1:0] node979;
	wire [3-1:0] node980;
	wire [3-1:0] node986;
	wire [3-1:0] node987;
	wire [3-1:0] node988;
	wire [3-1:0] node991;
	wire [3-1:0] node994;
	wire [3-1:0] node995;
	wire [3-1:0] node999;
	wire [3-1:0] node1000;
	wire [3-1:0] node1001;
	wire [3-1:0] node1002;
	wire [3-1:0] node1003;
	wire [3-1:0] node1005;
	wire [3-1:0] node1006;
	wire [3-1:0] node1009;
	wire [3-1:0] node1012;
	wire [3-1:0] node1013;
	wire [3-1:0] node1014;
	wire [3-1:0] node1017;
	wire [3-1:0] node1021;
	wire [3-1:0] node1022;
	wire [3-1:0] node1023;
	wire [3-1:0] node1025;
	wire [3-1:0] node1026;
	wire [3-1:0] node1029;
	wire [3-1:0] node1032;
	wire [3-1:0] node1034;
	wire [3-1:0] node1037;
	wire [3-1:0] node1038;
	wire [3-1:0] node1039;
	wire [3-1:0] node1040;
	wire [3-1:0] node1046;
	wire [3-1:0] node1047;
	wire [3-1:0] node1048;
	wire [3-1:0] node1050;
	wire [3-1:0] node1051;
	wire [3-1:0] node1052;
	wire [3-1:0] node1054;
	wire [3-1:0] node1057;
	wire [3-1:0] node1060;
	wire [3-1:0] node1063;
	wire [3-1:0] node1064;
	wire [3-1:0] node1065;
	wire [3-1:0] node1066;
	wire [3-1:0] node1072;
	wire [3-1:0] node1073;
	wire [3-1:0] node1074;
	wire [3-1:0] node1076;
	wire [3-1:0] node1079;
	wire [3-1:0] node1080;
	wire [3-1:0] node1081;
	wire [3-1:0] node1086;
	wire [3-1:0] node1087;
	wire [3-1:0] node1089;
	wire [3-1:0] node1092;
	wire [3-1:0] node1093;
	wire [3-1:0] node1094;
	wire [3-1:0] node1097;
	wire [3-1:0] node1101;
	wire [3-1:0] node1102;
	wire [3-1:0] node1103;
	wire [3-1:0] node1104;
	wire [3-1:0] node1105;
	wire [3-1:0] node1109;
	wire [3-1:0] node1110;
	wire [3-1:0] node1112;
	wire [3-1:0] node1116;
	wire [3-1:0] node1117;
	wire [3-1:0] node1119;
	wire [3-1:0] node1122;
	wire [3-1:0] node1123;
	wire [3-1:0] node1125;
	wire [3-1:0] node1128;
	wire [3-1:0] node1129;
	wire [3-1:0] node1133;
	wire [3-1:0] node1134;
	wire [3-1:0] node1135;
	wire [3-1:0] node1139;
	wire [3-1:0] node1140;
	wire [3-1:0] node1144;
	wire [3-1:0] node1145;
	wire [3-1:0] node1146;
	wire [3-1:0] node1147;
	wire [3-1:0] node1148;
	wire [3-1:0] node1149;
	wire [3-1:0] node1150;
	wire [3-1:0] node1153;
	wire [3-1:0] node1156;
	wire [3-1:0] node1157;
	wire [3-1:0] node1159;
	wire [3-1:0] node1162;
	wire [3-1:0] node1163;
	wire [3-1:0] node1166;
	wire [3-1:0] node1169;
	wire [3-1:0] node1170;
	wire [3-1:0] node1173;
	wire [3-1:0] node1176;
	wire [3-1:0] node1177;
	wire [3-1:0] node1178;
	wire [3-1:0] node1180;
	wire [3-1:0] node1181;
	wire [3-1:0] node1185;
	wire [3-1:0] node1186;
	wire [3-1:0] node1187;
	wire [3-1:0] node1192;
	wire [3-1:0] node1193;
	wire [3-1:0] node1194;
	wire [3-1:0] node1198;
	wire [3-1:0] node1199;
	wire [3-1:0] node1203;
	wire [3-1:0] node1204;
	wire [3-1:0] node1205;
	wire [3-1:0] node1206;
	wire [3-1:0] node1209;
	wire [3-1:0] node1212;
	wire [3-1:0] node1213;
	wire [3-1:0] node1214;
	wire [3-1:0] node1217;
	wire [3-1:0] node1219;
	wire [3-1:0] node1220;
	wire [3-1:0] node1223;
	wire [3-1:0] node1226;
	wire [3-1:0] node1227;
	wire [3-1:0] node1228;
	wire [3-1:0] node1232;
	wire [3-1:0] node1234;
	wire [3-1:0] node1236;
	wire [3-1:0] node1239;
	wire [3-1:0] node1240;
	wire [3-1:0] node1241;
	wire [3-1:0] node1245;
	wire [3-1:0] node1246;
	wire [3-1:0] node1250;
	wire [3-1:0] node1251;
	wire [3-1:0] node1252;
	wire [3-1:0] node1253;
	wire [3-1:0] node1254;
	wire [3-1:0] node1255;
	wire [3-1:0] node1257;
	wire [3-1:0] node1260;
	wire [3-1:0] node1263;
	wire [3-1:0] node1264;
	wire [3-1:0] node1266;
	wire [3-1:0] node1268;
	wire [3-1:0] node1269;
	wire [3-1:0] node1273;
	wire [3-1:0] node1276;
	wire [3-1:0] node1277;
	wire [3-1:0] node1279;
	wire [3-1:0] node1282;
	wire [3-1:0] node1283;
	wire [3-1:0] node1284;
	wire [3-1:0] node1287;
	wire [3-1:0] node1290;
	wire [3-1:0] node1291;
	wire [3-1:0] node1295;
	wire [3-1:0] node1296;
	wire [3-1:0] node1297;
	wire [3-1:0] node1298;
	wire [3-1:0] node1299;
	wire [3-1:0] node1305;
	wire [3-1:0] node1306;
	wire [3-1:0] node1310;
	wire [3-1:0] node1311;
	wire [3-1:0] node1312;
	wire [3-1:0] node1313;
	wire [3-1:0] node1314;
	wire [3-1:0] node1316;
	wire [3-1:0] node1317;
	wire [3-1:0] node1320;
	wire [3-1:0] node1323;
	wire [3-1:0] node1324;
	wire [3-1:0] node1325;
	wire [3-1:0] node1328;
	wire [3-1:0] node1332;
	wire [3-1:0] node1335;
	wire [3-1:0] node1336;
	wire [3-1:0] node1337;
	wire [3-1:0] node1338;
	wire [3-1:0] node1341;
	wire [3-1:0] node1344;
	wire [3-1:0] node1347;
	wire [3-1:0] node1348;
	wire [3-1:0] node1349;
	wire [3-1:0] node1352;
	wire [3-1:0] node1353;
	wire [3-1:0] node1358;
	wire [3-1:0] node1359;

	assign outp = (inp[4]) ? node834 : node1;
		assign node1 = (inp[6]) ? node457 : node2;
			assign node2 = (inp[5]) ? node228 : node3;
				assign node3 = (inp[8]) ? node141 : node4;
					assign node4 = (inp[1]) ? node72 : node5;
						assign node5 = (inp[9]) ? node39 : node6;
							assign node6 = (inp[7]) ? node26 : node7;
								assign node7 = (inp[0]) ? node21 : node8;
									assign node8 = (inp[10]) ? node12 : node9;
										assign node9 = (inp[3]) ? 3'b010 : 3'b000;
										assign node12 = (inp[3]) ? node16 : node13;
											assign node13 = (inp[11]) ? 3'b011 : 3'b010;
											assign node16 = (inp[11]) ? node18 : 3'b001;
												assign node18 = (inp[2]) ? 3'b000 : 3'b001;
									assign node21 = (inp[11]) ? node23 : 3'b011;
										assign node23 = (inp[10]) ? 3'b010 : 3'b011;
								assign node26 = (inp[0]) ? node30 : node27;
									assign node27 = (inp[3]) ? 3'b011 : 3'b010;
									assign node30 = (inp[10]) ? node32 : 3'b001;
										assign node32 = (inp[11]) ? node36 : node33;
											assign node33 = (inp[3]) ? 3'b001 : 3'b011;
											assign node36 = (inp[3]) ? 3'b010 : 3'b001;
							assign node39 = (inp[11]) ? node57 : node40;
								assign node40 = (inp[0]) ? node48 : node41;
									assign node41 = (inp[3]) ? node45 : node42;
										assign node42 = (inp[10]) ? 3'b011 : 3'b001;
										assign node45 = (inp[10]) ? 3'b000 : 3'b010;
									assign node48 = (inp[3]) ? node52 : node49;
										assign node49 = (inp[10]) ? 3'b010 : 3'b000;
										assign node52 = (inp[2]) ? node54 : 3'b000;
											assign node54 = (inp[7]) ? 3'b000 : 3'b001;
								assign node57 = (inp[3]) ? node63 : node58;
									assign node58 = (inp[2]) ? 3'b010 : node59;
										assign node59 = (inp[10]) ? 3'b010 : 3'b011;
									assign node63 = (inp[10]) ? node67 : node64;
										assign node64 = (inp[7]) ? 3'b000 : 3'b010;
										assign node67 = (inp[7]) ? node69 : 3'b001;
											assign node69 = (inp[0]) ? 3'b011 : 3'b010;
						assign node72 = (inp[7]) ? node104 : node73;
							assign node73 = (inp[0]) ? node83 : node74;
								assign node74 = (inp[2]) ? node76 : 3'b000;
									assign node76 = (inp[10]) ? node80 : node77;
										assign node77 = (inp[11]) ? 3'b010 : 3'b011;
										assign node80 = (inp[3]) ? 3'b001 : 3'b011;
								assign node83 = (inp[11]) ? node95 : node84;
									assign node84 = (inp[3]) ? node88 : node85;
										assign node85 = (inp[2]) ? 3'b001 : 3'b010;
										assign node88 = (inp[9]) ? node92 : node89;
											assign node89 = (inp[2]) ? 3'b010 : 3'b011;
											assign node92 = (inp[2]) ? 3'b011 : 3'b010;
									assign node95 = (inp[9]) ? 3'b011 : node96;
										assign node96 = (inp[10]) ? node100 : node97;
											assign node97 = (inp[2]) ? 3'b010 : 3'b011;
											assign node100 = (inp[2]) ? 3'b011 : 3'b010;
							assign node104 = (inp[11]) ? node124 : node105;
								assign node105 = (inp[0]) ? node115 : node106;
									assign node106 = (inp[9]) ? node108 : 3'b000;
										assign node108 = (inp[2]) ? node112 : node109;
											assign node109 = (inp[10]) ? 3'b011 : 3'b010;
											assign node112 = (inp[10]) ? 3'b010 : 3'b011;
									assign node115 = (inp[9]) ? node119 : node116;
										assign node116 = (inp[3]) ? 3'b001 : 3'b011;
										assign node119 = (inp[3]) ? 3'b000 : node120;
											assign node120 = (inp[2]) ? 3'b001 : 3'b000;
								assign node124 = (inp[0]) ? node136 : node125;
									assign node125 = (inp[10]) ? node129 : node126;
										assign node126 = (inp[3]) ? 3'b001 : 3'b011;
										assign node129 = (inp[3]) ? 3'b011 : node130;
											assign node130 = (inp[9]) ? node132 : 3'b001;
												assign node132 = (inp[2]) ? 3'b000 : 3'b001;
									assign node136 = (inp[2]) ? 3'b011 : node137;
										assign node137 = (inp[10]) ? 3'b010 : 3'b011;
					assign node141 = (inp[1]) ? node185 : node142;
						assign node142 = (inp[9]) ? node158 : node143;
							assign node143 = (inp[3]) ? node151 : node144;
								assign node144 = (inp[7]) ? node146 : 3'b100;
									assign node146 = (inp[0]) ? node148 : 3'b110;
										assign node148 = (inp[10]) ? 3'b111 : 3'b110;
								assign node151 = (inp[7]) ? node153 : 3'b110;
									assign node153 = (inp[0]) ? node155 : 3'b100;
										assign node155 = (inp[10]) ? 3'b100 : 3'b101;
							assign node158 = (inp[10]) ? node176 : node159;
								assign node159 = (inp[11]) ? 3'b101 : node160;
									assign node160 = (inp[2]) ? node166 : node161;
										assign node161 = (inp[3]) ? 3'b100 : node162;
											assign node162 = (inp[7]) ? 3'b111 : 3'b101;
										assign node166 = (inp[0]) ? node168 : 3'b111;
											assign node168 = (inp[3]) ? node172 : node169;
												assign node169 = (inp[7]) ? 3'b111 : 3'b101;
												assign node172 = (inp[7]) ? 3'b101 : 3'b111;
								assign node176 = (inp[2]) ? node178 : 3'b100;
									assign node178 = (inp[3]) ? node182 : node179;
										assign node179 = (inp[7]) ? 3'b110 : 3'b100;
										assign node182 = (inp[11]) ? 3'b111 : 3'b101;
						assign node185 = (inp[9]) ? node215 : node186;
							assign node186 = (inp[7]) ? node202 : node187;
								assign node187 = (inp[3]) ? node195 : node188;
									assign node188 = (inp[10]) ? node190 : 3'b101;
										assign node190 = (inp[0]) ? node192 : 3'b101;
											assign node192 = (inp[11]) ? 3'b100 : 3'b101;
									assign node195 = (inp[11]) ? node197 : 3'b111;
										assign node197 = (inp[2]) ? 3'b111 : node198;
											assign node198 = (inp[10]) ? 3'b110 : 3'b111;
								assign node202 = (inp[3]) ? node210 : node203;
									assign node203 = (inp[2]) ? node205 : 3'b111;
										assign node205 = (inp[11]) ? node207 : 3'b110;
											assign node207 = (inp[10]) ? 3'b111 : 3'b110;
									assign node210 = (inp[2]) ? 3'b101 : node211;
										assign node211 = (inp[11]) ? 3'b101 : 3'b100;
							assign node215 = (inp[7]) ? node219 : node216;
								assign node216 = (inp[3]) ? 3'b110 : 3'b100;
								assign node219 = (inp[3]) ? node223 : node220;
									assign node220 = (inp[2]) ? 3'b111 : 3'b110;
									assign node223 = (inp[2]) ? 3'b100 : node224;
										assign node224 = (inp[10]) ? 3'b101 : 3'b100;
				assign node228 = (inp[0]) ? node334 : node229;
					assign node229 = (inp[3]) ? node281 : node230;
						assign node230 = (inp[7]) ? node248 : node231;
							assign node231 = (inp[9]) ? node237 : node232;
								assign node232 = (inp[8]) ? 3'b100 : node233;
									assign node233 = (inp[2]) ? 3'b100 : 3'b110;
								assign node237 = (inp[2]) ? 3'b100 : node238;
									assign node238 = (inp[8]) ? node244 : node239;
										assign node239 = (inp[1]) ? 3'b101 : node240;
											assign node240 = (inp[11]) ? 3'b111 : 3'b101;
										assign node244 = (inp[1]) ? 3'b100 : 3'b101;
							assign node248 = (inp[8]) ? node262 : node249;
								assign node249 = (inp[10]) ? node257 : node250;
									assign node250 = (inp[11]) ? 3'b101 : node251;
										assign node251 = (inp[1]) ? 3'b100 : node252;
											assign node252 = (inp[9]) ? 3'b100 : 3'b101;
									assign node257 = (inp[2]) ? node259 : 3'b110;
										assign node259 = (inp[11]) ? 3'b110 : 3'b111;
								assign node262 = (inp[1]) ? node276 : node263;
									assign node263 = (inp[9]) ? node269 : node264;
										assign node264 = (inp[10]) ? 3'b110 : node265;
											assign node265 = (inp[2]) ? 3'b111 : 3'b110;
										assign node269 = (inp[10]) ? 3'b111 : node270;
											assign node270 = (inp[11]) ? node272 : 3'b110;
												assign node272 = (inp[2]) ? 3'b111 : 3'b110;
									assign node276 = (inp[2]) ? node278 : 3'b111;
										assign node278 = (inp[9]) ? 3'b110 : 3'b111;
						assign node281 = (inp[7]) ? node309 : node282;
							assign node282 = (inp[8]) ? node298 : node283;
								assign node283 = (inp[9]) ? node291 : node284;
									assign node284 = (inp[11]) ? node288 : node285;
										assign node285 = (inp[2]) ? 3'b110 : 3'b111;
										assign node288 = (inp[2]) ? 3'b111 : 3'b110;
									assign node291 = (inp[10]) ? node295 : node292;
										assign node292 = (inp[2]) ? 3'b101 : 3'b100;
										assign node295 = (inp[2]) ? 3'b100 : 3'b111;
								assign node298 = (inp[10]) ? 3'b111 : node299;
									assign node299 = (inp[9]) ? node303 : node300;
										assign node300 = (inp[2]) ? 3'b110 : 3'b111;
										assign node303 = (inp[1]) ? 3'b110 : node304;
											assign node304 = (inp[2]) ? 3'b111 : 3'b110;
							assign node309 = (inp[10]) ? node323 : node310;
								assign node310 = (inp[8]) ? node320 : node311;
									assign node311 = (inp[1]) ? node313 : 3'b111;
										assign node313 = (inp[11]) ? 3'b110 : node314;
											assign node314 = (inp[9]) ? 3'b111 : node315;
												assign node315 = (inp[2]) ? 3'b111 : 3'b110;
									assign node320 = (inp[2]) ? 3'b101 : 3'b100;
								assign node323 = (inp[11]) ? node329 : node324;
									assign node324 = (inp[9]) ? node326 : 3'b100;
										assign node326 = (inp[2]) ? 3'b100 : 3'b101;
									assign node329 = (inp[2]) ? 3'b101 : node330;
										assign node330 = (inp[8]) ? 3'b100 : 3'b101;
					assign node334 = (inp[8]) ? node406 : node335;
						assign node335 = (inp[9]) ? node377 : node336;
							assign node336 = (inp[3]) ? node362 : node337;
								assign node337 = (inp[10]) ? node351 : node338;
									assign node338 = (inp[7]) ? node342 : node339;
										assign node339 = (inp[11]) ? 3'b111 : 3'b101;
										assign node342 = (inp[11]) ? node348 : node343;
											assign node343 = (inp[1]) ? 3'b101 : node344;
												assign node344 = (inp[2]) ? 3'b100 : 3'b101;
											assign node348 = (inp[1]) ? 3'b100 : 3'b101;
									assign node351 = (inp[1]) ? node359 : node352;
										assign node352 = (inp[2]) ? 3'b110 : node353;
											assign node353 = (inp[11]) ? node355 : 3'b111;
												assign node355 = (inp[7]) ? 3'b111 : 3'b100;
										assign node359 = (inp[7]) ? 3'b111 : 3'b101;
								assign node362 = (inp[10]) ? node372 : node363;
									assign node363 = (inp[1]) ? node365 : 3'b111;
										assign node365 = (inp[11]) ? 3'b111 : node366;
											assign node366 = (inp[7]) ? node368 : 3'b110;
												assign node368 = (inp[2]) ? 3'b110 : 3'b111;
									assign node372 = (inp[2]) ? node374 : 3'b101;
										assign node374 = (inp[7]) ? 3'b100 : 3'b110;
							assign node377 = (inp[3]) ? node389 : node378;
								assign node378 = (inp[10]) ? node384 : node379;
									assign node379 = (inp[11]) ? node381 : 3'b100;
										assign node381 = (inp[1]) ? 3'b110 : 3'b100;
									assign node384 = (inp[1]) ? 3'b110 : node385;
										assign node385 = (inp[7]) ? 3'b111 : 3'b110;
								assign node389 = (inp[10]) ? node399 : node390;
									assign node390 = (inp[1]) ? node396 : node391;
										assign node391 = (inp[7]) ? node393 : 3'b110;
											assign node393 = (inp[11]) ? 3'b110 : 3'b111;
										assign node396 = (inp[11]) ? 3'b101 : 3'b111;
									assign node399 = (inp[7]) ? node401 : 3'b111;
										assign node401 = (inp[1]) ? 3'b100 : node402;
											assign node402 = (inp[11]) ? 3'b100 : 3'b101;
						assign node406 = (inp[7]) ? node434 : node407;
							assign node407 = (inp[3]) ? node425 : node408;
								assign node408 = (inp[1]) ? node414 : node409;
									assign node409 = (inp[9]) ? 3'b101 : node410;
										assign node410 = (inp[2]) ? 3'b101 : 3'b100;
									assign node414 = (inp[9]) ? node420 : node415;
										assign node415 = (inp[11]) ? node417 : 3'b101;
											assign node417 = (inp[10]) ? 3'b100 : 3'b101;
										assign node420 = (inp[2]) ? node422 : 3'b100;
											assign node422 = (inp[10]) ? 3'b101 : 3'b100;
								assign node425 = (inp[11]) ? node431 : node426;
									assign node426 = (inp[1]) ? 3'b110 : node427;
										assign node427 = (inp[9]) ? 3'b111 : 3'b110;
									assign node431 = (inp[9]) ? 3'b110 : 3'b111;
							assign node434 = (inp[3]) ? node446 : node435;
								assign node435 = (inp[1]) ? node443 : node436;
									assign node436 = (inp[11]) ? 3'b111 : node437;
										assign node437 = (inp[9]) ? node439 : 3'b110;
											assign node439 = (inp[2]) ? 3'b110 : 3'b111;
									assign node443 = (inp[2]) ? 3'b111 : 3'b110;
								assign node446 = (inp[2]) ? 3'b100 : node447;
									assign node447 = (inp[9]) ? 3'b101 : node448;
										assign node448 = (inp[1]) ? node450 : 3'b100;
											assign node450 = (inp[11]) ? node452 : 3'b101;
												assign node452 = (inp[10]) ? 3'b101 : 3'b100;
			assign node457 = (inp[5]) ? node667 : node458;
				assign node458 = (inp[8]) ? node570 : node459;
					assign node459 = (inp[10]) ? node521 : node460;
						assign node460 = (inp[3]) ? node488 : node461;
							assign node461 = (inp[11]) ? node467 : node462;
								assign node462 = (inp[7]) ? 3'b110 : node463;
									assign node463 = (inp[2]) ? 3'b100 : 3'b101;
								assign node467 = (inp[9]) ? node475 : node468;
									assign node468 = (inp[1]) ? 3'b100 : node469;
										assign node469 = (inp[7]) ? 3'b101 : node470;
											assign node470 = (inp[0]) ? 3'b101 : 3'b100;
									assign node475 = (inp[1]) ? node483 : node476;
										assign node476 = (inp[0]) ? node480 : node477;
											assign node477 = (inp[7]) ? 3'b100 : 3'b101;
											assign node480 = (inp[7]) ? 3'b101 : 3'b100;
										assign node483 = (inp[7]) ? 3'b101 : node484;
											assign node484 = (inp[0]) ? 3'b101 : 3'b100;
							assign node488 = (inp[7]) ? node506 : node489;
								assign node489 = (inp[11]) ? node497 : node490;
									assign node490 = (inp[0]) ? 3'b110 : node491;
										assign node491 = (inp[2]) ? node493 : 3'b111;
											assign node493 = (inp[1]) ? 3'b110 : 3'b111;
									assign node497 = (inp[2]) ? node499 : 3'b111;
										assign node499 = (inp[9]) ? node503 : node500;
											assign node500 = (inp[0]) ? 3'b111 : 3'b110;
											assign node503 = (inp[0]) ? 3'b110 : 3'b111;
								assign node506 = (inp[11]) ? node514 : node507;
									assign node507 = (inp[9]) ? 3'b101 : node508;
										assign node508 = (inp[0]) ? 3'b100 : node509;
											assign node509 = (inp[1]) ? 3'b101 : 3'b100;
									assign node514 = (inp[2]) ? 3'b110 : node515;
										assign node515 = (inp[1]) ? node517 : 3'b110;
											assign node517 = (inp[0]) ? 3'b111 : 3'b110;
						assign node521 = (inp[3]) ? node547 : node522;
							assign node522 = (inp[7]) ? node538 : node523;
								assign node523 = (inp[1]) ? node525 : 3'b110;
									assign node525 = (inp[0]) ? node533 : node526;
										assign node526 = (inp[2]) ? node528 : 3'b110;
											assign node528 = (inp[9]) ? 3'b110 : node529;
												assign node529 = (inp[11]) ? 3'b111 : 3'b110;
										assign node533 = (inp[11]) ? node535 : 3'b111;
											assign node535 = (inp[9]) ? 3'b111 : 3'b110;
								assign node538 = (inp[11]) ? node540 : 3'b101;
									assign node540 = (inp[2]) ? 3'b111 : node541;
										assign node541 = (inp[9]) ? node543 : 3'b110;
											assign node543 = (inp[0]) ? 3'b110 : 3'b111;
							assign node547 = (inp[7]) ? node559 : node548;
								assign node548 = (inp[0]) ? 3'b100 : node549;
									assign node549 = (inp[2]) ? 3'b100 : node550;
										assign node550 = (inp[9]) ? node552 : 3'b100;
											assign node552 = (inp[11]) ? 3'b101 : node553;
												assign node553 = (inp[1]) ? 3'b101 : 3'b100;
								assign node559 = (inp[11]) ? node565 : node560;
									assign node560 = (inp[9]) ? 3'b110 : node561;
										assign node561 = (inp[0]) ? 3'b111 : 3'b110;
									assign node565 = (inp[1]) ? node567 : 3'b100;
										assign node567 = (inp[0]) ? 3'b101 : 3'b100;
					assign node570 = (inp[10]) ? node614 : node571;
						assign node571 = (inp[9]) ? node595 : node572;
							assign node572 = (inp[2]) ? node584 : node573;
								assign node573 = (inp[7]) ? node577 : node574;
									assign node574 = (inp[3]) ? 3'b000 : 3'b010;
									assign node577 = (inp[0]) ? node581 : node578;
										assign node578 = (inp[1]) ? 3'b000 : 3'b011;
										assign node581 = (inp[11]) ? 3'b011 : 3'b000;
								assign node584 = (inp[1]) ? node588 : node585;
									assign node585 = (inp[3]) ? 3'b001 : 3'b011;
									assign node588 = (inp[7]) ? node592 : node589;
										assign node589 = (inp[0]) ? 3'b001 : 3'b010;
										assign node592 = (inp[3]) ? 3'b010 : 3'b001;
							assign node595 = (inp[3]) ? node605 : node596;
								assign node596 = (inp[11]) ? node602 : node597;
									assign node597 = (inp[2]) ? node599 : 3'b001;
										assign node599 = (inp[1]) ? 3'b001 : 3'b000;
									assign node602 = (inp[0]) ? 3'b011 : 3'b010;
								assign node605 = (inp[11]) ? node611 : node606;
									assign node606 = (inp[7]) ? node608 : 3'b011;
										assign node608 = (inp[2]) ? 3'b011 : 3'b010;
									assign node611 = (inp[2]) ? 3'b000 : 3'b001;
						assign node614 = (inp[0]) ? node640 : node615;
							assign node615 = (inp[2]) ? node631 : node616;
								assign node616 = (inp[1]) ? node622 : node617;
									assign node617 = (inp[11]) ? node619 : 3'b000;
										assign node619 = (inp[3]) ? 3'b001 : 3'b011;
									assign node622 = (inp[7]) ? node628 : node623;
										assign node623 = (inp[3]) ? 3'b011 : node624;
											assign node624 = (inp[9]) ? 3'b011 : 3'b010;
										assign node628 = (inp[9]) ? 3'b010 : 3'b000;
								assign node631 = (inp[9]) ? node633 : 3'b010;
									assign node633 = (inp[11]) ? node637 : node634;
										assign node634 = (inp[3]) ? 3'b010 : 3'b000;
										assign node637 = (inp[3]) ? 3'b000 : 3'b010;
							assign node640 = (inp[9]) ? node652 : node641;
								assign node641 = (inp[11]) ? node645 : node642;
									assign node642 = (inp[3]) ? 3'b011 : 3'b001;
									assign node645 = (inp[3]) ? node649 : node646;
										assign node646 = (inp[7]) ? 3'b011 : 3'b010;
										assign node649 = (inp[2]) ? 3'b001 : 3'b000;
								assign node652 = (inp[2]) ? node660 : node653;
									assign node653 = (inp[3]) ? node657 : node654;
										assign node654 = (inp[11]) ? 3'b011 : 3'b000;
										assign node657 = (inp[1]) ? 3'b011 : 3'b001;
									assign node660 = (inp[1]) ? node662 : 3'b000;
										assign node662 = (inp[11]) ? node664 : 3'b010;
											assign node664 = (inp[7]) ? 3'b010 : 3'b000;
				assign node667 = (inp[3]) ? node757 : node668;
					assign node668 = (inp[8]) ? node732 : node669;
						assign node669 = (inp[10]) ? node707 : node670;
							assign node670 = (inp[11]) ? node692 : node671;
								assign node671 = (inp[7]) ? node683 : node672;
									assign node672 = (inp[2]) ? node678 : node673;
										assign node673 = (inp[0]) ? node675 : 3'b010;
											assign node675 = (inp[1]) ? 3'b011 : 3'b010;
										assign node678 = (inp[0]) ? 3'b011 : node679;
											assign node679 = (inp[9]) ? 3'b010 : 3'b011;
									assign node683 = (inp[9]) ? node689 : node684;
										assign node684 = (inp[2]) ? 3'b000 : node685;
											assign node685 = (inp[0]) ? 3'b001 : 3'b000;
										assign node689 = (inp[2]) ? 3'b001 : 3'b000;
								assign node692 = (inp[0]) ? node704 : node693;
									assign node693 = (inp[1]) ? node695 : 3'b000;
										assign node695 = (inp[7]) ? node697 : 3'b001;
											assign node697 = (inp[2]) ? node701 : node698;
												assign node698 = (inp[9]) ? 3'b000 : 3'b001;
												assign node701 = (inp[9]) ? 3'b001 : 3'b000;
									assign node704 = (inp[1]) ? 3'b000 : 3'b001;
							assign node707 = (inp[11]) ? node721 : node708;
								assign node708 = (inp[7]) ? 3'b011 : node709;
									assign node709 = (inp[1]) ? node715 : node710;
										assign node710 = (inp[0]) ? node712 : 3'b001;
											assign node712 = (inp[9]) ? 3'b000 : 3'b001;
										assign node715 = (inp[0]) ? node717 : 3'b000;
											assign node717 = (inp[9]) ? 3'b000 : 3'b001;
								assign node721 = (inp[7]) ? node723 : 3'b011;
									assign node723 = (inp[0]) ? 3'b010 : node724;
										assign node724 = (inp[9]) ? 3'b011 : node725;
											assign node725 = (inp[1]) ? 3'b010 : node726;
												assign node726 = (inp[2]) ? 3'b010 : 3'b011;
						assign node732 = (inp[7]) ? node746 : node733;
							assign node733 = (inp[9]) ? node741 : node734;
								assign node734 = (inp[1]) ? 3'b010 : node735;
									assign node735 = (inp[0]) ? 3'b010 : node736;
										assign node736 = (inp[2]) ? 3'b011 : 3'b010;
								assign node741 = (inp[11]) ? 3'b011 : node742;
									assign node742 = (inp[1]) ? 3'b010 : 3'b011;
							assign node746 = (inp[9]) ? node752 : node747;
								assign node747 = (inp[11]) ? 3'b011 : node748;
									assign node748 = (inp[10]) ? 3'b011 : 3'b010;
								assign node752 = (inp[11]) ? 3'b010 : node753;
									assign node753 = (inp[10]) ? 3'b010 : 3'b011;
					assign node757 = (inp[8]) ? node807 : node758;
						assign node758 = (inp[10]) ? node780 : node759;
							assign node759 = (inp[1]) ? node773 : node760;
								assign node760 = (inp[7]) ? node764 : node761;
									assign node761 = (inp[0]) ? 3'b010 : 3'b000;
									assign node764 = (inp[11]) ? 3'b010 : node765;
										assign node765 = (inp[9]) ? 3'b011 : node766;
											assign node766 = (inp[2]) ? 3'b010 : node767;
												assign node767 = (inp[0]) ? 3'b011 : 3'b010;
								assign node773 = (inp[7]) ? node777 : node774;
									assign node774 = (inp[11]) ? 3'b011 : 3'b001;
									assign node777 = (inp[9]) ? 3'b010 : 3'b011;
							assign node780 = (inp[7]) ? node794 : node781;
								assign node781 = (inp[11]) ? node791 : node782;
									assign node782 = (inp[1]) ? node784 : 3'b011;
										assign node784 = (inp[0]) ? node788 : node785;
											assign node785 = (inp[9]) ? 3'b010 : 3'b011;
											assign node788 = (inp[9]) ? 3'b011 : 3'b010;
									assign node791 = (inp[9]) ? 3'b000 : 3'b001;
								assign node794 = (inp[1]) ? node802 : node795;
									assign node795 = (inp[2]) ? node797 : 3'b000;
										assign node797 = (inp[9]) ? node799 : 3'b000;
											assign node799 = (inp[0]) ? 3'b000 : 3'b001;
									assign node802 = (inp[0]) ? 3'b001 : node803;
										assign node803 = (inp[9]) ? 3'b001 : 3'b000;
						assign node807 = (inp[9]) ? node823 : node808;
							assign node808 = (inp[11]) ? 3'b001 : node809;
								assign node809 = (inp[0]) ? node815 : node810;
									assign node810 = (inp[10]) ? node812 : 3'b000;
										assign node812 = (inp[7]) ? 3'b001 : 3'b000;
									assign node815 = (inp[2]) ? node819 : node816;
										assign node816 = (inp[1]) ? 3'b000 : 3'b001;
										assign node819 = (inp[1]) ? 3'b001 : 3'b000;
							assign node823 = (inp[11]) ? 3'b000 : node824;
								assign node824 = (inp[0]) ? node826 : 3'b001;
									assign node826 = (inp[10]) ? node830 : node827;
										assign node827 = (inp[2]) ? 3'b001 : 3'b000;
										assign node830 = (inp[2]) ? 3'b000 : 3'b001;
		assign node834 = (inp[5]) ? node1144 : node835;
			assign node835 = (inp[8]) ? node999 : node836;
				assign node836 = (inp[10]) ? node920 : node837;
					assign node837 = (inp[11]) ? node879 : node838;
						assign node838 = (inp[6]) ? node858 : node839;
							assign node839 = (inp[1]) ? node851 : node840;
								assign node840 = (inp[7]) ? node842 : 3'b101;
									assign node842 = (inp[3]) ? 3'b100 : node843;
										assign node843 = (inp[0]) ? node847 : node844;
											assign node844 = (inp[2]) ? 3'b101 : 3'b100;
											assign node847 = (inp[2]) ? 3'b100 : 3'b101;
								assign node851 = (inp[0]) ? 3'b100 : node852;
									assign node852 = (inp[2]) ? 3'b101 : node853;
										assign node853 = (inp[3]) ? 3'b101 : 3'b100;
							assign node858 = (inp[0]) ? node870 : node859;
								assign node859 = (inp[7]) ? node861 : 3'b100;
									assign node861 = (inp[3]) ? node865 : node862;
										assign node862 = (inp[2]) ? 3'b101 : 3'b100;
										assign node865 = (inp[2]) ? 3'b100 : node866;
											assign node866 = (inp[1]) ? 3'b101 : 3'b100;
								assign node870 = (inp[3]) ? node874 : node871;
									assign node871 = (inp[1]) ? 3'b100 : 3'b101;
									assign node874 = (inp[2]) ? node876 : 3'b101;
										assign node876 = (inp[7]) ? 3'b101 : 3'b100;
						assign node879 = (inp[9]) ? node905 : node880;
							assign node880 = (inp[1]) ? node890 : node881;
								assign node881 = (inp[6]) ? 3'b110 : node882;
									assign node882 = (inp[2]) ? node886 : node883;
										assign node883 = (inp[0]) ? 3'b111 : 3'b110;
										assign node886 = (inp[0]) ? 3'b110 : 3'b111;
								assign node890 = (inp[6]) ? node900 : node891;
									assign node891 = (inp[2]) ? node893 : 3'b110;
										assign node893 = (inp[3]) ? 3'b110 : node894;
											assign node894 = (inp[0]) ? node896 : 3'b111;
												assign node896 = (inp[7]) ? 3'b111 : 3'b110;
									assign node900 = (inp[7]) ? node902 : 3'b111;
										assign node902 = (inp[2]) ? 3'b110 : 3'b111;
							assign node905 = (inp[3]) ? node911 : node906;
								assign node906 = (inp[6]) ? 3'b111 : node907;
									assign node907 = (inp[0]) ? 3'b110 : 3'b111;
								assign node911 = (inp[2]) ? 3'b110 : node912;
									assign node912 = (inp[0]) ? node914 : 3'b110;
										assign node914 = (inp[7]) ? 3'b111 : node915;
											assign node915 = (inp[6]) ? 3'b111 : 3'b110;
					assign node920 = (inp[11]) ? node960 : node921;
						assign node921 = (inp[0]) ? node947 : node922;
							assign node922 = (inp[2]) ? node940 : node923;
								assign node923 = (inp[1]) ? 3'b110 : node924;
									assign node924 = (inp[6]) ? node930 : node925;
										assign node925 = (inp[7]) ? node927 : 3'b110;
											assign node927 = (inp[3]) ? 3'b111 : 3'b110;
										assign node930 = (inp[9]) ? node934 : node931;
											assign node931 = (inp[3]) ? 3'b111 : 3'b110;
											assign node934 = (inp[7]) ? node936 : 3'b111;
												assign node936 = (inp[3]) ? 3'b110 : 3'b111;
								assign node940 = (inp[1]) ? 3'b111 : node941;
									assign node941 = (inp[9]) ? 3'b111 : node942;
										assign node942 = (inp[6]) ? 3'b111 : 3'b110;
							assign node947 = (inp[1]) ? 3'b111 : node948;
								assign node948 = (inp[6]) ? node954 : node949;
									assign node949 = (inp[2]) ? node951 : 3'b111;
										assign node951 = (inp[3]) ? 3'b111 : 3'b110;
									assign node954 = (inp[2]) ? 3'b111 : node955;
										assign node955 = (inp[3]) ? 3'b110 : 3'b111;
						assign node960 = (inp[2]) ? node976 : node961;
							assign node961 = (inp[0]) ? node967 : node962;
								assign node962 = (inp[3]) ? 3'b100 : node963;
									assign node963 = (inp[9]) ? 3'b100 : 3'b101;
								assign node967 = (inp[9]) ? 3'b101 : node968;
									assign node968 = (inp[6]) ? 3'b100 : node969;
										assign node969 = (inp[3]) ? node971 : 3'b101;
											assign node971 = (inp[7]) ? 3'b100 : 3'b101;
							assign node976 = (inp[0]) ? node986 : node977;
								assign node977 = (inp[9]) ? 3'b101 : node978;
									assign node978 = (inp[6]) ? 3'b100 : node979;
										assign node979 = (inp[1]) ? 3'b101 : node980;
											assign node980 = (inp[7]) ? 3'b101 : 3'b100;
								assign node986 = (inp[3]) ? node994 : node987;
									assign node987 = (inp[1]) ? node991 : node988;
										assign node988 = (inp[7]) ? 3'b101 : 3'b100;
										assign node991 = (inp[7]) ? 3'b100 : 3'b101;
									assign node994 = (inp[1]) ? 3'b100 : node995;
										assign node995 = (inp[7]) ? 3'b101 : 3'b100;
				assign node999 = (inp[11]) ? node1101 : node1000;
					assign node1000 = (inp[7]) ? node1046 : node1001;
						assign node1001 = (inp[6]) ? node1021 : node1002;
							assign node1002 = (inp[9]) ? node1012 : node1003;
								assign node1003 = (inp[2]) ? node1005 : 3'b001;
									assign node1005 = (inp[0]) ? node1009 : node1006;
										assign node1006 = (inp[3]) ? 3'b000 : 3'b001;
										assign node1009 = (inp[10]) ? 3'b001 : 3'b000;
								assign node1012 = (inp[3]) ? 3'b000 : node1013;
									assign node1013 = (inp[2]) ? node1017 : node1014;
										assign node1014 = (inp[1]) ? 3'b001 : 3'b000;
										assign node1017 = (inp[1]) ? 3'b000 : 3'b001;
							assign node1021 = (inp[9]) ? node1037 : node1022;
								assign node1022 = (inp[0]) ? node1032 : node1023;
									assign node1023 = (inp[3]) ? node1025 : 3'b011;
										assign node1025 = (inp[2]) ? node1029 : node1026;
											assign node1026 = (inp[10]) ? 3'b011 : 3'b010;
											assign node1029 = (inp[10]) ? 3'b010 : 3'b011;
									assign node1032 = (inp[10]) ? node1034 : 3'b010;
										assign node1034 = (inp[2]) ? 3'b010 : 3'b011;
								assign node1037 = (inp[3]) ? 3'b011 : node1038;
									assign node1038 = (inp[0]) ? 3'b011 : node1039;
										assign node1039 = (inp[1]) ? 3'b010 : node1040;
											assign node1040 = (inp[2]) ? 3'b011 : 3'b010;
						assign node1046 = (inp[0]) ? node1072 : node1047;
							assign node1047 = (inp[3]) ? node1063 : node1048;
								assign node1048 = (inp[9]) ? node1050 : 3'b010;
									assign node1050 = (inp[1]) ? node1060 : node1051;
										assign node1051 = (inp[2]) ? node1057 : node1052;
											assign node1052 = (inp[10]) ? node1054 : 3'b010;
												assign node1054 = (inp[6]) ? 3'b011 : 3'b010;
											assign node1057 = (inp[10]) ? 3'b010 : 3'b011;
										assign node1060 = (inp[2]) ? 3'b010 : 3'b011;
								assign node1063 = (inp[10]) ? 3'b010 : node1064;
									assign node1064 = (inp[2]) ? 3'b011 : node1065;
										assign node1065 = (inp[1]) ? 3'b010 : node1066;
											assign node1066 = (inp[6]) ? 3'b010 : 3'b011;
							assign node1072 = (inp[10]) ? node1086 : node1073;
								assign node1073 = (inp[2]) ? node1079 : node1074;
									assign node1074 = (inp[1]) ? node1076 : 3'b010;
										assign node1076 = (inp[6]) ? 3'b010 : 3'b011;
									assign node1079 = (inp[6]) ? 3'b011 : node1080;
										assign node1080 = (inp[9]) ? 3'b010 : node1081;
											assign node1081 = (inp[1]) ? 3'b010 : 3'b011;
								assign node1086 = (inp[9]) ? node1092 : node1087;
									assign node1087 = (inp[1]) ? node1089 : 3'b011;
										assign node1089 = (inp[2]) ? 3'b010 : 3'b011;
									assign node1092 = (inp[3]) ? 3'b010 : node1093;
										assign node1093 = (inp[2]) ? node1097 : node1094;
											assign node1094 = (inp[1]) ? 3'b011 : 3'b010;
											assign node1097 = (inp[6]) ? 3'b010 : 3'b011;
					assign node1101 = (inp[6]) ? node1133 : node1102;
						assign node1102 = (inp[7]) ? node1116 : node1103;
							assign node1103 = (inp[1]) ? node1109 : node1104;
								assign node1104 = (inp[2]) ? 3'b011 : node1105;
									assign node1105 = (inp[3]) ? 3'b010 : 3'b011;
								assign node1109 = (inp[2]) ? 3'b010 : node1110;
									assign node1110 = (inp[10]) ? node1112 : 3'b011;
										assign node1112 = (inp[9]) ? 3'b011 : 3'b010;
							assign node1116 = (inp[10]) ? node1122 : node1117;
								assign node1117 = (inp[9]) ? node1119 : 3'b001;
									assign node1119 = (inp[1]) ? 3'b000 : 3'b001;
								assign node1122 = (inp[9]) ? node1128 : node1123;
									assign node1123 = (inp[2]) ? node1125 : 3'b000;
										assign node1125 = (inp[1]) ? 3'b000 : 3'b001;
									assign node1128 = (inp[1]) ? 3'b001 : node1129;
										assign node1129 = (inp[2]) ? 3'b001 : 3'b000;
						assign node1133 = (inp[2]) ? node1139 : node1134;
							assign node1134 = (inp[3]) ? 3'b001 : node1135;
								assign node1135 = (inp[7]) ? 3'b001 : 3'b000;
							assign node1139 = (inp[7]) ? 3'b000 : node1140;
								assign node1140 = (inp[3]) ? 3'b000 : 3'b001;
			assign node1144 = (inp[6]) ? node1250 : node1145;
				assign node1145 = (inp[7]) ? node1203 : node1146;
					assign node1146 = (inp[10]) ? node1176 : node1147;
						assign node1147 = (inp[8]) ? node1169 : node1148;
							assign node1148 = (inp[1]) ? node1156 : node1149;
								assign node1149 = (inp[0]) ? node1153 : node1150;
									assign node1150 = (inp[3]) ? 3'b001 : 3'b000;
									assign node1153 = (inp[3]) ? 3'b000 : 3'b001;
								assign node1156 = (inp[11]) ? node1162 : node1157;
									assign node1157 = (inp[0]) ? node1159 : 3'b000;
										assign node1159 = (inp[2]) ? 3'b000 : 3'b001;
									assign node1162 = (inp[0]) ? node1166 : node1163;
										assign node1163 = (inp[3]) ? 3'b000 : 3'b001;
										assign node1166 = (inp[3]) ? 3'b001 : 3'b000;
							assign node1169 = (inp[3]) ? node1173 : node1170;
								assign node1170 = (inp[1]) ? 3'b011 : 3'b010;
								assign node1173 = (inp[1]) ? 3'b010 : 3'b011;
						assign node1176 = (inp[1]) ? node1192 : node1177;
							assign node1177 = (inp[3]) ? node1185 : node1178;
								assign node1178 = (inp[11]) ? node1180 : 3'b010;
									assign node1180 = (inp[8]) ? 3'b010 : node1181;
										assign node1181 = (inp[0]) ? 3'b010 : 3'b011;
								assign node1185 = (inp[8]) ? 3'b011 : node1186;
									assign node1186 = (inp[11]) ? 3'b010 : node1187;
										assign node1187 = (inp[0]) ? 3'b010 : 3'b011;
							assign node1192 = (inp[3]) ? node1198 : node1193;
								assign node1193 = (inp[8]) ? 3'b011 : node1194;
									assign node1194 = (inp[0]) ? 3'b011 : 3'b010;
								assign node1198 = (inp[8]) ? 3'b010 : node1199;
									assign node1199 = (inp[0]) ? 3'b010 : 3'b011;
					assign node1203 = (inp[8]) ? node1239 : node1204;
						assign node1204 = (inp[10]) ? node1212 : node1205;
							assign node1205 = (inp[11]) ? node1209 : node1206;
								assign node1206 = (inp[0]) ? 3'b011 : 3'b010;
								assign node1209 = (inp[0]) ? 3'b010 : 3'b011;
							assign node1212 = (inp[11]) ? node1226 : node1213;
								assign node1213 = (inp[2]) ? node1217 : node1214;
									assign node1214 = (inp[9]) ? 3'b001 : 3'b000;
									assign node1217 = (inp[3]) ? node1219 : 3'b001;
										assign node1219 = (inp[1]) ? node1223 : node1220;
											assign node1220 = (inp[9]) ? 3'b000 : 3'b001;
											assign node1223 = (inp[0]) ? 3'b000 : 3'b001;
								assign node1226 = (inp[3]) ? node1232 : node1227;
									assign node1227 = (inp[2]) ? 3'b000 : node1228;
										assign node1228 = (inp[0]) ? 3'b000 : 3'b001;
									assign node1232 = (inp[9]) ? node1234 : 3'b000;
										assign node1234 = (inp[1]) ? node1236 : 3'b001;
											assign node1236 = (inp[0]) ? 3'b000 : 3'b001;
						assign node1239 = (inp[1]) ? node1245 : node1240;
							assign node1240 = (inp[10]) ? 3'b001 : node1241;
								assign node1241 = (inp[11]) ? 3'b001 : 3'b000;
							assign node1245 = (inp[11]) ? 3'b000 : node1246;
								assign node1246 = (inp[10]) ? 3'b000 : 3'b001;
				assign node1250 = (inp[8]) ? node1310 : node1251;
					assign node1251 = (inp[10]) ? node1295 : node1252;
						assign node1252 = (inp[7]) ? node1276 : node1253;
							assign node1253 = (inp[2]) ? node1263 : node1254;
								assign node1254 = (inp[11]) ? node1260 : node1255;
									assign node1255 = (inp[3]) ? node1257 : 3'b010;
										assign node1257 = (inp[9]) ? 3'b011 : 3'b010;
									assign node1260 = (inp[1]) ? 3'b011 : 3'b010;
								assign node1263 = (inp[9]) ? node1273 : node1264;
									assign node1264 = (inp[1]) ? node1266 : 3'b011;
										assign node1266 = (inp[11]) ? node1268 : 3'b011;
											assign node1268 = (inp[3]) ? 3'b010 : node1269;
												assign node1269 = (inp[0]) ? 3'b011 : 3'b010;
									assign node1273 = (inp[3]) ? 3'b010 : 3'b011;
							assign node1276 = (inp[3]) ? node1282 : node1277;
								assign node1277 = (inp[0]) ? node1279 : 3'b011;
									assign node1279 = (inp[11]) ? 3'b010 : 3'b011;
								assign node1282 = (inp[2]) ? node1290 : node1283;
									assign node1283 = (inp[11]) ? node1287 : node1284;
										assign node1284 = (inp[0]) ? 3'b011 : 3'b010;
										assign node1287 = (inp[0]) ? 3'b010 : 3'b011;
									assign node1290 = (inp[11]) ? 3'b010 : node1291;
										assign node1291 = (inp[0]) ? 3'b011 : 3'b010;
						assign node1295 = (inp[0]) ? node1305 : node1296;
							assign node1296 = (inp[7]) ? 3'b001 : node1297;
								assign node1297 = (inp[3]) ? 3'b001 : node1298;
									assign node1298 = (inp[1]) ? 3'b000 : node1299;
										assign node1299 = (inp[11]) ? 3'b000 : 3'b001;
							assign node1305 = (inp[3]) ? 3'b000 : node1306;
								assign node1306 = (inp[11]) ? 3'b001 : 3'b000;
					assign node1310 = (inp[3]) ? node1358 : node1311;
						assign node1311 = (inp[9]) ? node1335 : node1312;
							assign node1312 = (inp[10]) ? node1332 : node1313;
								assign node1313 = (inp[0]) ? node1323 : node1314;
									assign node1314 = (inp[2]) ? node1316 : 3'b000;
										assign node1316 = (inp[7]) ? node1320 : node1317;
											assign node1317 = (inp[11]) ? 3'b001 : 3'b000;
											assign node1320 = (inp[11]) ? 3'b000 : 3'b001;
									assign node1323 = (inp[2]) ? 3'b001 : node1324;
										assign node1324 = (inp[7]) ? node1328 : node1325;
											assign node1325 = (inp[11]) ? 3'b001 : 3'b000;
											assign node1328 = (inp[11]) ? 3'b000 : 3'b001;
								assign node1332 = (inp[7]) ? 3'b000 : 3'b001;
							assign node1335 = (inp[2]) ? node1347 : node1336;
								assign node1336 = (inp[10]) ? node1344 : node1337;
									assign node1337 = (inp[11]) ? node1341 : node1338;
										assign node1338 = (inp[7]) ? 3'b001 : 3'b000;
										assign node1341 = (inp[7]) ? 3'b000 : 3'b001;
									assign node1344 = (inp[7]) ? 3'b000 : 3'b001;
								assign node1347 = (inp[10]) ? 3'b000 : node1348;
									assign node1348 = (inp[1]) ? node1352 : node1349;
										assign node1349 = (inp[0]) ? 3'b001 : 3'b000;
										assign node1352 = (inp[0]) ? 3'b000 : node1353;
											assign node1353 = (inp[7]) ? 3'b001 : 3'b000;
						assign node1358 = (inp[10]) ? 3'b000 : node1359;
							assign node1359 = (inp[11]) ? 3'b000 : 3'b001;

endmodule