module dtc_split5_bm97 (
	input  wire [12-1:0] inp,
	output wire [3-1:0] outp
);

	wire [3-1:0] node1;
	wire [3-1:0] node3;
	wire [3-1:0] node5;
	wire [3-1:0] node7;
	wire [3-1:0] node9;
	wire [3-1:0] node10;
	wire [3-1:0] node12;
	wire [3-1:0] node13;
	wire [3-1:0] node15;
	wire [3-1:0] node18;
	wire [3-1:0] node20;
	wire [3-1:0] node23;
	wire [3-1:0] node25;
	wire [3-1:0] node26;
	wire [3-1:0] node29;
	wire [3-1:0] node30;
	wire [3-1:0] node32;
	wire [3-1:0] node35;
	wire [3-1:0] node37;
	wire [3-1:0] node40;
	wire [3-1:0] node41;
	wire [3-1:0] node42;
	wire [3-1:0] node43;
	wire [3-1:0] node45;
	wire [3-1:0] node46;
	wire [3-1:0] node48;
	wire [3-1:0] node49;
	wire [3-1:0] node51;
	wire [3-1:0] node55;
	wire [3-1:0] node56;
	wire [3-1:0] node58;
	wire [3-1:0] node59;
	wire [3-1:0] node63;
	wire [3-1:0] node64;
	wire [3-1:0] node66;
	wire [3-1:0] node67;
	wire [3-1:0] node74;
	wire [3-1:0] node75;
	wire [3-1:0] node76;
	wire [3-1:0] node79;
	wire [3-1:0] node81;
	wire [3-1:0] node82;
	wire [3-1:0] node84;
	wire [3-1:0] node86;
	wire [3-1:0] node88;
	wire [3-1:0] node91;
	wire [3-1:0] node93;
	wire [3-1:0] node95;
	wire [3-1:0] node96;
	wire [3-1:0] node97;
	wire [3-1:0] node102;
	wire [3-1:0] node103;
	wire [3-1:0] node104;
	wire [3-1:0] node105;
	wire [3-1:0] node107;
	wire [3-1:0] node110;
	wire [3-1:0] node111;
	wire [3-1:0] node112;
	wire [3-1:0] node114;
	wire [3-1:0] node118;
	wire [3-1:0] node119;
	wire [3-1:0] node121;
	wire [3-1:0] node122;
	wire [3-1:0] node127;
	wire [3-1:0] node129;
	wire [3-1:0] node131;
	wire [3-1:0] node132;
	wire [3-1:0] node134;
	wire [3-1:0] node138;
	wire [3-1:0] node140;
	wire [3-1:0] node142;
	wire [3-1:0] node143;
	wire [3-1:0] node144;
	wire [3-1:0] node146;
	wire [3-1:0] node148;
	wire [3-1:0] node152;

	assign outp = (inp[3]) ? node40 : node1;
		assign node1 = (inp[6]) ? node3 : 3'b000;
			assign node3 = (inp[9]) ? node5 : 3'b000;
				assign node5 = (inp[7]) ? node7 : 3'b001;
					assign node7 = (inp[10]) ? node9 : 3'b000;
						assign node9 = (inp[4]) ? node23 : node10;
							assign node10 = (inp[11]) ? node12 : 3'b000;
								assign node12 = (inp[8]) ? node18 : node13;
									assign node13 = (inp[5]) ? node15 : 3'b000;
										assign node15 = (inp[1]) ? 3'b101 : 3'b001;
									assign node18 = (inp[5]) ? node20 : 3'b100;
										assign node20 = (inp[2]) ? 3'b100 : 3'b101;
							assign node23 = (inp[11]) ? node25 : 3'b100;
								assign node25 = (inp[5]) ? node29 : node26;
									assign node26 = (inp[8]) ? 3'b100 : 3'b000;
									assign node29 = (inp[8]) ? node35 : node30;
										assign node30 = (inp[0]) ? node32 : 3'b010;
											assign node32 = (inp[1]) ? 3'b110 : 3'b010;
										assign node35 = (inp[0]) ? node37 : 3'b100;
											assign node37 = (inp[1]) ? 3'b010 : 3'b110;
		assign node40 = (inp[9]) ? node74 : node41;
			assign node41 = (inp[6]) ? 3'b000 : node42;
				assign node42 = (inp[7]) ? 3'b000 : node43;
					assign node43 = (inp[4]) ? node45 : 3'b100;
						assign node45 = (inp[11]) ? node55 : node46;
							assign node46 = (inp[10]) ? node48 : 3'b100;
								assign node48 = (inp[8]) ? 3'b100 : node49;
									assign node49 = (inp[5]) ? node51 : 3'b000;
										assign node51 = (inp[2]) ? 3'b100 : 3'b000;
							assign node55 = (inp[5]) ? node63 : node56;
								assign node56 = (inp[10]) ? node58 : 3'b100;
									assign node58 = (inp[8]) ? 3'b000 : node59;
										assign node59 = (inp[0]) ? 3'b000 : 3'b100;
								assign node63 = (inp[0]) ? 3'b000 : node64;
									assign node64 = (inp[2]) ? node66 : 3'b000;
										assign node66 = (inp[1]) ? 3'b000 : node67;
											assign node67 = (inp[10]) ? 3'b000 : 3'b000;
			assign node74 = (inp[4]) ? node102 : node75;
				assign node75 = (inp[6]) ? node79 : node76;
					assign node76 = (inp[7]) ? 3'b110 : 3'b000;
					assign node79 = (inp[7]) ? node81 : 3'b110;
						assign node81 = (inp[5]) ? node91 : node82;
							assign node82 = (inp[10]) ? node84 : 3'b000;
								assign node84 = (inp[2]) ? node86 : 3'b010;
									assign node86 = (inp[8]) ? node88 : 3'b010;
										assign node88 = (inp[1]) ? 3'b100 : 3'b010;
							assign node91 = (inp[11]) ? node93 : 3'b000;
								assign node93 = (inp[10]) ? node95 : 3'b000;
									assign node95 = (inp[0]) ? 3'b100 : node96;
										assign node96 = (inp[1]) ? 3'b100 : node97;
											assign node97 = (inp[2]) ? 3'b010 : 3'b100;
				assign node102 = (inp[6]) ? node138 : node103;
					assign node103 = (inp[7]) ? node127 : node104;
						assign node104 = (inp[10]) ? node110 : node105;
							assign node105 = (inp[11]) ? node107 : 3'b010;
								assign node107 = (inp[5]) ? 3'b110 : 3'b010;
							assign node110 = (inp[11]) ? node118 : node111;
								assign node111 = (inp[8]) ? 3'b001 : node112;
									assign node112 = (inp[2]) ? node114 : 3'b101;
										assign node114 = (inp[0]) ? 3'b101 : 3'b001;
								assign node118 = (inp[8]) ? 3'b101 : node119;
									assign node119 = (inp[0]) ? node121 : 3'b011;
										assign node121 = (inp[5]) ? 3'b101 : node122;
											assign node122 = (inp[1]) ? 3'b101 : 3'b011;
						assign node127 = (inp[11]) ? node129 : 3'b001;
							assign node129 = (inp[10]) ? node131 : 3'b001;
								assign node131 = (inp[8]) ? 3'b110 : node132;
									assign node132 = (inp[0]) ? node134 : 3'b001;
										assign node134 = (inp[5]) ? 3'b110 : 3'b001;
					assign node138 = (inp[11]) ? node140 : 3'b000;
						assign node140 = (inp[10]) ? node142 : 3'b000;
							assign node142 = (inp[8]) ? node152 : node143;
								assign node143 = (inp[7]) ? 3'b000 : node144;
									assign node144 = (inp[5]) ? node146 : 3'b010;
										assign node146 = (inp[0]) ? node148 : 3'b010;
											assign node148 = (inp[1]) ? 3'b100 : 3'b010;
								assign node152 = (inp[7]) ? 3'b000 : 3'b100;

endmodule