module dtc_split33_bm91 (
	input  wire [12-1:0] inp,
	output wire [3-1:0] outp
);

	wire [3-1:0] node1;
	wire [3-1:0] node2;
	wire [3-1:0] node3;
	wire [3-1:0] node4;
	wire [3-1:0] node5;
	wire [3-1:0] node6;
	wire [3-1:0] node7;
	wire [3-1:0] node8;
	wire [3-1:0] node10;
	wire [3-1:0] node13;
	wire [3-1:0] node15;
	wire [3-1:0] node18;
	wire [3-1:0] node19;
	wire [3-1:0] node20;
	wire [3-1:0] node23;
	wire [3-1:0] node26;
	wire [3-1:0] node28;
	wire [3-1:0] node31;
	wire [3-1:0] node33;
	wire [3-1:0] node35;
	wire [3-1:0] node38;
	wire [3-1:0] node39;
	wire [3-1:0] node40;
	wire [3-1:0] node42;
	wire [3-1:0] node43;
	wire [3-1:0] node47;
	wire [3-1:0] node48;
	wire [3-1:0] node49;
	wire [3-1:0] node54;
	wire [3-1:0] node56;
	wire [3-1:0] node57;
	wire [3-1:0] node58;
	wire [3-1:0] node62;
	wire [3-1:0] node64;
	wire [3-1:0] node67;
	wire [3-1:0] node68;
	wire [3-1:0] node69;
	wire [3-1:0] node71;
	wire [3-1:0] node72;
	wire [3-1:0] node75;
	wire [3-1:0] node77;
	wire [3-1:0] node80;
	wire [3-1:0] node82;
	wire [3-1:0] node85;
	wire [3-1:0] node86;
	wire [3-1:0] node87;
	wire [3-1:0] node88;
	wire [3-1:0] node89;
	wire [3-1:0] node93;
	wire [3-1:0] node94;
	wire [3-1:0] node98;
	wire [3-1:0] node99;
	wire [3-1:0] node103;
	wire [3-1:0] node104;
	wire [3-1:0] node105;
	wire [3-1:0] node107;
	wire [3-1:0] node110;
	wire [3-1:0] node112;
	wire [3-1:0] node115;
	wire [3-1:0] node117;
	wire [3-1:0] node118;
	wire [3-1:0] node122;
	wire [3-1:0] node123;
	wire [3-1:0] node124;
	wire [3-1:0] node125;
	wire [3-1:0] node126;
	wire [3-1:0] node127;
	wire [3-1:0] node128;
	wire [3-1:0] node131;
	wire [3-1:0] node135;
	wire [3-1:0] node136;
	wire [3-1:0] node137;
	wire [3-1:0] node140;
	wire [3-1:0] node143;
	wire [3-1:0] node145;
	wire [3-1:0] node148;
	wire [3-1:0] node149;
	wire [3-1:0] node150;
	wire [3-1:0] node151;
	wire [3-1:0] node155;
	wire [3-1:0] node156;
	wire [3-1:0] node160;
	wire [3-1:0] node161;
	wire [3-1:0] node162;
	wire [3-1:0] node166;
	wire [3-1:0] node167;
	wire [3-1:0] node171;
	wire [3-1:0] node172;
	wire [3-1:0] node173;
	wire [3-1:0] node174;
	wire [3-1:0] node176;
	wire [3-1:0] node179;
	wire [3-1:0] node180;
	wire [3-1:0] node183;
	wire [3-1:0] node186;
	wire [3-1:0] node187;
	wire [3-1:0] node188;
	wire [3-1:0] node192;
	wire [3-1:0] node194;
	wire [3-1:0] node197;
	wire [3-1:0] node198;
	wire [3-1:0] node199;
	wire [3-1:0] node201;
	wire [3-1:0] node204;
	wire [3-1:0] node205;
	wire [3-1:0] node209;
	wire [3-1:0] node211;
	wire [3-1:0] node213;
	wire [3-1:0] node216;
	wire [3-1:0] node217;
	wire [3-1:0] node218;
	wire [3-1:0] node219;
	wire [3-1:0] node221;
	wire [3-1:0] node224;
	wire [3-1:0] node227;
	wire [3-1:0] node228;
	wire [3-1:0] node229;
	wire [3-1:0] node233;
	wire [3-1:0] node234;
	wire [3-1:0] node238;
	wire [3-1:0] node239;
	wire [3-1:0] node241;
	wire [3-1:0] node242;
	wire [3-1:0] node243;
	wire [3-1:0] node248;
	wire [3-1:0] node249;
	wire [3-1:0] node250;
	wire [3-1:0] node252;
	wire [3-1:0] node255;
	wire [3-1:0] node258;
	wire [3-1:0] node260;
	wire [3-1:0] node261;
	wire [3-1:0] node265;
	wire [3-1:0] node266;
	wire [3-1:0] node267;
	wire [3-1:0] node268;
	wire [3-1:0] node269;
	wire [3-1:0] node270;
	wire [3-1:0] node273;
	wire [3-1:0] node276;
	wire [3-1:0] node277;
	wire [3-1:0] node278;
	wire [3-1:0] node280;
	wire [3-1:0] node283;
	wire [3-1:0] node286;
	wire [3-1:0] node287;
	wire [3-1:0] node289;
	wire [3-1:0] node292;
	wire [3-1:0] node293;
	wire [3-1:0] node296;
	wire [3-1:0] node299;
	wire [3-1:0] node300;
	wire [3-1:0] node301;
	wire [3-1:0] node302;
	wire [3-1:0] node304;
	wire [3-1:0] node307;
	wire [3-1:0] node308;
	wire [3-1:0] node312;
	wire [3-1:0] node313;
	wire [3-1:0] node316;
	wire [3-1:0] node319;
	wire [3-1:0] node320;
	wire [3-1:0] node321;
	wire [3-1:0] node324;
	wire [3-1:0] node325;
	wire [3-1:0] node329;
	wire [3-1:0] node330;
	wire [3-1:0] node331;
	wire [3-1:0] node335;
	wire [3-1:0] node336;
	wire [3-1:0] node339;
	wire [3-1:0] node342;
	wire [3-1:0] node343;
	wire [3-1:0] node344;
	wire [3-1:0] node345;
	wire [3-1:0] node346;
	wire [3-1:0] node349;
	wire [3-1:0] node350;
	wire [3-1:0] node354;
	wire [3-1:0] node355;
	wire [3-1:0] node356;
	wire [3-1:0] node359;
	wire [3-1:0] node362;
	wire [3-1:0] node365;
	wire [3-1:0] node367;
	wire [3-1:0] node368;
	wire [3-1:0] node371;
	wire [3-1:0] node373;
	wire [3-1:0] node376;
	wire [3-1:0] node377;
	wire [3-1:0] node378;
	wire [3-1:0] node379;
	wire [3-1:0] node380;
	wire [3-1:0] node384;
	wire [3-1:0] node385;
	wire [3-1:0] node389;
	wire [3-1:0] node390;
	wire [3-1:0] node392;
	wire [3-1:0] node396;
	wire [3-1:0] node397;
	wire [3-1:0] node399;
	wire [3-1:0] node402;
	wire [3-1:0] node403;
	wire [3-1:0] node405;
	wire [3-1:0] node409;
	wire [3-1:0] node410;
	wire [3-1:0] node411;
	wire [3-1:0] node412;
	wire [3-1:0] node413;
	wire [3-1:0] node415;
	wire [3-1:0] node416;
	wire [3-1:0] node420;
	wire [3-1:0] node421;
	wire [3-1:0] node425;
	wire [3-1:0] node426;
	wire [3-1:0] node429;
	wire [3-1:0] node430;
	wire [3-1:0] node431;
	wire [3-1:0] node435;
	wire [3-1:0] node436;
	wire [3-1:0] node439;
	wire [3-1:0] node442;
	wire [3-1:0] node443;
	wire [3-1:0] node445;
	wire [3-1:0] node446;
	wire [3-1:0] node447;
	wire [3-1:0] node452;
	wire [3-1:0] node453;
	wire [3-1:0] node454;
	wire [3-1:0] node459;
	wire [3-1:0] node460;
	wire [3-1:0] node461;
	wire [3-1:0] node462;
	wire [3-1:0] node463;
	wire [3-1:0] node467;
	wire [3-1:0] node468;
	wire [3-1:0] node469;
	wire [3-1:0] node474;
	wire [3-1:0] node475;
	wire [3-1:0] node476;
	wire [3-1:0] node477;
	wire [3-1:0] node481;
	wire [3-1:0] node482;
	wire [3-1:0] node486;
	wire [3-1:0] node487;
	wire [3-1:0] node491;
	wire [3-1:0] node492;
	wire [3-1:0] node494;
	wire [3-1:0] node497;
	wire [3-1:0] node498;
	wire [3-1:0] node500;
	wire [3-1:0] node503;
	wire [3-1:0] node506;
	wire [3-1:0] node507;
	wire [3-1:0] node509;
	wire [3-1:0] node510;
	wire [3-1:0] node511;
	wire [3-1:0] node513;
	wire [3-1:0] node515;
	wire [3-1:0] node516;
	wire [3-1:0] node522;
	wire [3-1:0] node523;
	wire [3-1:0] node524;
	wire [3-1:0] node525;
	wire [3-1:0] node527;
	wire [3-1:0] node529;
	wire [3-1:0] node531;
	wire [3-1:0] node532;
	wire [3-1:0] node535;
	wire [3-1:0] node538;
	wire [3-1:0] node540;
	wire [3-1:0] node542;
	wire [3-1:0] node545;
	wire [3-1:0] node546;
	wire [3-1:0] node547;
	wire [3-1:0] node548;
	wire [3-1:0] node549;
	wire [3-1:0] node550;
	wire [3-1:0] node555;
	wire [3-1:0] node556;
	wire [3-1:0] node557;
	wire [3-1:0] node561;
	wire [3-1:0] node562;
	wire [3-1:0] node566;
	wire [3-1:0] node568;
	wire [3-1:0] node569;
	wire [3-1:0] node571;
	wire [3-1:0] node574;
	wire [3-1:0] node575;
	wire [3-1:0] node579;
	wire [3-1:0] node580;
	wire [3-1:0] node581;
	wire [3-1:0] node582;
	wire [3-1:0] node583;
	wire [3-1:0] node586;
	wire [3-1:0] node589;
	wire [3-1:0] node591;
	wire [3-1:0] node594;
	wire [3-1:0] node595;
	wire [3-1:0] node597;
	wire [3-1:0] node601;
	wire [3-1:0] node602;
	wire [3-1:0] node603;
	wire [3-1:0] node605;
	wire [3-1:0] node608;
	wire [3-1:0] node610;
	wire [3-1:0] node613;
	wire [3-1:0] node615;
	wire [3-1:0] node616;
	wire [3-1:0] node620;
	wire [3-1:0] node621;
	wire [3-1:0] node622;
	wire [3-1:0] node624;
	wire [3-1:0] node625;
	wire [3-1:0] node626;
	wire [3-1:0] node630;
	wire [3-1:0] node631;
	wire [3-1:0] node633;
	wire [3-1:0] node638;
	wire [3-1:0] node639;
	wire [3-1:0] node640;
	wire [3-1:0] node642;
	wire [3-1:0] node645;
	wire [3-1:0] node647;
	wire [3-1:0] node650;
	wire [3-1:0] node651;
	wire [3-1:0] node652;
	wire [3-1:0] node653;
	wire [3-1:0] node658;
	wire [3-1:0] node659;
	wire [3-1:0] node660;
	wire [3-1:0] node664;
	wire [3-1:0] node665;
	wire [3-1:0] node667;
	wire [3-1:0] node670;
	wire [3-1:0] node671;

	assign outp = (inp[3]) ? node506 : node1;
		assign node1 = (inp[9]) ? node265 : node2;
			assign node2 = (inp[8]) ? node122 : node3;
				assign node3 = (inp[5]) ? node67 : node4;
					assign node4 = (inp[1]) ? node38 : node5;
						assign node5 = (inp[6]) ? node31 : node6;
							assign node6 = (inp[2]) ? node18 : node7;
								assign node7 = (inp[11]) ? node13 : node8;
									assign node8 = (inp[4]) ? node10 : 3'b001;
										assign node10 = (inp[0]) ? 3'b001 : 3'b000;
									assign node13 = (inp[7]) ? node15 : 3'b000;
										assign node15 = (inp[4]) ? 3'b001 : 3'b000;
								assign node18 = (inp[10]) ? node26 : node19;
									assign node19 = (inp[11]) ? node23 : node20;
										assign node20 = (inp[7]) ? 3'b000 : 3'b000;
										assign node23 = (inp[7]) ? 3'b001 : 3'b000;
									assign node26 = (inp[0]) ? node28 : 3'b000;
										assign node28 = (inp[4]) ? 3'b001 : 3'b000;
							assign node31 = (inp[4]) ? node33 : 3'b000;
								assign node33 = (inp[7]) ? node35 : 3'b000;
									assign node35 = (inp[0]) ? 3'b000 : 3'b001;
						assign node38 = (inp[4]) ? node54 : node39;
							assign node39 = (inp[6]) ? node47 : node40;
								assign node40 = (inp[2]) ? node42 : 3'b000;
									assign node42 = (inp[0]) ? 3'b000 : node43;
										assign node43 = (inp[7]) ? 3'b000 : 3'b001;
								assign node47 = (inp[0]) ? 3'b001 : node48;
									assign node48 = (inp[2]) ? 3'b000 : node49;
										assign node49 = (inp[7]) ? 3'b001 : 3'b000;
							assign node54 = (inp[7]) ? node56 : 3'b001;
								assign node56 = (inp[10]) ? node62 : node57;
									assign node57 = (inp[0]) ? 3'b001 : node58;
										assign node58 = (inp[6]) ? 3'b001 : 3'b000;
									assign node62 = (inp[11]) ? node64 : 3'b000;
										assign node64 = (inp[0]) ? 3'b000 : 3'b001;
					assign node67 = (inp[1]) ? node85 : node68;
						assign node68 = (inp[4]) ? node80 : node69;
							assign node69 = (inp[10]) ? node71 : 3'b001;
								assign node71 = (inp[7]) ? node75 : node72;
									assign node72 = (inp[11]) ? 3'b000 : 3'b001;
									assign node75 = (inp[0]) ? node77 : 3'b001;
										assign node77 = (inp[6]) ? 3'b000 : 3'b001;
							assign node80 = (inp[0]) ? node82 : 3'b000;
								assign node82 = (inp[6]) ? 3'b001 : 3'b000;
						assign node85 = (inp[7]) ? node103 : node86;
							assign node86 = (inp[11]) ? node98 : node87;
								assign node87 = (inp[0]) ? node93 : node88;
									assign node88 = (inp[4]) ? 3'b000 : node89;
										assign node89 = (inp[6]) ? 3'b000 : 3'b001;
									assign node93 = (inp[4]) ? 3'b001 : node94;
										assign node94 = (inp[2]) ? 3'b001 : 3'b000;
								assign node98 = (inp[6]) ? 3'b000 : node99;
									assign node99 = (inp[4]) ? 3'b000 : 3'b001;
							assign node103 = (inp[0]) ? node115 : node104;
								assign node104 = (inp[11]) ? node110 : node105;
									assign node105 = (inp[4]) ? node107 : 3'b000;
										assign node107 = (inp[10]) ? 3'b001 : 3'b000;
									assign node110 = (inp[6]) ? node112 : 3'b001;
										assign node112 = (inp[4]) ? 3'b001 : 3'b000;
								assign node115 = (inp[10]) ? node117 : 3'b000;
									assign node117 = (inp[6]) ? 3'b000 : node118;
										assign node118 = (inp[4]) ? 3'b001 : 3'b000;
				assign node122 = (inp[0]) ? node216 : node123;
					assign node123 = (inp[2]) ? node171 : node124;
						assign node124 = (inp[1]) ? node148 : node125;
							assign node125 = (inp[11]) ? node135 : node126;
								assign node126 = (inp[5]) ? 3'b000 : node127;
									assign node127 = (inp[10]) ? node131 : node128;
										assign node128 = (inp[4]) ? 3'b001 : 3'b000;
										assign node131 = (inp[4]) ? 3'b000 : 3'b001;
								assign node135 = (inp[10]) ? node143 : node136;
									assign node136 = (inp[6]) ? node140 : node137;
										assign node137 = (inp[7]) ? 3'b001 : 3'b000;
										assign node140 = (inp[5]) ? 3'b000 : 3'b000;
									assign node143 = (inp[5]) ? node145 : 3'b001;
										assign node145 = (inp[4]) ? 3'b000 : 3'b001;
							assign node148 = (inp[4]) ? node160 : node149;
								assign node149 = (inp[5]) ? node155 : node150;
									assign node150 = (inp[6]) ? 3'b000 : node151;
										assign node151 = (inp[7]) ? 3'b001 : 3'b000;
									assign node155 = (inp[11]) ? 3'b001 : node156;
										assign node156 = (inp[10]) ? 3'b000 : 3'b001;
								assign node160 = (inp[6]) ? node166 : node161;
									assign node161 = (inp[10]) ? 3'b000 : node162;
										assign node162 = (inp[11]) ? 3'b001 : 3'b000;
									assign node166 = (inp[7]) ? 3'b001 : node167;
										assign node167 = (inp[5]) ? 3'b000 : 3'b001;
						assign node171 = (inp[11]) ? node197 : node172;
							assign node172 = (inp[7]) ? node186 : node173;
								assign node173 = (inp[10]) ? node179 : node174;
									assign node174 = (inp[1]) ? node176 : 3'b001;
										assign node176 = (inp[5]) ? 3'b001 : 3'b000;
									assign node179 = (inp[4]) ? node183 : node180;
										assign node180 = (inp[1]) ? 3'b000 : 3'b001;
										assign node183 = (inp[6]) ? 3'b000 : 3'b000;
								assign node186 = (inp[10]) ? node192 : node187;
									assign node187 = (inp[6]) ? 3'b000 : node188;
										assign node188 = (inp[1]) ? 3'b001 : 3'b000;
									assign node192 = (inp[1]) ? node194 : 3'b001;
										assign node194 = (inp[5]) ? 3'b000 : 3'b001;
							assign node197 = (inp[6]) ? node209 : node198;
								assign node198 = (inp[4]) ? node204 : node199;
									assign node199 = (inp[1]) ? node201 : 3'b001;
										assign node201 = (inp[5]) ? 3'b001 : 3'b000;
									assign node204 = (inp[10]) ? 3'b000 : node205;
										assign node205 = (inp[5]) ? 3'b000 : 3'b000;
								assign node209 = (inp[7]) ? node211 : 3'b000;
									assign node211 = (inp[10]) ? node213 : 3'b000;
										assign node213 = (inp[4]) ? 3'b001 : 3'b000;
					assign node216 = (inp[5]) ? node238 : node217;
						assign node217 = (inp[1]) ? node227 : node218;
							assign node218 = (inp[4]) ? node224 : node219;
								assign node219 = (inp[6]) ? node221 : 3'b000;
									assign node221 = (inp[2]) ? 3'b000 : 3'b001;
								assign node224 = (inp[6]) ? 3'b000 : 3'b001;
							assign node227 = (inp[4]) ? node233 : node228;
								assign node228 = (inp[6]) ? 3'b001 : node229;
									assign node229 = (inp[7]) ? 3'b001 : 3'b000;
								assign node233 = (inp[6]) ? 3'b000 : node234;
									assign node234 = (inp[7]) ? 3'b001 : 3'b000;
						assign node238 = (inp[2]) ? node248 : node239;
							assign node239 = (inp[10]) ? node241 : 3'b001;
								assign node241 = (inp[1]) ? 3'b001 : node242;
									assign node242 = (inp[11]) ? 3'b001 : node243;
										assign node243 = (inp[4]) ? 3'b001 : 3'b000;
							assign node248 = (inp[6]) ? node258 : node249;
								assign node249 = (inp[4]) ? node255 : node250;
									assign node250 = (inp[1]) ? node252 : 3'b001;
										assign node252 = (inp[10]) ? 3'b000 : 3'b001;
									assign node255 = (inp[1]) ? 3'b001 : 3'b000;
								assign node258 = (inp[7]) ? node260 : 3'b001;
									assign node260 = (inp[11]) ? 3'b001 : node261;
										assign node261 = (inp[1]) ? 3'b000 : 3'b000;
			assign node265 = (inp[4]) ? node409 : node266;
				assign node266 = (inp[6]) ? node342 : node267;
					assign node267 = (inp[0]) ? node299 : node268;
						assign node268 = (inp[1]) ? node276 : node269;
							assign node269 = (inp[7]) ? node273 : node270;
								assign node270 = (inp[5]) ? 3'b100 : 3'b010;
								assign node273 = (inp[5]) ? 3'b010 : 3'b110;
							assign node276 = (inp[5]) ? node286 : node277;
								assign node277 = (inp[7]) ? node283 : node278;
									assign node278 = (inp[2]) ? node280 : 3'b101;
										assign node280 = (inp[8]) ? 3'b110 : 3'b110;
									assign node283 = (inp[8]) ? 3'b001 : 3'b101;
								assign node286 = (inp[8]) ? node292 : node287;
									assign node287 = (inp[2]) ? node289 : 3'b010;
										assign node289 = (inp[7]) ? 3'b110 : 3'b010;
									assign node292 = (inp[7]) ? node296 : node293;
										assign node293 = (inp[11]) ? 3'b010 : 3'b001;
										assign node296 = (inp[10]) ? 3'b101 : 3'b110;
						assign node299 = (inp[5]) ? node319 : node300;
							assign node300 = (inp[7]) ? node312 : node301;
								assign node301 = (inp[2]) ? node307 : node302;
									assign node302 = (inp[1]) ? node304 : 3'b110;
										assign node304 = (inp[11]) ? 3'b000 : 3'b101;
									assign node307 = (inp[11]) ? 3'b001 : node308;
										assign node308 = (inp[1]) ? 3'b100 : 3'b001;
								assign node312 = (inp[8]) ? node316 : node313;
									assign node313 = (inp[1]) ? 3'b101 : 3'b001;
									assign node316 = (inp[1]) ? 3'b011 : 3'b001;
							assign node319 = (inp[1]) ? node329 : node320;
								assign node320 = (inp[11]) ? node324 : node321;
									assign node321 = (inp[8]) ? 3'b010 : 3'b110;
									assign node324 = (inp[2]) ? 3'b110 : node325;
										assign node325 = (inp[8]) ? 3'b110 : 3'b010;
								assign node329 = (inp[7]) ? node335 : node330;
									assign node330 = (inp[8]) ? 3'b111 : node331;
										assign node331 = (inp[11]) ? 3'b110 : 3'b111;
									assign node335 = (inp[11]) ? node339 : node336;
										assign node336 = (inp[2]) ? 3'b111 : 3'b101;
										assign node339 = (inp[8]) ? 3'b101 : 3'b001;
					assign node342 = (inp[1]) ? node376 : node343;
						assign node343 = (inp[0]) ? node365 : node344;
							assign node344 = (inp[5]) ? node354 : node345;
								assign node345 = (inp[2]) ? node349 : node346;
									assign node346 = (inp[10]) ? 3'b001 : 3'b101;
									assign node349 = (inp[8]) ? 3'b101 : node350;
										assign node350 = (inp[7]) ? 3'b001 : 3'b101;
								assign node354 = (inp[8]) ? node362 : node355;
									assign node355 = (inp[7]) ? node359 : node356;
										assign node356 = (inp[10]) ? 3'b010 : 3'b110;
										assign node359 = (inp[2]) ? 3'b010 : 3'b110;
									assign node362 = (inp[7]) ? 3'b001 : 3'b110;
							assign node365 = (inp[7]) ? node367 : 3'b101;
								assign node367 = (inp[10]) ? node371 : node368;
									assign node368 = (inp[8]) ? 3'b101 : 3'b001;
									assign node371 = (inp[5]) ? node373 : 3'b011;
										assign node373 = (inp[2]) ? 3'b011 : 3'b101;
						assign node376 = (inp[5]) ? node396 : node377;
							assign node377 = (inp[0]) ? node389 : node378;
								assign node378 = (inp[11]) ? node384 : node379;
									assign node379 = (inp[2]) ? 3'b011 : node380;
										assign node380 = (inp[10]) ? 3'b001 : 3'b001;
									assign node384 = (inp[2]) ? 3'b101 : node385;
										assign node385 = (inp[10]) ? 3'b011 : 3'b001;
								assign node389 = (inp[7]) ? 3'b111 : node390;
									assign node390 = (inp[10]) ? node392 : 3'b011;
										assign node392 = (inp[2]) ? 3'b111 : 3'b011;
							assign node396 = (inp[8]) ? node402 : node397;
								assign node397 = (inp[2]) ? node399 : 3'b001;
									assign node399 = (inp[11]) ? 3'b101 : 3'b001;
								assign node402 = (inp[0]) ? 3'b011 : node403;
									assign node403 = (inp[7]) ? node405 : 3'b001;
										assign node405 = (inp[10]) ? 3'b101 : 3'b001;
				assign node409 = (inp[6]) ? node459 : node410;
					assign node410 = (inp[0]) ? node442 : node411;
						assign node411 = (inp[1]) ? node425 : node412;
							assign node412 = (inp[5]) ? node420 : node413;
								assign node413 = (inp[10]) ? node415 : 3'b100;
									assign node415 = (inp[2]) ? 3'b100 : node416;
										assign node416 = (inp[8]) ? 3'b000 : 3'b100;
								assign node420 = (inp[8]) ? 3'b000 : node421;
									assign node421 = (inp[7]) ? 3'b000 : 3'b100;
							assign node425 = (inp[7]) ? node429 : node426;
								assign node426 = (inp[5]) ? 3'b000 : 3'b100;
								assign node429 = (inp[5]) ? node435 : node430;
									assign node430 = (inp[8]) ? 3'b010 : node431;
										assign node431 = (inp[10]) ? 3'b000 : 3'b010;
									assign node435 = (inp[2]) ? node439 : node436;
										assign node436 = (inp[11]) ? 3'b010 : 3'b110;
										assign node439 = (inp[10]) ? 3'b100 : 3'b110;
						assign node442 = (inp[1]) ? node452 : node443;
							assign node443 = (inp[5]) ? node445 : 3'b010;
								assign node445 = (inp[7]) ? 3'b100 : node446;
									assign node446 = (inp[2]) ? 3'b100 : node447;
										assign node447 = (inp[8]) ? 3'b110 : 3'b000;
							assign node452 = (inp[5]) ? 3'b010 : node453;
								assign node453 = (inp[7]) ? 3'b110 : node454;
									assign node454 = (inp[8]) ? 3'b100 : 3'b010;
					assign node459 = (inp[0]) ? node491 : node460;
						assign node460 = (inp[7]) ? node474 : node461;
							assign node461 = (inp[5]) ? node467 : node462;
								assign node462 = (inp[1]) ? 3'b110 : node463;
									assign node463 = (inp[8]) ? 3'b010 : 3'b100;
								assign node467 = (inp[1]) ? 3'b100 : node468;
									assign node468 = (inp[11]) ? 3'b100 : node469;
										assign node469 = (inp[8]) ? 3'b010 : 3'b100;
							assign node474 = (inp[5]) ? node486 : node475;
								assign node475 = (inp[2]) ? node481 : node476;
									assign node476 = (inp[1]) ? 3'b110 : node477;
										assign node477 = (inp[10]) ? 3'b010 : 3'b000;
									assign node481 = (inp[8]) ? 3'b001 : node482;
										assign node482 = (inp[11]) ? 3'b010 : 3'b110;
								assign node486 = (inp[10]) ? 3'b010 : node487;
									assign node487 = (inp[1]) ? 3'b010 : 3'b000;
						assign node491 = (inp[5]) ? node497 : node492;
							assign node492 = (inp[7]) ? node494 : 3'b001;
								assign node494 = (inp[1]) ? 3'b101 : 3'b001;
							assign node497 = (inp[1]) ? node503 : node498;
								assign node498 = (inp[7]) ? node500 : 3'b010;
									assign node500 = (inp[10]) ? 3'b110 : 3'b010;
								assign node503 = (inp[7]) ? 3'b001 : 3'b110;
		assign node506 = (inp[6]) ? node522 : node507;
			assign node507 = (inp[1]) ? node509 : 3'b000;
				assign node509 = (inp[4]) ? 3'b000 : node510;
					assign node510 = (inp[5]) ? 3'b000 : node511;
						assign node511 = (inp[0]) ? node513 : 3'b000;
							assign node513 = (inp[9]) ? node515 : 3'b000;
								assign node515 = (inp[7]) ? 3'b100 : node516;
									assign node516 = (inp[8]) ? 3'b100 : 3'b000;
			assign node522 = (inp[9]) ? node620 : node523;
				assign node523 = (inp[4]) ? node545 : node524;
					assign node524 = (inp[0]) ? node538 : node525;
						assign node525 = (inp[1]) ? node527 : 3'b010;
							assign node527 = (inp[2]) ? node529 : 3'b010;
								assign node529 = (inp[7]) ? node531 : 3'b010;
									assign node531 = (inp[5]) ? node535 : node532;
										assign node532 = (inp[11]) ? 3'b010 : 3'b011;
										assign node535 = (inp[8]) ? 3'b010 : 3'b011;
						assign node538 = (inp[5]) ? node540 : 3'b011;
							assign node540 = (inp[1]) ? node542 : 3'b010;
								assign node542 = (inp[7]) ? 3'b011 : 3'b010;
					assign node545 = (inp[0]) ? node579 : node546;
						assign node546 = (inp[10]) ? node566 : node547;
							assign node547 = (inp[8]) ? node555 : node548;
								assign node548 = (inp[1]) ? 3'b000 : node549;
									assign node549 = (inp[11]) ? 3'b100 : node550;
										assign node550 = (inp[2]) ? 3'b100 : 3'b110;
								assign node555 = (inp[2]) ? node561 : node556;
									assign node556 = (inp[1]) ? 3'b000 : node557;
										assign node557 = (inp[5]) ? 3'b000 : 3'b010;
									assign node561 = (inp[5]) ? 3'b010 : node562;
										assign node562 = (inp[1]) ? 3'b100 : 3'b010;
							assign node566 = (inp[1]) ? node568 : 3'b000;
								assign node568 = (inp[5]) ? node574 : node569;
									assign node569 = (inp[11]) ? node571 : 3'b000;
										assign node571 = (inp[8]) ? 3'b000 : 3'b100;
									assign node574 = (inp[11]) ? 3'b100 : node575;
										assign node575 = (inp[7]) ? 3'b100 : 3'b000;
						assign node579 = (inp[7]) ? node601 : node580;
							assign node580 = (inp[10]) ? node594 : node581;
								assign node581 = (inp[1]) ? node589 : node582;
									assign node582 = (inp[8]) ? node586 : node583;
										assign node583 = (inp[2]) ? 3'b100 : 3'b000;
										assign node586 = (inp[11]) ? 3'b100 : 3'b010;
									assign node589 = (inp[5]) ? node591 : 3'b110;
										assign node591 = (inp[11]) ? 3'b010 : 3'b110;
								assign node594 = (inp[5]) ? 3'b100 : node595;
									assign node595 = (inp[1]) ? node597 : 3'b100;
										assign node597 = (inp[8]) ? 3'b010 : 3'b100;
							assign node601 = (inp[5]) ? node613 : node602;
								assign node602 = (inp[2]) ? node608 : node603;
									assign node603 = (inp[1]) ? node605 : 3'b010;
										assign node605 = (inp[8]) ? 3'b001 : 3'b101;
									assign node608 = (inp[8]) ? node610 : 3'b010;
										assign node610 = (inp[11]) ? 3'b110 : 3'b010;
								assign node613 = (inp[11]) ? node615 : 3'b110;
									assign node615 = (inp[1]) ? 3'b010 : node616;
										assign node616 = (inp[10]) ? 3'b100 : 3'b010;
				assign node620 = (inp[0]) ? node638 : node621;
					assign node621 = (inp[4]) ? 3'b000 : node622;
						assign node622 = (inp[10]) ? node624 : 3'b000;
							assign node624 = (inp[2]) ? node630 : node625;
								assign node625 = (inp[5]) ? 3'b000 : node626;
									assign node626 = (inp[7]) ? 3'b100 : 3'b000;
								assign node630 = (inp[1]) ? 3'b100 : node631;
									assign node631 = (inp[8]) ? node633 : 3'b000;
										assign node633 = (inp[11]) ? 3'b000 : 3'b100;
					assign node638 = (inp[4]) ? node650 : node639;
						assign node639 = (inp[5]) ? node645 : node640;
							assign node640 = (inp[7]) ? node642 : 3'b010;
								assign node642 = (inp[1]) ? 3'b110 : 3'b010;
							assign node645 = (inp[1]) ? node647 : 3'b100;
								assign node647 = (inp[7]) ? 3'b010 : 3'b100;
						assign node650 = (inp[7]) ? node658 : node651;
							assign node651 = (inp[5]) ? 3'b000 : node652;
								assign node652 = (inp[10]) ? 3'b000 : node653;
									assign node653 = (inp[1]) ? 3'b100 : 3'b000;
							assign node658 = (inp[1]) ? node664 : node659;
								assign node659 = (inp[5]) ? 3'b000 : node660;
									assign node660 = (inp[8]) ? 3'b100 : 3'b000;
								assign node664 = (inp[10]) ? node670 : node665;
									assign node665 = (inp[11]) ? node667 : 3'b010;
										assign node667 = (inp[5]) ? 3'b100 : 3'b010;
									assign node670 = (inp[8]) ? 3'b100 : node671;
										assign node671 = (inp[5]) ? 3'b000 : 3'b100;

endmodule