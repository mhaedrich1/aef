module dtc_split33_bm62 (
	input  wire [16-1:0] inp,
	output wire [4-1:0] outp
);

	wire [4-1:0] node1;
	wire [4-1:0] node2;
	wire [4-1:0] node3;
	wire [4-1:0] node4;
	wire [4-1:0] node5;
	wire [4-1:0] node6;
	wire [4-1:0] node7;
	wire [4-1:0] node8;
	wire [4-1:0] node9;
	wire [4-1:0] node10;
	wire [4-1:0] node11;
	wire [4-1:0] node12;
	wire [4-1:0] node15;
	wire [4-1:0] node16;
	wire [4-1:0] node20;
	wire [4-1:0] node21;
	wire [4-1:0] node22;
	wire [4-1:0] node27;
	wire [4-1:0] node28;
	wire [4-1:0] node29;
	wire [4-1:0] node31;
	wire [4-1:0] node34;
	wire [4-1:0] node36;
	wire [4-1:0] node39;
	wire [4-1:0] node42;
	wire [4-1:0] node43;
	wire [4-1:0] node44;
	wire [4-1:0] node46;
	wire [4-1:0] node48;
	wire [4-1:0] node51;
	wire [4-1:0] node53;
	wire [4-1:0] node54;
	wire [4-1:0] node57;
	wire [4-1:0] node60;
	wire [4-1:0] node61;
	wire [4-1:0] node62;
	wire [4-1:0] node63;
	wire [4-1:0] node66;
	wire [4-1:0] node70;
	wire [4-1:0] node71;
	wire [4-1:0] node73;
	wire [4-1:0] node76;
	wire [4-1:0] node77;
	wire [4-1:0] node81;
	wire [4-1:0] node82;
	wire [4-1:0] node83;
	wire [4-1:0] node84;
	wire [4-1:0] node85;
	wire [4-1:0] node86;
	wire [4-1:0] node89;
	wire [4-1:0] node92;
	wire [4-1:0] node94;
	wire [4-1:0] node97;
	wire [4-1:0] node98;
	wire [4-1:0] node99;
	wire [4-1:0] node102;
	wire [4-1:0] node106;
	wire [4-1:0] node107;
	wire [4-1:0] node108;
	wire [4-1:0] node109;
	wire [4-1:0] node112;
	wire [4-1:0] node115;
	wire [4-1:0] node116;
	wire [4-1:0] node120;
	wire [4-1:0] node121;
	wire [4-1:0] node122;
	wire [4-1:0] node126;
	wire [4-1:0] node128;
	wire [4-1:0] node131;
	wire [4-1:0] node132;
	wire [4-1:0] node133;
	wire [4-1:0] node134;
	wire [4-1:0] node137;
	wire [4-1:0] node140;
	wire [4-1:0] node141;
	wire [4-1:0] node142;
	wire [4-1:0] node145;
	wire [4-1:0] node148;
	wire [4-1:0] node149;
	wire [4-1:0] node153;
	wire [4-1:0] node154;
	wire [4-1:0] node155;
	wire [4-1:0] node157;
	wire [4-1:0] node160;
	wire [4-1:0] node163;
	wire [4-1:0] node164;
	wire [4-1:0] node165;
	wire [4-1:0] node168;
	wire [4-1:0] node171;
	wire [4-1:0] node172;
	wire [4-1:0] node175;
	wire [4-1:0] node178;
	wire [4-1:0] node179;
	wire [4-1:0] node180;
	wire [4-1:0] node181;
	wire [4-1:0] node182;
	wire [4-1:0] node183;
	wire [4-1:0] node185;
	wire [4-1:0] node188;
	wire [4-1:0] node189;
	wire [4-1:0] node193;
	wire [4-1:0] node194;
	wire [4-1:0] node195;
	wire [4-1:0] node198;
	wire [4-1:0] node201;
	wire [4-1:0] node203;
	wire [4-1:0] node206;
	wire [4-1:0] node207;
	wire [4-1:0] node208;
	wire [4-1:0] node209;
	wire [4-1:0] node212;
	wire [4-1:0] node215;
	wire [4-1:0] node217;
	wire [4-1:0] node220;
	wire [4-1:0] node221;
	wire [4-1:0] node222;
	wire [4-1:0] node225;
	wire [4-1:0] node228;
	wire [4-1:0] node230;
	wire [4-1:0] node233;
	wire [4-1:0] node234;
	wire [4-1:0] node235;
	wire [4-1:0] node236;
	wire [4-1:0] node237;
	wire [4-1:0] node242;
	wire [4-1:0] node243;
	wire [4-1:0] node245;
	wire [4-1:0] node248;
	wire [4-1:0] node249;
	wire [4-1:0] node253;
	wire [4-1:0] node254;
	wire [4-1:0] node255;
	wire [4-1:0] node258;
	wire [4-1:0] node259;
	wire [4-1:0] node263;
	wire [4-1:0] node265;
	wire [4-1:0] node266;
	wire [4-1:0] node270;
	wire [4-1:0] node271;
	wire [4-1:0] node272;
	wire [4-1:0] node273;
	wire [4-1:0] node274;
	wire [4-1:0] node276;
	wire [4-1:0] node279;
	wire [4-1:0] node280;
	wire [4-1:0] node283;
	wire [4-1:0] node286;
	wire [4-1:0] node287;
	wire [4-1:0] node290;
	wire [4-1:0] node291;
	wire [4-1:0] node294;
	wire [4-1:0] node297;
	wire [4-1:0] node298;
	wire [4-1:0] node299;
	wire [4-1:0] node301;
	wire [4-1:0] node304;
	wire [4-1:0] node306;
	wire [4-1:0] node309;
	wire [4-1:0] node310;
	wire [4-1:0] node311;
	wire [4-1:0] node314;
	wire [4-1:0] node317;
	wire [4-1:0] node318;
	wire [4-1:0] node322;
	wire [4-1:0] node323;
	wire [4-1:0] node324;
	wire [4-1:0] node325;
	wire [4-1:0] node328;
	wire [4-1:0] node329;
	wire [4-1:0] node332;
	wire [4-1:0] node335;
	wire [4-1:0] node336;
	wire [4-1:0] node339;
	wire [4-1:0] node342;
	wire [4-1:0] node343;
	wire [4-1:0] node345;
	wire [4-1:0] node347;
	wire [4-1:0] node350;
	wire [4-1:0] node351;
	wire [4-1:0] node352;
	wire [4-1:0] node357;
	wire [4-1:0] node358;
	wire [4-1:0] node359;
	wire [4-1:0] node360;
	wire [4-1:0] node361;
	wire [4-1:0] node362;
	wire [4-1:0] node363;
	wire [4-1:0] node366;
	wire [4-1:0] node368;
	wire [4-1:0] node371;
	wire [4-1:0] node372;
	wire [4-1:0] node375;
	wire [4-1:0] node378;
	wire [4-1:0] node379;
	wire [4-1:0] node380;
	wire [4-1:0] node382;
	wire [4-1:0] node385;
	wire [4-1:0] node387;
	wire [4-1:0] node390;
	wire [4-1:0] node391;
	wire [4-1:0] node394;
	wire [4-1:0] node397;
	wire [4-1:0] node398;
	wire [4-1:0] node399;
	wire [4-1:0] node400;
	wire [4-1:0] node401;
	wire [4-1:0] node405;
	wire [4-1:0] node406;
	wire [4-1:0] node410;
	wire [4-1:0] node411;
	wire [4-1:0] node412;
	wire [4-1:0] node415;
	wire [4-1:0] node418;
	wire [4-1:0] node419;
	wire [4-1:0] node423;
	wire [4-1:0] node424;
	wire [4-1:0] node425;
	wire [4-1:0] node426;
	wire [4-1:0] node429;
	wire [4-1:0] node433;
	wire [4-1:0] node434;
	wire [4-1:0] node435;
	wire [4-1:0] node439;
	wire [4-1:0] node440;
	wire [4-1:0] node444;
	wire [4-1:0] node445;
	wire [4-1:0] node446;
	wire [4-1:0] node447;
	wire [4-1:0] node448;
	wire [4-1:0] node450;
	wire [4-1:0] node454;
	wire [4-1:0] node455;
	wire [4-1:0] node456;
	wire [4-1:0] node459;
	wire [4-1:0] node463;
	wire [4-1:0] node464;
	wire [4-1:0] node465;
	wire [4-1:0] node466;
	wire [4-1:0] node471;
	wire [4-1:0] node473;
	wire [4-1:0] node476;
	wire [4-1:0] node477;
	wire [4-1:0] node478;
	wire [4-1:0] node479;
	wire [4-1:0] node481;
	wire [4-1:0] node484;
	wire [4-1:0] node485;
	wire [4-1:0] node489;
	wire [4-1:0] node490;
	wire [4-1:0] node494;
	wire [4-1:0] node495;
	wire [4-1:0] node498;
	wire [4-1:0] node499;
	wire [4-1:0] node500;
	wire [4-1:0] node504;
	wire [4-1:0] node507;
	wire [4-1:0] node508;
	wire [4-1:0] node509;
	wire [4-1:0] node510;
	wire [4-1:0] node511;
	wire [4-1:0] node512;
	wire [4-1:0] node513;
	wire [4-1:0] node517;
	wire [4-1:0] node519;
	wire [4-1:0] node522;
	wire [4-1:0] node523;
	wire [4-1:0] node524;
	wire [4-1:0] node527;
	wire [4-1:0] node530;
	wire [4-1:0] node533;
	wire [4-1:0] node534;
	wire [4-1:0] node535;
	wire [4-1:0] node536;
	wire [4-1:0] node540;
	wire [4-1:0] node541;
	wire [4-1:0] node545;
	wire [4-1:0] node547;
	wire [4-1:0] node550;
	wire [4-1:0] node551;
	wire [4-1:0] node552;
	wire [4-1:0] node553;
	wire [4-1:0] node554;
	wire [4-1:0] node557;
	wire [4-1:0] node561;
	wire [4-1:0] node564;
	wire [4-1:0] node565;
	wire [4-1:0] node566;
	wire [4-1:0] node567;
	wire [4-1:0] node571;
	wire [4-1:0] node574;
	wire [4-1:0] node575;
	wire [4-1:0] node578;
	wire [4-1:0] node580;
	wire [4-1:0] node583;
	wire [4-1:0] node584;
	wire [4-1:0] node585;
	wire [4-1:0] node586;
	wire [4-1:0] node587;
	wire [4-1:0] node590;
	wire [4-1:0] node591;
	wire [4-1:0] node594;
	wire [4-1:0] node597;
	wire [4-1:0] node598;
	wire [4-1:0] node599;
	wire [4-1:0] node602;
	wire [4-1:0] node605;
	wire [4-1:0] node606;
	wire [4-1:0] node609;
	wire [4-1:0] node612;
	wire [4-1:0] node613;
	wire [4-1:0] node614;
	wire [4-1:0] node615;
	wire [4-1:0] node618;
	wire [4-1:0] node621;
	wire [4-1:0] node622;
	wire [4-1:0] node626;
	wire [4-1:0] node627;
	wire [4-1:0] node628;
	wire [4-1:0] node632;
	wire [4-1:0] node633;
	wire [4-1:0] node636;
	wire [4-1:0] node639;
	wire [4-1:0] node640;
	wire [4-1:0] node641;
	wire [4-1:0] node642;
	wire [4-1:0] node644;
	wire [4-1:0] node648;
	wire [4-1:0] node649;
	wire [4-1:0] node651;
	wire [4-1:0] node654;
	wire [4-1:0] node655;
	wire [4-1:0] node659;
	wire [4-1:0] node660;
	wire [4-1:0] node661;
	wire [4-1:0] node662;
	wire [4-1:0] node665;
	wire [4-1:0] node668;
	wire [4-1:0] node671;
	wire [4-1:0] node672;
	wire [4-1:0] node673;
	wire [4-1:0] node676;
	wire [4-1:0] node679;
	wire [4-1:0] node680;
	wire [4-1:0] node683;
	wire [4-1:0] node686;
	wire [4-1:0] node687;
	wire [4-1:0] node688;
	wire [4-1:0] node689;
	wire [4-1:0] node690;
	wire [4-1:0] node691;
	wire [4-1:0] node692;
	wire [4-1:0] node693;
	wire [4-1:0] node694;
	wire [4-1:0] node698;
	wire [4-1:0] node701;
	wire [4-1:0] node702;
	wire [4-1:0] node703;
	wire [4-1:0] node707;
	wire [4-1:0] node710;
	wire [4-1:0] node711;
	wire [4-1:0] node712;
	wire [4-1:0] node714;
	wire [4-1:0] node718;
	wire [4-1:0] node719;
	wire [4-1:0] node722;
	wire [4-1:0] node723;
	wire [4-1:0] node727;
	wire [4-1:0] node728;
	wire [4-1:0] node729;
	wire [4-1:0] node730;
	wire [4-1:0] node731;
	wire [4-1:0] node734;
	wire [4-1:0] node737;
	wire [4-1:0] node739;
	wire [4-1:0] node742;
	wire [4-1:0] node743;
	wire [4-1:0] node744;
	wire [4-1:0] node748;
	wire [4-1:0] node751;
	wire [4-1:0] node752;
	wire [4-1:0] node753;
	wire [4-1:0] node754;
	wire [4-1:0] node758;
	wire [4-1:0] node761;
	wire [4-1:0] node762;
	wire [4-1:0] node763;
	wire [4-1:0] node767;
	wire [4-1:0] node770;
	wire [4-1:0] node771;
	wire [4-1:0] node772;
	wire [4-1:0] node773;
	wire [4-1:0] node774;
	wire [4-1:0] node777;
	wire [4-1:0] node779;
	wire [4-1:0] node782;
	wire [4-1:0] node785;
	wire [4-1:0] node786;
	wire [4-1:0] node787;
	wire [4-1:0] node788;
	wire [4-1:0] node792;
	wire [4-1:0] node793;
	wire [4-1:0] node797;
	wire [4-1:0] node798;
	wire [4-1:0] node799;
	wire [4-1:0] node802;
	wire [4-1:0] node805;
	wire [4-1:0] node806;
	wire [4-1:0] node809;
	wire [4-1:0] node812;
	wire [4-1:0] node813;
	wire [4-1:0] node814;
	wire [4-1:0] node815;
	wire [4-1:0] node816;
	wire [4-1:0] node819;
	wire [4-1:0] node822;
	wire [4-1:0] node824;
	wire [4-1:0] node827;
	wire [4-1:0] node828;
	wire [4-1:0] node829;
	wire [4-1:0] node833;
	wire [4-1:0] node835;
	wire [4-1:0] node838;
	wire [4-1:0] node839;
	wire [4-1:0] node840;
	wire [4-1:0] node841;
	wire [4-1:0] node844;
	wire [4-1:0] node847;
	wire [4-1:0] node850;
	wire [4-1:0] node851;
	wire [4-1:0] node853;
	wire [4-1:0] node856;
	wire [4-1:0] node858;
	wire [4-1:0] node861;
	wire [4-1:0] node862;
	wire [4-1:0] node863;
	wire [4-1:0] node864;
	wire [4-1:0] node865;
	wire [4-1:0] node867;
	wire [4-1:0] node869;
	wire [4-1:0] node872;
	wire [4-1:0] node873;
	wire [4-1:0] node875;
	wire [4-1:0] node878;
	wire [4-1:0] node880;
	wire [4-1:0] node883;
	wire [4-1:0] node884;
	wire [4-1:0] node885;
	wire [4-1:0] node886;
	wire [4-1:0] node889;
	wire [4-1:0] node892;
	wire [4-1:0] node894;
	wire [4-1:0] node897;
	wire [4-1:0] node898;
	wire [4-1:0] node899;
	wire [4-1:0] node903;
	wire [4-1:0] node906;
	wire [4-1:0] node907;
	wire [4-1:0] node908;
	wire [4-1:0] node909;
	wire [4-1:0] node910;
	wire [4-1:0] node913;
	wire [4-1:0] node916;
	wire [4-1:0] node918;
	wire [4-1:0] node921;
	wire [4-1:0] node922;
	wire [4-1:0] node923;
	wire [4-1:0] node927;
	wire [4-1:0] node928;
	wire [4-1:0] node931;
	wire [4-1:0] node934;
	wire [4-1:0] node935;
	wire [4-1:0] node936;
	wire [4-1:0] node937;
	wire [4-1:0] node942;
	wire [4-1:0] node944;
	wire [4-1:0] node945;
	wire [4-1:0] node949;
	wire [4-1:0] node950;
	wire [4-1:0] node951;
	wire [4-1:0] node952;
	wire [4-1:0] node953;
	wire [4-1:0] node954;
	wire [4-1:0] node958;
	wire [4-1:0] node961;
	wire [4-1:0] node963;
	wire [4-1:0] node964;
	wire [4-1:0] node968;
	wire [4-1:0] node969;
	wire [4-1:0] node970;
	wire [4-1:0] node971;
	wire [4-1:0] node975;
	wire [4-1:0] node978;
	wire [4-1:0] node980;
	wire [4-1:0] node983;
	wire [4-1:0] node984;
	wire [4-1:0] node985;
	wire [4-1:0] node986;
	wire [4-1:0] node988;
	wire [4-1:0] node991;
	wire [4-1:0] node993;
	wire [4-1:0] node996;
	wire [4-1:0] node998;
	wire [4-1:0] node999;
	wire [4-1:0] node1003;
	wire [4-1:0] node1004;
	wire [4-1:0] node1005;
	wire [4-1:0] node1007;
	wire [4-1:0] node1010;
	wire [4-1:0] node1012;
	wire [4-1:0] node1015;
	wire [4-1:0] node1016;
	wire [4-1:0] node1017;
	wire [4-1:0] node1022;
	wire [4-1:0] node1023;
	wire [4-1:0] node1024;
	wire [4-1:0] node1025;
	wire [4-1:0] node1026;
	wire [4-1:0] node1027;
	wire [4-1:0] node1028;
	wire [4-1:0] node1030;
	wire [4-1:0] node1033;
	wire [4-1:0] node1035;
	wire [4-1:0] node1038;
	wire [4-1:0] node1039;
	wire [4-1:0] node1041;
	wire [4-1:0] node1044;
	wire [4-1:0] node1045;
	wire [4-1:0] node1048;
	wire [4-1:0] node1051;
	wire [4-1:0] node1052;
	wire [4-1:0] node1053;
	wire [4-1:0] node1054;
	wire [4-1:0] node1058;
	wire [4-1:0] node1060;
	wire [4-1:0] node1063;
	wire [4-1:0] node1064;
	wire [4-1:0] node1065;
	wire [4-1:0] node1069;
	wire [4-1:0] node1070;
	wire [4-1:0] node1074;
	wire [4-1:0] node1075;
	wire [4-1:0] node1076;
	wire [4-1:0] node1077;
	wire [4-1:0] node1078;
	wire [4-1:0] node1081;
	wire [4-1:0] node1084;
	wire [4-1:0] node1085;
	wire [4-1:0] node1089;
	wire [4-1:0] node1090;
	wire [4-1:0] node1091;
	wire [4-1:0] node1096;
	wire [4-1:0] node1097;
	wire [4-1:0] node1098;
	wire [4-1:0] node1100;
	wire [4-1:0] node1103;
	wire [4-1:0] node1106;
	wire [4-1:0] node1107;
	wire [4-1:0] node1108;
	wire [4-1:0] node1111;
	wire [4-1:0] node1114;
	wire [4-1:0] node1116;
	wire [4-1:0] node1119;
	wire [4-1:0] node1120;
	wire [4-1:0] node1121;
	wire [4-1:0] node1122;
	wire [4-1:0] node1123;
	wire [4-1:0] node1125;
	wire [4-1:0] node1128;
	wire [4-1:0] node1129;
	wire [4-1:0] node1133;
	wire [4-1:0] node1134;
	wire [4-1:0] node1136;
	wire [4-1:0] node1139;
	wire [4-1:0] node1141;
	wire [4-1:0] node1144;
	wire [4-1:0] node1145;
	wire [4-1:0] node1146;
	wire [4-1:0] node1148;
	wire [4-1:0] node1151;
	wire [4-1:0] node1153;
	wire [4-1:0] node1156;
	wire [4-1:0] node1157;
	wire [4-1:0] node1158;
	wire [4-1:0] node1161;
	wire [4-1:0] node1164;
	wire [4-1:0] node1166;
	wire [4-1:0] node1169;
	wire [4-1:0] node1170;
	wire [4-1:0] node1171;
	wire [4-1:0] node1172;
	wire [4-1:0] node1174;
	wire [4-1:0] node1177;
	wire [4-1:0] node1178;
	wire [4-1:0] node1182;
	wire [4-1:0] node1183;
	wire [4-1:0] node1186;
	wire [4-1:0] node1188;
	wire [4-1:0] node1191;
	wire [4-1:0] node1192;
	wire [4-1:0] node1193;
	wire [4-1:0] node1194;
	wire [4-1:0] node1198;
	wire [4-1:0] node1201;
	wire [4-1:0] node1202;
	wire [4-1:0] node1204;
	wire [4-1:0] node1207;
	wire [4-1:0] node1208;
	wire [4-1:0] node1211;
	wire [4-1:0] node1214;
	wire [4-1:0] node1215;
	wire [4-1:0] node1216;
	wire [4-1:0] node1217;
	wire [4-1:0] node1218;
	wire [4-1:0] node1219;
	wire [4-1:0] node1222;
	wire [4-1:0] node1224;
	wire [4-1:0] node1227;
	wire [4-1:0] node1228;
	wire [4-1:0] node1229;
	wire [4-1:0] node1233;
	wire [4-1:0] node1234;
	wire [4-1:0] node1237;
	wire [4-1:0] node1240;
	wire [4-1:0] node1241;
	wire [4-1:0] node1242;
	wire [4-1:0] node1244;
	wire [4-1:0] node1247;
	wire [4-1:0] node1248;
	wire [4-1:0] node1252;
	wire [4-1:0] node1254;
	wire [4-1:0] node1257;
	wire [4-1:0] node1258;
	wire [4-1:0] node1259;
	wire [4-1:0] node1260;
	wire [4-1:0] node1261;
	wire [4-1:0] node1264;
	wire [4-1:0] node1267;
	wire [4-1:0] node1268;
	wire [4-1:0] node1272;
	wire [4-1:0] node1273;
	wire [4-1:0] node1275;
	wire [4-1:0] node1278;
	wire [4-1:0] node1280;
	wire [4-1:0] node1283;
	wire [4-1:0] node1284;
	wire [4-1:0] node1285;
	wire [4-1:0] node1286;
	wire [4-1:0] node1289;
	wire [4-1:0] node1292;
	wire [4-1:0] node1294;
	wire [4-1:0] node1297;
	wire [4-1:0] node1298;
	wire [4-1:0] node1299;
	wire [4-1:0] node1302;
	wire [4-1:0] node1306;
	wire [4-1:0] node1307;
	wire [4-1:0] node1308;
	wire [4-1:0] node1309;
	wire [4-1:0] node1310;
	wire [4-1:0] node1313;
	wire [4-1:0] node1314;
	wire [4-1:0] node1317;
	wire [4-1:0] node1320;
	wire [4-1:0] node1321;
	wire [4-1:0] node1323;
	wire [4-1:0] node1326;
	wire [4-1:0] node1327;
	wire [4-1:0] node1330;
	wire [4-1:0] node1333;
	wire [4-1:0] node1335;
	wire [4-1:0] node1336;
	wire [4-1:0] node1337;
	wire [4-1:0] node1340;
	wire [4-1:0] node1343;
	wire [4-1:0] node1344;
	wire [4-1:0] node1347;
	wire [4-1:0] node1350;
	wire [4-1:0] node1351;
	wire [4-1:0] node1352;
	wire [4-1:0] node1353;
	wire [4-1:0] node1354;
	wire [4-1:0] node1358;
	wire [4-1:0] node1359;
	wire [4-1:0] node1363;
	wire [4-1:0] node1365;
	wire [4-1:0] node1366;
	wire [4-1:0] node1370;
	wire [4-1:0] node1371;
	wire [4-1:0] node1372;
	wire [4-1:0] node1375;
	wire [4-1:0] node1376;
	wire [4-1:0] node1380;
	wire [4-1:0] node1381;
	wire [4-1:0] node1382;
	wire [4-1:0] node1386;
	wire [4-1:0] node1387;
	wire [4-1:0] node1391;
	wire [4-1:0] node1392;
	wire [4-1:0] node1393;
	wire [4-1:0] node1394;
	wire [4-1:0] node1395;
	wire [4-1:0] node1396;
	wire [4-1:0] node1397;
	wire [4-1:0] node1398;
	wire [4-1:0] node1399;
	wire [4-1:0] node1400;
	wire [4-1:0] node1404;
	wire [4-1:0] node1406;
	wire [4-1:0] node1409;
	wire [4-1:0] node1410;
	wire [4-1:0] node1411;
	wire [4-1:0] node1414;
	wire [4-1:0] node1417;
	wire [4-1:0] node1420;
	wire [4-1:0] node1421;
	wire [4-1:0] node1422;
	wire [4-1:0] node1424;
	wire [4-1:0] node1428;
	wire [4-1:0] node1429;
	wire [4-1:0] node1430;
	wire [4-1:0] node1434;
	wire [4-1:0] node1435;
	wire [4-1:0] node1438;
	wire [4-1:0] node1441;
	wire [4-1:0] node1442;
	wire [4-1:0] node1443;
	wire [4-1:0] node1444;
	wire [4-1:0] node1445;
	wire [4-1:0] node1449;
	wire [4-1:0] node1450;
	wire [4-1:0] node1454;
	wire [4-1:0] node1455;
	wire [4-1:0] node1456;
	wire [4-1:0] node1459;
	wire [4-1:0] node1462;
	wire [4-1:0] node1464;
	wire [4-1:0] node1467;
	wire [4-1:0] node1468;
	wire [4-1:0] node1470;
	wire [4-1:0] node1473;
	wire [4-1:0] node1474;
	wire [4-1:0] node1475;
	wire [4-1:0] node1478;
	wire [4-1:0] node1481;
	wire [4-1:0] node1483;
	wire [4-1:0] node1486;
	wire [4-1:0] node1487;
	wire [4-1:0] node1488;
	wire [4-1:0] node1489;
	wire [4-1:0] node1490;
	wire [4-1:0] node1492;
	wire [4-1:0] node1495;
	wire [4-1:0] node1498;
	wire [4-1:0] node1499;
	wire [4-1:0] node1500;
	wire [4-1:0] node1503;
	wire [4-1:0] node1506;
	wire [4-1:0] node1508;
	wire [4-1:0] node1511;
	wire [4-1:0] node1512;
	wire [4-1:0] node1514;
	wire [4-1:0] node1515;
	wire [4-1:0] node1518;
	wire [4-1:0] node1521;
	wire [4-1:0] node1523;
	wire [4-1:0] node1524;
	wire [4-1:0] node1527;
	wire [4-1:0] node1530;
	wire [4-1:0] node1531;
	wire [4-1:0] node1532;
	wire [4-1:0] node1533;
	wire [4-1:0] node1535;
	wire [4-1:0] node1538;
	wire [4-1:0] node1539;
	wire [4-1:0] node1543;
	wire [4-1:0] node1544;
	wire [4-1:0] node1546;
	wire [4-1:0] node1549;
	wire [4-1:0] node1550;
	wire [4-1:0] node1554;
	wire [4-1:0] node1555;
	wire [4-1:0] node1556;
	wire [4-1:0] node1557;
	wire [4-1:0] node1561;
	wire [4-1:0] node1563;
	wire [4-1:0] node1566;
	wire [4-1:0] node1567;
	wire [4-1:0] node1568;
	wire [4-1:0] node1572;
	wire [4-1:0] node1574;
	wire [4-1:0] node1577;
	wire [4-1:0] node1578;
	wire [4-1:0] node1579;
	wire [4-1:0] node1580;
	wire [4-1:0] node1581;
	wire [4-1:0] node1582;
	wire [4-1:0] node1584;
	wire [4-1:0] node1587;
	wire [4-1:0] node1589;
	wire [4-1:0] node1592;
	wire [4-1:0] node1594;
	wire [4-1:0] node1596;
	wire [4-1:0] node1599;
	wire [4-1:0] node1600;
	wire [4-1:0] node1601;
	wire [4-1:0] node1603;
	wire [4-1:0] node1606;
	wire [4-1:0] node1607;
	wire [4-1:0] node1611;
	wire [4-1:0] node1612;
	wire [4-1:0] node1614;
	wire [4-1:0] node1617;
	wire [4-1:0] node1618;
	wire [4-1:0] node1622;
	wire [4-1:0] node1623;
	wire [4-1:0] node1624;
	wire [4-1:0] node1625;
	wire [4-1:0] node1628;
	wire [4-1:0] node1630;
	wire [4-1:0] node1633;
	wire [4-1:0] node1634;
	wire [4-1:0] node1635;
	wire [4-1:0] node1638;
	wire [4-1:0] node1641;
	wire [4-1:0] node1642;
	wire [4-1:0] node1646;
	wire [4-1:0] node1647;
	wire [4-1:0] node1648;
	wire [4-1:0] node1650;
	wire [4-1:0] node1653;
	wire [4-1:0] node1654;
	wire [4-1:0] node1657;
	wire [4-1:0] node1660;
	wire [4-1:0] node1661;
	wire [4-1:0] node1664;
	wire [4-1:0] node1665;
	wire [4-1:0] node1669;
	wire [4-1:0] node1670;
	wire [4-1:0] node1671;
	wire [4-1:0] node1672;
	wire [4-1:0] node1673;
	wire [4-1:0] node1675;
	wire [4-1:0] node1678;
	wire [4-1:0] node1681;
	wire [4-1:0] node1682;
	wire [4-1:0] node1683;
	wire [4-1:0] node1688;
	wire [4-1:0] node1689;
	wire [4-1:0] node1690;
	wire [4-1:0] node1692;
	wire [4-1:0] node1695;
	wire [4-1:0] node1696;
	wire [4-1:0] node1700;
	wire [4-1:0] node1701;
	wire [4-1:0] node1702;
	wire [4-1:0] node1705;
	wire [4-1:0] node1708;
	wire [4-1:0] node1709;
	wire [4-1:0] node1713;
	wire [4-1:0] node1714;
	wire [4-1:0] node1715;
	wire [4-1:0] node1716;
	wire [4-1:0] node1717;
	wire [4-1:0] node1722;
	wire [4-1:0] node1723;
	wire [4-1:0] node1724;
	wire [4-1:0] node1729;
	wire [4-1:0] node1730;
	wire [4-1:0] node1731;
	wire [4-1:0] node1734;
	wire [4-1:0] node1735;
	wire [4-1:0] node1738;
	wire [4-1:0] node1741;
	wire [4-1:0] node1742;
	wire [4-1:0] node1744;
	wire [4-1:0] node1747;
	wire [4-1:0] node1748;
	wire [4-1:0] node1751;
	wire [4-1:0] node1754;
	wire [4-1:0] node1755;
	wire [4-1:0] node1756;
	wire [4-1:0] node1757;
	wire [4-1:0] node1758;
	wire [4-1:0] node1759;
	wire [4-1:0] node1760;
	wire [4-1:0] node1761;
	wire [4-1:0] node1765;
	wire [4-1:0] node1768;
	wire [4-1:0] node1769;
	wire [4-1:0] node1770;
	wire [4-1:0] node1774;
	wire [4-1:0] node1777;
	wire [4-1:0] node1778;
	wire [4-1:0] node1779;
	wire [4-1:0] node1781;
	wire [4-1:0] node1784;
	wire [4-1:0] node1787;
	wire [4-1:0] node1788;
	wire [4-1:0] node1789;
	wire [4-1:0] node1793;
	wire [4-1:0] node1795;
	wire [4-1:0] node1798;
	wire [4-1:0] node1799;
	wire [4-1:0] node1800;
	wire [4-1:0] node1801;
	wire [4-1:0] node1802;
	wire [4-1:0] node1807;
	wire [4-1:0] node1808;
	wire [4-1:0] node1809;
	wire [4-1:0] node1814;
	wire [4-1:0] node1815;
	wire [4-1:0] node1816;
	wire [4-1:0] node1818;
	wire [4-1:0] node1821;
	wire [4-1:0] node1822;
	wire [4-1:0] node1826;
	wire [4-1:0] node1828;
	wire [4-1:0] node1830;
	wire [4-1:0] node1833;
	wire [4-1:0] node1834;
	wire [4-1:0] node1835;
	wire [4-1:0] node1836;
	wire [4-1:0] node1837;
	wire [4-1:0] node1839;
	wire [4-1:0] node1842;
	wire [4-1:0] node1843;
	wire [4-1:0] node1847;
	wire [4-1:0] node1848;
	wire [4-1:0] node1850;
	wire [4-1:0] node1853;
	wire [4-1:0] node1855;
	wire [4-1:0] node1858;
	wire [4-1:0] node1859;
	wire [4-1:0] node1860;
	wire [4-1:0] node1862;
	wire [4-1:0] node1865;
	wire [4-1:0] node1866;
	wire [4-1:0] node1870;
	wire [4-1:0] node1871;
	wire [4-1:0] node1874;
	wire [4-1:0] node1875;
	wire [4-1:0] node1879;
	wire [4-1:0] node1880;
	wire [4-1:0] node1881;
	wire [4-1:0] node1882;
	wire [4-1:0] node1883;
	wire [4-1:0] node1887;
	wire [4-1:0] node1889;
	wire [4-1:0] node1892;
	wire [4-1:0] node1893;
	wire [4-1:0] node1896;
	wire [4-1:0] node1898;
	wire [4-1:0] node1901;
	wire [4-1:0] node1902;
	wire [4-1:0] node1903;
	wire [4-1:0] node1905;
	wire [4-1:0] node1908;
	wire [4-1:0] node1909;
	wire [4-1:0] node1912;
	wire [4-1:0] node1915;
	wire [4-1:0] node1916;
	wire [4-1:0] node1918;
	wire [4-1:0] node1921;
	wire [4-1:0] node1923;
	wire [4-1:0] node1926;
	wire [4-1:0] node1927;
	wire [4-1:0] node1928;
	wire [4-1:0] node1929;
	wire [4-1:0] node1930;
	wire [4-1:0] node1932;
	wire [4-1:0] node1934;
	wire [4-1:0] node1937;
	wire [4-1:0] node1938;
	wire [4-1:0] node1939;
	wire [4-1:0] node1942;
	wire [4-1:0] node1945;
	wire [4-1:0] node1947;
	wire [4-1:0] node1950;
	wire [4-1:0] node1951;
	wire [4-1:0] node1952;
	wire [4-1:0] node1953;
	wire [4-1:0] node1957;
	wire [4-1:0] node1959;
	wire [4-1:0] node1962;
	wire [4-1:0] node1963;
	wire [4-1:0] node1967;
	wire [4-1:0] node1968;
	wire [4-1:0] node1969;
	wire [4-1:0] node1970;
	wire [4-1:0] node1971;
	wire [4-1:0] node1974;
	wire [4-1:0] node1977;
	wire [4-1:0] node1980;
	wire [4-1:0] node1981;
	wire [4-1:0] node1982;
	wire [4-1:0] node1985;
	wire [4-1:0] node1988;
	wire [4-1:0] node1989;
	wire [4-1:0] node1992;
	wire [4-1:0] node1995;
	wire [4-1:0] node1996;
	wire [4-1:0] node1997;
	wire [4-1:0] node1998;
	wire [4-1:0] node2001;
	wire [4-1:0] node2004;
	wire [4-1:0] node2006;
	wire [4-1:0] node2009;
	wire [4-1:0] node2010;
	wire [4-1:0] node2011;
	wire [4-1:0] node2014;
	wire [4-1:0] node2017;
	wire [4-1:0] node2018;
	wire [4-1:0] node2021;
	wire [4-1:0] node2024;
	wire [4-1:0] node2025;
	wire [4-1:0] node2026;
	wire [4-1:0] node2027;
	wire [4-1:0] node2028;
	wire [4-1:0] node2031;
	wire [4-1:0] node2032;
	wire [4-1:0] node2035;
	wire [4-1:0] node2038;
	wire [4-1:0] node2039;
	wire [4-1:0] node2040;
	wire [4-1:0] node2043;
	wire [4-1:0] node2046;
	wire [4-1:0] node2048;
	wire [4-1:0] node2051;
	wire [4-1:0] node2052;
	wire [4-1:0] node2053;
	wire [4-1:0] node2055;
	wire [4-1:0] node2059;
	wire [4-1:0] node2060;
	wire [4-1:0] node2061;
	wire [4-1:0] node2065;
	wire [4-1:0] node2066;
	wire [4-1:0] node2069;
	wire [4-1:0] node2072;
	wire [4-1:0] node2073;
	wire [4-1:0] node2074;
	wire [4-1:0] node2075;
	wire [4-1:0] node2076;
	wire [4-1:0] node2079;
	wire [4-1:0] node2083;
	wire [4-1:0] node2084;
	wire [4-1:0] node2085;
	wire [4-1:0] node2088;
	wire [4-1:0] node2091;
	wire [4-1:0] node2093;
	wire [4-1:0] node2096;
	wire [4-1:0] node2097;
	wire [4-1:0] node2098;
	wire [4-1:0] node2099;
	wire [4-1:0] node2103;
	wire [4-1:0] node2105;
	wire [4-1:0] node2108;
	wire [4-1:0] node2109;
	wire [4-1:0] node2110;
	wire [4-1:0] node2114;
	wire [4-1:0] node2115;
	wire [4-1:0] node2119;
	wire [4-1:0] node2120;
	wire [4-1:0] node2121;
	wire [4-1:0] node2122;
	wire [4-1:0] node2123;
	wire [4-1:0] node2124;
	wire [4-1:0] node2125;
	wire [4-1:0] node2126;
	wire [4-1:0] node2127;
	wire [4-1:0] node2132;
	wire [4-1:0] node2133;
	wire [4-1:0] node2134;
	wire [4-1:0] node2138;
	wire [4-1:0] node2139;
	wire [4-1:0] node2142;
	wire [4-1:0] node2145;
	wire [4-1:0] node2146;
	wire [4-1:0] node2147;
	wire [4-1:0] node2148;
	wire [4-1:0] node2152;
	wire [4-1:0] node2153;
	wire [4-1:0] node2157;
	wire [4-1:0] node2158;
	wire [4-1:0] node2159;
	wire [4-1:0] node2162;
	wire [4-1:0] node2165;
	wire [4-1:0] node2166;
	wire [4-1:0] node2169;
	wire [4-1:0] node2172;
	wire [4-1:0] node2173;
	wire [4-1:0] node2174;
	wire [4-1:0] node2175;
	wire [4-1:0] node2177;
	wire [4-1:0] node2180;
	wire [4-1:0] node2182;
	wire [4-1:0] node2185;
	wire [4-1:0] node2186;
	wire [4-1:0] node2188;
	wire [4-1:0] node2191;
	wire [4-1:0] node2194;
	wire [4-1:0] node2195;
	wire [4-1:0] node2196;
	wire [4-1:0] node2197;
	wire [4-1:0] node2202;
	wire [4-1:0] node2203;
	wire [4-1:0] node2205;
	wire [4-1:0] node2208;
	wire [4-1:0] node2209;
	wire [4-1:0] node2213;
	wire [4-1:0] node2214;
	wire [4-1:0] node2215;
	wire [4-1:0] node2216;
	wire [4-1:0] node2217;
	wire [4-1:0] node2218;
	wire [4-1:0] node2221;
	wire [4-1:0] node2224;
	wire [4-1:0] node2226;
	wire [4-1:0] node2229;
	wire [4-1:0] node2231;
	wire [4-1:0] node2232;
	wire [4-1:0] node2236;
	wire [4-1:0] node2237;
	wire [4-1:0] node2238;
	wire [4-1:0] node2240;
	wire [4-1:0] node2243;
	wire [4-1:0] node2245;
	wire [4-1:0] node2248;
	wire [4-1:0] node2250;
	wire [4-1:0] node2253;
	wire [4-1:0] node2254;
	wire [4-1:0] node2255;
	wire [4-1:0] node2256;
	wire [4-1:0] node2259;
	wire [4-1:0] node2261;
	wire [4-1:0] node2264;
	wire [4-1:0] node2265;
	wire [4-1:0] node2266;
	wire [4-1:0] node2269;
	wire [4-1:0] node2273;
	wire [4-1:0] node2274;
	wire [4-1:0] node2275;
	wire [4-1:0] node2277;
	wire [4-1:0] node2280;
	wire [4-1:0] node2282;
	wire [4-1:0] node2285;
	wire [4-1:0] node2286;
	wire [4-1:0] node2287;
	wire [4-1:0] node2290;
	wire [4-1:0] node2293;
	wire [4-1:0] node2294;
	wire [4-1:0] node2298;
	wire [4-1:0] node2299;
	wire [4-1:0] node2300;
	wire [4-1:0] node2301;
	wire [4-1:0] node2302;
	wire [4-1:0] node2303;
	wire [4-1:0] node2304;
	wire [4-1:0] node2308;
	wire [4-1:0] node2309;
	wire [4-1:0] node2312;
	wire [4-1:0] node2315;
	wire [4-1:0] node2316;
	wire [4-1:0] node2317;
	wire [4-1:0] node2320;
	wire [4-1:0] node2323;
	wire [4-1:0] node2324;
	wire [4-1:0] node2327;
	wire [4-1:0] node2330;
	wire [4-1:0] node2331;
	wire [4-1:0] node2332;
	wire [4-1:0] node2333;
	wire [4-1:0] node2338;
	wire [4-1:0] node2339;
	wire [4-1:0] node2340;
	wire [4-1:0] node2345;
	wire [4-1:0] node2346;
	wire [4-1:0] node2347;
	wire [4-1:0] node2348;
	wire [4-1:0] node2349;
	wire [4-1:0] node2352;
	wire [4-1:0] node2355;
	wire [4-1:0] node2357;
	wire [4-1:0] node2360;
	wire [4-1:0] node2361;
	wire [4-1:0] node2363;
	wire [4-1:0] node2366;
	wire [4-1:0] node2367;
	wire [4-1:0] node2370;
	wire [4-1:0] node2373;
	wire [4-1:0] node2374;
	wire [4-1:0] node2375;
	wire [4-1:0] node2376;
	wire [4-1:0] node2380;
	wire [4-1:0] node2381;
	wire [4-1:0] node2384;
	wire [4-1:0] node2387;
	wire [4-1:0] node2388;
	wire [4-1:0] node2391;
	wire [4-1:0] node2394;
	wire [4-1:0] node2395;
	wire [4-1:0] node2396;
	wire [4-1:0] node2397;
	wire [4-1:0] node2398;
	wire [4-1:0] node2400;
	wire [4-1:0] node2403;
	wire [4-1:0] node2405;
	wire [4-1:0] node2408;
	wire [4-1:0] node2409;
	wire [4-1:0] node2412;
	wire [4-1:0] node2413;
	wire [4-1:0] node2417;
	wire [4-1:0] node2418;
	wire [4-1:0] node2419;
	wire [4-1:0] node2421;
	wire [4-1:0] node2424;
	wire [4-1:0] node2425;
	wire [4-1:0] node2428;
	wire [4-1:0] node2431;
	wire [4-1:0] node2432;
	wire [4-1:0] node2433;
	wire [4-1:0] node2437;
	wire [4-1:0] node2438;
	wire [4-1:0] node2442;
	wire [4-1:0] node2443;
	wire [4-1:0] node2444;
	wire [4-1:0] node2445;
	wire [4-1:0] node2446;
	wire [4-1:0] node2450;
	wire [4-1:0] node2451;
	wire [4-1:0] node2455;
	wire [4-1:0] node2456;
	wire [4-1:0] node2457;
	wire [4-1:0] node2460;
	wire [4-1:0] node2463;
	wire [4-1:0] node2464;
	wire [4-1:0] node2467;
	wire [4-1:0] node2470;
	wire [4-1:0] node2471;
	wire [4-1:0] node2473;
	wire [4-1:0] node2475;
	wire [4-1:0] node2478;
	wire [4-1:0] node2480;
	wire [4-1:0] node2481;
	wire [4-1:0] node2485;
	wire [4-1:0] node2486;
	wire [4-1:0] node2487;
	wire [4-1:0] node2488;
	wire [4-1:0] node2489;
	wire [4-1:0] node2490;
	wire [4-1:0] node2491;
	wire [4-1:0] node2493;
	wire [4-1:0] node2496;
	wire [4-1:0] node2497;
	wire [4-1:0] node2501;
	wire [4-1:0] node2502;
	wire [4-1:0] node2503;
	wire [4-1:0] node2506;
	wire [4-1:0] node2509;
	wire [4-1:0] node2512;
	wire [4-1:0] node2513;
	wire [4-1:0] node2514;
	wire [4-1:0] node2515;
	wire [4-1:0] node2519;
	wire [4-1:0] node2520;
	wire [4-1:0] node2524;
	wire [4-1:0] node2525;
	wire [4-1:0] node2526;
	wire [4-1:0] node2529;
	wire [4-1:0] node2532;
	wire [4-1:0] node2533;
	wire [4-1:0] node2536;
	wire [4-1:0] node2539;
	wire [4-1:0] node2540;
	wire [4-1:0] node2541;
	wire [4-1:0] node2542;
	wire [4-1:0] node2544;
	wire [4-1:0] node2547;
	wire [4-1:0] node2550;
	wire [4-1:0] node2551;
	wire [4-1:0] node2553;
	wire [4-1:0] node2556;
	wire [4-1:0] node2559;
	wire [4-1:0] node2560;
	wire [4-1:0] node2561;
	wire [4-1:0] node2563;
	wire [4-1:0] node2566;
	wire [4-1:0] node2568;
	wire [4-1:0] node2571;
	wire [4-1:0] node2572;
	wire [4-1:0] node2573;
	wire [4-1:0] node2578;
	wire [4-1:0] node2579;
	wire [4-1:0] node2580;
	wire [4-1:0] node2581;
	wire [4-1:0] node2582;
	wire [4-1:0] node2583;
	wire [4-1:0] node2588;
	wire [4-1:0] node2589;
	wire [4-1:0] node2591;
	wire [4-1:0] node2594;
	wire [4-1:0] node2595;
	wire [4-1:0] node2599;
	wire [4-1:0] node2600;
	wire [4-1:0] node2601;
	wire [4-1:0] node2602;
	wire [4-1:0] node2605;
	wire [4-1:0] node2609;
	wire [4-1:0] node2610;
	wire [4-1:0] node2612;
	wire [4-1:0] node2615;
	wire [4-1:0] node2616;
	wire [4-1:0] node2620;
	wire [4-1:0] node2621;
	wire [4-1:0] node2622;
	wire [4-1:0] node2623;
	wire [4-1:0] node2624;
	wire [4-1:0] node2629;
	wire [4-1:0] node2630;
	wire [4-1:0] node2633;
	wire [4-1:0] node2634;
	wire [4-1:0] node2638;
	wire [4-1:0] node2639;
	wire [4-1:0] node2641;
	wire [4-1:0] node2643;
	wire [4-1:0] node2646;
	wire [4-1:0] node2647;
	wire [4-1:0] node2649;
	wire [4-1:0] node2653;
	wire [4-1:0] node2654;
	wire [4-1:0] node2655;
	wire [4-1:0] node2656;
	wire [4-1:0] node2657;
	wire [4-1:0] node2658;
	wire [4-1:0] node2660;
	wire [4-1:0] node2663;
	wire [4-1:0] node2665;
	wire [4-1:0] node2668;
	wire [4-1:0] node2669;
	wire [4-1:0] node2672;
	wire [4-1:0] node2673;
	wire [4-1:0] node2676;
	wire [4-1:0] node2679;
	wire [4-1:0] node2680;
	wire [4-1:0] node2681;
	wire [4-1:0] node2683;
	wire [4-1:0] node2686;
	wire [4-1:0] node2689;
	wire [4-1:0] node2690;
	wire [4-1:0] node2691;
	wire [4-1:0] node2695;
	wire [4-1:0] node2698;
	wire [4-1:0] node2699;
	wire [4-1:0] node2700;
	wire [4-1:0] node2701;
	wire [4-1:0] node2704;
	wire [4-1:0] node2706;
	wire [4-1:0] node2709;
	wire [4-1:0] node2710;
	wire [4-1:0] node2711;
	wire [4-1:0] node2715;
	wire [4-1:0] node2716;
	wire [4-1:0] node2720;
	wire [4-1:0] node2721;
	wire [4-1:0] node2722;
	wire [4-1:0] node2723;
	wire [4-1:0] node2726;
	wire [4-1:0] node2729;
	wire [4-1:0] node2730;
	wire [4-1:0] node2734;
	wire [4-1:0] node2736;
	wire [4-1:0] node2737;
	wire [4-1:0] node2740;
	wire [4-1:0] node2743;
	wire [4-1:0] node2744;
	wire [4-1:0] node2745;
	wire [4-1:0] node2746;
	wire [4-1:0] node2749;
	wire [4-1:0] node2750;
	wire [4-1:0] node2754;
	wire [4-1:0] node2755;
	wire [4-1:0] node2756;
	wire [4-1:0] node2757;
	wire [4-1:0] node2761;
	wire [4-1:0] node2762;
	wire [4-1:0] node2766;
	wire [4-1:0] node2767;
	wire [4-1:0] node2768;
	wire [4-1:0] node2771;
	wire [4-1:0] node2774;
	wire [4-1:0] node2775;
	wire [4-1:0] node2778;
	wire [4-1:0] node2781;
	wire [4-1:0] node2782;
	wire [4-1:0] node2783;
	wire [4-1:0] node2784;
	wire [4-1:0] node2785;
	wire [4-1:0] node2788;
	wire [4-1:0] node2791;
	wire [4-1:0] node2793;
	wire [4-1:0] node2796;
	wire [4-1:0] node2797;
	wire [4-1:0] node2800;
	wire [4-1:0] node2801;
	wire [4-1:0] node2805;
	wire [4-1:0] node2806;
	wire [4-1:0] node2807;
	wire [4-1:0] node2808;
	wire [4-1:0] node2811;
	wire [4-1:0] node2814;
	wire [4-1:0] node2817;
	wire [4-1:0] node2818;
	wire [4-1:0] node2821;
	wire [4-1:0] node2824;
	wire [4-1:0] node2825;
	wire [4-1:0] node2826;
	wire [4-1:0] node2827;
	wire [4-1:0] node2828;
	wire [4-1:0] node2829;
	wire [4-1:0] node2830;
	wire [4-1:0] node2831;
	wire [4-1:0] node2832;
	wire [4-1:0] node2833;
	wire [4-1:0] node2834;
	wire [4-1:0] node2838;
	wire [4-1:0] node2840;
	wire [4-1:0] node2843;
	wire [4-1:0] node2844;
	wire [4-1:0] node2845;
	wire [4-1:0] node2850;
	wire [4-1:0] node2851;
	wire [4-1:0] node2852;
	wire [4-1:0] node2855;
	wire [4-1:0] node2858;
	wire [4-1:0] node2859;
	wire [4-1:0] node2860;
	wire [4-1:0] node2865;
	wire [4-1:0] node2866;
	wire [4-1:0] node2867;
	wire [4-1:0] node2868;
	wire [4-1:0] node2870;
	wire [4-1:0] node2873;
	wire [4-1:0] node2875;
	wire [4-1:0] node2878;
	wire [4-1:0] node2879;
	wire [4-1:0] node2880;
	wire [4-1:0] node2885;
	wire [4-1:0] node2886;
	wire [4-1:0] node2887;
	wire [4-1:0] node2891;
	wire [4-1:0] node2892;
	wire [4-1:0] node2894;
	wire [4-1:0] node2897;
	wire [4-1:0] node2898;
	wire [4-1:0] node2902;
	wire [4-1:0] node2903;
	wire [4-1:0] node2904;
	wire [4-1:0] node2905;
	wire [4-1:0] node2906;
	wire [4-1:0] node2909;
	wire [4-1:0] node2912;
	wire [4-1:0] node2913;
	wire [4-1:0] node2917;
	wire [4-1:0] node2918;
	wire [4-1:0] node2919;
	wire [4-1:0] node2920;
	wire [4-1:0] node2924;
	wire [4-1:0] node2927;
	wire [4-1:0] node2929;
	wire [4-1:0] node2930;
	wire [4-1:0] node2934;
	wire [4-1:0] node2935;
	wire [4-1:0] node2936;
	wire [4-1:0] node2937;
	wire [4-1:0] node2938;
	wire [4-1:0] node2942;
	wire [4-1:0] node2945;
	wire [4-1:0] node2946;
	wire [4-1:0] node2949;
	wire [4-1:0] node2950;
	wire [4-1:0] node2954;
	wire [4-1:0] node2955;
	wire [4-1:0] node2957;
	wire [4-1:0] node2958;
	wire [4-1:0] node2961;
	wire [4-1:0] node2964;
	wire [4-1:0] node2965;
	wire [4-1:0] node2966;
	wire [4-1:0] node2969;
	wire [4-1:0] node2972;
	wire [4-1:0] node2973;
	wire [4-1:0] node2977;
	wire [4-1:0] node2978;
	wire [4-1:0] node2979;
	wire [4-1:0] node2980;
	wire [4-1:0] node2981;
	wire [4-1:0] node2982;
	wire [4-1:0] node2985;
	wire [4-1:0] node2986;
	wire [4-1:0] node2990;
	wire [4-1:0] node2991;
	wire [4-1:0] node2993;
	wire [4-1:0] node2997;
	wire [4-1:0] node2998;
	wire [4-1:0] node2999;
	wire [4-1:0] node3003;
	wire [4-1:0] node3004;
	wire [4-1:0] node3008;
	wire [4-1:0] node3009;
	wire [4-1:0] node3010;
	wire [4-1:0] node3011;
	wire [4-1:0] node3014;
	wire [4-1:0] node3016;
	wire [4-1:0] node3019;
	wire [4-1:0] node3021;
	wire [4-1:0] node3022;
	wire [4-1:0] node3025;
	wire [4-1:0] node3028;
	wire [4-1:0] node3029;
	wire [4-1:0] node3030;
	wire [4-1:0] node3031;
	wire [4-1:0] node3035;
	wire [4-1:0] node3037;
	wire [4-1:0] node3040;
	wire [4-1:0] node3041;
	wire [4-1:0] node3042;
	wire [4-1:0] node3046;
	wire [4-1:0] node3048;
	wire [4-1:0] node3051;
	wire [4-1:0] node3052;
	wire [4-1:0] node3053;
	wire [4-1:0] node3054;
	wire [4-1:0] node3056;
	wire [4-1:0] node3058;
	wire [4-1:0] node3061;
	wire [4-1:0] node3062;
	wire [4-1:0] node3064;
	wire [4-1:0] node3067;
	wire [4-1:0] node3069;
	wire [4-1:0] node3072;
	wire [4-1:0] node3073;
	wire [4-1:0] node3074;
	wire [4-1:0] node3075;
	wire [4-1:0] node3079;
	wire [4-1:0] node3081;
	wire [4-1:0] node3084;
	wire [4-1:0] node3085;
	wire [4-1:0] node3086;
	wire [4-1:0] node3089;
	wire [4-1:0] node3092;
	wire [4-1:0] node3093;
	wire [4-1:0] node3097;
	wire [4-1:0] node3098;
	wire [4-1:0] node3099;
	wire [4-1:0] node3100;
	wire [4-1:0] node3101;
	wire [4-1:0] node3105;
	wire [4-1:0] node3106;
	wire [4-1:0] node3109;
	wire [4-1:0] node3112;
	wire [4-1:0] node3113;
	wire [4-1:0] node3114;
	wire [4-1:0] node3117;
	wire [4-1:0] node3120;
	wire [4-1:0] node3122;
	wire [4-1:0] node3125;
	wire [4-1:0] node3126;
	wire [4-1:0] node3127;
	wire [4-1:0] node3130;
	wire [4-1:0] node3131;
	wire [4-1:0] node3135;
	wire [4-1:0] node3136;
	wire [4-1:0] node3137;
	wire [4-1:0] node3140;
	wire [4-1:0] node3143;
	wire [4-1:0] node3144;
	wire [4-1:0] node3147;
	wire [4-1:0] node3150;
	wire [4-1:0] node3151;
	wire [4-1:0] node3152;
	wire [4-1:0] node3153;
	wire [4-1:0] node3154;
	wire [4-1:0] node3155;
	wire [4-1:0] node3156;
	wire [4-1:0] node3158;
	wire [4-1:0] node3162;
	wire [4-1:0] node3163;
	wire [4-1:0] node3164;
	wire [4-1:0] node3168;
	wire [4-1:0] node3169;
	wire [4-1:0] node3173;
	wire [4-1:0] node3174;
	wire [4-1:0] node3176;
	wire [4-1:0] node3177;
	wire [4-1:0] node3181;
	wire [4-1:0] node3182;
	wire [4-1:0] node3185;
	wire [4-1:0] node3188;
	wire [4-1:0] node3189;
	wire [4-1:0] node3190;
	wire [4-1:0] node3191;
	wire [4-1:0] node3192;
	wire [4-1:0] node3196;
	wire [4-1:0] node3199;
	wire [4-1:0] node3200;
	wire [4-1:0] node3202;
	wire [4-1:0] node3205;
	wire [4-1:0] node3207;
	wire [4-1:0] node3210;
	wire [4-1:0] node3211;
	wire [4-1:0] node3212;
	wire [4-1:0] node3214;
	wire [4-1:0] node3217;
	wire [4-1:0] node3219;
	wire [4-1:0] node3222;
	wire [4-1:0] node3223;
	wire [4-1:0] node3225;
	wire [4-1:0] node3228;
	wire [4-1:0] node3231;
	wire [4-1:0] node3232;
	wire [4-1:0] node3233;
	wire [4-1:0] node3234;
	wire [4-1:0] node3235;
	wire [4-1:0] node3236;
	wire [4-1:0] node3241;
	wire [4-1:0] node3242;
	wire [4-1:0] node3244;
	wire [4-1:0] node3247;
	wire [4-1:0] node3249;
	wire [4-1:0] node3252;
	wire [4-1:0] node3253;
	wire [4-1:0] node3254;
	wire [4-1:0] node3255;
	wire [4-1:0] node3259;
	wire [4-1:0] node3260;
	wire [4-1:0] node3264;
	wire [4-1:0] node3265;
	wire [4-1:0] node3269;
	wire [4-1:0] node3270;
	wire [4-1:0] node3271;
	wire [4-1:0] node3272;
	wire [4-1:0] node3273;
	wire [4-1:0] node3276;
	wire [4-1:0] node3279;
	wire [4-1:0] node3280;
	wire [4-1:0] node3284;
	wire [4-1:0] node3285;
	wire [4-1:0] node3286;
	wire [4-1:0] node3290;
	wire [4-1:0] node3292;
	wire [4-1:0] node3295;
	wire [4-1:0] node3296;
	wire [4-1:0] node3297;
	wire [4-1:0] node3299;
	wire [4-1:0] node3302;
	wire [4-1:0] node3305;
	wire [4-1:0] node3306;
	wire [4-1:0] node3309;
	wire [4-1:0] node3310;
	wire [4-1:0] node3313;
	wire [4-1:0] node3316;
	wire [4-1:0] node3317;
	wire [4-1:0] node3318;
	wire [4-1:0] node3319;
	wire [4-1:0] node3320;
	wire [4-1:0] node3321;
	wire [4-1:0] node3323;
	wire [4-1:0] node3326;
	wire [4-1:0] node3327;
	wire [4-1:0] node3331;
	wire [4-1:0] node3332;
	wire [4-1:0] node3333;
	wire [4-1:0] node3337;
	wire [4-1:0] node3338;
	wire [4-1:0] node3341;
	wire [4-1:0] node3344;
	wire [4-1:0] node3345;
	wire [4-1:0] node3346;
	wire [4-1:0] node3349;
	wire [4-1:0] node3350;
	wire [4-1:0] node3354;
	wire [4-1:0] node3355;
	wire [4-1:0] node3357;
	wire [4-1:0] node3361;
	wire [4-1:0] node3362;
	wire [4-1:0] node3363;
	wire [4-1:0] node3364;
	wire [4-1:0] node3365;
	wire [4-1:0] node3368;
	wire [4-1:0] node3371;
	wire [4-1:0] node3373;
	wire [4-1:0] node3376;
	wire [4-1:0] node3377;
	wire [4-1:0] node3378;
	wire [4-1:0] node3382;
	wire [4-1:0] node3383;
	wire [4-1:0] node3387;
	wire [4-1:0] node3388;
	wire [4-1:0] node3389;
	wire [4-1:0] node3390;
	wire [4-1:0] node3395;
	wire [4-1:0] node3396;
	wire [4-1:0] node3399;
	wire [4-1:0] node3400;
	wire [4-1:0] node3404;
	wire [4-1:0] node3405;
	wire [4-1:0] node3406;
	wire [4-1:0] node3407;
	wire [4-1:0] node3408;
	wire [4-1:0] node3409;
	wire [4-1:0] node3413;
	wire [4-1:0] node3416;
	wire [4-1:0] node3417;
	wire [4-1:0] node3421;
	wire [4-1:0] node3422;
	wire [4-1:0] node3423;
	wire [4-1:0] node3426;
	wire [4-1:0] node3428;
	wire [4-1:0] node3431;
	wire [4-1:0] node3432;
	wire [4-1:0] node3433;
	wire [4-1:0] node3436;
	wire [4-1:0] node3439;
	wire [4-1:0] node3440;
	wire [4-1:0] node3443;
	wire [4-1:0] node3446;
	wire [4-1:0] node3447;
	wire [4-1:0] node3448;
	wire [4-1:0] node3450;
	wire [4-1:0] node3451;
	wire [4-1:0] node3455;
	wire [4-1:0] node3457;
	wire [4-1:0] node3460;
	wire [4-1:0] node3461;
	wire [4-1:0] node3462;
	wire [4-1:0] node3464;
	wire [4-1:0] node3467;
	wire [4-1:0] node3469;
	wire [4-1:0] node3472;
	wire [4-1:0] node3473;
	wire [4-1:0] node3474;
	wire [4-1:0] node3478;
	wire [4-1:0] node3481;
	wire [4-1:0] node3482;
	wire [4-1:0] node3483;
	wire [4-1:0] node3484;
	wire [4-1:0] node3485;
	wire [4-1:0] node3486;
	wire [4-1:0] node3487;
	wire [4-1:0] node3488;
	wire [4-1:0] node3490;
	wire [4-1:0] node3493;
	wire [4-1:0] node3495;
	wire [4-1:0] node3498;
	wire [4-1:0] node3499;
	wire [4-1:0] node3500;
	wire [4-1:0] node3504;
	wire [4-1:0] node3506;
	wire [4-1:0] node3509;
	wire [4-1:0] node3510;
	wire [4-1:0] node3511;
	wire [4-1:0] node3512;
	wire [4-1:0] node3515;
	wire [4-1:0] node3518;
	wire [4-1:0] node3520;
	wire [4-1:0] node3523;
	wire [4-1:0] node3524;
	wire [4-1:0] node3525;
	wire [4-1:0] node3530;
	wire [4-1:0] node3531;
	wire [4-1:0] node3532;
	wire [4-1:0] node3533;
	wire [4-1:0] node3535;
	wire [4-1:0] node3538;
	wire [4-1:0] node3540;
	wire [4-1:0] node3543;
	wire [4-1:0] node3544;
	wire [4-1:0] node3545;
	wire [4-1:0] node3550;
	wire [4-1:0] node3551;
	wire [4-1:0] node3552;
	wire [4-1:0] node3554;
	wire [4-1:0] node3557;
	wire [4-1:0] node3559;
	wire [4-1:0] node3562;
	wire [4-1:0] node3564;
	wire [4-1:0] node3565;
	wire [4-1:0] node3568;
	wire [4-1:0] node3571;
	wire [4-1:0] node3572;
	wire [4-1:0] node3573;
	wire [4-1:0] node3574;
	wire [4-1:0] node3575;
	wire [4-1:0] node3576;
	wire [4-1:0] node3579;
	wire [4-1:0] node3582;
	wire [4-1:0] node3583;
	wire [4-1:0] node3586;
	wire [4-1:0] node3589;
	wire [4-1:0] node3591;
	wire [4-1:0] node3592;
	wire [4-1:0] node3595;
	wire [4-1:0] node3598;
	wire [4-1:0] node3599;
	wire [4-1:0] node3600;
	wire [4-1:0] node3601;
	wire [4-1:0] node3605;
	wire [4-1:0] node3606;
	wire [4-1:0] node3610;
	wire [4-1:0] node3611;
	wire [4-1:0] node3613;
	wire [4-1:0] node3616;
	wire [4-1:0] node3618;
	wire [4-1:0] node3621;
	wire [4-1:0] node3622;
	wire [4-1:0] node3623;
	wire [4-1:0] node3625;
	wire [4-1:0] node3628;
	wire [4-1:0] node3629;
	wire [4-1:0] node3631;
	wire [4-1:0] node3634;
	wire [4-1:0] node3636;
	wire [4-1:0] node3639;
	wire [4-1:0] node3640;
	wire [4-1:0] node3642;
	wire [4-1:0] node3644;
	wire [4-1:0] node3647;
	wire [4-1:0] node3648;
	wire [4-1:0] node3651;
	wire [4-1:0] node3652;
	wire [4-1:0] node3655;
	wire [4-1:0] node3658;
	wire [4-1:0] node3659;
	wire [4-1:0] node3660;
	wire [4-1:0] node3661;
	wire [4-1:0] node3662;
	wire [4-1:0] node3663;
	wire [4-1:0] node3665;
	wire [4-1:0] node3669;
	wire [4-1:0] node3670;
	wire [4-1:0] node3673;
	wire [4-1:0] node3676;
	wire [4-1:0] node3677;
	wire [4-1:0] node3678;
	wire [4-1:0] node3679;
	wire [4-1:0] node3684;
	wire [4-1:0] node3685;
	wire [4-1:0] node3687;
	wire [4-1:0] node3690;
	wire [4-1:0] node3691;
	wire [4-1:0] node3694;
	wire [4-1:0] node3697;
	wire [4-1:0] node3698;
	wire [4-1:0] node3699;
	wire [4-1:0] node3700;
	wire [4-1:0] node3702;
	wire [4-1:0] node3706;
	wire [4-1:0] node3707;
	wire [4-1:0] node3710;
	wire [4-1:0] node3711;
	wire [4-1:0] node3714;
	wire [4-1:0] node3717;
	wire [4-1:0] node3718;
	wire [4-1:0] node3719;
	wire [4-1:0] node3721;
	wire [4-1:0] node3725;
	wire [4-1:0] node3726;
	wire [4-1:0] node3728;
	wire [4-1:0] node3731;
	wire [4-1:0] node3732;
	wire [4-1:0] node3736;
	wire [4-1:0] node3737;
	wire [4-1:0] node3738;
	wire [4-1:0] node3739;
	wire [4-1:0] node3740;
	wire [4-1:0] node3741;
	wire [4-1:0] node3745;
	wire [4-1:0] node3748;
	wire [4-1:0] node3749;
	wire [4-1:0] node3751;
	wire [4-1:0] node3754;
	wire [4-1:0] node3757;
	wire [4-1:0] node3758;
	wire [4-1:0] node3759;
	wire [4-1:0] node3761;
	wire [4-1:0] node3765;
	wire [4-1:0] node3767;
	wire [4-1:0] node3768;
	wire [4-1:0] node3771;
	wire [4-1:0] node3774;
	wire [4-1:0] node3775;
	wire [4-1:0] node3776;
	wire [4-1:0] node3777;
	wire [4-1:0] node3779;
	wire [4-1:0] node3782;
	wire [4-1:0] node3783;
	wire [4-1:0] node3786;
	wire [4-1:0] node3789;
	wire [4-1:0] node3790;
	wire [4-1:0] node3792;
	wire [4-1:0] node3795;
	wire [4-1:0] node3796;
	wire [4-1:0] node3799;
	wire [4-1:0] node3802;
	wire [4-1:0] node3803;
	wire [4-1:0] node3804;
	wire [4-1:0] node3805;
	wire [4-1:0] node3809;
	wire [4-1:0] node3810;
	wire [4-1:0] node3813;
	wire [4-1:0] node3816;
	wire [4-1:0] node3817;
	wire [4-1:0] node3819;
	wire [4-1:0] node3822;
	wire [4-1:0] node3823;
	wire [4-1:0] node3826;
	wire [4-1:0] node3829;
	wire [4-1:0] node3830;
	wire [4-1:0] node3831;
	wire [4-1:0] node3832;
	wire [4-1:0] node3833;
	wire [4-1:0] node3834;
	wire [4-1:0] node3836;
	wire [4-1:0] node3837;
	wire [4-1:0] node3840;
	wire [4-1:0] node3843;
	wire [4-1:0] node3844;
	wire [4-1:0] node3847;
	wire [4-1:0] node3849;
	wire [4-1:0] node3852;
	wire [4-1:0] node3853;
	wire [4-1:0] node3855;
	wire [4-1:0] node3856;
	wire [4-1:0] node3859;
	wire [4-1:0] node3862;
	wire [4-1:0] node3863;
	wire [4-1:0] node3864;
	wire [4-1:0] node3867;
	wire [4-1:0] node3871;
	wire [4-1:0] node3872;
	wire [4-1:0] node3873;
	wire [4-1:0] node3874;
	wire [4-1:0] node3876;
	wire [4-1:0] node3880;
	wire [4-1:0] node3881;
	wire [4-1:0] node3883;
	wire [4-1:0] node3886;
	wire [4-1:0] node3887;
	wire [4-1:0] node3890;
	wire [4-1:0] node3893;
	wire [4-1:0] node3894;
	wire [4-1:0] node3895;
	wire [4-1:0] node3896;
	wire [4-1:0] node3899;
	wire [4-1:0] node3902;
	wire [4-1:0] node3904;
	wire [4-1:0] node3907;
	wire [4-1:0] node3909;
	wire [4-1:0] node3910;
	wire [4-1:0] node3913;
	wire [4-1:0] node3916;
	wire [4-1:0] node3917;
	wire [4-1:0] node3918;
	wire [4-1:0] node3919;
	wire [4-1:0] node3920;
	wire [4-1:0] node3921;
	wire [4-1:0] node3925;
	wire [4-1:0] node3927;
	wire [4-1:0] node3930;
	wire [4-1:0] node3932;
	wire [4-1:0] node3933;
	wire [4-1:0] node3937;
	wire [4-1:0] node3938;
	wire [4-1:0] node3939;
	wire [4-1:0] node3942;
	wire [4-1:0] node3945;
	wire [4-1:0] node3946;
	wire [4-1:0] node3947;
	wire [4-1:0] node3951;
	wire [4-1:0] node3954;
	wire [4-1:0] node3955;
	wire [4-1:0] node3956;
	wire [4-1:0] node3957;
	wire [4-1:0] node3958;
	wire [4-1:0] node3961;
	wire [4-1:0] node3964;
	wire [4-1:0] node3965;
	wire [4-1:0] node3969;
	wire [4-1:0] node3970;
	wire [4-1:0] node3974;
	wire [4-1:0] node3975;
	wire [4-1:0] node3976;
	wire [4-1:0] node3977;
	wire [4-1:0] node3980;
	wire [4-1:0] node3983;
	wire [4-1:0] node3985;
	wire [4-1:0] node3988;
	wire [4-1:0] node3989;
	wire [4-1:0] node3990;
	wire [4-1:0] node3994;
	wire [4-1:0] node3995;
	wire [4-1:0] node3999;
	wire [4-1:0] node4000;
	wire [4-1:0] node4001;
	wire [4-1:0] node4002;
	wire [4-1:0] node4003;
	wire [4-1:0] node4004;
	wire [4-1:0] node4006;
	wire [4-1:0] node4009;
	wire [4-1:0] node4012;
	wire [4-1:0] node4013;
	wire [4-1:0] node4015;
	wire [4-1:0] node4018;
	wire [4-1:0] node4020;
	wire [4-1:0] node4023;
	wire [4-1:0] node4024;
	wire [4-1:0] node4025;
	wire [4-1:0] node4027;
	wire [4-1:0] node4030;
	wire [4-1:0] node4032;
	wire [4-1:0] node4035;
	wire [4-1:0] node4036;
	wire [4-1:0] node4038;
	wire [4-1:0] node4041;
	wire [4-1:0] node4043;
	wire [4-1:0] node4046;
	wire [4-1:0] node4047;
	wire [4-1:0] node4048;
	wire [4-1:0] node4049;
	wire [4-1:0] node4050;
	wire [4-1:0] node4054;
	wire [4-1:0] node4056;
	wire [4-1:0] node4059;
	wire [4-1:0] node4060;
	wire [4-1:0] node4061;
	wire [4-1:0] node4065;
	wire [4-1:0] node4066;
	wire [4-1:0] node4070;
	wire [4-1:0] node4071;
	wire [4-1:0] node4072;
	wire [4-1:0] node4073;
	wire [4-1:0] node4077;
	wire [4-1:0] node4079;
	wire [4-1:0] node4082;
	wire [4-1:0] node4083;
	wire [4-1:0] node4084;
	wire [4-1:0] node4087;
	wire [4-1:0] node4090;
	wire [4-1:0] node4092;
	wire [4-1:0] node4095;
	wire [4-1:0] node4096;
	wire [4-1:0] node4097;
	wire [4-1:0] node4098;
	wire [4-1:0] node4100;
	wire [4-1:0] node4103;
	wire [4-1:0] node4105;
	wire [4-1:0] node4107;
	wire [4-1:0] node4110;
	wire [4-1:0] node4111;
	wire [4-1:0] node4112;
	wire [4-1:0] node4113;
	wire [4-1:0] node4116;
	wire [4-1:0] node4119;
	wire [4-1:0] node4120;
	wire [4-1:0] node4124;
	wire [4-1:0] node4125;
	wire [4-1:0] node4128;
	wire [4-1:0] node4129;
	wire [4-1:0] node4132;
	wire [4-1:0] node4135;
	wire [4-1:0] node4136;
	wire [4-1:0] node4137;
	wire [4-1:0] node4138;
	wire [4-1:0] node4139;
	wire [4-1:0] node4142;
	wire [4-1:0] node4146;
	wire [4-1:0] node4147;
	wire [4-1:0] node4148;
	wire [4-1:0] node4153;
	wire [4-1:0] node4154;
	wire [4-1:0] node4155;
	wire [4-1:0] node4156;
	wire [4-1:0] node4159;
	wire [4-1:0] node4162;
	wire [4-1:0] node4163;
	wire [4-1:0] node4166;
	wire [4-1:0] node4169;
	wire [4-1:0] node4170;
	wire [4-1:0] node4171;
	wire [4-1:0] node4174;
	wire [4-1:0] node4177;
	wire [4-1:0] node4179;
	wire [4-1:0] node4182;
	wire [4-1:0] node4183;
	wire [4-1:0] node4184;
	wire [4-1:0] node4185;
	wire [4-1:0] node4186;
	wire [4-1:0] node4187;
	wire [4-1:0] node4188;
	wire [4-1:0] node4189;
	wire [4-1:0] node4190;
	wire [4-1:0] node4192;
	wire [4-1:0] node4195;
	wire [4-1:0] node4197;
	wire [4-1:0] node4200;
	wire [4-1:0] node4201;
	wire [4-1:0] node4202;
	wire [4-1:0] node4206;
	wire [4-1:0] node4207;
	wire [4-1:0] node4211;
	wire [4-1:0] node4212;
	wire [4-1:0] node4213;
	wire [4-1:0] node4214;
	wire [4-1:0] node4218;
	wire [4-1:0] node4220;
	wire [4-1:0] node4223;
	wire [4-1:0] node4224;
	wire [4-1:0] node4225;
	wire [4-1:0] node4228;
	wire [4-1:0] node4231;
	wire [4-1:0] node4232;
	wire [4-1:0] node4236;
	wire [4-1:0] node4237;
	wire [4-1:0] node4238;
	wire [4-1:0] node4239;
	wire [4-1:0] node4240;
	wire [4-1:0] node4244;
	wire [4-1:0] node4245;
	wire [4-1:0] node4249;
	wire [4-1:0] node4250;
	wire [4-1:0] node4251;
	wire [4-1:0] node4254;
	wire [4-1:0] node4257;
	wire [4-1:0] node4258;
	wire [4-1:0] node4262;
	wire [4-1:0] node4263;
	wire [4-1:0] node4264;
	wire [4-1:0] node4266;
	wire [4-1:0] node4269;
	wire [4-1:0] node4272;
	wire [4-1:0] node4273;
	wire [4-1:0] node4274;
	wire [4-1:0] node4277;
	wire [4-1:0] node4280;
	wire [4-1:0] node4281;
	wire [4-1:0] node4284;
	wire [4-1:0] node4287;
	wire [4-1:0] node4288;
	wire [4-1:0] node4289;
	wire [4-1:0] node4290;
	wire [4-1:0] node4291;
	wire [4-1:0] node4292;
	wire [4-1:0] node4296;
	wire [4-1:0] node4298;
	wire [4-1:0] node4301;
	wire [4-1:0] node4302;
	wire [4-1:0] node4303;
	wire [4-1:0] node4306;
	wire [4-1:0] node4309;
	wire [4-1:0] node4310;
	wire [4-1:0] node4314;
	wire [4-1:0] node4315;
	wire [4-1:0] node4316;
	wire [4-1:0] node4317;
	wire [4-1:0] node4320;
	wire [4-1:0] node4323;
	wire [4-1:0] node4324;
	wire [4-1:0] node4327;
	wire [4-1:0] node4330;
	wire [4-1:0] node4331;
	wire [4-1:0] node4334;
	wire [4-1:0] node4337;
	wire [4-1:0] node4338;
	wire [4-1:0] node4339;
	wire [4-1:0] node4340;
	wire [4-1:0] node4341;
	wire [4-1:0] node4345;
	wire [4-1:0] node4346;
	wire [4-1:0] node4350;
	wire [4-1:0] node4351;
	wire [4-1:0] node4352;
	wire [4-1:0] node4356;
	wire [4-1:0] node4357;
	wire [4-1:0] node4360;
	wire [4-1:0] node4363;
	wire [4-1:0] node4364;
	wire [4-1:0] node4365;
	wire [4-1:0] node4366;
	wire [4-1:0] node4369;
	wire [4-1:0] node4372;
	wire [4-1:0] node4374;
	wire [4-1:0] node4377;
	wire [4-1:0] node4378;
	wire [4-1:0] node4379;
	wire [4-1:0] node4383;
	wire [4-1:0] node4384;
	wire [4-1:0] node4388;
	wire [4-1:0] node4389;
	wire [4-1:0] node4390;
	wire [4-1:0] node4391;
	wire [4-1:0] node4392;
	wire [4-1:0] node4393;
	wire [4-1:0] node4394;
	wire [4-1:0] node4398;
	wire [4-1:0] node4399;
	wire [4-1:0] node4402;
	wire [4-1:0] node4405;
	wire [4-1:0] node4406;
	wire [4-1:0] node4408;
	wire [4-1:0] node4411;
	wire [4-1:0] node4412;
	wire [4-1:0] node4415;
	wire [4-1:0] node4418;
	wire [4-1:0] node4419;
	wire [4-1:0] node4420;
	wire [4-1:0] node4421;
	wire [4-1:0] node4425;
	wire [4-1:0] node4427;
	wire [4-1:0] node4430;
	wire [4-1:0] node4431;
	wire [4-1:0] node4432;
	wire [4-1:0] node4436;
	wire [4-1:0] node4439;
	wire [4-1:0] node4440;
	wire [4-1:0] node4441;
	wire [4-1:0] node4443;
	wire [4-1:0] node4445;
	wire [4-1:0] node4448;
	wire [4-1:0] node4449;
	wire [4-1:0] node4451;
	wire [4-1:0] node4454;
	wire [4-1:0] node4455;
	wire [4-1:0] node4458;
	wire [4-1:0] node4461;
	wire [4-1:0] node4462;
	wire [4-1:0] node4463;
	wire [4-1:0] node4464;
	wire [4-1:0] node4468;
	wire [4-1:0] node4469;
	wire [4-1:0] node4473;
	wire [4-1:0] node4474;
	wire [4-1:0] node4475;
	wire [4-1:0] node4478;
	wire [4-1:0] node4481;
	wire [4-1:0] node4483;
	wire [4-1:0] node4486;
	wire [4-1:0] node4487;
	wire [4-1:0] node4488;
	wire [4-1:0] node4489;
	wire [4-1:0] node4490;
	wire [4-1:0] node4491;
	wire [4-1:0] node4495;
	wire [4-1:0] node4496;
	wire [4-1:0] node4499;
	wire [4-1:0] node4502;
	wire [4-1:0] node4503;
	wire [4-1:0] node4504;
	wire [4-1:0] node4508;
	wire [4-1:0] node4509;
	wire [4-1:0] node4512;
	wire [4-1:0] node4515;
	wire [4-1:0] node4516;
	wire [4-1:0] node4517;
	wire [4-1:0] node4518;
	wire [4-1:0] node4521;
	wire [4-1:0] node4524;
	wire [4-1:0] node4525;
	wire [4-1:0] node4529;
	wire [4-1:0] node4530;
	wire [4-1:0] node4531;
	wire [4-1:0] node4534;
	wire [4-1:0] node4537;
	wire [4-1:0] node4540;
	wire [4-1:0] node4541;
	wire [4-1:0] node4542;
	wire [4-1:0] node4543;
	wire [4-1:0] node4545;
	wire [4-1:0] node4548;
	wire [4-1:0] node4549;
	wire [4-1:0] node4553;
	wire [4-1:0] node4554;
	wire [4-1:0] node4557;
	wire [4-1:0] node4560;
	wire [4-1:0] node4561;
	wire [4-1:0] node4562;
	wire [4-1:0] node4564;
	wire [4-1:0] node4568;
	wire [4-1:0] node4569;
	wire [4-1:0] node4571;
	wire [4-1:0] node4574;
	wire [4-1:0] node4575;
	wire [4-1:0] node4579;
	wire [4-1:0] node4580;
	wire [4-1:0] node4581;
	wire [4-1:0] node4582;
	wire [4-1:0] node4583;
	wire [4-1:0] node4584;
	wire [4-1:0] node4585;
	wire [4-1:0] node4588;
	wire [4-1:0] node4589;
	wire [4-1:0] node4593;
	wire [4-1:0] node4594;
	wire [4-1:0] node4595;
	wire [4-1:0] node4599;
	wire [4-1:0] node4600;
	wire [4-1:0] node4604;
	wire [4-1:0] node4605;
	wire [4-1:0] node4606;
	wire [4-1:0] node4607;
	wire [4-1:0] node4611;
	wire [4-1:0] node4612;
	wire [4-1:0] node4616;
	wire [4-1:0] node4617;
	wire [4-1:0] node4619;
	wire [4-1:0] node4622;
	wire [4-1:0] node4624;
	wire [4-1:0] node4627;
	wire [4-1:0] node4628;
	wire [4-1:0] node4629;
	wire [4-1:0] node4630;
	wire [4-1:0] node4631;
	wire [4-1:0] node4634;
	wire [4-1:0] node4637;
	wire [4-1:0] node4639;
	wire [4-1:0] node4642;
	wire [4-1:0] node4643;
	wire [4-1:0] node4646;
	wire [4-1:0] node4647;
	wire [4-1:0] node4651;
	wire [4-1:0] node4652;
	wire [4-1:0] node4653;
	wire [4-1:0] node4654;
	wire [4-1:0] node4657;
	wire [4-1:0] node4660;
	wire [4-1:0] node4661;
	wire [4-1:0] node4664;
	wire [4-1:0] node4667;
	wire [4-1:0] node4668;
	wire [4-1:0] node4670;
	wire [4-1:0] node4673;
	wire [4-1:0] node4674;
	wire [4-1:0] node4678;
	wire [4-1:0] node4679;
	wire [4-1:0] node4680;
	wire [4-1:0] node4681;
	wire [4-1:0] node4682;
	wire [4-1:0] node4683;
	wire [4-1:0] node4687;
	wire [4-1:0] node4689;
	wire [4-1:0] node4692;
	wire [4-1:0] node4694;
	wire [4-1:0] node4696;
	wire [4-1:0] node4699;
	wire [4-1:0] node4700;
	wire [4-1:0] node4701;
	wire [4-1:0] node4702;
	wire [4-1:0] node4706;
	wire [4-1:0] node4709;
	wire [4-1:0] node4710;
	wire [4-1:0] node4711;
	wire [4-1:0] node4714;
	wire [4-1:0] node4717;
	wire [4-1:0] node4719;
	wire [4-1:0] node4722;
	wire [4-1:0] node4723;
	wire [4-1:0] node4724;
	wire [4-1:0] node4725;
	wire [4-1:0] node4728;
	wire [4-1:0] node4729;
	wire [4-1:0] node4732;
	wire [4-1:0] node4735;
	wire [4-1:0] node4736;
	wire [4-1:0] node4739;
	wire [4-1:0] node4741;
	wire [4-1:0] node4744;
	wire [4-1:0] node4745;
	wire [4-1:0] node4746;
	wire [4-1:0] node4747;
	wire [4-1:0] node4750;
	wire [4-1:0] node4753;
	wire [4-1:0] node4756;
	wire [4-1:0] node4757;
	wire [4-1:0] node4759;
	wire [4-1:0] node4762;
	wire [4-1:0] node4763;
	wire [4-1:0] node4767;
	wire [4-1:0] node4768;
	wire [4-1:0] node4769;
	wire [4-1:0] node4770;
	wire [4-1:0] node4771;
	wire [4-1:0] node4772;
	wire [4-1:0] node4774;
	wire [4-1:0] node4777;
	wire [4-1:0] node4779;
	wire [4-1:0] node4782;
	wire [4-1:0] node4783;
	wire [4-1:0] node4786;
	wire [4-1:0] node4787;
	wire [4-1:0] node4790;
	wire [4-1:0] node4793;
	wire [4-1:0] node4794;
	wire [4-1:0] node4795;
	wire [4-1:0] node4796;
	wire [4-1:0] node4800;
	wire [4-1:0] node4801;
	wire [4-1:0] node4805;
	wire [4-1:0] node4806;
	wire [4-1:0] node4808;
	wire [4-1:0] node4811;
	wire [4-1:0] node4814;
	wire [4-1:0] node4815;
	wire [4-1:0] node4816;
	wire [4-1:0] node4817;
	wire [4-1:0] node4820;
	wire [4-1:0] node4821;
	wire [4-1:0] node4824;
	wire [4-1:0] node4827;
	wire [4-1:0] node4828;
	wire [4-1:0] node4829;
	wire [4-1:0] node4833;
	wire [4-1:0] node4834;
	wire [4-1:0] node4837;
	wire [4-1:0] node4840;
	wire [4-1:0] node4841;
	wire [4-1:0] node4842;
	wire [4-1:0] node4843;
	wire [4-1:0] node4847;
	wire [4-1:0] node4850;
	wire [4-1:0] node4852;
	wire [4-1:0] node4854;
	wire [4-1:0] node4857;
	wire [4-1:0] node4858;
	wire [4-1:0] node4859;
	wire [4-1:0] node4860;
	wire [4-1:0] node4861;
	wire [4-1:0] node4862;
	wire [4-1:0] node4865;
	wire [4-1:0] node4868;
	wire [4-1:0] node4869;
	wire [4-1:0] node4873;
	wire [4-1:0] node4874;
	wire [4-1:0] node4877;
	wire [4-1:0] node4879;
	wire [4-1:0] node4882;
	wire [4-1:0] node4883;
	wire [4-1:0] node4885;
	wire [4-1:0] node4886;
	wire [4-1:0] node4889;
	wire [4-1:0] node4892;
	wire [4-1:0] node4893;
	wire [4-1:0] node4895;
	wire [4-1:0] node4898;
	wire [4-1:0] node4899;
	wire [4-1:0] node4902;
	wire [4-1:0] node4905;
	wire [4-1:0] node4906;
	wire [4-1:0] node4907;
	wire [4-1:0] node4908;
	wire [4-1:0] node4910;
	wire [4-1:0] node4913;
	wire [4-1:0] node4916;
	wire [4-1:0] node4917;
	wire [4-1:0] node4918;
	wire [4-1:0] node4921;
	wire [4-1:0] node4924;
	wire [4-1:0] node4925;
	wire [4-1:0] node4928;
	wire [4-1:0] node4931;
	wire [4-1:0] node4932;
	wire [4-1:0] node4933;
	wire [4-1:0] node4934;
	wire [4-1:0] node4937;
	wire [4-1:0] node4941;
	wire [4-1:0] node4942;
	wire [4-1:0] node4943;
	wire [4-1:0] node4947;
	wire [4-1:0] node4949;
	wire [4-1:0] node4952;
	wire [4-1:0] node4953;
	wire [4-1:0] node4954;
	wire [4-1:0] node4955;
	wire [4-1:0] node4956;
	wire [4-1:0] node4957;
	wire [4-1:0] node4958;
	wire [4-1:0] node4959;
	wire [4-1:0] node4960;
	wire [4-1:0] node4964;
	wire [4-1:0] node4967;
	wire [4-1:0] node4968;
	wire [4-1:0] node4970;
	wire [4-1:0] node4973;
	wire [4-1:0] node4974;
	wire [4-1:0] node4978;
	wire [4-1:0] node4979;
	wire [4-1:0] node4980;
	wire [4-1:0] node4981;
	wire [4-1:0] node4984;
	wire [4-1:0] node4987;
	wire [4-1:0] node4989;
	wire [4-1:0] node4992;
	wire [4-1:0] node4993;
	wire [4-1:0] node4996;
	wire [4-1:0] node4998;
	wire [4-1:0] node5001;
	wire [4-1:0] node5002;
	wire [4-1:0] node5003;
	wire [4-1:0] node5004;
	wire [4-1:0] node5006;
	wire [4-1:0] node5009;
	wire [4-1:0] node5012;
	wire [4-1:0] node5013;
	wire [4-1:0] node5014;
	wire [4-1:0] node5019;
	wire [4-1:0] node5020;
	wire [4-1:0] node5021;
	wire [4-1:0] node5023;
	wire [4-1:0] node5026;
	wire [4-1:0] node5027;
	wire [4-1:0] node5030;
	wire [4-1:0] node5033;
	wire [4-1:0] node5034;
	wire [4-1:0] node5035;
	wire [4-1:0] node5040;
	wire [4-1:0] node5041;
	wire [4-1:0] node5042;
	wire [4-1:0] node5043;
	wire [4-1:0] node5044;
	wire [4-1:0] node5045;
	wire [4-1:0] node5048;
	wire [4-1:0] node5051;
	wire [4-1:0] node5054;
	wire [4-1:0] node5055;
	wire [4-1:0] node5057;
	wire [4-1:0] node5060;
	wire [4-1:0] node5061;
	wire [4-1:0] node5065;
	wire [4-1:0] node5066;
	wire [4-1:0] node5067;
	wire [4-1:0] node5069;
	wire [4-1:0] node5072;
	wire [4-1:0] node5074;
	wire [4-1:0] node5077;
	wire [4-1:0] node5078;
	wire [4-1:0] node5081;
	wire [4-1:0] node5082;
	wire [4-1:0] node5086;
	wire [4-1:0] node5087;
	wire [4-1:0] node5088;
	wire [4-1:0] node5089;
	wire [4-1:0] node5091;
	wire [4-1:0] node5094;
	wire [4-1:0] node5095;
	wire [4-1:0] node5099;
	wire [4-1:0] node5100;
	wire [4-1:0] node5101;
	wire [4-1:0] node5105;
	wire [4-1:0] node5108;
	wire [4-1:0] node5109;
	wire [4-1:0] node5110;
	wire [4-1:0] node5114;
	wire [4-1:0] node5115;
	wire [4-1:0] node5116;
	wire [4-1:0] node5119;
	wire [4-1:0] node5122;
	wire [4-1:0] node5125;
	wire [4-1:0] node5126;
	wire [4-1:0] node5127;
	wire [4-1:0] node5128;
	wire [4-1:0] node5129;
	wire [4-1:0] node5130;
	wire [4-1:0] node5131;
	wire [4-1:0] node5135;
	wire [4-1:0] node5137;
	wire [4-1:0] node5140;
	wire [4-1:0] node5141;
	wire [4-1:0] node5143;
	wire [4-1:0] node5146;
	wire [4-1:0] node5149;
	wire [4-1:0] node5150;
	wire [4-1:0] node5152;
	wire [4-1:0] node5153;
	wire [4-1:0] node5157;
	wire [4-1:0] node5159;
	wire [4-1:0] node5162;
	wire [4-1:0] node5163;
	wire [4-1:0] node5164;
	wire [4-1:0] node5165;
	wire [4-1:0] node5168;
	wire [4-1:0] node5170;
	wire [4-1:0] node5173;
	wire [4-1:0] node5174;
	wire [4-1:0] node5175;
	wire [4-1:0] node5179;
	wire [4-1:0] node5180;
	wire [4-1:0] node5183;
	wire [4-1:0] node5186;
	wire [4-1:0] node5187;
	wire [4-1:0] node5188;
	wire [4-1:0] node5189;
	wire [4-1:0] node5193;
	wire [4-1:0] node5194;
	wire [4-1:0] node5198;
	wire [4-1:0] node5200;
	wire [4-1:0] node5202;
	wire [4-1:0] node5205;
	wire [4-1:0] node5206;
	wire [4-1:0] node5207;
	wire [4-1:0] node5208;
	wire [4-1:0] node5209;
	wire [4-1:0] node5210;
	wire [4-1:0] node5214;
	wire [4-1:0] node5216;
	wire [4-1:0] node5219;
	wire [4-1:0] node5220;
	wire [4-1:0] node5223;
	wire [4-1:0] node5224;
	wire [4-1:0] node5228;
	wire [4-1:0] node5229;
	wire [4-1:0] node5230;
	wire [4-1:0] node5231;
	wire [4-1:0] node5235;
	wire [4-1:0] node5236;
	wire [4-1:0] node5239;
	wire [4-1:0] node5242;
	wire [4-1:0] node5243;
	wire [4-1:0] node5244;
	wire [4-1:0] node5248;
	wire [4-1:0] node5249;
	wire [4-1:0] node5252;
	wire [4-1:0] node5255;
	wire [4-1:0] node5256;
	wire [4-1:0] node5257;
	wire [4-1:0] node5258;
	wire [4-1:0] node5261;
	wire [4-1:0] node5263;
	wire [4-1:0] node5266;
	wire [4-1:0] node5267;
	wire [4-1:0] node5268;
	wire [4-1:0] node5271;
	wire [4-1:0] node5275;
	wire [4-1:0] node5276;
	wire [4-1:0] node5277;
	wire [4-1:0] node5280;
	wire [4-1:0] node5281;
	wire [4-1:0] node5284;
	wire [4-1:0] node5287;
	wire [4-1:0] node5288;
	wire [4-1:0] node5291;
	wire [4-1:0] node5293;
	wire [4-1:0] node5296;
	wire [4-1:0] node5297;
	wire [4-1:0] node5298;
	wire [4-1:0] node5299;
	wire [4-1:0] node5300;
	wire [4-1:0] node5301;
	wire [4-1:0] node5302;
	wire [4-1:0] node5304;
	wire [4-1:0] node5307;
	wire [4-1:0] node5308;
	wire [4-1:0] node5311;
	wire [4-1:0] node5314;
	wire [4-1:0] node5315;
	wire [4-1:0] node5316;
	wire [4-1:0] node5319;
	wire [4-1:0] node5322;
	wire [4-1:0] node5323;
	wire [4-1:0] node5327;
	wire [4-1:0] node5328;
	wire [4-1:0] node5329;
	wire [4-1:0] node5330;
	wire [4-1:0] node5333;
	wire [4-1:0] node5336;
	wire [4-1:0] node5337;
	wire [4-1:0] node5341;
	wire [4-1:0] node5343;
	wire [4-1:0] node5344;
	wire [4-1:0] node5348;
	wire [4-1:0] node5349;
	wire [4-1:0] node5350;
	wire [4-1:0] node5351;
	wire [4-1:0] node5352;
	wire [4-1:0] node5356;
	wire [4-1:0] node5358;
	wire [4-1:0] node5361;
	wire [4-1:0] node5362;
	wire [4-1:0] node5365;
	wire [4-1:0] node5366;
	wire [4-1:0] node5370;
	wire [4-1:0] node5371;
	wire [4-1:0] node5373;
	wire [4-1:0] node5375;
	wire [4-1:0] node5378;
	wire [4-1:0] node5379;
	wire [4-1:0] node5383;
	wire [4-1:0] node5384;
	wire [4-1:0] node5385;
	wire [4-1:0] node5386;
	wire [4-1:0] node5387;
	wire [4-1:0] node5388;
	wire [4-1:0] node5391;
	wire [4-1:0] node5394;
	wire [4-1:0] node5396;
	wire [4-1:0] node5399;
	wire [4-1:0] node5400;
	wire [4-1:0] node5401;
	wire [4-1:0] node5405;
	wire [4-1:0] node5408;
	wire [4-1:0] node5409;
	wire [4-1:0] node5411;
	wire [4-1:0] node5412;
	wire [4-1:0] node5415;
	wire [4-1:0] node5418;
	wire [4-1:0] node5419;
	wire [4-1:0] node5420;
	wire [4-1:0] node5423;
	wire [4-1:0] node5426;
	wire [4-1:0] node5428;
	wire [4-1:0] node5431;
	wire [4-1:0] node5432;
	wire [4-1:0] node5433;
	wire [4-1:0] node5434;
	wire [4-1:0] node5435;
	wire [4-1:0] node5438;
	wire [4-1:0] node5441;
	wire [4-1:0] node5442;
	wire [4-1:0] node5445;
	wire [4-1:0] node5448;
	wire [4-1:0] node5449;
	wire [4-1:0] node5451;
	wire [4-1:0] node5454;
	wire [4-1:0] node5455;
	wire [4-1:0] node5459;
	wire [4-1:0] node5460;
	wire [4-1:0] node5461;
	wire [4-1:0] node5464;
	wire [4-1:0] node5465;
	wire [4-1:0] node5469;
	wire [4-1:0] node5471;
	wire [4-1:0] node5474;
	wire [4-1:0] node5475;
	wire [4-1:0] node5476;
	wire [4-1:0] node5477;
	wire [4-1:0] node5478;
	wire [4-1:0] node5479;
	wire [4-1:0] node5481;
	wire [4-1:0] node5484;
	wire [4-1:0] node5486;
	wire [4-1:0] node5489;
	wire [4-1:0] node5490;
	wire [4-1:0] node5491;
	wire [4-1:0] node5494;
	wire [4-1:0] node5497;
	wire [4-1:0] node5498;
	wire [4-1:0] node5502;
	wire [4-1:0] node5503;
	wire [4-1:0] node5504;
	wire [4-1:0] node5506;
	wire [4-1:0] node5509;
	wire [4-1:0] node5511;
	wire [4-1:0] node5514;
	wire [4-1:0] node5515;
	wire [4-1:0] node5516;
	wire [4-1:0] node5520;
	wire [4-1:0] node5522;
	wire [4-1:0] node5525;
	wire [4-1:0] node5526;
	wire [4-1:0] node5527;
	wire [4-1:0] node5528;
	wire [4-1:0] node5530;
	wire [4-1:0] node5533;
	wire [4-1:0] node5535;
	wire [4-1:0] node5538;
	wire [4-1:0] node5539;
	wire [4-1:0] node5541;
	wire [4-1:0] node5544;
	wire [4-1:0] node5546;
	wire [4-1:0] node5549;
	wire [4-1:0] node5550;
	wire [4-1:0] node5551;
	wire [4-1:0] node5552;
	wire [4-1:0] node5556;
	wire [4-1:0] node5559;
	wire [4-1:0] node5560;
	wire [4-1:0] node5562;
	wire [4-1:0] node5565;
	wire [4-1:0] node5567;
	wire [4-1:0] node5570;
	wire [4-1:0] node5571;
	wire [4-1:0] node5572;
	wire [4-1:0] node5573;
	wire [4-1:0] node5574;
	wire [4-1:0] node5575;
	wire [4-1:0] node5579;
	wire [4-1:0] node5581;
	wire [4-1:0] node5584;
	wire [4-1:0] node5585;
	wire [4-1:0] node5588;
	wire [4-1:0] node5589;
	wire [4-1:0] node5592;
	wire [4-1:0] node5595;
	wire [4-1:0] node5596;
	wire [4-1:0] node5597;
	wire [4-1:0] node5598;
	wire [4-1:0] node5601;
	wire [4-1:0] node5604;
	wire [4-1:0] node5607;
	wire [4-1:0] node5609;
	wire [4-1:0] node5610;
	wire [4-1:0] node5614;
	wire [4-1:0] node5615;
	wire [4-1:0] node5616;
	wire [4-1:0] node5617;
	wire [4-1:0] node5620;
	wire [4-1:0] node5621;
	wire [4-1:0] node5625;
	wire [4-1:0] node5626;
	wire [4-1:0] node5627;
	wire [4-1:0] node5630;
	wire [4-1:0] node5633;
	wire [4-1:0] node5636;
	wire [4-1:0] node5637;
	wire [4-1:0] node5638;
	wire [4-1:0] node5641;
	wire [4-1:0] node5642;
	wire [4-1:0] node5645;
	wire [4-1:0] node5648;
	wire [4-1:0] node5650;
	wire [4-1:0] node5653;
	wire [4-1:0] node5654;
	wire [4-1:0] node5655;
	wire [4-1:0] node5656;
	wire [4-1:0] node5657;
	wire [4-1:0] node5658;
	wire [4-1:0] node5659;
	wire [4-1:0] node5660;
	wire [4-1:0] node5661;
	wire [4-1:0] node5662;
	wire [4-1:0] node5663;
	wire [4-1:0] node5664;
	wire [4-1:0] node5667;
	wire [4-1:0] node5670;
	wire [4-1:0] node5671;
	wire [4-1:0] node5674;
	wire [4-1:0] node5677;
	wire [4-1:0] node5678;
	wire [4-1:0] node5679;
	wire [4-1:0] node5682;
	wire [4-1:0] node5685;
	wire [4-1:0] node5687;
	wire [4-1:0] node5690;
	wire [4-1:0] node5691;
	wire [4-1:0] node5692;
	wire [4-1:0] node5693;
	wire [4-1:0] node5696;
	wire [4-1:0] node5699;
	wire [4-1:0] node5701;
	wire [4-1:0] node5704;
	wire [4-1:0] node5707;
	wire [4-1:0] node5708;
	wire [4-1:0] node5709;
	wire [4-1:0] node5710;
	wire [4-1:0] node5712;
	wire [4-1:0] node5716;
	wire [4-1:0] node5717;
	wire [4-1:0] node5719;
	wire [4-1:0] node5722;
	wire [4-1:0] node5725;
	wire [4-1:0] node5726;
	wire [4-1:0] node5727;
	wire [4-1:0] node5728;
	wire [4-1:0] node5731;
	wire [4-1:0] node5735;
	wire [4-1:0] node5736;
	wire [4-1:0] node5737;
	wire [4-1:0] node5740;
	wire [4-1:0] node5744;
	wire [4-1:0] node5745;
	wire [4-1:0] node5746;
	wire [4-1:0] node5747;
	wire [4-1:0] node5748;
	wire [4-1:0] node5749;
	wire [4-1:0] node5753;
	wire [4-1:0] node5756;
	wire [4-1:0] node5757;
	wire [4-1:0] node5758;
	wire [4-1:0] node5761;
	wire [4-1:0] node5764;
	wire [4-1:0] node5765;
	wire [4-1:0] node5769;
	wire [4-1:0] node5770;
	wire [4-1:0] node5771;
	wire [4-1:0] node5773;
	wire [4-1:0] node5776;
	wire [4-1:0] node5777;
	wire [4-1:0] node5781;
	wire [4-1:0] node5782;
	wire [4-1:0] node5785;
	wire [4-1:0] node5786;
	wire [4-1:0] node5789;
	wire [4-1:0] node5792;
	wire [4-1:0] node5793;
	wire [4-1:0] node5794;
	wire [4-1:0] node5795;
	wire [4-1:0] node5797;
	wire [4-1:0] node5800;
	wire [4-1:0] node5803;
	wire [4-1:0] node5804;
	wire [4-1:0] node5805;
	wire [4-1:0] node5809;
	wire [4-1:0] node5810;
	wire [4-1:0] node5814;
	wire [4-1:0] node5815;
	wire [4-1:0] node5816;
	wire [4-1:0] node5819;
	wire [4-1:0] node5820;
	wire [4-1:0] node5823;
	wire [4-1:0] node5826;
	wire [4-1:0] node5827;
	wire [4-1:0] node5831;
	wire [4-1:0] node5832;
	wire [4-1:0] node5833;
	wire [4-1:0] node5834;
	wire [4-1:0] node5835;
	wire [4-1:0] node5836;
	wire [4-1:0] node5837;
	wire [4-1:0] node5840;
	wire [4-1:0] node5843;
	wire [4-1:0] node5844;
	wire [4-1:0] node5847;
	wire [4-1:0] node5850;
	wire [4-1:0] node5851;
	wire [4-1:0] node5852;
	wire [4-1:0] node5856;
	wire [4-1:0] node5857;
	wire [4-1:0] node5860;
	wire [4-1:0] node5863;
	wire [4-1:0] node5864;
	wire [4-1:0] node5865;
	wire [4-1:0] node5868;
	wire [4-1:0] node5869;
	wire [4-1:0] node5872;
	wire [4-1:0] node5875;
	wire [4-1:0] node5876;
	wire [4-1:0] node5878;
	wire [4-1:0] node5881;
	wire [4-1:0] node5882;
	wire [4-1:0] node5885;
	wire [4-1:0] node5888;
	wire [4-1:0] node5889;
	wire [4-1:0] node5890;
	wire [4-1:0] node5891;
	wire [4-1:0] node5892;
	wire [4-1:0] node5896;
	wire [4-1:0] node5898;
	wire [4-1:0] node5901;
	wire [4-1:0] node5902;
	wire [4-1:0] node5903;
	wire [4-1:0] node5907;
	wire [4-1:0] node5910;
	wire [4-1:0] node5911;
	wire [4-1:0] node5914;
	wire [4-1:0] node5915;
	wire [4-1:0] node5917;
	wire [4-1:0] node5920;
	wire [4-1:0] node5923;
	wire [4-1:0] node5924;
	wire [4-1:0] node5925;
	wire [4-1:0] node5926;
	wire [4-1:0] node5927;
	wire [4-1:0] node5929;
	wire [4-1:0] node5932;
	wire [4-1:0] node5935;
	wire [4-1:0] node5936;
	wire [4-1:0] node5937;
	wire [4-1:0] node5940;
	wire [4-1:0] node5943;
	wire [4-1:0] node5944;
	wire [4-1:0] node5948;
	wire [4-1:0] node5949;
	wire [4-1:0] node5951;
	wire [4-1:0] node5952;
	wire [4-1:0] node5956;
	wire [4-1:0] node5958;
	wire [4-1:0] node5959;
	wire [4-1:0] node5962;
	wire [4-1:0] node5965;
	wire [4-1:0] node5966;
	wire [4-1:0] node5967;
	wire [4-1:0] node5968;
	wire [4-1:0] node5969;
	wire [4-1:0] node5973;
	wire [4-1:0] node5974;
	wire [4-1:0] node5977;
	wire [4-1:0] node5980;
	wire [4-1:0] node5981;
	wire [4-1:0] node5982;
	wire [4-1:0] node5986;
	wire [4-1:0] node5987;
	wire [4-1:0] node5990;
	wire [4-1:0] node5993;
	wire [4-1:0] node5994;
	wire [4-1:0] node5996;
	wire [4-1:0] node5997;
	wire [4-1:0] node6001;
	wire [4-1:0] node6002;
	wire [4-1:0] node6004;
	wire [4-1:0] node6007;
	wire [4-1:0] node6008;
	wire [4-1:0] node6012;
	wire [4-1:0] node6013;
	wire [4-1:0] node6014;
	wire [4-1:0] node6015;
	wire [4-1:0] node6016;
	wire [4-1:0] node6017;
	wire [4-1:0] node6019;
	wire [4-1:0] node6020;
	wire [4-1:0] node6023;
	wire [4-1:0] node6026;
	wire [4-1:0] node6027;
	wire [4-1:0] node6031;
	wire [4-1:0] node6032;
	wire [4-1:0] node6033;
	wire [4-1:0] node6034;
	wire [4-1:0] node6038;
	wire [4-1:0] node6040;
	wire [4-1:0] node6043;
	wire [4-1:0] node6044;
	wire [4-1:0] node6046;
	wire [4-1:0] node6049;
	wire [4-1:0] node6050;
	wire [4-1:0] node6054;
	wire [4-1:0] node6055;
	wire [4-1:0] node6056;
	wire [4-1:0] node6057;
	wire [4-1:0] node6059;
	wire [4-1:0] node6062;
	wire [4-1:0] node6065;
	wire [4-1:0] node6066;
	wire [4-1:0] node6067;
	wire [4-1:0] node6071;
	wire [4-1:0] node6072;
	wire [4-1:0] node6076;
	wire [4-1:0] node6077;
	wire [4-1:0] node6078;
	wire [4-1:0] node6079;
	wire [4-1:0] node6083;
	wire [4-1:0] node6086;
	wire [4-1:0] node6087;
	wire [4-1:0] node6089;
	wire [4-1:0] node6092;
	wire [4-1:0] node6094;
	wire [4-1:0] node6097;
	wire [4-1:0] node6098;
	wire [4-1:0] node6099;
	wire [4-1:0] node6100;
	wire [4-1:0] node6101;
	wire [4-1:0] node6105;
	wire [4-1:0] node6106;
	wire [4-1:0] node6108;
	wire [4-1:0] node6111;
	wire [4-1:0] node6112;
	wire [4-1:0] node6116;
	wire [4-1:0] node6117;
	wire [4-1:0] node6118;
	wire [4-1:0] node6119;
	wire [4-1:0] node6123;
	wire [4-1:0] node6124;
	wire [4-1:0] node6128;
	wire [4-1:0] node6129;
	wire [4-1:0] node6133;
	wire [4-1:0] node6134;
	wire [4-1:0] node6135;
	wire [4-1:0] node6136;
	wire [4-1:0] node6139;
	wire [4-1:0] node6142;
	wire [4-1:0] node6143;
	wire [4-1:0] node6145;
	wire [4-1:0] node6148;
	wire [4-1:0] node6151;
	wire [4-1:0] node6152;
	wire [4-1:0] node6154;
	wire [4-1:0] node6156;
	wire [4-1:0] node6159;
	wire [4-1:0] node6160;
	wire [4-1:0] node6162;
	wire [4-1:0] node6165;
	wire [4-1:0] node6166;
	wire [4-1:0] node6170;
	wire [4-1:0] node6171;
	wire [4-1:0] node6172;
	wire [4-1:0] node6173;
	wire [4-1:0] node6174;
	wire [4-1:0] node6175;
	wire [4-1:0] node6176;
	wire [4-1:0] node6180;
	wire [4-1:0] node6183;
	wire [4-1:0] node6184;
	wire [4-1:0] node6186;
	wire [4-1:0] node6189;
	wire [4-1:0] node6190;
	wire [4-1:0] node6194;
	wire [4-1:0] node6195;
	wire [4-1:0] node6196;
	wire [4-1:0] node6198;
	wire [4-1:0] node6201;
	wire [4-1:0] node6204;
	wire [4-1:0] node6205;
	wire [4-1:0] node6208;
	wire [4-1:0] node6210;
	wire [4-1:0] node6213;
	wire [4-1:0] node6214;
	wire [4-1:0] node6215;
	wire [4-1:0] node6216;
	wire [4-1:0] node6218;
	wire [4-1:0] node6221;
	wire [4-1:0] node6223;
	wire [4-1:0] node6226;
	wire [4-1:0] node6227;
	wire [4-1:0] node6228;
	wire [4-1:0] node6231;
	wire [4-1:0] node6234;
	wire [4-1:0] node6236;
	wire [4-1:0] node6239;
	wire [4-1:0] node6240;
	wire [4-1:0] node6241;
	wire [4-1:0] node6244;
	wire [4-1:0] node6245;
	wire [4-1:0] node6248;
	wire [4-1:0] node6251;
	wire [4-1:0] node6252;
	wire [4-1:0] node6254;
	wire [4-1:0] node6257;
	wire [4-1:0] node6260;
	wire [4-1:0] node6261;
	wire [4-1:0] node6262;
	wire [4-1:0] node6263;
	wire [4-1:0] node6264;
	wire [4-1:0] node6265;
	wire [4-1:0] node6269;
	wire [4-1:0] node6270;
	wire [4-1:0] node6273;
	wire [4-1:0] node6276;
	wire [4-1:0] node6277;
	wire [4-1:0] node6278;
	wire [4-1:0] node6281;
	wire [4-1:0] node6285;
	wire [4-1:0] node6286;
	wire [4-1:0] node6287;
	wire [4-1:0] node6288;
	wire [4-1:0] node6291;
	wire [4-1:0] node6294;
	wire [4-1:0] node6296;
	wire [4-1:0] node6299;
	wire [4-1:0] node6300;
	wire [4-1:0] node6302;
	wire [4-1:0] node6305;
	wire [4-1:0] node6306;
	wire [4-1:0] node6310;
	wire [4-1:0] node6311;
	wire [4-1:0] node6312;
	wire [4-1:0] node6313;
	wire [4-1:0] node6314;
	wire [4-1:0] node6317;
	wire [4-1:0] node6320;
	wire [4-1:0] node6321;
	wire [4-1:0] node6325;
	wire [4-1:0] node6327;
	wire [4-1:0] node6328;
	wire [4-1:0] node6331;
	wire [4-1:0] node6334;
	wire [4-1:0] node6335;
	wire [4-1:0] node6336;
	wire [4-1:0] node6337;
	wire [4-1:0] node6340;
	wire [4-1:0] node6343;
	wire [4-1:0] node6345;
	wire [4-1:0] node6348;
	wire [4-1:0] node6350;
	wire [4-1:0] node6351;
	wire [4-1:0] node6354;
	wire [4-1:0] node6357;
	wire [4-1:0] node6358;
	wire [4-1:0] node6359;
	wire [4-1:0] node6360;
	wire [4-1:0] node6361;
	wire [4-1:0] node6362;
	wire [4-1:0] node6363;
	wire [4-1:0] node6365;
	wire [4-1:0] node6366;
	wire [4-1:0] node6369;
	wire [4-1:0] node6372;
	wire [4-1:0] node6375;
	wire [4-1:0] node6376;
	wire [4-1:0] node6377;
	wire [4-1:0] node6378;
	wire [4-1:0] node6382;
	wire [4-1:0] node6383;
	wire [4-1:0] node6387;
	wire [4-1:0] node6388;
	wire [4-1:0] node6389;
	wire [4-1:0] node6393;
	wire [4-1:0] node6394;
	wire [4-1:0] node6397;
	wire [4-1:0] node6400;
	wire [4-1:0] node6401;
	wire [4-1:0] node6402;
	wire [4-1:0] node6403;
	wire [4-1:0] node6405;
	wire [4-1:0] node6408;
	wire [4-1:0] node6410;
	wire [4-1:0] node6413;
	wire [4-1:0] node6414;
	wire [4-1:0] node6415;
	wire [4-1:0] node6418;
	wire [4-1:0] node6422;
	wire [4-1:0] node6423;
	wire [4-1:0] node6424;
	wire [4-1:0] node6425;
	wire [4-1:0] node6429;
	wire [4-1:0] node6430;
	wire [4-1:0] node6434;
	wire [4-1:0] node6435;
	wire [4-1:0] node6437;
	wire [4-1:0] node6441;
	wire [4-1:0] node6442;
	wire [4-1:0] node6443;
	wire [4-1:0] node6444;
	wire [4-1:0] node6445;
	wire [4-1:0] node6447;
	wire [4-1:0] node6450;
	wire [4-1:0] node6453;
	wire [4-1:0] node6454;
	wire [4-1:0] node6455;
	wire [4-1:0] node6458;
	wire [4-1:0] node6461;
	wire [4-1:0] node6463;
	wire [4-1:0] node6466;
	wire [4-1:0] node6467;
	wire [4-1:0] node6468;
	wire [4-1:0] node6469;
	wire [4-1:0] node6473;
	wire [4-1:0] node6474;
	wire [4-1:0] node6477;
	wire [4-1:0] node6480;
	wire [4-1:0] node6481;
	wire [4-1:0] node6482;
	wire [4-1:0] node6485;
	wire [4-1:0] node6489;
	wire [4-1:0] node6490;
	wire [4-1:0] node6491;
	wire [4-1:0] node6492;
	wire [4-1:0] node6493;
	wire [4-1:0] node6496;
	wire [4-1:0] node6500;
	wire [4-1:0] node6501;
	wire [4-1:0] node6503;
	wire [4-1:0] node6506;
	wire [4-1:0] node6509;
	wire [4-1:0] node6510;
	wire [4-1:0] node6511;
	wire [4-1:0] node6512;
	wire [4-1:0] node6515;
	wire [4-1:0] node6519;
	wire [4-1:0] node6521;
	wire [4-1:0] node6523;
	wire [4-1:0] node6526;
	wire [4-1:0] node6527;
	wire [4-1:0] node6528;
	wire [4-1:0] node6529;
	wire [4-1:0] node6530;
	wire [4-1:0] node6531;
	wire [4-1:0] node6532;
	wire [4-1:0] node6535;
	wire [4-1:0] node6538;
	wire [4-1:0] node6539;
	wire [4-1:0] node6542;
	wire [4-1:0] node6545;
	wire [4-1:0] node6546;
	wire [4-1:0] node6547;
	wire [4-1:0] node6550;
	wire [4-1:0] node6553;
	wire [4-1:0] node6555;
	wire [4-1:0] node6558;
	wire [4-1:0] node6559;
	wire [4-1:0] node6560;
	wire [4-1:0] node6561;
	wire [4-1:0] node6564;
	wire [4-1:0] node6567;
	wire [4-1:0] node6568;
	wire [4-1:0] node6572;
	wire [4-1:0] node6574;
	wire [4-1:0] node6576;
	wire [4-1:0] node6579;
	wire [4-1:0] node6580;
	wire [4-1:0] node6581;
	wire [4-1:0] node6582;
	wire [4-1:0] node6584;
	wire [4-1:0] node6587;
	wire [4-1:0] node6589;
	wire [4-1:0] node6592;
	wire [4-1:0] node6594;
	wire [4-1:0] node6597;
	wire [4-1:0] node6598;
	wire [4-1:0] node6599;
	wire [4-1:0] node6601;
	wire [4-1:0] node6604;
	wire [4-1:0] node6607;
	wire [4-1:0] node6608;
	wire [4-1:0] node6610;
	wire [4-1:0] node6613;
	wire [4-1:0] node6615;
	wire [4-1:0] node6618;
	wire [4-1:0] node6619;
	wire [4-1:0] node6620;
	wire [4-1:0] node6621;
	wire [4-1:0] node6624;
	wire [4-1:0] node6625;
	wire [4-1:0] node6626;
	wire [4-1:0] node6629;
	wire [4-1:0] node6632;
	wire [4-1:0] node6633;
	wire [4-1:0] node6636;
	wire [4-1:0] node6639;
	wire [4-1:0] node6640;
	wire [4-1:0] node6641;
	wire [4-1:0] node6642;
	wire [4-1:0] node6646;
	wire [4-1:0] node6649;
	wire [4-1:0] node6650;
	wire [4-1:0] node6652;
	wire [4-1:0] node6656;
	wire [4-1:0] node6657;
	wire [4-1:0] node6658;
	wire [4-1:0] node6659;
	wire [4-1:0] node6662;
	wire [4-1:0] node6665;
	wire [4-1:0] node6666;
	wire [4-1:0] node6668;
	wire [4-1:0] node6671;
	wire [4-1:0] node6672;
	wire [4-1:0] node6675;
	wire [4-1:0] node6678;
	wire [4-1:0] node6679;
	wire [4-1:0] node6680;
	wire [4-1:0] node6682;
	wire [4-1:0] node6685;
	wire [4-1:0] node6686;
	wire [4-1:0] node6690;
	wire [4-1:0] node6691;
	wire [4-1:0] node6692;
	wire [4-1:0] node6696;
	wire [4-1:0] node6697;
	wire [4-1:0] node6701;
	wire [4-1:0] node6702;
	wire [4-1:0] node6703;
	wire [4-1:0] node6704;
	wire [4-1:0] node6705;
	wire [4-1:0] node6706;
	wire [4-1:0] node6707;
	wire [4-1:0] node6710;
	wire [4-1:0] node6712;
	wire [4-1:0] node6715;
	wire [4-1:0] node6716;
	wire [4-1:0] node6717;
	wire [4-1:0] node6720;
	wire [4-1:0] node6723;
	wire [4-1:0] node6724;
	wire [4-1:0] node6728;
	wire [4-1:0] node6729;
	wire [4-1:0] node6730;
	wire [4-1:0] node6731;
	wire [4-1:0] node6734;
	wire [4-1:0] node6737;
	wire [4-1:0] node6738;
	wire [4-1:0] node6742;
	wire [4-1:0] node6743;
	wire [4-1:0] node6745;
	wire [4-1:0] node6748;
	wire [4-1:0] node6751;
	wire [4-1:0] node6752;
	wire [4-1:0] node6753;
	wire [4-1:0] node6754;
	wire [4-1:0] node6755;
	wire [4-1:0] node6758;
	wire [4-1:0] node6761;
	wire [4-1:0] node6763;
	wire [4-1:0] node6766;
	wire [4-1:0] node6767;
	wire [4-1:0] node6768;
	wire [4-1:0] node6772;
	wire [4-1:0] node6773;
	wire [4-1:0] node6776;
	wire [4-1:0] node6779;
	wire [4-1:0] node6780;
	wire [4-1:0] node6781;
	wire [4-1:0] node6784;
	wire [4-1:0] node6786;
	wire [4-1:0] node6789;
	wire [4-1:0] node6790;
	wire [4-1:0] node6794;
	wire [4-1:0] node6795;
	wire [4-1:0] node6796;
	wire [4-1:0] node6797;
	wire [4-1:0] node6798;
	wire [4-1:0] node6799;
	wire [4-1:0] node6803;
	wire [4-1:0] node6804;
	wire [4-1:0] node6807;
	wire [4-1:0] node6810;
	wire [4-1:0] node6811;
	wire [4-1:0] node6812;
	wire [4-1:0] node6815;
	wire [4-1:0] node6819;
	wire [4-1:0] node6820;
	wire [4-1:0] node6821;
	wire [4-1:0] node6823;
	wire [4-1:0] node6826;
	wire [4-1:0] node6827;
	wire [4-1:0] node6830;
	wire [4-1:0] node6833;
	wire [4-1:0] node6834;
	wire [4-1:0] node6835;
	wire [4-1:0] node6839;
	wire [4-1:0] node6842;
	wire [4-1:0] node6843;
	wire [4-1:0] node6844;
	wire [4-1:0] node6846;
	wire [4-1:0] node6849;
	wire [4-1:0] node6850;
	wire [4-1:0] node6851;
	wire [4-1:0] node6854;
	wire [4-1:0] node6857;
	wire [4-1:0] node6858;
	wire [4-1:0] node6862;
	wire [4-1:0] node6863;
	wire [4-1:0] node6864;
	wire [4-1:0] node6865;
	wire [4-1:0] node6869;
	wire [4-1:0] node6870;
	wire [4-1:0] node6874;
	wire [4-1:0] node6875;
	wire [4-1:0] node6876;
	wire [4-1:0] node6879;
	wire [4-1:0] node6882;
	wire [4-1:0] node6883;
	wire [4-1:0] node6886;
	wire [4-1:0] node6889;
	wire [4-1:0] node6890;
	wire [4-1:0] node6891;
	wire [4-1:0] node6892;
	wire [4-1:0] node6893;
	wire [4-1:0] node6894;
	wire [4-1:0] node6896;
	wire [4-1:0] node6899;
	wire [4-1:0] node6900;
	wire [4-1:0] node6903;
	wire [4-1:0] node6906;
	wire [4-1:0] node6908;
	wire [4-1:0] node6909;
	wire [4-1:0] node6913;
	wire [4-1:0] node6914;
	wire [4-1:0] node6915;
	wire [4-1:0] node6918;
	wire [4-1:0] node6920;
	wire [4-1:0] node6923;
	wire [4-1:0] node6924;
	wire [4-1:0] node6925;
	wire [4-1:0] node6928;
	wire [4-1:0] node6931;
	wire [4-1:0] node6934;
	wire [4-1:0] node6935;
	wire [4-1:0] node6936;
	wire [4-1:0] node6937;
	wire [4-1:0] node6940;
	wire [4-1:0] node6941;
	wire [4-1:0] node6945;
	wire [4-1:0] node6946;
	wire [4-1:0] node6947;
	wire [4-1:0] node6951;
	wire [4-1:0] node6952;
	wire [4-1:0] node6955;
	wire [4-1:0] node6958;
	wire [4-1:0] node6959;
	wire [4-1:0] node6960;
	wire [4-1:0] node6962;
	wire [4-1:0] node6965;
	wire [4-1:0] node6968;
	wire [4-1:0] node6970;
	wire [4-1:0] node6971;
	wire [4-1:0] node6975;
	wire [4-1:0] node6976;
	wire [4-1:0] node6977;
	wire [4-1:0] node6978;
	wire [4-1:0] node6979;
	wire [4-1:0] node6980;
	wire [4-1:0] node6983;
	wire [4-1:0] node6986;
	wire [4-1:0] node6987;
	wire [4-1:0] node6990;
	wire [4-1:0] node6993;
	wire [4-1:0] node6994;
	wire [4-1:0] node6996;
	wire [4-1:0] node6999;
	wire [4-1:0] node7000;
	wire [4-1:0] node7003;
	wire [4-1:0] node7006;
	wire [4-1:0] node7007;
	wire [4-1:0] node7008;
	wire [4-1:0] node7009;
	wire [4-1:0] node7013;
	wire [4-1:0] node7016;
	wire [4-1:0] node7017;
	wire [4-1:0] node7018;
	wire [4-1:0] node7022;
	wire [4-1:0] node7023;
	wire [4-1:0] node7026;
	wire [4-1:0] node7029;
	wire [4-1:0] node7030;
	wire [4-1:0] node7031;
	wire [4-1:0] node7032;
	wire [4-1:0] node7033;
	wire [4-1:0] node7036;
	wire [4-1:0] node7040;
	wire [4-1:0] node7041;
	wire [4-1:0] node7042;
	wire [4-1:0] node7046;
	wire [4-1:0] node7049;
	wire [4-1:0] node7050;
	wire [4-1:0] node7051;
	wire [4-1:0] node7054;
	wire [4-1:0] node7056;
	wire [4-1:0] node7059;
	wire [4-1:0] node7060;
	wire [4-1:0] node7061;
	wire [4-1:0] node7065;
	wire [4-1:0] node7067;
	wire [4-1:0] node7070;
	wire [4-1:0] node7071;
	wire [4-1:0] node7072;
	wire [4-1:0] node7073;
	wire [4-1:0] node7074;
	wire [4-1:0] node7075;
	wire [4-1:0] node7076;
	wire [4-1:0] node7077;
	wire [4-1:0] node7078;
	wire [4-1:0] node7081;
	wire [4-1:0] node7084;
	wire [4-1:0] node7085;
	wire [4-1:0] node7086;
	wire [4-1:0] node7091;
	wire [4-1:0] node7092;
	wire [4-1:0] node7093;
	wire [4-1:0] node7094;
	wire [4-1:0] node7098;
	wire [4-1:0] node7099;
	wire [4-1:0] node7103;
	wire [4-1:0] node7104;
	wire [4-1:0] node7107;
	wire [4-1:0] node7110;
	wire [4-1:0] node7111;
	wire [4-1:0] node7112;
	wire [4-1:0] node7113;
	wire [4-1:0] node7116;
	wire [4-1:0] node7118;
	wire [4-1:0] node7121;
	wire [4-1:0] node7122;
	wire [4-1:0] node7123;
	wire [4-1:0] node7127;
	wire [4-1:0] node7129;
	wire [4-1:0] node7132;
	wire [4-1:0] node7133;
	wire [4-1:0] node7134;
	wire [4-1:0] node7136;
	wire [4-1:0] node7139;
	wire [4-1:0] node7141;
	wire [4-1:0] node7144;
	wire [4-1:0] node7145;
	wire [4-1:0] node7146;
	wire [4-1:0] node7149;
	wire [4-1:0] node7152;
	wire [4-1:0] node7154;
	wire [4-1:0] node7157;
	wire [4-1:0] node7158;
	wire [4-1:0] node7159;
	wire [4-1:0] node7160;
	wire [4-1:0] node7161;
	wire [4-1:0] node7162;
	wire [4-1:0] node7166;
	wire [4-1:0] node7168;
	wire [4-1:0] node7171;
	wire [4-1:0] node7172;
	wire [4-1:0] node7173;
	wire [4-1:0] node7176;
	wire [4-1:0] node7180;
	wire [4-1:0] node7181;
	wire [4-1:0] node7182;
	wire [4-1:0] node7183;
	wire [4-1:0] node7186;
	wire [4-1:0] node7189;
	wire [4-1:0] node7192;
	wire [4-1:0] node7193;
	wire [4-1:0] node7194;
	wire [4-1:0] node7197;
	wire [4-1:0] node7200;
	wire [4-1:0] node7202;
	wire [4-1:0] node7205;
	wire [4-1:0] node7206;
	wire [4-1:0] node7207;
	wire [4-1:0] node7208;
	wire [4-1:0] node7209;
	wire [4-1:0] node7212;
	wire [4-1:0] node7215;
	wire [4-1:0] node7216;
	wire [4-1:0] node7219;
	wire [4-1:0] node7222;
	wire [4-1:0] node7223;
	wire [4-1:0] node7227;
	wire [4-1:0] node7228;
	wire [4-1:0] node7229;
	wire [4-1:0] node7230;
	wire [4-1:0] node7233;
	wire [4-1:0] node7236;
	wire [4-1:0] node7239;
	wire [4-1:0] node7240;
	wire [4-1:0] node7241;
	wire [4-1:0] node7244;
	wire [4-1:0] node7248;
	wire [4-1:0] node7249;
	wire [4-1:0] node7250;
	wire [4-1:0] node7251;
	wire [4-1:0] node7252;
	wire [4-1:0] node7253;
	wire [4-1:0] node7254;
	wire [4-1:0] node7257;
	wire [4-1:0] node7260;
	wire [4-1:0] node7261;
	wire [4-1:0] node7264;
	wire [4-1:0] node7267;
	wire [4-1:0] node7268;
	wire [4-1:0] node7269;
	wire [4-1:0] node7272;
	wire [4-1:0] node7275;
	wire [4-1:0] node7278;
	wire [4-1:0] node7279;
	wire [4-1:0] node7280;
	wire [4-1:0] node7281;
	wire [4-1:0] node7285;
	wire [4-1:0] node7286;
	wire [4-1:0] node7290;
	wire [4-1:0] node7292;
	wire [4-1:0] node7295;
	wire [4-1:0] node7296;
	wire [4-1:0] node7297;
	wire [4-1:0] node7298;
	wire [4-1:0] node7299;
	wire [4-1:0] node7302;
	wire [4-1:0] node7306;
	wire [4-1:0] node7307;
	wire [4-1:0] node7308;
	wire [4-1:0] node7312;
	wire [4-1:0] node7313;
	wire [4-1:0] node7317;
	wire [4-1:0] node7318;
	wire [4-1:0] node7319;
	wire [4-1:0] node7320;
	wire [4-1:0] node7323;
	wire [4-1:0] node7326;
	wire [4-1:0] node7328;
	wire [4-1:0] node7331;
	wire [4-1:0] node7332;
	wire [4-1:0] node7334;
	wire [4-1:0] node7337;
	wire [4-1:0] node7338;
	wire [4-1:0] node7341;
	wire [4-1:0] node7344;
	wire [4-1:0] node7345;
	wire [4-1:0] node7346;
	wire [4-1:0] node7347;
	wire [4-1:0] node7348;
	wire [4-1:0] node7350;
	wire [4-1:0] node7353;
	wire [4-1:0] node7354;
	wire [4-1:0] node7358;
	wire [4-1:0] node7359;
	wire [4-1:0] node7360;
	wire [4-1:0] node7364;
	wire [4-1:0] node7365;
	wire [4-1:0] node7368;
	wire [4-1:0] node7371;
	wire [4-1:0] node7372;
	wire [4-1:0] node7373;
	wire [4-1:0] node7376;
	wire [4-1:0] node7379;
	wire [4-1:0] node7380;
	wire [4-1:0] node7382;
	wire [4-1:0] node7385;
	wire [4-1:0] node7387;
	wire [4-1:0] node7390;
	wire [4-1:0] node7391;
	wire [4-1:0] node7392;
	wire [4-1:0] node7393;
	wire [4-1:0] node7394;
	wire [4-1:0] node7397;
	wire [4-1:0] node7400;
	wire [4-1:0] node7402;
	wire [4-1:0] node7405;
	wire [4-1:0] node7406;
	wire [4-1:0] node7407;
	wire [4-1:0] node7411;
	wire [4-1:0] node7412;
	wire [4-1:0] node7416;
	wire [4-1:0] node7417;
	wire [4-1:0] node7418;
	wire [4-1:0] node7419;
	wire [4-1:0] node7423;
	wire [4-1:0] node7424;
	wire [4-1:0] node7427;
	wire [4-1:0] node7430;
	wire [4-1:0] node7431;
	wire [4-1:0] node7432;
	wire [4-1:0] node7435;
	wire [4-1:0] node7438;
	wire [4-1:0] node7441;
	wire [4-1:0] node7442;
	wire [4-1:0] node7443;
	wire [4-1:0] node7444;
	wire [4-1:0] node7445;
	wire [4-1:0] node7446;
	wire [4-1:0] node7447;
	wire [4-1:0] node7448;
	wire [4-1:0] node7451;
	wire [4-1:0] node7454;
	wire [4-1:0] node7455;
	wire [4-1:0] node7459;
	wire [4-1:0] node7460;
	wire [4-1:0] node7462;
	wire [4-1:0] node7465;
	wire [4-1:0] node7467;
	wire [4-1:0] node7470;
	wire [4-1:0] node7471;
	wire [4-1:0] node7472;
	wire [4-1:0] node7474;
	wire [4-1:0] node7477;
	wire [4-1:0] node7478;
	wire [4-1:0] node7481;
	wire [4-1:0] node7484;
	wire [4-1:0] node7485;
	wire [4-1:0] node7486;
	wire [4-1:0] node7490;
	wire [4-1:0] node7493;
	wire [4-1:0] node7494;
	wire [4-1:0] node7495;
	wire [4-1:0] node7496;
	wire [4-1:0] node7498;
	wire [4-1:0] node7501;
	wire [4-1:0] node7504;
	wire [4-1:0] node7505;
	wire [4-1:0] node7506;
	wire [4-1:0] node7509;
	wire [4-1:0] node7512;
	wire [4-1:0] node7513;
	wire [4-1:0] node7516;
	wire [4-1:0] node7519;
	wire [4-1:0] node7520;
	wire [4-1:0] node7522;
	wire [4-1:0] node7525;
	wire [4-1:0] node7526;
	wire [4-1:0] node7527;
	wire [4-1:0] node7531;
	wire [4-1:0] node7532;
	wire [4-1:0] node7535;
	wire [4-1:0] node7538;
	wire [4-1:0] node7539;
	wire [4-1:0] node7540;
	wire [4-1:0] node7541;
	wire [4-1:0] node7542;
	wire [4-1:0] node7544;
	wire [4-1:0] node7547;
	wire [4-1:0] node7549;
	wire [4-1:0] node7552;
	wire [4-1:0] node7553;
	wire [4-1:0] node7554;
	wire [4-1:0] node7557;
	wire [4-1:0] node7560;
	wire [4-1:0] node7562;
	wire [4-1:0] node7565;
	wire [4-1:0] node7566;
	wire [4-1:0] node7567;
	wire [4-1:0] node7568;
	wire [4-1:0] node7572;
	wire [4-1:0] node7574;
	wire [4-1:0] node7577;
	wire [4-1:0] node7578;
	wire [4-1:0] node7580;
	wire [4-1:0] node7583;
	wire [4-1:0] node7584;
	wire [4-1:0] node7587;
	wire [4-1:0] node7590;
	wire [4-1:0] node7591;
	wire [4-1:0] node7592;
	wire [4-1:0] node7593;
	wire [4-1:0] node7595;
	wire [4-1:0] node7598;
	wire [4-1:0] node7599;
	wire [4-1:0] node7603;
	wire [4-1:0] node7604;
	wire [4-1:0] node7605;
	wire [4-1:0] node7608;
	wire [4-1:0] node7611;
	wire [4-1:0] node7614;
	wire [4-1:0] node7615;
	wire [4-1:0] node7616;
	wire [4-1:0] node7618;
	wire [4-1:0] node7622;
	wire [4-1:0] node7623;
	wire [4-1:0] node7626;
	wire [4-1:0] node7627;
	wire [4-1:0] node7631;
	wire [4-1:0] node7632;
	wire [4-1:0] node7633;
	wire [4-1:0] node7634;
	wire [4-1:0] node7635;
	wire [4-1:0] node7636;
	wire [4-1:0] node7638;
	wire [4-1:0] node7641;
	wire [4-1:0] node7644;
	wire [4-1:0] node7645;
	wire [4-1:0] node7646;
	wire [4-1:0] node7649;
	wire [4-1:0] node7653;
	wire [4-1:0] node7654;
	wire [4-1:0] node7655;
	wire [4-1:0] node7656;
	wire [4-1:0] node7660;
	wire [4-1:0] node7661;
	wire [4-1:0] node7664;
	wire [4-1:0] node7667;
	wire [4-1:0] node7668;
	wire [4-1:0] node7671;
	wire [4-1:0] node7672;
	wire [4-1:0] node7676;
	wire [4-1:0] node7677;
	wire [4-1:0] node7678;
	wire [4-1:0] node7680;
	wire [4-1:0] node7682;
	wire [4-1:0] node7685;
	wire [4-1:0] node7686;
	wire [4-1:0] node7688;
	wire [4-1:0] node7691;
	wire [4-1:0] node7693;
	wire [4-1:0] node7696;
	wire [4-1:0] node7697;
	wire [4-1:0] node7699;
	wire [4-1:0] node7700;
	wire [4-1:0] node7703;
	wire [4-1:0] node7706;
	wire [4-1:0] node7707;
	wire [4-1:0] node7709;
	wire [4-1:0] node7713;
	wire [4-1:0] node7714;
	wire [4-1:0] node7715;
	wire [4-1:0] node7716;
	wire [4-1:0] node7717;
	wire [4-1:0] node7718;
	wire [4-1:0] node7721;
	wire [4-1:0] node7724;
	wire [4-1:0] node7725;
	wire [4-1:0] node7729;
	wire [4-1:0] node7730;
	wire [4-1:0] node7733;
	wire [4-1:0] node7734;
	wire [4-1:0] node7738;
	wire [4-1:0] node7739;
	wire [4-1:0] node7740;
	wire [4-1:0] node7742;
	wire [4-1:0] node7745;
	wire [4-1:0] node7746;
	wire [4-1:0] node7750;
	wire [4-1:0] node7751;
	wire [4-1:0] node7753;
	wire [4-1:0] node7756;
	wire [4-1:0] node7757;
	wire [4-1:0] node7760;
	wire [4-1:0] node7763;
	wire [4-1:0] node7764;
	wire [4-1:0] node7765;
	wire [4-1:0] node7766;
	wire [4-1:0] node7768;
	wire [4-1:0] node7771;
	wire [4-1:0] node7772;
	wire [4-1:0] node7775;
	wire [4-1:0] node7778;
	wire [4-1:0] node7779;
	wire [4-1:0] node7780;
	wire [4-1:0] node7783;
	wire [4-1:0] node7786;
	wire [4-1:0] node7787;
	wire [4-1:0] node7791;
	wire [4-1:0] node7792;
	wire [4-1:0] node7793;
	wire [4-1:0] node7794;
	wire [4-1:0] node7797;
	wire [4-1:0] node7800;
	wire [4-1:0] node7801;
	wire [4-1:0] node7805;
	wire [4-1:0] node7808;
	wire [4-1:0] node7809;
	wire [4-1:0] node7810;
	wire [4-1:0] node7811;
	wire [4-1:0] node7812;
	wire [4-1:0] node7813;
	wire [4-1:0] node7814;
	wire [4-1:0] node7815;
	wire [4-1:0] node7819;
	wire [4-1:0] node7820;
	wire [4-1:0] node7821;
	wire [4-1:0] node7825;
	wire [4-1:0] node7826;
	wire [4-1:0] node7830;
	wire [4-1:0] node7831;
	wire [4-1:0] node7832;
	wire [4-1:0] node7833;
	wire [4-1:0] node7837;
	wire [4-1:0] node7838;
	wire [4-1:0] node7842;
	wire [4-1:0] node7843;
	wire [4-1:0] node7846;
	wire [4-1:0] node7847;
	wire [4-1:0] node7851;
	wire [4-1:0] node7852;
	wire [4-1:0] node7853;
	wire [4-1:0] node7854;
	wire [4-1:0] node7855;
	wire [4-1:0] node7858;
	wire [4-1:0] node7861;
	wire [4-1:0] node7864;
	wire [4-1:0] node7865;
	wire [4-1:0] node7867;
	wire [4-1:0] node7870;
	wire [4-1:0] node7873;
	wire [4-1:0] node7874;
	wire [4-1:0] node7875;
	wire [4-1:0] node7878;
	wire [4-1:0] node7879;
	wire [4-1:0] node7883;
	wire [4-1:0] node7884;
	wire [4-1:0] node7885;
	wire [4-1:0] node7888;
	wire [4-1:0] node7891;
	wire [4-1:0] node7892;
	wire [4-1:0] node7896;
	wire [4-1:0] node7897;
	wire [4-1:0] node7898;
	wire [4-1:0] node7899;
	wire [4-1:0] node7900;
	wire [4-1:0] node7903;
	wire [4-1:0] node7906;
	wire [4-1:0] node7907;
	wire [4-1:0] node7908;
	wire [4-1:0] node7911;
	wire [4-1:0] node7914;
	wire [4-1:0] node7916;
	wire [4-1:0] node7919;
	wire [4-1:0] node7920;
	wire [4-1:0] node7921;
	wire [4-1:0] node7922;
	wire [4-1:0] node7925;
	wire [4-1:0] node7928;
	wire [4-1:0] node7929;
	wire [4-1:0] node7933;
	wire [4-1:0] node7935;
	wire [4-1:0] node7936;
	wire [4-1:0] node7940;
	wire [4-1:0] node7941;
	wire [4-1:0] node7942;
	wire [4-1:0] node7943;
	wire [4-1:0] node7944;
	wire [4-1:0] node7949;
	wire [4-1:0] node7951;
	wire [4-1:0] node7952;
	wire [4-1:0] node7956;
	wire [4-1:0] node7957;
	wire [4-1:0] node7958;
	wire [4-1:0] node7961;
	wire [4-1:0] node7962;
	wire [4-1:0] node7966;
	wire [4-1:0] node7968;
	wire [4-1:0] node7971;
	wire [4-1:0] node7972;
	wire [4-1:0] node7973;
	wire [4-1:0] node7974;
	wire [4-1:0] node7975;
	wire [4-1:0] node7977;
	wire [4-1:0] node7978;
	wire [4-1:0] node7982;
	wire [4-1:0] node7983;
	wire [4-1:0] node7984;
	wire [4-1:0] node7987;
	wire [4-1:0] node7990;
	wire [4-1:0] node7993;
	wire [4-1:0] node7994;
	wire [4-1:0] node7995;
	wire [4-1:0] node7998;
	wire [4-1:0] node8000;
	wire [4-1:0] node8003;
	wire [4-1:0] node8004;
	wire [4-1:0] node8006;
	wire [4-1:0] node8009;
	wire [4-1:0] node8010;
	wire [4-1:0] node8014;
	wire [4-1:0] node8015;
	wire [4-1:0] node8016;
	wire [4-1:0] node8017;
	wire [4-1:0] node8018;
	wire [4-1:0] node8022;
	wire [4-1:0] node8023;
	wire [4-1:0] node8027;
	wire [4-1:0] node8029;
	wire [4-1:0] node8031;
	wire [4-1:0] node8034;
	wire [4-1:0] node8035;
	wire [4-1:0] node8036;
	wire [4-1:0] node8037;
	wire [4-1:0] node8040;
	wire [4-1:0] node8043;
	wire [4-1:0] node8046;
	wire [4-1:0] node8047;
	wire [4-1:0] node8050;
	wire [4-1:0] node8051;
	wire [4-1:0] node8055;
	wire [4-1:0] node8056;
	wire [4-1:0] node8057;
	wire [4-1:0] node8058;
	wire [4-1:0] node8059;
	wire [4-1:0] node8060;
	wire [4-1:0] node8063;
	wire [4-1:0] node8066;
	wire [4-1:0] node8069;
	wire [4-1:0] node8070;
	wire [4-1:0] node8071;
	wire [4-1:0] node8075;
	wire [4-1:0] node8078;
	wire [4-1:0] node8079;
	wire [4-1:0] node8080;
	wire [4-1:0] node8082;
	wire [4-1:0] node8085;
	wire [4-1:0] node8087;
	wire [4-1:0] node8090;
	wire [4-1:0] node8091;
	wire [4-1:0] node8093;
	wire [4-1:0] node8096;
	wire [4-1:0] node8097;
	wire [4-1:0] node8100;
	wire [4-1:0] node8103;
	wire [4-1:0] node8104;
	wire [4-1:0] node8105;
	wire [4-1:0] node8106;
	wire [4-1:0] node8107;
	wire [4-1:0] node8110;
	wire [4-1:0] node8113;
	wire [4-1:0] node8114;
	wire [4-1:0] node8118;
	wire [4-1:0] node8119;
	wire [4-1:0] node8121;
	wire [4-1:0] node8124;
	wire [4-1:0] node8125;
	wire [4-1:0] node8129;
	wire [4-1:0] node8130;
	wire [4-1:0] node8131;
	wire [4-1:0] node8132;
	wire [4-1:0] node8137;
	wire [4-1:0] node8138;
	wire [4-1:0] node8139;
	wire [4-1:0] node8142;
	wire [4-1:0] node8145;
	wire [4-1:0] node8147;
	wire [4-1:0] node8150;
	wire [4-1:0] node8151;
	wire [4-1:0] node8152;
	wire [4-1:0] node8153;
	wire [4-1:0] node8154;
	wire [4-1:0] node8155;
	wire [4-1:0] node8156;
	wire [4-1:0] node8157;
	wire [4-1:0] node8162;
	wire [4-1:0] node8163;
	wire [4-1:0] node8165;
	wire [4-1:0] node8168;
	wire [4-1:0] node8171;
	wire [4-1:0] node8172;
	wire [4-1:0] node8173;
	wire [4-1:0] node8176;
	wire [4-1:0] node8177;
	wire [4-1:0] node8181;
	wire [4-1:0] node8182;
	wire [4-1:0] node8183;
	wire [4-1:0] node8186;
	wire [4-1:0] node8189;
	wire [4-1:0] node8190;
	wire [4-1:0] node8194;
	wire [4-1:0] node8195;
	wire [4-1:0] node8196;
	wire [4-1:0] node8197;
	wire [4-1:0] node8198;
	wire [4-1:0] node8201;
	wire [4-1:0] node8204;
	wire [4-1:0] node8205;
	wire [4-1:0] node8209;
	wire [4-1:0] node8211;
	wire [4-1:0] node8214;
	wire [4-1:0] node8215;
	wire [4-1:0] node8216;
	wire [4-1:0] node8217;
	wire [4-1:0] node8221;
	wire [4-1:0] node8222;
	wire [4-1:0] node8225;
	wire [4-1:0] node8228;
	wire [4-1:0] node8230;
	wire [4-1:0] node8231;
	wire [4-1:0] node8234;
	wire [4-1:0] node8237;
	wire [4-1:0] node8238;
	wire [4-1:0] node8239;
	wire [4-1:0] node8240;
	wire [4-1:0] node8241;
	wire [4-1:0] node8242;
	wire [4-1:0] node8245;
	wire [4-1:0] node8248;
	wire [4-1:0] node8250;
	wire [4-1:0] node8253;
	wire [4-1:0] node8254;
	wire [4-1:0] node8255;
	wire [4-1:0] node8258;
	wire [4-1:0] node8261;
	wire [4-1:0] node8264;
	wire [4-1:0] node8265;
	wire [4-1:0] node8266;
	wire [4-1:0] node8269;
	wire [4-1:0] node8270;
	wire [4-1:0] node8274;
	wire [4-1:0] node8275;
	wire [4-1:0] node8276;
	wire [4-1:0] node8280;
	wire [4-1:0] node8283;
	wire [4-1:0] node8284;
	wire [4-1:0] node8285;
	wire [4-1:0] node8286;
	wire [4-1:0] node8288;
	wire [4-1:0] node8291;
	wire [4-1:0] node8292;
	wire [4-1:0] node8296;
	wire [4-1:0] node8298;
	wire [4-1:0] node8300;
	wire [4-1:0] node8303;
	wire [4-1:0] node8304;
	wire [4-1:0] node8306;
	wire [4-1:0] node8307;
	wire [4-1:0] node8311;
	wire [4-1:0] node8312;
	wire [4-1:0] node8313;
	wire [4-1:0] node8317;
	wire [4-1:0] node8318;
	wire [4-1:0] node8322;
	wire [4-1:0] node8323;
	wire [4-1:0] node8324;
	wire [4-1:0] node8325;
	wire [4-1:0] node8326;
	wire [4-1:0] node8327;
	wire [4-1:0] node8328;
	wire [4-1:0] node8332;
	wire [4-1:0] node8334;
	wire [4-1:0] node8337;
	wire [4-1:0] node8338;
	wire [4-1:0] node8341;
	wire [4-1:0] node8342;
	wire [4-1:0] node8346;
	wire [4-1:0] node8347;
	wire [4-1:0] node8348;
	wire [4-1:0] node8352;
	wire [4-1:0] node8353;
	wire [4-1:0] node8357;
	wire [4-1:0] node8358;
	wire [4-1:0] node8359;
	wire [4-1:0] node8360;
	wire [4-1:0] node8362;
	wire [4-1:0] node8366;
	wire [4-1:0] node8367;
	wire [4-1:0] node8369;
	wire [4-1:0] node8372;
	wire [4-1:0] node8374;
	wire [4-1:0] node8377;
	wire [4-1:0] node8378;
	wire [4-1:0] node8379;
	wire [4-1:0] node8380;
	wire [4-1:0] node8383;
	wire [4-1:0] node8386;
	wire [4-1:0] node8387;
	wire [4-1:0] node8390;
	wire [4-1:0] node8393;
	wire [4-1:0] node8394;
	wire [4-1:0] node8395;
	wire [4-1:0] node8398;
	wire [4-1:0] node8401;
	wire [4-1:0] node8402;
	wire [4-1:0] node8406;
	wire [4-1:0] node8407;
	wire [4-1:0] node8408;
	wire [4-1:0] node8409;
	wire [4-1:0] node8410;
	wire [4-1:0] node8412;
	wire [4-1:0] node8415;
	wire [4-1:0] node8416;
	wire [4-1:0] node8420;
	wire [4-1:0] node8421;
	wire [4-1:0] node8425;
	wire [4-1:0] node8426;
	wire [4-1:0] node8427;
	wire [4-1:0] node8428;
	wire [4-1:0] node8434;
	wire [4-1:0] node8435;
	wire [4-1:0] node8436;
	wire [4-1:0] node8437;
	wire [4-1:0] node8438;
	wire [4-1:0] node8442;
	wire [4-1:0] node8445;
	wire [4-1:0] node8447;
	wire [4-1:0] node8448;
	wire [4-1:0] node8451;
	wire [4-1:0] node8454;
	wire [4-1:0] node8455;
	wire [4-1:0] node8456;
	wire [4-1:0] node8457;
	wire [4-1:0] node8461;
	wire [4-1:0] node8464;
	wire [4-1:0] node8465;
	wire [4-1:0] node8466;
	wire [4-1:0] node8470;
	wire [4-1:0] node8471;
	wire [4-1:0] node8474;
	wire [4-1:0] node8477;
	wire [4-1:0] node8478;
	wire [4-1:0] node8479;
	wire [4-1:0] node8480;
	wire [4-1:0] node8481;
	wire [4-1:0] node8482;
	wire [4-1:0] node8483;
	wire [4-1:0] node8484;
	wire [4-1:0] node8485;
	wire [4-1:0] node8486;
	wire [4-1:0] node8487;
	wire [4-1:0] node8491;
	wire [4-1:0] node8492;
	wire [4-1:0] node8496;
	wire [4-1:0] node8497;
	wire [4-1:0] node8498;
	wire [4-1:0] node8501;
	wire [4-1:0] node8505;
	wire [4-1:0] node8506;
	wire [4-1:0] node8507;
	wire [4-1:0] node8508;
	wire [4-1:0] node8512;
	wire [4-1:0] node8513;
	wire [4-1:0] node8517;
	wire [4-1:0] node8518;
	wire [4-1:0] node8519;
	wire [4-1:0] node8524;
	wire [4-1:0] node8525;
	wire [4-1:0] node8526;
	wire [4-1:0] node8529;
	wire [4-1:0] node8530;
	wire [4-1:0] node8531;
	wire [4-1:0] node8535;
	wire [4-1:0] node8536;
	wire [4-1:0] node8539;
	wire [4-1:0] node8542;
	wire [4-1:0] node8543;
	wire [4-1:0] node8544;
	wire [4-1:0] node8548;
	wire [4-1:0] node8550;
	wire [4-1:0] node8553;
	wire [4-1:0] node8554;
	wire [4-1:0] node8555;
	wire [4-1:0] node8556;
	wire [4-1:0] node8557;
	wire [4-1:0] node8558;
	wire [4-1:0] node8562;
	wire [4-1:0] node8564;
	wire [4-1:0] node8567;
	wire [4-1:0] node8568;
	wire [4-1:0] node8569;
	wire [4-1:0] node8573;
	wire [4-1:0] node8575;
	wire [4-1:0] node8578;
	wire [4-1:0] node8579;
	wire [4-1:0] node8580;
	wire [4-1:0] node8581;
	wire [4-1:0] node8585;
	wire [4-1:0] node8588;
	wire [4-1:0] node8590;
	wire [4-1:0] node8591;
	wire [4-1:0] node8595;
	wire [4-1:0] node8596;
	wire [4-1:0] node8597;
	wire [4-1:0] node8598;
	wire [4-1:0] node8599;
	wire [4-1:0] node8602;
	wire [4-1:0] node8605;
	wire [4-1:0] node8606;
	wire [4-1:0] node8609;
	wire [4-1:0] node8612;
	wire [4-1:0] node8613;
	wire [4-1:0] node8615;
	wire [4-1:0] node8618;
	wire [4-1:0] node8619;
	wire [4-1:0] node8623;
	wire [4-1:0] node8624;
	wire [4-1:0] node8625;
	wire [4-1:0] node8627;
	wire [4-1:0] node8630;
	wire [4-1:0] node8633;
	wire [4-1:0] node8635;
	wire [4-1:0] node8637;
	wire [4-1:0] node8640;
	wire [4-1:0] node8641;
	wire [4-1:0] node8642;
	wire [4-1:0] node8643;
	wire [4-1:0] node8644;
	wire [4-1:0] node8646;
	wire [4-1:0] node8649;
	wire [4-1:0] node8650;
	wire [4-1:0] node8653;
	wire [4-1:0] node8655;
	wire [4-1:0] node8658;
	wire [4-1:0] node8659;
	wire [4-1:0] node8660;
	wire [4-1:0] node8661;
	wire [4-1:0] node8665;
	wire [4-1:0] node8666;
	wire [4-1:0] node8669;
	wire [4-1:0] node8672;
	wire [4-1:0] node8673;
	wire [4-1:0] node8674;
	wire [4-1:0] node8678;
	wire [4-1:0] node8681;
	wire [4-1:0] node8682;
	wire [4-1:0] node8683;
	wire [4-1:0] node8685;
	wire [4-1:0] node8686;
	wire [4-1:0] node8689;
	wire [4-1:0] node8692;
	wire [4-1:0] node8693;
	wire [4-1:0] node8696;
	wire [4-1:0] node8698;
	wire [4-1:0] node8701;
	wire [4-1:0] node8702;
	wire [4-1:0] node8705;
	wire [4-1:0] node8706;
	wire [4-1:0] node8709;
	wire [4-1:0] node8710;
	wire [4-1:0] node8714;
	wire [4-1:0] node8715;
	wire [4-1:0] node8716;
	wire [4-1:0] node8717;
	wire [4-1:0] node8718;
	wire [4-1:0] node8719;
	wire [4-1:0] node8724;
	wire [4-1:0] node8726;
	wire [4-1:0] node8729;
	wire [4-1:0] node8730;
	wire [4-1:0] node8731;
	wire [4-1:0] node8732;
	wire [4-1:0] node8735;
	wire [4-1:0] node8738;
	wire [4-1:0] node8740;
	wire [4-1:0] node8743;
	wire [4-1:0] node8744;
	wire [4-1:0] node8745;
	wire [4-1:0] node8749;
	wire [4-1:0] node8751;
	wire [4-1:0] node8754;
	wire [4-1:0] node8755;
	wire [4-1:0] node8756;
	wire [4-1:0] node8757;
	wire [4-1:0] node8759;
	wire [4-1:0] node8762;
	wire [4-1:0] node8763;
	wire [4-1:0] node8767;
	wire [4-1:0] node8768;
	wire [4-1:0] node8770;
	wire [4-1:0] node8773;
	wire [4-1:0] node8775;
	wire [4-1:0] node8778;
	wire [4-1:0] node8779;
	wire [4-1:0] node8780;
	wire [4-1:0] node8782;
	wire [4-1:0] node8785;
	wire [4-1:0] node8786;
	wire [4-1:0] node8790;
	wire [4-1:0] node8791;
	wire [4-1:0] node8793;
	wire [4-1:0] node8797;
	wire [4-1:0] node8798;
	wire [4-1:0] node8799;
	wire [4-1:0] node8800;
	wire [4-1:0] node8801;
	wire [4-1:0] node8802;
	wire [4-1:0] node8803;
	wire [4-1:0] node8805;
	wire [4-1:0] node8809;
	wire [4-1:0] node8810;
	wire [4-1:0] node8811;
	wire [4-1:0] node8816;
	wire [4-1:0] node8817;
	wire [4-1:0] node8818;
	wire [4-1:0] node8820;
	wire [4-1:0] node8823;
	wire [4-1:0] node8824;
	wire [4-1:0] node8828;
	wire [4-1:0] node8829;
	wire [4-1:0] node8830;
	wire [4-1:0] node8833;
	wire [4-1:0] node8836;
	wire [4-1:0] node8839;
	wire [4-1:0] node8840;
	wire [4-1:0] node8841;
	wire [4-1:0] node8842;
	wire [4-1:0] node8845;
	wire [4-1:0] node8848;
	wire [4-1:0] node8849;
	wire [4-1:0] node8851;
	wire [4-1:0] node8854;
	wire [4-1:0] node8855;
	wire [4-1:0] node8859;
	wire [4-1:0] node8860;
	wire [4-1:0] node8861;
	wire [4-1:0] node8863;
	wire [4-1:0] node8866;
	wire [4-1:0] node8867;
	wire [4-1:0] node8871;
	wire [4-1:0] node8872;
	wire [4-1:0] node8873;
	wire [4-1:0] node8878;
	wire [4-1:0] node8879;
	wire [4-1:0] node8880;
	wire [4-1:0] node8881;
	wire [4-1:0] node8882;
	wire [4-1:0] node8884;
	wire [4-1:0] node8887;
	wire [4-1:0] node8889;
	wire [4-1:0] node8892;
	wire [4-1:0] node8893;
	wire [4-1:0] node8895;
	wire [4-1:0] node8898;
	wire [4-1:0] node8901;
	wire [4-1:0] node8902;
	wire [4-1:0] node8903;
	wire [4-1:0] node8906;
	wire [4-1:0] node8908;
	wire [4-1:0] node8911;
	wire [4-1:0] node8912;
	wire [4-1:0] node8913;
	wire [4-1:0] node8916;
	wire [4-1:0] node8920;
	wire [4-1:0] node8921;
	wire [4-1:0] node8922;
	wire [4-1:0] node8923;
	wire [4-1:0] node8924;
	wire [4-1:0] node8928;
	wire [4-1:0] node8930;
	wire [4-1:0] node8933;
	wire [4-1:0] node8934;
	wire [4-1:0] node8935;
	wire [4-1:0] node8938;
	wire [4-1:0] node8941;
	wire [4-1:0] node8943;
	wire [4-1:0] node8946;
	wire [4-1:0] node8947;
	wire [4-1:0] node8948;
	wire [4-1:0] node8949;
	wire [4-1:0] node8952;
	wire [4-1:0] node8955;
	wire [4-1:0] node8956;
	wire [4-1:0] node8960;
	wire [4-1:0] node8962;
	wire [4-1:0] node8964;
	wire [4-1:0] node8967;
	wire [4-1:0] node8968;
	wire [4-1:0] node8969;
	wire [4-1:0] node8970;
	wire [4-1:0] node8971;
	wire [4-1:0] node8972;
	wire [4-1:0] node8974;
	wire [4-1:0] node8977;
	wire [4-1:0] node8978;
	wire [4-1:0] node8981;
	wire [4-1:0] node8984;
	wire [4-1:0] node8985;
	wire [4-1:0] node8986;
	wire [4-1:0] node8989;
	wire [4-1:0] node8992;
	wire [4-1:0] node8993;
	wire [4-1:0] node8997;
	wire [4-1:0] node8998;
	wire [4-1:0] node8999;
	wire [4-1:0] node9000;
	wire [4-1:0] node9003;
	wire [4-1:0] node9006;
	wire [4-1:0] node9009;
	wire [4-1:0] node9010;
	wire [4-1:0] node9011;
	wire [4-1:0] node9015;
	wire [4-1:0] node9016;
	wire [4-1:0] node9019;
	wire [4-1:0] node9022;
	wire [4-1:0] node9023;
	wire [4-1:0] node9024;
	wire [4-1:0] node9026;
	wire [4-1:0] node9028;
	wire [4-1:0] node9031;
	wire [4-1:0] node9033;
	wire [4-1:0] node9034;
	wire [4-1:0] node9037;
	wire [4-1:0] node9040;
	wire [4-1:0] node9041;
	wire [4-1:0] node9042;
	wire [4-1:0] node9043;
	wire [4-1:0] node9046;
	wire [4-1:0] node9049;
	wire [4-1:0] node9051;
	wire [4-1:0] node9054;
	wire [4-1:0] node9055;
	wire [4-1:0] node9056;
	wire [4-1:0] node9060;
	wire [4-1:0] node9061;
	wire [4-1:0] node9065;
	wire [4-1:0] node9066;
	wire [4-1:0] node9067;
	wire [4-1:0] node9068;
	wire [4-1:0] node9069;
	wire [4-1:0] node9070;
	wire [4-1:0] node9074;
	wire [4-1:0] node9075;
	wire [4-1:0] node9078;
	wire [4-1:0] node9081;
	wire [4-1:0] node9082;
	wire [4-1:0] node9083;
	wire [4-1:0] node9087;
	wire [4-1:0] node9088;
	wire [4-1:0] node9092;
	wire [4-1:0] node9093;
	wire [4-1:0] node9095;
	wire [4-1:0] node9098;
	wire [4-1:0] node9100;
	wire [4-1:0] node9101;
	wire [4-1:0] node9104;
	wire [4-1:0] node9107;
	wire [4-1:0] node9108;
	wire [4-1:0] node9109;
	wire [4-1:0] node9110;
	wire [4-1:0] node9113;
	wire [4-1:0] node9114;
	wire [4-1:0] node9117;
	wire [4-1:0] node9120;
	wire [4-1:0] node9121;
	wire [4-1:0] node9122;
	wire [4-1:0] node9125;
	wire [4-1:0] node9128;
	wire [4-1:0] node9130;
	wire [4-1:0] node9133;
	wire [4-1:0] node9134;
	wire [4-1:0] node9135;
	wire [4-1:0] node9136;
	wire [4-1:0] node9139;
	wire [4-1:0] node9142;
	wire [4-1:0] node9143;
	wire [4-1:0] node9146;
	wire [4-1:0] node9149;
	wire [4-1:0] node9150;
	wire [4-1:0] node9152;
	wire [4-1:0] node9155;
	wire [4-1:0] node9157;
	wire [4-1:0] node9160;
	wire [4-1:0] node9161;
	wire [4-1:0] node9162;
	wire [4-1:0] node9163;
	wire [4-1:0] node9164;
	wire [4-1:0] node9165;
	wire [4-1:0] node9166;
	wire [4-1:0] node9167;
	wire [4-1:0] node9170;
	wire [4-1:0] node9171;
	wire [4-1:0] node9174;
	wire [4-1:0] node9177;
	wire [4-1:0] node9178;
	wire [4-1:0] node9179;
	wire [4-1:0] node9182;
	wire [4-1:0] node9185;
	wire [4-1:0] node9186;
	wire [4-1:0] node9190;
	wire [4-1:0] node9191;
	wire [4-1:0] node9192;
	wire [4-1:0] node9193;
	wire [4-1:0] node9196;
	wire [4-1:0] node9199;
	wire [4-1:0] node9202;
	wire [4-1:0] node9203;
	wire [4-1:0] node9204;
	wire [4-1:0] node9207;
	wire [4-1:0] node9210;
	wire [4-1:0] node9211;
	wire [4-1:0] node9214;
	wire [4-1:0] node9217;
	wire [4-1:0] node9218;
	wire [4-1:0] node9219;
	wire [4-1:0] node9220;
	wire [4-1:0] node9221;
	wire [4-1:0] node9225;
	wire [4-1:0] node9227;
	wire [4-1:0] node9230;
	wire [4-1:0] node9231;
	wire [4-1:0] node9232;
	wire [4-1:0] node9236;
	wire [4-1:0] node9239;
	wire [4-1:0] node9240;
	wire [4-1:0] node9241;
	wire [4-1:0] node9243;
	wire [4-1:0] node9246;
	wire [4-1:0] node9247;
	wire [4-1:0] node9251;
	wire [4-1:0] node9252;
	wire [4-1:0] node9253;
	wire [4-1:0] node9257;
	wire [4-1:0] node9258;
	wire [4-1:0] node9262;
	wire [4-1:0] node9263;
	wire [4-1:0] node9264;
	wire [4-1:0] node9265;
	wire [4-1:0] node9266;
	wire [4-1:0] node9267;
	wire [4-1:0] node9270;
	wire [4-1:0] node9273;
	wire [4-1:0] node9274;
	wire [4-1:0] node9278;
	wire [4-1:0] node9279;
	wire [4-1:0] node9280;
	wire [4-1:0] node9285;
	wire [4-1:0] node9286;
	wire [4-1:0] node9287;
	wire [4-1:0] node9289;
	wire [4-1:0] node9292;
	wire [4-1:0] node9293;
	wire [4-1:0] node9297;
	wire [4-1:0] node9298;
	wire [4-1:0] node9300;
	wire [4-1:0] node9303;
	wire [4-1:0] node9306;
	wire [4-1:0] node9307;
	wire [4-1:0] node9308;
	wire [4-1:0] node9309;
	wire [4-1:0] node9310;
	wire [4-1:0] node9313;
	wire [4-1:0] node9316;
	wire [4-1:0] node9318;
	wire [4-1:0] node9321;
	wire [4-1:0] node9322;
	wire [4-1:0] node9325;
	wire [4-1:0] node9327;
	wire [4-1:0] node9330;
	wire [4-1:0] node9331;
	wire [4-1:0] node9332;
	wire [4-1:0] node9333;
	wire [4-1:0] node9338;
	wire [4-1:0] node9339;
	wire [4-1:0] node9342;
	wire [4-1:0] node9345;
	wire [4-1:0] node9346;
	wire [4-1:0] node9347;
	wire [4-1:0] node9348;
	wire [4-1:0] node9349;
	wire [4-1:0] node9350;
	wire [4-1:0] node9351;
	wire [4-1:0] node9354;
	wire [4-1:0] node9357;
	wire [4-1:0] node9358;
	wire [4-1:0] node9361;
	wire [4-1:0] node9364;
	wire [4-1:0] node9365;
	wire [4-1:0] node9367;
	wire [4-1:0] node9370;
	wire [4-1:0] node9372;
	wire [4-1:0] node9375;
	wire [4-1:0] node9376;
	wire [4-1:0] node9377;
	wire [4-1:0] node9378;
	wire [4-1:0] node9382;
	wire [4-1:0] node9384;
	wire [4-1:0] node9387;
	wire [4-1:0] node9388;
	wire [4-1:0] node9391;
	wire [4-1:0] node9392;
	wire [4-1:0] node9395;
	wire [4-1:0] node9398;
	wire [4-1:0] node9399;
	wire [4-1:0] node9400;
	wire [4-1:0] node9401;
	wire [4-1:0] node9402;
	wire [4-1:0] node9406;
	wire [4-1:0] node9409;
	wire [4-1:0] node9410;
	wire [4-1:0] node9411;
	wire [4-1:0] node9415;
	wire [4-1:0] node9418;
	wire [4-1:0] node9419;
	wire [4-1:0] node9420;
	wire [4-1:0] node9421;
	wire [4-1:0] node9424;
	wire [4-1:0] node9427;
	wire [4-1:0] node9430;
	wire [4-1:0] node9431;
	wire [4-1:0] node9432;
	wire [4-1:0] node9435;
	wire [4-1:0] node9438;
	wire [4-1:0] node9439;
	wire [4-1:0] node9443;
	wire [4-1:0] node9444;
	wire [4-1:0] node9445;
	wire [4-1:0] node9446;
	wire [4-1:0] node9447;
	wire [4-1:0] node9448;
	wire [4-1:0] node9452;
	wire [4-1:0] node9455;
	wire [4-1:0] node9456;
	wire [4-1:0] node9457;
	wire [4-1:0] node9461;
	wire [4-1:0] node9463;
	wire [4-1:0] node9466;
	wire [4-1:0] node9467;
	wire [4-1:0] node9468;
	wire [4-1:0] node9471;
	wire [4-1:0] node9474;
	wire [4-1:0] node9475;
	wire [4-1:0] node9476;
	wire [4-1:0] node9480;
	wire [4-1:0] node9483;
	wire [4-1:0] node9484;
	wire [4-1:0] node9485;
	wire [4-1:0] node9486;
	wire [4-1:0] node9488;
	wire [4-1:0] node9491;
	wire [4-1:0] node9493;
	wire [4-1:0] node9496;
	wire [4-1:0] node9498;
	wire [4-1:0] node9500;
	wire [4-1:0] node9503;
	wire [4-1:0] node9504;
	wire [4-1:0] node9505;
	wire [4-1:0] node9506;
	wire [4-1:0] node9510;
	wire [4-1:0] node9513;
	wire [4-1:0] node9514;
	wire [4-1:0] node9515;
	wire [4-1:0] node9518;
	wire [4-1:0] node9522;
	wire [4-1:0] node9523;
	wire [4-1:0] node9524;
	wire [4-1:0] node9525;
	wire [4-1:0] node9526;
	wire [4-1:0] node9527;
	wire [4-1:0] node9528;
	wire [4-1:0] node9530;
	wire [4-1:0] node9533;
	wire [4-1:0] node9536;
	wire [4-1:0] node9537;
	wire [4-1:0] node9538;
	wire [4-1:0] node9542;
	wire [4-1:0] node9543;
	wire [4-1:0] node9547;
	wire [4-1:0] node9548;
	wire [4-1:0] node9549;
	wire [4-1:0] node9552;
	wire [4-1:0] node9553;
	wire [4-1:0] node9557;
	wire [4-1:0] node9558;
	wire [4-1:0] node9559;
	wire [4-1:0] node9563;
	wire [4-1:0] node9564;
	wire [4-1:0] node9568;
	wire [4-1:0] node9569;
	wire [4-1:0] node9570;
	wire [4-1:0] node9571;
	wire [4-1:0] node9573;
	wire [4-1:0] node9577;
	wire [4-1:0] node9578;
	wire [4-1:0] node9579;
	wire [4-1:0] node9583;
	wire [4-1:0] node9584;
	wire [4-1:0] node9588;
	wire [4-1:0] node9589;
	wire [4-1:0] node9590;
	wire [4-1:0] node9592;
	wire [4-1:0] node9596;
	wire [4-1:0] node9598;
	wire [4-1:0] node9600;
	wire [4-1:0] node9603;
	wire [4-1:0] node9604;
	wire [4-1:0] node9605;
	wire [4-1:0] node9606;
	wire [4-1:0] node9607;
	wire [4-1:0] node9609;
	wire [4-1:0] node9612;
	wire [4-1:0] node9614;
	wire [4-1:0] node9617;
	wire [4-1:0] node9618;
	wire [4-1:0] node9620;
	wire [4-1:0] node9623;
	wire [4-1:0] node9625;
	wire [4-1:0] node9628;
	wire [4-1:0] node9629;
	wire [4-1:0] node9630;
	wire [4-1:0] node9631;
	wire [4-1:0] node9635;
	wire [4-1:0] node9636;
	wire [4-1:0] node9640;
	wire [4-1:0] node9641;
	wire [4-1:0] node9642;
	wire [4-1:0] node9645;
	wire [4-1:0] node9648;
	wire [4-1:0] node9649;
	wire [4-1:0] node9652;
	wire [4-1:0] node9655;
	wire [4-1:0] node9656;
	wire [4-1:0] node9657;
	wire [4-1:0] node9658;
	wire [4-1:0] node9661;
	wire [4-1:0] node9664;
	wire [4-1:0] node9665;
	wire [4-1:0] node9668;
	wire [4-1:0] node9669;
	wire [4-1:0] node9673;
	wire [4-1:0] node9674;
	wire [4-1:0] node9676;
	wire [4-1:0] node9677;
	wire [4-1:0] node9681;
	wire [4-1:0] node9682;
	wire [4-1:0] node9685;
	wire [4-1:0] node9688;
	wire [4-1:0] node9689;
	wire [4-1:0] node9690;
	wire [4-1:0] node9691;
	wire [4-1:0] node9692;
	wire [4-1:0] node9693;
	wire [4-1:0] node9696;
	wire [4-1:0] node9698;
	wire [4-1:0] node9701;
	wire [4-1:0] node9702;
	wire [4-1:0] node9705;
	wire [4-1:0] node9707;
	wire [4-1:0] node9710;
	wire [4-1:0] node9711;
	wire [4-1:0] node9712;
	wire [4-1:0] node9713;
	wire [4-1:0] node9716;
	wire [4-1:0] node9719;
	wire [4-1:0] node9720;
	wire [4-1:0] node9724;
	wire [4-1:0] node9725;
	wire [4-1:0] node9727;
	wire [4-1:0] node9730;
	wire [4-1:0] node9732;
	wire [4-1:0] node9735;
	wire [4-1:0] node9736;
	wire [4-1:0] node9737;
	wire [4-1:0] node9738;
	wire [4-1:0] node9739;
	wire [4-1:0] node9743;
	wire [4-1:0] node9744;
	wire [4-1:0] node9748;
	wire [4-1:0] node9749;
	wire [4-1:0] node9750;
	wire [4-1:0] node9753;
	wire [4-1:0] node9756;
	wire [4-1:0] node9757;
	wire [4-1:0] node9761;
	wire [4-1:0] node9762;
	wire [4-1:0] node9763;
	wire [4-1:0] node9764;
	wire [4-1:0] node9767;
	wire [4-1:0] node9770;
	wire [4-1:0] node9772;
	wire [4-1:0] node9775;
	wire [4-1:0] node9777;
	wire [4-1:0] node9780;
	wire [4-1:0] node9781;
	wire [4-1:0] node9782;
	wire [4-1:0] node9783;
	wire [4-1:0] node9784;
	wire [4-1:0] node9785;
	wire [4-1:0] node9790;
	wire [4-1:0] node9792;
	wire [4-1:0] node9793;
	wire [4-1:0] node9796;
	wire [4-1:0] node9799;
	wire [4-1:0] node9800;
	wire [4-1:0] node9801;
	wire [4-1:0] node9803;
	wire [4-1:0] node9806;
	wire [4-1:0] node9807;
	wire [4-1:0] node9810;
	wire [4-1:0] node9813;
	wire [4-1:0] node9814;
	wire [4-1:0] node9817;
	wire [4-1:0] node9818;
	wire [4-1:0] node9821;
	wire [4-1:0] node9824;
	wire [4-1:0] node9825;
	wire [4-1:0] node9826;
	wire [4-1:0] node9827;
	wire [4-1:0] node9829;
	wire [4-1:0] node9832;
	wire [4-1:0] node9834;
	wire [4-1:0] node9837;
	wire [4-1:0] node9838;
	wire [4-1:0] node9839;
	wire [4-1:0] node9843;
	wire [4-1:0] node9844;
	wire [4-1:0] node9847;
	wire [4-1:0] node9850;
	wire [4-1:0] node9851;
	wire [4-1:0] node9852;
	wire [4-1:0] node9853;
	wire [4-1:0] node9856;
	wire [4-1:0] node9859;
	wire [4-1:0] node9860;
	wire [4-1:0] node9863;
	wire [4-1:0] node9866;
	wire [4-1:0] node9867;
	wire [4-1:0] node9868;
	wire [4-1:0] node9872;
	wire [4-1:0] node9875;
	wire [4-1:0] node9876;
	wire [4-1:0] node9877;
	wire [4-1:0] node9878;
	wire [4-1:0] node9879;
	wire [4-1:0] node9880;
	wire [4-1:0] node9881;
	wire [4-1:0] node9882;
	wire [4-1:0] node9883;
	wire [4-1:0] node9885;
	wire [4-1:0] node9888;
	wire [4-1:0] node9889;
	wire [4-1:0] node9893;
	wire [4-1:0] node9894;
	wire [4-1:0] node9895;
	wire [4-1:0] node9898;
	wire [4-1:0] node9901;
	wire [4-1:0] node9902;
	wire [4-1:0] node9906;
	wire [4-1:0] node9907;
	wire [4-1:0] node9908;
	wire [4-1:0] node9910;
	wire [4-1:0] node9913;
	wire [4-1:0] node9915;
	wire [4-1:0] node9918;
	wire [4-1:0] node9919;
	wire [4-1:0] node9920;
	wire [4-1:0] node9923;
	wire [4-1:0] node9926;
	wire [4-1:0] node9927;
	wire [4-1:0] node9930;
	wire [4-1:0] node9933;
	wire [4-1:0] node9934;
	wire [4-1:0] node9935;
	wire [4-1:0] node9936;
	wire [4-1:0] node9937;
	wire [4-1:0] node9941;
	wire [4-1:0] node9942;
	wire [4-1:0] node9946;
	wire [4-1:0] node9947;
	wire [4-1:0] node9950;
	wire [4-1:0] node9952;
	wire [4-1:0] node9955;
	wire [4-1:0] node9956;
	wire [4-1:0] node9957;
	wire [4-1:0] node9960;
	wire [4-1:0] node9962;
	wire [4-1:0] node9965;
	wire [4-1:0] node9966;
	wire [4-1:0] node9969;
	wire [4-1:0] node9971;
	wire [4-1:0] node9974;
	wire [4-1:0] node9975;
	wire [4-1:0] node9976;
	wire [4-1:0] node9977;
	wire [4-1:0] node9978;
	wire [4-1:0] node9981;
	wire [4-1:0] node9983;
	wire [4-1:0] node9986;
	wire [4-1:0] node9987;
	wire [4-1:0] node9989;
	wire [4-1:0] node9992;
	wire [4-1:0] node9993;
	wire [4-1:0] node9997;
	wire [4-1:0] node9998;
	wire [4-1:0] node9999;
	wire [4-1:0] node10000;
	wire [4-1:0] node10004;
	wire [4-1:0] node10007;
	wire [4-1:0] node10008;
	wire [4-1:0] node10011;
	wire [4-1:0] node10012;
	wire [4-1:0] node10015;
	wire [4-1:0] node10018;
	wire [4-1:0] node10019;
	wire [4-1:0] node10020;
	wire [4-1:0] node10021;
	wire [4-1:0] node10022;
	wire [4-1:0] node10025;
	wire [4-1:0] node10028;
	wire [4-1:0] node10030;
	wire [4-1:0] node10033;
	wire [4-1:0] node10034;
	wire [4-1:0] node10035;
	wire [4-1:0] node10038;
	wire [4-1:0] node10041;
	wire [4-1:0] node10043;
	wire [4-1:0] node10046;
	wire [4-1:0] node10047;
	wire [4-1:0] node10048;
	wire [4-1:0] node10049;
	wire [4-1:0] node10053;
	wire [4-1:0] node10054;
	wire [4-1:0] node10058;
	wire [4-1:0] node10059;
	wire [4-1:0] node10062;
	wire [4-1:0] node10064;
	wire [4-1:0] node10067;
	wire [4-1:0] node10068;
	wire [4-1:0] node10069;
	wire [4-1:0] node10070;
	wire [4-1:0] node10071;
	wire [4-1:0] node10072;
	wire [4-1:0] node10073;
	wire [4-1:0] node10078;
	wire [4-1:0] node10080;
	wire [4-1:0] node10081;
	wire [4-1:0] node10085;
	wire [4-1:0] node10086;
	wire [4-1:0] node10087;
	wire [4-1:0] node10089;
	wire [4-1:0] node10092;
	wire [4-1:0] node10093;
	wire [4-1:0] node10096;
	wire [4-1:0] node10099;
	wire [4-1:0] node10100;
	wire [4-1:0] node10101;
	wire [4-1:0] node10105;
	wire [4-1:0] node10108;
	wire [4-1:0] node10109;
	wire [4-1:0] node10110;
	wire [4-1:0] node10111;
	wire [4-1:0] node10112;
	wire [4-1:0] node10116;
	wire [4-1:0] node10117;
	wire [4-1:0] node10120;
	wire [4-1:0] node10123;
	wire [4-1:0] node10124;
	wire [4-1:0] node10127;
	wire [4-1:0] node10128;
	wire [4-1:0] node10131;
	wire [4-1:0] node10134;
	wire [4-1:0] node10135;
	wire [4-1:0] node10136;
	wire [4-1:0] node10137;
	wire [4-1:0] node10140;
	wire [4-1:0] node10143;
	wire [4-1:0] node10146;
	wire [4-1:0] node10147;
	wire [4-1:0] node10148;
	wire [4-1:0] node10151;
	wire [4-1:0] node10154;
	wire [4-1:0] node10157;
	wire [4-1:0] node10158;
	wire [4-1:0] node10159;
	wire [4-1:0] node10160;
	wire [4-1:0] node10161;
	wire [4-1:0] node10163;
	wire [4-1:0] node10166;
	wire [4-1:0] node10167;
	wire [4-1:0] node10171;
	wire [4-1:0] node10172;
	wire [4-1:0] node10175;
	wire [4-1:0] node10176;
	wire [4-1:0] node10179;
	wire [4-1:0] node10182;
	wire [4-1:0] node10183;
	wire [4-1:0] node10184;
	wire [4-1:0] node10185;
	wire [4-1:0] node10188;
	wire [4-1:0] node10192;
	wire [4-1:0] node10193;
	wire [4-1:0] node10194;
	wire [4-1:0] node10198;
	wire [4-1:0] node10199;
	wire [4-1:0] node10203;
	wire [4-1:0] node10204;
	wire [4-1:0] node10205;
	wire [4-1:0] node10206;
	wire [4-1:0] node10207;
	wire [4-1:0] node10210;
	wire [4-1:0] node10213;
	wire [4-1:0] node10214;
	wire [4-1:0] node10217;
	wire [4-1:0] node10220;
	wire [4-1:0] node10221;
	wire [4-1:0] node10222;
	wire [4-1:0] node10226;
	wire [4-1:0] node10227;
	wire [4-1:0] node10231;
	wire [4-1:0] node10232;
	wire [4-1:0] node10233;
	wire [4-1:0] node10235;
	wire [4-1:0] node10238;
	wire [4-1:0] node10239;
	wire [4-1:0] node10242;
	wire [4-1:0] node10245;
	wire [4-1:0] node10246;
	wire [4-1:0] node10248;
	wire [4-1:0] node10252;
	wire [4-1:0] node10253;
	wire [4-1:0] node10254;
	wire [4-1:0] node10255;
	wire [4-1:0] node10256;
	wire [4-1:0] node10257;
	wire [4-1:0] node10258;
	wire [4-1:0] node10259;
	wire [4-1:0] node10263;
	wire [4-1:0] node10264;
	wire [4-1:0] node10267;
	wire [4-1:0] node10270;
	wire [4-1:0] node10271;
	wire [4-1:0] node10273;
	wire [4-1:0] node10276;
	wire [4-1:0] node10277;
	wire [4-1:0] node10281;
	wire [4-1:0] node10282;
	wire [4-1:0] node10283;
	wire [4-1:0] node10284;
	wire [4-1:0] node10287;
	wire [4-1:0] node10290;
	wire [4-1:0] node10291;
	wire [4-1:0] node10294;
	wire [4-1:0] node10297;
	wire [4-1:0] node10299;
	wire [4-1:0] node10300;
	wire [4-1:0] node10304;
	wire [4-1:0] node10305;
	wire [4-1:0] node10306;
	wire [4-1:0] node10307;
	wire [4-1:0] node10308;
	wire [4-1:0] node10312;
	wire [4-1:0] node10313;
	wire [4-1:0] node10316;
	wire [4-1:0] node10319;
	wire [4-1:0] node10320;
	wire [4-1:0] node10323;
	wire [4-1:0] node10324;
	wire [4-1:0] node10328;
	wire [4-1:0] node10329;
	wire [4-1:0] node10330;
	wire [4-1:0] node10332;
	wire [4-1:0] node10335;
	wire [4-1:0] node10336;
	wire [4-1:0] node10339;
	wire [4-1:0] node10342;
	wire [4-1:0] node10343;
	wire [4-1:0] node10344;
	wire [4-1:0] node10347;
	wire [4-1:0] node10350;
	wire [4-1:0] node10352;
	wire [4-1:0] node10355;
	wire [4-1:0] node10356;
	wire [4-1:0] node10357;
	wire [4-1:0] node10358;
	wire [4-1:0] node10360;
	wire [4-1:0] node10362;
	wire [4-1:0] node10365;
	wire [4-1:0] node10366;
	wire [4-1:0] node10367;
	wire [4-1:0] node10370;
	wire [4-1:0] node10373;
	wire [4-1:0] node10376;
	wire [4-1:0] node10377;
	wire [4-1:0] node10378;
	wire [4-1:0] node10379;
	wire [4-1:0] node10382;
	wire [4-1:0] node10385;
	wire [4-1:0] node10388;
	wire [4-1:0] node10389;
	wire [4-1:0] node10391;
	wire [4-1:0] node10394;
	wire [4-1:0] node10395;
	wire [4-1:0] node10398;
	wire [4-1:0] node10401;
	wire [4-1:0] node10402;
	wire [4-1:0] node10403;
	wire [4-1:0] node10405;
	wire [4-1:0] node10408;
	wire [4-1:0] node10409;
	wire [4-1:0] node10411;
	wire [4-1:0] node10414;
	wire [4-1:0] node10416;
	wire [4-1:0] node10419;
	wire [4-1:0] node10420;
	wire [4-1:0] node10421;
	wire [4-1:0] node10423;
	wire [4-1:0] node10426;
	wire [4-1:0] node10427;
	wire [4-1:0] node10430;
	wire [4-1:0] node10433;
	wire [4-1:0] node10434;
	wire [4-1:0] node10436;
	wire [4-1:0] node10439;
	wire [4-1:0] node10440;
	wire [4-1:0] node10444;
	wire [4-1:0] node10445;
	wire [4-1:0] node10446;
	wire [4-1:0] node10447;
	wire [4-1:0] node10448;
	wire [4-1:0] node10450;
	wire [4-1:0] node10451;
	wire [4-1:0] node10455;
	wire [4-1:0] node10456;
	wire [4-1:0] node10457;
	wire [4-1:0] node10462;
	wire [4-1:0] node10463;
	wire [4-1:0] node10464;
	wire [4-1:0] node10466;
	wire [4-1:0] node10469;
	wire [4-1:0] node10471;
	wire [4-1:0] node10474;
	wire [4-1:0] node10476;
	wire [4-1:0] node10477;
	wire [4-1:0] node10481;
	wire [4-1:0] node10482;
	wire [4-1:0] node10483;
	wire [4-1:0] node10484;
	wire [4-1:0] node10485;
	wire [4-1:0] node10489;
	wire [4-1:0] node10490;
	wire [4-1:0] node10494;
	wire [4-1:0] node10495;
	wire [4-1:0] node10496;
	wire [4-1:0] node10501;
	wire [4-1:0] node10502;
	wire [4-1:0] node10503;
	wire [4-1:0] node10505;
	wire [4-1:0] node10508;
	wire [4-1:0] node10509;
	wire [4-1:0] node10513;
	wire [4-1:0] node10514;
	wire [4-1:0] node10515;
	wire [4-1:0] node10518;
	wire [4-1:0] node10521;
	wire [4-1:0] node10522;
	wire [4-1:0] node10525;
	wire [4-1:0] node10528;
	wire [4-1:0] node10529;
	wire [4-1:0] node10530;
	wire [4-1:0] node10531;
	wire [4-1:0] node10532;
	wire [4-1:0] node10533;
	wire [4-1:0] node10537;
	wire [4-1:0] node10540;
	wire [4-1:0] node10541;
	wire [4-1:0] node10545;
	wire [4-1:0] node10546;
	wire [4-1:0] node10547;
	wire [4-1:0] node10548;
	wire [4-1:0] node10552;
	wire [4-1:0] node10553;
	wire [4-1:0] node10557;
	wire [4-1:0] node10559;
	wire [4-1:0] node10560;
	wire [4-1:0] node10564;
	wire [4-1:0] node10565;
	wire [4-1:0] node10566;
	wire [4-1:0] node10567;
	wire [4-1:0] node10568;
	wire [4-1:0] node10572;
	wire [4-1:0] node10575;
	wire [4-1:0] node10576;
	wire [4-1:0] node10577;
	wire [4-1:0] node10581;
	wire [4-1:0] node10582;
	wire [4-1:0] node10586;
	wire [4-1:0] node10587;
	wire [4-1:0] node10588;
	wire [4-1:0] node10589;
	wire [4-1:0] node10593;
	wire [4-1:0] node10594;
	wire [4-1:0] node10598;
	wire [4-1:0] node10599;
	wire [4-1:0] node10603;
	wire [4-1:0] node10604;
	wire [4-1:0] node10605;
	wire [4-1:0] node10606;
	wire [4-1:0] node10607;
	wire [4-1:0] node10608;
	wire [4-1:0] node10609;
	wire [4-1:0] node10610;
	wire [4-1:0] node10611;
	wire [4-1:0] node10614;
	wire [4-1:0] node10617;
	wire [4-1:0] node10620;
	wire [4-1:0] node10621;
	wire [4-1:0] node10623;
	wire [4-1:0] node10626;
	wire [4-1:0] node10628;
	wire [4-1:0] node10631;
	wire [4-1:0] node10632;
	wire [4-1:0] node10635;
	wire [4-1:0] node10636;
	wire [4-1:0] node10638;
	wire [4-1:0] node10641;
	wire [4-1:0] node10643;
	wire [4-1:0] node10646;
	wire [4-1:0] node10647;
	wire [4-1:0] node10648;
	wire [4-1:0] node10649;
	wire [4-1:0] node10651;
	wire [4-1:0] node10654;
	wire [4-1:0] node10655;
	wire [4-1:0] node10659;
	wire [4-1:0] node10660;
	wire [4-1:0] node10661;
	wire [4-1:0] node10665;
	wire [4-1:0] node10667;
	wire [4-1:0] node10670;
	wire [4-1:0] node10671;
	wire [4-1:0] node10672;
	wire [4-1:0] node10674;
	wire [4-1:0] node10677;
	wire [4-1:0] node10679;
	wire [4-1:0] node10682;
	wire [4-1:0] node10683;
	wire [4-1:0] node10686;
	wire [4-1:0] node10687;
	wire [4-1:0] node10690;
	wire [4-1:0] node10693;
	wire [4-1:0] node10694;
	wire [4-1:0] node10695;
	wire [4-1:0] node10696;
	wire [4-1:0] node10697;
	wire [4-1:0] node10700;
	wire [4-1:0] node10701;
	wire [4-1:0] node10705;
	wire [4-1:0] node10706;
	wire [4-1:0] node10707;
	wire [4-1:0] node10710;
	wire [4-1:0] node10713;
	wire [4-1:0] node10714;
	wire [4-1:0] node10717;
	wire [4-1:0] node10720;
	wire [4-1:0] node10721;
	wire [4-1:0] node10722;
	wire [4-1:0] node10723;
	wire [4-1:0] node10727;
	wire [4-1:0] node10729;
	wire [4-1:0] node10732;
	wire [4-1:0] node10733;
	wire [4-1:0] node10734;
	wire [4-1:0] node10738;
	wire [4-1:0] node10740;
	wire [4-1:0] node10743;
	wire [4-1:0] node10744;
	wire [4-1:0] node10745;
	wire [4-1:0] node10746;
	wire [4-1:0] node10747;
	wire [4-1:0] node10751;
	wire [4-1:0] node10752;
	wire [4-1:0] node10756;
	wire [4-1:0] node10757;
	wire [4-1:0] node10758;
	wire [4-1:0] node10762;
	wire [4-1:0] node10763;
	wire [4-1:0] node10767;
	wire [4-1:0] node10768;
	wire [4-1:0] node10769;
	wire [4-1:0] node10772;
	wire [4-1:0] node10773;
	wire [4-1:0] node10777;
	wire [4-1:0] node10778;
	wire [4-1:0] node10779;
	wire [4-1:0] node10782;
	wire [4-1:0] node10785;
	wire [4-1:0] node10786;
	wire [4-1:0] node10790;
	wire [4-1:0] node10791;
	wire [4-1:0] node10792;
	wire [4-1:0] node10793;
	wire [4-1:0] node10794;
	wire [4-1:0] node10795;
	wire [4-1:0] node10796;
	wire [4-1:0] node10799;
	wire [4-1:0] node10802;
	wire [4-1:0] node10803;
	wire [4-1:0] node10807;
	wire [4-1:0] node10808;
	wire [4-1:0] node10809;
	wire [4-1:0] node10813;
	wire [4-1:0] node10816;
	wire [4-1:0] node10817;
	wire [4-1:0] node10818;
	wire [4-1:0] node10819;
	wire [4-1:0] node10822;
	wire [4-1:0] node10825;
	wire [4-1:0] node10828;
	wire [4-1:0] node10829;
	wire [4-1:0] node10830;
	wire [4-1:0] node10833;
	wire [4-1:0] node10836;
	wire [4-1:0] node10837;
	wire [4-1:0] node10840;
	wire [4-1:0] node10843;
	wire [4-1:0] node10844;
	wire [4-1:0] node10845;
	wire [4-1:0] node10846;
	wire [4-1:0] node10849;
	wire [4-1:0] node10850;
	wire [4-1:0] node10853;
	wire [4-1:0] node10856;
	wire [4-1:0] node10857;
	wire [4-1:0] node10858;
	wire [4-1:0] node10863;
	wire [4-1:0] node10864;
	wire [4-1:0] node10866;
	wire [4-1:0] node10867;
	wire [4-1:0] node10871;
	wire [4-1:0] node10873;
	wire [4-1:0] node10874;
	wire [4-1:0] node10877;
	wire [4-1:0] node10880;
	wire [4-1:0] node10881;
	wire [4-1:0] node10882;
	wire [4-1:0] node10883;
	wire [4-1:0] node10884;
	wire [4-1:0] node10885;
	wire [4-1:0] node10889;
	wire [4-1:0] node10890;
	wire [4-1:0] node10894;
	wire [4-1:0] node10895;
	wire [4-1:0] node10897;
	wire [4-1:0] node10900;
	wire [4-1:0] node10903;
	wire [4-1:0] node10904;
	wire [4-1:0] node10905;
	wire [4-1:0] node10906;
	wire [4-1:0] node10909;
	wire [4-1:0] node10912;
	wire [4-1:0] node10915;
	wire [4-1:0] node10918;
	wire [4-1:0] node10919;
	wire [4-1:0] node10920;
	wire [4-1:0] node10921;
	wire [4-1:0] node10922;
	wire [4-1:0] node10927;
	wire [4-1:0] node10928;
	wire [4-1:0] node10929;
	wire [4-1:0] node10934;
	wire [4-1:0] node10935;
	wire [4-1:0] node10936;
	wire [4-1:0] node10937;
	wire [4-1:0] node10940;
	wire [4-1:0] node10943;
	wire [4-1:0] node10946;
	wire [4-1:0] node10947;
	wire [4-1:0] node10948;
	wire [4-1:0] node10952;
	wire [4-1:0] node10953;
	wire [4-1:0] node10957;
	wire [4-1:0] node10958;
	wire [4-1:0] node10959;
	wire [4-1:0] node10960;
	wire [4-1:0] node10961;
	wire [4-1:0] node10962;
	wire [4-1:0] node10963;
	wire [4-1:0] node10964;
	wire [4-1:0] node10968;
	wire [4-1:0] node10971;
	wire [4-1:0] node10972;
	wire [4-1:0] node10974;
	wire [4-1:0] node10978;
	wire [4-1:0] node10979;
	wire [4-1:0] node10980;
	wire [4-1:0] node10983;
	wire [4-1:0] node10984;
	wire [4-1:0] node10988;
	wire [4-1:0] node10989;
	wire [4-1:0] node10991;
	wire [4-1:0] node10994;
	wire [4-1:0] node10995;
	wire [4-1:0] node10999;
	wire [4-1:0] node11000;
	wire [4-1:0] node11001;
	wire [4-1:0] node11002;
	wire [4-1:0] node11004;
	wire [4-1:0] node11007;
	wire [4-1:0] node11008;
	wire [4-1:0] node11012;
	wire [4-1:0] node11013;
	wire [4-1:0] node11015;
	wire [4-1:0] node11018;
	wire [4-1:0] node11021;
	wire [4-1:0] node11022;
	wire [4-1:0] node11023;
	wire [4-1:0] node11024;
	wire [4-1:0] node11028;
	wire [4-1:0] node11029;
	wire [4-1:0] node11033;
	wire [4-1:0] node11034;
	wire [4-1:0] node11035;
	wire [4-1:0] node11039;
	wire [4-1:0] node11040;
	wire [4-1:0] node11044;
	wire [4-1:0] node11045;
	wire [4-1:0] node11046;
	wire [4-1:0] node11047;
	wire [4-1:0] node11049;
	wire [4-1:0] node11052;
	wire [4-1:0] node11053;
	wire [4-1:0] node11054;
	wire [4-1:0] node11058;
	wire [4-1:0] node11059;
	wire [4-1:0] node11063;
	wire [4-1:0] node11064;
	wire [4-1:0] node11065;
	wire [4-1:0] node11067;
	wire [4-1:0] node11071;
	wire [4-1:0] node11072;
	wire [4-1:0] node11076;
	wire [4-1:0] node11077;
	wire [4-1:0] node11078;
	wire [4-1:0] node11079;
	wire [4-1:0] node11080;
	wire [4-1:0] node11083;
	wire [4-1:0] node11086;
	wire [4-1:0] node11087;
	wire [4-1:0] node11091;
	wire [4-1:0] node11092;
	wire [4-1:0] node11093;
	wire [4-1:0] node11097;
	wire [4-1:0] node11098;
	wire [4-1:0] node11101;
	wire [4-1:0] node11104;
	wire [4-1:0] node11105;
	wire [4-1:0] node11107;
	wire [4-1:0] node11108;
	wire [4-1:0] node11111;
	wire [4-1:0] node11114;
	wire [4-1:0] node11115;
	wire [4-1:0] node11116;
	wire [4-1:0] node11121;
	wire [4-1:0] node11122;
	wire [4-1:0] node11123;
	wire [4-1:0] node11124;
	wire [4-1:0] node11125;
	wire [4-1:0] node11126;
	wire [4-1:0] node11128;
	wire [4-1:0] node11132;
	wire [4-1:0] node11134;
	wire [4-1:0] node11135;
	wire [4-1:0] node11139;
	wire [4-1:0] node11140;
	wire [4-1:0] node11142;
	wire [4-1:0] node11143;
	wire [4-1:0] node11147;
	wire [4-1:0] node11148;
	wire [4-1:0] node11151;
	wire [4-1:0] node11153;
	wire [4-1:0] node11156;
	wire [4-1:0] node11157;
	wire [4-1:0] node11158;
	wire [4-1:0] node11160;
	wire [4-1:0] node11161;
	wire [4-1:0] node11165;
	wire [4-1:0] node11166;
	wire [4-1:0] node11167;
	wire [4-1:0] node11170;
	wire [4-1:0] node11173;
	wire [4-1:0] node11174;
	wire [4-1:0] node11178;
	wire [4-1:0] node11179;
	wire [4-1:0] node11180;
	wire [4-1:0] node11181;
	wire [4-1:0] node11184;
	wire [4-1:0] node11187;
	wire [4-1:0] node11188;
	wire [4-1:0] node11192;
	wire [4-1:0] node11193;
	wire [4-1:0] node11196;
	wire [4-1:0] node11199;
	wire [4-1:0] node11200;
	wire [4-1:0] node11201;
	wire [4-1:0] node11202;
	wire [4-1:0] node11203;
	wire [4-1:0] node11205;
	wire [4-1:0] node11208;
	wire [4-1:0] node11209;
	wire [4-1:0] node11212;
	wire [4-1:0] node11215;
	wire [4-1:0] node11216;
	wire [4-1:0] node11219;
	wire [4-1:0] node11220;
	wire [4-1:0] node11224;
	wire [4-1:0] node11225;
	wire [4-1:0] node11226;
	wire [4-1:0] node11229;
	wire [4-1:0] node11232;
	wire [4-1:0] node11234;
	wire [4-1:0] node11235;
	wire [4-1:0] node11239;
	wire [4-1:0] node11240;
	wire [4-1:0] node11241;
	wire [4-1:0] node11242;
	wire [4-1:0] node11246;
	wire [4-1:0] node11247;
	wire [4-1:0] node11248;
	wire [4-1:0] node11251;
	wire [4-1:0] node11255;
	wire [4-1:0] node11256;
	wire [4-1:0] node11258;
	wire [4-1:0] node11261;
	wire [4-1:0] node11262;
	wire [4-1:0] node11263;
	wire [4-1:0] node11267;
	wire [4-1:0] node11270;
	wire [4-1:0] node11271;
	wire [4-1:0] node11272;
	wire [4-1:0] node11273;
	wire [4-1:0] node11274;
	wire [4-1:0] node11275;
	wire [4-1:0] node11276;
	wire [4-1:0] node11277;
	wire [4-1:0] node11278;
	wire [4-1:0] node11279;
	wire [4-1:0] node11280;
	wire [4-1:0] node11281;
	wire [4-1:0] node11282;
	wire [4-1:0] node11286;
	wire [4-1:0] node11288;
	wire [4-1:0] node11291;
	wire [4-1:0] node11292;
	wire [4-1:0] node11293;
	wire [4-1:0] node11297;
	wire [4-1:0] node11298;
	wire [4-1:0] node11301;
	wire [4-1:0] node11304;
	wire [4-1:0] node11305;
	wire [4-1:0] node11306;
	wire [4-1:0] node11307;
	wire [4-1:0] node11311;
	wire [4-1:0] node11313;
	wire [4-1:0] node11316;
	wire [4-1:0] node11317;
	wire [4-1:0] node11318;
	wire [4-1:0] node11323;
	wire [4-1:0] node11324;
	wire [4-1:0] node11325;
	wire [4-1:0] node11326;
	wire [4-1:0] node11327;
	wire [4-1:0] node11331;
	wire [4-1:0] node11333;
	wire [4-1:0] node11336;
	wire [4-1:0] node11337;
	wire [4-1:0] node11339;
	wire [4-1:0] node11342;
	wire [4-1:0] node11345;
	wire [4-1:0] node11346;
	wire [4-1:0] node11347;
	wire [4-1:0] node11348;
	wire [4-1:0] node11352;
	wire [4-1:0] node11355;
	wire [4-1:0] node11356;
	wire [4-1:0] node11358;
	wire [4-1:0] node11362;
	wire [4-1:0] node11363;
	wire [4-1:0] node11364;
	wire [4-1:0] node11365;
	wire [4-1:0] node11366;
	wire [4-1:0] node11369;
	wire [4-1:0] node11371;
	wire [4-1:0] node11374;
	wire [4-1:0] node11375;
	wire [4-1:0] node11376;
	wire [4-1:0] node11380;
	wire [4-1:0] node11381;
	wire [4-1:0] node11384;
	wire [4-1:0] node11387;
	wire [4-1:0] node11388;
	wire [4-1:0] node11389;
	wire [4-1:0] node11391;
	wire [4-1:0] node11394;
	wire [4-1:0] node11396;
	wire [4-1:0] node11399;
	wire [4-1:0] node11400;
	wire [4-1:0] node11402;
	wire [4-1:0] node11405;
	wire [4-1:0] node11408;
	wire [4-1:0] node11409;
	wire [4-1:0] node11410;
	wire [4-1:0] node11411;
	wire [4-1:0] node11414;
	wire [4-1:0] node11415;
	wire [4-1:0] node11419;
	wire [4-1:0] node11421;
	wire [4-1:0] node11424;
	wire [4-1:0] node11425;
	wire [4-1:0] node11426;
	wire [4-1:0] node11427;
	wire [4-1:0] node11431;
	wire [4-1:0] node11432;
	wire [4-1:0] node11436;
	wire [4-1:0] node11437;
	wire [4-1:0] node11438;
	wire [4-1:0] node11441;
	wire [4-1:0] node11444;
	wire [4-1:0] node11445;
	wire [4-1:0] node11449;
	wire [4-1:0] node11450;
	wire [4-1:0] node11451;
	wire [4-1:0] node11452;
	wire [4-1:0] node11453;
	wire [4-1:0] node11454;
	wire [4-1:0] node11455;
	wire [4-1:0] node11459;
	wire [4-1:0] node11460;
	wire [4-1:0] node11464;
	wire [4-1:0] node11465;
	wire [4-1:0] node11467;
	wire [4-1:0] node11470;
	wire [4-1:0] node11471;
	wire [4-1:0] node11474;
	wire [4-1:0] node11477;
	wire [4-1:0] node11478;
	wire [4-1:0] node11479;
	wire [4-1:0] node11481;
	wire [4-1:0] node11484;
	wire [4-1:0] node11485;
	wire [4-1:0] node11489;
	wire [4-1:0] node11491;
	wire [4-1:0] node11493;
	wire [4-1:0] node11496;
	wire [4-1:0] node11497;
	wire [4-1:0] node11498;
	wire [4-1:0] node11499;
	wire [4-1:0] node11500;
	wire [4-1:0] node11503;
	wire [4-1:0] node11506;
	wire [4-1:0] node11508;
	wire [4-1:0] node11511;
	wire [4-1:0] node11512;
	wire [4-1:0] node11513;
	wire [4-1:0] node11518;
	wire [4-1:0] node11519;
	wire [4-1:0] node11520;
	wire [4-1:0] node11521;
	wire [4-1:0] node11525;
	wire [4-1:0] node11528;
	wire [4-1:0] node11529;
	wire [4-1:0] node11531;
	wire [4-1:0] node11534;
	wire [4-1:0] node11535;
	wire [4-1:0] node11539;
	wire [4-1:0] node11540;
	wire [4-1:0] node11541;
	wire [4-1:0] node11542;
	wire [4-1:0] node11543;
	wire [4-1:0] node11544;
	wire [4-1:0] node11547;
	wire [4-1:0] node11550;
	wire [4-1:0] node11553;
	wire [4-1:0] node11554;
	wire [4-1:0] node11556;
	wire [4-1:0] node11559;
	wire [4-1:0] node11560;
	wire [4-1:0] node11564;
	wire [4-1:0] node11565;
	wire [4-1:0] node11567;
	wire [4-1:0] node11569;
	wire [4-1:0] node11572;
	wire [4-1:0] node11573;
	wire [4-1:0] node11576;
	wire [4-1:0] node11578;
	wire [4-1:0] node11581;
	wire [4-1:0] node11582;
	wire [4-1:0] node11583;
	wire [4-1:0] node11584;
	wire [4-1:0] node11585;
	wire [4-1:0] node11589;
	wire [4-1:0] node11591;
	wire [4-1:0] node11594;
	wire [4-1:0] node11595;
	wire [4-1:0] node11597;
	wire [4-1:0] node11600;
	wire [4-1:0] node11601;
	wire [4-1:0] node11605;
	wire [4-1:0] node11606;
	wire [4-1:0] node11607;
	wire [4-1:0] node11608;
	wire [4-1:0] node11612;
	wire [4-1:0] node11613;
	wire [4-1:0] node11617;
	wire [4-1:0] node11618;
	wire [4-1:0] node11619;
	wire [4-1:0] node11624;
	wire [4-1:0] node11625;
	wire [4-1:0] node11626;
	wire [4-1:0] node11627;
	wire [4-1:0] node11628;
	wire [4-1:0] node11629;
	wire [4-1:0] node11630;
	wire [4-1:0] node11631;
	wire [4-1:0] node11634;
	wire [4-1:0] node11637;
	wire [4-1:0] node11638;
	wire [4-1:0] node11641;
	wire [4-1:0] node11644;
	wire [4-1:0] node11645;
	wire [4-1:0] node11648;
	wire [4-1:0] node11650;
	wire [4-1:0] node11653;
	wire [4-1:0] node11654;
	wire [4-1:0] node11655;
	wire [4-1:0] node11656;
	wire [4-1:0] node11659;
	wire [4-1:0] node11662;
	wire [4-1:0] node11663;
	wire [4-1:0] node11667;
	wire [4-1:0] node11668;
	wire [4-1:0] node11671;
	wire [4-1:0] node11673;
	wire [4-1:0] node11676;
	wire [4-1:0] node11677;
	wire [4-1:0] node11678;
	wire [4-1:0] node11679;
	wire [4-1:0] node11682;
	wire [4-1:0] node11684;
	wire [4-1:0] node11687;
	wire [4-1:0] node11688;
	wire [4-1:0] node11689;
	wire [4-1:0] node11692;
	wire [4-1:0] node11695;
	wire [4-1:0] node11696;
	wire [4-1:0] node11699;
	wire [4-1:0] node11702;
	wire [4-1:0] node11703;
	wire [4-1:0] node11704;
	wire [4-1:0] node11706;
	wire [4-1:0] node11709;
	wire [4-1:0] node11711;
	wire [4-1:0] node11714;
	wire [4-1:0] node11715;
	wire [4-1:0] node11716;
	wire [4-1:0] node11719;
	wire [4-1:0] node11722;
	wire [4-1:0] node11723;
	wire [4-1:0] node11726;
	wire [4-1:0] node11729;
	wire [4-1:0] node11730;
	wire [4-1:0] node11731;
	wire [4-1:0] node11732;
	wire [4-1:0] node11733;
	wire [4-1:0] node11734;
	wire [4-1:0] node11738;
	wire [4-1:0] node11740;
	wire [4-1:0] node11743;
	wire [4-1:0] node11744;
	wire [4-1:0] node11746;
	wire [4-1:0] node11749;
	wire [4-1:0] node11751;
	wire [4-1:0] node11754;
	wire [4-1:0] node11755;
	wire [4-1:0] node11756;
	wire [4-1:0] node11757;
	wire [4-1:0] node11760;
	wire [4-1:0] node11763;
	wire [4-1:0] node11764;
	wire [4-1:0] node11767;
	wire [4-1:0] node11770;
	wire [4-1:0] node11771;
	wire [4-1:0] node11772;
	wire [4-1:0] node11776;
	wire [4-1:0] node11777;
	wire [4-1:0] node11780;
	wire [4-1:0] node11783;
	wire [4-1:0] node11784;
	wire [4-1:0] node11785;
	wire [4-1:0] node11786;
	wire [4-1:0] node11787;
	wire [4-1:0] node11791;
	wire [4-1:0] node11793;
	wire [4-1:0] node11796;
	wire [4-1:0] node11797;
	wire [4-1:0] node11798;
	wire [4-1:0] node11802;
	wire [4-1:0] node11803;
	wire [4-1:0] node11807;
	wire [4-1:0] node11808;
	wire [4-1:0] node11809;
	wire [4-1:0] node11810;
	wire [4-1:0] node11814;
	wire [4-1:0] node11815;
	wire [4-1:0] node11819;
	wire [4-1:0] node11820;
	wire [4-1:0] node11821;
	wire [4-1:0] node11825;
	wire [4-1:0] node11828;
	wire [4-1:0] node11829;
	wire [4-1:0] node11830;
	wire [4-1:0] node11831;
	wire [4-1:0] node11832;
	wire [4-1:0] node11833;
	wire [4-1:0] node11835;
	wire [4-1:0] node11838;
	wire [4-1:0] node11840;
	wire [4-1:0] node11843;
	wire [4-1:0] node11844;
	wire [4-1:0] node11847;
	wire [4-1:0] node11849;
	wire [4-1:0] node11852;
	wire [4-1:0] node11853;
	wire [4-1:0] node11854;
	wire [4-1:0] node11855;
	wire [4-1:0] node11859;
	wire [4-1:0] node11860;
	wire [4-1:0] node11864;
	wire [4-1:0] node11865;
	wire [4-1:0] node11869;
	wire [4-1:0] node11870;
	wire [4-1:0] node11871;
	wire [4-1:0] node11872;
	wire [4-1:0] node11874;
	wire [4-1:0] node11877;
	wire [4-1:0] node11878;
	wire [4-1:0] node11882;
	wire [4-1:0] node11883;
	wire [4-1:0] node11886;
	wire [4-1:0] node11887;
	wire [4-1:0] node11890;
	wire [4-1:0] node11893;
	wire [4-1:0] node11894;
	wire [4-1:0] node11895;
	wire [4-1:0] node11897;
	wire [4-1:0] node11900;
	wire [4-1:0] node11901;
	wire [4-1:0] node11904;
	wire [4-1:0] node11907;
	wire [4-1:0] node11908;
	wire [4-1:0] node11909;
	wire [4-1:0] node11913;
	wire [4-1:0] node11914;
	wire [4-1:0] node11918;
	wire [4-1:0] node11919;
	wire [4-1:0] node11920;
	wire [4-1:0] node11921;
	wire [4-1:0] node11922;
	wire [4-1:0] node11924;
	wire [4-1:0] node11927;
	wire [4-1:0] node11928;
	wire [4-1:0] node11932;
	wire [4-1:0] node11933;
	wire [4-1:0] node11936;
	wire [4-1:0] node11939;
	wire [4-1:0] node11940;
	wire [4-1:0] node11941;
	wire [4-1:0] node11944;
	wire [4-1:0] node11947;
	wire [4-1:0] node11948;
	wire [4-1:0] node11949;
	wire [4-1:0] node11952;
	wire [4-1:0] node11955;
	wire [4-1:0] node11956;
	wire [4-1:0] node11960;
	wire [4-1:0] node11961;
	wire [4-1:0] node11962;
	wire [4-1:0] node11963;
	wire [4-1:0] node11964;
	wire [4-1:0] node11968;
	wire [4-1:0] node11971;
	wire [4-1:0] node11972;
	wire [4-1:0] node11975;
	wire [4-1:0] node11976;
	wire [4-1:0] node11980;
	wire [4-1:0] node11981;
	wire [4-1:0] node11982;
	wire [4-1:0] node11983;
	wire [4-1:0] node11987;
	wire [4-1:0] node11988;
	wire [4-1:0] node11992;
	wire [4-1:0] node11993;
	wire [4-1:0] node11994;
	wire [4-1:0] node11998;
	wire [4-1:0] node12001;
	wire [4-1:0] node12002;
	wire [4-1:0] node12003;
	wire [4-1:0] node12004;
	wire [4-1:0] node12005;
	wire [4-1:0] node12006;
	wire [4-1:0] node12007;
	wire [4-1:0] node12008;
	wire [4-1:0] node12011;
	wire [4-1:0] node12013;
	wire [4-1:0] node12016;
	wire [4-1:0] node12017;
	wire [4-1:0] node12019;
	wire [4-1:0] node12023;
	wire [4-1:0] node12024;
	wire [4-1:0] node12025;
	wire [4-1:0] node12026;
	wire [4-1:0] node12029;
	wire [4-1:0] node12032;
	wire [4-1:0] node12033;
	wire [4-1:0] node12036;
	wire [4-1:0] node12039;
	wire [4-1:0] node12040;
	wire [4-1:0] node12041;
	wire [4-1:0] node12044;
	wire [4-1:0] node12047;
	wire [4-1:0] node12050;
	wire [4-1:0] node12051;
	wire [4-1:0] node12052;
	wire [4-1:0] node12054;
	wire [4-1:0] node12055;
	wire [4-1:0] node12058;
	wire [4-1:0] node12061;
	wire [4-1:0] node12062;
	wire [4-1:0] node12064;
	wire [4-1:0] node12067;
	wire [4-1:0] node12069;
	wire [4-1:0] node12072;
	wire [4-1:0] node12073;
	wire [4-1:0] node12075;
	wire [4-1:0] node12078;
	wire [4-1:0] node12079;
	wire [4-1:0] node12081;
	wire [4-1:0] node12085;
	wire [4-1:0] node12086;
	wire [4-1:0] node12087;
	wire [4-1:0] node12088;
	wire [4-1:0] node12089;
	wire [4-1:0] node12090;
	wire [4-1:0] node12094;
	wire [4-1:0] node12097;
	wire [4-1:0] node12098;
	wire [4-1:0] node12099;
	wire [4-1:0] node12102;
	wire [4-1:0] node12105;
	wire [4-1:0] node12107;
	wire [4-1:0] node12110;
	wire [4-1:0] node12111;
	wire [4-1:0] node12112;
	wire [4-1:0] node12113;
	wire [4-1:0] node12116;
	wire [4-1:0] node12119;
	wire [4-1:0] node12122;
	wire [4-1:0] node12123;
	wire [4-1:0] node12125;
	wire [4-1:0] node12128;
	wire [4-1:0] node12129;
	wire [4-1:0] node12132;
	wire [4-1:0] node12135;
	wire [4-1:0] node12136;
	wire [4-1:0] node12137;
	wire [4-1:0] node12138;
	wire [4-1:0] node12139;
	wire [4-1:0] node12143;
	wire [4-1:0] node12144;
	wire [4-1:0] node12148;
	wire [4-1:0] node12149;
	wire [4-1:0] node12150;
	wire [4-1:0] node12154;
	wire [4-1:0] node12156;
	wire [4-1:0] node12159;
	wire [4-1:0] node12160;
	wire [4-1:0] node12161;
	wire [4-1:0] node12163;
	wire [4-1:0] node12166;
	wire [4-1:0] node12167;
	wire [4-1:0] node12170;
	wire [4-1:0] node12173;
	wire [4-1:0] node12174;
	wire [4-1:0] node12175;
	wire [4-1:0] node12179;
	wire [4-1:0] node12182;
	wire [4-1:0] node12183;
	wire [4-1:0] node12184;
	wire [4-1:0] node12185;
	wire [4-1:0] node12186;
	wire [4-1:0] node12187;
	wire [4-1:0] node12188;
	wire [4-1:0] node12191;
	wire [4-1:0] node12194;
	wire [4-1:0] node12195;
	wire [4-1:0] node12199;
	wire [4-1:0] node12200;
	wire [4-1:0] node12201;
	wire [4-1:0] node12204;
	wire [4-1:0] node12207;
	wire [4-1:0] node12209;
	wire [4-1:0] node12212;
	wire [4-1:0] node12213;
	wire [4-1:0] node12214;
	wire [4-1:0] node12215;
	wire [4-1:0] node12218;
	wire [4-1:0] node12221;
	wire [4-1:0] node12223;
	wire [4-1:0] node12226;
	wire [4-1:0] node12227;
	wire [4-1:0] node12228;
	wire [4-1:0] node12231;
	wire [4-1:0] node12234;
	wire [4-1:0] node12236;
	wire [4-1:0] node12239;
	wire [4-1:0] node12240;
	wire [4-1:0] node12241;
	wire [4-1:0] node12242;
	wire [4-1:0] node12245;
	wire [4-1:0] node12246;
	wire [4-1:0] node12250;
	wire [4-1:0] node12251;
	wire [4-1:0] node12254;
	wire [4-1:0] node12256;
	wire [4-1:0] node12259;
	wire [4-1:0] node12260;
	wire [4-1:0] node12261;
	wire [4-1:0] node12263;
	wire [4-1:0] node12266;
	wire [4-1:0] node12267;
	wire [4-1:0] node12270;
	wire [4-1:0] node12273;
	wire [4-1:0] node12275;
	wire [4-1:0] node12278;
	wire [4-1:0] node12279;
	wire [4-1:0] node12280;
	wire [4-1:0] node12281;
	wire [4-1:0] node12283;
	wire [4-1:0] node12285;
	wire [4-1:0] node12288;
	wire [4-1:0] node12290;
	wire [4-1:0] node12291;
	wire [4-1:0] node12294;
	wire [4-1:0] node12297;
	wire [4-1:0] node12298;
	wire [4-1:0] node12299;
	wire [4-1:0] node12301;
	wire [4-1:0] node12304;
	wire [4-1:0] node12305;
	wire [4-1:0] node12308;
	wire [4-1:0] node12311;
	wire [4-1:0] node12312;
	wire [4-1:0] node12315;
	wire [4-1:0] node12316;
	wire [4-1:0] node12320;
	wire [4-1:0] node12321;
	wire [4-1:0] node12322;
	wire [4-1:0] node12324;
	wire [4-1:0] node12326;
	wire [4-1:0] node12329;
	wire [4-1:0] node12330;
	wire [4-1:0] node12333;
	wire [4-1:0] node12334;
	wire [4-1:0] node12337;
	wire [4-1:0] node12340;
	wire [4-1:0] node12341;
	wire [4-1:0] node12342;
	wire [4-1:0] node12344;
	wire [4-1:0] node12347;
	wire [4-1:0] node12348;
	wire [4-1:0] node12352;
	wire [4-1:0] node12353;
	wire [4-1:0] node12355;
	wire [4-1:0] node12358;
	wire [4-1:0] node12361;
	wire [4-1:0] node12362;
	wire [4-1:0] node12363;
	wire [4-1:0] node12364;
	wire [4-1:0] node12365;
	wire [4-1:0] node12366;
	wire [4-1:0] node12367;
	wire [4-1:0] node12368;
	wire [4-1:0] node12372;
	wire [4-1:0] node12373;
	wire [4-1:0] node12377;
	wire [4-1:0] node12378;
	wire [4-1:0] node12380;
	wire [4-1:0] node12384;
	wire [4-1:0] node12385;
	wire [4-1:0] node12386;
	wire [4-1:0] node12389;
	wire [4-1:0] node12390;
	wire [4-1:0] node12394;
	wire [4-1:0] node12396;
	wire [4-1:0] node12397;
	wire [4-1:0] node12400;
	wire [4-1:0] node12403;
	wire [4-1:0] node12404;
	wire [4-1:0] node12405;
	wire [4-1:0] node12407;
	wire [4-1:0] node12408;
	wire [4-1:0] node12411;
	wire [4-1:0] node12414;
	wire [4-1:0] node12415;
	wire [4-1:0] node12416;
	wire [4-1:0] node12420;
	wire [4-1:0] node12421;
	wire [4-1:0] node12424;
	wire [4-1:0] node12427;
	wire [4-1:0] node12428;
	wire [4-1:0] node12429;
	wire [4-1:0] node12430;
	wire [4-1:0] node12434;
	wire [4-1:0] node12436;
	wire [4-1:0] node12439;
	wire [4-1:0] node12440;
	wire [4-1:0] node12441;
	wire [4-1:0] node12445;
	wire [4-1:0] node12447;
	wire [4-1:0] node12450;
	wire [4-1:0] node12451;
	wire [4-1:0] node12452;
	wire [4-1:0] node12453;
	wire [4-1:0] node12454;
	wire [4-1:0] node12457;
	wire [4-1:0] node12458;
	wire [4-1:0] node12462;
	wire [4-1:0] node12464;
	wire [4-1:0] node12467;
	wire [4-1:0] node12468;
	wire [4-1:0] node12469;
	wire [4-1:0] node12470;
	wire [4-1:0] node12474;
	wire [4-1:0] node12475;
	wire [4-1:0] node12479;
	wire [4-1:0] node12481;
	wire [4-1:0] node12484;
	wire [4-1:0] node12485;
	wire [4-1:0] node12486;
	wire [4-1:0] node12488;
	wire [4-1:0] node12490;
	wire [4-1:0] node12493;
	wire [4-1:0] node12494;
	wire [4-1:0] node12496;
	wire [4-1:0] node12499;
	wire [4-1:0] node12502;
	wire [4-1:0] node12503;
	wire [4-1:0] node12504;
	wire [4-1:0] node12505;
	wire [4-1:0] node12509;
	wire [4-1:0] node12510;
	wire [4-1:0] node12514;
	wire [4-1:0] node12516;
	wire [4-1:0] node12517;
	wire [4-1:0] node12521;
	wire [4-1:0] node12522;
	wire [4-1:0] node12523;
	wire [4-1:0] node12524;
	wire [4-1:0] node12525;
	wire [4-1:0] node12526;
	wire [4-1:0] node12527;
	wire [4-1:0] node12530;
	wire [4-1:0] node12533;
	wire [4-1:0] node12536;
	wire [4-1:0] node12537;
	wire [4-1:0] node12538;
	wire [4-1:0] node12542;
	wire [4-1:0] node12544;
	wire [4-1:0] node12547;
	wire [4-1:0] node12548;
	wire [4-1:0] node12549;
	wire [4-1:0] node12550;
	wire [4-1:0] node12553;
	wire [4-1:0] node12556;
	wire [4-1:0] node12558;
	wire [4-1:0] node12561;
	wire [4-1:0] node12562;
	wire [4-1:0] node12565;
	wire [4-1:0] node12566;
	wire [4-1:0] node12570;
	wire [4-1:0] node12571;
	wire [4-1:0] node12572;
	wire [4-1:0] node12573;
	wire [4-1:0] node12575;
	wire [4-1:0] node12579;
	wire [4-1:0] node12580;
	wire [4-1:0] node12583;
	wire [4-1:0] node12584;
	wire [4-1:0] node12587;
	wire [4-1:0] node12590;
	wire [4-1:0] node12591;
	wire [4-1:0] node12592;
	wire [4-1:0] node12595;
	wire [4-1:0] node12597;
	wire [4-1:0] node12600;
	wire [4-1:0] node12601;
	wire [4-1:0] node12602;
	wire [4-1:0] node12605;
	wire [4-1:0] node12609;
	wire [4-1:0] node12610;
	wire [4-1:0] node12611;
	wire [4-1:0] node12612;
	wire [4-1:0] node12613;
	wire [4-1:0] node12614;
	wire [4-1:0] node12618;
	wire [4-1:0] node12620;
	wire [4-1:0] node12623;
	wire [4-1:0] node12624;
	wire [4-1:0] node12626;
	wire [4-1:0] node12629;
	wire [4-1:0] node12631;
	wire [4-1:0] node12634;
	wire [4-1:0] node12635;
	wire [4-1:0] node12636;
	wire [4-1:0] node12639;
	wire [4-1:0] node12642;
	wire [4-1:0] node12643;
	wire [4-1:0] node12646;
	wire [4-1:0] node12648;
	wire [4-1:0] node12651;
	wire [4-1:0] node12652;
	wire [4-1:0] node12653;
	wire [4-1:0] node12654;
	wire [4-1:0] node12655;
	wire [4-1:0] node12659;
	wire [4-1:0] node12661;
	wire [4-1:0] node12664;
	wire [4-1:0] node12665;
	wire [4-1:0] node12666;
	wire [4-1:0] node12669;
	wire [4-1:0] node12672;
	wire [4-1:0] node12674;
	wire [4-1:0] node12677;
	wire [4-1:0] node12678;
	wire [4-1:0] node12679;
	wire [4-1:0] node12680;
	wire [4-1:0] node12685;
	wire [4-1:0] node12686;
	wire [4-1:0] node12688;
	wire [4-1:0] node12692;
	wire [4-1:0] node12693;
	wire [4-1:0] node12694;
	wire [4-1:0] node12695;
	wire [4-1:0] node12696;
	wire [4-1:0] node12697;
	wire [4-1:0] node12698;
	wire [4-1:0] node12699;
	wire [4-1:0] node12700;
	wire [4-1:0] node12701;
	wire [4-1:0] node12704;
	wire [4-1:0] node12707;
	wire [4-1:0] node12709;
	wire [4-1:0] node12712;
	wire [4-1:0] node12713;
	wire [4-1:0] node12714;
	wire [4-1:0] node12717;
	wire [4-1:0] node12720;
	wire [4-1:0] node12721;
	wire [4-1:0] node12725;
	wire [4-1:0] node12726;
	wire [4-1:0] node12727;
	wire [4-1:0] node12728;
	wire [4-1:0] node12731;
	wire [4-1:0] node12734;
	wire [4-1:0] node12735;
	wire [4-1:0] node12739;
	wire [4-1:0] node12740;
	wire [4-1:0] node12741;
	wire [4-1:0] node12744;
	wire [4-1:0] node12747;
	wire [4-1:0] node12749;
	wire [4-1:0] node12752;
	wire [4-1:0] node12753;
	wire [4-1:0] node12754;
	wire [4-1:0] node12755;
	wire [4-1:0] node12756;
	wire [4-1:0] node12759;
	wire [4-1:0] node12762;
	wire [4-1:0] node12764;
	wire [4-1:0] node12767;
	wire [4-1:0] node12768;
	wire [4-1:0] node12770;
	wire [4-1:0] node12773;
	wire [4-1:0] node12776;
	wire [4-1:0] node12777;
	wire [4-1:0] node12778;
	wire [4-1:0] node12781;
	wire [4-1:0] node12784;
	wire [4-1:0] node12785;
	wire [4-1:0] node12788;
	wire [4-1:0] node12790;
	wire [4-1:0] node12793;
	wire [4-1:0] node12794;
	wire [4-1:0] node12795;
	wire [4-1:0] node12796;
	wire [4-1:0] node12797;
	wire [4-1:0] node12799;
	wire [4-1:0] node12802;
	wire [4-1:0] node12804;
	wire [4-1:0] node12807;
	wire [4-1:0] node12808;
	wire [4-1:0] node12809;
	wire [4-1:0] node12812;
	wire [4-1:0] node12815;
	wire [4-1:0] node12817;
	wire [4-1:0] node12820;
	wire [4-1:0] node12821;
	wire [4-1:0] node12822;
	wire [4-1:0] node12823;
	wire [4-1:0] node12827;
	wire [4-1:0] node12828;
	wire [4-1:0] node12832;
	wire [4-1:0] node12834;
	wire [4-1:0] node12837;
	wire [4-1:0] node12838;
	wire [4-1:0] node12839;
	wire [4-1:0] node12841;
	wire [4-1:0] node12843;
	wire [4-1:0] node12846;
	wire [4-1:0] node12848;
	wire [4-1:0] node12849;
	wire [4-1:0] node12852;
	wire [4-1:0] node12855;
	wire [4-1:0] node12856;
	wire [4-1:0] node12857;
	wire [4-1:0] node12860;
	wire [4-1:0] node12863;
	wire [4-1:0] node12864;
	wire [4-1:0] node12868;
	wire [4-1:0] node12869;
	wire [4-1:0] node12870;
	wire [4-1:0] node12871;
	wire [4-1:0] node12872;
	wire [4-1:0] node12873;
	wire [4-1:0] node12874;
	wire [4-1:0] node12878;
	wire [4-1:0] node12881;
	wire [4-1:0] node12882;
	wire [4-1:0] node12885;
	wire [4-1:0] node12887;
	wire [4-1:0] node12890;
	wire [4-1:0] node12891;
	wire [4-1:0] node12892;
	wire [4-1:0] node12894;
	wire [4-1:0] node12897;
	wire [4-1:0] node12898;
	wire [4-1:0] node12901;
	wire [4-1:0] node12904;
	wire [4-1:0] node12906;
	wire [4-1:0] node12908;
	wire [4-1:0] node12911;
	wire [4-1:0] node12912;
	wire [4-1:0] node12913;
	wire [4-1:0] node12914;
	wire [4-1:0] node12916;
	wire [4-1:0] node12919;
	wire [4-1:0] node12921;
	wire [4-1:0] node12924;
	wire [4-1:0] node12925;
	wire [4-1:0] node12927;
	wire [4-1:0] node12930;
	wire [4-1:0] node12932;
	wire [4-1:0] node12935;
	wire [4-1:0] node12936;
	wire [4-1:0] node12937;
	wire [4-1:0] node12940;
	wire [4-1:0] node12941;
	wire [4-1:0] node12945;
	wire [4-1:0] node12946;
	wire [4-1:0] node12947;
	wire [4-1:0] node12950;
	wire [4-1:0] node12953;
	wire [4-1:0] node12956;
	wire [4-1:0] node12957;
	wire [4-1:0] node12958;
	wire [4-1:0] node12959;
	wire [4-1:0] node12960;
	wire [4-1:0] node12962;
	wire [4-1:0] node12965;
	wire [4-1:0] node12968;
	wire [4-1:0] node12969;
	wire [4-1:0] node12970;
	wire [4-1:0] node12974;
	wire [4-1:0] node12975;
	wire [4-1:0] node12978;
	wire [4-1:0] node12981;
	wire [4-1:0] node12982;
	wire [4-1:0] node12983;
	wire [4-1:0] node12986;
	wire [4-1:0] node12989;
	wire [4-1:0] node12990;
	wire [4-1:0] node12993;
	wire [4-1:0] node12995;
	wire [4-1:0] node12998;
	wire [4-1:0] node12999;
	wire [4-1:0] node13000;
	wire [4-1:0] node13001;
	wire [4-1:0] node13003;
	wire [4-1:0] node13006;
	wire [4-1:0] node13008;
	wire [4-1:0] node13011;
	wire [4-1:0] node13012;
	wire [4-1:0] node13015;
	wire [4-1:0] node13016;
	wire [4-1:0] node13019;
	wire [4-1:0] node13022;
	wire [4-1:0] node13023;
	wire [4-1:0] node13024;
	wire [4-1:0] node13025;
	wire [4-1:0] node13028;
	wire [4-1:0] node13032;
	wire [4-1:0] node13034;
	wire [4-1:0] node13037;
	wire [4-1:0] node13038;
	wire [4-1:0] node13039;
	wire [4-1:0] node13040;
	wire [4-1:0] node13041;
	wire [4-1:0] node13042;
	wire [4-1:0] node13043;
	wire [4-1:0] node13045;
	wire [4-1:0] node13048;
	wire [4-1:0] node13050;
	wire [4-1:0] node13053;
	wire [4-1:0] node13054;
	wire [4-1:0] node13057;
	wire [4-1:0] node13060;
	wire [4-1:0] node13061;
	wire [4-1:0] node13062;
	wire [4-1:0] node13063;
	wire [4-1:0] node13066;
	wire [4-1:0] node13069;
	wire [4-1:0] node13070;
	wire [4-1:0] node13074;
	wire [4-1:0] node13075;
	wire [4-1:0] node13076;
	wire [4-1:0] node13079;
	wire [4-1:0] node13082;
	wire [4-1:0] node13083;
	wire [4-1:0] node13086;
	wire [4-1:0] node13089;
	wire [4-1:0] node13090;
	wire [4-1:0] node13091;
	wire [4-1:0] node13093;
	wire [4-1:0] node13095;
	wire [4-1:0] node13098;
	wire [4-1:0] node13099;
	wire [4-1:0] node13102;
	wire [4-1:0] node13103;
	wire [4-1:0] node13106;
	wire [4-1:0] node13109;
	wire [4-1:0] node13110;
	wire [4-1:0] node13111;
	wire [4-1:0] node13113;
	wire [4-1:0] node13116;
	wire [4-1:0] node13117;
	wire [4-1:0] node13121;
	wire [4-1:0] node13122;
	wire [4-1:0] node13123;
	wire [4-1:0] node13127;
	wire [4-1:0] node13129;
	wire [4-1:0] node13132;
	wire [4-1:0] node13133;
	wire [4-1:0] node13134;
	wire [4-1:0] node13135;
	wire [4-1:0] node13136;
	wire [4-1:0] node13139;
	wire [4-1:0] node13141;
	wire [4-1:0] node13144;
	wire [4-1:0] node13145;
	wire [4-1:0] node13146;
	wire [4-1:0] node13150;
	wire [4-1:0] node13152;
	wire [4-1:0] node13155;
	wire [4-1:0] node13156;
	wire [4-1:0] node13157;
	wire [4-1:0] node13159;
	wire [4-1:0] node13162;
	wire [4-1:0] node13163;
	wire [4-1:0] node13167;
	wire [4-1:0] node13168;
	wire [4-1:0] node13169;
	wire [4-1:0] node13174;
	wire [4-1:0] node13175;
	wire [4-1:0] node13176;
	wire [4-1:0] node13177;
	wire [4-1:0] node13178;
	wire [4-1:0] node13182;
	wire [4-1:0] node13184;
	wire [4-1:0] node13187;
	wire [4-1:0] node13188;
	wire [4-1:0] node13191;
	wire [4-1:0] node13192;
	wire [4-1:0] node13196;
	wire [4-1:0] node13197;
	wire [4-1:0] node13198;
	wire [4-1:0] node13199;
	wire [4-1:0] node13202;
	wire [4-1:0] node13205;
	wire [4-1:0] node13206;
	wire [4-1:0] node13209;
	wire [4-1:0] node13212;
	wire [4-1:0] node13213;
	wire [4-1:0] node13214;
	wire [4-1:0] node13218;
	wire [4-1:0] node13220;
	wire [4-1:0] node13223;
	wire [4-1:0] node13224;
	wire [4-1:0] node13225;
	wire [4-1:0] node13226;
	wire [4-1:0] node13227;
	wire [4-1:0] node13228;
	wire [4-1:0] node13231;
	wire [4-1:0] node13234;
	wire [4-1:0] node13237;
	wire [4-1:0] node13238;
	wire [4-1:0] node13239;
	wire [4-1:0] node13240;
	wire [4-1:0] node13244;
	wire [4-1:0] node13246;
	wire [4-1:0] node13249;
	wire [4-1:0] node13250;
	wire [4-1:0] node13252;
	wire [4-1:0] node13255;
	wire [4-1:0] node13256;
	wire [4-1:0] node13260;
	wire [4-1:0] node13261;
	wire [4-1:0] node13262;
	wire [4-1:0] node13263;
	wire [4-1:0] node13266;
	wire [4-1:0] node13268;
	wire [4-1:0] node13271;
	wire [4-1:0] node13272;
	wire [4-1:0] node13275;
	wire [4-1:0] node13277;
	wire [4-1:0] node13280;
	wire [4-1:0] node13281;
	wire [4-1:0] node13282;
	wire [4-1:0] node13283;
	wire [4-1:0] node13286;
	wire [4-1:0] node13289;
	wire [4-1:0] node13292;
	wire [4-1:0] node13293;
	wire [4-1:0] node13294;
	wire [4-1:0] node13298;
	wire [4-1:0] node13300;
	wire [4-1:0] node13303;
	wire [4-1:0] node13304;
	wire [4-1:0] node13305;
	wire [4-1:0] node13306;
	wire [4-1:0] node13307;
	wire [4-1:0] node13309;
	wire [4-1:0] node13312;
	wire [4-1:0] node13314;
	wire [4-1:0] node13317;
	wire [4-1:0] node13319;
	wire [4-1:0] node13322;
	wire [4-1:0] node13323;
	wire [4-1:0] node13324;
	wire [4-1:0] node13325;
	wire [4-1:0] node13328;
	wire [4-1:0] node13331;
	wire [4-1:0] node13332;
	wire [4-1:0] node13335;
	wire [4-1:0] node13338;
	wire [4-1:0] node13339;
	wire [4-1:0] node13340;
	wire [4-1:0] node13344;
	wire [4-1:0] node13345;
	wire [4-1:0] node13349;
	wire [4-1:0] node13350;
	wire [4-1:0] node13351;
	wire [4-1:0] node13353;
	wire [4-1:0] node13354;
	wire [4-1:0] node13357;
	wire [4-1:0] node13360;
	wire [4-1:0] node13362;
	wire [4-1:0] node13364;
	wire [4-1:0] node13367;
	wire [4-1:0] node13368;
	wire [4-1:0] node13369;
	wire [4-1:0] node13370;
	wire [4-1:0] node13374;
	wire [4-1:0] node13375;
	wire [4-1:0] node13378;
	wire [4-1:0] node13381;
	wire [4-1:0] node13383;
	wire [4-1:0] node13384;
	wire [4-1:0] node13387;
	wire [4-1:0] node13390;
	wire [4-1:0] node13391;
	wire [4-1:0] node13392;
	wire [4-1:0] node13393;
	wire [4-1:0] node13394;
	wire [4-1:0] node13395;
	wire [4-1:0] node13396;
	wire [4-1:0] node13398;
	wire [4-1:0] node13399;
	wire [4-1:0] node13403;
	wire [4-1:0] node13404;
	wire [4-1:0] node13407;
	wire [4-1:0] node13409;
	wire [4-1:0] node13412;
	wire [4-1:0] node13413;
	wire [4-1:0] node13414;
	wire [4-1:0] node13416;
	wire [4-1:0] node13419;
	wire [4-1:0] node13421;
	wire [4-1:0] node13424;
	wire [4-1:0] node13425;
	wire [4-1:0] node13427;
	wire [4-1:0] node13430;
	wire [4-1:0] node13431;
	wire [4-1:0] node13435;
	wire [4-1:0] node13436;
	wire [4-1:0] node13437;
	wire [4-1:0] node13438;
	wire [4-1:0] node13439;
	wire [4-1:0] node13443;
	wire [4-1:0] node13445;
	wire [4-1:0] node13448;
	wire [4-1:0] node13449;
	wire [4-1:0] node13450;
	wire [4-1:0] node13454;
	wire [4-1:0] node13456;
	wire [4-1:0] node13459;
	wire [4-1:0] node13460;
	wire [4-1:0] node13461;
	wire [4-1:0] node13462;
	wire [4-1:0] node13465;
	wire [4-1:0] node13468;
	wire [4-1:0] node13470;
	wire [4-1:0] node13473;
	wire [4-1:0] node13474;
	wire [4-1:0] node13475;
	wire [4-1:0] node13479;
	wire [4-1:0] node13481;
	wire [4-1:0] node13484;
	wire [4-1:0] node13485;
	wire [4-1:0] node13486;
	wire [4-1:0] node13487;
	wire [4-1:0] node13488;
	wire [4-1:0] node13492;
	wire [4-1:0] node13493;
	wire [4-1:0] node13494;
	wire [4-1:0] node13498;
	wire [4-1:0] node13499;
	wire [4-1:0] node13503;
	wire [4-1:0] node13504;
	wire [4-1:0] node13505;
	wire [4-1:0] node13506;
	wire [4-1:0] node13509;
	wire [4-1:0] node13512;
	wire [4-1:0] node13513;
	wire [4-1:0] node13517;
	wire [4-1:0] node13518;
	wire [4-1:0] node13521;
	wire [4-1:0] node13522;
	wire [4-1:0] node13526;
	wire [4-1:0] node13527;
	wire [4-1:0] node13528;
	wire [4-1:0] node13529;
	wire [4-1:0] node13530;
	wire [4-1:0] node13534;
	wire [4-1:0] node13535;
	wire [4-1:0] node13538;
	wire [4-1:0] node13541;
	wire [4-1:0] node13542;
	wire [4-1:0] node13543;
	wire [4-1:0] node13547;
	wire [4-1:0] node13548;
	wire [4-1:0] node13551;
	wire [4-1:0] node13554;
	wire [4-1:0] node13555;
	wire [4-1:0] node13557;
	wire [4-1:0] node13558;
	wire [4-1:0] node13561;
	wire [4-1:0] node13564;
	wire [4-1:0] node13565;
	wire [4-1:0] node13566;
	wire [4-1:0] node13570;
	wire [4-1:0] node13572;
	wire [4-1:0] node13575;
	wire [4-1:0] node13576;
	wire [4-1:0] node13577;
	wire [4-1:0] node13578;
	wire [4-1:0] node13579;
	wire [4-1:0] node13580;
	wire [4-1:0] node13581;
	wire [4-1:0] node13585;
	wire [4-1:0] node13586;
	wire [4-1:0] node13590;
	wire [4-1:0] node13591;
	wire [4-1:0] node13594;
	wire [4-1:0] node13595;
	wire [4-1:0] node13599;
	wire [4-1:0] node13600;
	wire [4-1:0] node13601;
	wire [4-1:0] node13602;
	wire [4-1:0] node13606;
	wire [4-1:0] node13607;
	wire [4-1:0] node13611;
	wire [4-1:0] node13612;
	wire [4-1:0] node13613;
	wire [4-1:0] node13617;
	wire [4-1:0] node13618;
	wire [4-1:0] node13622;
	wire [4-1:0] node13623;
	wire [4-1:0] node13624;
	wire [4-1:0] node13625;
	wire [4-1:0] node13627;
	wire [4-1:0] node13630;
	wire [4-1:0] node13631;
	wire [4-1:0] node13635;
	wire [4-1:0] node13636;
	wire [4-1:0] node13638;
	wire [4-1:0] node13641;
	wire [4-1:0] node13642;
	wire [4-1:0] node13645;
	wire [4-1:0] node13648;
	wire [4-1:0] node13649;
	wire [4-1:0] node13650;
	wire [4-1:0] node13652;
	wire [4-1:0] node13655;
	wire [4-1:0] node13656;
	wire [4-1:0] node13660;
	wire [4-1:0] node13661;
	wire [4-1:0] node13663;
	wire [4-1:0] node13666;
	wire [4-1:0] node13667;
	wire [4-1:0] node13671;
	wire [4-1:0] node13672;
	wire [4-1:0] node13673;
	wire [4-1:0] node13674;
	wire [4-1:0] node13675;
	wire [4-1:0] node13677;
	wire [4-1:0] node13680;
	wire [4-1:0] node13682;
	wire [4-1:0] node13685;
	wire [4-1:0] node13686;
	wire [4-1:0] node13688;
	wire [4-1:0] node13691;
	wire [4-1:0] node13692;
	wire [4-1:0] node13696;
	wire [4-1:0] node13697;
	wire [4-1:0] node13698;
	wire [4-1:0] node13701;
	wire [4-1:0] node13702;
	wire [4-1:0] node13706;
	wire [4-1:0] node13707;
	wire [4-1:0] node13708;
	wire [4-1:0] node13713;
	wire [4-1:0] node13714;
	wire [4-1:0] node13715;
	wire [4-1:0] node13716;
	wire [4-1:0] node13717;
	wire [4-1:0] node13721;
	wire [4-1:0] node13722;
	wire [4-1:0] node13726;
	wire [4-1:0] node13728;
	wire [4-1:0] node13731;
	wire [4-1:0] node13732;
	wire [4-1:0] node13733;
	wire [4-1:0] node13734;
	wire [4-1:0] node13737;
	wire [4-1:0] node13740;
	wire [4-1:0] node13741;
	wire [4-1:0] node13745;
	wire [4-1:0] node13746;
	wire [4-1:0] node13747;
	wire [4-1:0] node13751;
	wire [4-1:0] node13754;
	wire [4-1:0] node13755;
	wire [4-1:0] node13756;
	wire [4-1:0] node13757;
	wire [4-1:0] node13758;
	wire [4-1:0] node13759;
	wire [4-1:0] node13760;
	wire [4-1:0] node13762;
	wire [4-1:0] node13766;
	wire [4-1:0] node13768;
	wire [4-1:0] node13769;
	wire [4-1:0] node13773;
	wire [4-1:0] node13774;
	wire [4-1:0] node13775;
	wire [4-1:0] node13776;
	wire [4-1:0] node13780;
	wire [4-1:0] node13783;
	wire [4-1:0] node13785;
	wire [4-1:0] node13786;
	wire [4-1:0] node13789;
	wire [4-1:0] node13792;
	wire [4-1:0] node13793;
	wire [4-1:0] node13794;
	wire [4-1:0] node13795;
	wire [4-1:0] node13796;
	wire [4-1:0] node13800;
	wire [4-1:0] node13801;
	wire [4-1:0] node13804;
	wire [4-1:0] node13807;
	wire [4-1:0] node13810;
	wire [4-1:0] node13811;
	wire [4-1:0] node13812;
	wire [4-1:0] node13814;
	wire [4-1:0] node13817;
	wire [4-1:0] node13818;
	wire [4-1:0] node13821;
	wire [4-1:0] node13824;
	wire [4-1:0] node13825;
	wire [4-1:0] node13828;
	wire [4-1:0] node13831;
	wire [4-1:0] node13832;
	wire [4-1:0] node13833;
	wire [4-1:0] node13834;
	wire [4-1:0] node13835;
	wire [4-1:0] node13838;
	wire [4-1:0] node13839;
	wire [4-1:0] node13842;
	wire [4-1:0] node13845;
	wire [4-1:0] node13847;
	wire [4-1:0] node13848;
	wire [4-1:0] node13851;
	wire [4-1:0] node13854;
	wire [4-1:0] node13855;
	wire [4-1:0] node13856;
	wire [4-1:0] node13857;
	wire [4-1:0] node13861;
	wire [4-1:0] node13862;
	wire [4-1:0] node13866;
	wire [4-1:0] node13867;
	wire [4-1:0] node13870;
	wire [4-1:0] node13871;
	wire [4-1:0] node13875;
	wire [4-1:0] node13876;
	wire [4-1:0] node13877;
	wire [4-1:0] node13878;
	wire [4-1:0] node13879;
	wire [4-1:0] node13882;
	wire [4-1:0] node13885;
	wire [4-1:0] node13888;
	wire [4-1:0] node13889;
	wire [4-1:0] node13891;
	wire [4-1:0] node13894;
	wire [4-1:0] node13896;
	wire [4-1:0] node13899;
	wire [4-1:0] node13900;
	wire [4-1:0] node13901;
	wire [4-1:0] node13903;
	wire [4-1:0] node13906;
	wire [4-1:0] node13908;
	wire [4-1:0] node13911;
	wire [4-1:0] node13912;
	wire [4-1:0] node13913;
	wire [4-1:0] node13916;
	wire [4-1:0] node13919;
	wire [4-1:0] node13921;
	wire [4-1:0] node13924;
	wire [4-1:0] node13925;
	wire [4-1:0] node13926;
	wire [4-1:0] node13927;
	wire [4-1:0] node13928;
	wire [4-1:0] node13929;
	wire [4-1:0] node13930;
	wire [4-1:0] node13934;
	wire [4-1:0] node13936;
	wire [4-1:0] node13939;
	wire [4-1:0] node13940;
	wire [4-1:0] node13942;
	wire [4-1:0] node13945;
	wire [4-1:0] node13947;
	wire [4-1:0] node13950;
	wire [4-1:0] node13951;
	wire [4-1:0] node13952;
	wire [4-1:0] node13955;
	wire [4-1:0] node13956;
	wire [4-1:0] node13959;
	wire [4-1:0] node13962;
	wire [4-1:0] node13963;
	wire [4-1:0] node13967;
	wire [4-1:0] node13968;
	wire [4-1:0] node13969;
	wire [4-1:0] node13970;
	wire [4-1:0] node13971;
	wire [4-1:0] node13975;
	wire [4-1:0] node13976;
	wire [4-1:0] node13979;
	wire [4-1:0] node13982;
	wire [4-1:0] node13983;
	wire [4-1:0] node13984;
	wire [4-1:0] node13988;
	wire [4-1:0] node13989;
	wire [4-1:0] node13993;
	wire [4-1:0] node13994;
	wire [4-1:0] node13996;
	wire [4-1:0] node13997;
	wire [4-1:0] node14001;
	wire [4-1:0] node14002;
	wire [4-1:0] node14003;
	wire [4-1:0] node14006;
	wire [4-1:0] node14009;
	wire [4-1:0] node14010;
	wire [4-1:0] node14013;
	wire [4-1:0] node14016;
	wire [4-1:0] node14017;
	wire [4-1:0] node14018;
	wire [4-1:0] node14019;
	wire [4-1:0] node14021;
	wire [4-1:0] node14022;
	wire [4-1:0] node14026;
	wire [4-1:0] node14027;
	wire [4-1:0] node14031;
	wire [4-1:0] node14032;
	wire [4-1:0] node14033;
	wire [4-1:0] node14034;
	wire [4-1:0] node14037;
	wire [4-1:0] node14040;
	wire [4-1:0] node14042;
	wire [4-1:0] node14045;
	wire [4-1:0] node14046;
	wire [4-1:0] node14047;
	wire [4-1:0] node14051;
	wire [4-1:0] node14054;
	wire [4-1:0] node14055;
	wire [4-1:0] node14056;
	wire [4-1:0] node14058;
	wire [4-1:0] node14059;
	wire [4-1:0] node14063;
	wire [4-1:0] node14064;
	wire [4-1:0] node14065;
	wire [4-1:0] node14069;
	wire [4-1:0] node14071;
	wire [4-1:0] node14074;
	wire [4-1:0] node14075;
	wire [4-1:0] node14077;
	wire [4-1:0] node14079;
	wire [4-1:0] node14082;
	wire [4-1:0] node14083;
	wire [4-1:0] node14086;
	wire [4-1:0] node14087;
	wire [4-1:0] node14091;
	wire [4-1:0] node14092;
	wire [4-1:0] node14093;
	wire [4-1:0] node14094;
	wire [4-1:0] node14095;
	wire [4-1:0] node14096;
	wire [4-1:0] node14097;
	wire [4-1:0] node14098;
	wire [4-1:0] node14099;
	wire [4-1:0] node14100;
	wire [4-1:0] node14101;
	wire [4-1:0] node14104;
	wire [4-1:0] node14107;
	wire [4-1:0] node14109;
	wire [4-1:0] node14112;
	wire [4-1:0] node14113;
	wire [4-1:0] node14114;
	wire [4-1:0] node14118;
	wire [4-1:0] node14119;
	wire [4-1:0] node14122;
	wire [4-1:0] node14125;
	wire [4-1:0] node14126;
	wire [4-1:0] node14128;
	wire [4-1:0] node14130;
	wire [4-1:0] node14133;
	wire [4-1:0] node14134;
	wire [4-1:0] node14137;
	wire [4-1:0] node14140;
	wire [4-1:0] node14141;
	wire [4-1:0] node14142;
	wire [4-1:0] node14143;
	wire [4-1:0] node14144;
	wire [4-1:0] node14148;
	wire [4-1:0] node14149;
	wire [4-1:0] node14153;
	wire [4-1:0] node14154;
	wire [4-1:0] node14157;
	wire [4-1:0] node14160;
	wire [4-1:0] node14161;
	wire [4-1:0] node14162;
	wire [4-1:0] node14163;
	wire [4-1:0] node14167;
	wire [4-1:0] node14170;
	wire [4-1:0] node14171;
	wire [4-1:0] node14173;
	wire [4-1:0] node14176;
	wire [4-1:0] node14178;
	wire [4-1:0] node14181;
	wire [4-1:0] node14182;
	wire [4-1:0] node14183;
	wire [4-1:0] node14184;
	wire [4-1:0] node14186;
	wire [4-1:0] node14187;
	wire [4-1:0] node14190;
	wire [4-1:0] node14193;
	wire [4-1:0] node14194;
	wire [4-1:0] node14197;
	wire [4-1:0] node14199;
	wire [4-1:0] node14202;
	wire [4-1:0] node14203;
	wire [4-1:0] node14204;
	wire [4-1:0] node14205;
	wire [4-1:0] node14209;
	wire [4-1:0] node14210;
	wire [4-1:0] node14214;
	wire [4-1:0] node14215;
	wire [4-1:0] node14219;
	wire [4-1:0] node14220;
	wire [4-1:0] node14221;
	wire [4-1:0] node14222;
	wire [4-1:0] node14224;
	wire [4-1:0] node14227;
	wire [4-1:0] node14228;
	wire [4-1:0] node14232;
	wire [4-1:0] node14233;
	wire [4-1:0] node14234;
	wire [4-1:0] node14238;
	wire [4-1:0] node14241;
	wire [4-1:0] node14242;
	wire [4-1:0] node14244;
	wire [4-1:0] node14245;
	wire [4-1:0] node14249;
	wire [4-1:0] node14250;
	wire [4-1:0] node14253;
	wire [4-1:0] node14256;
	wire [4-1:0] node14257;
	wire [4-1:0] node14258;
	wire [4-1:0] node14259;
	wire [4-1:0] node14260;
	wire [4-1:0] node14262;
	wire [4-1:0] node14264;
	wire [4-1:0] node14267;
	wire [4-1:0] node14268;
	wire [4-1:0] node14271;
	wire [4-1:0] node14273;
	wire [4-1:0] node14276;
	wire [4-1:0] node14277;
	wire [4-1:0] node14278;
	wire [4-1:0] node14280;
	wire [4-1:0] node14283;
	wire [4-1:0] node14286;
	wire [4-1:0] node14287;
	wire [4-1:0] node14289;
	wire [4-1:0] node14292;
	wire [4-1:0] node14295;
	wire [4-1:0] node14296;
	wire [4-1:0] node14297;
	wire [4-1:0] node14298;
	wire [4-1:0] node14299;
	wire [4-1:0] node14303;
	wire [4-1:0] node14305;
	wire [4-1:0] node14308;
	wire [4-1:0] node14309;
	wire [4-1:0] node14311;
	wire [4-1:0] node14314;
	wire [4-1:0] node14316;
	wire [4-1:0] node14319;
	wire [4-1:0] node14320;
	wire [4-1:0] node14322;
	wire [4-1:0] node14325;
	wire [4-1:0] node14326;
	wire [4-1:0] node14328;
	wire [4-1:0] node14331;
	wire [4-1:0] node14334;
	wire [4-1:0] node14335;
	wire [4-1:0] node14336;
	wire [4-1:0] node14337;
	wire [4-1:0] node14338;
	wire [4-1:0] node14339;
	wire [4-1:0] node14344;
	wire [4-1:0] node14345;
	wire [4-1:0] node14346;
	wire [4-1:0] node14349;
	wire [4-1:0] node14352;
	wire [4-1:0] node14353;
	wire [4-1:0] node14356;
	wire [4-1:0] node14359;
	wire [4-1:0] node14360;
	wire [4-1:0] node14361;
	wire [4-1:0] node14364;
	wire [4-1:0] node14365;
	wire [4-1:0] node14369;
	wire [4-1:0] node14370;
	wire [4-1:0] node14372;
	wire [4-1:0] node14376;
	wire [4-1:0] node14377;
	wire [4-1:0] node14378;
	wire [4-1:0] node14379;
	wire [4-1:0] node14380;
	wire [4-1:0] node14383;
	wire [4-1:0] node14386;
	wire [4-1:0] node14388;
	wire [4-1:0] node14391;
	wire [4-1:0] node14392;
	wire [4-1:0] node14393;
	wire [4-1:0] node14396;
	wire [4-1:0] node14399;
	wire [4-1:0] node14400;
	wire [4-1:0] node14404;
	wire [4-1:0] node14405;
	wire [4-1:0] node14406;
	wire [4-1:0] node14407;
	wire [4-1:0] node14410;
	wire [4-1:0] node14413;
	wire [4-1:0] node14415;
	wire [4-1:0] node14418;
	wire [4-1:0] node14419;
	wire [4-1:0] node14420;
	wire [4-1:0] node14424;
	wire [4-1:0] node14427;
	wire [4-1:0] node14428;
	wire [4-1:0] node14429;
	wire [4-1:0] node14430;
	wire [4-1:0] node14431;
	wire [4-1:0] node14432;
	wire [4-1:0] node14433;
	wire [4-1:0] node14435;
	wire [4-1:0] node14438;
	wire [4-1:0] node14439;
	wire [4-1:0] node14443;
	wire [4-1:0] node14444;
	wire [4-1:0] node14445;
	wire [4-1:0] node14448;
	wire [4-1:0] node14451;
	wire [4-1:0] node14453;
	wire [4-1:0] node14456;
	wire [4-1:0] node14457;
	wire [4-1:0] node14458;
	wire [4-1:0] node14462;
	wire [4-1:0] node14463;
	wire [4-1:0] node14465;
	wire [4-1:0] node14468;
	wire [4-1:0] node14471;
	wire [4-1:0] node14472;
	wire [4-1:0] node14473;
	wire [4-1:0] node14474;
	wire [4-1:0] node14475;
	wire [4-1:0] node14479;
	wire [4-1:0] node14480;
	wire [4-1:0] node14483;
	wire [4-1:0] node14486;
	wire [4-1:0] node14487;
	wire [4-1:0] node14488;
	wire [4-1:0] node14491;
	wire [4-1:0] node14494;
	wire [4-1:0] node14495;
	wire [4-1:0] node14499;
	wire [4-1:0] node14500;
	wire [4-1:0] node14501;
	wire [4-1:0] node14503;
	wire [4-1:0] node14506;
	wire [4-1:0] node14509;
	wire [4-1:0] node14510;
	wire [4-1:0] node14511;
	wire [4-1:0] node14515;
	wire [4-1:0] node14516;
	wire [4-1:0] node14520;
	wire [4-1:0] node14521;
	wire [4-1:0] node14522;
	wire [4-1:0] node14523;
	wire [4-1:0] node14524;
	wire [4-1:0] node14525;
	wire [4-1:0] node14529;
	wire [4-1:0] node14530;
	wire [4-1:0] node14533;
	wire [4-1:0] node14536;
	wire [4-1:0] node14537;
	wire [4-1:0] node14538;
	wire [4-1:0] node14542;
	wire [4-1:0] node14544;
	wire [4-1:0] node14547;
	wire [4-1:0] node14548;
	wire [4-1:0] node14549;
	wire [4-1:0] node14552;
	wire [4-1:0] node14553;
	wire [4-1:0] node14557;
	wire [4-1:0] node14558;
	wire [4-1:0] node14559;
	wire [4-1:0] node14564;
	wire [4-1:0] node14565;
	wire [4-1:0] node14566;
	wire [4-1:0] node14567;
	wire [4-1:0] node14569;
	wire [4-1:0] node14572;
	wire [4-1:0] node14573;
	wire [4-1:0] node14577;
	wire [4-1:0] node14579;
	wire [4-1:0] node14580;
	wire [4-1:0] node14584;
	wire [4-1:0] node14585;
	wire [4-1:0] node14586;
	wire [4-1:0] node14588;
	wire [4-1:0] node14592;
	wire [4-1:0] node14593;
	wire [4-1:0] node14594;
	wire [4-1:0] node14598;
	wire [4-1:0] node14599;
	wire [4-1:0] node14602;
	wire [4-1:0] node14605;
	wire [4-1:0] node14606;
	wire [4-1:0] node14607;
	wire [4-1:0] node14608;
	wire [4-1:0] node14609;
	wire [4-1:0] node14610;
	wire [4-1:0] node14611;
	wire [4-1:0] node14614;
	wire [4-1:0] node14617;
	wire [4-1:0] node14618;
	wire [4-1:0] node14622;
	wire [4-1:0] node14623;
	wire [4-1:0] node14624;
	wire [4-1:0] node14628;
	wire [4-1:0] node14629;
	wire [4-1:0] node14633;
	wire [4-1:0] node14634;
	wire [4-1:0] node14635;
	wire [4-1:0] node14637;
	wire [4-1:0] node14640;
	wire [4-1:0] node14641;
	wire [4-1:0] node14645;
	wire [4-1:0] node14646;
	wire [4-1:0] node14647;
	wire [4-1:0] node14651;
	wire [4-1:0] node14654;
	wire [4-1:0] node14655;
	wire [4-1:0] node14656;
	wire [4-1:0] node14657;
	wire [4-1:0] node14659;
	wire [4-1:0] node14663;
	wire [4-1:0] node14664;
	wire [4-1:0] node14666;
	wire [4-1:0] node14669;
	wire [4-1:0] node14672;
	wire [4-1:0] node14673;
	wire [4-1:0] node14674;
	wire [4-1:0] node14675;
	wire [4-1:0] node14678;
	wire [4-1:0] node14681;
	wire [4-1:0] node14682;
	wire [4-1:0] node14686;
	wire [4-1:0] node14687;
	wire [4-1:0] node14690;
	wire [4-1:0] node14691;
	wire [4-1:0] node14695;
	wire [4-1:0] node14696;
	wire [4-1:0] node14697;
	wire [4-1:0] node14698;
	wire [4-1:0] node14699;
	wire [4-1:0] node14700;
	wire [4-1:0] node14704;
	wire [4-1:0] node14705;
	wire [4-1:0] node14708;
	wire [4-1:0] node14711;
	wire [4-1:0] node14712;
	wire [4-1:0] node14714;
	wire [4-1:0] node14717;
	wire [4-1:0] node14718;
	wire [4-1:0] node14721;
	wire [4-1:0] node14724;
	wire [4-1:0] node14725;
	wire [4-1:0] node14726;
	wire [4-1:0] node14728;
	wire [4-1:0] node14731;
	wire [4-1:0] node14733;
	wire [4-1:0] node14736;
	wire [4-1:0] node14737;
	wire [4-1:0] node14738;
	wire [4-1:0] node14742;
	wire [4-1:0] node14743;
	wire [4-1:0] node14746;
	wire [4-1:0] node14749;
	wire [4-1:0] node14750;
	wire [4-1:0] node14751;
	wire [4-1:0] node14753;
	wire [4-1:0] node14754;
	wire [4-1:0] node14758;
	wire [4-1:0] node14759;
	wire [4-1:0] node14760;
	wire [4-1:0] node14763;
	wire [4-1:0] node14766;
	wire [4-1:0] node14768;
	wire [4-1:0] node14771;
	wire [4-1:0] node14772;
	wire [4-1:0] node14773;
	wire [4-1:0] node14774;
	wire [4-1:0] node14777;
	wire [4-1:0] node14780;
	wire [4-1:0] node14782;
	wire [4-1:0] node14785;
	wire [4-1:0] node14786;
	wire [4-1:0] node14788;
	wire [4-1:0] node14792;
	wire [4-1:0] node14793;
	wire [4-1:0] node14794;
	wire [4-1:0] node14795;
	wire [4-1:0] node14796;
	wire [4-1:0] node14797;
	wire [4-1:0] node14798;
	wire [4-1:0] node14799;
	wire [4-1:0] node14801;
	wire [4-1:0] node14804;
	wire [4-1:0] node14807;
	wire [4-1:0] node14808;
	wire [4-1:0] node14809;
	wire [4-1:0] node14812;
	wire [4-1:0] node14815;
	wire [4-1:0] node14817;
	wire [4-1:0] node14820;
	wire [4-1:0] node14821;
	wire [4-1:0] node14823;
	wire [4-1:0] node14824;
	wire [4-1:0] node14828;
	wire [4-1:0] node14829;
	wire [4-1:0] node14831;
	wire [4-1:0] node14834;
	wire [4-1:0] node14835;
	wire [4-1:0] node14838;
	wire [4-1:0] node14841;
	wire [4-1:0] node14842;
	wire [4-1:0] node14843;
	wire [4-1:0] node14844;
	wire [4-1:0] node14846;
	wire [4-1:0] node14850;
	wire [4-1:0] node14851;
	wire [4-1:0] node14853;
	wire [4-1:0] node14856;
	wire [4-1:0] node14858;
	wire [4-1:0] node14861;
	wire [4-1:0] node14862;
	wire [4-1:0] node14863;
	wire [4-1:0] node14864;
	wire [4-1:0] node14867;
	wire [4-1:0] node14870;
	wire [4-1:0] node14872;
	wire [4-1:0] node14875;
	wire [4-1:0] node14876;
	wire [4-1:0] node14877;
	wire [4-1:0] node14880;
	wire [4-1:0] node14883;
	wire [4-1:0] node14884;
	wire [4-1:0] node14887;
	wire [4-1:0] node14890;
	wire [4-1:0] node14891;
	wire [4-1:0] node14892;
	wire [4-1:0] node14893;
	wire [4-1:0] node14894;
	wire [4-1:0] node14895;
	wire [4-1:0] node14898;
	wire [4-1:0] node14901;
	wire [4-1:0] node14903;
	wire [4-1:0] node14906;
	wire [4-1:0] node14907;
	wire [4-1:0] node14910;
	wire [4-1:0] node14913;
	wire [4-1:0] node14914;
	wire [4-1:0] node14915;
	wire [4-1:0] node14916;
	wire [4-1:0] node14919;
	wire [4-1:0] node14922;
	wire [4-1:0] node14923;
	wire [4-1:0] node14927;
	wire [4-1:0] node14928;
	wire [4-1:0] node14931;
	wire [4-1:0] node14933;
	wire [4-1:0] node14936;
	wire [4-1:0] node14937;
	wire [4-1:0] node14938;
	wire [4-1:0] node14939;
	wire [4-1:0] node14940;
	wire [4-1:0] node14943;
	wire [4-1:0] node14946;
	wire [4-1:0] node14947;
	wire [4-1:0] node14950;
	wire [4-1:0] node14953;
	wire [4-1:0] node14954;
	wire [4-1:0] node14955;
	wire [4-1:0] node14958;
	wire [4-1:0] node14961;
	wire [4-1:0] node14962;
	wire [4-1:0] node14966;
	wire [4-1:0] node14967;
	wire [4-1:0] node14968;
	wire [4-1:0] node14969;
	wire [4-1:0] node14972;
	wire [4-1:0] node14975;
	wire [4-1:0] node14977;
	wire [4-1:0] node14980;
	wire [4-1:0] node14981;
	wire [4-1:0] node14982;
	wire [4-1:0] node14985;
	wire [4-1:0] node14988;
	wire [4-1:0] node14991;
	wire [4-1:0] node14992;
	wire [4-1:0] node14993;
	wire [4-1:0] node14994;
	wire [4-1:0] node14995;
	wire [4-1:0] node14996;
	wire [4-1:0] node14997;
	wire [4-1:0] node15001;
	wire [4-1:0] node15002;
	wire [4-1:0] node15005;
	wire [4-1:0] node15008;
	wire [4-1:0] node15009;
	wire [4-1:0] node15010;
	wire [4-1:0] node15013;
	wire [4-1:0] node15016;
	wire [4-1:0] node15018;
	wire [4-1:0] node15021;
	wire [4-1:0] node15022;
	wire [4-1:0] node15023;
	wire [4-1:0] node15024;
	wire [4-1:0] node15027;
	wire [4-1:0] node15030;
	wire [4-1:0] node15031;
	wire [4-1:0] node15034;
	wire [4-1:0] node15037;
	wire [4-1:0] node15038;
	wire [4-1:0] node15039;
	wire [4-1:0] node15043;
	wire [4-1:0] node15044;
	wire [4-1:0] node15048;
	wire [4-1:0] node15049;
	wire [4-1:0] node15050;
	wire [4-1:0] node15051;
	wire [4-1:0] node15054;
	wire [4-1:0] node15056;
	wire [4-1:0] node15059;
	wire [4-1:0] node15060;
	wire [4-1:0] node15062;
	wire [4-1:0] node15065;
	wire [4-1:0] node15066;
	wire [4-1:0] node15069;
	wire [4-1:0] node15072;
	wire [4-1:0] node15073;
	wire [4-1:0] node15074;
	wire [4-1:0] node15077;
	wire [4-1:0] node15079;
	wire [4-1:0] node15082;
	wire [4-1:0] node15084;
	wire [4-1:0] node15085;
	wire [4-1:0] node15089;
	wire [4-1:0] node15090;
	wire [4-1:0] node15091;
	wire [4-1:0] node15092;
	wire [4-1:0] node15093;
	wire [4-1:0] node15094;
	wire [4-1:0] node15097;
	wire [4-1:0] node15100;
	wire [4-1:0] node15101;
	wire [4-1:0] node15104;
	wire [4-1:0] node15107;
	wire [4-1:0] node15108;
	wire [4-1:0] node15109;
	wire [4-1:0] node15112;
	wire [4-1:0] node15115;
	wire [4-1:0] node15116;
	wire [4-1:0] node15119;
	wire [4-1:0] node15122;
	wire [4-1:0] node15123;
	wire [4-1:0] node15125;
	wire [4-1:0] node15126;
	wire [4-1:0] node15129;
	wire [4-1:0] node15132;
	wire [4-1:0] node15133;
	wire [4-1:0] node15134;
	wire [4-1:0] node15138;
	wire [4-1:0] node15139;
	wire [4-1:0] node15142;
	wire [4-1:0] node15145;
	wire [4-1:0] node15146;
	wire [4-1:0] node15147;
	wire [4-1:0] node15148;
	wire [4-1:0] node15149;
	wire [4-1:0] node15152;
	wire [4-1:0] node15155;
	wire [4-1:0] node15158;
	wire [4-1:0] node15159;
	wire [4-1:0] node15162;
	wire [4-1:0] node15164;
	wire [4-1:0] node15167;
	wire [4-1:0] node15168;
	wire [4-1:0] node15169;
	wire [4-1:0] node15170;
	wire [4-1:0] node15175;
	wire [4-1:0] node15176;
	wire [4-1:0] node15179;
	wire [4-1:0] node15180;
	wire [4-1:0] node15184;
	wire [4-1:0] node15185;
	wire [4-1:0] node15186;
	wire [4-1:0] node15187;
	wire [4-1:0] node15188;
	wire [4-1:0] node15189;
	wire [4-1:0] node15190;
	wire [4-1:0] node15191;
	wire [4-1:0] node15196;
	wire [4-1:0] node15197;
	wire [4-1:0] node15199;
	wire [4-1:0] node15202;
	wire [4-1:0] node15205;
	wire [4-1:0] node15206;
	wire [4-1:0] node15207;
	wire [4-1:0] node15208;
	wire [4-1:0] node15212;
	wire [4-1:0] node15214;
	wire [4-1:0] node15217;
	wire [4-1:0] node15218;
	wire [4-1:0] node15219;
	wire [4-1:0] node15222;
	wire [4-1:0] node15226;
	wire [4-1:0] node15227;
	wire [4-1:0] node15228;
	wire [4-1:0] node15229;
	wire [4-1:0] node15232;
	wire [4-1:0] node15234;
	wire [4-1:0] node15237;
	wire [4-1:0] node15238;
	wire [4-1:0] node15239;
	wire [4-1:0] node15244;
	wire [4-1:0] node15245;
	wire [4-1:0] node15246;
	wire [4-1:0] node15247;
	wire [4-1:0] node15251;
	wire [4-1:0] node15252;
	wire [4-1:0] node15255;
	wire [4-1:0] node15258;
	wire [4-1:0] node15259;
	wire [4-1:0] node15260;
	wire [4-1:0] node15263;
	wire [4-1:0] node15266;
	wire [4-1:0] node15267;
	wire [4-1:0] node15271;
	wire [4-1:0] node15272;
	wire [4-1:0] node15273;
	wire [4-1:0] node15274;
	wire [4-1:0] node15275;
	wire [4-1:0] node15276;
	wire [4-1:0] node15280;
	wire [4-1:0] node15282;
	wire [4-1:0] node15285;
	wire [4-1:0] node15286;
	wire [4-1:0] node15288;
	wire [4-1:0] node15291;
	wire [4-1:0] node15293;
	wire [4-1:0] node15296;
	wire [4-1:0] node15297;
	wire [4-1:0] node15298;
	wire [4-1:0] node15299;
	wire [4-1:0] node15303;
	wire [4-1:0] node15305;
	wire [4-1:0] node15308;
	wire [4-1:0] node15309;
	wire [4-1:0] node15310;
	wire [4-1:0] node15313;
	wire [4-1:0] node15316;
	wire [4-1:0] node15319;
	wire [4-1:0] node15320;
	wire [4-1:0] node15321;
	wire [4-1:0] node15322;
	wire [4-1:0] node15325;
	wire [4-1:0] node15326;
	wire [4-1:0] node15330;
	wire [4-1:0] node15331;
	wire [4-1:0] node15332;
	wire [4-1:0] node15336;
	wire [4-1:0] node15337;
	wire [4-1:0] node15341;
	wire [4-1:0] node15342;
	wire [4-1:0] node15343;
	wire [4-1:0] node15347;
	wire [4-1:0] node15348;
	wire [4-1:0] node15351;
	wire [4-1:0] node15352;
	wire [4-1:0] node15356;
	wire [4-1:0] node15357;
	wire [4-1:0] node15358;
	wire [4-1:0] node15359;
	wire [4-1:0] node15360;
	wire [4-1:0] node15361;
	wire [4-1:0] node15363;
	wire [4-1:0] node15366;
	wire [4-1:0] node15367;
	wire [4-1:0] node15371;
	wire [4-1:0] node15372;
	wire [4-1:0] node15373;
	wire [4-1:0] node15377;
	wire [4-1:0] node15379;
	wire [4-1:0] node15382;
	wire [4-1:0] node15383;
	wire [4-1:0] node15384;
	wire [4-1:0] node15385;
	wire [4-1:0] node15389;
	wire [4-1:0] node15391;
	wire [4-1:0] node15394;
	wire [4-1:0] node15395;
	wire [4-1:0] node15397;
	wire [4-1:0] node15400;
	wire [4-1:0] node15403;
	wire [4-1:0] node15404;
	wire [4-1:0] node15405;
	wire [4-1:0] node15406;
	wire [4-1:0] node15407;
	wire [4-1:0] node15411;
	wire [4-1:0] node15412;
	wire [4-1:0] node15415;
	wire [4-1:0] node15418;
	wire [4-1:0] node15419;
	wire [4-1:0] node15420;
	wire [4-1:0] node15424;
	wire [4-1:0] node15426;
	wire [4-1:0] node15429;
	wire [4-1:0] node15430;
	wire [4-1:0] node15432;
	wire [4-1:0] node15433;
	wire [4-1:0] node15437;
	wire [4-1:0] node15440;
	wire [4-1:0] node15441;
	wire [4-1:0] node15442;
	wire [4-1:0] node15443;
	wire [4-1:0] node15444;
	wire [4-1:0] node15447;
	wire [4-1:0] node15450;
	wire [4-1:0] node15451;
	wire [4-1:0] node15452;
	wire [4-1:0] node15456;
	wire [4-1:0] node15459;
	wire [4-1:0] node15460;
	wire [4-1:0] node15461;
	wire [4-1:0] node15462;
	wire [4-1:0] node15467;
	wire [4-1:0] node15468;
	wire [4-1:0] node15471;
	wire [4-1:0] node15472;
	wire [4-1:0] node15476;
	wire [4-1:0] node15477;
	wire [4-1:0] node15478;
	wire [4-1:0] node15479;
	wire [4-1:0] node15482;
	wire [4-1:0] node15483;
	wire [4-1:0] node15487;
	wire [4-1:0] node15488;
	wire [4-1:0] node15489;
	wire [4-1:0] node15493;
	wire [4-1:0] node15494;
	wire [4-1:0] node15497;
	wire [4-1:0] node15500;
	wire [4-1:0] node15501;
	wire [4-1:0] node15503;
	wire [4-1:0] node15506;
	wire [4-1:0] node15507;
	wire [4-1:0] node15508;
	wire [4-1:0] node15512;
	wire [4-1:0] node15514;
	wire [4-1:0] node15517;
	wire [4-1:0] node15518;
	wire [4-1:0] node15519;
	wire [4-1:0] node15520;
	wire [4-1:0] node15521;
	wire [4-1:0] node15522;
	wire [4-1:0] node15523;
	wire [4-1:0] node15524;
	wire [4-1:0] node15525;
	wire [4-1:0] node15526;
	wire [4-1:0] node15530;
	wire [4-1:0] node15531;
	wire [4-1:0] node15535;
	wire [4-1:0] node15536;
	wire [4-1:0] node15540;
	wire [4-1:0] node15541;
	wire [4-1:0] node15543;
	wire [4-1:0] node15544;
	wire [4-1:0] node15548;
	wire [4-1:0] node15549;
	wire [4-1:0] node15551;
	wire [4-1:0] node15554;
	wire [4-1:0] node15555;
	wire [4-1:0] node15558;
	wire [4-1:0] node15561;
	wire [4-1:0] node15562;
	wire [4-1:0] node15563;
	wire [4-1:0] node15565;
	wire [4-1:0] node15568;
	wire [4-1:0] node15570;
	wire [4-1:0] node15573;
	wire [4-1:0] node15574;
	wire [4-1:0] node15575;
	wire [4-1:0] node15576;
	wire [4-1:0] node15579;
	wire [4-1:0] node15582;
	wire [4-1:0] node15585;
	wire [4-1:0] node15586;
	wire [4-1:0] node15588;
	wire [4-1:0] node15591;
	wire [4-1:0] node15592;
	wire [4-1:0] node15596;
	wire [4-1:0] node15597;
	wire [4-1:0] node15598;
	wire [4-1:0] node15599;
	wire [4-1:0] node15600;
	wire [4-1:0] node15603;
	wire [4-1:0] node15604;
	wire [4-1:0] node15607;
	wire [4-1:0] node15610;
	wire [4-1:0] node15611;
	wire [4-1:0] node15613;
	wire [4-1:0] node15616;
	wire [4-1:0] node15619;
	wire [4-1:0] node15620;
	wire [4-1:0] node15621;
	wire [4-1:0] node15624;
	wire [4-1:0] node15625;
	wire [4-1:0] node15629;
	wire [4-1:0] node15630;
	wire [4-1:0] node15631;
	wire [4-1:0] node15634;
	wire [4-1:0] node15637;
	wire [4-1:0] node15638;
	wire [4-1:0] node15641;
	wire [4-1:0] node15644;
	wire [4-1:0] node15645;
	wire [4-1:0] node15646;
	wire [4-1:0] node15647;
	wire [4-1:0] node15649;
	wire [4-1:0] node15652;
	wire [4-1:0] node15654;
	wire [4-1:0] node15657;
	wire [4-1:0] node15658;
	wire [4-1:0] node15660;
	wire [4-1:0] node15663;
	wire [4-1:0] node15664;
	wire [4-1:0] node15667;
	wire [4-1:0] node15670;
	wire [4-1:0] node15671;
	wire [4-1:0] node15672;
	wire [4-1:0] node15673;
	wire [4-1:0] node15677;
	wire [4-1:0] node15678;
	wire [4-1:0] node15681;
	wire [4-1:0] node15684;
	wire [4-1:0] node15685;
	wire [4-1:0] node15686;
	wire [4-1:0] node15690;
	wire [4-1:0] node15691;
	wire [4-1:0] node15694;
	wire [4-1:0] node15697;
	wire [4-1:0] node15698;
	wire [4-1:0] node15699;
	wire [4-1:0] node15700;
	wire [4-1:0] node15701;
	wire [4-1:0] node15702;
	wire [4-1:0] node15703;
	wire [4-1:0] node15707;
	wire [4-1:0] node15710;
	wire [4-1:0] node15712;
	wire [4-1:0] node15713;
	wire [4-1:0] node15716;
	wire [4-1:0] node15719;
	wire [4-1:0] node15720;
	wire [4-1:0] node15721;
	wire [4-1:0] node15722;
	wire [4-1:0] node15726;
	wire [4-1:0] node15728;
	wire [4-1:0] node15731;
	wire [4-1:0] node15732;
	wire [4-1:0] node15733;
	wire [4-1:0] node15737;
	wire [4-1:0] node15739;
	wire [4-1:0] node15742;
	wire [4-1:0] node15743;
	wire [4-1:0] node15744;
	wire [4-1:0] node15745;
	wire [4-1:0] node15747;
	wire [4-1:0] node15750;
	wire [4-1:0] node15752;
	wire [4-1:0] node15755;
	wire [4-1:0] node15757;
	wire [4-1:0] node15758;
	wire [4-1:0] node15761;
	wire [4-1:0] node15764;
	wire [4-1:0] node15765;
	wire [4-1:0] node15766;
	wire [4-1:0] node15769;
	wire [4-1:0] node15771;
	wire [4-1:0] node15774;
	wire [4-1:0] node15775;
	wire [4-1:0] node15777;
	wire [4-1:0] node15781;
	wire [4-1:0] node15782;
	wire [4-1:0] node15783;
	wire [4-1:0] node15784;
	wire [4-1:0] node15785;
	wire [4-1:0] node15786;
	wire [4-1:0] node15790;
	wire [4-1:0] node15791;
	wire [4-1:0] node15795;
	wire [4-1:0] node15796;
	wire [4-1:0] node15797;
	wire [4-1:0] node15800;
	wire [4-1:0] node15803;
	wire [4-1:0] node15804;
	wire [4-1:0] node15807;
	wire [4-1:0] node15810;
	wire [4-1:0] node15811;
	wire [4-1:0] node15812;
	wire [4-1:0] node15813;
	wire [4-1:0] node15817;
	wire [4-1:0] node15818;
	wire [4-1:0] node15821;
	wire [4-1:0] node15824;
	wire [4-1:0] node15825;
	wire [4-1:0] node15827;
	wire [4-1:0] node15830;
	wire [4-1:0] node15831;
	wire [4-1:0] node15835;
	wire [4-1:0] node15836;
	wire [4-1:0] node15837;
	wire [4-1:0] node15838;
	wire [4-1:0] node15839;
	wire [4-1:0] node15842;
	wire [4-1:0] node15845;
	wire [4-1:0] node15846;
	wire [4-1:0] node15849;
	wire [4-1:0] node15852;
	wire [4-1:0] node15853;
	wire [4-1:0] node15854;
	wire [4-1:0] node15857;
	wire [4-1:0] node15860;
	wire [4-1:0] node15862;
	wire [4-1:0] node15865;
	wire [4-1:0] node15866;
	wire [4-1:0] node15868;
	wire [4-1:0] node15870;
	wire [4-1:0] node15873;
	wire [4-1:0] node15874;
	wire [4-1:0] node15875;
	wire [4-1:0] node15879;
	wire [4-1:0] node15882;
	wire [4-1:0] node15883;
	wire [4-1:0] node15884;
	wire [4-1:0] node15885;
	wire [4-1:0] node15886;
	wire [4-1:0] node15887;
	wire [4-1:0] node15888;
	wire [4-1:0] node15889;
	wire [4-1:0] node15893;
	wire [4-1:0] node15895;
	wire [4-1:0] node15898;
	wire [4-1:0] node15899;
	wire [4-1:0] node15902;
	wire [4-1:0] node15903;
	wire [4-1:0] node15906;
	wire [4-1:0] node15909;
	wire [4-1:0] node15910;
	wire [4-1:0] node15911;
	wire [4-1:0] node15913;
	wire [4-1:0] node15916;
	wire [4-1:0] node15917;
	wire [4-1:0] node15921;
	wire [4-1:0] node15922;
	wire [4-1:0] node15923;
	wire [4-1:0] node15927;
	wire [4-1:0] node15930;
	wire [4-1:0] node15931;
	wire [4-1:0] node15932;
	wire [4-1:0] node15933;
	wire [4-1:0] node15934;
	wire [4-1:0] node15937;
	wire [4-1:0] node15940;
	wire [4-1:0] node15943;
	wire [4-1:0] node15944;
	wire [4-1:0] node15945;
	wire [4-1:0] node15949;
	wire [4-1:0] node15950;
	wire [4-1:0] node15953;
	wire [4-1:0] node15956;
	wire [4-1:0] node15957;
	wire [4-1:0] node15958;
	wire [4-1:0] node15959;
	wire [4-1:0] node15963;
	wire [4-1:0] node15964;
	wire [4-1:0] node15967;
	wire [4-1:0] node15970;
	wire [4-1:0] node15971;
	wire [4-1:0] node15973;
	wire [4-1:0] node15976;
	wire [4-1:0] node15977;
	wire [4-1:0] node15981;
	wire [4-1:0] node15982;
	wire [4-1:0] node15983;
	wire [4-1:0] node15984;
	wire [4-1:0] node15985;
	wire [4-1:0] node15988;
	wire [4-1:0] node15989;
	wire [4-1:0] node15993;
	wire [4-1:0] node15994;
	wire [4-1:0] node15995;
	wire [4-1:0] node15998;
	wire [4-1:0] node16001;
	wire [4-1:0] node16004;
	wire [4-1:0] node16005;
	wire [4-1:0] node16006;
	wire [4-1:0] node16007;
	wire [4-1:0] node16011;
	wire [4-1:0] node16012;
	wire [4-1:0] node16016;
	wire [4-1:0] node16017;
	wire [4-1:0] node16018;
	wire [4-1:0] node16022;
	wire [4-1:0] node16024;
	wire [4-1:0] node16027;
	wire [4-1:0] node16028;
	wire [4-1:0] node16029;
	wire [4-1:0] node16031;
	wire [4-1:0] node16033;
	wire [4-1:0] node16036;
	wire [4-1:0] node16037;
	wire [4-1:0] node16038;
	wire [4-1:0] node16042;
	wire [4-1:0] node16045;
	wire [4-1:0] node16046;
	wire [4-1:0] node16047;
	wire [4-1:0] node16048;
	wire [4-1:0] node16051;
	wire [4-1:0] node16054;
	wire [4-1:0] node16055;
	wire [4-1:0] node16059;
	wire [4-1:0] node16060;
	wire [4-1:0] node16061;
	wire [4-1:0] node16066;
	wire [4-1:0] node16067;
	wire [4-1:0] node16068;
	wire [4-1:0] node16069;
	wire [4-1:0] node16070;
	wire [4-1:0] node16071;
	wire [4-1:0] node16072;
	wire [4-1:0] node16075;
	wire [4-1:0] node16078;
	wire [4-1:0] node16080;
	wire [4-1:0] node16083;
	wire [4-1:0] node16084;
	wire [4-1:0] node16085;
	wire [4-1:0] node16089;
	wire [4-1:0] node16090;
	wire [4-1:0] node16093;
	wire [4-1:0] node16096;
	wire [4-1:0] node16097;
	wire [4-1:0] node16098;
	wire [4-1:0] node16100;
	wire [4-1:0] node16103;
	wire [4-1:0] node16105;
	wire [4-1:0] node16108;
	wire [4-1:0] node16109;
	wire [4-1:0] node16110;
	wire [4-1:0] node16113;
	wire [4-1:0] node16116;
	wire [4-1:0] node16117;
	wire [4-1:0] node16121;
	wire [4-1:0] node16122;
	wire [4-1:0] node16123;
	wire [4-1:0] node16124;
	wire [4-1:0] node16127;
	wire [4-1:0] node16130;
	wire [4-1:0] node16131;
	wire [4-1:0] node16132;
	wire [4-1:0] node16135;
	wire [4-1:0] node16138;
	wire [4-1:0] node16139;
	wire [4-1:0] node16142;
	wire [4-1:0] node16145;
	wire [4-1:0] node16146;
	wire [4-1:0] node16147;
	wire [4-1:0] node16148;
	wire [4-1:0] node16152;
	wire [4-1:0] node16155;
	wire [4-1:0] node16156;
	wire [4-1:0] node16159;
	wire [4-1:0] node16160;
	wire [4-1:0] node16163;
	wire [4-1:0] node16166;
	wire [4-1:0] node16167;
	wire [4-1:0] node16168;
	wire [4-1:0] node16169;
	wire [4-1:0] node16170;
	wire [4-1:0] node16171;
	wire [4-1:0] node16175;
	wire [4-1:0] node16177;
	wire [4-1:0] node16180;
	wire [4-1:0] node16181;
	wire [4-1:0] node16182;
	wire [4-1:0] node16185;
	wire [4-1:0] node16188;
	wire [4-1:0] node16191;
	wire [4-1:0] node16192;
	wire [4-1:0] node16193;
	wire [4-1:0] node16196;
	wire [4-1:0] node16197;
	wire [4-1:0] node16201;
	wire [4-1:0] node16202;
	wire [4-1:0] node16203;
	wire [4-1:0] node16207;
	wire [4-1:0] node16210;
	wire [4-1:0] node16211;
	wire [4-1:0] node16212;
	wire [4-1:0] node16213;
	wire [4-1:0] node16214;
	wire [4-1:0] node16218;
	wire [4-1:0] node16220;
	wire [4-1:0] node16223;
	wire [4-1:0] node16224;
	wire [4-1:0] node16226;
	wire [4-1:0] node16229;
	wire [4-1:0] node16232;
	wire [4-1:0] node16233;
	wire [4-1:0] node16234;
	wire [4-1:0] node16237;
	wire [4-1:0] node16238;
	wire [4-1:0] node16242;
	wire [4-1:0] node16243;
	wire [4-1:0] node16244;
	wire [4-1:0] node16248;
	wire [4-1:0] node16249;
	wire [4-1:0] node16253;
	wire [4-1:0] node16254;
	wire [4-1:0] node16255;
	wire [4-1:0] node16256;
	wire [4-1:0] node16257;
	wire [4-1:0] node16258;
	wire [4-1:0] node16259;
	wire [4-1:0] node16260;
	wire [4-1:0] node16261;
	wire [4-1:0] node16265;
	wire [4-1:0] node16268;
	wire [4-1:0] node16269;
	wire [4-1:0] node16272;
	wire [4-1:0] node16273;
	wire [4-1:0] node16276;
	wire [4-1:0] node16279;
	wire [4-1:0] node16280;
	wire [4-1:0] node16281;
	wire [4-1:0] node16282;
	wire [4-1:0] node16285;
	wire [4-1:0] node16288;
	wire [4-1:0] node16289;
	wire [4-1:0] node16292;
	wire [4-1:0] node16295;
	wire [4-1:0] node16296;
	wire [4-1:0] node16298;
	wire [4-1:0] node16302;
	wire [4-1:0] node16303;
	wire [4-1:0] node16304;
	wire [4-1:0] node16305;
	wire [4-1:0] node16306;
	wire [4-1:0] node16309;
	wire [4-1:0] node16312;
	wire [4-1:0] node16313;
	wire [4-1:0] node16316;
	wire [4-1:0] node16319;
	wire [4-1:0] node16320;
	wire [4-1:0] node16321;
	wire [4-1:0] node16325;
	wire [4-1:0] node16328;
	wire [4-1:0] node16329;
	wire [4-1:0] node16330;
	wire [4-1:0] node16331;
	wire [4-1:0] node16334;
	wire [4-1:0] node16337;
	wire [4-1:0] node16338;
	wire [4-1:0] node16341;
	wire [4-1:0] node16344;
	wire [4-1:0] node16345;
	wire [4-1:0] node16348;
	wire [4-1:0] node16350;
	wire [4-1:0] node16353;
	wire [4-1:0] node16354;
	wire [4-1:0] node16355;
	wire [4-1:0] node16356;
	wire [4-1:0] node16357;
	wire [4-1:0] node16358;
	wire [4-1:0] node16361;
	wire [4-1:0] node16365;
	wire [4-1:0] node16366;
	wire [4-1:0] node16368;
	wire [4-1:0] node16371;
	wire [4-1:0] node16372;
	wire [4-1:0] node16376;
	wire [4-1:0] node16377;
	wire [4-1:0] node16378;
	wire [4-1:0] node16380;
	wire [4-1:0] node16383;
	wire [4-1:0] node16384;
	wire [4-1:0] node16388;
	wire [4-1:0] node16390;
	wire [4-1:0] node16392;
	wire [4-1:0] node16395;
	wire [4-1:0] node16396;
	wire [4-1:0] node16397;
	wire [4-1:0] node16399;
	wire [4-1:0] node16401;
	wire [4-1:0] node16404;
	wire [4-1:0] node16405;
	wire [4-1:0] node16408;
	wire [4-1:0] node16409;
	wire [4-1:0] node16413;
	wire [4-1:0] node16414;
	wire [4-1:0] node16415;
	wire [4-1:0] node16416;
	wire [4-1:0] node16420;
	wire [4-1:0] node16421;
	wire [4-1:0] node16425;
	wire [4-1:0] node16427;
	wire [4-1:0] node16429;
	wire [4-1:0] node16432;
	wire [4-1:0] node16433;
	wire [4-1:0] node16434;
	wire [4-1:0] node16435;
	wire [4-1:0] node16436;
	wire [4-1:0] node16437;
	wire [4-1:0] node16438;
	wire [4-1:0] node16441;
	wire [4-1:0] node16444;
	wire [4-1:0] node16445;
	wire [4-1:0] node16449;
	wire [4-1:0] node16450;
	wire [4-1:0] node16452;
	wire [4-1:0] node16456;
	wire [4-1:0] node16457;
	wire [4-1:0] node16458;
	wire [4-1:0] node16460;
	wire [4-1:0] node16463;
	wire [4-1:0] node16466;
	wire [4-1:0] node16467;
	wire [4-1:0] node16469;
	wire [4-1:0] node16472;
	wire [4-1:0] node16473;
	wire [4-1:0] node16477;
	wire [4-1:0] node16478;
	wire [4-1:0] node16479;
	wire [4-1:0] node16480;
	wire [4-1:0] node16481;
	wire [4-1:0] node16485;
	wire [4-1:0] node16486;
	wire [4-1:0] node16490;
	wire [4-1:0] node16491;
	wire [4-1:0] node16492;
	wire [4-1:0] node16496;
	wire [4-1:0] node16497;
	wire [4-1:0] node16500;
	wire [4-1:0] node16503;
	wire [4-1:0] node16504;
	wire [4-1:0] node16505;
	wire [4-1:0] node16506;
	wire [4-1:0] node16510;
	wire [4-1:0] node16511;
	wire [4-1:0] node16514;
	wire [4-1:0] node16517;
	wire [4-1:0] node16518;
	wire [4-1:0] node16519;
	wire [4-1:0] node16523;
	wire [4-1:0] node16525;
	wire [4-1:0] node16528;
	wire [4-1:0] node16529;
	wire [4-1:0] node16530;
	wire [4-1:0] node16531;
	wire [4-1:0] node16532;
	wire [4-1:0] node16534;
	wire [4-1:0] node16537;
	wire [4-1:0] node16538;
	wire [4-1:0] node16542;
	wire [4-1:0] node16543;
	wire [4-1:0] node16544;
	wire [4-1:0] node16547;
	wire [4-1:0] node16550;
	wire [4-1:0] node16551;
	wire [4-1:0] node16555;
	wire [4-1:0] node16556;
	wire [4-1:0] node16557;
	wire [4-1:0] node16558;
	wire [4-1:0] node16562;
	wire [4-1:0] node16564;
	wire [4-1:0] node16567;
	wire [4-1:0] node16568;
	wire [4-1:0] node16571;
	wire [4-1:0] node16573;
	wire [4-1:0] node16576;
	wire [4-1:0] node16577;
	wire [4-1:0] node16578;
	wire [4-1:0] node16579;
	wire [4-1:0] node16581;
	wire [4-1:0] node16584;
	wire [4-1:0] node16585;
	wire [4-1:0] node16588;
	wire [4-1:0] node16591;
	wire [4-1:0] node16592;
	wire [4-1:0] node16594;
	wire [4-1:0] node16598;
	wire [4-1:0] node16599;
	wire [4-1:0] node16600;
	wire [4-1:0] node16601;
	wire [4-1:0] node16605;
	wire [4-1:0] node16606;
	wire [4-1:0] node16610;
	wire [4-1:0] node16611;
	wire [4-1:0] node16612;
	wire [4-1:0] node16615;
	wire [4-1:0] node16618;
	wire [4-1:0] node16620;
	wire [4-1:0] node16623;
	wire [4-1:0] node16624;
	wire [4-1:0] node16625;
	wire [4-1:0] node16626;
	wire [4-1:0] node16627;
	wire [4-1:0] node16628;
	wire [4-1:0] node16629;
	wire [4-1:0] node16631;
	wire [4-1:0] node16634;
	wire [4-1:0] node16635;
	wire [4-1:0] node16639;
	wire [4-1:0] node16640;
	wire [4-1:0] node16641;
	wire [4-1:0] node16645;
	wire [4-1:0] node16646;
	wire [4-1:0] node16649;
	wire [4-1:0] node16652;
	wire [4-1:0] node16653;
	wire [4-1:0] node16654;
	wire [4-1:0] node16655;
	wire [4-1:0] node16658;
	wire [4-1:0] node16661;
	wire [4-1:0] node16662;
	wire [4-1:0] node16665;
	wire [4-1:0] node16668;
	wire [4-1:0] node16669;
	wire [4-1:0] node16670;
	wire [4-1:0] node16673;
	wire [4-1:0] node16676;
	wire [4-1:0] node16677;
	wire [4-1:0] node16681;
	wire [4-1:0] node16682;
	wire [4-1:0] node16683;
	wire [4-1:0] node16684;
	wire [4-1:0] node16686;
	wire [4-1:0] node16690;
	wire [4-1:0] node16691;
	wire [4-1:0] node16692;
	wire [4-1:0] node16695;
	wire [4-1:0] node16698;
	wire [4-1:0] node16699;
	wire [4-1:0] node16703;
	wire [4-1:0] node16704;
	wire [4-1:0] node16705;
	wire [4-1:0] node16707;
	wire [4-1:0] node16711;
	wire [4-1:0] node16712;
	wire [4-1:0] node16713;
	wire [4-1:0] node16716;
	wire [4-1:0] node16719;
	wire [4-1:0] node16720;
	wire [4-1:0] node16723;
	wire [4-1:0] node16726;
	wire [4-1:0] node16727;
	wire [4-1:0] node16728;
	wire [4-1:0] node16729;
	wire [4-1:0] node16730;
	wire [4-1:0] node16731;
	wire [4-1:0] node16734;
	wire [4-1:0] node16737;
	wire [4-1:0] node16739;
	wire [4-1:0] node16742;
	wire [4-1:0] node16743;
	wire [4-1:0] node16744;
	wire [4-1:0] node16748;
	wire [4-1:0] node16751;
	wire [4-1:0] node16752;
	wire [4-1:0] node16754;
	wire [4-1:0] node16757;
	wire [4-1:0] node16759;
	wire [4-1:0] node16760;
	wire [4-1:0] node16763;
	wire [4-1:0] node16766;
	wire [4-1:0] node16767;
	wire [4-1:0] node16768;
	wire [4-1:0] node16769;
	wire [4-1:0] node16770;
	wire [4-1:0] node16774;
	wire [4-1:0] node16777;
	wire [4-1:0] node16778;
	wire [4-1:0] node16780;
	wire [4-1:0] node16783;
	wire [4-1:0] node16784;
	wire [4-1:0] node16788;
	wire [4-1:0] node16789;
	wire [4-1:0] node16790;
	wire [4-1:0] node16791;
	wire [4-1:0] node16794;
	wire [4-1:0] node16797;
	wire [4-1:0] node16800;
	wire [4-1:0] node16801;
	wire [4-1:0] node16804;
	wire [4-1:0] node16807;
	wire [4-1:0] node16808;
	wire [4-1:0] node16809;
	wire [4-1:0] node16810;
	wire [4-1:0] node16811;
	wire [4-1:0] node16812;
	wire [4-1:0] node16813;
	wire [4-1:0] node16817;
	wire [4-1:0] node16818;
	wire [4-1:0] node16822;
	wire [4-1:0] node16823;
	wire [4-1:0] node16825;
	wire [4-1:0] node16828;
	wire [4-1:0] node16829;
	wire [4-1:0] node16833;
	wire [4-1:0] node16834;
	wire [4-1:0] node16835;
	wire [4-1:0] node16836;
	wire [4-1:0] node16840;
	wire [4-1:0] node16842;
	wire [4-1:0] node16845;
	wire [4-1:0] node16846;
	wire [4-1:0] node16849;
	wire [4-1:0] node16850;
	wire [4-1:0] node16854;
	wire [4-1:0] node16855;
	wire [4-1:0] node16856;
	wire [4-1:0] node16857;
	wire [4-1:0] node16860;
	wire [4-1:0] node16861;
	wire [4-1:0] node16864;
	wire [4-1:0] node16867;
	wire [4-1:0] node16868;
	wire [4-1:0] node16869;
	wire [4-1:0] node16873;
	wire [4-1:0] node16875;
	wire [4-1:0] node16878;
	wire [4-1:0] node16879;
	wire [4-1:0] node16880;
	wire [4-1:0] node16882;
	wire [4-1:0] node16885;
	wire [4-1:0] node16886;
	wire [4-1:0] node16890;
	wire [4-1:0] node16891;
	wire [4-1:0] node16893;
	wire [4-1:0] node16896;
	wire [4-1:0] node16897;
	wire [4-1:0] node16901;
	wire [4-1:0] node16902;
	wire [4-1:0] node16903;
	wire [4-1:0] node16904;
	wire [4-1:0] node16906;
	wire [4-1:0] node16909;
	wire [4-1:0] node16910;
	wire [4-1:0] node16911;
	wire [4-1:0] node16915;
	wire [4-1:0] node16916;
	wire [4-1:0] node16919;
	wire [4-1:0] node16922;
	wire [4-1:0] node16923;
	wire [4-1:0] node16924;
	wire [4-1:0] node16926;
	wire [4-1:0] node16929;
	wire [4-1:0] node16931;
	wire [4-1:0] node16934;
	wire [4-1:0] node16935;
	wire [4-1:0] node16937;
	wire [4-1:0] node16940;
	wire [4-1:0] node16942;
	wire [4-1:0] node16945;
	wire [4-1:0] node16946;
	wire [4-1:0] node16947;
	wire [4-1:0] node16948;
	wire [4-1:0] node16949;
	wire [4-1:0] node16952;
	wire [4-1:0] node16955;
	wire [4-1:0] node16956;
	wire [4-1:0] node16959;
	wire [4-1:0] node16962;
	wire [4-1:0] node16963;
	wire [4-1:0] node16964;
	wire [4-1:0] node16967;
	wire [4-1:0] node16970;
	wire [4-1:0] node16971;
	wire [4-1:0] node16975;
	wire [4-1:0] node16976;
	wire [4-1:0] node16977;
	wire [4-1:0] node16979;
	wire [4-1:0] node16982;
	wire [4-1:0] node16984;
	wire [4-1:0] node16987;
	wire [4-1:0] node16988;
	wire [4-1:0] node16989;
	wire [4-1:0] node16993;
	wire [4-1:0] node16994;
	wire [4-1:0] node16998;
	wire [4-1:0] node16999;
	wire [4-1:0] node17000;
	wire [4-1:0] node17001;
	wire [4-1:0] node17002;
	wire [4-1:0] node17003;
	wire [4-1:0] node17004;
	wire [4-1:0] node17005;
	wire [4-1:0] node17006;
	wire [4-1:0] node17007;
	wire [4-1:0] node17008;
	wire [4-1:0] node17009;
	wire [4-1:0] node17012;
	wire [4-1:0] node17016;
	wire [4-1:0] node17017;
	wire [4-1:0] node17020;
	wire [4-1:0] node17022;
	wire [4-1:0] node17025;
	wire [4-1:0] node17026;
	wire [4-1:0] node17027;
	wire [4-1:0] node17028;
	wire [4-1:0] node17031;
	wire [4-1:0] node17034;
	wire [4-1:0] node17036;
	wire [4-1:0] node17039;
	wire [4-1:0] node17040;
	wire [4-1:0] node17042;
	wire [4-1:0] node17045;
	wire [4-1:0] node17046;
	wire [4-1:0] node17050;
	wire [4-1:0] node17051;
	wire [4-1:0] node17052;
	wire [4-1:0] node17053;
	wire [4-1:0] node17054;
	wire [4-1:0] node17057;
	wire [4-1:0] node17060;
	wire [4-1:0] node17061;
	wire [4-1:0] node17064;
	wire [4-1:0] node17067;
	wire [4-1:0] node17068;
	wire [4-1:0] node17069;
	wire [4-1:0] node17073;
	wire [4-1:0] node17074;
	wire [4-1:0] node17078;
	wire [4-1:0] node17079;
	wire [4-1:0] node17080;
	wire [4-1:0] node17082;
	wire [4-1:0] node17085;
	wire [4-1:0] node17087;
	wire [4-1:0] node17090;
	wire [4-1:0] node17091;
	wire [4-1:0] node17092;
	wire [4-1:0] node17096;
	wire [4-1:0] node17097;
	wire [4-1:0] node17101;
	wire [4-1:0] node17102;
	wire [4-1:0] node17103;
	wire [4-1:0] node17104;
	wire [4-1:0] node17105;
	wire [4-1:0] node17106;
	wire [4-1:0] node17110;
	wire [4-1:0] node17111;
	wire [4-1:0] node17114;
	wire [4-1:0] node17117;
	wire [4-1:0] node17118;
	wire [4-1:0] node17121;
	wire [4-1:0] node17122;
	wire [4-1:0] node17125;
	wire [4-1:0] node17128;
	wire [4-1:0] node17129;
	wire [4-1:0] node17130;
	wire [4-1:0] node17131;
	wire [4-1:0] node17135;
	wire [4-1:0] node17136;
	wire [4-1:0] node17139;
	wire [4-1:0] node17142;
	wire [4-1:0] node17143;
	wire [4-1:0] node17146;
	wire [4-1:0] node17147;
	wire [4-1:0] node17151;
	wire [4-1:0] node17152;
	wire [4-1:0] node17153;
	wire [4-1:0] node17154;
	wire [4-1:0] node17155;
	wire [4-1:0] node17159;
	wire [4-1:0] node17161;
	wire [4-1:0] node17164;
	wire [4-1:0] node17166;
	wire [4-1:0] node17168;
	wire [4-1:0] node17171;
	wire [4-1:0] node17172;
	wire [4-1:0] node17173;
	wire [4-1:0] node17174;
	wire [4-1:0] node17178;
	wire [4-1:0] node17181;
	wire [4-1:0] node17182;
	wire [4-1:0] node17183;
	wire [4-1:0] node17186;
	wire [4-1:0] node17189;
	wire [4-1:0] node17192;
	wire [4-1:0] node17193;
	wire [4-1:0] node17194;
	wire [4-1:0] node17195;
	wire [4-1:0] node17196;
	wire [4-1:0] node17197;
	wire [4-1:0] node17199;
	wire [4-1:0] node17202;
	wire [4-1:0] node17204;
	wire [4-1:0] node17207;
	wire [4-1:0] node17208;
	wire [4-1:0] node17209;
	wire [4-1:0] node17212;
	wire [4-1:0] node17216;
	wire [4-1:0] node17217;
	wire [4-1:0] node17218;
	wire [4-1:0] node17219;
	wire [4-1:0] node17224;
	wire [4-1:0] node17225;
	wire [4-1:0] node17228;
	wire [4-1:0] node17229;
	wire [4-1:0] node17233;
	wire [4-1:0] node17234;
	wire [4-1:0] node17235;
	wire [4-1:0] node17236;
	wire [4-1:0] node17238;
	wire [4-1:0] node17241;
	wire [4-1:0] node17242;
	wire [4-1:0] node17246;
	wire [4-1:0] node17247;
	wire [4-1:0] node17249;
	wire [4-1:0] node17252;
	wire [4-1:0] node17253;
	wire [4-1:0] node17256;
	wire [4-1:0] node17259;
	wire [4-1:0] node17260;
	wire [4-1:0] node17261;
	wire [4-1:0] node17262;
	wire [4-1:0] node17266;
	wire [4-1:0] node17267;
	wire [4-1:0] node17270;
	wire [4-1:0] node17273;
	wire [4-1:0] node17274;
	wire [4-1:0] node17275;
	wire [4-1:0] node17279;
	wire [4-1:0] node17280;
	wire [4-1:0] node17283;
	wire [4-1:0] node17286;
	wire [4-1:0] node17287;
	wire [4-1:0] node17288;
	wire [4-1:0] node17289;
	wire [4-1:0] node17290;
	wire [4-1:0] node17291;
	wire [4-1:0] node17294;
	wire [4-1:0] node17297;
	wire [4-1:0] node17298;
	wire [4-1:0] node17301;
	wire [4-1:0] node17304;
	wire [4-1:0] node17305;
	wire [4-1:0] node17306;
	wire [4-1:0] node17309;
	wire [4-1:0] node17312;
	wire [4-1:0] node17313;
	wire [4-1:0] node17317;
	wire [4-1:0] node17318;
	wire [4-1:0] node17319;
	wire [4-1:0] node17321;
	wire [4-1:0] node17325;
	wire [4-1:0] node17326;
	wire [4-1:0] node17330;
	wire [4-1:0] node17331;
	wire [4-1:0] node17332;
	wire [4-1:0] node17333;
	wire [4-1:0] node17335;
	wire [4-1:0] node17338;
	wire [4-1:0] node17340;
	wire [4-1:0] node17343;
	wire [4-1:0] node17344;
	wire [4-1:0] node17345;
	wire [4-1:0] node17349;
	wire [4-1:0] node17351;
	wire [4-1:0] node17354;
	wire [4-1:0] node17355;
	wire [4-1:0] node17356;
	wire [4-1:0] node17358;
	wire [4-1:0] node17362;
	wire [4-1:0] node17363;
	wire [4-1:0] node17364;
	wire [4-1:0] node17368;
	wire [4-1:0] node17370;
	wire [4-1:0] node17373;
	wire [4-1:0] node17374;
	wire [4-1:0] node17375;
	wire [4-1:0] node17376;
	wire [4-1:0] node17377;
	wire [4-1:0] node17378;
	wire [4-1:0] node17379;
	wire [4-1:0] node17380;
	wire [4-1:0] node17383;
	wire [4-1:0] node17386;
	wire [4-1:0] node17389;
	wire [4-1:0] node17390;
	wire [4-1:0] node17391;
	wire [4-1:0] node17396;
	wire [4-1:0] node17397;
	wire [4-1:0] node17398;
	wire [4-1:0] node17400;
	wire [4-1:0] node17403;
	wire [4-1:0] node17404;
	wire [4-1:0] node17407;
	wire [4-1:0] node17410;
	wire [4-1:0] node17411;
	wire [4-1:0] node17412;
	wire [4-1:0] node17416;
	wire [4-1:0] node17417;
	wire [4-1:0] node17420;
	wire [4-1:0] node17423;
	wire [4-1:0] node17424;
	wire [4-1:0] node17425;
	wire [4-1:0] node17426;
	wire [4-1:0] node17427;
	wire [4-1:0] node17431;
	wire [4-1:0] node17433;
	wire [4-1:0] node17436;
	wire [4-1:0] node17437;
	wire [4-1:0] node17438;
	wire [4-1:0] node17441;
	wire [4-1:0] node17444;
	wire [4-1:0] node17445;
	wire [4-1:0] node17449;
	wire [4-1:0] node17450;
	wire [4-1:0] node17452;
	wire [4-1:0] node17455;
	wire [4-1:0] node17456;
	wire [4-1:0] node17457;
	wire [4-1:0] node17461;
	wire [4-1:0] node17463;
	wire [4-1:0] node17466;
	wire [4-1:0] node17467;
	wire [4-1:0] node17468;
	wire [4-1:0] node17469;
	wire [4-1:0] node17470;
	wire [4-1:0] node17471;
	wire [4-1:0] node17474;
	wire [4-1:0] node17477;
	wire [4-1:0] node17478;
	wire [4-1:0] node17482;
	wire [4-1:0] node17483;
	wire [4-1:0] node17484;
	wire [4-1:0] node17488;
	wire [4-1:0] node17489;
	wire [4-1:0] node17493;
	wire [4-1:0] node17494;
	wire [4-1:0] node17495;
	wire [4-1:0] node17497;
	wire [4-1:0] node17500;
	wire [4-1:0] node17501;
	wire [4-1:0] node17504;
	wire [4-1:0] node17507;
	wire [4-1:0] node17508;
	wire [4-1:0] node17509;
	wire [4-1:0] node17513;
	wire [4-1:0] node17514;
	wire [4-1:0] node17518;
	wire [4-1:0] node17519;
	wire [4-1:0] node17520;
	wire [4-1:0] node17521;
	wire [4-1:0] node17522;
	wire [4-1:0] node17525;
	wire [4-1:0] node17528;
	wire [4-1:0] node17529;
	wire [4-1:0] node17533;
	wire [4-1:0] node17534;
	wire [4-1:0] node17535;
	wire [4-1:0] node17539;
	wire [4-1:0] node17540;
	wire [4-1:0] node17544;
	wire [4-1:0] node17545;
	wire [4-1:0] node17546;
	wire [4-1:0] node17549;
	wire [4-1:0] node17551;
	wire [4-1:0] node17554;
	wire [4-1:0] node17555;
	wire [4-1:0] node17556;
	wire [4-1:0] node17559;
	wire [4-1:0] node17562;
	wire [4-1:0] node17564;
	wire [4-1:0] node17567;
	wire [4-1:0] node17568;
	wire [4-1:0] node17569;
	wire [4-1:0] node17570;
	wire [4-1:0] node17571;
	wire [4-1:0] node17573;
	wire [4-1:0] node17574;
	wire [4-1:0] node17577;
	wire [4-1:0] node17580;
	wire [4-1:0] node17581;
	wire [4-1:0] node17584;
	wire [4-1:0] node17585;
	wire [4-1:0] node17588;
	wire [4-1:0] node17591;
	wire [4-1:0] node17592;
	wire [4-1:0] node17594;
	wire [4-1:0] node17597;
	wire [4-1:0] node17598;
	wire [4-1:0] node17600;
	wire [4-1:0] node17603;
	wire [4-1:0] node17605;
	wire [4-1:0] node17608;
	wire [4-1:0] node17609;
	wire [4-1:0] node17610;
	wire [4-1:0] node17611;
	wire [4-1:0] node17612;
	wire [4-1:0] node17616;
	wire [4-1:0] node17617;
	wire [4-1:0] node17621;
	wire [4-1:0] node17622;
	wire [4-1:0] node17625;
	wire [4-1:0] node17626;
	wire [4-1:0] node17630;
	wire [4-1:0] node17631;
	wire [4-1:0] node17633;
	wire [4-1:0] node17634;
	wire [4-1:0] node17637;
	wire [4-1:0] node17640;
	wire [4-1:0] node17641;
	wire [4-1:0] node17644;
	wire [4-1:0] node17645;
	wire [4-1:0] node17649;
	wire [4-1:0] node17650;
	wire [4-1:0] node17651;
	wire [4-1:0] node17652;
	wire [4-1:0] node17653;
	wire [4-1:0] node17656;
	wire [4-1:0] node17657;
	wire [4-1:0] node17661;
	wire [4-1:0] node17662;
	wire [4-1:0] node17663;
	wire [4-1:0] node17666;
	wire [4-1:0] node17669;
	wire [4-1:0] node17671;
	wire [4-1:0] node17674;
	wire [4-1:0] node17675;
	wire [4-1:0] node17677;
	wire [4-1:0] node17679;
	wire [4-1:0] node17682;
	wire [4-1:0] node17683;
	wire [4-1:0] node17685;
	wire [4-1:0] node17688;
	wire [4-1:0] node17689;
	wire [4-1:0] node17693;
	wire [4-1:0] node17694;
	wire [4-1:0] node17695;
	wire [4-1:0] node17696;
	wire [4-1:0] node17698;
	wire [4-1:0] node17701;
	wire [4-1:0] node17702;
	wire [4-1:0] node17706;
	wire [4-1:0] node17707;
	wire [4-1:0] node17709;
	wire [4-1:0] node17712;
	wire [4-1:0] node17713;
	wire [4-1:0] node17716;
	wire [4-1:0] node17719;
	wire [4-1:0] node17720;
	wire [4-1:0] node17721;
	wire [4-1:0] node17722;
	wire [4-1:0] node17725;
	wire [4-1:0] node17728;
	wire [4-1:0] node17729;
	wire [4-1:0] node17733;
	wire [4-1:0] node17734;
	wire [4-1:0] node17735;
	wire [4-1:0] node17738;
	wire [4-1:0] node17742;
	wire [4-1:0] node17743;
	wire [4-1:0] node17744;
	wire [4-1:0] node17745;
	wire [4-1:0] node17746;
	wire [4-1:0] node17747;
	wire [4-1:0] node17748;
	wire [4-1:0] node17749;
	wire [4-1:0] node17750;
	wire [4-1:0] node17753;
	wire [4-1:0] node17756;
	wire [4-1:0] node17757;
	wire [4-1:0] node17761;
	wire [4-1:0] node17763;
	wire [4-1:0] node17764;
	wire [4-1:0] node17768;
	wire [4-1:0] node17769;
	wire [4-1:0] node17771;
	wire [4-1:0] node17772;
	wire [4-1:0] node17776;
	wire [4-1:0] node17778;
	wire [4-1:0] node17780;
	wire [4-1:0] node17783;
	wire [4-1:0] node17784;
	wire [4-1:0] node17785;
	wire [4-1:0] node17786;
	wire [4-1:0] node17788;
	wire [4-1:0] node17791;
	wire [4-1:0] node17793;
	wire [4-1:0] node17796;
	wire [4-1:0] node17797;
	wire [4-1:0] node17799;
	wire [4-1:0] node17802;
	wire [4-1:0] node17803;
	wire [4-1:0] node17806;
	wire [4-1:0] node17809;
	wire [4-1:0] node17810;
	wire [4-1:0] node17811;
	wire [4-1:0] node17813;
	wire [4-1:0] node17816;
	wire [4-1:0] node17818;
	wire [4-1:0] node17821;
	wire [4-1:0] node17822;
	wire [4-1:0] node17824;
	wire [4-1:0] node17828;
	wire [4-1:0] node17829;
	wire [4-1:0] node17830;
	wire [4-1:0] node17831;
	wire [4-1:0] node17832;
	wire [4-1:0] node17833;
	wire [4-1:0] node17837;
	wire [4-1:0] node17840;
	wire [4-1:0] node17842;
	wire [4-1:0] node17843;
	wire [4-1:0] node17846;
	wire [4-1:0] node17849;
	wire [4-1:0] node17850;
	wire [4-1:0] node17851;
	wire [4-1:0] node17853;
	wire [4-1:0] node17856;
	wire [4-1:0] node17857;
	wire [4-1:0] node17861;
	wire [4-1:0] node17862;
	wire [4-1:0] node17863;
	wire [4-1:0] node17866;
	wire [4-1:0] node17870;
	wire [4-1:0] node17871;
	wire [4-1:0] node17872;
	wire [4-1:0] node17873;
	wire [4-1:0] node17875;
	wire [4-1:0] node17878;
	wire [4-1:0] node17879;
	wire [4-1:0] node17883;
	wire [4-1:0] node17884;
	wire [4-1:0] node17886;
	wire [4-1:0] node17889;
	wire [4-1:0] node17890;
	wire [4-1:0] node17893;
	wire [4-1:0] node17896;
	wire [4-1:0] node17897;
	wire [4-1:0] node17898;
	wire [4-1:0] node17899;
	wire [4-1:0] node17903;
	wire [4-1:0] node17905;
	wire [4-1:0] node17908;
	wire [4-1:0] node17910;
	wire [4-1:0] node17912;
	wire [4-1:0] node17915;
	wire [4-1:0] node17916;
	wire [4-1:0] node17917;
	wire [4-1:0] node17918;
	wire [4-1:0] node17919;
	wire [4-1:0] node17920;
	wire [4-1:0] node17922;
	wire [4-1:0] node17925;
	wire [4-1:0] node17926;
	wire [4-1:0] node17930;
	wire [4-1:0] node17931;
	wire [4-1:0] node17934;
	wire [4-1:0] node17936;
	wire [4-1:0] node17939;
	wire [4-1:0] node17940;
	wire [4-1:0] node17941;
	wire [4-1:0] node17944;
	wire [4-1:0] node17945;
	wire [4-1:0] node17948;
	wire [4-1:0] node17951;
	wire [4-1:0] node17952;
	wire [4-1:0] node17953;
	wire [4-1:0] node17956;
	wire [4-1:0] node17959;
	wire [4-1:0] node17962;
	wire [4-1:0] node17963;
	wire [4-1:0] node17964;
	wire [4-1:0] node17965;
	wire [4-1:0] node17967;
	wire [4-1:0] node17970;
	wire [4-1:0] node17971;
	wire [4-1:0] node17974;
	wire [4-1:0] node17977;
	wire [4-1:0] node17978;
	wire [4-1:0] node17980;
	wire [4-1:0] node17984;
	wire [4-1:0] node17985;
	wire [4-1:0] node17986;
	wire [4-1:0] node17987;
	wire [4-1:0] node17990;
	wire [4-1:0] node17993;
	wire [4-1:0] node17995;
	wire [4-1:0] node17998;
	wire [4-1:0] node17999;
	wire [4-1:0] node18001;
	wire [4-1:0] node18004;
	wire [4-1:0] node18005;
	wire [4-1:0] node18008;
	wire [4-1:0] node18011;
	wire [4-1:0] node18012;
	wire [4-1:0] node18013;
	wire [4-1:0] node18014;
	wire [4-1:0] node18015;
	wire [4-1:0] node18018;
	wire [4-1:0] node18020;
	wire [4-1:0] node18023;
	wire [4-1:0] node18024;
	wire [4-1:0] node18025;
	wire [4-1:0] node18028;
	wire [4-1:0] node18031;
	wire [4-1:0] node18032;
	wire [4-1:0] node18036;
	wire [4-1:0] node18037;
	wire [4-1:0] node18038;
	wire [4-1:0] node18039;
	wire [4-1:0] node18043;
	wire [4-1:0] node18044;
	wire [4-1:0] node18047;
	wire [4-1:0] node18050;
	wire [4-1:0] node18053;
	wire [4-1:0] node18054;
	wire [4-1:0] node18055;
	wire [4-1:0] node18056;
	wire [4-1:0] node18058;
	wire [4-1:0] node18061;
	wire [4-1:0] node18064;
	wire [4-1:0] node18065;
	wire [4-1:0] node18066;
	wire [4-1:0] node18071;
	wire [4-1:0] node18072;
	wire [4-1:0] node18073;
	wire [4-1:0] node18074;
	wire [4-1:0] node18077;
	wire [4-1:0] node18080;
	wire [4-1:0] node18082;
	wire [4-1:0] node18085;
	wire [4-1:0] node18086;
	wire [4-1:0] node18089;
	wire [4-1:0] node18092;
	wire [4-1:0] node18093;
	wire [4-1:0] node18094;
	wire [4-1:0] node18095;
	wire [4-1:0] node18096;
	wire [4-1:0] node18097;
	wire [4-1:0] node18098;
	wire [4-1:0] node18099;
	wire [4-1:0] node18102;
	wire [4-1:0] node18105;
	wire [4-1:0] node18107;
	wire [4-1:0] node18110;
	wire [4-1:0] node18111;
	wire [4-1:0] node18112;
	wire [4-1:0] node18115;
	wire [4-1:0] node18118;
	wire [4-1:0] node18120;
	wire [4-1:0] node18123;
	wire [4-1:0] node18124;
	wire [4-1:0] node18125;
	wire [4-1:0] node18127;
	wire [4-1:0] node18131;
	wire [4-1:0] node18132;
	wire [4-1:0] node18134;
	wire [4-1:0] node18137;
	wire [4-1:0] node18139;
	wire [4-1:0] node18142;
	wire [4-1:0] node18143;
	wire [4-1:0] node18144;
	wire [4-1:0] node18145;
	wire [4-1:0] node18146;
	wire [4-1:0] node18150;
	wire [4-1:0] node18151;
	wire [4-1:0] node18154;
	wire [4-1:0] node18157;
	wire [4-1:0] node18158;
	wire [4-1:0] node18160;
	wire [4-1:0] node18163;
	wire [4-1:0] node18165;
	wire [4-1:0] node18168;
	wire [4-1:0] node18169;
	wire [4-1:0] node18170;
	wire [4-1:0] node18172;
	wire [4-1:0] node18176;
	wire [4-1:0] node18177;
	wire [4-1:0] node18178;
	wire [4-1:0] node18183;
	wire [4-1:0] node18184;
	wire [4-1:0] node18185;
	wire [4-1:0] node18186;
	wire [4-1:0] node18187;
	wire [4-1:0] node18189;
	wire [4-1:0] node18192;
	wire [4-1:0] node18194;
	wire [4-1:0] node18197;
	wire [4-1:0] node18198;
	wire [4-1:0] node18199;
	wire [4-1:0] node18202;
	wire [4-1:0] node18205;
	wire [4-1:0] node18206;
	wire [4-1:0] node18210;
	wire [4-1:0] node18211;
	wire [4-1:0] node18213;
	wire [4-1:0] node18215;
	wire [4-1:0] node18218;
	wire [4-1:0] node18219;
	wire [4-1:0] node18220;
	wire [4-1:0] node18224;
	wire [4-1:0] node18227;
	wire [4-1:0] node18228;
	wire [4-1:0] node18229;
	wire [4-1:0] node18230;
	wire [4-1:0] node18231;
	wire [4-1:0] node18236;
	wire [4-1:0] node18237;
	wire [4-1:0] node18239;
	wire [4-1:0] node18242;
	wire [4-1:0] node18243;
	wire [4-1:0] node18246;
	wire [4-1:0] node18249;
	wire [4-1:0] node18250;
	wire [4-1:0] node18251;
	wire [4-1:0] node18252;
	wire [4-1:0] node18256;
	wire [4-1:0] node18257;
	wire [4-1:0] node18261;
	wire [4-1:0] node18263;
	wire [4-1:0] node18264;
	wire [4-1:0] node18268;
	wire [4-1:0] node18269;
	wire [4-1:0] node18270;
	wire [4-1:0] node18271;
	wire [4-1:0] node18272;
	wire [4-1:0] node18273;
	wire [4-1:0] node18274;
	wire [4-1:0] node18278;
	wire [4-1:0] node18279;
	wire [4-1:0] node18283;
	wire [4-1:0] node18284;
	wire [4-1:0] node18286;
	wire [4-1:0] node18289;
	wire [4-1:0] node18290;
	wire [4-1:0] node18293;
	wire [4-1:0] node18296;
	wire [4-1:0] node18297;
	wire [4-1:0] node18298;
	wire [4-1:0] node18299;
	wire [4-1:0] node18304;
	wire [4-1:0] node18305;
	wire [4-1:0] node18306;
	wire [4-1:0] node18310;
	wire [4-1:0] node18311;
	wire [4-1:0] node18315;
	wire [4-1:0] node18316;
	wire [4-1:0] node18317;
	wire [4-1:0] node18318;
	wire [4-1:0] node18320;
	wire [4-1:0] node18323;
	wire [4-1:0] node18324;
	wire [4-1:0] node18328;
	wire [4-1:0] node18329;
	wire [4-1:0] node18332;
	wire [4-1:0] node18334;
	wire [4-1:0] node18337;
	wire [4-1:0] node18338;
	wire [4-1:0] node18340;
	wire [4-1:0] node18342;
	wire [4-1:0] node18345;
	wire [4-1:0] node18346;
	wire [4-1:0] node18347;
	wire [4-1:0] node18351;
	wire [4-1:0] node18352;
	wire [4-1:0] node18356;
	wire [4-1:0] node18357;
	wire [4-1:0] node18358;
	wire [4-1:0] node18359;
	wire [4-1:0] node18360;
	wire [4-1:0] node18361;
	wire [4-1:0] node18365;
	wire [4-1:0] node18367;
	wire [4-1:0] node18370;
	wire [4-1:0] node18371;
	wire [4-1:0] node18372;
	wire [4-1:0] node18375;
	wire [4-1:0] node18378;
	wire [4-1:0] node18380;
	wire [4-1:0] node18383;
	wire [4-1:0] node18384;
	wire [4-1:0] node18385;
	wire [4-1:0] node18387;
	wire [4-1:0] node18390;
	wire [4-1:0] node18391;
	wire [4-1:0] node18395;
	wire [4-1:0] node18396;
	wire [4-1:0] node18397;
	wire [4-1:0] node18401;
	wire [4-1:0] node18402;
	wire [4-1:0] node18406;
	wire [4-1:0] node18407;
	wire [4-1:0] node18408;
	wire [4-1:0] node18410;
	wire [4-1:0] node18413;
	wire [4-1:0] node18415;
	wire [4-1:0] node18416;
	wire [4-1:0] node18419;
	wire [4-1:0] node18422;
	wire [4-1:0] node18423;
	wire [4-1:0] node18424;
	wire [4-1:0] node18426;
	wire [4-1:0] node18429;
	wire [4-1:0] node18432;
	wire [4-1:0] node18433;
	wire [4-1:0] node18434;
	wire [4-1:0] node18438;
	wire [4-1:0] node18439;
	wire [4-1:0] node18443;
	wire [4-1:0] node18444;
	wire [4-1:0] node18445;
	wire [4-1:0] node18446;
	wire [4-1:0] node18447;
	wire [4-1:0] node18448;
	wire [4-1:0] node18449;
	wire [4-1:0] node18450;
	wire [4-1:0] node18452;
	wire [4-1:0] node18453;
	wire [4-1:0] node18456;
	wire [4-1:0] node18459;
	wire [4-1:0] node18460;
	wire [4-1:0] node18461;
	wire [4-1:0] node18465;
	wire [4-1:0] node18468;
	wire [4-1:0] node18469;
	wire [4-1:0] node18471;
	wire [4-1:0] node18473;
	wire [4-1:0] node18476;
	wire [4-1:0] node18477;
	wire [4-1:0] node18479;
	wire [4-1:0] node18482;
	wire [4-1:0] node18484;
	wire [4-1:0] node18487;
	wire [4-1:0] node18488;
	wire [4-1:0] node18489;
	wire [4-1:0] node18490;
	wire [4-1:0] node18491;
	wire [4-1:0] node18495;
	wire [4-1:0] node18497;
	wire [4-1:0] node18500;
	wire [4-1:0] node18501;
	wire [4-1:0] node18503;
	wire [4-1:0] node18506;
	wire [4-1:0] node18507;
	wire [4-1:0] node18511;
	wire [4-1:0] node18512;
	wire [4-1:0] node18514;
	wire [4-1:0] node18516;
	wire [4-1:0] node18519;
	wire [4-1:0] node18520;
	wire [4-1:0] node18521;
	wire [4-1:0] node18525;
	wire [4-1:0] node18528;
	wire [4-1:0] node18529;
	wire [4-1:0] node18530;
	wire [4-1:0] node18531;
	wire [4-1:0] node18532;
	wire [4-1:0] node18534;
	wire [4-1:0] node18537;
	wire [4-1:0] node18539;
	wire [4-1:0] node18542;
	wire [4-1:0] node18543;
	wire [4-1:0] node18544;
	wire [4-1:0] node18547;
	wire [4-1:0] node18550;
	wire [4-1:0] node18552;
	wire [4-1:0] node18555;
	wire [4-1:0] node18556;
	wire [4-1:0] node18557;
	wire [4-1:0] node18560;
	wire [4-1:0] node18563;
	wire [4-1:0] node18564;
	wire [4-1:0] node18565;
	wire [4-1:0] node18568;
	wire [4-1:0] node18571;
	wire [4-1:0] node18572;
	wire [4-1:0] node18575;
	wire [4-1:0] node18578;
	wire [4-1:0] node18579;
	wire [4-1:0] node18580;
	wire [4-1:0] node18581;
	wire [4-1:0] node18582;
	wire [4-1:0] node18586;
	wire [4-1:0] node18588;
	wire [4-1:0] node18591;
	wire [4-1:0] node18592;
	wire [4-1:0] node18593;
	wire [4-1:0] node18596;
	wire [4-1:0] node18599;
	wire [4-1:0] node18601;
	wire [4-1:0] node18604;
	wire [4-1:0] node18605;
	wire [4-1:0] node18606;
	wire [4-1:0] node18607;
	wire [4-1:0] node18610;
	wire [4-1:0] node18613;
	wire [4-1:0] node18614;
	wire [4-1:0] node18618;
	wire [4-1:0] node18619;
	wire [4-1:0] node18622;
	wire [4-1:0] node18623;
	wire [4-1:0] node18626;
	wire [4-1:0] node18629;
	wire [4-1:0] node18630;
	wire [4-1:0] node18631;
	wire [4-1:0] node18632;
	wire [4-1:0] node18633;
	wire [4-1:0] node18634;
	wire [4-1:0] node18635;
	wire [4-1:0] node18639;
	wire [4-1:0] node18642;
	wire [4-1:0] node18643;
	wire [4-1:0] node18644;
	wire [4-1:0] node18647;
	wire [4-1:0] node18650;
	wire [4-1:0] node18651;
	wire [4-1:0] node18655;
	wire [4-1:0] node18656;
	wire [4-1:0] node18657;
	wire [4-1:0] node18658;
	wire [4-1:0] node18661;
	wire [4-1:0] node18664;
	wire [4-1:0] node18665;
	wire [4-1:0] node18668;
	wire [4-1:0] node18671;
	wire [4-1:0] node18672;
	wire [4-1:0] node18673;
	wire [4-1:0] node18677;
	wire [4-1:0] node18679;
	wire [4-1:0] node18682;
	wire [4-1:0] node18683;
	wire [4-1:0] node18684;
	wire [4-1:0] node18686;
	wire [4-1:0] node18687;
	wire [4-1:0] node18691;
	wire [4-1:0] node18692;
	wire [4-1:0] node18693;
	wire [4-1:0] node18698;
	wire [4-1:0] node18699;
	wire [4-1:0] node18701;
	wire [4-1:0] node18702;
	wire [4-1:0] node18706;
	wire [4-1:0] node18708;
	wire [4-1:0] node18710;
	wire [4-1:0] node18713;
	wire [4-1:0] node18714;
	wire [4-1:0] node18715;
	wire [4-1:0] node18716;
	wire [4-1:0] node18717;
	wire [4-1:0] node18719;
	wire [4-1:0] node18723;
	wire [4-1:0] node18724;
	wire [4-1:0] node18725;
	wire [4-1:0] node18729;
	wire [4-1:0] node18732;
	wire [4-1:0] node18733;
	wire [4-1:0] node18734;
	wire [4-1:0] node18735;
	wire [4-1:0] node18740;
	wire [4-1:0] node18741;
	wire [4-1:0] node18742;
	wire [4-1:0] node18746;
	wire [4-1:0] node18749;
	wire [4-1:0] node18750;
	wire [4-1:0] node18751;
	wire [4-1:0] node18752;
	wire [4-1:0] node18753;
	wire [4-1:0] node18757;
	wire [4-1:0] node18759;
	wire [4-1:0] node18762;
	wire [4-1:0] node18763;
	wire [4-1:0] node18766;
	wire [4-1:0] node18769;
	wire [4-1:0] node18770;
	wire [4-1:0] node18771;
	wire [4-1:0] node18774;
	wire [4-1:0] node18775;
	wire [4-1:0] node18778;
	wire [4-1:0] node18781;
	wire [4-1:0] node18782;
	wire [4-1:0] node18784;
	wire [4-1:0] node18788;
	wire [4-1:0] node18789;
	wire [4-1:0] node18790;
	wire [4-1:0] node18791;
	wire [4-1:0] node18792;
	wire [4-1:0] node18793;
	wire [4-1:0] node18794;
	wire [4-1:0] node18795;
	wire [4-1:0] node18798;
	wire [4-1:0] node18801;
	wire [4-1:0] node18802;
	wire [4-1:0] node18805;
	wire [4-1:0] node18808;
	wire [4-1:0] node18809;
	wire [4-1:0] node18810;
	wire [4-1:0] node18814;
	wire [4-1:0] node18817;
	wire [4-1:0] node18818;
	wire [4-1:0] node18819;
	wire [4-1:0] node18820;
	wire [4-1:0] node18823;
	wire [4-1:0] node18826;
	wire [4-1:0] node18827;
	wire [4-1:0] node18830;
	wire [4-1:0] node18833;
	wire [4-1:0] node18834;
	wire [4-1:0] node18836;
	wire [4-1:0] node18839;
	wire [4-1:0] node18840;
	wire [4-1:0] node18843;
	wire [4-1:0] node18846;
	wire [4-1:0] node18847;
	wire [4-1:0] node18848;
	wire [4-1:0] node18849;
	wire [4-1:0] node18850;
	wire [4-1:0] node18853;
	wire [4-1:0] node18856;
	wire [4-1:0] node18858;
	wire [4-1:0] node18861;
	wire [4-1:0] node18862;
	wire [4-1:0] node18863;
	wire [4-1:0] node18866;
	wire [4-1:0] node18869;
	wire [4-1:0] node18870;
	wire [4-1:0] node18874;
	wire [4-1:0] node18875;
	wire [4-1:0] node18876;
	wire [4-1:0] node18877;
	wire [4-1:0] node18880;
	wire [4-1:0] node18883;
	wire [4-1:0] node18884;
	wire [4-1:0] node18888;
	wire [4-1:0] node18889;
	wire [4-1:0] node18890;
	wire [4-1:0] node18894;
	wire [4-1:0] node18896;
	wire [4-1:0] node18899;
	wire [4-1:0] node18900;
	wire [4-1:0] node18901;
	wire [4-1:0] node18902;
	wire [4-1:0] node18903;
	wire [4-1:0] node18905;
	wire [4-1:0] node18908;
	wire [4-1:0] node18909;
	wire [4-1:0] node18912;
	wire [4-1:0] node18915;
	wire [4-1:0] node18916;
	wire [4-1:0] node18917;
	wire [4-1:0] node18920;
	wire [4-1:0] node18923;
	wire [4-1:0] node18926;
	wire [4-1:0] node18927;
	wire [4-1:0] node18929;
	wire [4-1:0] node18930;
	wire [4-1:0] node18933;
	wire [4-1:0] node18936;
	wire [4-1:0] node18938;
	wire [4-1:0] node18939;
	wire [4-1:0] node18942;
	wire [4-1:0] node18945;
	wire [4-1:0] node18946;
	wire [4-1:0] node18947;
	wire [4-1:0] node18948;
	wire [4-1:0] node18951;
	wire [4-1:0] node18952;
	wire [4-1:0] node18956;
	wire [4-1:0] node18957;
	wire [4-1:0] node18959;
	wire [4-1:0] node18962;
	wire [4-1:0] node18963;
	wire [4-1:0] node18967;
	wire [4-1:0] node18968;
	wire [4-1:0] node18969;
	wire [4-1:0] node18970;
	wire [4-1:0] node18974;
	wire [4-1:0] node18976;
	wire [4-1:0] node18979;
	wire [4-1:0] node18980;
	wire [4-1:0] node18981;
	wire [4-1:0] node18984;
	wire [4-1:0] node18987;
	wire [4-1:0] node18988;
	wire [4-1:0] node18992;
	wire [4-1:0] node18993;
	wire [4-1:0] node18994;
	wire [4-1:0] node18995;
	wire [4-1:0] node18996;
	wire [4-1:0] node18997;
	wire [4-1:0] node18998;
	wire [4-1:0] node19001;
	wire [4-1:0] node19004;
	wire [4-1:0] node19005;
	wire [4-1:0] node19008;
	wire [4-1:0] node19011;
	wire [4-1:0] node19012;
	wire [4-1:0] node19014;
	wire [4-1:0] node19017;
	wire [4-1:0] node19018;
	wire [4-1:0] node19022;
	wire [4-1:0] node19023;
	wire [4-1:0] node19024;
	wire [4-1:0] node19026;
	wire [4-1:0] node19029;
	wire [4-1:0] node19030;
	wire [4-1:0] node19034;
	wire [4-1:0] node19035;
	wire [4-1:0] node19036;
	wire [4-1:0] node19039;
	wire [4-1:0] node19042;
	wire [4-1:0] node19044;
	wire [4-1:0] node19047;
	wire [4-1:0] node19048;
	wire [4-1:0] node19049;
	wire [4-1:0] node19050;
	wire [4-1:0] node19052;
	wire [4-1:0] node19055;
	wire [4-1:0] node19056;
	wire [4-1:0] node19060;
	wire [4-1:0] node19061;
	wire [4-1:0] node19064;
	wire [4-1:0] node19067;
	wire [4-1:0] node19068;
	wire [4-1:0] node19069;
	wire [4-1:0] node19071;
	wire [4-1:0] node19074;
	wire [4-1:0] node19077;
	wire [4-1:0] node19078;
	wire [4-1:0] node19079;
	wire [4-1:0] node19083;
	wire [4-1:0] node19084;
	wire [4-1:0] node19087;
	wire [4-1:0] node19090;
	wire [4-1:0] node19091;
	wire [4-1:0] node19092;
	wire [4-1:0] node19093;
	wire [4-1:0] node19094;
	wire [4-1:0] node19096;
	wire [4-1:0] node19099;
	wire [4-1:0] node19101;
	wire [4-1:0] node19104;
	wire [4-1:0] node19105;
	wire [4-1:0] node19106;
	wire [4-1:0] node19109;
	wire [4-1:0] node19112;
	wire [4-1:0] node19115;
	wire [4-1:0] node19116;
	wire [4-1:0] node19117;
	wire [4-1:0] node19118;
	wire [4-1:0] node19123;
	wire [4-1:0] node19124;
	wire [4-1:0] node19125;
	wire [4-1:0] node19129;
	wire [4-1:0] node19132;
	wire [4-1:0] node19133;
	wire [4-1:0] node19134;
	wire [4-1:0] node19136;
	wire [4-1:0] node19137;
	wire [4-1:0] node19141;
	wire [4-1:0] node19142;
	wire [4-1:0] node19144;
	wire [4-1:0] node19147;
	wire [4-1:0] node19148;
	wire [4-1:0] node19152;
	wire [4-1:0] node19153;
	wire [4-1:0] node19154;
	wire [4-1:0] node19155;
	wire [4-1:0] node19159;
	wire [4-1:0] node19162;
	wire [4-1:0] node19163;
	wire [4-1:0] node19164;
	wire [4-1:0] node19168;
	wire [4-1:0] node19169;
	wire [4-1:0] node19173;
	wire [4-1:0] node19174;
	wire [4-1:0] node19175;
	wire [4-1:0] node19176;
	wire [4-1:0] node19177;
	wire [4-1:0] node19178;
	wire [4-1:0] node19179;
	wire [4-1:0] node19180;
	wire [4-1:0] node19181;
	wire [4-1:0] node19184;
	wire [4-1:0] node19187;
	wire [4-1:0] node19190;
	wire [4-1:0] node19191;
	wire [4-1:0] node19194;
	wire [4-1:0] node19196;
	wire [4-1:0] node19199;
	wire [4-1:0] node19200;
	wire [4-1:0] node19201;
	wire [4-1:0] node19202;
	wire [4-1:0] node19205;
	wire [4-1:0] node19208;
	wire [4-1:0] node19209;
	wire [4-1:0] node19213;
	wire [4-1:0] node19214;
	wire [4-1:0] node19216;
	wire [4-1:0] node19219;
	wire [4-1:0] node19220;
	wire [4-1:0] node19224;
	wire [4-1:0] node19225;
	wire [4-1:0] node19226;
	wire [4-1:0] node19227;
	wire [4-1:0] node19228;
	wire [4-1:0] node19231;
	wire [4-1:0] node19234;
	wire [4-1:0] node19236;
	wire [4-1:0] node19239;
	wire [4-1:0] node19241;
	wire [4-1:0] node19242;
	wire [4-1:0] node19246;
	wire [4-1:0] node19247;
	wire [4-1:0] node19248;
	wire [4-1:0] node19250;
	wire [4-1:0] node19253;
	wire [4-1:0] node19255;
	wire [4-1:0] node19258;
	wire [4-1:0] node19259;
	wire [4-1:0] node19260;
	wire [4-1:0] node19263;
	wire [4-1:0] node19266;
	wire [4-1:0] node19268;
	wire [4-1:0] node19271;
	wire [4-1:0] node19272;
	wire [4-1:0] node19273;
	wire [4-1:0] node19274;
	wire [4-1:0] node19275;
	wire [4-1:0] node19277;
	wire [4-1:0] node19280;
	wire [4-1:0] node19282;
	wire [4-1:0] node19285;
	wire [4-1:0] node19286;
	wire [4-1:0] node19287;
	wire [4-1:0] node19291;
	wire [4-1:0] node19292;
	wire [4-1:0] node19295;
	wire [4-1:0] node19298;
	wire [4-1:0] node19299;
	wire [4-1:0] node19300;
	wire [4-1:0] node19302;
	wire [4-1:0] node19306;
	wire [4-1:0] node19307;
	wire [4-1:0] node19308;
	wire [4-1:0] node19312;
	wire [4-1:0] node19313;
	wire [4-1:0] node19317;
	wire [4-1:0] node19318;
	wire [4-1:0] node19319;
	wire [4-1:0] node19320;
	wire [4-1:0] node19323;
	wire [4-1:0] node19325;
	wire [4-1:0] node19328;
	wire [4-1:0] node19329;
	wire [4-1:0] node19330;
	wire [4-1:0] node19334;
	wire [4-1:0] node19335;
	wire [4-1:0] node19338;
	wire [4-1:0] node19341;
	wire [4-1:0] node19342;
	wire [4-1:0] node19343;
	wire [4-1:0] node19344;
	wire [4-1:0] node19348;
	wire [4-1:0] node19351;
	wire [4-1:0] node19352;
	wire [4-1:0] node19354;
	wire [4-1:0] node19357;
	wire [4-1:0] node19360;
	wire [4-1:0] node19361;
	wire [4-1:0] node19362;
	wire [4-1:0] node19363;
	wire [4-1:0] node19364;
	wire [4-1:0] node19366;
	wire [4-1:0] node19368;
	wire [4-1:0] node19371;
	wire [4-1:0] node19372;
	wire [4-1:0] node19374;
	wire [4-1:0] node19377;
	wire [4-1:0] node19378;
	wire [4-1:0] node19381;
	wire [4-1:0] node19384;
	wire [4-1:0] node19385;
	wire [4-1:0] node19386;
	wire [4-1:0] node19387;
	wire [4-1:0] node19391;
	wire [4-1:0] node19392;
	wire [4-1:0] node19396;
	wire [4-1:0] node19397;
	wire [4-1:0] node19398;
	wire [4-1:0] node19402;
	wire [4-1:0] node19405;
	wire [4-1:0] node19406;
	wire [4-1:0] node19407;
	wire [4-1:0] node19409;
	wire [4-1:0] node19412;
	wire [4-1:0] node19413;
	wire [4-1:0] node19414;
	wire [4-1:0] node19417;
	wire [4-1:0] node19420;
	wire [4-1:0] node19421;
	wire [4-1:0] node19425;
	wire [4-1:0] node19426;
	wire [4-1:0] node19427;
	wire [4-1:0] node19429;
	wire [4-1:0] node19432;
	wire [4-1:0] node19433;
	wire [4-1:0] node19437;
	wire [4-1:0] node19438;
	wire [4-1:0] node19440;
	wire [4-1:0] node19443;
	wire [4-1:0] node19444;
	wire [4-1:0] node19447;
	wire [4-1:0] node19450;
	wire [4-1:0] node19451;
	wire [4-1:0] node19452;
	wire [4-1:0] node19453;
	wire [4-1:0] node19454;
	wire [4-1:0] node19455;
	wire [4-1:0] node19458;
	wire [4-1:0] node19461;
	wire [4-1:0] node19462;
	wire [4-1:0] node19465;
	wire [4-1:0] node19468;
	wire [4-1:0] node19469;
	wire [4-1:0] node19470;
	wire [4-1:0] node19474;
	wire [4-1:0] node19475;
	wire [4-1:0] node19478;
	wire [4-1:0] node19481;
	wire [4-1:0] node19482;
	wire [4-1:0] node19483;
	wire [4-1:0] node19487;
	wire [4-1:0] node19488;
	wire [4-1:0] node19490;
	wire [4-1:0] node19493;
	wire [4-1:0] node19494;
	wire [4-1:0] node19498;
	wire [4-1:0] node19499;
	wire [4-1:0] node19500;
	wire [4-1:0] node19501;
	wire [4-1:0] node19502;
	wire [4-1:0] node19506;
	wire [4-1:0] node19507;
	wire [4-1:0] node19511;
	wire [4-1:0] node19513;
	wire [4-1:0] node19514;
	wire [4-1:0] node19517;
	wire [4-1:0] node19520;
	wire [4-1:0] node19521;
	wire [4-1:0] node19522;
	wire [4-1:0] node19524;
	wire [4-1:0] node19527;
	wire [4-1:0] node19530;
	wire [4-1:0] node19532;
	wire [4-1:0] node19533;
	wire [4-1:0] node19537;
	wire [4-1:0] node19538;
	wire [4-1:0] node19539;
	wire [4-1:0] node19540;
	wire [4-1:0] node19541;
	wire [4-1:0] node19542;
	wire [4-1:0] node19543;
	wire [4-1:0] node19546;
	wire [4-1:0] node19549;
	wire [4-1:0] node19551;
	wire [4-1:0] node19552;
	wire [4-1:0] node19555;
	wire [4-1:0] node19558;
	wire [4-1:0] node19559;
	wire [4-1:0] node19560;
	wire [4-1:0] node19561;
	wire [4-1:0] node19565;
	wire [4-1:0] node19566;
	wire [4-1:0] node19570;
	wire [4-1:0] node19571;
	wire [4-1:0] node19572;
	wire [4-1:0] node19576;
	wire [4-1:0] node19578;
	wire [4-1:0] node19581;
	wire [4-1:0] node19582;
	wire [4-1:0] node19583;
	wire [4-1:0] node19584;
	wire [4-1:0] node19585;
	wire [4-1:0] node19590;
	wire [4-1:0] node19591;
	wire [4-1:0] node19592;
	wire [4-1:0] node19596;
	wire [4-1:0] node19597;
	wire [4-1:0] node19601;
	wire [4-1:0] node19602;
	wire [4-1:0] node19603;
	wire [4-1:0] node19605;
	wire [4-1:0] node19608;
	wire [4-1:0] node19610;
	wire [4-1:0] node19613;
	wire [4-1:0] node19614;
	wire [4-1:0] node19615;
	wire [4-1:0] node19619;
	wire [4-1:0] node19621;
	wire [4-1:0] node19624;
	wire [4-1:0] node19625;
	wire [4-1:0] node19626;
	wire [4-1:0] node19627;
	wire [4-1:0] node19628;
	wire [4-1:0] node19631;
	wire [4-1:0] node19634;
	wire [4-1:0] node19635;
	wire [4-1:0] node19637;
	wire [4-1:0] node19640;
	wire [4-1:0] node19642;
	wire [4-1:0] node19645;
	wire [4-1:0] node19646;
	wire [4-1:0] node19647;
	wire [4-1:0] node19648;
	wire [4-1:0] node19651;
	wire [4-1:0] node19654;
	wire [4-1:0] node19655;
	wire [4-1:0] node19659;
	wire [4-1:0] node19660;
	wire [4-1:0] node19661;
	wire [4-1:0] node19664;
	wire [4-1:0] node19667;
	wire [4-1:0] node19669;
	wire [4-1:0] node19672;
	wire [4-1:0] node19673;
	wire [4-1:0] node19674;
	wire [4-1:0] node19675;
	wire [4-1:0] node19676;
	wire [4-1:0] node19680;
	wire [4-1:0] node19683;
	wire [4-1:0] node19684;
	wire [4-1:0] node19687;
	wire [4-1:0] node19689;
	wire [4-1:0] node19692;
	wire [4-1:0] node19693;
	wire [4-1:0] node19694;
	wire [4-1:0] node19695;
	wire [4-1:0] node19699;
	wire [4-1:0] node19702;
	wire [4-1:0] node19703;
	wire [4-1:0] node19705;
	wire [4-1:0] node19708;
	wire [4-1:0] node19710;
	wire [4-1:0] node19713;
	wire [4-1:0] node19714;
	wire [4-1:0] node19715;
	wire [4-1:0] node19716;
	wire [4-1:0] node19717;
	wire [4-1:0] node19718;
	wire [4-1:0] node19719;
	wire [4-1:0] node19723;
	wire [4-1:0] node19726;
	wire [4-1:0] node19728;
	wire [4-1:0] node19729;
	wire [4-1:0] node19732;
	wire [4-1:0] node19735;
	wire [4-1:0] node19736;
	wire [4-1:0] node19737;
	wire [4-1:0] node19739;
	wire [4-1:0] node19742;
	wire [4-1:0] node19744;
	wire [4-1:0] node19747;
	wire [4-1:0] node19749;
	wire [4-1:0] node19750;
	wire [4-1:0] node19753;
	wire [4-1:0] node19756;
	wire [4-1:0] node19757;
	wire [4-1:0] node19758;
	wire [4-1:0] node19759;
	wire [4-1:0] node19760;
	wire [4-1:0] node19764;
	wire [4-1:0] node19765;
	wire [4-1:0] node19769;
	wire [4-1:0] node19770;
	wire [4-1:0] node19772;
	wire [4-1:0] node19775;
	wire [4-1:0] node19776;
	wire [4-1:0] node19780;
	wire [4-1:0] node19781;
	wire [4-1:0] node19782;
	wire [4-1:0] node19785;
	wire [4-1:0] node19786;
	wire [4-1:0] node19790;
	wire [4-1:0] node19791;
	wire [4-1:0] node19793;
	wire [4-1:0] node19796;
	wire [4-1:0] node19798;
	wire [4-1:0] node19801;
	wire [4-1:0] node19802;
	wire [4-1:0] node19803;
	wire [4-1:0] node19804;
	wire [4-1:0] node19805;
	wire [4-1:0] node19807;
	wire [4-1:0] node19810;
	wire [4-1:0] node19812;
	wire [4-1:0] node19815;
	wire [4-1:0] node19816;
	wire [4-1:0] node19817;
	wire [4-1:0] node19820;
	wire [4-1:0] node19824;
	wire [4-1:0] node19825;
	wire [4-1:0] node19826;
	wire [4-1:0] node19827;
	wire [4-1:0] node19830;
	wire [4-1:0] node19833;
	wire [4-1:0] node19836;
	wire [4-1:0] node19838;
	wire [4-1:0] node19841;
	wire [4-1:0] node19842;
	wire [4-1:0] node19843;
	wire [4-1:0] node19844;
	wire [4-1:0] node19846;
	wire [4-1:0] node19849;
	wire [4-1:0] node19850;
	wire [4-1:0] node19854;
	wire [4-1:0] node19855;
	wire [4-1:0] node19857;
	wire [4-1:0] node19861;
	wire [4-1:0] node19862;
	wire [4-1:0] node19863;
	wire [4-1:0] node19867;
	wire [4-1:0] node19869;
	wire [4-1:0] node19870;
	wire [4-1:0] node19874;
	wire [4-1:0] node19875;
	wire [4-1:0] node19876;
	wire [4-1:0] node19877;
	wire [4-1:0] node19878;
	wire [4-1:0] node19879;
	wire [4-1:0] node19880;
	wire [4-1:0] node19881;
	wire [4-1:0] node19882;
	wire [4-1:0] node19883;
	wire [4-1:0] node19884;
	wire [4-1:0] node19887;
	wire [4-1:0] node19891;
	wire [4-1:0] node19892;
	wire [4-1:0] node19893;
	wire [4-1:0] node19896;
	wire [4-1:0] node19899;
	wire [4-1:0] node19902;
	wire [4-1:0] node19903;
	wire [4-1:0] node19905;
	wire [4-1:0] node19906;
	wire [4-1:0] node19909;
	wire [4-1:0] node19912;
	wire [4-1:0] node19913;
	wire [4-1:0] node19914;
	wire [4-1:0] node19917;
	wire [4-1:0] node19920;
	wire [4-1:0] node19921;
	wire [4-1:0] node19925;
	wire [4-1:0] node19926;
	wire [4-1:0] node19927;
	wire [4-1:0] node19928;
	wire [4-1:0] node19930;
	wire [4-1:0] node19933;
	wire [4-1:0] node19934;
	wire [4-1:0] node19937;
	wire [4-1:0] node19940;
	wire [4-1:0] node19941;
	wire [4-1:0] node19942;
	wire [4-1:0] node19946;
	wire [4-1:0] node19947;
	wire [4-1:0] node19951;
	wire [4-1:0] node19952;
	wire [4-1:0] node19953;
	wire [4-1:0] node19956;
	wire [4-1:0] node19957;
	wire [4-1:0] node19961;
	wire [4-1:0] node19962;
	wire [4-1:0] node19965;
	wire [4-1:0] node19966;
	wire [4-1:0] node19970;
	wire [4-1:0] node19971;
	wire [4-1:0] node19972;
	wire [4-1:0] node19973;
	wire [4-1:0] node19974;
	wire [4-1:0] node19975;
	wire [4-1:0] node19979;
	wire [4-1:0] node19982;
	wire [4-1:0] node19983;
	wire [4-1:0] node19984;
	wire [4-1:0] node19988;
	wire [4-1:0] node19989;
	wire [4-1:0] node19992;
	wire [4-1:0] node19995;
	wire [4-1:0] node19996;
	wire [4-1:0] node19997;
	wire [4-1:0] node19998;
	wire [4-1:0] node20002;
	wire [4-1:0] node20005;
	wire [4-1:0] node20007;
	wire [4-1:0] node20008;
	wire [4-1:0] node20011;
	wire [4-1:0] node20014;
	wire [4-1:0] node20015;
	wire [4-1:0] node20016;
	wire [4-1:0] node20017;
	wire [4-1:0] node20019;
	wire [4-1:0] node20023;
	wire [4-1:0] node20024;
	wire [4-1:0] node20027;
	wire [4-1:0] node20028;
	wire [4-1:0] node20032;
	wire [4-1:0] node20033;
	wire [4-1:0] node20034;
	wire [4-1:0] node20036;
	wire [4-1:0] node20039;
	wire [4-1:0] node20042;
	wire [4-1:0] node20043;
	wire [4-1:0] node20045;
	wire [4-1:0] node20048;
	wire [4-1:0] node20049;
	wire [4-1:0] node20052;
	wire [4-1:0] node20055;
	wire [4-1:0] node20056;
	wire [4-1:0] node20057;
	wire [4-1:0] node20058;
	wire [4-1:0] node20059;
	wire [4-1:0] node20060;
	wire [4-1:0] node20061;
	wire [4-1:0] node20065;
	wire [4-1:0] node20068;
	wire [4-1:0] node20069;
	wire [4-1:0] node20070;
	wire [4-1:0] node20074;
	wire [4-1:0] node20075;
	wire [4-1:0] node20079;
	wire [4-1:0] node20080;
	wire [4-1:0] node20082;
	wire [4-1:0] node20085;
	wire [4-1:0] node20087;
	wire [4-1:0] node20090;
	wire [4-1:0] node20091;
	wire [4-1:0] node20092;
	wire [4-1:0] node20093;
	wire [4-1:0] node20094;
	wire [4-1:0] node20097;
	wire [4-1:0] node20100;
	wire [4-1:0] node20102;
	wire [4-1:0] node20105;
	wire [4-1:0] node20106;
	wire [4-1:0] node20107;
	wire [4-1:0] node20111;
	wire [4-1:0] node20112;
	wire [4-1:0] node20115;
	wire [4-1:0] node20118;
	wire [4-1:0] node20119;
	wire [4-1:0] node20120;
	wire [4-1:0] node20121;
	wire [4-1:0] node20124;
	wire [4-1:0] node20127;
	wire [4-1:0] node20128;
	wire [4-1:0] node20132;
	wire [4-1:0] node20133;
	wire [4-1:0] node20136;
	wire [4-1:0] node20137;
	wire [4-1:0] node20141;
	wire [4-1:0] node20142;
	wire [4-1:0] node20143;
	wire [4-1:0] node20144;
	wire [4-1:0] node20146;
	wire [4-1:0] node20148;
	wire [4-1:0] node20151;
	wire [4-1:0] node20153;
	wire [4-1:0] node20154;
	wire [4-1:0] node20157;
	wire [4-1:0] node20160;
	wire [4-1:0] node20161;
	wire [4-1:0] node20162;
	wire [4-1:0] node20164;
	wire [4-1:0] node20167;
	wire [4-1:0] node20169;
	wire [4-1:0] node20172;
	wire [4-1:0] node20173;
	wire [4-1:0] node20174;
	wire [4-1:0] node20178;
	wire [4-1:0] node20179;
	wire [4-1:0] node20182;
	wire [4-1:0] node20185;
	wire [4-1:0] node20186;
	wire [4-1:0] node20187;
	wire [4-1:0] node20189;
	wire [4-1:0] node20190;
	wire [4-1:0] node20194;
	wire [4-1:0] node20195;
	wire [4-1:0] node20196;
	wire [4-1:0] node20200;
	wire [4-1:0] node20202;
	wire [4-1:0] node20205;
	wire [4-1:0] node20206;
	wire [4-1:0] node20207;
	wire [4-1:0] node20209;
	wire [4-1:0] node20212;
	wire [4-1:0] node20214;
	wire [4-1:0] node20217;
	wire [4-1:0] node20218;
	wire [4-1:0] node20219;
	wire [4-1:0] node20223;
	wire [4-1:0] node20224;
	wire [4-1:0] node20227;
	wire [4-1:0] node20230;
	wire [4-1:0] node20231;
	wire [4-1:0] node20232;
	wire [4-1:0] node20233;
	wire [4-1:0] node20234;
	wire [4-1:0] node20235;
	wire [4-1:0] node20236;
	wire [4-1:0] node20237;
	wire [4-1:0] node20240;
	wire [4-1:0] node20243;
	wire [4-1:0] node20244;
	wire [4-1:0] node20247;
	wire [4-1:0] node20250;
	wire [4-1:0] node20251;
	wire [4-1:0] node20252;
	wire [4-1:0] node20256;
	wire [4-1:0] node20257;
	wire [4-1:0] node20260;
	wire [4-1:0] node20263;
	wire [4-1:0] node20264;
	wire [4-1:0] node20265;
	wire [4-1:0] node20266;
	wire [4-1:0] node20270;
	wire [4-1:0] node20273;
	wire [4-1:0] node20274;
	wire [4-1:0] node20275;
	wire [4-1:0] node20278;
	wire [4-1:0] node20281;
	wire [4-1:0] node20284;
	wire [4-1:0] node20285;
	wire [4-1:0] node20286;
	wire [4-1:0] node20287;
	wire [4-1:0] node20290;
	wire [4-1:0] node20293;
	wire [4-1:0] node20294;
	wire [4-1:0] node20298;
	wire [4-1:0] node20299;
	wire [4-1:0] node20300;
	wire [4-1:0] node20301;
	wire [4-1:0] node20304;
	wire [4-1:0] node20307;
	wire [4-1:0] node20309;
	wire [4-1:0] node20312;
	wire [4-1:0] node20313;
	wire [4-1:0] node20314;
	wire [4-1:0] node20317;
	wire [4-1:0] node20320;
	wire [4-1:0] node20321;
	wire [4-1:0] node20324;
	wire [4-1:0] node20327;
	wire [4-1:0] node20328;
	wire [4-1:0] node20329;
	wire [4-1:0] node20330;
	wire [4-1:0] node20331;
	wire [4-1:0] node20333;
	wire [4-1:0] node20336;
	wire [4-1:0] node20338;
	wire [4-1:0] node20341;
	wire [4-1:0] node20342;
	wire [4-1:0] node20343;
	wire [4-1:0] node20346;
	wire [4-1:0] node20350;
	wire [4-1:0] node20351;
	wire [4-1:0] node20352;
	wire [4-1:0] node20353;
	wire [4-1:0] node20358;
	wire [4-1:0] node20359;
	wire [4-1:0] node20360;
	wire [4-1:0] node20364;
	wire [4-1:0] node20366;
	wire [4-1:0] node20369;
	wire [4-1:0] node20370;
	wire [4-1:0] node20371;
	wire [4-1:0] node20372;
	wire [4-1:0] node20374;
	wire [4-1:0] node20377;
	wire [4-1:0] node20379;
	wire [4-1:0] node20382;
	wire [4-1:0] node20383;
	wire [4-1:0] node20384;
	wire [4-1:0] node20387;
	wire [4-1:0] node20390;
	wire [4-1:0] node20391;
	wire [4-1:0] node20395;
	wire [4-1:0] node20396;
	wire [4-1:0] node20397;
	wire [4-1:0] node20398;
	wire [4-1:0] node20402;
	wire [4-1:0] node20405;
	wire [4-1:0] node20406;
	wire [4-1:0] node20407;
	wire [4-1:0] node20410;
	wire [4-1:0] node20413;
	wire [4-1:0] node20415;
	wire [4-1:0] node20418;
	wire [4-1:0] node20419;
	wire [4-1:0] node20420;
	wire [4-1:0] node20421;
	wire [4-1:0] node20422;
	wire [4-1:0] node20423;
	wire [4-1:0] node20424;
	wire [4-1:0] node20427;
	wire [4-1:0] node20430;
	wire [4-1:0] node20431;
	wire [4-1:0] node20435;
	wire [4-1:0] node20436;
	wire [4-1:0] node20438;
	wire [4-1:0] node20441;
	wire [4-1:0] node20443;
	wire [4-1:0] node20446;
	wire [4-1:0] node20447;
	wire [4-1:0] node20448;
	wire [4-1:0] node20451;
	wire [4-1:0] node20454;
	wire [4-1:0] node20456;
	wire [4-1:0] node20459;
	wire [4-1:0] node20460;
	wire [4-1:0] node20461;
	wire [4-1:0] node20462;
	wire [4-1:0] node20464;
	wire [4-1:0] node20467;
	wire [4-1:0] node20468;
	wire [4-1:0] node20471;
	wire [4-1:0] node20474;
	wire [4-1:0] node20475;
	wire [4-1:0] node20477;
	wire [4-1:0] node20480;
	wire [4-1:0] node20481;
	wire [4-1:0] node20484;
	wire [4-1:0] node20487;
	wire [4-1:0] node20488;
	wire [4-1:0] node20489;
	wire [4-1:0] node20490;
	wire [4-1:0] node20495;
	wire [4-1:0] node20497;
	wire [4-1:0] node20498;
	wire [4-1:0] node20501;
	wire [4-1:0] node20504;
	wire [4-1:0] node20505;
	wire [4-1:0] node20506;
	wire [4-1:0] node20507;
	wire [4-1:0] node20508;
	wire [4-1:0] node20511;
	wire [4-1:0] node20512;
	wire [4-1:0] node20516;
	wire [4-1:0] node20517;
	wire [4-1:0] node20518;
	wire [4-1:0] node20522;
	wire [4-1:0] node20524;
	wire [4-1:0] node20527;
	wire [4-1:0] node20528;
	wire [4-1:0] node20530;
	wire [4-1:0] node20532;
	wire [4-1:0] node20535;
	wire [4-1:0] node20536;
	wire [4-1:0] node20538;
	wire [4-1:0] node20541;
	wire [4-1:0] node20542;
	wire [4-1:0] node20546;
	wire [4-1:0] node20547;
	wire [4-1:0] node20548;
	wire [4-1:0] node20549;
	wire [4-1:0] node20551;
	wire [4-1:0] node20554;
	wire [4-1:0] node20557;
	wire [4-1:0] node20558;
	wire [4-1:0] node20560;
	wire [4-1:0] node20563;
	wire [4-1:0] node20564;
	wire [4-1:0] node20567;
	wire [4-1:0] node20570;
	wire [4-1:0] node20571;
	wire [4-1:0] node20572;
	wire [4-1:0] node20573;
	wire [4-1:0] node20576;
	wire [4-1:0] node20579;
	wire [4-1:0] node20580;
	wire [4-1:0] node20583;
	wire [4-1:0] node20586;
	wire [4-1:0] node20587;
	wire [4-1:0] node20589;
	wire [4-1:0] node20592;
	wire [4-1:0] node20593;
	wire [4-1:0] node20597;
	wire [4-1:0] node20598;
	wire [4-1:0] node20599;
	wire [4-1:0] node20600;
	wire [4-1:0] node20601;
	wire [4-1:0] node20602;
	wire [4-1:0] node20603;
	wire [4-1:0] node20604;
	wire [4-1:0] node20605;
	wire [4-1:0] node20609;
	wire [4-1:0] node20610;
	wire [4-1:0] node20614;
	wire [4-1:0] node20615;
	wire [4-1:0] node20616;
	wire [4-1:0] node20620;
	wire [4-1:0] node20622;
	wire [4-1:0] node20625;
	wire [4-1:0] node20626;
	wire [4-1:0] node20627;
	wire [4-1:0] node20628;
	wire [4-1:0] node20632;
	wire [4-1:0] node20633;
	wire [4-1:0] node20637;
	wire [4-1:0] node20638;
	wire [4-1:0] node20639;
	wire [4-1:0] node20643;
	wire [4-1:0] node20644;
	wire [4-1:0] node20648;
	wire [4-1:0] node20649;
	wire [4-1:0] node20650;
	wire [4-1:0] node20651;
	wire [4-1:0] node20652;
	wire [4-1:0] node20656;
	wire [4-1:0] node20657;
	wire [4-1:0] node20660;
	wire [4-1:0] node20663;
	wire [4-1:0] node20664;
	wire [4-1:0] node20665;
	wire [4-1:0] node20669;
	wire [4-1:0] node20671;
	wire [4-1:0] node20674;
	wire [4-1:0] node20675;
	wire [4-1:0] node20676;
	wire [4-1:0] node20679;
	wire [4-1:0] node20680;
	wire [4-1:0] node20683;
	wire [4-1:0] node20686;
	wire [4-1:0] node20687;
	wire [4-1:0] node20688;
	wire [4-1:0] node20692;
	wire [4-1:0] node20693;
	wire [4-1:0] node20696;
	wire [4-1:0] node20699;
	wire [4-1:0] node20700;
	wire [4-1:0] node20701;
	wire [4-1:0] node20702;
	wire [4-1:0] node20703;
	wire [4-1:0] node20704;
	wire [4-1:0] node20708;
	wire [4-1:0] node20709;
	wire [4-1:0] node20712;
	wire [4-1:0] node20715;
	wire [4-1:0] node20716;
	wire [4-1:0] node20717;
	wire [4-1:0] node20720;
	wire [4-1:0] node20723;
	wire [4-1:0] node20726;
	wire [4-1:0] node20727;
	wire [4-1:0] node20728;
	wire [4-1:0] node20730;
	wire [4-1:0] node20734;
	wire [4-1:0] node20736;
	wire [4-1:0] node20739;
	wire [4-1:0] node20740;
	wire [4-1:0] node20741;
	wire [4-1:0] node20743;
	wire [4-1:0] node20744;
	wire [4-1:0] node20748;
	wire [4-1:0] node20749;
	wire [4-1:0] node20751;
	wire [4-1:0] node20755;
	wire [4-1:0] node20756;
	wire [4-1:0] node20757;
	wire [4-1:0] node20759;
	wire [4-1:0] node20762;
	wire [4-1:0] node20764;
	wire [4-1:0] node20767;
	wire [4-1:0] node20768;
	wire [4-1:0] node20770;
	wire [4-1:0] node20773;
	wire [4-1:0] node20776;
	wire [4-1:0] node20777;
	wire [4-1:0] node20778;
	wire [4-1:0] node20779;
	wire [4-1:0] node20780;
	wire [4-1:0] node20781;
	wire [4-1:0] node20782;
	wire [4-1:0] node20787;
	wire [4-1:0] node20788;
	wire [4-1:0] node20789;
	wire [4-1:0] node20793;
	wire [4-1:0] node20794;
	wire [4-1:0] node20797;
	wire [4-1:0] node20800;
	wire [4-1:0] node20801;
	wire [4-1:0] node20802;
	wire [4-1:0] node20804;
	wire [4-1:0] node20807;
	wire [4-1:0] node20808;
	wire [4-1:0] node20812;
	wire [4-1:0] node20813;
	wire [4-1:0] node20814;
	wire [4-1:0] node20817;
	wire [4-1:0] node20820;
	wire [4-1:0] node20821;
	wire [4-1:0] node20824;
	wire [4-1:0] node20827;
	wire [4-1:0] node20828;
	wire [4-1:0] node20829;
	wire [4-1:0] node20830;
	wire [4-1:0] node20832;
	wire [4-1:0] node20835;
	wire [4-1:0] node20837;
	wire [4-1:0] node20840;
	wire [4-1:0] node20841;
	wire [4-1:0] node20842;
	wire [4-1:0] node20846;
	wire [4-1:0] node20847;
	wire [4-1:0] node20851;
	wire [4-1:0] node20852;
	wire [4-1:0] node20853;
	wire [4-1:0] node20856;
	wire [4-1:0] node20859;
	wire [4-1:0] node20860;
	wire [4-1:0] node20861;
	wire [4-1:0] node20864;
	wire [4-1:0] node20867;
	wire [4-1:0] node20869;
	wire [4-1:0] node20872;
	wire [4-1:0] node20873;
	wire [4-1:0] node20874;
	wire [4-1:0] node20875;
	wire [4-1:0] node20876;
	wire [4-1:0] node20878;
	wire [4-1:0] node20881;
	wire [4-1:0] node20882;
	wire [4-1:0] node20886;
	wire [4-1:0] node20888;
	wire [4-1:0] node20890;
	wire [4-1:0] node20893;
	wire [4-1:0] node20894;
	wire [4-1:0] node20895;
	wire [4-1:0] node20897;
	wire [4-1:0] node20900;
	wire [4-1:0] node20901;
	wire [4-1:0] node20904;
	wire [4-1:0] node20907;
	wire [4-1:0] node20908;
	wire [4-1:0] node20909;
	wire [4-1:0] node20913;
	wire [4-1:0] node20916;
	wire [4-1:0] node20917;
	wire [4-1:0] node20918;
	wire [4-1:0] node20919;
	wire [4-1:0] node20922;
	wire [4-1:0] node20923;
	wire [4-1:0] node20926;
	wire [4-1:0] node20929;
	wire [4-1:0] node20930;
	wire [4-1:0] node20931;
	wire [4-1:0] node20934;
	wire [4-1:0] node20937;
	wire [4-1:0] node20940;
	wire [4-1:0] node20941;
	wire [4-1:0] node20942;
	wire [4-1:0] node20945;
	wire [4-1:0] node20947;
	wire [4-1:0] node20950;
	wire [4-1:0] node20951;
	wire [4-1:0] node20952;
	wire [4-1:0] node20955;
	wire [4-1:0] node20958;
	wire [4-1:0] node20960;
	wire [4-1:0] node20963;
	wire [4-1:0] node20964;
	wire [4-1:0] node20965;
	wire [4-1:0] node20966;
	wire [4-1:0] node20967;
	wire [4-1:0] node20968;
	wire [4-1:0] node20969;
	wire [4-1:0] node20971;
	wire [4-1:0] node20974;
	wire [4-1:0] node20975;
	wire [4-1:0] node20978;
	wire [4-1:0] node20981;
	wire [4-1:0] node20982;
	wire [4-1:0] node20984;
	wire [4-1:0] node20987;
	wire [4-1:0] node20988;
	wire [4-1:0] node20991;
	wire [4-1:0] node20994;
	wire [4-1:0] node20995;
	wire [4-1:0] node20996;
	wire [4-1:0] node20997;
	wire [4-1:0] node21000;
	wire [4-1:0] node21003;
	wire [4-1:0] node21004;
	wire [4-1:0] node21007;
	wire [4-1:0] node21010;
	wire [4-1:0] node21012;
	wire [4-1:0] node21015;
	wire [4-1:0] node21016;
	wire [4-1:0] node21017;
	wire [4-1:0] node21018;
	wire [4-1:0] node21019;
	wire [4-1:0] node21023;
	wire [4-1:0] node21024;
	wire [4-1:0] node21027;
	wire [4-1:0] node21030;
	wire [4-1:0] node21031;
	wire [4-1:0] node21032;
	wire [4-1:0] node21036;
	wire [4-1:0] node21037;
	wire [4-1:0] node21041;
	wire [4-1:0] node21042;
	wire [4-1:0] node21043;
	wire [4-1:0] node21046;
	wire [4-1:0] node21047;
	wire [4-1:0] node21050;
	wire [4-1:0] node21053;
	wire [4-1:0] node21056;
	wire [4-1:0] node21057;
	wire [4-1:0] node21058;
	wire [4-1:0] node21059;
	wire [4-1:0] node21060;
	wire [4-1:0] node21061;
	wire [4-1:0] node21065;
	wire [4-1:0] node21067;
	wire [4-1:0] node21070;
	wire [4-1:0] node21071;
	wire [4-1:0] node21073;
	wire [4-1:0] node21076;
	wire [4-1:0] node21078;
	wire [4-1:0] node21081;
	wire [4-1:0] node21082;
	wire [4-1:0] node21083;
	wire [4-1:0] node21086;
	wire [4-1:0] node21087;
	wire [4-1:0] node21090;
	wire [4-1:0] node21093;
	wire [4-1:0] node21095;
	wire [4-1:0] node21096;
	wire [4-1:0] node21100;
	wire [4-1:0] node21101;
	wire [4-1:0] node21102;
	wire [4-1:0] node21103;
	wire [4-1:0] node21104;
	wire [4-1:0] node21107;
	wire [4-1:0] node21110;
	wire [4-1:0] node21111;
	wire [4-1:0] node21116;
	wire [4-1:0] node21117;
	wire [4-1:0] node21118;
	wire [4-1:0] node21120;
	wire [4-1:0] node21123;
	wire [4-1:0] node21125;
	wire [4-1:0] node21128;
	wire [4-1:0] node21129;
	wire [4-1:0] node21130;
	wire [4-1:0] node21134;
	wire [4-1:0] node21135;
	wire [4-1:0] node21139;
	wire [4-1:0] node21140;
	wire [4-1:0] node21141;
	wire [4-1:0] node21142;
	wire [4-1:0] node21143;
	wire [4-1:0] node21144;
	wire [4-1:0] node21145;
	wire [4-1:0] node21149;
	wire [4-1:0] node21152;
	wire [4-1:0] node21153;
	wire [4-1:0] node21154;
	wire [4-1:0] node21158;
	wire [4-1:0] node21160;
	wire [4-1:0] node21163;
	wire [4-1:0] node21164;
	wire [4-1:0] node21165;
	wire [4-1:0] node21166;
	wire [4-1:0] node21170;
	wire [4-1:0] node21171;
	wire [4-1:0] node21175;
	wire [4-1:0] node21176;
	wire [4-1:0] node21178;
	wire [4-1:0] node21181;
	wire [4-1:0] node21182;
	wire [4-1:0] node21186;
	wire [4-1:0] node21187;
	wire [4-1:0] node21188;
	wire [4-1:0] node21189;
	wire [4-1:0] node21190;
	wire [4-1:0] node21194;
	wire [4-1:0] node21196;
	wire [4-1:0] node21199;
	wire [4-1:0] node21201;
	wire [4-1:0] node21202;
	wire [4-1:0] node21205;
	wire [4-1:0] node21208;
	wire [4-1:0] node21209;
	wire [4-1:0] node21210;
	wire [4-1:0] node21211;
	wire [4-1:0] node21215;
	wire [4-1:0] node21219;
	wire [4-1:0] node21220;
	wire [4-1:0] node21221;
	wire [4-1:0] node21222;
	wire [4-1:0] node21223;
	wire [4-1:0] node21224;
	wire [4-1:0] node21227;
	wire [4-1:0] node21230;
	wire [4-1:0] node21231;
	wire [4-1:0] node21235;
	wire [4-1:0] node21236;
	wire [4-1:0] node21238;
	wire [4-1:0] node21241;
	wire [4-1:0] node21244;
	wire [4-1:0] node21245;
	wire [4-1:0] node21246;
	wire [4-1:0] node21247;
	wire [4-1:0] node21251;
	wire [4-1:0] node21254;
	wire [4-1:0] node21255;
	wire [4-1:0] node21256;
	wire [4-1:0] node21259;
	wire [4-1:0] node21262;
	wire [4-1:0] node21264;
	wire [4-1:0] node21267;
	wire [4-1:0] node21268;
	wire [4-1:0] node21269;
	wire [4-1:0] node21270;
	wire [4-1:0] node21272;
	wire [4-1:0] node21275;
	wire [4-1:0] node21277;
	wire [4-1:0] node21280;
	wire [4-1:0] node21281;
	wire [4-1:0] node21282;
	wire [4-1:0] node21285;
	wire [4-1:0] node21288;
	wire [4-1:0] node21289;
	wire [4-1:0] node21293;
	wire [4-1:0] node21294;
	wire [4-1:0] node21295;
	wire [4-1:0] node21296;
	wire [4-1:0] node21299;
	wire [4-1:0] node21302;
	wire [4-1:0] node21303;
	wire [4-1:0] node21307;
	wire [4-1:0] node21308;
	wire [4-1:0] node21309;
	wire [4-1:0] node21312;
	wire [4-1:0] node21315;
	wire [4-1:0] node21316;
	wire [4-1:0] node21320;
	wire [4-1:0] node21321;
	wire [4-1:0] node21322;
	wire [4-1:0] node21323;
	wire [4-1:0] node21324;
	wire [4-1:0] node21325;
	wire [4-1:0] node21326;
	wire [4-1:0] node21327;
	wire [4-1:0] node21328;
	wire [4-1:0] node21329;
	wire [4-1:0] node21333;
	wire [4-1:0] node21334;
	wire [4-1:0] node21337;
	wire [4-1:0] node21340;
	wire [4-1:0] node21341;
	wire [4-1:0] node21342;
	wire [4-1:0] node21345;
	wire [4-1:0] node21348;
	wire [4-1:0] node21351;
	wire [4-1:0] node21352;
	wire [4-1:0] node21353;
	wire [4-1:0] node21356;
	wire [4-1:0] node21358;
	wire [4-1:0] node21361;
	wire [4-1:0] node21362;
	wire [4-1:0] node21363;
	wire [4-1:0] node21366;
	wire [4-1:0] node21369;
	wire [4-1:0] node21370;
	wire [4-1:0] node21373;
	wire [4-1:0] node21376;
	wire [4-1:0] node21377;
	wire [4-1:0] node21378;
	wire [4-1:0] node21380;
	wire [4-1:0] node21382;
	wire [4-1:0] node21385;
	wire [4-1:0] node21386;
	wire [4-1:0] node21387;
	wire [4-1:0] node21390;
	wire [4-1:0] node21393;
	wire [4-1:0] node21394;
	wire [4-1:0] node21398;
	wire [4-1:0] node21399;
	wire [4-1:0] node21400;
	wire [4-1:0] node21401;
	wire [4-1:0] node21406;
	wire [4-1:0] node21407;
	wire [4-1:0] node21408;
	wire [4-1:0] node21411;
	wire [4-1:0] node21414;
	wire [4-1:0] node21416;
	wire [4-1:0] node21419;
	wire [4-1:0] node21420;
	wire [4-1:0] node21421;
	wire [4-1:0] node21422;
	wire [4-1:0] node21424;
	wire [4-1:0] node21425;
	wire [4-1:0] node21428;
	wire [4-1:0] node21431;
	wire [4-1:0] node21432;
	wire [4-1:0] node21433;
	wire [4-1:0] node21437;
	wire [4-1:0] node21439;
	wire [4-1:0] node21442;
	wire [4-1:0] node21443;
	wire [4-1:0] node21444;
	wire [4-1:0] node21446;
	wire [4-1:0] node21449;
	wire [4-1:0] node21452;
	wire [4-1:0] node21453;
	wire [4-1:0] node21455;
	wire [4-1:0] node21458;
	wire [4-1:0] node21460;
	wire [4-1:0] node21463;
	wire [4-1:0] node21464;
	wire [4-1:0] node21465;
	wire [4-1:0] node21466;
	wire [4-1:0] node21468;
	wire [4-1:0] node21471;
	wire [4-1:0] node21473;
	wire [4-1:0] node21476;
	wire [4-1:0] node21477;
	wire [4-1:0] node21478;
	wire [4-1:0] node21481;
	wire [4-1:0] node21485;
	wire [4-1:0] node21486;
	wire [4-1:0] node21487;
	wire [4-1:0] node21488;
	wire [4-1:0] node21492;
	wire [4-1:0] node21493;
	wire [4-1:0] node21497;
	wire [4-1:0] node21498;
	wire [4-1:0] node21500;
	wire [4-1:0] node21503;
	wire [4-1:0] node21504;
	wire [4-1:0] node21507;
	wire [4-1:0] node21510;
	wire [4-1:0] node21511;
	wire [4-1:0] node21512;
	wire [4-1:0] node21513;
	wire [4-1:0] node21514;
	wire [4-1:0] node21515;
	wire [4-1:0] node21516;
	wire [4-1:0] node21519;
	wire [4-1:0] node21523;
	wire [4-1:0] node21524;
	wire [4-1:0] node21525;
	wire [4-1:0] node21528;
	wire [4-1:0] node21531;
	wire [4-1:0] node21534;
	wire [4-1:0] node21535;
	wire [4-1:0] node21536;
	wire [4-1:0] node21537;
	wire [4-1:0] node21541;
	wire [4-1:0] node21542;
	wire [4-1:0] node21545;
	wire [4-1:0] node21548;
	wire [4-1:0] node21549;
	wire [4-1:0] node21551;
	wire [4-1:0] node21554;
	wire [4-1:0] node21556;
	wire [4-1:0] node21559;
	wire [4-1:0] node21560;
	wire [4-1:0] node21561;
	wire [4-1:0] node21562;
	wire [4-1:0] node21563;
	wire [4-1:0] node21567;
	wire [4-1:0] node21568;
	wire [4-1:0] node21572;
	wire [4-1:0] node21573;
	wire [4-1:0] node21575;
	wire [4-1:0] node21578;
	wire [4-1:0] node21580;
	wire [4-1:0] node21583;
	wire [4-1:0] node21584;
	wire [4-1:0] node21585;
	wire [4-1:0] node21586;
	wire [4-1:0] node21589;
	wire [4-1:0] node21592;
	wire [4-1:0] node21595;
	wire [4-1:0] node21596;
	wire [4-1:0] node21598;
	wire [4-1:0] node21602;
	wire [4-1:0] node21603;
	wire [4-1:0] node21604;
	wire [4-1:0] node21605;
	wire [4-1:0] node21607;
	wire [4-1:0] node21608;
	wire [4-1:0] node21611;
	wire [4-1:0] node21614;
	wire [4-1:0] node21615;
	wire [4-1:0] node21616;
	wire [4-1:0] node21619;
	wire [4-1:0] node21622;
	wire [4-1:0] node21623;
	wire [4-1:0] node21626;
	wire [4-1:0] node21629;
	wire [4-1:0] node21630;
	wire [4-1:0] node21631;
	wire [4-1:0] node21633;
	wire [4-1:0] node21636;
	wire [4-1:0] node21638;
	wire [4-1:0] node21641;
	wire [4-1:0] node21642;
	wire [4-1:0] node21643;
	wire [4-1:0] node21646;
	wire [4-1:0] node21649;
	wire [4-1:0] node21651;
	wire [4-1:0] node21654;
	wire [4-1:0] node21655;
	wire [4-1:0] node21656;
	wire [4-1:0] node21657;
	wire [4-1:0] node21659;
	wire [4-1:0] node21663;
	wire [4-1:0] node21664;
	wire [4-1:0] node21667;
	wire [4-1:0] node21670;
	wire [4-1:0] node21671;
	wire [4-1:0] node21672;
	wire [4-1:0] node21673;
	wire [4-1:0] node21677;
	wire [4-1:0] node21680;
	wire [4-1:0] node21681;
	wire [4-1:0] node21682;
	wire [4-1:0] node21686;
	wire [4-1:0] node21687;
	wire [4-1:0] node21690;
	wire [4-1:0] node21693;
	wire [4-1:0] node21694;
	wire [4-1:0] node21695;
	wire [4-1:0] node21696;
	wire [4-1:0] node21697;
	wire [4-1:0] node21698;
	wire [4-1:0] node21699;
	wire [4-1:0] node21701;
	wire [4-1:0] node21704;
	wire [4-1:0] node21707;
	wire [4-1:0] node21708;
	wire [4-1:0] node21709;
	wire [4-1:0] node21713;
	wire [4-1:0] node21716;
	wire [4-1:0] node21717;
	wire [4-1:0] node21718;
	wire [4-1:0] node21720;
	wire [4-1:0] node21723;
	wire [4-1:0] node21724;
	wire [4-1:0] node21728;
	wire [4-1:0] node21729;
	wire [4-1:0] node21732;
	wire [4-1:0] node21734;
	wire [4-1:0] node21737;
	wire [4-1:0] node21738;
	wire [4-1:0] node21739;
	wire [4-1:0] node21740;
	wire [4-1:0] node21742;
	wire [4-1:0] node21746;
	wire [4-1:0] node21747;
	wire [4-1:0] node21748;
	wire [4-1:0] node21752;
	wire [4-1:0] node21753;
	wire [4-1:0] node21756;
	wire [4-1:0] node21759;
	wire [4-1:0] node21760;
	wire [4-1:0] node21761;
	wire [4-1:0] node21763;
	wire [4-1:0] node21766;
	wire [4-1:0] node21767;
	wire [4-1:0] node21771;
	wire [4-1:0] node21772;
	wire [4-1:0] node21773;
	wire [4-1:0] node21776;
	wire [4-1:0] node21780;
	wire [4-1:0] node21781;
	wire [4-1:0] node21782;
	wire [4-1:0] node21783;
	wire [4-1:0] node21784;
	wire [4-1:0] node21785;
	wire [4-1:0] node21789;
	wire [4-1:0] node21791;
	wire [4-1:0] node21794;
	wire [4-1:0] node21795;
	wire [4-1:0] node21797;
	wire [4-1:0] node21800;
	wire [4-1:0] node21801;
	wire [4-1:0] node21804;
	wire [4-1:0] node21807;
	wire [4-1:0] node21808;
	wire [4-1:0] node21809;
	wire [4-1:0] node21812;
	wire [4-1:0] node21813;
	wire [4-1:0] node21817;
	wire [4-1:0] node21818;
	wire [4-1:0] node21819;
	wire [4-1:0] node21823;
	wire [4-1:0] node21826;
	wire [4-1:0] node21827;
	wire [4-1:0] node21828;
	wire [4-1:0] node21829;
	wire [4-1:0] node21831;
	wire [4-1:0] node21836;
	wire [4-1:0] node21837;
	wire [4-1:0] node21838;
	wire [4-1:0] node21840;
	wire [4-1:0] node21843;
	wire [4-1:0] node21845;
	wire [4-1:0] node21848;
	wire [4-1:0] node21850;
	wire [4-1:0] node21851;
	wire [4-1:0] node21854;
	wire [4-1:0] node21857;
	wire [4-1:0] node21858;
	wire [4-1:0] node21859;
	wire [4-1:0] node21860;
	wire [4-1:0] node21861;
	wire [4-1:0] node21863;
	wire [4-1:0] node21864;
	wire [4-1:0] node21867;
	wire [4-1:0] node21870;
	wire [4-1:0] node21871;
	wire [4-1:0] node21872;
	wire [4-1:0] node21875;
	wire [4-1:0] node21878;
	wire [4-1:0] node21879;
	wire [4-1:0] node21883;
	wire [4-1:0] node21884;
	wire [4-1:0] node21885;
	wire [4-1:0] node21886;
	wire [4-1:0] node21889;
	wire [4-1:0] node21892;
	wire [4-1:0] node21895;
	wire [4-1:0] node21896;
	wire [4-1:0] node21897;
	wire [4-1:0] node21901;
	wire [4-1:0] node21904;
	wire [4-1:0] node21905;
	wire [4-1:0] node21906;
	wire [4-1:0] node21908;
	wire [4-1:0] node21910;
	wire [4-1:0] node21913;
	wire [4-1:0] node21914;
	wire [4-1:0] node21917;
	wire [4-1:0] node21919;
	wire [4-1:0] node21922;
	wire [4-1:0] node21923;
	wire [4-1:0] node21924;
	wire [4-1:0] node21925;
	wire [4-1:0] node21929;
	wire [4-1:0] node21930;
	wire [4-1:0] node21933;
	wire [4-1:0] node21936;
	wire [4-1:0] node21937;
	wire [4-1:0] node21940;
	wire [4-1:0] node21941;
	wire [4-1:0] node21944;
	wire [4-1:0] node21947;
	wire [4-1:0] node21948;
	wire [4-1:0] node21949;
	wire [4-1:0] node21950;
	wire [4-1:0] node21951;
	wire [4-1:0] node21952;
	wire [4-1:0] node21956;
	wire [4-1:0] node21957;
	wire [4-1:0] node21961;
	wire [4-1:0] node21962;
	wire [4-1:0] node21964;
	wire [4-1:0] node21968;
	wire [4-1:0] node21969;
	wire [4-1:0] node21970;
	wire [4-1:0] node21973;
	wire [4-1:0] node21975;
	wire [4-1:0] node21978;
	wire [4-1:0] node21979;
	wire [4-1:0] node21980;
	wire [4-1:0] node21985;
	wire [4-1:0] node21986;
	wire [4-1:0] node21987;
	wire [4-1:0] node21988;
	wire [4-1:0] node21989;
	wire [4-1:0] node21993;
	wire [4-1:0] node21996;
	wire [4-1:0] node21997;
	wire [4-1:0] node21998;
	wire [4-1:0] node22001;
	wire [4-1:0] node22004;
	wire [4-1:0] node22007;
	wire [4-1:0] node22008;
	wire [4-1:0] node22009;
	wire [4-1:0] node22010;
	wire [4-1:0] node22014;
	wire [4-1:0] node22017;
	wire [4-1:0] node22019;
	wire [4-1:0] node22022;
	wire [4-1:0] node22023;
	wire [4-1:0] node22024;
	wire [4-1:0] node22025;
	wire [4-1:0] node22026;
	wire [4-1:0] node22027;
	wire [4-1:0] node22028;
	wire [4-1:0] node22029;
	wire [4-1:0] node22030;
	wire [4-1:0] node22033;
	wire [4-1:0] node22037;
	wire [4-1:0] node22038;
	wire [4-1:0] node22040;
	wire [4-1:0] node22043;
	wire [4-1:0] node22045;
	wire [4-1:0] node22048;
	wire [4-1:0] node22049;
	wire [4-1:0] node22050;
	wire [4-1:0] node22053;
	wire [4-1:0] node22055;
	wire [4-1:0] node22058;
	wire [4-1:0] node22059;
	wire [4-1:0] node22062;
	wire [4-1:0] node22063;
	wire [4-1:0] node22067;
	wire [4-1:0] node22068;
	wire [4-1:0] node22069;
	wire [4-1:0] node22070;
	wire [4-1:0] node22071;
	wire [4-1:0] node22076;
	wire [4-1:0] node22078;
	wire [4-1:0] node22080;
	wire [4-1:0] node22083;
	wire [4-1:0] node22084;
	wire [4-1:0] node22085;
	wire [4-1:0] node22087;
	wire [4-1:0] node22091;
	wire [4-1:0] node22092;
	wire [4-1:0] node22095;
	wire [4-1:0] node22096;
	wire [4-1:0] node22100;
	wire [4-1:0] node22101;
	wire [4-1:0] node22102;
	wire [4-1:0] node22103;
	wire [4-1:0] node22104;
	wire [4-1:0] node22105;
	wire [4-1:0] node22108;
	wire [4-1:0] node22111;
	wire [4-1:0] node22113;
	wire [4-1:0] node22116;
	wire [4-1:0] node22118;
	wire [4-1:0] node22119;
	wire [4-1:0] node22122;
	wire [4-1:0] node22125;
	wire [4-1:0] node22126;
	wire [4-1:0] node22127;
	wire [4-1:0] node22130;
	wire [4-1:0] node22131;
	wire [4-1:0] node22135;
	wire [4-1:0] node22136;
	wire [4-1:0] node22138;
	wire [4-1:0] node22141;
	wire [4-1:0] node22142;
	wire [4-1:0] node22146;
	wire [4-1:0] node22147;
	wire [4-1:0] node22148;
	wire [4-1:0] node22149;
	wire [4-1:0] node22152;
	wire [4-1:0] node22155;
	wire [4-1:0] node22156;
	wire [4-1:0] node22158;
	wire [4-1:0] node22161;
	wire [4-1:0] node22163;
	wire [4-1:0] node22166;
	wire [4-1:0] node22167;
	wire [4-1:0] node22168;
	wire [4-1:0] node22170;
	wire [4-1:0] node22174;
	wire [4-1:0] node22175;
	wire [4-1:0] node22176;
	wire [4-1:0] node22180;
	wire [4-1:0] node22183;
	wire [4-1:0] node22184;
	wire [4-1:0] node22185;
	wire [4-1:0] node22186;
	wire [4-1:0] node22187;
	wire [4-1:0] node22188;
	wire [4-1:0] node22190;
	wire [4-1:0] node22193;
	wire [4-1:0] node22194;
	wire [4-1:0] node22198;
	wire [4-1:0] node22199;
	wire [4-1:0] node22201;
	wire [4-1:0] node22204;
	wire [4-1:0] node22205;
	wire [4-1:0] node22208;
	wire [4-1:0] node22211;
	wire [4-1:0] node22212;
	wire [4-1:0] node22213;
	wire [4-1:0] node22214;
	wire [4-1:0] node22218;
	wire [4-1:0] node22220;
	wire [4-1:0] node22223;
	wire [4-1:0] node22224;
	wire [4-1:0] node22225;
	wire [4-1:0] node22228;
	wire [4-1:0] node22232;
	wire [4-1:0] node22233;
	wire [4-1:0] node22234;
	wire [4-1:0] node22236;
	wire [4-1:0] node22237;
	wire [4-1:0] node22240;
	wire [4-1:0] node22243;
	wire [4-1:0] node22244;
	wire [4-1:0] node22248;
	wire [4-1:0] node22249;
	wire [4-1:0] node22250;
	wire [4-1:0] node22252;
	wire [4-1:0] node22255;
	wire [4-1:0] node22257;
	wire [4-1:0] node22260;
	wire [4-1:0] node22261;
	wire [4-1:0] node22262;
	wire [4-1:0] node22266;
	wire [4-1:0] node22267;
	wire [4-1:0] node22270;
	wire [4-1:0] node22273;
	wire [4-1:0] node22274;
	wire [4-1:0] node22275;
	wire [4-1:0] node22276;
	wire [4-1:0] node22277;
	wire [4-1:0] node22278;
	wire [4-1:0] node22281;
	wire [4-1:0] node22284;
	wire [4-1:0] node22285;
	wire [4-1:0] node22288;
	wire [4-1:0] node22291;
	wire [4-1:0] node22292;
	wire [4-1:0] node22294;
	wire [4-1:0] node22297;
	wire [4-1:0] node22298;
	wire [4-1:0] node22302;
	wire [4-1:0] node22303;
	wire [4-1:0] node22304;
	wire [4-1:0] node22305;
	wire [4-1:0] node22309;
	wire [4-1:0] node22310;
	wire [4-1:0] node22313;
	wire [4-1:0] node22316;
	wire [4-1:0] node22317;
	wire [4-1:0] node22320;
	wire [4-1:0] node22321;
	wire [4-1:0] node22324;
	wire [4-1:0] node22327;
	wire [4-1:0] node22328;
	wire [4-1:0] node22329;
	wire [4-1:0] node22330;
	wire [4-1:0] node22331;
	wire [4-1:0] node22334;
	wire [4-1:0] node22337;
	wire [4-1:0] node22338;
	wire [4-1:0] node22342;
	wire [4-1:0] node22343;
	wire [4-1:0] node22344;
	wire [4-1:0] node22347;
	wire [4-1:0] node22350;
	wire [4-1:0] node22351;
	wire [4-1:0] node22354;
	wire [4-1:0] node22357;
	wire [4-1:0] node22358;
	wire [4-1:0] node22359;
	wire [4-1:0] node22360;
	wire [4-1:0] node22363;
	wire [4-1:0] node22366;
	wire [4-1:0] node22367;
	wire [4-1:0] node22370;
	wire [4-1:0] node22373;
	wire [4-1:0] node22374;
	wire [4-1:0] node22375;
	wire [4-1:0] node22379;
	wire [4-1:0] node22380;
	wire [4-1:0] node22383;
	wire [4-1:0] node22386;
	wire [4-1:0] node22387;
	wire [4-1:0] node22388;
	wire [4-1:0] node22389;
	wire [4-1:0] node22390;
	wire [4-1:0] node22391;
	wire [4-1:0] node22392;
	wire [4-1:0] node22395;
	wire [4-1:0] node22396;
	wire [4-1:0] node22400;
	wire [4-1:0] node22401;
	wire [4-1:0] node22403;
	wire [4-1:0] node22406;
	wire [4-1:0] node22407;
	wire [4-1:0] node22411;
	wire [4-1:0] node22412;
	wire [4-1:0] node22413;
	wire [4-1:0] node22414;
	wire [4-1:0] node22417;
	wire [4-1:0] node22421;
	wire [4-1:0] node22422;
	wire [4-1:0] node22423;
	wire [4-1:0] node22426;
	wire [4-1:0] node22429;
	wire [4-1:0] node22430;
	wire [4-1:0] node22434;
	wire [4-1:0] node22435;
	wire [4-1:0] node22436;
	wire [4-1:0] node22437;
	wire [4-1:0] node22438;
	wire [4-1:0] node22442;
	wire [4-1:0] node22443;
	wire [4-1:0] node22446;
	wire [4-1:0] node22449;
	wire [4-1:0] node22450;
	wire [4-1:0] node22451;
	wire [4-1:0] node22455;
	wire [4-1:0] node22456;
	wire [4-1:0] node22460;
	wire [4-1:0] node22461;
	wire [4-1:0] node22462;
	wire [4-1:0] node22463;
	wire [4-1:0] node22467;
	wire [4-1:0] node22468;
	wire [4-1:0] node22471;
	wire [4-1:0] node22474;
	wire [4-1:0] node22475;
	wire [4-1:0] node22476;
	wire [4-1:0] node22479;
	wire [4-1:0] node22482;
	wire [4-1:0] node22483;
	wire [4-1:0] node22486;
	wire [4-1:0] node22489;
	wire [4-1:0] node22490;
	wire [4-1:0] node22491;
	wire [4-1:0] node22492;
	wire [4-1:0] node22493;
	wire [4-1:0] node22495;
	wire [4-1:0] node22498;
	wire [4-1:0] node22501;
	wire [4-1:0] node22503;
	wire [4-1:0] node22504;
	wire [4-1:0] node22507;
	wire [4-1:0] node22510;
	wire [4-1:0] node22511;
	wire [4-1:0] node22512;
	wire [4-1:0] node22513;
	wire [4-1:0] node22516;
	wire [4-1:0] node22519;
	wire [4-1:0] node22521;
	wire [4-1:0] node22524;
	wire [4-1:0] node22525;
	wire [4-1:0] node22526;
	wire [4-1:0] node22530;
	wire [4-1:0] node22531;
	wire [4-1:0] node22534;
	wire [4-1:0] node22537;
	wire [4-1:0] node22538;
	wire [4-1:0] node22539;
	wire [4-1:0] node22540;
	wire [4-1:0] node22542;
	wire [4-1:0] node22545;
	wire [4-1:0] node22546;
	wire [4-1:0] node22550;
	wire [4-1:0] node22551;
	wire [4-1:0] node22553;
	wire [4-1:0] node22556;
	wire [4-1:0] node22557;
	wire [4-1:0] node22560;
	wire [4-1:0] node22563;
	wire [4-1:0] node22564;
	wire [4-1:0] node22565;
	wire [4-1:0] node22566;
	wire [4-1:0] node22569;
	wire [4-1:0] node22572;
	wire [4-1:0] node22574;
	wire [4-1:0] node22577;
	wire [4-1:0] node22578;
	wire [4-1:0] node22580;
	wire [4-1:0] node22584;
	wire [4-1:0] node22585;
	wire [4-1:0] node22586;
	wire [4-1:0] node22587;
	wire [4-1:0] node22588;
	wire [4-1:0] node22589;
	wire [4-1:0] node22591;
	wire [4-1:0] node22594;
	wire [4-1:0] node22595;
	wire [4-1:0] node22599;
	wire [4-1:0] node22600;
	wire [4-1:0] node22602;
	wire [4-1:0] node22606;
	wire [4-1:0] node22607;
	wire [4-1:0] node22609;
	wire [4-1:0] node22610;
	wire [4-1:0] node22614;
	wire [4-1:0] node22615;
	wire [4-1:0] node22616;
	wire [4-1:0] node22619;
	wire [4-1:0] node22622;
	wire [4-1:0] node22623;
	wire [4-1:0] node22627;
	wire [4-1:0] node22628;
	wire [4-1:0] node22629;
	wire [4-1:0] node22632;
	wire [4-1:0] node22634;
	wire [4-1:0] node22635;
	wire [4-1:0] node22638;
	wire [4-1:0] node22641;
	wire [4-1:0] node22642;
	wire [4-1:0] node22643;
	wire [4-1:0] node22644;
	wire [4-1:0] node22647;
	wire [4-1:0] node22650;
	wire [4-1:0] node22651;
	wire [4-1:0] node22655;
	wire [4-1:0] node22656;
	wire [4-1:0] node22657;
	wire [4-1:0] node22661;
	wire [4-1:0] node22662;
	wire [4-1:0] node22665;
	wire [4-1:0] node22668;
	wire [4-1:0] node22669;
	wire [4-1:0] node22670;
	wire [4-1:0] node22671;
	wire [4-1:0] node22672;
	wire [4-1:0] node22673;
	wire [4-1:0] node22676;
	wire [4-1:0] node22679;
	wire [4-1:0] node22680;
	wire [4-1:0] node22683;
	wire [4-1:0] node22686;
	wire [4-1:0] node22687;
	wire [4-1:0] node22689;
	wire [4-1:0] node22692;
	wire [4-1:0] node22693;
	wire [4-1:0] node22696;
	wire [4-1:0] node22699;
	wire [4-1:0] node22700;
	wire [4-1:0] node22701;
	wire [4-1:0] node22703;
	wire [4-1:0] node22706;
	wire [4-1:0] node22707;
	wire [4-1:0] node22711;
	wire [4-1:0] node22712;
	wire [4-1:0] node22714;
	wire [4-1:0] node22717;
	wire [4-1:0] node22719;
	wire [4-1:0] node22722;
	wire [4-1:0] node22723;
	wire [4-1:0] node22724;
	wire [4-1:0] node22725;
	wire [4-1:0] node22726;
	wire [4-1:0] node22730;
	wire [4-1:0] node22731;
	wire [4-1:0] node22734;
	wire [4-1:0] node22737;
	wire [4-1:0] node22738;
	wire [4-1:0] node22739;
	wire [4-1:0] node22742;
	wire [4-1:0] node22745;
	wire [4-1:0] node22747;
	wire [4-1:0] node22750;
	wire [4-1:0] node22751;
	wire [4-1:0] node22752;
	wire [4-1:0] node22753;
	wire [4-1:0] node22757;
	wire [4-1:0] node22760;
	wire [4-1:0] node22761;
	wire [4-1:0] node22762;
	wire [4-1:0] node22766;
	wire [4-1:0] node22767;
	wire [4-1:0] node22770;

	assign outp = (inp[0]) ? node11270 : node1;
		assign node1 = (inp[4]) ? node5653 : node2;
			assign node2 = (inp[15]) ? node2824 : node3;
				assign node3 = (inp[5]) ? node1391 : node4;
					assign node4 = (inp[9]) ? node686 : node5;
						assign node5 = (inp[12]) ? node357 : node6;
							assign node6 = (inp[10]) ? node178 : node7;
								assign node7 = (inp[7]) ? node81 : node8;
									assign node8 = (inp[8]) ? node42 : node9;
										assign node9 = (inp[14]) ? node27 : node10;
											assign node10 = (inp[2]) ? node20 : node11;
												assign node11 = (inp[3]) ? node15 : node12;
													assign node12 = (inp[6]) ? 4'b0111 : 4'b1111;
													assign node15 = (inp[1]) ? 4'b1111 : node16;
														assign node16 = (inp[11]) ? 4'b0111 : 4'b0111;
												assign node20 = (inp[3]) ? 4'b1110 : node21;
													assign node21 = (inp[13]) ? 4'b1110 : node22;
														assign node22 = (inp[1]) ? 4'b0110 : 4'b1110;
											assign node27 = (inp[11]) ? node39 : node28;
												assign node28 = (inp[6]) ? node34 : node29;
													assign node29 = (inp[13]) ? node31 : 4'b1110;
														assign node31 = (inp[1]) ? 4'b0110 : 4'b1110;
													assign node34 = (inp[13]) ? node36 : 4'b0110;
														assign node36 = (inp[1]) ? 4'b1110 : 4'b0110;
												assign node39 = (inp[6]) ? 4'b1110 : 4'b0110;
										assign node42 = (inp[2]) ? node60 : node43;
											assign node43 = (inp[14]) ? node51 : node44;
												assign node44 = (inp[1]) ? node46 : 4'b1110;
													assign node46 = (inp[11]) ? node48 : 4'b0110;
														assign node48 = (inp[13]) ? 4'b0110 : 4'b0110;
												assign node51 = (inp[13]) ? node53 : 4'b0111;
													assign node53 = (inp[3]) ? node57 : node54;
														assign node54 = (inp[1]) ? 4'b1111 : 4'b0111;
														assign node57 = (inp[6]) ? 4'b0111 : 4'b1111;
											assign node60 = (inp[3]) ? node70 : node61;
												assign node61 = (inp[11]) ? 4'b1111 : node62;
													assign node62 = (inp[6]) ? node66 : node63;
														assign node63 = (inp[1]) ? 4'b0111 : 4'b1111;
														assign node66 = (inp[1]) ? 4'b1111 : 4'b0111;
												assign node70 = (inp[11]) ? node76 : node71;
													assign node71 = (inp[1]) ? node73 : 4'b1111;
														assign node73 = (inp[6]) ? 4'b1111 : 4'b0111;
													assign node76 = (inp[6]) ? 4'b0111 : node77;
														assign node77 = (inp[13]) ? 4'b1111 : 4'b0111;
									assign node81 = (inp[8]) ? node131 : node82;
										assign node82 = (inp[14]) ? node106 : node83;
											assign node83 = (inp[2]) ? node97 : node84;
												assign node84 = (inp[1]) ? node92 : node85;
													assign node85 = (inp[11]) ? node89 : node86;
														assign node86 = (inp[6]) ? 4'b0110 : 4'b1110;
														assign node89 = (inp[6]) ? 4'b1110 : 4'b0110;
													assign node92 = (inp[13]) ? node94 : 4'b0110;
														assign node94 = (inp[11]) ? 4'b1110 : 4'b0110;
												assign node97 = (inp[3]) ? 4'b0111 : node98;
													assign node98 = (inp[13]) ? node102 : node99;
														assign node99 = (inp[1]) ? 4'b1111 : 4'b0111;
														assign node102 = (inp[6]) ? 4'b1111 : 4'b0111;
											assign node106 = (inp[3]) ? node120 : node107;
												assign node107 = (inp[1]) ? node115 : node108;
													assign node108 = (inp[11]) ? node112 : node109;
														assign node109 = (inp[2]) ? 4'b0111 : 4'b0111;
														assign node112 = (inp[6]) ? 4'b0111 : 4'b1111;
													assign node115 = (inp[2]) ? 4'b0111 : node116;
														assign node116 = (inp[11]) ? 4'b1111 : 4'b0111;
												assign node120 = (inp[6]) ? node126 : node121;
													assign node121 = (inp[11]) ? 4'b1111 : node122;
														assign node122 = (inp[13]) ? 4'b0111 : 4'b0111;
													assign node126 = (inp[11]) ? node128 : 4'b1111;
														assign node128 = (inp[1]) ? 4'b0111 : 4'b0111;
										assign node131 = (inp[14]) ? node153 : node132;
											assign node132 = (inp[2]) ? node140 : node133;
												assign node133 = (inp[13]) ? node137 : node134;
													assign node134 = (inp[3]) ? 4'b1111 : 4'b0111;
													assign node137 = (inp[3]) ? 4'b0111 : 4'b1111;
												assign node140 = (inp[13]) ? node148 : node141;
													assign node141 = (inp[1]) ? node145 : node142;
														assign node142 = (inp[11]) ? 4'b0110 : 4'b1110;
														assign node145 = (inp[11]) ? 4'b1110 : 4'b0110;
													assign node148 = (inp[11]) ? 4'b0110 : node149;
														assign node149 = (inp[6]) ? 4'b1110 : 4'b0110;
											assign node153 = (inp[3]) ? node163 : node154;
												assign node154 = (inp[11]) ? node160 : node155;
													assign node155 = (inp[6]) ? node157 : 4'b0110;
														assign node157 = (inp[13]) ? 4'b1110 : 4'b0110;
													assign node160 = (inp[6]) ? 4'b0110 : 4'b1110;
												assign node163 = (inp[1]) ? node171 : node164;
													assign node164 = (inp[11]) ? node168 : node165;
														assign node165 = (inp[13]) ? 4'b0110 : 4'b1110;
														assign node168 = (inp[13]) ? 4'b0110 : 4'b0110;
													assign node171 = (inp[2]) ? node175 : node172;
														assign node172 = (inp[6]) ? 4'b0110 : 4'b1110;
														assign node175 = (inp[11]) ? 4'b1110 : 4'b1110;
								assign node178 = (inp[11]) ? node270 : node179;
									assign node179 = (inp[6]) ? node233 : node180;
										assign node180 = (inp[13]) ? node206 : node181;
											assign node181 = (inp[1]) ? node193 : node182;
												assign node182 = (inp[2]) ? node188 : node183;
													assign node183 = (inp[14]) ? node185 : 4'b1111;
														assign node185 = (inp[7]) ? 4'b1110 : 4'b1111;
													assign node188 = (inp[3]) ? 4'b1110 : node189;
														assign node189 = (inp[8]) ? 4'b1110 : 4'b1111;
												assign node193 = (inp[14]) ? node201 : node194;
													assign node194 = (inp[7]) ? node198 : node195;
														assign node195 = (inp[2]) ? 4'b1110 : 4'b1110;
														assign node198 = (inp[8]) ? 4'b0110 : 4'b1110;
													assign node201 = (inp[3]) ? node203 : 4'b0111;
														assign node203 = (inp[7]) ? 4'b0110 : 4'b0110;
											assign node206 = (inp[1]) ? node220 : node207;
												assign node207 = (inp[2]) ? node215 : node208;
													assign node208 = (inp[8]) ? node212 : node209;
														assign node209 = (inp[14]) ? 4'b1110 : 4'b1111;
														assign node212 = (inp[14]) ? 4'b0111 : 4'b1110;
													assign node215 = (inp[8]) ? node217 : 4'b0111;
														assign node217 = (inp[7]) ? 4'b0110 : 4'b0111;
												assign node220 = (inp[8]) ? node228 : node221;
													assign node221 = (inp[7]) ? node225 : node222;
														assign node222 = (inp[2]) ? 4'b0110 : 4'b0110;
														assign node225 = (inp[2]) ? 4'b0111 : 4'b0111;
													assign node228 = (inp[7]) ? node230 : 4'b0111;
														assign node230 = (inp[14]) ? 4'b0110 : 4'b0110;
										assign node233 = (inp[7]) ? node253 : node234;
											assign node234 = (inp[8]) ? node242 : node235;
												assign node235 = (inp[14]) ? 4'b0110 : node236;
													assign node236 = (inp[2]) ? 4'b0110 : node237;
														assign node237 = (inp[1]) ? 4'b0011 : 4'b0111;
												assign node242 = (inp[1]) ? node248 : node243;
													assign node243 = (inp[13]) ? node245 : 4'b0111;
														assign node245 = (inp[3]) ? 4'b0110 : 4'b1011;
													assign node248 = (inp[3]) ? 4'b1011 : node249;
														assign node249 = (inp[14]) ? 4'b1011 : 4'b0110;
											assign node253 = (inp[8]) ? node263 : node254;
												assign node254 = (inp[14]) ? node258 : node255;
													assign node255 = (inp[2]) ? 4'b1011 : 4'b0110;
													assign node258 = (inp[1]) ? 4'b1011 : node259;
														assign node259 = (inp[13]) ? 4'b1011 : 4'b0111;
												assign node263 = (inp[14]) ? node265 : 4'b1011;
													assign node265 = (inp[1]) ? 4'b1010 : node266;
														assign node266 = (inp[13]) ? 4'b1010 : 4'b0110;
									assign node270 = (inp[6]) ? node322 : node271;
										assign node271 = (inp[13]) ? node297 : node272;
											assign node272 = (inp[1]) ? node286 : node273;
												assign node273 = (inp[7]) ? node279 : node274;
													assign node274 = (inp[8]) ? node276 : 4'b0110;
														assign node276 = (inp[2]) ? 4'b0111 : 4'b0110;
													assign node279 = (inp[8]) ? node283 : node280;
														assign node280 = (inp[14]) ? 4'b0111 : 4'b0110;
														assign node283 = (inp[14]) ? 4'b0110 : 4'b0110;
												assign node286 = (inp[7]) ? node290 : node287;
													assign node287 = (inp[3]) ? 4'b0111 : 4'b0110;
													assign node290 = (inp[8]) ? node294 : node291;
														assign node291 = (inp[3]) ? 4'b0110 : 4'b1011;
														assign node294 = (inp[2]) ? 4'b1010 : 4'b1010;
											assign node297 = (inp[14]) ? node309 : node298;
												assign node298 = (inp[1]) ? node304 : node299;
													assign node299 = (inp[2]) ? node301 : 4'b0110;
														assign node301 = (inp[7]) ? 4'b1010 : 4'b0110;
													assign node304 = (inp[8]) ? node306 : 4'b1010;
														assign node306 = (inp[7]) ? 4'b1011 : 4'b1010;
												assign node309 = (inp[3]) ? node317 : node310;
													assign node310 = (inp[7]) ? node314 : node311;
														assign node311 = (inp[8]) ? 4'b1011 : 4'b1010;
														assign node314 = (inp[8]) ? 4'b1010 : 4'b1011;
													assign node317 = (inp[8]) ? 4'b1011 : node318;
														assign node318 = (inp[7]) ? 4'b1011 : 4'b1010;
										assign node322 = (inp[1]) ? node342 : node323;
											assign node323 = (inp[8]) ? node335 : node324;
												assign node324 = (inp[7]) ? node328 : node325;
													assign node325 = (inp[2]) ? 4'b1010 : 4'b1011;
													assign node328 = (inp[14]) ? node332 : node329;
														assign node329 = (inp[2]) ? 4'b1011 : 4'b1010;
														assign node332 = (inp[13]) ? 4'b0011 : 4'b1011;
												assign node335 = (inp[13]) ? node339 : node336;
													assign node336 = (inp[7]) ? 4'b1010 : 4'b1011;
													assign node339 = (inp[7]) ? 4'b0010 : 4'b0011;
											assign node342 = (inp[7]) ? node350 : node343;
												assign node343 = (inp[13]) ? node345 : 4'b1010;
													assign node345 = (inp[8]) ? node347 : 4'b0010;
														assign node347 = (inp[2]) ? 4'b0011 : 4'b0010;
												assign node350 = (inp[14]) ? 4'b0011 : node351;
													assign node351 = (inp[8]) ? 4'b0011 : node352;
														assign node352 = (inp[2]) ? 4'b0011 : 4'b0010;
							assign node357 = (inp[10]) ? node507 : node358;
								assign node358 = (inp[11]) ? node444 : node359;
									assign node359 = (inp[6]) ? node397 : node360;
										assign node360 = (inp[8]) ? node378 : node361;
											assign node361 = (inp[7]) ? node371 : node362;
												assign node362 = (inp[14]) ? node366 : node363;
													assign node363 = (inp[2]) ? 4'b1110 : 4'b1111;
													assign node366 = (inp[1]) ? node368 : 4'b1110;
														assign node368 = (inp[13]) ? 4'b0110 : 4'b1110;
												assign node371 = (inp[13]) ? node375 : node372;
													assign node372 = (inp[1]) ? 4'b1110 : 4'b1111;
													assign node375 = (inp[2]) ? 4'b0111 : 4'b0110;
											assign node378 = (inp[13]) ? node390 : node379;
												assign node379 = (inp[1]) ? node385 : node380;
													assign node380 = (inp[7]) ? node382 : 4'b1111;
														assign node382 = (inp[3]) ? 4'b1110 : 4'b1111;
													assign node385 = (inp[7]) ? node387 : 4'b0111;
														assign node387 = (inp[2]) ? 4'b0110 : 4'b0111;
												assign node390 = (inp[7]) ? node394 : node391;
													assign node391 = (inp[2]) ? 4'b0111 : 4'b0110;
													assign node394 = (inp[2]) ? 4'b0110 : 4'b0111;
										assign node397 = (inp[13]) ? node423 : node398;
											assign node398 = (inp[1]) ? node410 : node399;
												assign node399 = (inp[8]) ? node405 : node400;
													assign node400 = (inp[7]) ? 4'b0111 : node401;
														assign node401 = (inp[3]) ? 4'b0110 : 4'b0110;
													assign node405 = (inp[14]) ? 4'b0110 : node406;
														assign node406 = (inp[2]) ? 4'b0110 : 4'b0110;
												assign node410 = (inp[7]) ? node418 : node411;
													assign node411 = (inp[2]) ? node415 : node412;
														assign node412 = (inp[8]) ? 4'b0110 : 4'b0110;
														assign node415 = (inp[8]) ? 4'b1011 : 4'b0110;
													assign node418 = (inp[3]) ? 4'b1010 : node419;
														assign node419 = (inp[2]) ? 4'b1010 : 4'b1011;
											assign node423 = (inp[8]) ? node433 : node424;
												assign node424 = (inp[7]) ? 4'b1011 : node425;
													assign node425 = (inp[1]) ? node429 : node426;
														assign node426 = (inp[14]) ? 4'b0110 : 4'b0111;
														assign node429 = (inp[2]) ? 4'b1010 : 4'b1011;
												assign node433 = (inp[7]) ? node439 : node434;
													assign node434 = (inp[14]) ? 4'b1011 : node435;
														assign node435 = (inp[2]) ? 4'b1011 : 4'b1010;
													assign node439 = (inp[14]) ? 4'b1010 : node440;
														assign node440 = (inp[2]) ? 4'b1010 : 4'b1011;
									assign node444 = (inp[6]) ? node476 : node445;
										assign node445 = (inp[1]) ? node463 : node446;
											assign node446 = (inp[13]) ? node454 : node447;
												assign node447 = (inp[2]) ? 4'b0110 : node448;
													assign node448 = (inp[14]) ? node450 : 4'b0111;
														assign node450 = (inp[8]) ? 4'b0110 : 4'b0111;
												assign node454 = (inp[14]) ? 4'b1011 : node455;
													assign node455 = (inp[2]) ? node459 : node456;
														assign node456 = (inp[3]) ? 4'b0110 : 4'b1011;
														assign node459 = (inp[8]) ? 4'b1010 : 4'b1011;
											assign node463 = (inp[2]) ? node471 : node464;
												assign node464 = (inp[13]) ? 4'b1011 : node465;
													assign node465 = (inp[14]) ? 4'b1011 : node466;
														assign node466 = (inp[8]) ? 4'b0010 : 4'b0110;
												assign node471 = (inp[7]) ? node473 : 4'b1011;
													assign node473 = (inp[8]) ? 4'b1010 : 4'b1011;
										assign node476 = (inp[13]) ? node494 : node477;
											assign node477 = (inp[1]) ? node489 : node478;
												assign node478 = (inp[3]) ? node484 : node479;
													assign node479 = (inp[2]) ? node481 : 4'b1010;
														assign node481 = (inp[8]) ? 4'b1010 : 4'b1010;
													assign node484 = (inp[2]) ? 4'b1011 : node485;
														assign node485 = (inp[7]) ? 4'b1010 : 4'b1011;
												assign node489 = (inp[2]) ? 4'b0011 : node490;
													assign node490 = (inp[7]) ? 4'b0011 : 4'b1010;
											assign node494 = (inp[7]) ? node498 : node495;
												assign node495 = (inp[8]) ? 4'b0011 : 4'b0010;
												assign node498 = (inp[8]) ? node504 : node499;
													assign node499 = (inp[14]) ? 4'b0011 : node500;
														assign node500 = (inp[2]) ? 4'b0011 : 4'b0010;
													assign node504 = (inp[2]) ? 4'b0010 : 4'b0011;
								assign node507 = (inp[13]) ? node583 : node508;
									assign node508 = (inp[6]) ? node550 : node509;
										assign node509 = (inp[11]) ? node533 : node510;
											assign node510 = (inp[1]) ? node522 : node511;
												assign node511 = (inp[2]) ? node517 : node512;
													assign node512 = (inp[3]) ? 4'b1010 : node513;
														assign node513 = (inp[8]) ? 4'b1010 : 4'b1010;
													assign node517 = (inp[14]) ? node519 : 4'b1011;
														assign node519 = (inp[8]) ? 4'b1010 : 4'b1010;
												assign node522 = (inp[7]) ? node530 : node523;
													assign node523 = (inp[8]) ? node527 : node524;
														assign node524 = (inp[14]) ? 4'b1010 : 4'b1011;
														assign node527 = (inp[14]) ? 4'b0011 : 4'b1010;
													assign node530 = (inp[2]) ? 4'b0010 : 4'b0011;
											assign node533 = (inp[7]) ? node545 : node534;
												assign node534 = (inp[8]) ? node540 : node535;
													assign node535 = (inp[2]) ? 4'b0010 : node536;
														assign node536 = (inp[14]) ? 4'b0010 : 4'b0011;
													assign node540 = (inp[14]) ? 4'b1011 : node541;
														assign node541 = (inp[2]) ? 4'b0011 : 4'b0010;
												assign node545 = (inp[1]) ? node547 : 4'b0011;
													assign node547 = (inp[8]) ? 4'b1010 : 4'b1011;
										assign node550 = (inp[8]) ? node564 : node551;
											assign node551 = (inp[11]) ? node561 : node552;
												assign node552 = (inp[14]) ? 4'b0010 : node553;
													assign node553 = (inp[2]) ? node557 : node554;
														assign node554 = (inp[7]) ? 4'b0010 : 4'b0011;
														assign node557 = (inp[7]) ? 4'b1011 : 4'b0010;
												assign node561 = (inp[7]) ? 4'b0011 : 4'b1010;
											assign node564 = (inp[14]) ? node574 : node565;
												assign node565 = (inp[11]) ? node571 : node566;
													assign node566 = (inp[7]) ? 4'b1011 : node567;
														assign node567 = (inp[2]) ? 4'b0011 : 4'b0010;
													assign node571 = (inp[1]) ? 4'b0011 : 4'b1011;
												assign node574 = (inp[7]) ? node578 : node575;
													assign node575 = (inp[1]) ? 4'b1011 : 4'b0011;
													assign node578 = (inp[3]) ? node580 : 4'b0010;
														assign node580 = (inp[11]) ? 4'b0010 : 4'b1010;
									assign node583 = (inp[1]) ? node639 : node584;
										assign node584 = (inp[14]) ? node612 : node585;
											assign node585 = (inp[3]) ? node597 : node586;
												assign node586 = (inp[8]) ? node590 : node587;
													assign node587 = (inp[2]) ? 4'b1011 : 4'b1010;
													assign node590 = (inp[11]) ? node594 : node591;
														assign node591 = (inp[6]) ? 4'b0010 : 4'b0010;
														assign node594 = (inp[2]) ? 4'b1011 : 4'b0010;
												assign node597 = (inp[2]) ? node605 : node598;
													assign node598 = (inp[11]) ? node602 : node599;
														assign node599 = (inp[6]) ? 4'b0010 : 4'b1011;
														assign node602 = (inp[6]) ? 4'b0010 : 4'b0010;
													assign node605 = (inp[7]) ? node609 : node606;
														assign node606 = (inp[8]) ? 4'b1011 : 4'b0010;
														assign node609 = (inp[8]) ? 4'b0010 : 4'b0011;
											assign node612 = (inp[6]) ? node626 : node613;
												assign node613 = (inp[11]) ? node621 : node614;
													assign node614 = (inp[3]) ? node618 : node615;
														assign node615 = (inp[8]) ? 4'b0010 : 4'b0011;
														assign node618 = (inp[8]) ? 4'b0011 : 4'b1010;
													assign node621 = (inp[8]) ? 4'b1011 : node622;
														assign node622 = (inp[7]) ? 4'b1011 : 4'b0010;
												assign node626 = (inp[11]) ? node632 : node627;
													assign node627 = (inp[8]) ? 4'b1010 : node628;
														assign node628 = (inp[7]) ? 4'b1011 : 4'b0010;
													assign node632 = (inp[8]) ? node636 : node633;
														assign node633 = (inp[2]) ? 4'b1010 : 4'b0011;
														assign node636 = (inp[7]) ? 4'b0010 : 4'b0011;
										assign node639 = (inp[8]) ? node659 : node640;
											assign node640 = (inp[7]) ? node648 : node641;
												assign node641 = (inp[2]) ? 4'b1010 : node642;
													assign node642 = (inp[3]) ? node644 : 4'b1010;
														assign node644 = (inp[11]) ? 4'b0011 : 4'b0011;
												assign node648 = (inp[3]) ? node654 : node649;
													assign node649 = (inp[14]) ? node651 : 4'b0011;
														assign node651 = (inp[6]) ? 4'b1011 : 4'b0011;
													assign node654 = (inp[14]) ? 4'b1011 : node655;
														assign node655 = (inp[2]) ? 4'b1011 : 4'b1010;
											assign node659 = (inp[7]) ? node671 : node660;
												assign node660 = (inp[6]) ? node668 : node661;
													assign node661 = (inp[11]) ? node665 : node662;
														assign node662 = (inp[2]) ? 4'b0011 : 4'b0010;
														assign node665 = (inp[3]) ? 4'b1010 : 4'b1011;
													assign node668 = (inp[11]) ? 4'b0011 : 4'b1011;
												assign node671 = (inp[14]) ? node679 : node672;
													assign node672 = (inp[2]) ? node676 : node673;
														assign node673 = (inp[3]) ? 4'b0011 : 4'b1011;
														assign node676 = (inp[6]) ? 4'b0010 : 4'b1010;
													assign node679 = (inp[3]) ? node683 : node680;
														assign node680 = (inp[11]) ? 4'b0010 : 4'b0010;
														assign node683 = (inp[11]) ? 4'b1010 : 4'b0010;
						assign node686 = (inp[12]) ? node1022 : node687;
							assign node687 = (inp[10]) ? node861 : node688;
								assign node688 = (inp[6]) ? node770 : node689;
									assign node689 = (inp[7]) ? node727 : node690;
										assign node690 = (inp[8]) ? node710 : node691;
											assign node691 = (inp[11]) ? node701 : node692;
												assign node692 = (inp[13]) ? node698 : node693;
													assign node693 = (inp[2]) ? 4'b1010 : node694;
														assign node694 = (inp[14]) ? 4'b1010 : 4'b1011;
													assign node698 = (inp[1]) ? 4'b0010 : 4'b1010;
												assign node701 = (inp[13]) ? node707 : node702;
													assign node702 = (inp[14]) ? 4'b0010 : node703;
														assign node703 = (inp[2]) ? 4'b0010 : 4'b0011;
													assign node707 = (inp[14]) ? 4'b1010 : 4'b0011;
											assign node710 = (inp[14]) ? node718 : node711;
												assign node711 = (inp[2]) ? 4'b1011 : node712;
													assign node712 = (inp[11]) ? node714 : 4'b1010;
														assign node714 = (inp[13]) ? 4'b0010 : 4'b0010;
												assign node718 = (inp[11]) ? node722 : node719;
													assign node719 = (inp[1]) ? 4'b0011 : 4'b1011;
													assign node722 = (inp[13]) ? 4'b1011 : node723;
														assign node723 = (inp[3]) ? 4'b0011 : 4'b1011;
										assign node727 = (inp[8]) ? node751 : node728;
											assign node728 = (inp[2]) ? node742 : node729;
												assign node729 = (inp[14]) ? node737 : node730;
													assign node730 = (inp[13]) ? node734 : node731;
														assign node731 = (inp[11]) ? 4'b0010 : 4'b1010;
														assign node734 = (inp[11]) ? 4'b1010 : 4'b0010;
													assign node737 = (inp[3]) ? node739 : 4'b1011;
														assign node739 = (inp[13]) ? 4'b0011 : 4'b1011;
												assign node742 = (inp[11]) ? node748 : node743;
													assign node743 = (inp[13]) ? 4'b0011 : node744;
														assign node744 = (inp[14]) ? 4'b0011 : 4'b1011;
													assign node748 = (inp[13]) ? 4'b1011 : 4'b0011;
											assign node751 = (inp[2]) ? node761 : node752;
												assign node752 = (inp[14]) ? node758 : node753;
													assign node753 = (inp[3]) ? 4'b1011 : node754;
														assign node754 = (inp[1]) ? 4'b0011 : 4'b0011;
													assign node758 = (inp[1]) ? 4'b0010 : 4'b1010;
												assign node761 = (inp[11]) ? node767 : node762;
													assign node762 = (inp[13]) ? 4'b0010 : node763;
														assign node763 = (inp[1]) ? 4'b0010 : 4'b1010;
													assign node767 = (inp[13]) ? 4'b1010 : 4'b0010;
									assign node770 = (inp[3]) ? node812 : node771;
										assign node771 = (inp[7]) ? node785 : node772;
											assign node772 = (inp[8]) ? node782 : node773;
												assign node773 = (inp[2]) ? node777 : node774;
													assign node774 = (inp[14]) ? 4'b0010 : 4'b0011;
													assign node777 = (inp[13]) ? node779 : 4'b1010;
														assign node779 = (inp[11]) ? 4'b0010 : 4'b0010;
												assign node782 = (inp[2]) ? 4'b0011 : 4'b0010;
											assign node785 = (inp[8]) ? node797 : node786;
												assign node786 = (inp[2]) ? node792 : node787;
													assign node787 = (inp[14]) ? 4'b1011 : node788;
														assign node788 = (inp[1]) ? 4'b1010 : 4'b0010;
													assign node792 = (inp[13]) ? 4'b0011 : node793;
														assign node793 = (inp[11]) ? 4'b0011 : 4'b1011;
												assign node797 = (inp[11]) ? node805 : node798;
													assign node798 = (inp[13]) ? node802 : node799;
														assign node799 = (inp[1]) ? 4'b1010 : 4'b0010;
														assign node802 = (inp[2]) ? 4'b1010 : 4'b1011;
													assign node805 = (inp[1]) ? node809 : node806;
														assign node806 = (inp[13]) ? 4'b0010 : 4'b1010;
														assign node809 = (inp[2]) ? 4'b0010 : 4'b0010;
										assign node812 = (inp[2]) ? node838 : node813;
											assign node813 = (inp[14]) ? node827 : node814;
												assign node814 = (inp[8]) ? node822 : node815;
													assign node815 = (inp[7]) ? node819 : node816;
														assign node816 = (inp[13]) ? 4'b0011 : 4'b0011;
														assign node819 = (inp[1]) ? 4'b1010 : 4'b0010;
													assign node822 = (inp[7]) ? node824 : 4'b1010;
														assign node824 = (inp[13]) ? 4'b1011 : 4'b0011;
												assign node827 = (inp[1]) ? node833 : node828;
													assign node828 = (inp[11]) ? 4'b0010 : node829;
														assign node829 = (inp[13]) ? 4'b1011 : 4'b0010;
													assign node833 = (inp[11]) ? node835 : 4'b1010;
														assign node835 = (inp[13]) ? 4'b0011 : 4'b0010;
											assign node838 = (inp[7]) ? node850 : node839;
												assign node839 = (inp[8]) ? node847 : node840;
													assign node840 = (inp[11]) ? node844 : node841;
														assign node841 = (inp[1]) ? 4'b1010 : 4'b0010;
														assign node844 = (inp[13]) ? 4'b0010 : 4'b1010;
													assign node847 = (inp[1]) ? 4'b1011 : 4'b0011;
												assign node850 = (inp[8]) ? node856 : node851;
													assign node851 = (inp[14]) ? node853 : 4'b0011;
														assign node853 = (inp[13]) ? 4'b0011 : 4'b1011;
													assign node856 = (inp[1]) ? node858 : 4'b1010;
														assign node858 = (inp[11]) ? 4'b0010 : 4'b1010;
								assign node861 = (inp[11]) ? node949 : node862;
									assign node862 = (inp[6]) ? node906 : node863;
										assign node863 = (inp[1]) ? node883 : node864;
											assign node864 = (inp[8]) ? node872 : node865;
												assign node865 = (inp[7]) ? node867 : 4'b1010;
													assign node867 = (inp[3]) ? node869 : 4'b0011;
														assign node869 = (inp[2]) ? 4'b1011 : 4'b1010;
												assign node872 = (inp[13]) ? node878 : node873;
													assign node873 = (inp[2]) ? node875 : 4'b1010;
														assign node875 = (inp[7]) ? 4'b1010 : 4'b1011;
													assign node878 = (inp[3]) ? node880 : 4'b0011;
														assign node880 = (inp[7]) ? 4'b0010 : 4'b1010;
											assign node883 = (inp[8]) ? node897 : node884;
												assign node884 = (inp[13]) ? node892 : node885;
													assign node885 = (inp[2]) ? node889 : node886;
														assign node886 = (inp[7]) ? 4'b1010 : 4'b1010;
														assign node889 = (inp[14]) ? 4'b1010 : 4'b0011;
													assign node892 = (inp[7]) ? node894 : 4'b0010;
														assign node894 = (inp[2]) ? 4'b0011 : 4'b0010;
												assign node897 = (inp[2]) ? node903 : node898;
													assign node898 = (inp[14]) ? 4'b0011 : node899;
														assign node899 = (inp[7]) ? 4'b0011 : 4'b0010;
													assign node903 = (inp[7]) ? 4'b0010 : 4'b0011;
										assign node906 = (inp[13]) ? node934 : node907;
											assign node907 = (inp[1]) ? node921 : node908;
												assign node908 = (inp[14]) ? node916 : node909;
													assign node909 = (inp[7]) ? node913 : node910;
														assign node910 = (inp[2]) ? 4'b0010 : 4'b0010;
														assign node913 = (inp[8]) ? 4'b0010 : 4'b0011;
													assign node916 = (inp[8]) ? node918 : 4'b0010;
														assign node918 = (inp[7]) ? 4'b0010 : 4'b0011;
												assign node921 = (inp[7]) ? node927 : node922;
													assign node922 = (inp[8]) ? 4'b1111 : node923;
														assign node923 = (inp[2]) ? 4'b0010 : 4'b0010;
													assign node927 = (inp[3]) ? node931 : node928;
														assign node928 = (inp[14]) ? 4'b1110 : 4'b0010;
														assign node931 = (inp[8]) ? 4'b1100 : 4'b1101;
											assign node934 = (inp[3]) ? node942 : node935;
												assign node935 = (inp[8]) ? 4'b1111 : node936;
													assign node936 = (inp[7]) ? 4'b1111 : node937;
														assign node937 = (inp[2]) ? 4'b0010 : 4'b1110;
												assign node942 = (inp[8]) ? node944 : 4'b1101;
													assign node944 = (inp[2]) ? 4'b1100 : node945;
														assign node945 = (inp[7]) ? 4'b1101 : 4'b1100;
									assign node949 = (inp[3]) ? node983 : node950;
										assign node950 = (inp[6]) ? node968 : node951;
											assign node951 = (inp[13]) ? node961 : node952;
												assign node952 = (inp[7]) ? node958 : node953;
													assign node953 = (inp[1]) ? 4'b0010 : node954;
														assign node954 = (inp[8]) ? 4'b0011 : 4'b0010;
													assign node958 = (inp[1]) ? 4'b1111 : 4'b0010;
												assign node961 = (inp[7]) ? node963 : 4'b1111;
													assign node963 = (inp[8]) ? 4'b1110 : node964;
														assign node964 = (inp[2]) ? 4'b1111 : 4'b1110;
											assign node968 = (inp[13]) ? node978 : node969;
												assign node969 = (inp[7]) ? node975 : node970;
													assign node970 = (inp[1]) ? 4'b1110 : node971;
														assign node971 = (inp[2]) ? 4'b1111 : 4'b1110;
													assign node975 = (inp[1]) ? 4'b0111 : 4'b1111;
												assign node978 = (inp[7]) ? node980 : 4'b0111;
													assign node980 = (inp[8]) ? 4'b0110 : 4'b0111;
										assign node983 = (inp[6]) ? node1003 : node984;
											assign node984 = (inp[13]) ? node996 : node985;
												assign node985 = (inp[1]) ? node991 : node986;
													assign node986 = (inp[14]) ? node988 : 4'b0010;
														assign node988 = (inp[2]) ? 4'b0011 : 4'b0010;
													assign node991 = (inp[7]) ? node993 : 4'b0010;
														assign node993 = (inp[2]) ? 4'b1101 : 4'b0000;
												assign node996 = (inp[1]) ? node998 : 4'b1101;
													assign node998 = (inp[2]) ? 4'b1100 : node999;
														assign node999 = (inp[14]) ? 4'b1100 : 4'b1101;
											assign node1003 = (inp[13]) ? node1015 : node1004;
												assign node1004 = (inp[7]) ? node1010 : node1005;
													assign node1005 = (inp[1]) ? node1007 : 4'b1101;
														assign node1007 = (inp[2]) ? 4'b1100 : 4'b1101;
													assign node1010 = (inp[14]) ? node1012 : 4'b1100;
														assign node1012 = (inp[2]) ? 4'b1100 : 4'b0100;
												assign node1015 = (inp[2]) ? 4'b0101 : node1016;
													assign node1016 = (inp[8]) ? 4'b0100 : node1017;
														assign node1017 = (inp[14]) ? 4'b0100 : 4'b0101;
							assign node1022 = (inp[3]) ? node1214 : node1023;
								assign node1023 = (inp[10]) ? node1119 : node1024;
									assign node1024 = (inp[6]) ? node1074 : node1025;
										assign node1025 = (inp[1]) ? node1051 : node1026;
											assign node1026 = (inp[11]) ? node1038 : node1027;
												assign node1027 = (inp[8]) ? node1033 : node1028;
													assign node1028 = (inp[13]) ? node1030 : 4'b1010;
														assign node1030 = (inp[2]) ? 4'b1010 : 4'b1011;
													assign node1033 = (inp[13]) ? node1035 : 4'b1011;
														assign node1035 = (inp[7]) ? 4'b0010 : 4'b0011;
												assign node1038 = (inp[7]) ? node1044 : node1039;
													assign node1039 = (inp[13]) ? node1041 : 4'b0010;
														assign node1041 = (inp[2]) ? 4'b0010 : 4'b0010;
													assign node1044 = (inp[13]) ? node1048 : node1045;
														assign node1045 = (inp[8]) ? 4'b0010 : 4'b0011;
														assign node1048 = (inp[2]) ? 4'b1111 : 4'b0010;
											assign node1051 = (inp[11]) ? node1063 : node1052;
												assign node1052 = (inp[13]) ? node1058 : node1053;
													assign node1053 = (inp[7]) ? 4'b0010 : node1054;
														assign node1054 = (inp[8]) ? 4'b1010 : 4'b1010;
													assign node1058 = (inp[2]) ? node1060 : 4'b0011;
														assign node1060 = (inp[7]) ? 4'b0011 : 4'b0010;
												assign node1063 = (inp[2]) ? node1069 : node1064;
													assign node1064 = (inp[7]) ? 4'b1111 : node1065;
														assign node1065 = (inp[13]) ? 4'b1111 : 4'b0010;
													assign node1069 = (inp[13]) ? 4'b1110 : node1070;
														assign node1070 = (inp[14]) ? 4'b1111 : 4'b1110;
										assign node1074 = (inp[11]) ? node1096 : node1075;
											assign node1075 = (inp[7]) ? node1089 : node1076;
												assign node1076 = (inp[8]) ? node1084 : node1077;
													assign node1077 = (inp[13]) ? node1081 : node1078;
														assign node1078 = (inp[2]) ? 4'b0010 : 4'b0010;
														assign node1081 = (inp[1]) ? 4'b1110 : 4'b0010;
													assign node1084 = (inp[2]) ? 4'b1111 : node1085;
														assign node1085 = (inp[14]) ? 4'b1111 : 4'b0010;
												assign node1089 = (inp[8]) ? 4'b1110 : node1090;
													assign node1090 = (inp[13]) ? 4'b1111 : node1091;
														assign node1091 = (inp[1]) ? 4'b1111 : 4'b0011;
											assign node1096 = (inp[1]) ? node1106 : node1097;
												assign node1097 = (inp[7]) ? node1103 : node1098;
													assign node1098 = (inp[8]) ? node1100 : 4'b1110;
														assign node1100 = (inp[14]) ? 4'b1111 : 4'b1110;
													assign node1103 = (inp[13]) ? 4'b0110 : 4'b1110;
												assign node1106 = (inp[7]) ? node1114 : node1107;
													assign node1107 = (inp[13]) ? node1111 : node1108;
														assign node1108 = (inp[14]) ? 4'b1110 : 4'b1111;
														assign node1111 = (inp[14]) ? 4'b0110 : 4'b0111;
													assign node1114 = (inp[8]) ? node1116 : 4'b0111;
														assign node1116 = (inp[2]) ? 4'b0110 : 4'b0110;
									assign node1119 = (inp[2]) ? node1169 : node1120;
										assign node1120 = (inp[14]) ? node1144 : node1121;
											assign node1121 = (inp[1]) ? node1133 : node1122;
												assign node1122 = (inp[7]) ? node1128 : node1123;
													assign node1123 = (inp[8]) ? node1125 : 4'b0111;
														assign node1125 = (inp[13]) ? 4'b1110 : 4'b0110;
													assign node1128 = (inp[8]) ? 4'b1111 : node1129;
														assign node1129 = (inp[6]) ? 4'b1110 : 4'b0110;
												assign node1133 = (inp[6]) ? node1139 : node1134;
													assign node1134 = (inp[7]) ? node1136 : 4'b0110;
														assign node1136 = (inp[8]) ? 4'b0111 : 4'b0110;
													assign node1139 = (inp[11]) ? node1141 : 4'b1110;
														assign node1141 = (inp[13]) ? 4'b0110 : 4'b1111;
											assign node1144 = (inp[7]) ? node1156 : node1145;
												assign node1145 = (inp[8]) ? node1151 : node1146;
													assign node1146 = (inp[1]) ? node1148 : 4'b0110;
														assign node1148 = (inp[6]) ? 4'b1110 : 4'b0110;
													assign node1151 = (inp[13]) ? node1153 : 4'b0111;
														assign node1153 = (inp[6]) ? 4'b1111 : 4'b0111;
												assign node1156 = (inp[8]) ? node1164 : node1157;
													assign node1157 = (inp[11]) ? node1161 : node1158;
														assign node1158 = (inp[6]) ? 4'b1111 : 4'b0111;
														assign node1161 = (inp[6]) ? 4'b0111 : 4'b1111;
													assign node1164 = (inp[11]) ? node1166 : 4'b1110;
														assign node1166 = (inp[6]) ? 4'b0110 : 4'b1110;
										assign node1169 = (inp[6]) ? node1191 : node1170;
											assign node1170 = (inp[11]) ? node1182 : node1171;
												assign node1171 = (inp[1]) ? node1177 : node1172;
													assign node1172 = (inp[8]) ? node1174 : 4'b1110;
														assign node1174 = (inp[13]) ? 4'b0111 : 4'b1111;
													assign node1177 = (inp[13]) ? 4'b0111 : node1178;
														assign node1178 = (inp[7]) ? 4'b0110 : 4'b0111;
												assign node1182 = (inp[13]) ? node1186 : node1183;
													assign node1183 = (inp[1]) ? 4'b1111 : 4'b0111;
													assign node1186 = (inp[8]) ? node1188 : 4'b1111;
														assign node1188 = (inp[7]) ? 4'b1110 : 4'b1111;
											assign node1191 = (inp[11]) ? node1201 : node1192;
												assign node1192 = (inp[7]) ? node1198 : node1193;
													assign node1193 = (inp[8]) ? 4'b1111 : node1194;
														assign node1194 = (inp[14]) ? 4'b1110 : 4'b0110;
													assign node1198 = (inp[8]) ? 4'b1110 : 4'b1111;
												assign node1201 = (inp[13]) ? node1207 : node1202;
													assign node1202 = (inp[1]) ? node1204 : 4'b1110;
														assign node1204 = (inp[7]) ? 4'b0111 : 4'b1110;
													assign node1207 = (inp[1]) ? node1211 : node1208;
														assign node1208 = (inp[8]) ? 4'b0111 : 4'b1110;
														assign node1211 = (inp[14]) ? 4'b0110 : 4'b0110;
								assign node1214 = (inp[10]) ? node1306 : node1215;
									assign node1215 = (inp[11]) ? node1257 : node1216;
										assign node1216 = (inp[6]) ? node1240 : node1217;
											assign node1217 = (inp[13]) ? node1227 : node1218;
												assign node1218 = (inp[2]) ? node1222 : node1219;
													assign node1219 = (inp[7]) ? 4'b0011 : 4'b1011;
													assign node1222 = (inp[8]) ? node1224 : 4'b1010;
														assign node1224 = (inp[7]) ? 4'b1010 : 4'b1011;
												assign node1227 = (inp[14]) ? node1233 : node1228;
													assign node1228 = (inp[1]) ? 4'b0010 : node1229;
														assign node1229 = (inp[2]) ? 4'b0010 : 4'b0011;
													assign node1233 = (inp[7]) ? node1237 : node1234;
														assign node1234 = (inp[8]) ? 4'b0011 : 4'b1010;
														assign node1237 = (inp[8]) ? 4'b0010 : 4'b0011;
											assign node1240 = (inp[1]) ? node1252 : node1241;
												assign node1241 = (inp[13]) ? node1247 : node1242;
													assign node1242 = (inp[7]) ? node1244 : 4'b0010;
														assign node1244 = (inp[8]) ? 4'b0010 : 4'b0011;
													assign node1247 = (inp[8]) ? 4'b1101 : node1248;
														assign node1248 = (inp[2]) ? 4'b0000 : 4'b0010;
												assign node1252 = (inp[2]) ? node1254 : 4'b0010;
													assign node1254 = (inp[13]) ? 4'b1100 : 4'b1101;
										assign node1257 = (inp[6]) ? node1283 : node1258;
											assign node1258 = (inp[2]) ? node1272 : node1259;
												assign node1259 = (inp[14]) ? node1267 : node1260;
													assign node1260 = (inp[8]) ? node1264 : node1261;
														assign node1261 = (inp[7]) ? 4'b0010 : 4'b0011;
														assign node1264 = (inp[7]) ? 4'b0001 : 4'b0010;
													assign node1267 = (inp[13]) ? 4'b1101 : node1268;
														assign node1268 = (inp[8]) ? 4'b1100 : 4'b0010;
												assign node1272 = (inp[1]) ? node1278 : node1273;
													assign node1273 = (inp[8]) ? node1275 : 4'b0010;
														assign node1275 = (inp[7]) ? 4'b1100 : 4'b1101;
													assign node1278 = (inp[7]) ? node1280 : 4'b1101;
														assign node1280 = (inp[8]) ? 4'b1100 : 4'b1101;
											assign node1283 = (inp[13]) ? node1297 : node1284;
												assign node1284 = (inp[2]) ? node1292 : node1285;
													assign node1285 = (inp[7]) ? node1289 : node1286;
														assign node1286 = (inp[8]) ? 4'b0101 : 4'b1100;
														assign node1289 = (inp[1]) ? 4'b1100 : 4'b1101;
													assign node1292 = (inp[7]) ? node1294 : 4'b1100;
														assign node1294 = (inp[14]) ? 4'b0101 : 4'b0100;
												assign node1297 = (inp[8]) ? 4'b0101 : node1298;
													assign node1298 = (inp[1]) ? node1302 : node1299;
														assign node1299 = (inp[7]) ? 4'b0101 : 4'b1100;
														assign node1302 = (inp[2]) ? 4'b0100 : 4'b0101;
									assign node1306 = (inp[14]) ? node1350 : node1307;
										assign node1307 = (inp[13]) ? node1333 : node1308;
											assign node1308 = (inp[1]) ? node1320 : node1309;
												assign node1309 = (inp[11]) ? node1313 : node1310;
													assign node1310 = (inp[6]) ? 4'b0101 : 4'b1101;
													assign node1313 = (inp[6]) ? node1317 : node1314;
														assign node1314 = (inp[7]) ? 4'b0100 : 4'b0101;
														assign node1317 = (inp[2]) ? 4'b1100 : 4'b1100;
												assign node1320 = (inp[8]) ? node1326 : node1321;
													assign node1321 = (inp[6]) ? node1323 : 4'b0100;
														assign node1323 = (inp[11]) ? 4'b0101 : 4'b0100;
													assign node1326 = (inp[6]) ? node1330 : node1327;
														assign node1327 = (inp[2]) ? 4'b0100 : 4'b1100;
														assign node1330 = (inp[2]) ? 4'b1100 : 4'b1100;
											assign node1333 = (inp[8]) ? node1335 : 4'b1100;
												assign node1335 = (inp[7]) ? node1343 : node1336;
													assign node1336 = (inp[2]) ? node1340 : node1337;
														assign node1337 = (inp[1]) ? 4'b0100 : 4'b0100;
														assign node1340 = (inp[6]) ? 4'b1101 : 4'b0101;
													assign node1343 = (inp[2]) ? node1347 : node1344;
														assign node1344 = (inp[11]) ? 4'b0101 : 4'b1101;
														assign node1347 = (inp[1]) ? 4'b1100 : 4'b1100;
										assign node1350 = (inp[1]) ? node1370 : node1351;
											assign node1351 = (inp[8]) ? node1363 : node1352;
												assign node1352 = (inp[7]) ? node1358 : node1353;
													assign node1353 = (inp[6]) ? 4'b1100 : node1354;
														assign node1354 = (inp[11]) ? 4'b0100 : 4'b1100;
													assign node1358 = (inp[6]) ? 4'b1101 : node1359;
														assign node1359 = (inp[13]) ? 4'b1101 : 4'b0101;
												assign node1363 = (inp[7]) ? node1365 : 4'b0101;
													assign node1365 = (inp[11]) ? 4'b0100 : node1366;
														assign node1366 = (inp[13]) ? 4'b1100 : 4'b0100;
											assign node1370 = (inp[8]) ? node1380 : node1371;
												assign node1371 = (inp[7]) ? node1375 : node1372;
													assign node1372 = (inp[11]) ? 4'b0100 : 4'b1100;
													assign node1375 = (inp[13]) ? 4'b1101 : node1376;
														assign node1376 = (inp[11]) ? 4'b1101 : 4'b0101;
												assign node1380 = (inp[7]) ? node1386 : node1381;
													assign node1381 = (inp[6]) ? 4'b1101 : node1382;
														assign node1382 = (inp[13]) ? 4'b0101 : 4'b1101;
													assign node1386 = (inp[13]) ? 4'b1100 : node1387;
														assign node1387 = (inp[6]) ? 4'b1100 : 4'b1100;
					assign node1391 = (inp[3]) ? node2119 : node1392;
						assign node1392 = (inp[9]) ? node1754 : node1393;
							assign node1393 = (inp[12]) ? node1577 : node1394;
								assign node1394 = (inp[10]) ? node1486 : node1395;
									assign node1395 = (inp[13]) ? node1441 : node1396;
										assign node1396 = (inp[1]) ? node1420 : node1397;
											assign node1397 = (inp[7]) ? node1409 : node1398;
												assign node1398 = (inp[8]) ? node1404 : node1399;
													assign node1399 = (inp[2]) ? 4'b0110 : node1400;
														assign node1400 = (inp[11]) ? 4'b0111 : 4'b0111;
													assign node1404 = (inp[11]) ? node1406 : 4'b1111;
														assign node1406 = (inp[6]) ? 4'b1111 : 4'b0111;
												assign node1409 = (inp[14]) ? node1417 : node1410;
													assign node1410 = (inp[2]) ? node1414 : node1411;
														assign node1411 = (inp[8]) ? 4'b0111 : 4'b1110;
														assign node1414 = (inp[6]) ? 4'b1111 : 4'b0111;
													assign node1417 = (inp[8]) ? 4'b0110 : 4'b0111;
											assign node1420 = (inp[8]) ? node1428 : node1421;
												assign node1421 = (inp[7]) ? 4'b1111 : node1422;
													assign node1422 = (inp[6]) ? node1424 : 4'b0110;
														assign node1424 = (inp[11]) ? 4'b1110 : 4'b0110;
												assign node1428 = (inp[6]) ? node1434 : node1429;
													assign node1429 = (inp[11]) ? 4'b1110 : node1430;
														assign node1430 = (inp[2]) ? 4'b0111 : 4'b1110;
													assign node1434 = (inp[11]) ? node1438 : node1435;
														assign node1435 = (inp[14]) ? 4'b1111 : 4'b0110;
														assign node1438 = (inp[14]) ? 4'b0110 : 4'b0111;
										assign node1441 = (inp[6]) ? node1467 : node1442;
											assign node1442 = (inp[11]) ? node1454 : node1443;
												assign node1443 = (inp[2]) ? node1449 : node1444;
													assign node1444 = (inp[8]) ? 4'b0111 : node1445;
														assign node1445 = (inp[1]) ? 4'b0110 : 4'b1110;
													assign node1449 = (inp[8]) ? 4'b0110 : node1450;
														assign node1450 = (inp[7]) ? 4'b0111 : 4'b0110;
												assign node1454 = (inp[8]) ? node1462 : node1455;
													assign node1455 = (inp[1]) ? node1459 : node1456;
														assign node1456 = (inp[2]) ? 4'b1111 : 4'b0110;
														assign node1459 = (inp[14]) ? 4'b1110 : 4'b1110;
													assign node1462 = (inp[7]) ? node1464 : 4'b1111;
														assign node1464 = (inp[2]) ? 4'b1110 : 4'b1111;
											assign node1467 = (inp[11]) ? node1473 : node1468;
												assign node1468 = (inp[1]) ? node1470 : 4'b0110;
													assign node1470 = (inp[7]) ? 4'b1110 : 4'b1111;
												assign node1473 = (inp[1]) ? node1481 : node1474;
													assign node1474 = (inp[8]) ? node1478 : node1475;
														assign node1475 = (inp[2]) ? 4'b0110 : 4'b1110;
														assign node1478 = (inp[7]) ? 4'b0110 : 4'b0111;
													assign node1481 = (inp[7]) ? node1483 : 4'b0110;
														assign node1483 = (inp[8]) ? 4'b0110 : 4'b0111;
									assign node1486 = (inp[6]) ? node1530 : node1487;
										assign node1487 = (inp[11]) ? node1511 : node1488;
											assign node1488 = (inp[1]) ? node1498 : node1489;
												assign node1489 = (inp[13]) ? node1495 : node1490;
													assign node1490 = (inp[8]) ? node1492 : 4'b1110;
														assign node1492 = (inp[7]) ? 4'b1110 : 4'b1111;
													assign node1495 = (inp[8]) ? 4'b0110 : 4'b1110;
												assign node1498 = (inp[13]) ? node1506 : node1499;
													assign node1499 = (inp[8]) ? node1503 : node1500;
														assign node1500 = (inp[7]) ? 4'b0111 : 4'b1110;
														assign node1503 = (inp[7]) ? 4'b0110 : 4'b0111;
													assign node1506 = (inp[14]) ? node1508 : 4'b0110;
														assign node1508 = (inp[2]) ? 4'b0110 : 4'b0110;
											assign node1511 = (inp[13]) ? node1521 : node1512;
												assign node1512 = (inp[8]) ? node1514 : 4'b0110;
													assign node1514 = (inp[1]) ? node1518 : node1515;
														assign node1515 = (inp[2]) ? 4'b0110 : 4'b0111;
														assign node1518 = (inp[14]) ? 4'b1010 : 4'b0010;
												assign node1521 = (inp[7]) ? node1523 : 4'b1010;
													assign node1523 = (inp[8]) ? node1527 : node1524;
														assign node1524 = (inp[14]) ? 4'b1011 : 4'b1010;
														assign node1527 = (inp[14]) ? 4'b1010 : 4'b1011;
										assign node1530 = (inp[1]) ? node1554 : node1531;
											assign node1531 = (inp[11]) ? node1543 : node1532;
												assign node1532 = (inp[7]) ? node1538 : node1533;
													assign node1533 = (inp[2]) ? node1535 : 4'b0110;
														assign node1535 = (inp[8]) ? 4'b0111 : 4'b0110;
													assign node1538 = (inp[13]) ? 4'b1011 : node1539;
														assign node1539 = (inp[8]) ? 4'b0110 : 4'b0111;
												assign node1543 = (inp[13]) ? node1549 : node1544;
													assign node1544 = (inp[7]) ? node1546 : 4'b1010;
														assign node1546 = (inp[14]) ? 4'b1010 : 4'b1010;
													assign node1549 = (inp[14]) ? 4'b0011 : node1550;
														assign node1550 = (inp[8]) ? 4'b0010 : 4'b1010;
											assign node1554 = (inp[11]) ? node1566 : node1555;
												assign node1555 = (inp[14]) ? node1561 : node1556;
													assign node1556 = (inp[8]) ? 4'b1011 : node1557;
														assign node1557 = (inp[2]) ? 4'b1010 : 4'b1011;
													assign node1561 = (inp[2]) ? node1563 : 4'b1010;
														assign node1563 = (inp[13]) ? 4'b1010 : 4'b1010;
												assign node1566 = (inp[8]) ? node1572 : node1567;
													assign node1567 = (inp[14]) ? 4'b1010 : node1568;
														assign node1568 = (inp[2]) ? 4'b0011 : 4'b1011;
													assign node1572 = (inp[7]) ? node1574 : 4'b0011;
														assign node1574 = (inp[2]) ? 4'b0010 : 4'b0011;
								assign node1577 = (inp[10]) ? node1669 : node1578;
									assign node1578 = (inp[11]) ? node1622 : node1579;
										assign node1579 = (inp[6]) ? node1599 : node1580;
											assign node1580 = (inp[1]) ? node1592 : node1581;
												assign node1581 = (inp[2]) ? node1587 : node1582;
													assign node1582 = (inp[8]) ? node1584 : 4'b1111;
														assign node1584 = (inp[7]) ? 4'b1111 : 4'b1110;
													assign node1587 = (inp[13]) ? node1589 : 4'b1110;
														assign node1589 = (inp[7]) ? 4'b0110 : 4'b0111;
												assign node1592 = (inp[13]) ? node1594 : 4'b0111;
													assign node1594 = (inp[14]) ? node1596 : 4'b0111;
														assign node1596 = (inp[2]) ? 4'b0110 : 4'b0110;
											assign node1599 = (inp[1]) ? node1611 : node1600;
												assign node1600 = (inp[7]) ? node1606 : node1601;
													assign node1601 = (inp[2]) ? node1603 : 4'b0110;
														assign node1603 = (inp[8]) ? 4'b0111 : 4'b0110;
													assign node1606 = (inp[2]) ? 4'b1011 : node1607;
														assign node1607 = (inp[13]) ? 4'b0010 : 4'b0110;
												assign node1611 = (inp[13]) ? node1617 : node1612;
													assign node1612 = (inp[2]) ? node1614 : 4'b0110;
														assign node1614 = (inp[7]) ? 4'b1010 : 4'b1011;
													assign node1617 = (inp[7]) ? 4'b1011 : node1618;
														assign node1618 = (inp[8]) ? 4'b1011 : 4'b1010;
										assign node1622 = (inp[6]) ? node1646 : node1623;
											assign node1623 = (inp[1]) ? node1633 : node1624;
												assign node1624 = (inp[13]) ? node1628 : node1625;
													assign node1625 = (inp[7]) ? 4'b0110 : 4'b0111;
													assign node1628 = (inp[14]) ? node1630 : 4'b0110;
														assign node1630 = (inp[7]) ? 4'b1010 : 4'b1011;
												assign node1633 = (inp[13]) ? node1641 : node1634;
													assign node1634 = (inp[7]) ? node1638 : node1635;
														assign node1635 = (inp[2]) ? 4'b1011 : 4'b0110;
														assign node1638 = (inp[8]) ? 4'b1010 : 4'b1011;
													assign node1641 = (inp[2]) ? 4'b1010 : node1642;
														assign node1642 = (inp[7]) ? 4'b1010 : 4'b1010;
											assign node1646 = (inp[1]) ? node1660 : node1647;
												assign node1647 = (inp[13]) ? node1653 : node1648;
													assign node1648 = (inp[14]) ? node1650 : 4'b1011;
														assign node1650 = (inp[8]) ? 4'b1010 : 4'b1011;
													assign node1653 = (inp[2]) ? node1657 : node1654;
														assign node1654 = (inp[14]) ? 4'b0010 : 4'b1010;
														assign node1657 = (inp[7]) ? 4'b0010 : 4'b0011;
												assign node1660 = (inp[8]) ? node1664 : node1661;
													assign node1661 = (inp[7]) ? 4'b0011 : 4'b0010;
													assign node1664 = (inp[7]) ? 4'b0010 : node1665;
														assign node1665 = (inp[13]) ? 4'b0010 : 4'b1010;
									assign node1669 = (inp[7]) ? node1713 : node1670;
										assign node1670 = (inp[8]) ? node1688 : node1671;
											assign node1671 = (inp[14]) ? node1681 : node1672;
												assign node1672 = (inp[2]) ? node1678 : node1673;
													assign node1673 = (inp[1]) ? node1675 : 4'b0011;
														assign node1675 = (inp[6]) ? 4'b0011 : 4'b0011;
													assign node1678 = (inp[11]) ? 4'b1010 : 4'b0010;
												assign node1681 = (inp[1]) ? 4'b1010 : node1682;
													assign node1682 = (inp[11]) ? 4'b0010 : node1683;
														assign node1683 = (inp[13]) ? 4'b0010 : 4'b1010;
											assign node1688 = (inp[2]) ? node1700 : node1689;
												assign node1689 = (inp[14]) ? node1695 : node1690;
													assign node1690 = (inp[13]) ? node1692 : 4'b1010;
														assign node1692 = (inp[11]) ? 4'b1010 : 4'b0010;
													assign node1695 = (inp[11]) ? 4'b0011 : node1696;
														assign node1696 = (inp[1]) ? 4'b0011 : 4'b1011;
												assign node1700 = (inp[6]) ? node1708 : node1701;
													assign node1701 = (inp[11]) ? node1705 : node1702;
														assign node1702 = (inp[1]) ? 4'b0011 : 4'b1011;
														assign node1705 = (inp[13]) ? 4'b1011 : 4'b0011;
													assign node1708 = (inp[11]) ? 4'b0011 : node1709;
														assign node1709 = (inp[13]) ? 4'b1011 : 4'b0011;
										assign node1713 = (inp[8]) ? node1729 : node1714;
											assign node1714 = (inp[14]) ? node1722 : node1715;
												assign node1715 = (inp[2]) ? 4'b0011 : node1716;
													assign node1716 = (inp[1]) ? 4'b0010 : node1717;
														assign node1717 = (inp[13]) ? 4'b0010 : 4'b1010;
												assign node1722 = (inp[13]) ? 4'b1011 : node1723;
													assign node1723 = (inp[1]) ? 4'b1011 : node1724;
														assign node1724 = (inp[2]) ? 4'b0011 : 4'b0011;
											assign node1729 = (inp[14]) ? node1741 : node1730;
												assign node1730 = (inp[2]) ? node1734 : node1731;
													assign node1731 = (inp[6]) ? 4'b1011 : 4'b0011;
													assign node1734 = (inp[13]) ? node1738 : node1735;
														assign node1735 = (inp[11]) ? 4'b0010 : 4'b1010;
														assign node1738 = (inp[6]) ? 4'b0010 : 4'b0010;
												assign node1741 = (inp[6]) ? node1747 : node1742;
													assign node1742 = (inp[13]) ? node1744 : 4'b0010;
														assign node1744 = (inp[2]) ? 4'b0010 : 4'b1010;
													assign node1747 = (inp[11]) ? node1751 : node1748;
														assign node1748 = (inp[1]) ? 4'b1010 : 4'b0010;
														assign node1751 = (inp[13]) ? 4'b0010 : 4'b1010;
							assign node1754 = (inp[12]) ? node1926 : node1755;
								assign node1755 = (inp[10]) ? node1833 : node1756;
									assign node1756 = (inp[8]) ? node1798 : node1757;
										assign node1757 = (inp[7]) ? node1777 : node1758;
											assign node1758 = (inp[14]) ? node1768 : node1759;
												assign node1759 = (inp[2]) ? node1765 : node1760;
													assign node1760 = (inp[1]) ? 4'b0011 : node1761;
														assign node1761 = (inp[6]) ? 4'b0011 : 4'b1011;
													assign node1765 = (inp[13]) ? 4'b0010 : 4'b1010;
												assign node1768 = (inp[11]) ? node1774 : node1769;
													assign node1769 = (inp[6]) ? 4'b0010 : node1770;
														assign node1770 = (inp[13]) ? 4'b0010 : 4'b1010;
													assign node1774 = (inp[6]) ? 4'b1010 : 4'b0010;
											assign node1777 = (inp[2]) ? node1787 : node1778;
												assign node1778 = (inp[14]) ? node1784 : node1779;
													assign node1779 = (inp[6]) ? node1781 : 4'b0010;
														assign node1781 = (inp[11]) ? 4'b1010 : 4'b0010;
													assign node1784 = (inp[13]) ? 4'b0011 : 4'b1011;
												assign node1787 = (inp[13]) ? node1793 : node1788;
													assign node1788 = (inp[11]) ? 4'b0011 : node1789;
														assign node1789 = (inp[1]) ? 4'b0011 : 4'b0011;
													assign node1793 = (inp[14]) ? node1795 : 4'b1011;
														assign node1795 = (inp[11]) ? 4'b1011 : 4'b0011;
										assign node1798 = (inp[7]) ? node1814 : node1799;
											assign node1799 = (inp[14]) ? node1807 : node1800;
												assign node1800 = (inp[2]) ? 4'b1011 : node1801;
													assign node1801 = (inp[1]) ? 4'b1010 : node1802;
														assign node1802 = (inp[13]) ? 4'b1010 : 4'b0010;
												assign node1807 = (inp[13]) ? 4'b1011 : node1808;
													assign node1808 = (inp[6]) ? 4'b0011 : node1809;
														assign node1809 = (inp[1]) ? 4'b0011 : 4'b1011;
											assign node1814 = (inp[14]) ? node1826 : node1815;
												assign node1815 = (inp[2]) ? node1821 : node1816;
													assign node1816 = (inp[1]) ? node1818 : 4'b1011;
														assign node1818 = (inp[6]) ? 4'b0011 : 4'b0011;
													assign node1821 = (inp[6]) ? 4'b0010 : node1822;
														assign node1822 = (inp[13]) ? 4'b0010 : 4'b1010;
												assign node1826 = (inp[6]) ? node1828 : 4'b0010;
													assign node1828 = (inp[11]) ? node1830 : 4'b1010;
														assign node1830 = (inp[13]) ? 4'b0010 : 4'b0010;
									assign node1833 = (inp[11]) ? node1879 : node1834;
										assign node1834 = (inp[6]) ? node1858 : node1835;
											assign node1835 = (inp[13]) ? node1847 : node1836;
												assign node1836 = (inp[1]) ? node1842 : node1837;
													assign node1837 = (inp[8]) ? node1839 : 4'b1010;
														assign node1839 = (inp[2]) ? 4'b1011 : 4'b1010;
													assign node1842 = (inp[2]) ? 4'b0011 : node1843;
														assign node1843 = (inp[8]) ? 4'b0010 : 4'b1010;
												assign node1847 = (inp[7]) ? node1853 : node1848;
													assign node1848 = (inp[1]) ? node1850 : 4'b1011;
														assign node1850 = (inp[8]) ? 4'b0011 : 4'b0010;
													assign node1853 = (inp[8]) ? node1855 : 4'b0011;
														assign node1855 = (inp[2]) ? 4'b0010 : 4'b0010;
											assign node1858 = (inp[1]) ? node1870 : node1859;
												assign node1859 = (inp[14]) ? node1865 : node1860;
													assign node1860 = (inp[7]) ? node1862 : 4'b0010;
														assign node1862 = (inp[13]) ? 4'b0010 : 4'b0011;
													assign node1865 = (inp[13]) ? 4'b1101 : node1866;
														assign node1866 = (inp[7]) ? 4'b0010 : 4'b0011;
												assign node1870 = (inp[8]) ? node1874 : node1871;
													assign node1871 = (inp[7]) ? 4'b1101 : 4'b0010;
													assign node1874 = (inp[7]) ? 4'b1100 : node1875;
														assign node1875 = (inp[13]) ? 4'b1100 : 4'b1101;
										assign node1879 = (inp[6]) ? node1901 : node1880;
											assign node1880 = (inp[13]) ? node1892 : node1881;
												assign node1881 = (inp[1]) ? node1887 : node1882;
													assign node1882 = (inp[7]) ? 4'b0011 : node1883;
														assign node1883 = (inp[8]) ? 4'b0010 : 4'b0010;
													assign node1887 = (inp[8]) ? node1889 : 4'b0010;
														assign node1889 = (inp[14]) ? 4'b1101 : 4'b0000;
												assign node1892 = (inp[14]) ? node1896 : node1893;
													assign node1893 = (inp[2]) ? 4'b1101 : 4'b0011;
													assign node1896 = (inp[7]) ? node1898 : 4'b1101;
														assign node1898 = (inp[8]) ? 4'b1100 : 4'b1101;
											assign node1901 = (inp[1]) ? node1915 : node1902;
												assign node1902 = (inp[13]) ? node1908 : node1903;
													assign node1903 = (inp[2]) ? node1905 : 4'b1100;
														assign node1905 = (inp[8]) ? 4'b1101 : 4'b1100;
													assign node1908 = (inp[8]) ? node1912 : node1909;
														assign node1909 = (inp[14]) ? 4'b1100 : 4'b0100;
														assign node1912 = (inp[14]) ? 4'b0101 : 4'b0100;
												assign node1915 = (inp[7]) ? node1921 : node1916;
													assign node1916 = (inp[13]) ? node1918 : 4'b1101;
														assign node1918 = (inp[2]) ? 4'b0100 : 4'b0100;
													assign node1921 = (inp[14]) ? node1923 : 4'b0101;
														assign node1923 = (inp[2]) ? 4'b0101 : 4'b0100;
								assign node1926 = (inp[10]) ? node2024 : node1927;
									assign node1927 = (inp[11]) ? node1967 : node1928;
										assign node1928 = (inp[6]) ? node1950 : node1929;
											assign node1929 = (inp[1]) ? node1937 : node1930;
												assign node1930 = (inp[13]) ? node1932 : 4'b1010;
													assign node1932 = (inp[8]) ? node1934 : 4'b1010;
														assign node1934 = (inp[14]) ? 4'b0010 : 4'b0011;
												assign node1937 = (inp[8]) ? node1945 : node1938;
													assign node1938 = (inp[7]) ? node1942 : node1939;
														assign node1939 = (inp[14]) ? 4'b0010 : 4'b1011;
														assign node1942 = (inp[2]) ? 4'b0011 : 4'b0010;
													assign node1945 = (inp[14]) ? node1947 : 4'b0010;
														assign node1947 = (inp[7]) ? 4'b0010 : 4'b0011;
											assign node1950 = (inp[1]) ? node1962 : node1951;
												assign node1951 = (inp[13]) ? node1957 : node1952;
													assign node1952 = (inp[7]) ? 4'b0011 : node1953;
														assign node1953 = (inp[8]) ? 4'b0011 : 4'b0010;
													assign node1957 = (inp[8]) ? node1959 : 4'b0010;
														assign node1959 = (inp[2]) ? 4'b1100 : 4'b0000;
												assign node1962 = (inp[7]) ? 4'b1101 : node1963;
													assign node1963 = (inp[8]) ? 4'b1101 : 4'b0010;
										assign node1967 = (inp[6]) ? node1995 : node1968;
											assign node1968 = (inp[1]) ? node1980 : node1969;
												assign node1969 = (inp[13]) ? node1977 : node1970;
													assign node1970 = (inp[14]) ? node1974 : node1971;
														assign node1971 = (inp[7]) ? 4'b0011 : 4'b0010;
														assign node1974 = (inp[7]) ? 4'b0010 : 4'b0010;
													assign node1977 = (inp[2]) ? 4'b1101 : 4'b0010;
												assign node1980 = (inp[13]) ? node1988 : node1981;
													assign node1981 = (inp[8]) ? node1985 : node1982;
														assign node1982 = (inp[2]) ? 4'b1101 : 4'b0010;
														assign node1985 = (inp[2]) ? 4'b1100 : 4'b1101;
													assign node1988 = (inp[14]) ? node1992 : node1989;
														assign node1989 = (inp[7]) ? 4'b1101 : 4'b1100;
														assign node1992 = (inp[7]) ? 4'b1101 : 4'b1101;
											assign node1995 = (inp[1]) ? node2009 : node1996;
												assign node1996 = (inp[13]) ? node2004 : node1997;
													assign node1997 = (inp[14]) ? node2001 : node1998;
														assign node1998 = (inp[7]) ? 4'b1101 : 4'b1100;
														assign node2001 = (inp[7]) ? 4'b1100 : 4'b1100;
													assign node2004 = (inp[7]) ? node2006 : 4'b1100;
														assign node2006 = (inp[14]) ? 4'b0101 : 4'b0100;
												assign node2009 = (inp[13]) ? node2017 : node2010;
													assign node2010 = (inp[8]) ? node2014 : node2011;
														assign node2011 = (inp[2]) ? 4'b0100 : 4'b1100;
														assign node2014 = (inp[7]) ? 4'b0100 : 4'b0101;
													assign node2017 = (inp[7]) ? node2021 : node2018;
														assign node2018 = (inp[8]) ? 4'b0101 : 4'b0100;
														assign node2021 = (inp[8]) ? 4'b0100 : 4'b0101;
									assign node2024 = (inp[2]) ? node2072 : node2025;
										assign node2025 = (inp[6]) ? node2051 : node2026;
											assign node2026 = (inp[14]) ? node2038 : node2027;
												assign node2027 = (inp[7]) ? node2031 : node2028;
													assign node2028 = (inp[8]) ? 4'b0100 : 4'b0101;
													assign node2031 = (inp[8]) ? node2035 : node2032;
														assign node2032 = (inp[11]) ? 4'b0100 : 4'b1100;
														assign node2035 = (inp[13]) ? 4'b0101 : 4'b0101;
												assign node2038 = (inp[1]) ? node2046 : node2039;
													assign node2039 = (inp[7]) ? node2043 : node2040;
														assign node2040 = (inp[8]) ? 4'b1101 : 4'b1100;
														assign node2043 = (inp[11]) ? 4'b0101 : 4'b0101;
													assign node2046 = (inp[13]) ? node2048 : 4'b0100;
														assign node2048 = (inp[7]) ? 4'b1100 : 4'b1100;
											assign node2051 = (inp[11]) ? node2059 : node2052;
												assign node2052 = (inp[13]) ? 4'b1100 : node2053;
													assign node2053 = (inp[7]) ? node2055 : 4'b0100;
														assign node2055 = (inp[1]) ? 4'b1101 : 4'b0100;
												assign node2059 = (inp[13]) ? node2065 : node2060;
													assign node2060 = (inp[8]) ? 4'b0101 : node2061;
														assign node2061 = (inp[14]) ? 4'b1100 : 4'b1100;
													assign node2065 = (inp[7]) ? node2069 : node2066;
														assign node2066 = (inp[8]) ? 4'b1100 : 4'b0101;
														assign node2069 = (inp[1]) ? 4'b0100 : 4'b0100;
										assign node2072 = (inp[7]) ? node2096 : node2073;
											assign node2073 = (inp[8]) ? node2083 : node2074;
												assign node2074 = (inp[11]) ? 4'b0100 : node2075;
													assign node2075 = (inp[6]) ? node2079 : node2076;
														assign node2076 = (inp[14]) ? 4'b0100 : 4'b1100;
														assign node2079 = (inp[1]) ? 4'b1100 : 4'b0100;
												assign node2083 = (inp[1]) ? node2091 : node2084;
													assign node2084 = (inp[6]) ? node2088 : node2085;
														assign node2085 = (inp[14]) ? 4'b0101 : 4'b1101;
														assign node2088 = (inp[14]) ? 4'b0101 : 4'b0101;
													assign node2091 = (inp[14]) ? node2093 : 4'b1101;
														assign node2093 = (inp[11]) ? 4'b0101 : 4'b1101;
											assign node2096 = (inp[8]) ? node2108 : node2097;
												assign node2097 = (inp[13]) ? node2103 : node2098;
													assign node2098 = (inp[1]) ? 4'b0101 : node2099;
														assign node2099 = (inp[6]) ? 4'b0101 : 4'b1101;
													assign node2103 = (inp[11]) ? node2105 : 4'b1101;
														assign node2105 = (inp[6]) ? 4'b0101 : 4'b1101;
												assign node2108 = (inp[1]) ? node2114 : node2109;
													assign node2109 = (inp[11]) ? 4'b1100 : node2110;
														assign node2110 = (inp[6]) ? 4'b0100 : 4'b1100;
													assign node2114 = (inp[14]) ? 4'b0100 : node2115;
														assign node2115 = (inp[13]) ? 4'b0100 : 4'b1100;
						assign node2119 = (inp[12]) ? node2485 : node2120;
							assign node2120 = (inp[9]) ? node2298 : node2121;
								assign node2121 = (inp[10]) ? node2213 : node2122;
									assign node2122 = (inp[13]) ? node2172 : node2123;
										assign node2123 = (inp[7]) ? node2145 : node2124;
											assign node2124 = (inp[8]) ? node2132 : node2125;
												assign node2125 = (inp[14]) ? 4'b0100 : node2126;
													assign node2126 = (inp[2]) ? 4'b1100 : node2127;
														assign node2127 = (inp[6]) ? 4'b0101 : 4'b0101;
												assign node2132 = (inp[11]) ? node2138 : node2133;
													assign node2133 = (inp[2]) ? 4'b1101 : node2134;
														assign node2134 = (inp[1]) ? 4'b0101 : 4'b1101;
													assign node2138 = (inp[14]) ? node2142 : node2139;
														assign node2139 = (inp[1]) ? 4'b0101 : 4'b0100;
														assign node2142 = (inp[1]) ? 4'b0101 : 4'b0101;
											assign node2145 = (inp[8]) ? node2157 : node2146;
												assign node2146 = (inp[2]) ? node2152 : node2147;
													assign node2147 = (inp[14]) ? 4'b1101 : node2148;
														assign node2148 = (inp[6]) ? 4'b0100 : 4'b1100;
													assign node2152 = (inp[1]) ? 4'b1101 : node2153;
														assign node2153 = (inp[11]) ? 4'b0101 : 4'b1101;
												assign node2157 = (inp[14]) ? node2165 : node2158;
													assign node2158 = (inp[2]) ? node2162 : node2159;
														assign node2159 = (inp[6]) ? 4'b0101 : 4'b0101;
														assign node2162 = (inp[11]) ? 4'b1100 : 4'b0100;
													assign node2165 = (inp[2]) ? node2169 : node2166;
														assign node2166 = (inp[11]) ? 4'b0100 : 4'b1100;
														assign node2169 = (inp[6]) ? 4'b0100 : 4'b0100;
										assign node2172 = (inp[11]) ? node2194 : node2173;
											assign node2173 = (inp[6]) ? node2185 : node2174;
												assign node2174 = (inp[2]) ? node2180 : node2175;
													assign node2175 = (inp[8]) ? node2177 : 4'b1100;
														assign node2177 = (inp[1]) ? 4'b0100 : 4'b0101;
													assign node2180 = (inp[7]) ? node2182 : 4'b0101;
														assign node2182 = (inp[8]) ? 4'b0100 : 4'b0101;
												assign node2185 = (inp[7]) ? node2191 : node2186;
													assign node2186 = (inp[1]) ? node2188 : 4'b0100;
														assign node2188 = (inp[8]) ? 4'b1100 : 4'b1100;
													assign node2191 = (inp[8]) ? 4'b1100 : 4'b1101;
											assign node2194 = (inp[6]) ? node2202 : node2195;
												assign node2195 = (inp[2]) ? 4'b1100 : node2196;
													assign node2196 = (inp[7]) ? 4'b1100 : node2197;
														assign node2197 = (inp[1]) ? 4'b1100 : 4'b0100;
												assign node2202 = (inp[7]) ? node2208 : node2203;
													assign node2203 = (inp[1]) ? node2205 : 4'b1100;
														assign node2205 = (inp[8]) ? 4'b0101 : 4'b0100;
													assign node2208 = (inp[8]) ? 4'b0100 : node2209;
														assign node2209 = (inp[1]) ? 4'b0100 : 4'b0101;
									assign node2213 = (inp[11]) ? node2253 : node2214;
										assign node2214 = (inp[6]) ? node2236 : node2215;
											assign node2215 = (inp[1]) ? node2229 : node2216;
												assign node2216 = (inp[13]) ? node2224 : node2217;
													assign node2217 = (inp[2]) ? node2221 : node2218;
														assign node2218 = (inp[14]) ? 4'b1100 : 4'b1100;
														assign node2221 = (inp[7]) ? 4'b1100 : 4'b1101;
													assign node2224 = (inp[14]) ? node2226 : 4'b1100;
														assign node2226 = (inp[8]) ? 4'b0100 : 4'b0101;
												assign node2229 = (inp[7]) ? node2231 : 4'b0101;
													assign node2231 = (inp[14]) ? 4'b0100 : node2232;
														assign node2232 = (inp[2]) ? 4'b0100 : 4'b0101;
											assign node2236 = (inp[1]) ? node2248 : node2237;
												assign node2237 = (inp[13]) ? node2243 : node2238;
													assign node2238 = (inp[2]) ? node2240 : 4'b0100;
														assign node2240 = (inp[14]) ? 4'b0101 : 4'b0100;
													assign node2243 = (inp[7]) ? node2245 : 4'b0101;
														assign node2245 = (inp[8]) ? 4'b1000 : 4'b1001;
												assign node2248 = (inp[14]) ? node2250 : 4'b1001;
													assign node2250 = (inp[13]) ? 4'b1000 : 4'b1001;
										assign node2253 = (inp[6]) ? node2273 : node2254;
											assign node2254 = (inp[1]) ? node2264 : node2255;
												assign node2255 = (inp[13]) ? node2259 : node2256;
													assign node2256 = (inp[8]) ? 4'b0100 : 4'b0101;
													assign node2259 = (inp[7]) ? node2261 : 4'b0100;
														assign node2261 = (inp[8]) ? 4'b1000 : 4'b0000;
												assign node2264 = (inp[7]) ? 4'b1000 : node2265;
													assign node2265 = (inp[8]) ? node2269 : node2266;
														assign node2266 = (inp[13]) ? 4'b1000 : 4'b0100;
														assign node2269 = (inp[14]) ? 4'b1001 : 4'b1000;
											assign node2273 = (inp[14]) ? node2285 : node2274;
												assign node2274 = (inp[13]) ? node2280 : node2275;
													assign node2275 = (inp[8]) ? node2277 : 4'b1000;
														assign node2277 = (inp[1]) ? 4'b1000 : 4'b1001;
													assign node2280 = (inp[7]) ? node2282 : 4'b1000;
														assign node2282 = (inp[8]) ? 4'b0001 : 4'b0000;
												assign node2285 = (inp[13]) ? node2293 : node2286;
													assign node2286 = (inp[1]) ? node2290 : node2287;
														assign node2287 = (inp[7]) ? 4'b1000 : 4'b1000;
														assign node2290 = (inp[7]) ? 4'b0000 : 4'b0001;
													assign node2293 = (inp[1]) ? 4'b0000 : node2294;
														assign node2294 = (inp[8]) ? 4'b0000 : 4'b0001;
								assign node2298 = (inp[10]) ? node2394 : node2299;
									assign node2299 = (inp[11]) ? node2345 : node2300;
										assign node2300 = (inp[2]) ? node2330 : node2301;
											assign node2301 = (inp[13]) ? node2315 : node2302;
												assign node2302 = (inp[6]) ? node2308 : node2303;
													assign node2303 = (inp[1]) ? 4'b0001 : node2304;
														assign node2304 = (inp[7]) ? 4'b1001 : 4'b1000;
													assign node2308 = (inp[1]) ? node2312 : node2309;
														assign node2309 = (inp[14]) ? 4'b0000 : 4'b0001;
														assign node2312 = (inp[14]) ? 4'b1000 : 4'b0000;
												assign node2315 = (inp[6]) ? node2323 : node2316;
													assign node2316 = (inp[1]) ? node2320 : node2317;
														assign node2317 = (inp[14]) ? 4'b0001 : 4'b1001;
														assign node2320 = (inp[8]) ? 4'b0000 : 4'b0000;
													assign node2323 = (inp[1]) ? node2327 : node2324;
														assign node2324 = (inp[14]) ? 4'b1000 : 4'b0000;
														assign node2327 = (inp[7]) ? 4'b1001 : 4'b1000;
											assign node2330 = (inp[8]) ? node2338 : node2331;
												assign node2331 = (inp[7]) ? 4'b1001 : node2332;
													assign node2332 = (inp[14]) ? 4'b1000 : node2333;
														assign node2333 = (inp[6]) ? 4'b0000 : 4'b1000;
												assign node2338 = (inp[7]) ? 4'b0000 : node2339;
													assign node2339 = (inp[13]) ? 4'b1001 : node2340;
														assign node2340 = (inp[6]) ? 4'b0001 : 4'b1001;
										assign node2345 = (inp[1]) ? node2373 : node2346;
											assign node2346 = (inp[6]) ? node2360 : node2347;
												assign node2347 = (inp[2]) ? node2355 : node2348;
													assign node2348 = (inp[13]) ? node2352 : node2349;
														assign node2349 = (inp[14]) ? 4'b0000 : 4'b0001;
														assign node2352 = (inp[8]) ? 4'b0000 : 4'b0000;
													assign node2355 = (inp[13]) ? node2357 : 4'b0001;
														assign node2357 = (inp[8]) ? 4'b1001 : 4'b0000;
												assign node2360 = (inp[13]) ? node2366 : node2361;
													assign node2361 = (inp[14]) ? node2363 : 4'b1001;
														assign node2363 = (inp[7]) ? 4'b1000 : 4'b1001;
													assign node2366 = (inp[14]) ? node2370 : node2367;
														assign node2367 = (inp[2]) ? 4'b1000 : 4'b1001;
														assign node2370 = (inp[2]) ? 4'b0001 : 4'b0001;
											assign node2373 = (inp[6]) ? node2387 : node2374;
												assign node2374 = (inp[14]) ? node2380 : node2375;
													assign node2375 = (inp[7]) ? 4'b1001 : node2376;
														assign node2376 = (inp[2]) ? 4'b1000 : 4'b0001;
													assign node2380 = (inp[8]) ? node2384 : node2381;
														assign node2381 = (inp[7]) ? 4'b1001 : 4'b1000;
														assign node2384 = (inp[7]) ? 4'b1000 : 4'b1001;
												assign node2387 = (inp[8]) ? node2391 : node2388;
													assign node2388 = (inp[14]) ? 4'b1000 : 4'b1001;
													assign node2391 = (inp[7]) ? 4'b0000 : 4'b0001;
									assign node2394 = (inp[11]) ? node2442 : node2395;
										assign node2395 = (inp[6]) ? node2417 : node2396;
											assign node2396 = (inp[13]) ? node2408 : node2397;
												assign node2397 = (inp[14]) ? node2403 : node2398;
													assign node2398 = (inp[1]) ? node2400 : 4'b1001;
														assign node2400 = (inp[2]) ? 4'b0000 : 4'b1000;
													assign node2403 = (inp[1]) ? node2405 : 4'b1000;
														assign node2405 = (inp[8]) ? 4'b0000 : 4'b1000;
												assign node2408 = (inp[1]) ? node2412 : node2409;
													assign node2409 = (inp[14]) ? 4'b0000 : 4'b1000;
													assign node2412 = (inp[7]) ? 4'b0001 : node2413;
														assign node2413 = (inp[8]) ? 4'b0001 : 4'b0000;
											assign node2417 = (inp[1]) ? node2431 : node2418;
												assign node2418 = (inp[13]) ? node2424 : node2419;
													assign node2419 = (inp[7]) ? node2421 : 4'b0000;
														assign node2421 = (inp[8]) ? 4'b0001 : 4'b0000;
													assign node2424 = (inp[8]) ? node2428 : node2425;
														assign node2425 = (inp[14]) ? 4'b0000 : 4'b0000;
														assign node2428 = (inp[7]) ? 4'b1100 : 4'b1101;
												assign node2431 = (inp[8]) ? node2437 : node2432;
													assign node2432 = (inp[7]) ? 4'b1101 : node2433;
														assign node2433 = (inp[14]) ? 4'b0000 : 4'b1101;
													assign node2437 = (inp[13]) ? 4'b1100 : node2438;
														assign node2438 = (inp[7]) ? 4'b1100 : 4'b1101;
										assign node2442 = (inp[6]) ? node2470 : node2443;
											assign node2443 = (inp[13]) ? node2455 : node2444;
												assign node2444 = (inp[1]) ? node2450 : node2445;
													assign node2445 = (inp[14]) ? 4'b0000 : node2446;
														assign node2446 = (inp[2]) ? 4'b0000 : 4'b0001;
													assign node2450 = (inp[7]) ? 4'b1101 : node2451;
														assign node2451 = (inp[8]) ? 4'b1101 : 4'b0000;
												assign node2455 = (inp[1]) ? node2463 : node2456;
													assign node2456 = (inp[7]) ? node2460 : node2457;
														assign node2457 = (inp[8]) ? 4'b1101 : 4'b0000;
														assign node2460 = (inp[8]) ? 4'b1100 : 4'b1101;
													assign node2463 = (inp[7]) ? node2467 : node2464;
														assign node2464 = (inp[14]) ? 4'b1101 : 4'b1100;
														assign node2467 = (inp[8]) ? 4'b1100 : 4'b1100;
											assign node2470 = (inp[1]) ? node2478 : node2471;
												assign node2471 = (inp[2]) ? node2473 : 4'b0101;
													assign node2473 = (inp[8]) ? node2475 : 4'b1100;
														assign node2475 = (inp[7]) ? 4'b0100 : 4'b0101;
												assign node2478 = (inp[7]) ? node2480 : 4'b0101;
													assign node2480 = (inp[14]) ? 4'b0101 : node2481;
														assign node2481 = (inp[8]) ? 4'b0100 : 4'b1100;
							assign node2485 = (inp[9]) ? node2653 : node2486;
								assign node2486 = (inp[10]) ? node2578 : node2487;
									assign node2487 = (inp[11]) ? node2539 : node2488;
										assign node2488 = (inp[6]) ? node2512 : node2489;
											assign node2489 = (inp[7]) ? node2501 : node2490;
												assign node2490 = (inp[8]) ? node2496 : node2491;
													assign node2491 = (inp[2]) ? node2493 : 4'b1101;
														assign node2493 = (inp[1]) ? 4'b0100 : 4'b1100;
													assign node2496 = (inp[14]) ? 4'b0101 : node2497;
														assign node2497 = (inp[2]) ? 4'b0101 : 4'b1100;
												assign node2501 = (inp[2]) ? node2509 : node2502;
													assign node2502 = (inp[1]) ? node2506 : node2503;
														assign node2503 = (inp[13]) ? 4'b0100 : 4'b1101;
														assign node2506 = (inp[8]) ? 4'b0101 : 4'b0100;
													assign node2509 = (inp[8]) ? 4'b0100 : 4'b0101;
											assign node2512 = (inp[1]) ? node2524 : node2513;
												assign node2513 = (inp[13]) ? node2519 : node2514;
													assign node2514 = (inp[2]) ? 4'b0101 : node2515;
														assign node2515 = (inp[7]) ? 4'b0100 : 4'b0101;
													assign node2519 = (inp[7]) ? 4'b1001 : node2520;
														assign node2520 = (inp[2]) ? 4'b0100 : 4'b0101;
												assign node2524 = (inp[13]) ? node2532 : node2525;
													assign node2525 = (inp[8]) ? node2529 : node2526;
														assign node2526 = (inp[14]) ? 4'b0100 : 4'b0100;
														assign node2529 = (inp[2]) ? 4'b1000 : 4'b1001;
													assign node2532 = (inp[2]) ? node2536 : node2533;
														assign node2533 = (inp[7]) ? 4'b1000 : 4'b1000;
														assign node2536 = (inp[8]) ? 4'b1000 : 4'b1001;
										assign node2539 = (inp[6]) ? node2559 : node2540;
											assign node2540 = (inp[7]) ? node2550 : node2541;
												assign node2541 = (inp[1]) ? node2547 : node2542;
													assign node2542 = (inp[13]) ? node2544 : 4'b0101;
														assign node2544 = (inp[2]) ? 4'b0100 : 4'b0100;
													assign node2547 = (inp[13]) ? 4'b1000 : 4'b0100;
												assign node2550 = (inp[2]) ? node2556 : node2551;
													assign node2551 = (inp[13]) ? node2553 : 4'b0101;
														assign node2553 = (inp[8]) ? 4'b1000 : 4'b0000;
													assign node2556 = (inp[8]) ? 4'b1000 : 4'b1001;
											assign node2559 = (inp[1]) ? node2571 : node2560;
												assign node2560 = (inp[14]) ? node2566 : node2561;
													assign node2561 = (inp[13]) ? node2563 : 4'b1000;
														assign node2563 = (inp[2]) ? 4'b0000 : 4'b1000;
													assign node2566 = (inp[13]) ? node2568 : 4'b1001;
														assign node2568 = (inp[2]) ? 4'b0000 : 4'b0001;
												assign node2571 = (inp[2]) ? 4'b0000 : node2572;
													assign node2572 = (inp[14]) ? 4'b0001 : node2573;
														assign node2573 = (inp[13]) ? 4'b0001 : 4'b1001;
									assign node2578 = (inp[7]) ? node2620 : node2579;
										assign node2579 = (inp[8]) ? node2599 : node2580;
											assign node2580 = (inp[2]) ? node2588 : node2581;
												assign node2581 = (inp[14]) ? 4'b1000 : node2582;
													assign node2582 = (inp[1]) ? 4'b1001 : node2583;
														assign node2583 = (inp[13]) ? 4'b1001 : 4'b0001;
												assign node2588 = (inp[14]) ? node2594 : node2589;
													assign node2589 = (inp[1]) ? node2591 : 4'b0000;
														assign node2591 = (inp[13]) ? 4'b0000 : 4'b1000;
													assign node2594 = (inp[13]) ? 4'b1000 : node2595;
														assign node2595 = (inp[11]) ? 4'b0000 : 4'b1000;
											assign node2599 = (inp[14]) ? node2609 : node2600;
												assign node2600 = (inp[2]) ? 4'b0001 : node2601;
													assign node2601 = (inp[6]) ? node2605 : node2602;
														assign node2602 = (inp[11]) ? 4'b0000 : 4'b1000;
														assign node2605 = (inp[11]) ? 4'b1000 : 4'b0000;
												assign node2609 = (inp[2]) ? node2615 : node2610;
													assign node2610 = (inp[13]) ? node2612 : 4'b1001;
														assign node2612 = (inp[11]) ? 4'b0001 : 4'b1001;
													assign node2615 = (inp[11]) ? 4'b0001 : node2616;
														assign node2616 = (inp[6]) ? 4'b0001 : 4'b0001;
										assign node2620 = (inp[8]) ? node2638 : node2621;
											assign node2621 = (inp[2]) ? node2629 : node2622;
												assign node2622 = (inp[14]) ? 4'b0001 : node2623;
													assign node2623 = (inp[1]) ? 4'b0000 : node2624;
														assign node2624 = (inp[6]) ? 4'b0000 : 4'b1000;
												assign node2629 = (inp[6]) ? node2633 : node2630;
													assign node2630 = (inp[14]) ? 4'b0001 : 4'b1001;
													assign node2633 = (inp[13]) ? 4'b0001 : node2634;
														assign node2634 = (inp[1]) ? 4'b0001 : 4'b1001;
											assign node2638 = (inp[2]) ? node2646 : node2639;
												assign node2639 = (inp[14]) ? node2641 : 4'b0001;
													assign node2641 = (inp[13]) ? node2643 : 4'b1000;
														assign node2643 = (inp[11]) ? 4'b0000 : 4'b0000;
												assign node2646 = (inp[13]) ? 4'b1000 : node2647;
													assign node2647 = (inp[1]) ? node2649 : 4'b0000;
														assign node2649 = (inp[6]) ? 4'b0000 : 4'b1000;
								assign node2653 = (inp[10]) ? node2743 : node2654;
									assign node2654 = (inp[6]) ? node2698 : node2655;
										assign node2655 = (inp[11]) ? node2679 : node2656;
											assign node2656 = (inp[13]) ? node2668 : node2657;
												assign node2657 = (inp[1]) ? node2663 : node2658;
													assign node2658 = (inp[8]) ? node2660 : 4'b1001;
														assign node2660 = (inp[7]) ? 4'b1000 : 4'b1001;
													assign node2663 = (inp[14]) ? node2665 : 4'b1000;
														assign node2665 = (inp[2]) ? 4'b1000 : 4'b0001;
												assign node2668 = (inp[14]) ? node2672 : node2669;
													assign node2669 = (inp[8]) ? 4'b0000 : 4'b1000;
													assign node2672 = (inp[8]) ? node2676 : node2673;
														assign node2673 = (inp[7]) ? 4'b0001 : 4'b0000;
														assign node2676 = (inp[7]) ? 4'b0000 : 4'b0001;
											assign node2679 = (inp[8]) ? node2689 : node2680;
												assign node2680 = (inp[14]) ? node2686 : node2681;
													assign node2681 = (inp[13]) ? node2683 : 4'b0001;
														assign node2683 = (inp[2]) ? 4'b1101 : 4'b0000;
													assign node2686 = (inp[7]) ? 4'b0001 : 4'b0000;
												assign node2689 = (inp[14]) ? node2695 : node2690;
													assign node2690 = (inp[7]) ? 4'b1101 : node2691;
														assign node2691 = (inp[2]) ? 4'b0001 : 4'b0000;
													assign node2695 = (inp[7]) ? 4'b1100 : 4'b1101;
										assign node2698 = (inp[11]) ? node2720 : node2699;
											assign node2699 = (inp[13]) ? node2709 : node2700;
												assign node2700 = (inp[1]) ? node2704 : node2701;
													assign node2701 = (inp[8]) ? 4'b0000 : 4'b0001;
													assign node2704 = (inp[7]) ? node2706 : 4'b0000;
														assign node2706 = (inp[8]) ? 4'b1100 : 4'b1101;
												assign node2709 = (inp[7]) ? node2715 : node2710;
													assign node2710 = (inp[1]) ? 4'b1101 : node2711;
														assign node2711 = (inp[14]) ? 4'b1101 : 4'b0000;
													assign node2715 = (inp[14]) ? 4'b1100 : node2716;
														assign node2716 = (inp[1]) ? 4'b1100 : 4'b1100;
											assign node2720 = (inp[1]) ? node2734 : node2721;
												assign node2721 = (inp[7]) ? node2729 : node2722;
													assign node2722 = (inp[8]) ? node2726 : node2723;
														assign node2723 = (inp[2]) ? 4'b1100 : 4'b1100;
														assign node2726 = (inp[14]) ? 4'b0101 : 4'b1100;
													assign node2729 = (inp[13]) ? 4'b0101 : node2730;
														assign node2730 = (inp[2]) ? 4'b1101 : 4'b1100;
												assign node2734 = (inp[2]) ? node2736 : 4'b0101;
													assign node2736 = (inp[14]) ? node2740 : node2737;
														assign node2737 = (inp[8]) ? 4'b0100 : 4'b0100;
														assign node2740 = (inp[13]) ? 4'b0100 : 4'b1100;
									assign node2743 = (inp[2]) ? node2781 : node2744;
										assign node2744 = (inp[13]) ? node2754 : node2745;
											assign node2745 = (inp[11]) ? node2749 : node2746;
												assign node2746 = (inp[6]) ? 4'b0100 : 4'b1100;
												assign node2749 = (inp[6]) ? 4'b1100 : node2750;
													assign node2750 = (inp[1]) ? 4'b0100 : 4'b0101;
											assign node2754 = (inp[11]) ? node2766 : node2755;
												assign node2755 = (inp[6]) ? node2761 : node2756;
													assign node2756 = (inp[14]) ? 4'b0101 : node2757;
														assign node2757 = (inp[7]) ? 4'b0100 : 4'b0100;
													assign node2761 = (inp[7]) ? 4'b1101 : node2762;
														assign node2762 = (inp[1]) ? 4'b1100 : 4'b0100;
												assign node2766 = (inp[6]) ? node2774 : node2767;
													assign node2767 = (inp[14]) ? node2771 : node2768;
														assign node2768 = (inp[1]) ? 4'b1100 : 4'b0100;
														assign node2771 = (inp[1]) ? 4'b1100 : 4'b1100;
													assign node2774 = (inp[14]) ? node2778 : node2775;
														assign node2775 = (inp[7]) ? 4'b0101 : 4'b1100;
														assign node2778 = (inp[1]) ? 4'b0100 : 4'b0100;
										assign node2781 = (inp[13]) ? node2805 : node2782;
											assign node2782 = (inp[6]) ? node2796 : node2783;
												assign node2783 = (inp[14]) ? node2791 : node2784;
													assign node2784 = (inp[11]) ? node2788 : node2785;
														assign node2785 = (inp[8]) ? 4'b1100 : 4'b1100;
														assign node2788 = (inp[8]) ? 4'b1100 : 4'b0100;
													assign node2791 = (inp[1]) ? node2793 : 4'b1101;
														assign node2793 = (inp[11]) ? 4'b1101 : 4'b0100;
												assign node2796 = (inp[7]) ? node2800 : node2797;
													assign node2797 = (inp[8]) ? 4'b0101 : 4'b0100;
													assign node2800 = (inp[8]) ? 4'b1100 : node2801;
														assign node2801 = (inp[14]) ? 4'b0101 : 4'b0101;
											assign node2805 = (inp[11]) ? node2817 : node2806;
												assign node2806 = (inp[6]) ? node2814 : node2807;
													assign node2807 = (inp[1]) ? node2811 : node2808;
														assign node2808 = (inp[7]) ? 4'b0100 : 4'b1100;
														assign node2811 = (inp[8]) ? 4'b0100 : 4'b0100;
													assign node2814 = (inp[14]) ? 4'b0100 : 4'b1100;
												assign node2817 = (inp[8]) ? node2821 : node2818;
													assign node2818 = (inp[7]) ? 4'b0101 : 4'b0100;
													assign node2821 = (inp[6]) ? 4'b0101 : 4'b1101;
				assign node2824 = (inp[3]) ? node4182 : node2825;
					assign node2825 = (inp[9]) ? node3481 : node2826;
						assign node2826 = (inp[10]) ? node3150 : node2827;
							assign node2827 = (inp[12]) ? node2977 : node2828;
								assign node2828 = (inp[8]) ? node2902 : node2829;
									assign node2829 = (inp[7]) ? node2865 : node2830;
										assign node2830 = (inp[2]) ? node2850 : node2831;
											assign node2831 = (inp[14]) ? node2843 : node2832;
												assign node2832 = (inp[1]) ? node2838 : node2833;
													assign node2833 = (inp[13]) ? 4'b1101 : node2834;
														assign node2834 = (inp[11]) ? 4'b1101 : 4'b0101;
													assign node2838 = (inp[6]) ? node2840 : 4'b0101;
														assign node2840 = (inp[5]) ? 4'b1101 : 4'b0101;
												assign node2843 = (inp[1]) ? 4'b0100 : node2844;
													assign node2844 = (inp[6]) ? 4'b1100 : node2845;
														assign node2845 = (inp[11]) ? 4'b0100 : 4'b1100;
											assign node2850 = (inp[13]) ? node2858 : node2851;
												assign node2851 = (inp[6]) ? node2855 : node2852;
													assign node2852 = (inp[11]) ? 4'b0100 : 4'b1100;
													assign node2855 = (inp[11]) ? 4'b1100 : 4'b0100;
												assign node2858 = (inp[11]) ? 4'b1100 : node2859;
													assign node2859 = (inp[5]) ? 4'b0100 : node2860;
														assign node2860 = (inp[1]) ? 4'b1100 : 4'b0100;
										assign node2865 = (inp[2]) ? node2885 : node2866;
											assign node2866 = (inp[14]) ? node2878 : node2867;
												assign node2867 = (inp[1]) ? node2873 : node2868;
													assign node2868 = (inp[5]) ? node2870 : 4'b0100;
														assign node2870 = (inp[6]) ? 4'b1100 : 4'b0100;
													assign node2873 = (inp[5]) ? node2875 : 4'b1100;
														assign node2875 = (inp[6]) ? 4'b1100 : 4'b0100;
												assign node2878 = (inp[13]) ? 4'b0101 : node2879;
													assign node2879 = (inp[6]) ? 4'b1101 : node2880;
														assign node2880 = (inp[11]) ? 4'b0101 : 4'b0101;
											assign node2885 = (inp[14]) ? node2891 : node2886;
												assign node2886 = (inp[5]) ? 4'b0101 : node2887;
													assign node2887 = (inp[6]) ? 4'b1101 : 4'b0101;
												assign node2891 = (inp[1]) ? node2897 : node2892;
													assign node2892 = (inp[13]) ? node2894 : 4'b1101;
														assign node2894 = (inp[11]) ? 4'b1101 : 4'b0101;
													assign node2897 = (inp[13]) ? 4'b0101 : node2898;
														assign node2898 = (inp[5]) ? 4'b1101 : 4'b0101;
									assign node2902 = (inp[7]) ? node2934 : node2903;
										assign node2903 = (inp[14]) ? node2917 : node2904;
											assign node2904 = (inp[2]) ? node2912 : node2905;
												assign node2905 = (inp[11]) ? node2909 : node2906;
													assign node2906 = (inp[6]) ? 4'b0100 : 4'b1100;
													assign node2909 = (inp[6]) ? 4'b1100 : 4'b0100;
												assign node2912 = (inp[1]) ? 4'b1101 : node2913;
													assign node2913 = (inp[5]) ? 4'b0101 : 4'b1101;
											assign node2917 = (inp[6]) ? node2927 : node2918;
												assign node2918 = (inp[11]) ? node2924 : node2919;
													assign node2919 = (inp[13]) ? 4'b0101 : node2920;
														assign node2920 = (inp[1]) ? 4'b0101 : 4'b1101;
													assign node2924 = (inp[1]) ? 4'b1101 : 4'b0101;
												assign node2927 = (inp[11]) ? node2929 : 4'b1101;
													assign node2929 = (inp[2]) ? 4'b0101 : node2930;
														assign node2930 = (inp[5]) ? 4'b0101 : 4'b1101;
										assign node2934 = (inp[2]) ? node2954 : node2935;
											assign node2935 = (inp[14]) ? node2945 : node2936;
												assign node2936 = (inp[13]) ? node2942 : node2937;
													assign node2937 = (inp[11]) ? 4'b0101 : node2938;
														assign node2938 = (inp[1]) ? 4'b1101 : 4'b0101;
													assign node2942 = (inp[11]) ? 4'b1101 : 4'b0101;
												assign node2945 = (inp[6]) ? node2949 : node2946;
													assign node2946 = (inp[11]) ? 4'b1100 : 4'b0100;
													assign node2949 = (inp[13]) ? 4'b1100 : node2950;
														assign node2950 = (inp[1]) ? 4'b1100 : 4'b0100;
											assign node2954 = (inp[5]) ? node2964 : node2955;
												assign node2955 = (inp[11]) ? node2957 : 4'b1100;
													assign node2957 = (inp[13]) ? node2961 : node2958;
														assign node2958 = (inp[14]) ? 4'b1100 : 4'b1100;
														assign node2961 = (inp[6]) ? 4'b0100 : 4'b1100;
												assign node2964 = (inp[11]) ? node2972 : node2965;
													assign node2965 = (inp[6]) ? node2969 : node2966;
														assign node2966 = (inp[13]) ? 4'b0100 : 4'b0100;
														assign node2969 = (inp[1]) ? 4'b1100 : 4'b0100;
													assign node2972 = (inp[6]) ? 4'b0100 : node2973;
														assign node2973 = (inp[13]) ? 4'b1100 : 4'b0100;
								assign node2977 = (inp[6]) ? node3051 : node2978;
									assign node2978 = (inp[11]) ? node3008 : node2979;
										assign node2979 = (inp[8]) ? node2997 : node2980;
											assign node2980 = (inp[13]) ? node2990 : node2981;
												assign node2981 = (inp[7]) ? node2985 : node2982;
													assign node2982 = (inp[14]) ? 4'b1100 : 4'b1101;
													assign node2985 = (inp[1]) ? 4'b0101 : node2986;
														assign node2986 = (inp[2]) ? 4'b1101 : 4'b1100;
												assign node2990 = (inp[1]) ? 4'b0100 : node2991;
													assign node2991 = (inp[7]) ? node2993 : 4'b1100;
														assign node2993 = (inp[2]) ? 4'b0101 : 4'b1100;
											assign node2997 = (inp[7]) ? node3003 : node2998;
												assign node2998 = (inp[1]) ? 4'b0101 : node2999;
													assign node2999 = (inp[13]) ? 4'b0101 : 4'b1101;
												assign node3003 = (inp[2]) ? 4'b0100 : node3004;
													assign node3004 = (inp[14]) ? 4'b1100 : 4'b0101;
										assign node3008 = (inp[1]) ? node3028 : node3009;
											assign node3009 = (inp[13]) ? node3019 : node3010;
												assign node3010 = (inp[5]) ? node3014 : node3011;
													assign node3011 = (inp[2]) ? 4'b0100 : 4'b0101;
													assign node3014 = (inp[14]) ? node3016 : 4'b0100;
														assign node3016 = (inp[7]) ? 4'b0100 : 4'b0100;
												assign node3019 = (inp[2]) ? node3021 : 4'b0100;
													assign node3021 = (inp[7]) ? node3025 : node3022;
														assign node3022 = (inp[8]) ? 4'b1001 : 4'b0100;
														assign node3025 = (inp[8]) ? 4'b1000 : 4'b1001;
											assign node3028 = (inp[13]) ? node3040 : node3029;
												assign node3029 = (inp[7]) ? node3035 : node3030;
													assign node3030 = (inp[8]) ? 4'b1001 : node3031;
														assign node3031 = (inp[14]) ? 4'b0100 : 4'b0101;
													assign node3035 = (inp[8]) ? node3037 : 4'b1001;
														assign node3037 = (inp[14]) ? 4'b1000 : 4'b1001;
												assign node3040 = (inp[14]) ? node3046 : node3041;
													assign node3041 = (inp[7]) ? 4'b1000 : node3042;
														assign node3042 = (inp[5]) ? 4'b1000 : 4'b1001;
													assign node3046 = (inp[7]) ? node3048 : 4'b1000;
														assign node3048 = (inp[8]) ? 4'b1000 : 4'b1001;
									assign node3051 = (inp[11]) ? node3097 : node3052;
										assign node3052 = (inp[1]) ? node3072 : node3053;
											assign node3053 = (inp[13]) ? node3061 : node3054;
												assign node3054 = (inp[5]) ? node3056 : 4'b0101;
													assign node3056 = (inp[2]) ? node3058 : 4'b0101;
														assign node3058 = (inp[14]) ? 4'b0101 : 4'b0100;
												assign node3061 = (inp[8]) ? node3067 : node3062;
													assign node3062 = (inp[2]) ? node3064 : 4'b0100;
														assign node3064 = (inp[7]) ? 4'b1001 : 4'b0100;
													assign node3067 = (inp[7]) ? node3069 : 4'b1001;
														assign node3069 = (inp[2]) ? 4'b1000 : 4'b1001;
											assign node3072 = (inp[13]) ? node3084 : node3073;
												assign node3073 = (inp[2]) ? node3079 : node3074;
													assign node3074 = (inp[7]) ? 4'b1001 : node3075;
														assign node3075 = (inp[5]) ? 4'b0101 : 4'b0100;
													assign node3079 = (inp[7]) ? node3081 : 4'b1001;
														assign node3081 = (inp[8]) ? 4'b1000 : 4'b1001;
												assign node3084 = (inp[7]) ? node3092 : node3085;
													assign node3085 = (inp[5]) ? node3089 : node3086;
														assign node3086 = (inp[14]) ? 4'b1000 : 4'b1001;
														assign node3089 = (inp[8]) ? 4'b1001 : 4'b1000;
													assign node3092 = (inp[8]) ? 4'b1000 : node3093;
														assign node3093 = (inp[2]) ? 4'b1001 : 4'b1000;
										assign node3097 = (inp[13]) ? node3125 : node3098;
											assign node3098 = (inp[1]) ? node3112 : node3099;
												assign node3099 = (inp[8]) ? node3105 : node3100;
													assign node3100 = (inp[2]) ? 4'b1001 : node3101;
														assign node3101 = (inp[14]) ? 4'b1001 : 4'b1000;
													assign node3105 = (inp[2]) ? node3109 : node3106;
														assign node3106 = (inp[5]) ? 4'b1001 : 4'b1000;
														assign node3109 = (inp[7]) ? 4'b1000 : 4'b1001;
												assign node3112 = (inp[8]) ? node3120 : node3113;
													assign node3113 = (inp[7]) ? node3117 : node3114;
														assign node3114 = (inp[2]) ? 4'b1000 : 4'b1000;
														assign node3117 = (inp[2]) ? 4'b0001 : 4'b0000;
													assign node3120 = (inp[7]) ? node3122 : 4'b0001;
														assign node3122 = (inp[2]) ? 4'b0000 : 4'b0000;
											assign node3125 = (inp[14]) ? node3135 : node3126;
												assign node3126 = (inp[5]) ? node3130 : node3127;
													assign node3127 = (inp[2]) ? 4'b0001 : 4'b1001;
													assign node3130 = (inp[2]) ? 4'b0001 : node3131;
														assign node3131 = (inp[8]) ? 4'b0001 : 4'b0000;
												assign node3135 = (inp[2]) ? node3143 : node3136;
													assign node3136 = (inp[7]) ? node3140 : node3137;
														assign node3137 = (inp[1]) ? 4'b0000 : 4'b1000;
														assign node3140 = (inp[8]) ? 4'b0000 : 4'b0001;
													assign node3143 = (inp[7]) ? node3147 : node3144;
														assign node3144 = (inp[8]) ? 4'b0001 : 4'b0000;
														assign node3147 = (inp[8]) ? 4'b0000 : 4'b0001;
							assign node3150 = (inp[12]) ? node3316 : node3151;
								assign node3151 = (inp[6]) ? node3231 : node3152;
									assign node3152 = (inp[11]) ? node3188 : node3153;
										assign node3153 = (inp[1]) ? node3173 : node3154;
											assign node3154 = (inp[13]) ? node3162 : node3155;
												assign node3155 = (inp[5]) ? 4'b1101 : node3156;
													assign node3156 = (inp[7]) ? node3158 : 4'b1101;
														assign node3158 = (inp[2]) ? 4'b1100 : 4'b1100;
												assign node3162 = (inp[5]) ? node3168 : node3163;
													assign node3163 = (inp[7]) ? 4'b0100 : node3164;
														assign node3164 = (inp[14]) ? 4'b1100 : 4'b1100;
													assign node3168 = (inp[2]) ? 4'b0101 : node3169;
														assign node3169 = (inp[8]) ? 4'b0100 : 4'b0101;
											assign node3173 = (inp[8]) ? node3181 : node3174;
												assign node3174 = (inp[13]) ? node3176 : 4'b1100;
													assign node3176 = (inp[14]) ? 4'b0100 : node3177;
														assign node3177 = (inp[2]) ? 4'b0100 : 4'b0101;
												assign node3181 = (inp[7]) ? node3185 : node3182;
													assign node3182 = (inp[14]) ? 4'b0101 : 4'b0100;
													assign node3185 = (inp[2]) ? 4'b0100 : 4'b0101;
										assign node3188 = (inp[1]) ? node3210 : node3189;
											assign node3189 = (inp[13]) ? node3199 : node3190;
												assign node3190 = (inp[8]) ? node3196 : node3191;
													assign node3191 = (inp[2]) ? 4'b0100 : node3192;
														assign node3192 = (inp[14]) ? 4'b0101 : 4'b0100;
													assign node3196 = (inp[14]) ? 4'b0100 : 4'b0101;
												assign node3199 = (inp[2]) ? node3205 : node3200;
													assign node3200 = (inp[8]) ? node3202 : 4'b0100;
														assign node3202 = (inp[14]) ? 4'b1001 : 4'b0000;
													assign node3205 = (inp[7]) ? node3207 : 4'b0100;
														assign node3207 = (inp[8]) ? 4'b1000 : 4'b1001;
											assign node3210 = (inp[2]) ? node3222 : node3211;
												assign node3211 = (inp[14]) ? node3217 : node3212;
													assign node3212 = (inp[13]) ? node3214 : 4'b0100;
														assign node3214 = (inp[7]) ? 4'b1000 : 4'b1000;
													assign node3217 = (inp[8]) ? node3219 : 4'b1001;
														assign node3219 = (inp[7]) ? 4'b1000 : 4'b1001;
												assign node3222 = (inp[14]) ? node3228 : node3223;
													assign node3223 = (inp[5]) ? node3225 : 4'b1001;
														assign node3225 = (inp[13]) ? 4'b1000 : 4'b1001;
													assign node3228 = (inp[7]) ? 4'b1000 : 4'b1001;
									assign node3231 = (inp[11]) ? node3269 : node3232;
										assign node3232 = (inp[13]) ? node3252 : node3233;
											assign node3233 = (inp[1]) ? node3241 : node3234;
												assign node3234 = (inp[14]) ? 4'b0101 : node3235;
													assign node3235 = (inp[2]) ? 4'b0100 : node3236;
														assign node3236 = (inp[7]) ? 4'b0100 : 4'b0101;
												assign node3241 = (inp[7]) ? node3247 : node3242;
													assign node3242 = (inp[2]) ? node3244 : 4'b0100;
														assign node3244 = (inp[8]) ? 4'b1001 : 4'b0100;
													assign node3247 = (inp[5]) ? node3249 : 4'b1001;
														assign node3249 = (inp[2]) ? 4'b1000 : 4'b1001;
											assign node3252 = (inp[7]) ? node3264 : node3253;
												assign node3253 = (inp[8]) ? node3259 : node3254;
													assign node3254 = (inp[1]) ? 4'b1001 : node3255;
														assign node3255 = (inp[5]) ? 4'b0100 : 4'b0101;
													assign node3259 = (inp[14]) ? 4'b1001 : node3260;
														assign node3260 = (inp[2]) ? 4'b1001 : 4'b0000;
												assign node3264 = (inp[8]) ? 4'b1000 : node3265;
													assign node3265 = (inp[2]) ? 4'b1001 : 4'b1000;
										assign node3269 = (inp[13]) ? node3295 : node3270;
											assign node3270 = (inp[1]) ? node3284 : node3271;
												assign node3271 = (inp[7]) ? node3279 : node3272;
													assign node3272 = (inp[8]) ? node3276 : node3273;
														assign node3273 = (inp[2]) ? 4'b1000 : 4'b1001;
														assign node3276 = (inp[14]) ? 4'b1001 : 4'b1000;
													assign node3279 = (inp[14]) ? 4'b1000 : node3280;
														assign node3280 = (inp[5]) ? 4'b1001 : 4'b1000;
												assign node3284 = (inp[8]) ? node3290 : node3285;
													assign node3285 = (inp[2]) ? 4'b1000 : node3286;
														assign node3286 = (inp[14]) ? 4'b1000 : 4'b1000;
													assign node3290 = (inp[7]) ? node3292 : 4'b0001;
														assign node3292 = (inp[2]) ? 4'b0000 : 4'b0000;
											assign node3295 = (inp[1]) ? node3305 : node3296;
												assign node3296 = (inp[8]) ? node3302 : node3297;
													assign node3297 = (inp[7]) ? node3299 : 4'b1000;
														assign node3299 = (inp[14]) ? 4'b0001 : 4'b1000;
													assign node3302 = (inp[2]) ? 4'b0001 : 4'b0000;
												assign node3305 = (inp[14]) ? node3309 : node3306;
													assign node3306 = (inp[5]) ? 4'b0000 : 4'b0001;
													assign node3309 = (inp[2]) ? node3313 : node3310;
														assign node3310 = (inp[8]) ? 4'b0000 : 4'b0001;
														assign node3313 = (inp[5]) ? 4'b0001 : 4'b0000;
								assign node3316 = (inp[14]) ? node3404 : node3317;
									assign node3317 = (inp[7]) ? node3361 : node3318;
										assign node3318 = (inp[1]) ? node3344 : node3319;
											assign node3319 = (inp[8]) ? node3331 : node3320;
												assign node3320 = (inp[2]) ? node3326 : node3321;
													assign node3321 = (inp[5]) ? node3323 : 4'b1001;
														assign node3323 = (inp[6]) ? 4'b0001 : 4'b0001;
													assign node3326 = (inp[13]) ? 4'b0000 : node3327;
														assign node3327 = (inp[5]) ? 4'b0000 : 4'b1000;
												assign node3331 = (inp[2]) ? node3337 : node3332;
													assign node3332 = (inp[6]) ? 4'b1000 : node3333;
														assign node3333 = (inp[5]) ? 4'b1000 : 4'b0000;
													assign node3337 = (inp[5]) ? node3341 : node3338;
														assign node3338 = (inp[6]) ? 4'b1001 : 4'b0001;
														assign node3341 = (inp[13]) ? 4'b0001 : 4'b1001;
											assign node3344 = (inp[2]) ? node3354 : node3345;
												assign node3345 = (inp[8]) ? node3349 : node3346;
													assign node3346 = (inp[13]) ? 4'b0001 : 4'b1001;
													assign node3349 = (inp[13]) ? 4'b1000 : node3350;
														assign node3350 = (inp[6]) ? 4'b1000 : 4'b0000;
												assign node3354 = (inp[8]) ? 4'b0001 : node3355;
													assign node3355 = (inp[11]) ? node3357 : 4'b0000;
														assign node3357 = (inp[13]) ? 4'b0000 : 4'b1000;
										assign node3361 = (inp[13]) ? node3387 : node3362;
											assign node3362 = (inp[5]) ? node3376 : node3363;
												assign node3363 = (inp[8]) ? node3371 : node3364;
													assign node3364 = (inp[2]) ? node3368 : node3365;
														assign node3365 = (inp[6]) ? 4'b1000 : 4'b0000;
														assign node3368 = (inp[1]) ? 4'b0001 : 4'b0001;
													assign node3371 = (inp[11]) ? node3373 : 4'b0000;
														assign node3373 = (inp[2]) ? 4'b1000 : 4'b1001;
												assign node3376 = (inp[8]) ? node3382 : node3377;
													assign node3377 = (inp[2]) ? 4'b1001 : node3378;
														assign node3378 = (inp[11]) ? 4'b0000 : 4'b1000;
													assign node3382 = (inp[2]) ? 4'b1000 : node3383;
														assign node3383 = (inp[1]) ? 4'b1001 : 4'b0001;
											assign node3387 = (inp[8]) ? node3395 : node3388;
												assign node3388 = (inp[2]) ? 4'b1001 : node3389;
													assign node3389 = (inp[5]) ? 4'b1000 : node3390;
														assign node3390 = (inp[1]) ? 4'b1000 : 4'b1000;
												assign node3395 = (inp[2]) ? node3399 : node3396;
													assign node3396 = (inp[6]) ? 4'b0001 : 4'b1001;
													assign node3399 = (inp[1]) ? 4'b1000 : node3400;
														assign node3400 = (inp[11]) ? 4'b1000 : 4'b0000;
									assign node3404 = (inp[11]) ? node3446 : node3405;
										assign node3405 = (inp[6]) ? node3421 : node3406;
											assign node3406 = (inp[13]) ? node3416 : node3407;
												assign node3407 = (inp[7]) ? node3413 : node3408;
													assign node3408 = (inp[2]) ? 4'b0001 : node3409;
														assign node3409 = (inp[1]) ? 4'b1000 : 4'b1001;
													assign node3413 = (inp[1]) ? 4'b0000 : 4'b1000;
												assign node3416 = (inp[8]) ? 4'b0000 : node3417;
													assign node3417 = (inp[7]) ? 4'b0001 : 4'b0000;
											assign node3421 = (inp[1]) ? node3431 : node3422;
												assign node3422 = (inp[13]) ? node3426 : node3423;
													assign node3423 = (inp[2]) ? 4'b0001 : 4'b0000;
													assign node3426 = (inp[7]) ? node3428 : 4'b0000;
														assign node3428 = (inp[8]) ? 4'b1000 : 4'b1001;
												assign node3431 = (inp[13]) ? node3439 : node3432;
													assign node3432 = (inp[7]) ? node3436 : node3433;
														assign node3433 = (inp[8]) ? 4'b1001 : 4'b0000;
														assign node3436 = (inp[8]) ? 4'b1000 : 4'b1001;
													assign node3439 = (inp[7]) ? node3443 : node3440;
														assign node3440 = (inp[8]) ? 4'b1001 : 4'b1000;
														assign node3443 = (inp[8]) ? 4'b1000 : 4'b1001;
										assign node3446 = (inp[6]) ? node3460 : node3447;
											assign node3447 = (inp[7]) ? node3455 : node3448;
												assign node3448 = (inp[8]) ? node3450 : 4'b0000;
													assign node3450 = (inp[1]) ? 4'b1001 : node3451;
														assign node3451 = (inp[13]) ? 4'b1001 : 4'b0001;
												assign node3455 = (inp[8]) ? node3457 : 4'b1001;
													assign node3457 = (inp[5]) ? 4'b1000 : 4'b0000;
											assign node3460 = (inp[1]) ? node3472 : node3461;
												assign node3461 = (inp[13]) ? node3467 : node3462;
													assign node3462 = (inp[7]) ? node3464 : 4'b1001;
														assign node3464 = (inp[8]) ? 4'b1000 : 4'b1001;
													assign node3467 = (inp[8]) ? node3469 : 4'b1000;
														assign node3469 = (inp[7]) ? 4'b0000 : 4'b0001;
												assign node3472 = (inp[7]) ? node3478 : node3473;
													assign node3473 = (inp[8]) ? 4'b0001 : node3474;
														assign node3474 = (inp[13]) ? 4'b0000 : 4'b1000;
													assign node3478 = (inp[8]) ? 4'b0000 : 4'b0001;
						assign node3481 = (inp[10]) ? node3829 : node3482;
							assign node3482 = (inp[12]) ? node3658 : node3483;
								assign node3483 = (inp[7]) ? node3571 : node3484;
									assign node3484 = (inp[8]) ? node3530 : node3485;
										assign node3485 = (inp[2]) ? node3509 : node3486;
											assign node3486 = (inp[14]) ? node3498 : node3487;
												assign node3487 = (inp[11]) ? node3493 : node3488;
													assign node3488 = (inp[6]) ? node3490 : 4'b1001;
														assign node3490 = (inp[1]) ? 4'b1001 : 4'b0001;
													assign node3493 = (inp[1]) ? node3495 : 4'b1001;
														assign node3495 = (inp[13]) ? 4'b1001 : 4'b0001;
												assign node3498 = (inp[5]) ? node3504 : node3499;
													assign node3499 = (inp[1]) ? 4'b1000 : node3500;
														assign node3500 = (inp[13]) ? 4'b0000 : 4'b1000;
													assign node3504 = (inp[1]) ? node3506 : 4'b1000;
														assign node3506 = (inp[11]) ? 4'b0000 : 4'b1000;
											assign node3509 = (inp[1]) ? node3523 : node3510;
												assign node3510 = (inp[5]) ? node3518 : node3511;
													assign node3511 = (inp[11]) ? node3515 : node3512;
														assign node3512 = (inp[6]) ? 4'b0000 : 4'b1000;
														assign node3515 = (inp[6]) ? 4'b1000 : 4'b0000;
													assign node3518 = (inp[13]) ? node3520 : 4'b1000;
														assign node3520 = (inp[11]) ? 4'b0000 : 4'b1000;
												assign node3523 = (inp[13]) ? 4'b1000 : node3524;
													assign node3524 = (inp[14]) ? 4'b1000 : node3525;
														assign node3525 = (inp[11]) ? 4'b0000 : 4'b0000;
										assign node3530 = (inp[14]) ? node3550 : node3531;
											assign node3531 = (inp[2]) ? node3543 : node3532;
												assign node3532 = (inp[6]) ? node3538 : node3533;
													assign node3533 = (inp[13]) ? node3535 : 4'b1000;
														assign node3535 = (inp[1]) ? 4'b0000 : 4'b1000;
													assign node3538 = (inp[11]) ? node3540 : 4'b0000;
														assign node3540 = (inp[13]) ? 4'b0000 : 4'b1000;
												assign node3543 = (inp[6]) ? 4'b0001 : node3544;
													assign node3544 = (inp[13]) ? 4'b1001 : node3545;
														assign node3545 = (inp[11]) ? 4'b0001 : 4'b1001;
											assign node3550 = (inp[1]) ? node3562 : node3551;
												assign node3551 = (inp[5]) ? node3557 : node3552;
													assign node3552 = (inp[6]) ? node3554 : 4'b0001;
														assign node3554 = (inp[11]) ? 4'b0001 : 4'b1001;
													assign node3557 = (inp[13]) ? node3559 : 4'b1001;
														assign node3559 = (inp[11]) ? 4'b0001 : 4'b1001;
												assign node3562 = (inp[5]) ? node3564 : 4'b1001;
													assign node3564 = (inp[11]) ? node3568 : node3565;
														assign node3565 = (inp[6]) ? 4'b1001 : 4'b0001;
														assign node3568 = (inp[6]) ? 4'b0001 : 4'b1001;
									assign node3571 = (inp[8]) ? node3621 : node3572;
										assign node3572 = (inp[2]) ? node3598 : node3573;
											assign node3573 = (inp[14]) ? node3589 : node3574;
												assign node3574 = (inp[5]) ? node3582 : node3575;
													assign node3575 = (inp[11]) ? node3579 : node3576;
														assign node3576 = (inp[6]) ? 4'b0000 : 4'b1000;
														assign node3579 = (inp[6]) ? 4'b1000 : 4'b0000;
													assign node3582 = (inp[11]) ? node3586 : node3583;
														assign node3583 = (inp[6]) ? 4'b0000 : 4'b0000;
														assign node3586 = (inp[6]) ? 4'b1000 : 4'b0000;
												assign node3589 = (inp[1]) ? node3591 : 4'b1001;
													assign node3591 = (inp[5]) ? node3595 : node3592;
														assign node3592 = (inp[6]) ? 4'b0001 : 4'b1001;
														assign node3595 = (inp[6]) ? 4'b1001 : 4'b0001;
											assign node3598 = (inp[1]) ? node3610 : node3599;
												assign node3599 = (inp[14]) ? node3605 : node3600;
													assign node3600 = (inp[11]) ? 4'b1001 : node3601;
														assign node3601 = (inp[5]) ? 4'b1001 : 4'b0001;
													assign node3605 = (inp[6]) ? 4'b0001 : node3606;
														assign node3606 = (inp[11]) ? 4'b1001 : 4'b0001;
												assign node3610 = (inp[14]) ? node3616 : node3611;
													assign node3611 = (inp[13]) ? node3613 : 4'b0001;
														assign node3613 = (inp[6]) ? 4'b1001 : 4'b0001;
													assign node3616 = (inp[11]) ? node3618 : 4'b1001;
														assign node3618 = (inp[6]) ? 4'b0001 : 4'b1001;
										assign node3621 = (inp[2]) ? node3639 : node3622;
											assign node3622 = (inp[14]) ? node3628 : node3623;
												assign node3623 = (inp[6]) ? node3625 : 4'b0001;
													assign node3625 = (inp[11]) ? 4'b0001 : 4'b1001;
												assign node3628 = (inp[5]) ? node3634 : node3629;
													assign node3629 = (inp[11]) ? node3631 : 4'b1000;
														assign node3631 = (inp[6]) ? 4'b0000 : 4'b1000;
													assign node3634 = (inp[13]) ? node3636 : 4'b0000;
														assign node3636 = (inp[11]) ? 4'b0000 : 4'b1000;
											assign node3639 = (inp[5]) ? node3647 : node3640;
												assign node3640 = (inp[13]) ? node3642 : 4'b0000;
													assign node3642 = (inp[1]) ? node3644 : 4'b0000;
														assign node3644 = (inp[11]) ? 4'b0000 : 4'b1000;
												assign node3647 = (inp[11]) ? node3651 : node3648;
													assign node3648 = (inp[6]) ? 4'b1000 : 4'b0000;
													assign node3651 = (inp[6]) ? node3655 : node3652;
														assign node3652 = (inp[13]) ? 4'b1000 : 4'b0000;
														assign node3655 = (inp[14]) ? 4'b0000 : 4'b0000;
								assign node3658 = (inp[11]) ? node3736 : node3659;
									assign node3659 = (inp[6]) ? node3697 : node3660;
										assign node3660 = (inp[1]) ? node3676 : node3661;
											assign node3661 = (inp[13]) ? node3669 : node3662;
												assign node3662 = (inp[2]) ? 4'b1001 : node3663;
													assign node3663 = (inp[8]) ? node3665 : 4'b1001;
														assign node3665 = (inp[14]) ? 4'b1001 : 4'b1000;
												assign node3669 = (inp[8]) ? node3673 : node3670;
													assign node3670 = (inp[2]) ? 4'b0001 : 4'b1000;
													assign node3673 = (inp[2]) ? 4'b0000 : 4'b0001;
											assign node3676 = (inp[14]) ? node3684 : node3677;
												assign node3677 = (inp[8]) ? 4'b0001 : node3678;
													assign node3678 = (inp[13]) ? 4'b0001 : node3679;
														assign node3679 = (inp[2]) ? 4'b1000 : 4'b1001;
												assign node3684 = (inp[5]) ? node3690 : node3685;
													assign node3685 = (inp[2]) ? node3687 : 4'b0000;
														assign node3687 = (inp[7]) ? 4'b0001 : 4'b0000;
													assign node3690 = (inp[7]) ? node3694 : node3691;
														assign node3691 = (inp[8]) ? 4'b0001 : 4'b0000;
														assign node3694 = (inp[8]) ? 4'b0000 : 4'b0001;
										assign node3697 = (inp[13]) ? node3717 : node3698;
											assign node3698 = (inp[2]) ? node3706 : node3699;
												assign node3699 = (inp[1]) ? 4'b0000 : node3700;
													assign node3700 = (inp[14]) ? node3702 : 4'b0000;
														assign node3702 = (inp[5]) ? 4'b0000 : 4'b0001;
												assign node3706 = (inp[8]) ? node3710 : node3707;
													assign node3707 = (inp[7]) ? 4'b0001 : 4'b0000;
													assign node3710 = (inp[7]) ? node3714 : node3711;
														assign node3711 = (inp[14]) ? 4'b1111 : 4'b1101;
														assign node3714 = (inp[14]) ? 4'b1100 : 4'b1110;
											assign node3717 = (inp[5]) ? node3725 : node3718;
												assign node3718 = (inp[1]) ? 4'b1101 : node3719;
													assign node3719 = (inp[7]) ? node3721 : 4'b0000;
														assign node3721 = (inp[2]) ? 4'b1100 : 4'b1100;
												assign node3725 = (inp[1]) ? node3731 : node3726;
													assign node3726 = (inp[8]) ? node3728 : 4'b0000;
														assign node3728 = (inp[2]) ? 4'b1110 : 4'b0000;
													assign node3731 = (inp[2]) ? 4'b1111 : node3732;
														assign node3732 = (inp[7]) ? 4'b1111 : 4'b1110;
									assign node3736 = (inp[5]) ? node3774 : node3737;
										assign node3737 = (inp[6]) ? node3757 : node3738;
											assign node3738 = (inp[13]) ? node3748 : node3739;
												assign node3739 = (inp[1]) ? node3745 : node3740;
													assign node3740 = (inp[8]) ? 4'b0001 : node3741;
														assign node3741 = (inp[7]) ? 4'b0001 : 4'b0000;
													assign node3745 = (inp[7]) ? 4'b1100 : 4'b0000;
												assign node3748 = (inp[2]) ? node3754 : node3749;
													assign node3749 = (inp[7]) ? node3751 : 4'b0000;
														assign node3751 = (inp[14]) ? 4'b1101 : 4'b0000;
													assign node3754 = (inp[8]) ? 4'b1101 : 4'b1100;
											assign node3757 = (inp[1]) ? node3765 : node3758;
												assign node3758 = (inp[14]) ? 4'b1101 : node3759;
													assign node3759 = (inp[13]) ? node3761 : 4'b1100;
														assign node3761 = (inp[2]) ? 4'b0100 : 4'b1100;
												assign node3765 = (inp[13]) ? node3767 : 4'b0101;
													assign node3767 = (inp[7]) ? node3771 : node3768;
														assign node3768 = (inp[8]) ? 4'b0101 : 4'b0100;
														assign node3771 = (inp[8]) ? 4'b0100 : 4'b0101;
										assign node3774 = (inp[6]) ? node3802 : node3775;
											assign node3775 = (inp[1]) ? node3789 : node3776;
												assign node3776 = (inp[13]) ? node3782 : node3777;
													assign node3777 = (inp[7]) ? node3779 : 4'b0000;
														assign node3779 = (inp[14]) ? 4'b0001 : 4'b0000;
													assign node3782 = (inp[7]) ? node3786 : node3783;
														assign node3783 = (inp[8]) ? 4'b0000 : 4'b0000;
														assign node3786 = (inp[8]) ? 4'b1110 : 4'b1111;
												assign node3789 = (inp[2]) ? node3795 : node3790;
													assign node3790 = (inp[13]) ? node3792 : 4'b0001;
														assign node3792 = (inp[8]) ? 4'b1110 : 4'b1110;
													assign node3795 = (inp[8]) ? node3799 : node3796;
														assign node3796 = (inp[7]) ? 4'b1111 : 4'b1110;
														assign node3799 = (inp[7]) ? 4'b1110 : 4'b1111;
											assign node3802 = (inp[13]) ? node3816 : node3803;
												assign node3803 = (inp[2]) ? node3809 : node3804;
													assign node3804 = (inp[1]) ? 4'b1110 : node3805;
														assign node3805 = (inp[8]) ? 4'b1111 : 4'b1110;
													assign node3809 = (inp[7]) ? node3813 : node3810;
														assign node3810 = (inp[1]) ? 4'b1110 : 4'b1111;
														assign node3813 = (inp[1]) ? 4'b0111 : 4'b1111;
												assign node3816 = (inp[1]) ? node3822 : node3817;
													assign node3817 = (inp[7]) ? node3819 : 4'b1110;
														assign node3819 = (inp[8]) ? 4'b0110 : 4'b0111;
													assign node3822 = (inp[7]) ? node3826 : node3823;
														assign node3823 = (inp[14]) ? 4'b0111 : 4'b0110;
														assign node3826 = (inp[8]) ? 4'b0110 : 4'b0111;
							assign node3829 = (inp[5]) ? node3999 : node3830;
								assign node3830 = (inp[12]) ? node3916 : node3831;
									assign node3831 = (inp[11]) ? node3871 : node3832;
										assign node3832 = (inp[6]) ? node3852 : node3833;
											assign node3833 = (inp[1]) ? node3843 : node3834;
												assign node3834 = (inp[14]) ? node3836 : 4'b1001;
													assign node3836 = (inp[8]) ? node3840 : node3837;
														assign node3837 = (inp[7]) ? 4'b1001 : 4'b1000;
														assign node3840 = (inp[7]) ? 4'b1000 : 4'b0001;
												assign node3843 = (inp[13]) ? node3847 : node3844;
													assign node3844 = (inp[8]) ? 4'b0001 : 4'b1000;
													assign node3847 = (inp[7]) ? node3849 : 4'b0000;
														assign node3849 = (inp[8]) ? 4'b0000 : 4'b0001;
											assign node3852 = (inp[13]) ? node3862 : node3853;
												assign node3853 = (inp[1]) ? node3855 : 4'b0001;
													assign node3855 = (inp[14]) ? node3859 : node3856;
														assign node3856 = (inp[8]) ? 4'b1101 : 4'b0000;
														assign node3859 = (inp[8]) ? 4'b1100 : 4'b1101;
												assign node3862 = (inp[2]) ? 4'b1101 : node3863;
													assign node3863 = (inp[8]) ? node3867 : node3864;
														assign node3864 = (inp[7]) ? 4'b0000 : 4'b1100;
														assign node3867 = (inp[14]) ? 4'b1100 : 4'b1101;
										assign node3871 = (inp[6]) ? node3893 : node3872;
											assign node3872 = (inp[1]) ? node3880 : node3873;
												assign node3873 = (inp[13]) ? 4'b1101 : node3874;
													assign node3874 = (inp[2]) ? node3876 : 4'b0000;
														assign node3876 = (inp[7]) ? 4'b0000 : 4'b0001;
												assign node3880 = (inp[2]) ? node3886 : node3881;
													assign node3881 = (inp[8]) ? node3883 : 4'b1101;
														assign node3883 = (inp[14]) ? 4'b1101 : 4'b1100;
													assign node3886 = (inp[8]) ? node3890 : node3887;
														assign node3887 = (inp[13]) ? 4'b1100 : 4'b0000;
														assign node3890 = (inp[7]) ? 4'b1100 : 4'b1101;
											assign node3893 = (inp[1]) ? node3907 : node3894;
												assign node3894 = (inp[14]) ? node3902 : node3895;
													assign node3895 = (inp[2]) ? node3899 : node3896;
														assign node3896 = (inp[8]) ? 4'b1100 : 4'b1101;
														assign node3899 = (inp[8]) ? 4'b1101 : 4'b1100;
													assign node3902 = (inp[2]) ? node3904 : 4'b1100;
														assign node3904 = (inp[8]) ? 4'b0100 : 4'b1100;
												assign node3907 = (inp[13]) ? node3909 : 4'b0100;
													assign node3909 = (inp[14]) ? node3913 : node3910;
														assign node3910 = (inp[2]) ? 4'b0100 : 4'b0101;
														assign node3913 = (inp[2]) ? 4'b0101 : 4'b0100;
									assign node3916 = (inp[1]) ? node3954 : node3917;
										assign node3917 = (inp[6]) ? node3937 : node3918;
											assign node3918 = (inp[11]) ? node3930 : node3919;
												assign node3919 = (inp[14]) ? node3925 : node3920;
													assign node3920 = (inp[2]) ? 4'b1100 : node3921;
														assign node3921 = (inp[8]) ? 4'b1100 : 4'b1100;
													assign node3925 = (inp[13]) ? node3927 : 4'b1101;
														assign node3927 = (inp[8]) ? 4'b0100 : 4'b1100;
												assign node3930 = (inp[13]) ? node3932 : 4'b0100;
													assign node3932 = (inp[8]) ? 4'b1101 : node3933;
														assign node3933 = (inp[2]) ? 4'b1101 : 4'b0101;
											assign node3937 = (inp[11]) ? node3945 : node3938;
												assign node3938 = (inp[13]) ? node3942 : node3939;
													assign node3939 = (inp[2]) ? 4'b0100 : 4'b0101;
													assign node3942 = (inp[8]) ? 4'b1101 : 4'b0101;
												assign node3945 = (inp[13]) ? node3951 : node3946;
													assign node3946 = (inp[14]) ? 4'b1101 : node3947;
														assign node3947 = (inp[8]) ? 4'b1100 : 4'b1101;
													assign node3951 = (inp[2]) ? 4'b0101 : 4'b1100;
										assign node3954 = (inp[14]) ? node3974 : node3955;
											assign node3955 = (inp[11]) ? node3969 : node3956;
												assign node3956 = (inp[6]) ? node3964 : node3957;
													assign node3957 = (inp[7]) ? node3961 : node3958;
														assign node3958 = (inp[13]) ? 4'b0100 : 4'b1100;
														assign node3961 = (inp[8]) ? 4'b0101 : 4'b0100;
													assign node3964 = (inp[13]) ? 4'b1100 : node3965;
														assign node3965 = (inp[7]) ? 4'b0100 : 4'b0100;
												assign node3969 = (inp[2]) ? 4'b0100 : node3970;
													assign node3970 = (inp[8]) ? 4'b1100 : 4'b1101;
											assign node3974 = (inp[13]) ? node3988 : node3975;
												assign node3975 = (inp[7]) ? node3983 : node3976;
													assign node3976 = (inp[8]) ? node3980 : node3977;
														assign node3977 = (inp[2]) ? 4'b0100 : 4'b1100;
														assign node3980 = (inp[6]) ? 4'b1101 : 4'b0101;
													assign node3983 = (inp[2]) ? node3985 : 4'b1101;
														assign node3985 = (inp[6]) ? 4'b0101 : 4'b1101;
												assign node3988 = (inp[11]) ? node3994 : node3989;
													assign node3989 = (inp[8]) ? 4'b1100 : node3990;
														assign node3990 = (inp[7]) ? 4'b1101 : 4'b1100;
													assign node3994 = (inp[7]) ? 4'b0100 : node3995;
														assign node3995 = (inp[8]) ? 4'b1101 : 4'b1100;
								assign node3999 = (inp[12]) ? node4095 : node4000;
									assign node4000 = (inp[6]) ? node4046 : node4001;
										assign node4001 = (inp[11]) ? node4023 : node4002;
											assign node4002 = (inp[7]) ? node4012 : node4003;
												assign node4003 = (inp[8]) ? node4009 : node4004;
													assign node4004 = (inp[1]) ? node4006 : 4'b1000;
														assign node4006 = (inp[2]) ? 4'b1000 : 4'b1001;
													assign node4009 = (inp[13]) ? 4'b0001 : 4'b1001;
												assign node4012 = (inp[13]) ? node4018 : node4013;
													assign node4013 = (inp[1]) ? node4015 : 4'b1000;
														assign node4015 = (inp[2]) ? 4'b0001 : 4'b0000;
													assign node4018 = (inp[14]) ? node4020 : 4'b0001;
														assign node4020 = (inp[8]) ? 4'b0000 : 4'b0001;
											assign node4023 = (inp[1]) ? node4035 : node4024;
												assign node4024 = (inp[13]) ? node4030 : node4025;
													assign node4025 = (inp[8]) ? node4027 : 4'b0000;
														assign node4027 = (inp[7]) ? 4'b0000 : 4'b0001;
													assign node4030 = (inp[2]) ? node4032 : 4'b0000;
														assign node4032 = (inp[7]) ? 4'b1110 : 4'b1111;
												assign node4035 = (inp[8]) ? node4041 : node4036;
													assign node4036 = (inp[13]) ? node4038 : 4'b0000;
														assign node4038 = (inp[14]) ? 4'b1111 : 4'b1110;
													assign node4041 = (inp[7]) ? node4043 : 4'b1111;
														assign node4043 = (inp[13]) ? 4'b1110 : 4'b1110;
										assign node4046 = (inp[11]) ? node4070 : node4047;
											assign node4047 = (inp[1]) ? node4059 : node4048;
												assign node4048 = (inp[13]) ? node4054 : node4049;
													assign node4049 = (inp[14]) ? 4'b0001 : node4050;
														assign node4050 = (inp[2]) ? 4'b0000 : 4'b0001;
													assign node4054 = (inp[7]) ? node4056 : 4'b0000;
														assign node4056 = (inp[8]) ? 4'b1110 : 4'b0000;
												assign node4059 = (inp[13]) ? node4065 : node4060;
													assign node4060 = (inp[2]) ? 4'b1111 : node4061;
														assign node4061 = (inp[7]) ? 4'b1110 : 4'b0001;
													assign node4065 = (inp[7]) ? 4'b1110 : node4066;
														assign node4066 = (inp[8]) ? 4'b1110 : 4'b1110;
											assign node4070 = (inp[1]) ? node4082 : node4071;
												assign node4071 = (inp[14]) ? node4077 : node4072;
													assign node4072 = (inp[2]) ? 4'b1111 : node4073;
														assign node4073 = (inp[8]) ? 4'b1110 : 4'b1110;
													assign node4077 = (inp[8]) ? node4079 : 4'b1110;
														assign node4079 = (inp[7]) ? 4'b0110 : 4'b0111;
												assign node4082 = (inp[8]) ? node4090 : node4083;
													assign node4083 = (inp[2]) ? node4087 : node4084;
														assign node4084 = (inp[13]) ? 4'b0110 : 4'b0111;
														assign node4087 = (inp[14]) ? 4'b1110 : 4'b0110;
													assign node4090 = (inp[7]) ? node4092 : 4'b0111;
														assign node4092 = (inp[14]) ? 4'b0110 : 4'b0111;
									assign node4095 = (inp[6]) ? node4135 : node4096;
										assign node4096 = (inp[13]) ? node4110 : node4097;
											assign node4097 = (inp[11]) ? node4103 : node4098;
												assign node4098 = (inp[2]) ? node4100 : 4'b1110;
													assign node4100 = (inp[1]) ? 4'b0111 : 4'b1111;
												assign node4103 = (inp[1]) ? node4105 : 4'b0110;
													assign node4105 = (inp[7]) ? node4107 : 4'b0110;
														assign node4107 = (inp[2]) ? 4'b1110 : 4'b1111;
											assign node4110 = (inp[2]) ? node4124 : node4111;
												assign node4111 = (inp[8]) ? node4119 : node4112;
													assign node4112 = (inp[11]) ? node4116 : node4113;
														assign node4113 = (inp[1]) ? 4'b0111 : 4'b1110;
														assign node4116 = (inp[1]) ? 4'b1110 : 4'b0110;
													assign node4119 = (inp[11]) ? 4'b1111 : node4120;
														assign node4120 = (inp[14]) ? 4'b0110 : 4'b1110;
												assign node4124 = (inp[11]) ? node4128 : node4125;
													assign node4125 = (inp[7]) ? 4'b0110 : 4'b1110;
													assign node4128 = (inp[7]) ? node4132 : node4129;
														assign node4129 = (inp[14]) ? 4'b1110 : 4'b0110;
														assign node4132 = (inp[8]) ? 4'b1110 : 4'b1111;
										assign node4135 = (inp[11]) ? node4153 : node4136;
											assign node4136 = (inp[1]) ? node4146 : node4137;
												assign node4137 = (inp[8]) ? 4'b0110 : node4138;
													assign node4138 = (inp[7]) ? node4142 : node4139;
														assign node4139 = (inp[2]) ? 4'b0110 : 4'b0111;
														assign node4142 = (inp[2]) ? 4'b1111 : 4'b0110;
												assign node4146 = (inp[8]) ? 4'b1110 : node4147;
													assign node4147 = (inp[13]) ? 4'b1110 : node4148;
														assign node4148 = (inp[14]) ? 4'b0110 : 4'b0111;
											assign node4153 = (inp[1]) ? node4169 : node4154;
												assign node4154 = (inp[14]) ? node4162 : node4155;
													assign node4155 = (inp[8]) ? node4159 : node4156;
														assign node4156 = (inp[7]) ? 4'b1110 : 4'b1111;
														assign node4159 = (inp[7]) ? 4'b1111 : 4'b1110;
													assign node4162 = (inp[13]) ? node4166 : node4163;
														assign node4163 = (inp[8]) ? 4'b1111 : 4'b1110;
														assign node4166 = (inp[8]) ? 4'b0110 : 4'b0111;
												assign node4169 = (inp[7]) ? node4177 : node4170;
													assign node4170 = (inp[13]) ? node4174 : node4171;
														assign node4171 = (inp[14]) ? 4'b0111 : 4'b1110;
														assign node4174 = (inp[14]) ? 4'b0110 : 4'b0111;
													assign node4177 = (inp[8]) ? node4179 : 4'b0111;
														assign node4179 = (inp[13]) ? 4'b0111 : 4'b0110;
					assign node4182 = (inp[5]) ? node4952 : node4183;
						assign node4183 = (inp[9]) ? node4579 : node4184;
							assign node4184 = (inp[10]) ? node4388 : node4185;
								assign node4185 = (inp[12]) ? node4287 : node4186;
									assign node4186 = (inp[2]) ? node4236 : node4187;
										assign node4187 = (inp[11]) ? node4211 : node4188;
											assign node4188 = (inp[8]) ? node4200 : node4189;
												assign node4189 = (inp[13]) ? node4195 : node4190;
													assign node4190 = (inp[1]) ? node4192 : 4'b1101;
														assign node4192 = (inp[14]) ? 4'b0100 : 4'b0101;
													assign node4195 = (inp[7]) ? node4197 : 4'b1100;
														assign node4197 = (inp[14]) ? 4'b0101 : 4'b0100;
												assign node4200 = (inp[13]) ? node4206 : node4201;
													assign node4201 = (inp[6]) ? 4'b0100 : node4202;
														assign node4202 = (inp[14]) ? 4'b0100 : 4'b1100;
													assign node4206 = (inp[6]) ? 4'b0100 : node4207;
														assign node4207 = (inp[1]) ? 4'b0100 : 4'b0101;
											assign node4211 = (inp[1]) ? node4223 : node4212;
												assign node4212 = (inp[13]) ? node4218 : node4213;
													assign node4213 = (inp[6]) ? 4'b1101 : node4214;
														assign node4214 = (inp[14]) ? 4'b0101 : 4'b0100;
													assign node4218 = (inp[6]) ? node4220 : 4'b1101;
														assign node4220 = (inp[8]) ? 4'b1100 : 4'b1100;
												assign node4223 = (inp[6]) ? node4231 : node4224;
													assign node4224 = (inp[13]) ? node4228 : node4225;
														assign node4225 = (inp[8]) ? 4'b1101 : 4'b0100;
														assign node4228 = (inp[14]) ? 4'b1100 : 4'b1101;
													assign node4231 = (inp[8]) ? 4'b0100 : node4232;
														assign node4232 = (inp[7]) ? 4'b0101 : 4'b0100;
										assign node4236 = (inp[13]) ? node4262 : node4237;
											assign node4237 = (inp[14]) ? node4249 : node4238;
												assign node4238 = (inp[8]) ? node4244 : node4239;
													assign node4239 = (inp[7]) ? 4'b1101 : node4240;
														assign node4240 = (inp[11]) ? 4'b0100 : 4'b1100;
													assign node4244 = (inp[1]) ? 4'b0100 : node4245;
														assign node4245 = (inp[6]) ? 4'b0100 : 4'b0100;
												assign node4249 = (inp[6]) ? node4257 : node4250;
													assign node4250 = (inp[11]) ? node4254 : node4251;
														assign node4251 = (inp[8]) ? 4'b1100 : 4'b1100;
														assign node4254 = (inp[8]) ? 4'b1100 : 4'b0100;
													assign node4257 = (inp[7]) ? 4'b0101 : node4258;
														assign node4258 = (inp[1]) ? 4'b1101 : 4'b0101;
											assign node4262 = (inp[1]) ? node4272 : node4263;
												assign node4263 = (inp[7]) ? node4269 : node4264;
													assign node4264 = (inp[8]) ? node4266 : 4'b0100;
														assign node4266 = (inp[11]) ? 4'b0101 : 4'b0101;
													assign node4269 = (inp[8]) ? 4'b0100 : 4'b1101;
												assign node4272 = (inp[14]) ? node4280 : node4273;
													assign node4273 = (inp[8]) ? node4277 : node4274;
														assign node4274 = (inp[7]) ? 4'b0101 : 4'b0100;
														assign node4277 = (inp[7]) ? 4'b1100 : 4'b1101;
													assign node4280 = (inp[7]) ? node4284 : node4281;
														assign node4281 = (inp[8]) ? 4'b0101 : 4'b0100;
														assign node4284 = (inp[6]) ? 4'b1100 : 4'b0100;
									assign node4287 = (inp[11]) ? node4337 : node4288;
										assign node4288 = (inp[6]) ? node4314 : node4289;
											assign node4289 = (inp[1]) ? node4301 : node4290;
												assign node4290 = (inp[13]) ? node4296 : node4291;
													assign node4291 = (inp[14]) ? 4'b1101 : node4292;
														assign node4292 = (inp[7]) ? 4'b1100 : 4'b1100;
													assign node4296 = (inp[8]) ? node4298 : 4'b1100;
														assign node4298 = (inp[2]) ? 4'b0100 : 4'b0100;
												assign node4301 = (inp[13]) ? node4309 : node4302;
													assign node4302 = (inp[8]) ? node4306 : node4303;
														assign node4303 = (inp[14]) ? 4'b0101 : 4'b1100;
														assign node4306 = (inp[14]) ? 4'b0100 : 4'b0101;
													assign node4309 = (inp[7]) ? 4'b0100 : node4310;
														assign node4310 = (inp[14]) ? 4'b0100 : 4'b0101;
											assign node4314 = (inp[1]) ? node4330 : node4315;
												assign node4315 = (inp[13]) ? node4323 : node4316;
													assign node4316 = (inp[8]) ? node4320 : node4317;
														assign node4317 = (inp[7]) ? 4'b0100 : 4'b0100;
														assign node4320 = (inp[14]) ? 4'b0101 : 4'b0100;
													assign node4323 = (inp[2]) ? node4327 : node4324;
														assign node4324 = (inp[8]) ? 4'b0000 : 4'b0100;
														assign node4327 = (inp[14]) ? 4'b1000 : 4'b1001;
												assign node4330 = (inp[7]) ? node4334 : node4331;
													assign node4331 = (inp[8]) ? 4'b1001 : 4'b1000;
													assign node4334 = (inp[8]) ? 4'b1000 : 4'b1001;
										assign node4337 = (inp[6]) ? node4363 : node4338;
											assign node4338 = (inp[1]) ? node4350 : node4339;
												assign node4339 = (inp[13]) ? node4345 : node4340;
													assign node4340 = (inp[7]) ? 4'b0101 : node4341;
														assign node4341 = (inp[14]) ? 4'b0100 : 4'b0101;
													assign node4345 = (inp[8]) ? 4'b1001 : node4346;
														assign node4346 = (inp[7]) ? 4'b1001 : 4'b0100;
												assign node4350 = (inp[7]) ? node4356 : node4351;
													assign node4351 = (inp[13]) ? 4'b1000 : node4352;
														assign node4352 = (inp[2]) ? 4'b0000 : 4'b0100;
													assign node4356 = (inp[14]) ? node4360 : node4357;
														assign node4357 = (inp[2]) ? 4'b1000 : 4'b1000;
														assign node4360 = (inp[8]) ? 4'b1000 : 4'b1001;
											assign node4363 = (inp[13]) ? node4377 : node4364;
												assign node4364 = (inp[1]) ? node4372 : node4365;
													assign node4365 = (inp[8]) ? node4369 : node4366;
														assign node4366 = (inp[7]) ? 4'b1001 : 4'b1000;
														assign node4369 = (inp[7]) ? 4'b1000 : 4'b1001;
													assign node4372 = (inp[7]) ? node4374 : 4'b1000;
														assign node4374 = (inp[2]) ? 4'b0000 : 4'b0001;
												assign node4377 = (inp[8]) ? node4383 : node4378;
													assign node4378 = (inp[7]) ? 4'b0001 : node4379;
														assign node4379 = (inp[1]) ? 4'b0000 : 4'b1000;
													assign node4383 = (inp[2]) ? 4'b0001 : node4384;
														assign node4384 = (inp[1]) ? 4'b0000 : 4'b0001;
								assign node4388 = (inp[12]) ? node4486 : node4389;
									assign node4389 = (inp[13]) ? node4439 : node4390;
										assign node4390 = (inp[6]) ? node4418 : node4391;
											assign node4391 = (inp[11]) ? node4405 : node4392;
												assign node4392 = (inp[1]) ? node4398 : node4393;
													assign node4393 = (inp[7]) ? 4'b1101 : node4394;
														assign node4394 = (inp[14]) ? 4'b1100 : 4'b1101;
													assign node4398 = (inp[7]) ? node4402 : node4399;
														assign node4399 = (inp[14]) ? 4'b1100 : 4'b0100;
														assign node4402 = (inp[8]) ? 4'b0100 : 4'b0101;
												assign node4405 = (inp[1]) ? node4411 : node4406;
													assign node4406 = (inp[8]) ? node4408 : 4'b0101;
														assign node4408 = (inp[7]) ? 4'b0100 : 4'b0101;
													assign node4411 = (inp[8]) ? node4415 : node4412;
														assign node4412 = (inp[7]) ? 4'b0100 : 4'b0100;
														assign node4415 = (inp[7]) ? 4'b1000 : 4'b1001;
											assign node4418 = (inp[11]) ? node4430 : node4419;
												assign node4419 = (inp[1]) ? node4425 : node4420;
													assign node4420 = (inp[8]) ? 4'b0100 : node4421;
														assign node4421 = (inp[14]) ? 4'b0100 : 4'b0101;
													assign node4425 = (inp[8]) ? node4427 : 4'b0100;
														assign node4427 = (inp[7]) ? 4'b1000 : 4'b1001;
												assign node4430 = (inp[2]) ? node4436 : node4431;
													assign node4431 = (inp[8]) ? 4'b0000 : node4432;
														assign node4432 = (inp[14]) ? 4'b1000 : 4'b1000;
													assign node4436 = (inp[1]) ? 4'b0001 : 4'b1001;
										assign node4439 = (inp[6]) ? node4461 : node4440;
											assign node4440 = (inp[11]) ? node4448 : node4441;
												assign node4441 = (inp[8]) ? node4443 : 4'b1100;
													assign node4443 = (inp[14]) ? node4445 : 4'b1100;
														assign node4445 = (inp[7]) ? 4'b0100 : 4'b0101;
												assign node4448 = (inp[1]) ? node4454 : node4449;
													assign node4449 = (inp[7]) ? node4451 : 4'b0100;
														assign node4451 = (inp[14]) ? 4'b1001 : 4'b0000;
													assign node4454 = (inp[7]) ? node4458 : node4455;
														assign node4455 = (inp[2]) ? 4'b1000 : 4'b1000;
														assign node4458 = (inp[2]) ? 4'b1000 : 4'b1000;
											assign node4461 = (inp[11]) ? node4473 : node4462;
												assign node4462 = (inp[7]) ? node4468 : node4463;
													assign node4463 = (inp[8]) ? 4'b1001 : node4464;
														assign node4464 = (inp[1]) ? 4'b1000 : 4'b0100;
													assign node4468 = (inp[8]) ? 4'b1000 : node4469;
														assign node4469 = (inp[2]) ? 4'b1001 : 4'b1000;
												assign node4473 = (inp[14]) ? node4481 : node4474;
													assign node4474 = (inp[2]) ? node4478 : node4475;
														assign node4475 = (inp[1]) ? 4'b0000 : 4'b1000;
														assign node4478 = (inp[8]) ? 4'b0000 : 4'b0001;
													assign node4481 = (inp[1]) ? node4483 : 4'b0001;
														assign node4483 = (inp[2]) ? 4'b0000 : 4'b0001;
									assign node4486 = (inp[1]) ? node4540 : node4487;
										assign node4487 = (inp[7]) ? node4515 : node4488;
											assign node4488 = (inp[8]) ? node4502 : node4489;
												assign node4489 = (inp[14]) ? node4495 : node4490;
													assign node4490 = (inp[2]) ? 4'b0000 : node4491;
														assign node4491 = (inp[11]) ? 4'b0001 : 4'b0001;
													assign node4495 = (inp[11]) ? node4499 : node4496;
														assign node4496 = (inp[6]) ? 4'b0000 : 4'b1000;
														assign node4499 = (inp[6]) ? 4'b1000 : 4'b0000;
												assign node4502 = (inp[14]) ? node4508 : node4503;
													assign node4503 = (inp[11]) ? 4'b1000 : node4504;
														assign node4504 = (inp[6]) ? 4'b1001 : 4'b0001;
													assign node4508 = (inp[6]) ? node4512 : node4509;
														assign node4509 = (inp[11]) ? 4'b1001 : 4'b0001;
														assign node4512 = (inp[2]) ? 4'b1001 : 4'b0001;
											assign node4515 = (inp[8]) ? node4529 : node4516;
												assign node4516 = (inp[2]) ? node4524 : node4517;
													assign node4517 = (inp[13]) ? node4521 : node4518;
														assign node4518 = (inp[11]) ? 4'b1001 : 4'b1000;
														assign node4521 = (inp[6]) ? 4'b0001 : 4'b0000;
													assign node4524 = (inp[11]) ? 4'b0001 : node4525;
														assign node4525 = (inp[14]) ? 4'b0001 : 4'b0001;
												assign node4529 = (inp[14]) ? node4537 : node4530;
													assign node4530 = (inp[2]) ? node4534 : node4531;
														assign node4531 = (inp[11]) ? 4'b0001 : 4'b1001;
														assign node4534 = (inp[11]) ? 4'b0000 : 4'b0000;
													assign node4537 = (inp[2]) ? 4'b1000 : 4'b0000;
										assign node4540 = (inp[13]) ? node4560 : node4541;
											assign node4541 = (inp[6]) ? node4553 : node4542;
												assign node4542 = (inp[2]) ? node4548 : node4543;
													assign node4543 = (inp[14]) ? node4545 : 4'b0000;
														assign node4545 = (inp[11]) ? 4'b1001 : 4'b0001;
													assign node4548 = (inp[14]) ? 4'b1001 : node4549;
														assign node4549 = (inp[7]) ? 4'b1000 : 4'b1000;
												assign node4553 = (inp[11]) ? node4557 : node4554;
													assign node4554 = (inp[8]) ? 4'b1000 : 4'b0000;
													assign node4557 = (inp[8]) ? 4'b0001 : 4'b1000;
											assign node4560 = (inp[6]) ? node4568 : node4561;
												assign node4561 = (inp[11]) ? 4'b1000 : node4562;
													assign node4562 = (inp[8]) ? node4564 : 4'b0000;
														assign node4564 = (inp[7]) ? 4'b0000 : 4'b0001;
												assign node4568 = (inp[11]) ? node4574 : node4569;
													assign node4569 = (inp[14]) ? node4571 : 4'b1001;
														assign node4571 = (inp[7]) ? 4'b1001 : 4'b1000;
													assign node4574 = (inp[8]) ? 4'b0000 : node4575;
														assign node4575 = (inp[2]) ? 4'b0001 : 4'b0000;
							assign node4579 = (inp[10]) ? node4767 : node4580;
								assign node4580 = (inp[12]) ? node4678 : node4581;
									assign node4581 = (inp[1]) ? node4627 : node4582;
										assign node4582 = (inp[8]) ? node4604 : node4583;
											assign node4583 = (inp[7]) ? node4593 : node4584;
												assign node4584 = (inp[6]) ? node4588 : node4585;
													assign node4585 = (inp[11]) ? 4'b0000 : 4'b1000;
													assign node4588 = (inp[11]) ? 4'b1000 : node4589;
														assign node4589 = (inp[14]) ? 4'b0000 : 4'b0000;
												assign node4593 = (inp[2]) ? node4599 : node4594;
													assign node4594 = (inp[14]) ? 4'b0001 : node4595;
														assign node4595 = (inp[6]) ? 4'b1000 : 4'b0000;
													assign node4599 = (inp[11]) ? 4'b1001 : node4600;
														assign node4600 = (inp[13]) ? 4'b0001 : 4'b0001;
											assign node4604 = (inp[7]) ? node4616 : node4605;
												assign node4605 = (inp[2]) ? node4611 : node4606;
													assign node4606 = (inp[14]) ? 4'b1001 : node4607;
														assign node4607 = (inp[6]) ? 4'b1000 : 4'b0000;
													assign node4611 = (inp[11]) ? 4'b1001 : node4612;
														assign node4612 = (inp[6]) ? 4'b1001 : 4'b0001;
												assign node4616 = (inp[14]) ? node4622 : node4617;
													assign node4617 = (inp[2]) ? node4619 : 4'b0001;
														assign node4619 = (inp[6]) ? 4'b0000 : 4'b0000;
													assign node4622 = (inp[11]) ? node4624 : 4'b1000;
														assign node4624 = (inp[2]) ? 4'b1000 : 4'b0000;
										assign node4627 = (inp[7]) ? node4651 : node4628;
											assign node4628 = (inp[8]) ? node4642 : node4629;
												assign node4629 = (inp[13]) ? node4637 : node4630;
													assign node4630 = (inp[11]) ? node4634 : node4631;
														assign node4631 = (inp[6]) ? 4'b0000 : 4'b1000;
														assign node4634 = (inp[2]) ? 4'b1000 : 4'b1001;
													assign node4637 = (inp[2]) ? node4639 : 4'b0000;
														assign node4639 = (inp[11]) ? 4'b0000 : 4'b0000;
												assign node4642 = (inp[2]) ? node4646 : node4643;
													assign node4643 = (inp[14]) ? 4'b1001 : 4'b1000;
													assign node4646 = (inp[11]) ? 4'b0001 : node4647;
														assign node4647 = (inp[6]) ? 4'b1001 : 4'b0001;
											assign node4651 = (inp[8]) ? node4667 : node4652;
												assign node4652 = (inp[13]) ? node4660 : node4653;
													assign node4653 = (inp[11]) ? node4657 : node4654;
														assign node4654 = (inp[6]) ? 4'b1001 : 4'b0001;
														assign node4657 = (inp[6]) ? 4'b1000 : 4'b1001;
													assign node4660 = (inp[2]) ? node4664 : node4661;
														assign node4661 = (inp[14]) ? 4'b0001 : 4'b0000;
														assign node4664 = (inp[11]) ? 4'b0001 : 4'b1001;
												assign node4667 = (inp[6]) ? node4673 : node4668;
													assign node4668 = (inp[11]) ? node4670 : 4'b0001;
														assign node4670 = (inp[14]) ? 4'b1000 : 4'b1001;
													assign node4673 = (inp[2]) ? 4'b0000 : node4674;
														assign node4674 = (inp[14]) ? 4'b0000 : 4'b0001;
									assign node4678 = (inp[11]) ? node4722 : node4679;
										assign node4679 = (inp[6]) ? node4699 : node4680;
											assign node4680 = (inp[13]) ? node4692 : node4681;
												assign node4681 = (inp[1]) ? node4687 : node4682;
													assign node4682 = (inp[14]) ? 4'b1000 : node4683;
														assign node4683 = (inp[2]) ? 4'b1001 : 4'b1001;
													assign node4687 = (inp[8]) ? node4689 : 4'b1000;
														assign node4689 = (inp[2]) ? 4'b0000 : 4'b0000;
												assign node4692 = (inp[1]) ? node4694 : 4'b0001;
													assign node4694 = (inp[7]) ? node4696 : 4'b0000;
														assign node4696 = (inp[14]) ? 4'b0001 : 4'b0000;
											assign node4699 = (inp[13]) ? node4709 : node4700;
												assign node4700 = (inp[8]) ? node4706 : node4701;
													assign node4701 = (inp[1]) ? 4'b0000 : node4702;
														assign node4702 = (inp[7]) ? 4'b0000 : 4'b0001;
													assign node4706 = (inp[1]) ? 4'b1111 : 4'b0000;
												assign node4709 = (inp[1]) ? node4717 : node4710;
													assign node4710 = (inp[7]) ? node4714 : node4711;
														assign node4711 = (inp[14]) ? 4'b1111 : 4'b0000;
														assign node4714 = (inp[8]) ? 4'b1110 : 4'b1111;
													assign node4717 = (inp[8]) ? node4719 : 4'b1111;
														assign node4719 = (inp[14]) ? 4'b1110 : 4'b1111;
										assign node4722 = (inp[6]) ? node4744 : node4723;
											assign node4723 = (inp[1]) ? node4735 : node4724;
												assign node4724 = (inp[7]) ? node4728 : node4725;
													assign node4725 = (inp[8]) ? 4'b0001 : 4'b0000;
													assign node4728 = (inp[13]) ? node4732 : node4729;
														assign node4729 = (inp[14]) ? 4'b0001 : 4'b0000;
														assign node4732 = (inp[14]) ? 4'b1111 : 4'b1110;
												assign node4735 = (inp[8]) ? node4739 : node4736;
													assign node4736 = (inp[13]) ? 4'b1110 : 4'b0000;
													assign node4739 = (inp[7]) ? node4741 : 4'b1111;
														assign node4741 = (inp[14]) ? 4'b1110 : 4'b1110;
											assign node4744 = (inp[1]) ? node4756 : node4745;
												assign node4745 = (inp[7]) ? node4753 : node4746;
													assign node4746 = (inp[2]) ? node4750 : node4747;
														assign node4747 = (inp[8]) ? 4'b1110 : 4'b1110;
														assign node4750 = (inp[13]) ? 4'b0111 : 4'b1111;
													assign node4753 = (inp[2]) ? 4'b1111 : 4'b0111;
												assign node4756 = (inp[13]) ? node4762 : node4757;
													assign node4757 = (inp[8]) ? node4759 : 4'b1110;
														assign node4759 = (inp[7]) ? 4'b0110 : 4'b0111;
													assign node4762 = (inp[8]) ? 4'b0111 : node4763;
														assign node4763 = (inp[7]) ? 4'b0110 : 4'b0110;
								assign node4767 = (inp[12]) ? node4857 : node4768;
									assign node4768 = (inp[11]) ? node4814 : node4769;
										assign node4769 = (inp[6]) ? node4793 : node4770;
											assign node4770 = (inp[13]) ? node4782 : node4771;
												assign node4771 = (inp[1]) ? node4777 : node4772;
													assign node4772 = (inp[7]) ? node4774 : 4'b1001;
														assign node4774 = (inp[8]) ? 4'b1000 : 4'b1001;
													assign node4777 = (inp[8]) ? node4779 : 4'b1000;
														assign node4779 = (inp[14]) ? 4'b0000 : 4'b0001;
												assign node4782 = (inp[7]) ? node4786 : node4783;
													assign node4783 = (inp[1]) ? 4'b0000 : 4'b1000;
													assign node4786 = (inp[8]) ? node4790 : node4787;
														assign node4787 = (inp[2]) ? 4'b0001 : 4'b0000;
														assign node4790 = (inp[2]) ? 4'b0000 : 4'b0000;
											assign node4793 = (inp[1]) ? node4805 : node4794;
												assign node4794 = (inp[13]) ? node4800 : node4795;
													assign node4795 = (inp[8]) ? 4'b0000 : node4796;
														assign node4796 = (inp[14]) ? 4'b0001 : 4'b0000;
													assign node4800 = (inp[14]) ? 4'b1111 : node4801;
														assign node4801 = (inp[7]) ? 4'b1111 : 4'b0000;
												assign node4805 = (inp[7]) ? node4811 : node4806;
													assign node4806 = (inp[13]) ? node4808 : 4'b0000;
														assign node4808 = (inp[2]) ? 4'b1110 : 4'b1110;
													assign node4811 = (inp[8]) ? 4'b1110 : 4'b1111;
										assign node4814 = (inp[6]) ? node4840 : node4815;
											assign node4815 = (inp[1]) ? node4827 : node4816;
												assign node4816 = (inp[13]) ? node4820 : node4817;
													assign node4817 = (inp[14]) ? 4'b0000 : 4'b0001;
													assign node4820 = (inp[14]) ? node4824 : node4821;
														assign node4821 = (inp[7]) ? 4'b0000 : 4'b0000;
														assign node4824 = (inp[8]) ? 4'b1110 : 4'b1111;
												assign node4827 = (inp[7]) ? node4833 : node4828;
													assign node4828 = (inp[8]) ? 4'b1111 : node4829;
														assign node4829 = (inp[2]) ? 4'b1110 : 4'b1111;
													assign node4833 = (inp[14]) ? node4837 : node4834;
														assign node4834 = (inp[8]) ? 4'b1110 : 4'b0000;
														assign node4837 = (inp[8]) ? 4'b1110 : 4'b1111;
											assign node4840 = (inp[1]) ? node4850 : node4841;
												assign node4841 = (inp[13]) ? node4847 : node4842;
													assign node4842 = (inp[14]) ? 4'b1111 : node4843;
														assign node4843 = (inp[8]) ? 4'b1111 : 4'b1110;
													assign node4847 = (inp[2]) ? 4'b0110 : 4'b1110;
												assign node4850 = (inp[14]) ? node4852 : 4'b0111;
													assign node4852 = (inp[7]) ? node4854 : 4'b1110;
														assign node4854 = (inp[8]) ? 4'b0110 : 4'b0111;
									assign node4857 = (inp[2]) ? node4905 : node4858;
										assign node4858 = (inp[14]) ? node4882 : node4859;
											assign node4859 = (inp[6]) ? node4873 : node4860;
												assign node4860 = (inp[11]) ? node4868 : node4861;
													assign node4861 = (inp[1]) ? node4865 : node4862;
														assign node4862 = (inp[8]) ? 4'b1110 : 4'b1110;
														assign node4865 = (inp[13]) ? 4'b0111 : 4'b1110;
													assign node4868 = (inp[8]) ? 4'b0110 : node4869;
														assign node4869 = (inp[1]) ? 4'b1111 : 4'b0111;
												assign node4873 = (inp[13]) ? node4877 : node4874;
													assign node4874 = (inp[8]) ? 4'b0110 : 4'b1111;
													assign node4877 = (inp[1]) ? node4879 : 4'b1110;
														assign node4879 = (inp[8]) ? 4'b1111 : 4'b1110;
											assign node4882 = (inp[7]) ? node4892 : node4883;
												assign node4883 = (inp[8]) ? node4885 : 4'b1110;
													assign node4885 = (inp[11]) ? node4889 : node4886;
														assign node4886 = (inp[6]) ? 4'b1111 : 4'b0111;
														assign node4889 = (inp[6]) ? 4'b0111 : 4'b1111;
												assign node4892 = (inp[8]) ? node4898 : node4893;
													assign node4893 = (inp[13]) ? node4895 : 4'b1111;
														assign node4895 = (inp[11]) ? 4'b1111 : 4'b0111;
													assign node4898 = (inp[11]) ? node4902 : node4899;
														assign node4899 = (inp[1]) ? 4'b0110 : 4'b1110;
														assign node4902 = (inp[13]) ? 4'b0110 : 4'b0110;
										assign node4905 = (inp[1]) ? node4931 : node4906;
											assign node4906 = (inp[11]) ? node4916 : node4907;
												assign node4907 = (inp[6]) ? node4913 : node4908;
													assign node4908 = (inp[8]) ? node4910 : 4'b1110;
														assign node4910 = (inp[13]) ? 4'b0111 : 4'b1111;
													assign node4913 = (inp[7]) ? 4'b1110 : 4'b0110;
												assign node4916 = (inp[14]) ? node4924 : node4917;
													assign node4917 = (inp[6]) ? node4921 : node4918;
														assign node4918 = (inp[8]) ? 4'b0110 : 4'b0110;
														assign node4921 = (inp[13]) ? 4'b0110 : 4'b1110;
													assign node4924 = (inp[13]) ? node4928 : node4925;
														assign node4925 = (inp[6]) ? 4'b1111 : 4'b0110;
														assign node4928 = (inp[6]) ? 4'b0110 : 4'b1111;
											assign node4931 = (inp[13]) ? node4941 : node4932;
												assign node4932 = (inp[6]) ? 4'b0110 : node4933;
													assign node4933 = (inp[11]) ? node4937 : node4934;
														assign node4934 = (inp[8]) ? 4'b0110 : 4'b0111;
														assign node4937 = (inp[8]) ? 4'b1110 : 4'b0110;
												assign node4941 = (inp[6]) ? node4947 : node4942;
													assign node4942 = (inp[11]) ? 4'b1111 : node4943;
														assign node4943 = (inp[8]) ? 4'b0110 : 4'b0111;
													assign node4947 = (inp[11]) ? node4949 : 4'b1111;
														assign node4949 = (inp[8]) ? 4'b0111 : 4'b0110;
						assign node4952 = (inp[6]) ? node5296 : node4953;
							assign node4953 = (inp[9]) ? node5125 : node4954;
								assign node4954 = (inp[10]) ? node5040 : node4955;
									assign node4955 = (inp[12]) ? node5001 : node4956;
										assign node4956 = (inp[7]) ? node4978 : node4957;
											assign node4957 = (inp[11]) ? node4967 : node4958;
												assign node4958 = (inp[8]) ? node4964 : node4959;
													assign node4959 = (inp[14]) ? 4'b1110 : node4960;
														assign node4960 = (inp[2]) ? 4'b1110 : 4'b1111;
													assign node4964 = (inp[2]) ? 4'b0111 : 4'b1110;
												assign node4967 = (inp[8]) ? node4973 : node4968;
													assign node4968 = (inp[2]) ? node4970 : 4'b0111;
														assign node4970 = (inp[14]) ? 4'b0110 : 4'b0110;
													assign node4973 = (inp[14]) ? 4'b1111 : node4974;
														assign node4974 = (inp[1]) ? 4'b1110 : 4'b0110;
											assign node4978 = (inp[8]) ? node4992 : node4979;
												assign node4979 = (inp[14]) ? node4987 : node4980;
													assign node4980 = (inp[2]) ? node4984 : node4981;
														assign node4981 = (inp[13]) ? 4'b1110 : 4'b0110;
														assign node4984 = (inp[1]) ? 4'b0111 : 4'b1111;
													assign node4987 = (inp[11]) ? node4989 : 4'b0111;
														assign node4989 = (inp[1]) ? 4'b1111 : 4'b0111;
												assign node4992 = (inp[14]) ? node4996 : node4993;
													assign node4993 = (inp[11]) ? 4'b1111 : 4'b1110;
													assign node4996 = (inp[11]) ? node4998 : 4'b0110;
														assign node4998 = (inp[2]) ? 4'b0110 : 4'b1110;
										assign node5001 = (inp[11]) ? node5019 : node5002;
											assign node5002 = (inp[13]) ? node5012 : node5003;
												assign node5003 = (inp[7]) ? node5009 : node5004;
													assign node5004 = (inp[14]) ? node5006 : 4'b1110;
														assign node5006 = (inp[1]) ? 4'b1110 : 4'b1111;
													assign node5009 = (inp[2]) ? 4'b0111 : 4'b1110;
												assign node5012 = (inp[1]) ? 4'b0110 : node5013;
													assign node5013 = (inp[7]) ? 4'b0111 : node5014;
														assign node5014 = (inp[14]) ? 4'b0111 : 4'b1110;
											assign node5019 = (inp[13]) ? node5033 : node5020;
												assign node5020 = (inp[1]) ? node5026 : node5021;
													assign node5021 = (inp[8]) ? node5023 : 4'b0111;
														assign node5023 = (inp[2]) ? 4'b0110 : 4'b0110;
													assign node5026 = (inp[8]) ? node5030 : node5027;
														assign node5027 = (inp[7]) ? 4'b1011 : 4'b0110;
														assign node5030 = (inp[7]) ? 4'b1010 : 4'b1011;
												assign node5033 = (inp[7]) ? 4'b1010 : node5034;
													assign node5034 = (inp[2]) ? 4'b1011 : node5035;
														assign node5035 = (inp[1]) ? 4'b1011 : 4'b0110;
									assign node5040 = (inp[12]) ? node5086 : node5041;
										assign node5041 = (inp[11]) ? node5065 : node5042;
											assign node5042 = (inp[1]) ? node5054 : node5043;
												assign node5043 = (inp[13]) ? node5051 : node5044;
													assign node5044 = (inp[7]) ? node5048 : node5045;
														assign node5045 = (inp[8]) ? 4'b1111 : 4'b1110;
														assign node5048 = (inp[14]) ? 4'b1110 : 4'b1110;
													assign node5051 = (inp[8]) ? 4'b0110 : 4'b1110;
												assign node5054 = (inp[2]) ? node5060 : node5055;
													assign node5055 = (inp[14]) ? node5057 : 4'b1110;
														assign node5057 = (inp[13]) ? 4'b0111 : 4'b0110;
													assign node5060 = (inp[7]) ? 4'b0111 : node5061;
														assign node5061 = (inp[8]) ? 4'b0111 : 4'b1110;
											assign node5065 = (inp[1]) ? node5077 : node5066;
												assign node5066 = (inp[7]) ? node5072 : node5067;
													assign node5067 = (inp[13]) ? node5069 : 4'b0111;
														assign node5069 = (inp[8]) ? 4'b0010 : 4'b0110;
													assign node5072 = (inp[13]) ? node5074 : 4'b0110;
														assign node5074 = (inp[8]) ? 4'b1010 : 4'b1011;
												assign node5077 = (inp[8]) ? node5081 : node5078;
													assign node5078 = (inp[7]) ? 4'b1011 : 4'b1010;
													assign node5081 = (inp[7]) ? 4'b1010 : node5082;
														assign node5082 = (inp[2]) ? 4'b1011 : 4'b1010;
										assign node5086 = (inp[11]) ? node5108 : node5087;
											assign node5087 = (inp[2]) ? node5099 : node5088;
												assign node5088 = (inp[13]) ? node5094 : node5089;
													assign node5089 = (inp[14]) ? node5091 : 4'b1010;
														assign node5091 = (inp[7]) ? 4'b1011 : 4'b1010;
													assign node5094 = (inp[8]) ? 4'b0010 : node5095;
														assign node5095 = (inp[7]) ? 4'b0011 : 4'b1011;
												assign node5099 = (inp[7]) ? node5105 : node5100;
													assign node5100 = (inp[8]) ? 4'b0011 : node5101;
														assign node5101 = (inp[14]) ? 4'b0010 : 4'b1010;
													assign node5105 = (inp[8]) ? 4'b0010 : 4'b0011;
											assign node5108 = (inp[8]) ? node5114 : node5109;
												assign node5109 = (inp[1]) ? 4'b1011 : node5110;
													assign node5110 = (inp[13]) ? 4'b0010 : 4'b0011;
												assign node5114 = (inp[14]) ? node5122 : node5115;
													assign node5115 = (inp[2]) ? node5119 : node5116;
														assign node5116 = (inp[7]) ? 4'b1011 : 4'b0010;
														assign node5119 = (inp[7]) ? 4'b1010 : 4'b1011;
													assign node5122 = (inp[7]) ? 4'b1010 : 4'b1011;
								assign node5125 = (inp[10]) ? node5205 : node5126;
									assign node5126 = (inp[8]) ? node5162 : node5127;
										assign node5127 = (inp[7]) ? node5149 : node5128;
											assign node5128 = (inp[2]) ? node5140 : node5129;
												assign node5129 = (inp[14]) ? node5135 : node5130;
													assign node5130 = (inp[11]) ? 4'b0011 : node5131;
														assign node5131 = (inp[1]) ? 4'b0011 : 4'b1011;
													assign node5135 = (inp[13]) ? node5137 : 4'b1010;
														assign node5137 = (inp[11]) ? 4'b0010 : 4'b0010;
												assign node5140 = (inp[11]) ? node5146 : node5141;
													assign node5141 = (inp[1]) ? node5143 : 4'b1010;
														assign node5143 = (inp[13]) ? 4'b0010 : 4'b1010;
													assign node5146 = (inp[13]) ? 4'b1010 : 4'b0010;
											assign node5149 = (inp[2]) ? node5157 : node5150;
												assign node5150 = (inp[14]) ? node5152 : 4'b0010;
													assign node5152 = (inp[1]) ? 4'b0011 : node5153;
														assign node5153 = (inp[11]) ? 4'b0011 : 4'b1011;
												assign node5157 = (inp[11]) ? node5159 : 4'b0011;
													assign node5159 = (inp[12]) ? 4'b1111 : 4'b1011;
										assign node5162 = (inp[7]) ? node5186 : node5163;
											assign node5163 = (inp[14]) ? node5173 : node5164;
												assign node5164 = (inp[2]) ? node5168 : node5165;
													assign node5165 = (inp[11]) ? 4'b0010 : 4'b1010;
													assign node5168 = (inp[1]) ? node5170 : 4'b1011;
														assign node5170 = (inp[11]) ? 4'b1011 : 4'b0011;
												assign node5173 = (inp[11]) ? node5179 : node5174;
													assign node5174 = (inp[13]) ? 4'b0011 : node5175;
														assign node5175 = (inp[12]) ? 4'b1011 : 4'b0011;
													assign node5179 = (inp[1]) ? node5183 : node5180;
														assign node5180 = (inp[13]) ? 4'b1011 : 4'b0011;
														assign node5183 = (inp[12]) ? 4'b1111 : 4'b1011;
											assign node5186 = (inp[14]) ? node5198 : node5187;
												assign node5187 = (inp[2]) ? node5193 : node5188;
													assign node5188 = (inp[12]) ? 4'b0011 : node5189;
														assign node5189 = (inp[1]) ? 4'b0011 : 4'b1011;
													assign node5193 = (inp[1]) ? 4'b0010 : node5194;
														assign node5194 = (inp[11]) ? 4'b1110 : 4'b1010;
												assign node5198 = (inp[13]) ? node5200 : 4'b1010;
													assign node5200 = (inp[11]) ? node5202 : 4'b0010;
														assign node5202 = (inp[2]) ? 4'b1110 : 4'b1010;
									assign node5205 = (inp[12]) ? node5255 : node5206;
										assign node5206 = (inp[11]) ? node5228 : node5207;
											assign node5207 = (inp[7]) ? node5219 : node5208;
												assign node5208 = (inp[1]) ? node5214 : node5209;
													assign node5209 = (inp[2]) ? 4'b1010 : node5210;
														assign node5210 = (inp[8]) ? 4'b1010 : 4'b1011;
													assign node5214 = (inp[8]) ? node5216 : 4'b1010;
														assign node5216 = (inp[14]) ? 4'b0011 : 4'b0010;
												assign node5219 = (inp[8]) ? node5223 : node5220;
													assign node5220 = (inp[2]) ? 4'b0011 : 4'b0010;
													assign node5223 = (inp[2]) ? 4'b0010 : node5224;
														assign node5224 = (inp[13]) ? 4'b0010 : 4'b1010;
											assign node5228 = (inp[8]) ? node5242 : node5229;
												assign node5229 = (inp[1]) ? node5235 : node5230;
													assign node5230 = (inp[2]) ? 4'b0010 : node5231;
														assign node5231 = (inp[7]) ? 4'b0010 : 4'b0011;
													assign node5235 = (inp[13]) ? node5239 : node5236;
														assign node5236 = (inp[14]) ? 4'b0010 : 4'b0011;
														assign node5239 = (inp[14]) ? 4'b1110 : 4'b1111;
												assign node5242 = (inp[7]) ? node5248 : node5243;
													assign node5243 = (inp[2]) ? 4'b1111 : node5244;
														assign node5244 = (inp[13]) ? 4'b0010 : 4'b1111;
													assign node5248 = (inp[13]) ? node5252 : node5249;
														assign node5249 = (inp[1]) ? 4'b1110 : 4'b0010;
														assign node5252 = (inp[14]) ? 4'b1110 : 4'b1110;
										assign node5255 = (inp[2]) ? node5275 : node5256;
											assign node5256 = (inp[14]) ? node5266 : node5257;
												assign node5257 = (inp[8]) ? node5261 : node5258;
													assign node5258 = (inp[13]) ? 4'b0111 : 4'b0110;
													assign node5261 = (inp[7]) ? node5263 : 4'b1110;
														assign node5263 = (inp[11]) ? 4'b0111 : 4'b1111;
												assign node5266 = (inp[11]) ? 4'b0110 : node5267;
													assign node5267 = (inp[1]) ? node5271 : node5268;
														assign node5268 = (inp[7]) ? 4'b0111 : 4'b1110;
														assign node5271 = (inp[7]) ? 4'b0110 : 4'b0111;
											assign node5275 = (inp[13]) ? node5287 : node5276;
												assign node5276 = (inp[8]) ? node5280 : node5277;
													assign node5277 = (inp[11]) ? 4'b0110 : 4'b1110;
													assign node5280 = (inp[7]) ? node5284 : node5281;
														assign node5281 = (inp[11]) ? 4'b1111 : 4'b0111;
														assign node5284 = (inp[14]) ? 4'b0110 : 4'b1110;
												assign node5287 = (inp[11]) ? node5291 : node5288;
													assign node5288 = (inp[7]) ? 4'b0111 : 4'b0110;
													assign node5291 = (inp[7]) ? node5293 : 4'b1111;
														assign node5293 = (inp[8]) ? 4'b1110 : 4'b1111;
							assign node5296 = (inp[9]) ? node5474 : node5297;
								assign node5297 = (inp[12]) ? node5383 : node5298;
									assign node5298 = (inp[10]) ? node5348 : node5299;
										assign node5299 = (inp[13]) ? node5327 : node5300;
											assign node5300 = (inp[11]) ? node5314 : node5301;
												assign node5301 = (inp[8]) ? node5307 : node5302;
													assign node5302 = (inp[1]) ? node5304 : 4'b0111;
														assign node5304 = (inp[2]) ? 4'b0110 : 4'b0110;
													assign node5307 = (inp[1]) ? node5311 : node5308;
														assign node5308 = (inp[2]) ? 4'b0111 : 4'b0110;
														assign node5311 = (inp[14]) ? 4'b1110 : 4'b1111;
												assign node5314 = (inp[1]) ? node5322 : node5315;
													assign node5315 = (inp[14]) ? node5319 : node5316;
														assign node5316 = (inp[2]) ? 4'b1111 : 4'b1110;
														assign node5319 = (inp[2]) ? 4'b1110 : 4'b1110;
													assign node5322 = (inp[2]) ? 4'b0110 : node5323;
														assign node5323 = (inp[14]) ? 4'b0110 : 4'b1110;
											assign node5327 = (inp[11]) ? node5341 : node5328;
												assign node5328 = (inp[1]) ? node5336 : node5329;
													assign node5329 = (inp[7]) ? node5333 : node5330;
														assign node5330 = (inp[14]) ? 4'b0110 : 4'b0110;
														assign node5333 = (inp[2]) ? 4'b1110 : 4'b1111;
													assign node5336 = (inp[14]) ? 4'b1111 : node5337;
														assign node5337 = (inp[8]) ? 4'b1110 : 4'b1110;
												assign node5341 = (inp[8]) ? node5343 : 4'b0111;
													assign node5343 = (inp[14]) ? 4'b0110 : node5344;
														assign node5344 = (inp[7]) ? 4'b0111 : 4'b0110;
										assign node5348 = (inp[13]) ? node5370 : node5349;
											assign node5349 = (inp[11]) ? node5361 : node5350;
												assign node5350 = (inp[7]) ? node5356 : node5351;
													assign node5351 = (inp[8]) ? 4'b0111 : node5352;
														assign node5352 = (inp[2]) ? 4'b0110 : 4'b0110;
													assign node5356 = (inp[1]) ? node5358 : 4'b0110;
														assign node5358 = (inp[14]) ? 4'b1011 : 4'b0110;
												assign node5361 = (inp[1]) ? node5365 : node5362;
													assign node5362 = (inp[8]) ? 4'b1010 : 4'b1011;
													assign node5365 = (inp[2]) ? 4'b0010 : node5366;
														assign node5366 = (inp[8]) ? 4'b0011 : 4'b0011;
											assign node5370 = (inp[11]) ? node5378 : node5371;
												assign node5371 = (inp[1]) ? node5373 : 4'b1011;
													assign node5373 = (inp[8]) ? node5375 : 4'b1010;
														assign node5375 = (inp[7]) ? 4'b1010 : 4'b1011;
												assign node5378 = (inp[2]) ? 4'b0010 : node5379;
													assign node5379 = (inp[14]) ? 4'b0011 : 4'b1010;
									assign node5383 = (inp[11]) ? node5431 : node5384;
										assign node5384 = (inp[13]) ? node5408 : node5385;
											assign node5385 = (inp[10]) ? node5399 : node5386;
												assign node5386 = (inp[7]) ? node5394 : node5387;
													assign node5387 = (inp[8]) ? node5391 : node5388;
														assign node5388 = (inp[2]) ? 4'b0110 : 4'b0110;
														assign node5391 = (inp[2]) ? 4'b1011 : 4'b0110;
													assign node5394 = (inp[1]) ? node5396 : 4'b0111;
														assign node5396 = (inp[2]) ? 4'b1011 : 4'b0010;
												assign node5399 = (inp[8]) ? node5405 : node5400;
													assign node5400 = (inp[14]) ? 4'b1011 : node5401;
														assign node5401 = (inp[2]) ? 4'b0010 : 4'b0010;
													assign node5405 = (inp[1]) ? 4'b1011 : 4'b0011;
											assign node5408 = (inp[1]) ? node5418 : node5409;
												assign node5409 = (inp[10]) ? node5411 : 4'b0111;
													assign node5411 = (inp[7]) ? node5415 : node5412;
														assign node5412 = (inp[8]) ? 4'b1011 : 4'b0010;
														assign node5415 = (inp[2]) ? 4'b1010 : 4'b1011;
												assign node5418 = (inp[2]) ? node5426 : node5419;
													assign node5419 = (inp[8]) ? node5423 : node5420;
														assign node5420 = (inp[7]) ? 4'b1011 : 4'b1010;
														assign node5423 = (inp[10]) ? 4'b1010 : 4'b1010;
													assign node5426 = (inp[7]) ? node5428 : 4'b1011;
														assign node5428 = (inp[8]) ? 4'b1010 : 4'b1011;
										assign node5431 = (inp[1]) ? node5459 : node5432;
											assign node5432 = (inp[13]) ? node5448 : node5433;
												assign node5433 = (inp[2]) ? node5441 : node5434;
													assign node5434 = (inp[14]) ? node5438 : node5435;
														assign node5435 = (inp[8]) ? 4'b1010 : 4'b1010;
														assign node5438 = (inp[10]) ? 4'b1011 : 4'b1010;
													assign node5441 = (inp[8]) ? node5445 : node5442;
														assign node5442 = (inp[7]) ? 4'b1011 : 4'b1010;
														assign node5445 = (inp[7]) ? 4'b1010 : 4'b1011;
												assign node5448 = (inp[14]) ? node5454 : node5449;
													assign node5449 = (inp[8]) ? node5451 : 4'b1010;
														assign node5451 = (inp[7]) ? 4'b0010 : 4'b1010;
													assign node5454 = (inp[8]) ? 4'b0011 : node5455;
														assign node5455 = (inp[7]) ? 4'b0011 : 4'b1010;
											assign node5459 = (inp[14]) ? node5469 : node5460;
												assign node5460 = (inp[8]) ? node5464 : node5461;
													assign node5461 = (inp[13]) ? 4'b0010 : 4'b1010;
													assign node5464 = (inp[10]) ? 4'b0010 : node5465;
														assign node5465 = (inp[13]) ? 4'b0010 : 4'b0010;
												assign node5469 = (inp[7]) ? node5471 : 4'b0011;
													assign node5471 = (inp[8]) ? 4'b0010 : 4'b0011;
								assign node5474 = (inp[12]) ? node5570 : node5475;
									assign node5475 = (inp[10]) ? node5525 : node5476;
										assign node5476 = (inp[11]) ? node5502 : node5477;
											assign node5477 = (inp[1]) ? node5489 : node5478;
												assign node5478 = (inp[13]) ? node5484 : node5479;
													assign node5479 = (inp[2]) ? node5481 : 4'b0010;
														assign node5481 = (inp[14]) ? 4'b0011 : 4'b0010;
													assign node5484 = (inp[7]) ? node5486 : 4'b0010;
														assign node5486 = (inp[14]) ? 4'b1010 : 4'b1011;
												assign node5489 = (inp[13]) ? node5497 : node5490;
													assign node5490 = (inp[8]) ? node5494 : node5491;
														assign node5491 = (inp[7]) ? 4'b1011 : 4'b0010;
														assign node5494 = (inp[7]) ? 4'b1010 : 4'b1011;
													assign node5497 = (inp[14]) ? 4'b1011 : node5498;
														assign node5498 = (inp[7]) ? 4'b1011 : 4'b1010;
											assign node5502 = (inp[13]) ? node5514 : node5503;
												assign node5503 = (inp[8]) ? node5509 : node5504;
													assign node5504 = (inp[1]) ? node5506 : 4'b1011;
														assign node5506 = (inp[14]) ? 4'b1010 : 4'b1011;
													assign node5509 = (inp[1]) ? node5511 : 4'b1010;
														assign node5511 = (inp[14]) ? 4'b0011 : 4'b0010;
												assign node5514 = (inp[7]) ? node5520 : node5515;
													assign node5515 = (inp[2]) ? 4'b1010 : node5516;
														assign node5516 = (inp[1]) ? 4'b0010 : 4'b0011;
													assign node5520 = (inp[8]) ? node5522 : 4'b0011;
														assign node5522 = (inp[14]) ? 4'b0010 : 4'b0011;
										assign node5525 = (inp[11]) ? node5549 : node5526;
											assign node5526 = (inp[13]) ? node5538 : node5527;
												assign node5527 = (inp[8]) ? node5533 : node5528;
													assign node5528 = (inp[2]) ? node5530 : 4'b0010;
														assign node5530 = (inp[7]) ? 4'b0011 : 4'b0010;
													assign node5533 = (inp[7]) ? node5535 : 4'b1111;
														assign node5535 = (inp[2]) ? 4'b0010 : 4'b0011;
												assign node5538 = (inp[1]) ? node5544 : node5539;
													assign node5539 = (inp[7]) ? node5541 : 4'b0010;
														assign node5541 = (inp[2]) ? 4'b1111 : 4'b0010;
													assign node5544 = (inp[14]) ? node5546 : 4'b1110;
														assign node5546 = (inp[8]) ? 4'b1110 : 4'b1111;
											assign node5549 = (inp[13]) ? node5559 : node5550;
												assign node5550 = (inp[1]) ? node5556 : node5551;
													assign node5551 = (inp[8]) ? 4'b1110 : node5552;
														assign node5552 = (inp[7]) ? 4'b1111 : 4'b1110;
													assign node5556 = (inp[8]) ? 4'b0111 : 4'b1110;
												assign node5559 = (inp[1]) ? node5565 : node5560;
													assign node5560 = (inp[7]) ? node5562 : 4'b1110;
														assign node5562 = (inp[8]) ? 4'b0110 : 4'b0111;
													assign node5565 = (inp[8]) ? node5567 : 4'b0110;
														assign node5567 = (inp[7]) ? 4'b0110 : 4'b0111;
									assign node5570 = (inp[11]) ? node5614 : node5571;
										assign node5571 = (inp[1]) ? node5595 : node5572;
											assign node5572 = (inp[10]) ? node5584 : node5573;
												assign node5573 = (inp[14]) ? node5579 : node5574;
													assign node5574 = (inp[2]) ? 4'b0011 : node5575;
														assign node5575 = (inp[13]) ? 4'b0010 : 4'b0010;
													assign node5579 = (inp[13]) ? node5581 : 4'b0010;
														assign node5581 = (inp[7]) ? 4'b1110 : 4'b1111;
												assign node5584 = (inp[13]) ? node5588 : node5585;
													assign node5585 = (inp[2]) ? 4'b0110 : 4'b0111;
													assign node5588 = (inp[7]) ? node5592 : node5589;
														assign node5589 = (inp[8]) ? 4'b1111 : 4'b0110;
														assign node5592 = (inp[8]) ? 4'b1110 : 4'b1111;
											assign node5595 = (inp[7]) ? node5607 : node5596;
												assign node5596 = (inp[13]) ? node5604 : node5597;
													assign node5597 = (inp[8]) ? node5601 : node5598;
														assign node5598 = (inp[14]) ? 4'b0010 : 4'b0011;
														assign node5601 = (inp[14]) ? 4'b1111 : 4'b0010;
													assign node5604 = (inp[10]) ? 4'b1111 : 4'b1110;
												assign node5607 = (inp[8]) ? node5609 : 4'b1111;
													assign node5609 = (inp[2]) ? 4'b1110 : node5610;
														assign node5610 = (inp[14]) ? 4'b1110 : 4'b1111;
										assign node5614 = (inp[13]) ? node5636 : node5615;
											assign node5615 = (inp[1]) ? node5625 : node5616;
												assign node5616 = (inp[10]) ? node5620 : node5617;
													assign node5617 = (inp[7]) ? 4'b1110 : 4'b1111;
													assign node5620 = (inp[14]) ? 4'b1110 : node5621;
														assign node5621 = (inp[7]) ? 4'b1111 : 4'b1110;
												assign node5625 = (inp[7]) ? node5633 : node5626;
													assign node5626 = (inp[14]) ? node5630 : node5627;
														assign node5627 = (inp[10]) ? 4'b1111 : 4'b1110;
														assign node5630 = (inp[8]) ? 4'b0111 : 4'b1110;
													assign node5633 = (inp[8]) ? 4'b0110 : 4'b0111;
											assign node5636 = (inp[14]) ? node5648 : node5637;
												assign node5637 = (inp[1]) ? node5641 : node5638;
													assign node5638 = (inp[10]) ? 4'b0111 : 4'b1110;
													assign node5641 = (inp[2]) ? node5645 : node5642;
														assign node5642 = (inp[8]) ? 4'b0111 : 4'b0110;
														assign node5645 = (inp[7]) ? 4'b0110 : 4'b0110;
												assign node5648 = (inp[8]) ? node5650 : 4'b0111;
													assign node5650 = (inp[7]) ? 4'b0110 : 4'b0111;
			assign node5653 = (inp[15]) ? node8477 : node5654;
				assign node5654 = (inp[3]) ? node7070 : node5655;
					assign node5655 = (inp[5]) ? node6357 : node5656;
						assign node5656 = (inp[10]) ? node6012 : node5657;
							assign node5657 = (inp[9]) ? node5831 : node5658;
								assign node5658 = (inp[12]) ? node5744 : node5659;
									assign node5659 = (inp[13]) ? node5707 : node5660;
										assign node5660 = (inp[1]) ? node5690 : node5661;
											assign node5661 = (inp[7]) ? node5677 : node5662;
												assign node5662 = (inp[8]) ? node5670 : node5663;
													assign node5663 = (inp[2]) ? node5667 : node5664;
														assign node5664 = (inp[6]) ? 4'b1010 : 4'b0011;
														assign node5667 = (inp[14]) ? 4'b0010 : 4'b1010;
													assign node5670 = (inp[2]) ? node5674 : node5671;
														assign node5671 = (inp[14]) ? 4'b0011 : 4'b0010;
														assign node5674 = (inp[14]) ? 4'b1011 : 4'b0011;
												assign node5677 = (inp[8]) ? node5685 : node5678;
													assign node5678 = (inp[14]) ? node5682 : node5679;
														assign node5679 = (inp[2]) ? 4'b0011 : 4'b0010;
														assign node5682 = (inp[2]) ? 4'b1011 : 4'b0011;
													assign node5685 = (inp[11]) ? node5687 : 4'b1010;
														assign node5687 = (inp[2]) ? 4'b0010 : 4'b0011;
											assign node5690 = (inp[7]) ? node5704 : node5691;
												assign node5691 = (inp[6]) ? node5699 : node5692;
													assign node5692 = (inp[14]) ? node5696 : node5693;
														assign node5693 = (inp[11]) ? 4'b0010 : 4'b1011;
														assign node5696 = (inp[8]) ? 4'b1011 : 4'b0010;
													assign node5699 = (inp[2]) ? node5701 : 4'b1010;
														assign node5701 = (inp[8]) ? 4'b0011 : 4'b0010;
												assign node5704 = (inp[8]) ? 4'b1010 : 4'b1011;
										assign node5707 = (inp[11]) ? node5725 : node5708;
											assign node5708 = (inp[6]) ? node5716 : node5709;
												assign node5709 = (inp[2]) ? 4'b0011 : node5710;
													assign node5710 = (inp[8]) ? node5712 : 4'b0011;
														assign node5712 = (inp[14]) ? 4'b0010 : 4'b0011;
												assign node5716 = (inp[14]) ? node5722 : node5717;
													assign node5717 = (inp[1]) ? node5719 : 4'b1011;
														assign node5719 = (inp[2]) ? 4'b1010 : 4'b1011;
													assign node5722 = (inp[1]) ? 4'b1011 : 4'b0010;
											assign node5725 = (inp[6]) ? node5735 : node5726;
												assign node5726 = (inp[14]) ? 4'b1011 : node5727;
													assign node5727 = (inp[7]) ? node5731 : node5728;
														assign node5728 = (inp[2]) ? 4'b0010 : 4'b0010;
														assign node5731 = (inp[1]) ? 4'b1010 : 4'b1011;
												assign node5735 = (inp[8]) ? 4'b0011 : node5736;
													assign node5736 = (inp[1]) ? node5740 : node5737;
														assign node5737 = (inp[7]) ? 4'b1010 : 4'b1011;
														assign node5740 = (inp[7]) ? 4'b0011 : 4'b0010;
									assign node5744 = (inp[6]) ? node5792 : node5745;
										assign node5745 = (inp[11]) ? node5769 : node5746;
											assign node5746 = (inp[1]) ? node5756 : node5747;
												assign node5747 = (inp[14]) ? node5753 : node5748;
													assign node5748 = (inp[2]) ? 4'b0010 : node5749;
														assign node5749 = (inp[8]) ? 4'b1010 : 4'b1011;
													assign node5753 = (inp[13]) ? 4'b0011 : 4'b1010;
												assign node5756 = (inp[7]) ? node5764 : node5757;
													assign node5757 = (inp[13]) ? node5761 : node5758;
														assign node5758 = (inp[14]) ? 4'b0010 : 4'b1010;
														assign node5761 = (inp[2]) ? 4'b0011 : 4'b0010;
													assign node5764 = (inp[8]) ? 4'b0010 : node5765;
														assign node5765 = (inp[13]) ? 4'b0010 : 4'b0011;
											assign node5769 = (inp[1]) ? node5781 : node5770;
												assign node5770 = (inp[13]) ? node5776 : node5771;
													assign node5771 = (inp[7]) ? node5773 : 4'b0011;
														assign node5773 = (inp[8]) ? 4'b0011 : 4'b0011;
													assign node5776 = (inp[7]) ? 4'b1111 : node5777;
														assign node5777 = (inp[2]) ? 4'b0010 : 4'b0010;
												assign node5781 = (inp[7]) ? node5785 : node5782;
													assign node5782 = (inp[13]) ? 4'b1110 : 4'b0010;
													assign node5785 = (inp[8]) ? node5789 : node5786;
														assign node5786 = (inp[14]) ? 4'b1111 : 4'b1110;
														assign node5789 = (inp[2]) ? 4'b1110 : 4'b1111;
										assign node5792 = (inp[11]) ? node5814 : node5793;
											assign node5793 = (inp[1]) ? node5803 : node5794;
												assign node5794 = (inp[13]) ? node5800 : node5795;
													assign node5795 = (inp[7]) ? node5797 : 4'b0010;
														assign node5797 = (inp[8]) ? 4'b0010 : 4'b0011;
													assign node5800 = (inp[8]) ? 4'b1110 : 4'b1111;
												assign node5803 = (inp[7]) ? node5809 : node5804;
													assign node5804 = (inp[14]) ? 4'b1111 : node5805;
														assign node5805 = (inp[13]) ? 4'b1110 : 4'b0010;
													assign node5809 = (inp[8]) ? 4'b1110 : node5810;
														assign node5810 = (inp[13]) ? 4'b1110 : 4'b1111;
											assign node5814 = (inp[14]) ? node5826 : node5815;
												assign node5815 = (inp[1]) ? node5819 : node5816;
													assign node5816 = (inp[13]) ? 4'b1110 : 4'b1111;
													assign node5819 = (inp[2]) ? node5823 : node5820;
														assign node5820 = (inp[8]) ? 4'b0111 : 4'b0110;
														assign node5823 = (inp[7]) ? 4'b0110 : 4'b1110;
												assign node5826 = (inp[7]) ? 4'b0111 : node5827;
													assign node5827 = (inp[8]) ? 4'b0111 : 4'b1110;
								assign node5831 = (inp[12]) ? node5923 : node5832;
									assign node5832 = (inp[1]) ? node5888 : node5833;
										assign node5833 = (inp[14]) ? node5863 : node5834;
											assign node5834 = (inp[2]) ? node5850 : node5835;
												assign node5835 = (inp[7]) ? node5843 : node5836;
													assign node5836 = (inp[8]) ? node5840 : node5837;
														assign node5837 = (inp[6]) ? 4'b0111 : 4'b1111;
														assign node5840 = (inp[13]) ? 4'b1110 : 4'b0110;
													assign node5843 = (inp[8]) ? node5847 : node5844;
														assign node5844 = (inp[11]) ? 4'b0110 : 4'b0110;
														assign node5847 = (inp[6]) ? 4'b1111 : 4'b0111;
												assign node5850 = (inp[6]) ? node5856 : node5851;
													assign node5851 = (inp[8]) ? 4'b0111 : node5852;
														assign node5852 = (inp[11]) ? 4'b0111 : 4'b1111;
													assign node5856 = (inp[11]) ? node5860 : node5857;
														assign node5857 = (inp[13]) ? 4'b1110 : 4'b0110;
														assign node5860 = (inp[7]) ? 4'b0111 : 4'b1110;
											assign node5863 = (inp[2]) ? node5875 : node5864;
												assign node5864 = (inp[7]) ? node5868 : node5865;
													assign node5865 = (inp[8]) ? 4'b0111 : 4'b0110;
													assign node5868 = (inp[8]) ? node5872 : node5869;
														assign node5869 = (inp[6]) ? 4'b1111 : 4'b0111;
														assign node5872 = (inp[13]) ? 4'b0110 : 4'b0110;
												assign node5875 = (inp[6]) ? node5881 : node5876;
													assign node5876 = (inp[11]) ? node5878 : 4'b1110;
														assign node5878 = (inp[7]) ? 4'b0110 : 4'b0110;
													assign node5881 = (inp[8]) ? node5885 : node5882;
														assign node5882 = (inp[7]) ? 4'b0111 : 4'b0110;
														assign node5885 = (inp[7]) ? 4'b1110 : 4'b0111;
										assign node5888 = (inp[8]) ? node5910 : node5889;
											assign node5889 = (inp[7]) ? node5901 : node5890;
												assign node5890 = (inp[6]) ? node5896 : node5891;
													assign node5891 = (inp[13]) ? 4'b0110 : node5892;
														assign node5892 = (inp[11]) ? 4'b0110 : 4'b1110;
													assign node5896 = (inp[2]) ? node5898 : 4'b1110;
														assign node5898 = (inp[11]) ? 4'b1110 : 4'b0110;
												assign node5901 = (inp[2]) ? node5907 : node5902;
													assign node5902 = (inp[13]) ? 4'b1110 : node5903;
														assign node5903 = (inp[14]) ? 4'b0111 : 4'b0110;
													assign node5907 = (inp[11]) ? 4'b0111 : 4'b1111;
											assign node5910 = (inp[6]) ? node5914 : node5911;
												assign node5911 = (inp[11]) ? 4'b1111 : 4'b0111;
												assign node5914 = (inp[11]) ? node5920 : node5915;
													assign node5915 = (inp[13]) ? node5917 : 4'b1111;
														assign node5917 = (inp[7]) ? 4'b1110 : 4'b1110;
													assign node5920 = (inp[7]) ? 4'b0110 : 4'b0111;
									assign node5923 = (inp[6]) ? node5965 : node5924;
										assign node5924 = (inp[11]) ? node5948 : node5925;
											assign node5925 = (inp[1]) ? node5935 : node5926;
												assign node5926 = (inp[13]) ? node5932 : node5927;
													assign node5927 = (inp[7]) ? node5929 : 4'b1110;
														assign node5929 = (inp[8]) ? 4'b1110 : 4'b1111;
													assign node5932 = (inp[8]) ? 4'b0110 : 4'b1110;
												assign node5935 = (inp[7]) ? node5943 : node5936;
													assign node5936 = (inp[8]) ? node5940 : node5937;
														assign node5937 = (inp[13]) ? 4'b0110 : 4'b1110;
														assign node5940 = (inp[2]) ? 4'b0111 : 4'b0110;
													assign node5943 = (inp[13]) ? 4'b0110 : node5944;
														assign node5944 = (inp[8]) ? 4'b0110 : 4'b0111;
											assign node5948 = (inp[1]) ? node5956 : node5949;
												assign node5949 = (inp[7]) ? node5951 : 4'b0110;
													assign node5951 = (inp[13]) ? 4'b1011 : node5952;
														assign node5952 = (inp[2]) ? 4'b0110 : 4'b0111;
												assign node5956 = (inp[7]) ? node5958 : 4'b1010;
													assign node5958 = (inp[13]) ? node5962 : node5959;
														assign node5959 = (inp[8]) ? 4'b1011 : 4'b0110;
														assign node5962 = (inp[14]) ? 4'b1010 : 4'b1011;
										assign node5965 = (inp[11]) ? node5993 : node5966;
											assign node5966 = (inp[1]) ? node5980 : node5967;
												assign node5967 = (inp[13]) ? node5973 : node5968;
													assign node5968 = (inp[2]) ? 4'b0111 : node5969;
														assign node5969 = (inp[7]) ? 4'b0110 : 4'b0111;
													assign node5973 = (inp[2]) ? node5977 : node5974;
														assign node5974 = (inp[14]) ? 4'b0110 : 4'b0110;
														assign node5977 = (inp[7]) ? 4'b1010 : 4'b0110;
												assign node5980 = (inp[13]) ? node5986 : node5981;
													assign node5981 = (inp[8]) ? 4'b1011 : node5982;
														assign node5982 = (inp[2]) ? 4'b0110 : 4'b0111;
													assign node5986 = (inp[14]) ? node5990 : node5987;
														assign node5987 = (inp[2]) ? 4'b1010 : 4'b1011;
														assign node5990 = (inp[7]) ? 4'b1011 : 4'b1010;
											assign node5993 = (inp[13]) ? node6001 : node5994;
												assign node5994 = (inp[1]) ? node5996 : 4'b1011;
													assign node5996 = (inp[14]) ? 4'b0011 : node5997;
														assign node5997 = (inp[2]) ? 4'b0011 : 4'b1010;
												assign node6001 = (inp[1]) ? node6007 : node6002;
													assign node6002 = (inp[14]) ? node6004 : 4'b0011;
														assign node6004 = (inp[7]) ? 4'b0010 : 4'b0011;
													assign node6007 = (inp[8]) ? 4'b0010 : node6008;
														assign node6008 = (inp[7]) ? 4'b0010 : 4'b0010;
							assign node6012 = (inp[9]) ? node6170 : node6013;
								assign node6013 = (inp[12]) ? node6097 : node6014;
									assign node6014 = (inp[6]) ? node6054 : node6015;
										assign node6015 = (inp[11]) ? node6031 : node6016;
											assign node6016 = (inp[13]) ? node6026 : node6017;
												assign node6017 = (inp[1]) ? node6019 : 4'b1011;
													assign node6019 = (inp[7]) ? node6023 : node6020;
														assign node6020 = (inp[2]) ? 4'b1010 : 4'b1010;
														assign node6023 = (inp[8]) ? 4'b0010 : 4'b1010;
												assign node6026 = (inp[1]) ? 4'b0010 : node6027;
													assign node6027 = (inp[8]) ? 4'b0010 : 4'b1010;
											assign node6031 = (inp[7]) ? node6043 : node6032;
												assign node6032 = (inp[8]) ? node6038 : node6033;
													assign node6033 = (inp[2]) ? 4'b0010 : node6034;
														assign node6034 = (inp[14]) ? 4'b0010 : 4'b0011;
													assign node6038 = (inp[13]) ? node6040 : 4'b0011;
														assign node6040 = (inp[14]) ? 4'b1111 : 4'b0010;
												assign node6043 = (inp[8]) ? node6049 : node6044;
													assign node6044 = (inp[13]) ? node6046 : 4'b0011;
														assign node6046 = (inp[14]) ? 4'b1111 : 4'b1110;
													assign node6049 = (inp[14]) ? 4'b1110 : node6050;
														assign node6050 = (inp[2]) ? 4'b1110 : 4'b1111;
										assign node6054 = (inp[11]) ? node6076 : node6055;
											assign node6055 = (inp[13]) ? node6065 : node6056;
												assign node6056 = (inp[1]) ? node6062 : node6057;
													assign node6057 = (inp[8]) ? node6059 : 4'b0011;
														assign node6059 = (inp[14]) ? 4'b0010 : 4'b0010;
													assign node6062 = (inp[14]) ? 4'b1111 : 4'b0010;
												assign node6065 = (inp[14]) ? node6071 : node6066;
													assign node6066 = (inp[7]) ? 4'b1111 : node6067;
														assign node6067 = (inp[1]) ? 4'b1111 : 4'b0011;
													assign node6071 = (inp[8]) ? 4'b1110 : node6072;
														assign node6072 = (inp[7]) ? 4'b1111 : 4'b1110;
											assign node6076 = (inp[13]) ? node6086 : node6077;
												assign node6077 = (inp[8]) ? node6083 : node6078;
													assign node6078 = (inp[14]) ? 4'b1110 : node6079;
														assign node6079 = (inp[2]) ? 4'b1111 : 4'b1110;
													assign node6083 = (inp[1]) ? 4'b0110 : 4'b1110;
												assign node6086 = (inp[1]) ? node6092 : node6087;
													assign node6087 = (inp[7]) ? node6089 : 4'b0111;
														assign node6089 = (inp[2]) ? 4'b0110 : 4'b0111;
													assign node6092 = (inp[8]) ? node6094 : 4'b0110;
														assign node6094 = (inp[7]) ? 4'b0110 : 4'b0110;
									assign node6097 = (inp[8]) ? node6133 : node6098;
										assign node6098 = (inp[7]) ? node6116 : node6099;
											assign node6099 = (inp[11]) ? node6105 : node6100;
												assign node6100 = (inp[6]) ? 4'b0110 : node6101;
													assign node6101 = (inp[14]) ? 4'b1110 : 4'b0110;
												assign node6105 = (inp[2]) ? node6111 : node6106;
													assign node6106 = (inp[6]) ? node6108 : 4'b0111;
														assign node6108 = (inp[14]) ? 4'b1110 : 4'b1111;
													assign node6111 = (inp[13]) ? 4'b1110 : node6112;
														assign node6112 = (inp[1]) ? 4'b0110 : 4'b1110;
											assign node6116 = (inp[2]) ? node6128 : node6117;
												assign node6117 = (inp[14]) ? node6123 : node6118;
													assign node6118 = (inp[11]) ? 4'b0110 : node6119;
														assign node6119 = (inp[13]) ? 4'b1110 : 4'b0110;
													assign node6123 = (inp[13]) ? 4'b0111 : node6124;
														assign node6124 = (inp[1]) ? 4'b0111 : 4'b0111;
												assign node6128 = (inp[1]) ? 4'b0111 : node6129;
													assign node6129 = (inp[11]) ? 4'b0111 : 4'b1111;
										assign node6133 = (inp[7]) ? node6151 : node6134;
											assign node6134 = (inp[14]) ? node6142 : node6135;
												assign node6135 = (inp[2]) ? node6139 : node6136;
													assign node6136 = (inp[1]) ? 4'b0110 : 4'b1110;
													assign node6139 = (inp[6]) ? 4'b0111 : 4'b1111;
												assign node6142 = (inp[13]) ? node6148 : node6143;
													assign node6143 = (inp[2]) ? node6145 : 4'b1111;
														assign node6145 = (inp[1]) ? 4'b0111 : 4'b0111;
													assign node6148 = (inp[11]) ? 4'b0111 : 4'b1111;
											assign node6151 = (inp[2]) ? node6159 : node6152;
												assign node6152 = (inp[14]) ? node6154 : 4'b1111;
													assign node6154 = (inp[11]) ? node6156 : 4'b1110;
														assign node6156 = (inp[6]) ? 4'b0110 : 4'b1110;
												assign node6159 = (inp[1]) ? node6165 : node6160;
													assign node6160 = (inp[6]) ? node6162 : 4'b1110;
														assign node6162 = (inp[11]) ? 4'b1110 : 4'b0110;
													assign node6165 = (inp[11]) ? 4'b0110 : node6166;
														assign node6166 = (inp[6]) ? 4'b1110 : 4'b0110;
								assign node6170 = (inp[12]) ? node6260 : node6171;
									assign node6171 = (inp[11]) ? node6213 : node6172;
										assign node6172 = (inp[6]) ? node6194 : node6173;
											assign node6173 = (inp[1]) ? node6183 : node6174;
												assign node6174 = (inp[7]) ? node6180 : node6175;
													assign node6175 = (inp[13]) ? 4'b1110 : node6176;
														assign node6176 = (inp[14]) ? 4'b1110 : 4'b1110;
													assign node6180 = (inp[13]) ? 4'b0111 : 4'b1111;
												assign node6183 = (inp[8]) ? node6189 : node6184;
													assign node6184 = (inp[13]) ? node6186 : 4'b1111;
														assign node6186 = (inp[2]) ? 4'b0110 : 4'b0111;
													assign node6189 = (inp[2]) ? 4'b0110 : node6190;
														assign node6190 = (inp[14]) ? 4'b0110 : 4'b0111;
											assign node6194 = (inp[13]) ? node6204 : node6195;
												assign node6195 = (inp[8]) ? node6201 : node6196;
													assign node6196 = (inp[1]) ? node6198 : 4'b0111;
														assign node6198 = (inp[14]) ? 4'b0110 : 4'b0110;
													assign node6201 = (inp[2]) ? 4'b1010 : 4'b0110;
												assign node6204 = (inp[1]) ? node6208 : node6205;
													assign node6205 = (inp[7]) ? 4'b1010 : 4'b0110;
													assign node6208 = (inp[14]) ? node6210 : 4'b1011;
														assign node6210 = (inp[2]) ? 4'b1011 : 4'b1010;
										assign node6213 = (inp[6]) ? node6239 : node6214;
											assign node6214 = (inp[13]) ? node6226 : node6215;
												assign node6215 = (inp[1]) ? node6221 : node6216;
													assign node6216 = (inp[14]) ? node6218 : 4'b0110;
														assign node6218 = (inp[7]) ? 4'b0110 : 4'b0111;
													assign node6221 = (inp[8]) ? node6223 : 4'b0110;
														assign node6223 = (inp[14]) ? 4'b1010 : 4'b1011;
												assign node6226 = (inp[2]) ? node6234 : node6227;
													assign node6227 = (inp[8]) ? node6231 : node6228;
														assign node6228 = (inp[7]) ? 4'b1010 : 4'b0110;
														assign node6231 = (inp[7]) ? 4'b1010 : 4'b1010;
													assign node6234 = (inp[8]) ? node6236 : 4'b1011;
														assign node6236 = (inp[7]) ? 4'b1010 : 4'b1011;
											assign node6239 = (inp[13]) ? node6251 : node6240;
												assign node6240 = (inp[7]) ? node6244 : node6241;
													assign node6241 = (inp[8]) ? 4'b1011 : 4'b1010;
													assign node6244 = (inp[1]) ? node6248 : node6245;
														assign node6245 = (inp[8]) ? 4'b1010 : 4'b1011;
														assign node6248 = (inp[8]) ? 4'b0010 : 4'b0011;
												assign node6251 = (inp[14]) ? node6257 : node6252;
													assign node6252 = (inp[2]) ? node6254 : 4'b0011;
														assign node6254 = (inp[7]) ? 4'b0010 : 4'b0011;
													assign node6257 = (inp[2]) ? 4'b0010 : 4'b1010;
									assign node6260 = (inp[6]) ? node6310 : node6261;
										assign node6261 = (inp[2]) ? node6285 : node6262;
											assign node6262 = (inp[13]) ? node6276 : node6263;
												assign node6263 = (inp[1]) ? node6269 : node6264;
													assign node6264 = (inp[11]) ? 4'b0011 : node6265;
														assign node6265 = (inp[8]) ? 4'b1011 : 4'b1010;
													assign node6269 = (inp[7]) ? node6273 : node6270;
														assign node6270 = (inp[11]) ? 4'b0010 : 4'b1011;
														assign node6273 = (inp[11]) ? 4'b1011 : 4'b0010;
												assign node6276 = (inp[1]) ? 4'b0011 : node6277;
													assign node6277 = (inp[11]) ? node6281 : node6278;
														assign node6278 = (inp[14]) ? 4'b0010 : 4'b1010;
														assign node6281 = (inp[14]) ? 4'b0010 : 4'b0010;
											assign node6285 = (inp[11]) ? node6299 : node6286;
												assign node6286 = (inp[1]) ? node6294 : node6287;
													assign node6287 = (inp[13]) ? node6291 : node6288;
														assign node6288 = (inp[8]) ? 4'b1011 : 4'b1010;
														assign node6291 = (inp[14]) ? 4'b0010 : 4'b0011;
													assign node6294 = (inp[7]) ? node6296 : 4'b0011;
														assign node6296 = (inp[8]) ? 4'b0010 : 4'b0011;
												assign node6299 = (inp[1]) ? node6305 : node6300;
													assign node6300 = (inp[14]) ? node6302 : 4'b0010;
														assign node6302 = (inp[7]) ? 4'b0011 : 4'b0010;
													assign node6305 = (inp[8]) ? 4'b1010 : node6306;
														assign node6306 = (inp[14]) ? 4'b0010 : 4'b1010;
										assign node6310 = (inp[7]) ? node6334 : node6311;
											assign node6311 = (inp[2]) ? node6325 : node6312;
												assign node6312 = (inp[11]) ? node6320 : node6313;
													assign node6313 = (inp[8]) ? node6317 : node6314;
														assign node6314 = (inp[14]) ? 4'b0010 : 4'b0011;
														assign node6317 = (inp[13]) ? 4'b1010 : 4'b0010;
													assign node6320 = (inp[13]) ? 4'b1010 : node6321;
														assign node6321 = (inp[1]) ? 4'b1011 : 4'b1010;
												assign node6325 = (inp[8]) ? node6327 : 4'b1010;
													assign node6327 = (inp[11]) ? node6331 : node6328;
														assign node6328 = (inp[13]) ? 4'b1011 : 4'b0011;
														assign node6331 = (inp[13]) ? 4'b0011 : 4'b1011;
											assign node6334 = (inp[14]) ? node6348 : node6335;
												assign node6335 = (inp[1]) ? node6343 : node6336;
													assign node6336 = (inp[11]) ? node6340 : node6337;
														assign node6337 = (inp[13]) ? 4'b0010 : 4'b0010;
														assign node6340 = (inp[13]) ? 4'b0011 : 4'b1010;
													assign node6343 = (inp[11]) ? node6345 : 4'b1011;
														assign node6345 = (inp[13]) ? 4'b0010 : 4'b0011;
												assign node6348 = (inp[8]) ? node6350 : 4'b0011;
													assign node6350 = (inp[1]) ? node6354 : node6351;
														assign node6351 = (inp[2]) ? 4'b0010 : 4'b1010;
														assign node6354 = (inp[11]) ? 4'b0010 : 4'b1010;
						assign node6357 = (inp[9]) ? node6701 : node6358;
							assign node6358 = (inp[12]) ? node6526 : node6359;
								assign node6359 = (inp[10]) ? node6441 : node6360;
									assign node6360 = (inp[14]) ? node6400 : node6361;
										assign node6361 = (inp[7]) ? node6375 : node6362;
											assign node6362 = (inp[8]) ? node6372 : node6363;
												assign node6363 = (inp[2]) ? node6365 : 4'b1011;
													assign node6365 = (inp[13]) ? node6369 : node6366;
														assign node6366 = (inp[1]) ? 4'b0010 : 4'b0010;
														assign node6369 = (inp[11]) ? 4'b0010 : 4'b0010;
												assign node6372 = (inp[2]) ? 4'b0011 : 4'b0010;
											assign node6375 = (inp[1]) ? node6387 : node6376;
												assign node6376 = (inp[8]) ? node6382 : node6377;
													assign node6377 = (inp[2]) ? 4'b0011 : node6378;
														assign node6378 = (inp[13]) ? 4'b1010 : 4'b0010;
													assign node6382 = (inp[2]) ? 4'b0010 : node6383;
														assign node6383 = (inp[6]) ? 4'b0011 : 4'b0011;
												assign node6387 = (inp[6]) ? node6393 : node6388;
													assign node6388 = (inp[11]) ? 4'b1011 : node6389;
														assign node6389 = (inp[8]) ? 4'b0011 : 4'b1010;
													assign node6393 = (inp[11]) ? node6397 : node6394;
														assign node6394 = (inp[8]) ? 4'b1010 : 4'b1011;
														assign node6397 = (inp[13]) ? 4'b0010 : 4'b0011;
										assign node6400 = (inp[8]) ? node6422 : node6401;
											assign node6401 = (inp[7]) ? node6413 : node6402;
												assign node6402 = (inp[11]) ? node6408 : node6403;
													assign node6403 = (inp[6]) ? node6405 : 4'b1010;
														assign node6405 = (inp[1]) ? 4'b0010 : 4'b0010;
													assign node6408 = (inp[13]) ? node6410 : 4'b1010;
														assign node6410 = (inp[1]) ? 4'b0010 : 4'b0010;
												assign node6413 = (inp[6]) ? 4'b0011 : node6414;
													assign node6414 = (inp[11]) ? node6418 : node6415;
														assign node6415 = (inp[13]) ? 4'b0011 : 4'b1011;
														assign node6418 = (inp[2]) ? 4'b1011 : 4'b0011;
											assign node6422 = (inp[7]) ? node6434 : node6423;
												assign node6423 = (inp[1]) ? node6429 : node6424;
													assign node6424 = (inp[2]) ? 4'b0011 : node6425;
														assign node6425 = (inp[11]) ? 4'b0011 : 4'b1011;
													assign node6429 = (inp[13]) ? 4'b1011 : node6430;
														assign node6430 = (inp[2]) ? 4'b1011 : 4'b0011;
												assign node6434 = (inp[2]) ? 4'b1010 : node6435;
													assign node6435 = (inp[11]) ? node6437 : 4'b1010;
														assign node6437 = (inp[1]) ? 4'b1010 : 4'b0010;
									assign node6441 = (inp[11]) ? node6489 : node6442;
										assign node6442 = (inp[6]) ? node6466 : node6443;
											assign node6443 = (inp[1]) ? node6453 : node6444;
												assign node6444 = (inp[8]) ? node6450 : node6445;
													assign node6445 = (inp[7]) ? node6447 : 4'b1010;
														assign node6447 = (inp[2]) ? 4'b0011 : 4'b1010;
													assign node6450 = (inp[13]) ? 4'b0011 : 4'b1011;
												assign node6453 = (inp[7]) ? node6461 : node6454;
													assign node6454 = (inp[13]) ? node6458 : node6455;
														assign node6455 = (inp[2]) ? 4'b1010 : 4'b0010;
														assign node6458 = (inp[14]) ? 4'b0010 : 4'b0011;
													assign node6461 = (inp[8]) ? node6463 : 4'b0011;
														assign node6463 = (inp[2]) ? 4'b0010 : 4'b0011;
											assign node6466 = (inp[13]) ? node6480 : node6467;
												assign node6467 = (inp[7]) ? node6473 : node6468;
													assign node6468 = (inp[1]) ? 4'b0010 : node6469;
														assign node6469 = (inp[2]) ? 4'b0011 : 4'b0010;
													assign node6473 = (inp[1]) ? node6477 : node6474;
														assign node6474 = (inp[14]) ? 4'b0011 : 4'b0010;
														assign node6477 = (inp[8]) ? 4'b1101 : 4'b0000;
												assign node6480 = (inp[14]) ? 4'b1101 : node6481;
													assign node6481 = (inp[1]) ? node6485 : node6482;
														assign node6482 = (inp[8]) ? 4'b1100 : 4'b0010;
														assign node6485 = (inp[7]) ? 4'b1101 : 4'b1100;
										assign node6489 = (inp[6]) ? node6509 : node6490;
											assign node6490 = (inp[8]) ? node6500 : node6491;
												assign node6491 = (inp[13]) ? 4'b0010 : node6492;
													assign node6492 = (inp[14]) ? node6496 : node6493;
														assign node6493 = (inp[7]) ? 4'b0010 : 4'b0011;
														assign node6496 = (inp[2]) ? 4'b0011 : 4'b1101;
												assign node6500 = (inp[1]) ? node6506 : node6501;
													assign node6501 = (inp[13]) ? node6503 : 4'b0010;
														assign node6503 = (inp[7]) ? 4'b1100 : 4'b1101;
													assign node6506 = (inp[14]) ? 4'b1100 : 4'b1101;
											assign node6509 = (inp[13]) ? node6519 : node6510;
												assign node6510 = (inp[7]) ? 4'b0101 : node6511;
													assign node6511 = (inp[1]) ? node6515 : node6512;
														assign node6512 = (inp[8]) ? 4'b1101 : 4'b1100;
														assign node6515 = (inp[2]) ? 4'b1100 : 4'b1100;
												assign node6519 = (inp[8]) ? node6521 : 4'b1101;
													assign node6521 = (inp[7]) ? node6523 : 4'b0101;
														assign node6523 = (inp[14]) ? 4'b0100 : 4'b0101;
								assign node6526 = (inp[10]) ? node6618 : node6527;
									assign node6527 = (inp[6]) ? node6579 : node6528;
										assign node6528 = (inp[11]) ? node6558 : node6529;
											assign node6529 = (inp[1]) ? node6545 : node6530;
												assign node6530 = (inp[13]) ? node6538 : node6531;
													assign node6531 = (inp[7]) ? node6535 : node6532;
														assign node6532 = (inp[8]) ? 4'b1011 : 4'b1010;
														assign node6535 = (inp[8]) ? 4'b1010 : 4'b1011;
													assign node6538 = (inp[8]) ? node6542 : node6539;
														assign node6539 = (inp[7]) ? 4'b0011 : 4'b1010;
														assign node6542 = (inp[7]) ? 4'b0010 : 4'b0011;
												assign node6545 = (inp[2]) ? node6553 : node6546;
													assign node6546 = (inp[14]) ? node6550 : node6547;
														assign node6547 = (inp[13]) ? 4'b0010 : 4'b1010;
														assign node6550 = (inp[8]) ? 4'b0010 : 4'b0010;
													assign node6553 = (inp[8]) ? node6555 : 4'b0011;
														assign node6555 = (inp[7]) ? 4'b0010 : 4'b0011;
											assign node6558 = (inp[1]) ? node6572 : node6559;
												assign node6559 = (inp[13]) ? node6567 : node6560;
													assign node6560 = (inp[8]) ? node6564 : node6561;
														assign node6561 = (inp[7]) ? 4'b0010 : 4'b0010;
														assign node6564 = (inp[7]) ? 4'b0010 : 4'b0011;
													assign node6567 = (inp[7]) ? 4'b1101 : node6568;
														assign node6568 = (inp[8]) ? 4'b0000 : 4'b0010;
												assign node6572 = (inp[2]) ? node6574 : 4'b1101;
													assign node6574 = (inp[13]) ? node6576 : 4'b0010;
														assign node6576 = (inp[8]) ? 4'b1101 : 4'b1100;
										assign node6579 = (inp[11]) ? node6597 : node6580;
											assign node6580 = (inp[1]) ? node6592 : node6581;
												assign node6581 = (inp[8]) ? node6587 : node6582;
													assign node6582 = (inp[7]) ? node6584 : 4'b0010;
														assign node6584 = (inp[14]) ? 4'b0001 : 4'b0010;
													assign node6587 = (inp[13]) ? node6589 : 4'b0010;
														assign node6589 = (inp[7]) ? 4'b1100 : 4'b1101;
												assign node6592 = (inp[14]) ? node6594 : 4'b1101;
													assign node6594 = (inp[7]) ? 4'b1100 : 4'b1101;
											assign node6597 = (inp[13]) ? node6607 : node6598;
												assign node6598 = (inp[2]) ? node6604 : node6599;
													assign node6599 = (inp[14]) ? node6601 : 4'b1101;
														assign node6601 = (inp[7]) ? 4'b1101 : 4'b1100;
													assign node6604 = (inp[1]) ? 4'b0101 : 4'b1101;
												assign node6607 = (inp[8]) ? node6613 : node6608;
													assign node6608 = (inp[1]) ? node6610 : 4'b1100;
														assign node6610 = (inp[14]) ? 4'b0101 : 4'b0100;
													assign node6613 = (inp[7]) ? node6615 : 4'b0101;
														assign node6615 = (inp[14]) ? 4'b0100 : 4'b0101;
									assign node6618 = (inp[8]) ? node6656 : node6619;
										assign node6619 = (inp[7]) ? node6639 : node6620;
											assign node6620 = (inp[14]) ? node6624 : node6621;
												assign node6621 = (inp[2]) ? 4'b0100 : 4'b0101;
												assign node6624 = (inp[2]) ? node6632 : node6625;
													assign node6625 = (inp[11]) ? node6629 : node6626;
														assign node6626 = (inp[6]) ? 4'b0100 : 4'b0100;
														assign node6629 = (inp[13]) ? 4'b1100 : 4'b0100;
													assign node6632 = (inp[11]) ? node6636 : node6633;
														assign node6633 = (inp[6]) ? 4'b0100 : 4'b1100;
														assign node6636 = (inp[1]) ? 4'b1100 : 4'b0100;
											assign node6639 = (inp[14]) ? node6649 : node6640;
												assign node6640 = (inp[2]) ? node6646 : node6641;
													assign node6641 = (inp[6]) ? 4'b0100 : node6642;
														assign node6642 = (inp[11]) ? 4'b0100 : 4'b1100;
													assign node6646 = (inp[13]) ? 4'b0101 : 4'b1101;
												assign node6649 = (inp[1]) ? 4'b0101 : node6650;
													assign node6650 = (inp[13]) ? node6652 : 4'b1101;
														assign node6652 = (inp[2]) ? 4'b0101 : 4'b0101;
										assign node6656 = (inp[7]) ? node6678 : node6657;
											assign node6657 = (inp[14]) ? node6665 : node6658;
												assign node6658 = (inp[2]) ? node6662 : node6659;
													assign node6659 = (inp[1]) ? 4'b0100 : 4'b1100;
													assign node6662 = (inp[13]) ? 4'b1101 : 4'b0101;
												assign node6665 = (inp[6]) ? node6671 : node6666;
													assign node6666 = (inp[1]) ? node6668 : 4'b0101;
														assign node6668 = (inp[13]) ? 4'b0101 : 4'b1101;
													assign node6671 = (inp[11]) ? node6675 : node6672;
														assign node6672 = (inp[1]) ? 4'b1101 : 4'b0101;
														assign node6675 = (inp[13]) ? 4'b0101 : 4'b1101;
											assign node6678 = (inp[14]) ? node6690 : node6679;
												assign node6679 = (inp[2]) ? node6685 : node6680;
													assign node6680 = (inp[1]) ? node6682 : 4'b0101;
														assign node6682 = (inp[13]) ? 4'b0101 : 4'b1101;
													assign node6685 = (inp[11]) ? 4'b0100 : node6686;
														assign node6686 = (inp[1]) ? 4'b1100 : 4'b0100;
												assign node6690 = (inp[1]) ? node6696 : node6691;
													assign node6691 = (inp[13]) ? 4'b0100 : node6692;
														assign node6692 = (inp[2]) ? 4'b0100 : 4'b1100;
													assign node6696 = (inp[6]) ? 4'b1100 : node6697;
														assign node6697 = (inp[11]) ? 4'b1100 : 4'b0100;
							assign node6701 = (inp[10]) ? node6889 : node6702;
								assign node6702 = (inp[12]) ? node6794 : node6703;
									assign node6703 = (inp[13]) ? node6751 : node6704;
										assign node6704 = (inp[2]) ? node6728 : node6705;
											assign node6705 = (inp[6]) ? node6715 : node6706;
												assign node6706 = (inp[14]) ? node6710 : node6707;
													assign node6707 = (inp[11]) ? 4'b0100 : 4'b1100;
													assign node6710 = (inp[11]) ? node6712 : 4'b0101;
														assign node6712 = (inp[7]) ? 4'b0101 : 4'b0100;
												assign node6715 = (inp[11]) ? node6723 : node6716;
													assign node6716 = (inp[7]) ? node6720 : node6717;
														assign node6717 = (inp[8]) ? 4'b0100 : 4'b0101;
														assign node6720 = (inp[8]) ? 4'b1100 : 4'b0100;
													assign node6723 = (inp[14]) ? 4'b0101 : node6724;
														assign node6724 = (inp[8]) ? 4'b1101 : 4'b1100;
											assign node6728 = (inp[11]) ? node6742 : node6729;
												assign node6729 = (inp[14]) ? node6737 : node6730;
													assign node6730 = (inp[6]) ? node6734 : node6731;
														assign node6731 = (inp[7]) ? 4'b1100 : 4'b1100;
														assign node6734 = (inp[1]) ? 4'b1101 : 4'b0101;
													assign node6737 = (inp[7]) ? 4'b1100 : node6738;
														assign node6738 = (inp[6]) ? 4'b0100 : 4'b0101;
												assign node6742 = (inp[1]) ? node6748 : node6743;
													assign node6743 = (inp[7]) ? node6745 : 4'b1100;
														assign node6745 = (inp[8]) ? 4'b1100 : 4'b1101;
													assign node6748 = (inp[6]) ? 4'b0101 : 4'b1101;
										assign node6751 = (inp[2]) ? node6779 : node6752;
											assign node6752 = (inp[6]) ? node6766 : node6753;
												assign node6753 = (inp[11]) ? node6761 : node6754;
													assign node6754 = (inp[7]) ? node6758 : node6755;
														assign node6755 = (inp[1]) ? 4'b0100 : 4'b1100;
														assign node6758 = (inp[1]) ? 4'b0101 : 4'b0100;
													assign node6761 = (inp[7]) ? node6763 : 4'b0100;
														assign node6763 = (inp[8]) ? 4'b1100 : 4'b1100;
												assign node6766 = (inp[14]) ? node6772 : node6767;
													assign node6767 = (inp[8]) ? 4'b0101 : node6768;
														assign node6768 = (inp[7]) ? 4'b1100 : 4'b1101;
													assign node6772 = (inp[8]) ? node6776 : node6773;
														assign node6773 = (inp[7]) ? 4'b0101 : 4'b0100;
														assign node6776 = (inp[11]) ? 4'b0101 : 4'b1101;
											assign node6779 = (inp[8]) ? node6789 : node6780;
												assign node6780 = (inp[11]) ? node6784 : node6781;
													assign node6781 = (inp[7]) ? 4'b1101 : 4'b1100;
													assign node6784 = (inp[14]) ? node6786 : 4'b0100;
														assign node6786 = (inp[6]) ? 4'b0100 : 4'b0100;
												assign node6789 = (inp[7]) ? 4'b0100 : node6790;
													assign node6790 = (inp[1]) ? 4'b1101 : 4'b0101;
									assign node6794 = (inp[6]) ? node6842 : node6795;
										assign node6795 = (inp[11]) ? node6819 : node6796;
											assign node6796 = (inp[8]) ? node6810 : node6797;
												assign node6797 = (inp[1]) ? node6803 : node6798;
													assign node6798 = (inp[13]) ? 4'b1100 : node6799;
														assign node6799 = (inp[2]) ? 4'b1100 : 4'b1100;
													assign node6803 = (inp[2]) ? node6807 : node6804;
														assign node6804 = (inp[13]) ? 4'b0100 : 4'b1100;
														assign node6807 = (inp[7]) ? 4'b0101 : 4'b1100;
												assign node6810 = (inp[1]) ? 4'b0101 : node6811;
													assign node6811 = (inp[2]) ? node6815 : node6812;
														assign node6812 = (inp[7]) ? 4'b0100 : 4'b1100;
														assign node6815 = (inp[7]) ? 4'b0100 : 4'b0101;
											assign node6819 = (inp[1]) ? node6833 : node6820;
												assign node6820 = (inp[13]) ? node6826 : node6821;
													assign node6821 = (inp[2]) ? node6823 : 4'b0100;
														assign node6823 = (inp[8]) ? 4'b0100 : 4'b0101;
													assign node6826 = (inp[2]) ? node6830 : node6827;
														assign node6827 = (inp[14]) ? 4'b1000 : 4'b0100;
														assign node6830 = (inp[14]) ? 4'b0100 : 4'b1001;
												assign node6833 = (inp[13]) ? node6839 : node6834;
													assign node6834 = (inp[7]) ? 4'b1000 : node6835;
														assign node6835 = (inp[14]) ? 4'b0000 : 4'b0100;
													assign node6839 = (inp[14]) ? 4'b1001 : 4'b1000;
										assign node6842 = (inp[11]) ? node6862 : node6843;
											assign node6843 = (inp[13]) ? node6849 : node6844;
												assign node6844 = (inp[8]) ? node6846 : 4'b0100;
													assign node6846 = (inp[1]) ? 4'b0100 : 4'b0101;
												assign node6849 = (inp[2]) ? node6857 : node6850;
													assign node6850 = (inp[7]) ? node6854 : node6851;
														assign node6851 = (inp[14]) ? 4'b1001 : 4'b0000;
														assign node6854 = (inp[14]) ? 4'b1000 : 4'b1001;
													assign node6857 = (inp[1]) ? 4'b1000 : node6858;
														assign node6858 = (inp[8]) ? 4'b1000 : 4'b1001;
											assign node6862 = (inp[1]) ? node6874 : node6863;
												assign node6863 = (inp[2]) ? node6869 : node6864;
													assign node6864 = (inp[13]) ? 4'b1001 : node6865;
														assign node6865 = (inp[8]) ? 4'b1001 : 4'b1000;
													assign node6869 = (inp[7]) ? 4'b0000 : node6870;
														assign node6870 = (inp[8]) ? 4'b1001 : 4'b1000;
												assign node6874 = (inp[13]) ? node6882 : node6875;
													assign node6875 = (inp[8]) ? node6879 : node6876;
														assign node6876 = (inp[2]) ? 4'b1000 : 4'b1001;
														assign node6879 = (inp[7]) ? 4'b0000 : 4'b0001;
													assign node6882 = (inp[2]) ? node6886 : node6883;
														assign node6883 = (inp[7]) ? 4'b0000 : 4'b0000;
														assign node6886 = (inp[8]) ? 4'b0000 : 4'b0001;
								assign node6889 = (inp[12]) ? node6975 : node6890;
									assign node6890 = (inp[11]) ? node6934 : node6891;
										assign node6891 = (inp[6]) ? node6913 : node6892;
											assign node6892 = (inp[13]) ? node6906 : node6893;
												assign node6893 = (inp[8]) ? node6899 : node6894;
													assign node6894 = (inp[7]) ? node6896 : 4'b1100;
														assign node6896 = (inp[14]) ? 4'b1101 : 4'b1100;
													assign node6899 = (inp[1]) ? node6903 : node6900;
														assign node6900 = (inp[14]) ? 4'b1100 : 4'b1101;
														assign node6903 = (inp[14]) ? 4'b0100 : 4'b0101;
												assign node6906 = (inp[7]) ? node6908 : 4'b0101;
													assign node6908 = (inp[8]) ? 4'b0100 : node6909;
														assign node6909 = (inp[14]) ? 4'b0101 : 4'b0100;
											assign node6913 = (inp[1]) ? node6923 : node6914;
												assign node6914 = (inp[2]) ? node6918 : node6915;
													assign node6915 = (inp[8]) ? 4'b0101 : 4'b0100;
													assign node6918 = (inp[13]) ? node6920 : 4'b0101;
														assign node6920 = (inp[14]) ? 4'b1001 : 4'b0000;
												assign node6923 = (inp[13]) ? node6931 : node6924;
													assign node6924 = (inp[7]) ? node6928 : node6925;
														assign node6925 = (inp[8]) ? 4'b0000 : 4'b0100;
														assign node6928 = (inp[8]) ? 4'b1000 : 4'b0000;
													assign node6931 = (inp[2]) ? 4'b1000 : 4'b1001;
										assign node6934 = (inp[6]) ? node6958 : node6935;
											assign node6935 = (inp[1]) ? node6945 : node6936;
												assign node6936 = (inp[8]) ? node6940 : node6937;
													assign node6937 = (inp[7]) ? 4'b0101 : 4'b0100;
													assign node6940 = (inp[14]) ? 4'b1001 : node6941;
														assign node6941 = (inp[7]) ? 4'b1000 : 4'b0100;
												assign node6945 = (inp[13]) ? node6951 : node6946;
													assign node6946 = (inp[7]) ? 4'b1001 : node6947;
														assign node6947 = (inp[14]) ? 4'b1001 : 4'b0000;
													assign node6951 = (inp[7]) ? node6955 : node6952;
														assign node6952 = (inp[8]) ? 4'b1000 : 4'b1000;
														assign node6955 = (inp[2]) ? 4'b1001 : 4'b1000;
											assign node6958 = (inp[13]) ? node6968 : node6959;
												assign node6959 = (inp[8]) ? node6965 : node6960;
													assign node6960 = (inp[7]) ? node6962 : 4'b1001;
														assign node6962 = (inp[14]) ? 4'b1001 : 4'b1000;
													assign node6965 = (inp[1]) ? 4'b0001 : 4'b1001;
												assign node6968 = (inp[1]) ? node6970 : 4'b0001;
													assign node6970 = (inp[8]) ? 4'b0000 : node6971;
														assign node6971 = (inp[2]) ? 4'b0000 : 4'b0001;
									assign node6975 = (inp[1]) ? node7029 : node6976;
										assign node6976 = (inp[8]) ? node7006 : node6977;
											assign node6977 = (inp[7]) ? node6993 : node6978;
												assign node6978 = (inp[2]) ? node6986 : node6979;
													assign node6979 = (inp[14]) ? node6983 : node6980;
														assign node6980 = (inp[6]) ? 4'b1001 : 4'b0001;
														assign node6983 = (inp[13]) ? 4'b0000 : 4'b1000;
													assign node6986 = (inp[11]) ? node6990 : node6987;
														assign node6987 = (inp[6]) ? 4'b0000 : 4'b1000;
														assign node6990 = (inp[6]) ? 4'b1000 : 4'b0000;
												assign node6993 = (inp[2]) ? node6999 : node6994;
													assign node6994 = (inp[14]) ? node6996 : 4'b1000;
														assign node6996 = (inp[6]) ? 4'b0001 : 4'b1001;
													assign node6999 = (inp[14]) ? node7003 : node7000;
														assign node7000 = (inp[13]) ? 4'b0001 : 4'b1001;
														assign node7003 = (inp[6]) ? 4'b1001 : 4'b0001;
											assign node7006 = (inp[7]) ? node7016 : node7007;
												assign node7007 = (inp[2]) ? node7013 : node7008;
													assign node7008 = (inp[13]) ? 4'b1001 : node7009;
														assign node7009 = (inp[6]) ? 4'b1000 : 4'b0000;
													assign node7013 = (inp[14]) ? 4'b0001 : 4'b1001;
												assign node7016 = (inp[14]) ? node7022 : node7017;
													assign node7017 = (inp[6]) ? 4'b1000 : node7018;
														assign node7018 = (inp[11]) ? 4'b1000 : 4'b0000;
													assign node7022 = (inp[6]) ? node7026 : node7023;
														assign node7023 = (inp[11]) ? 4'b1000 : 4'b0000;
														assign node7026 = (inp[11]) ? 4'b0000 : 4'b1000;
										assign node7029 = (inp[6]) ? node7049 : node7030;
											assign node7030 = (inp[11]) ? node7040 : node7031;
												assign node7031 = (inp[2]) ? 4'b0001 : node7032;
													assign node7032 = (inp[13]) ? node7036 : node7033;
														assign node7033 = (inp[8]) ? 4'b0000 : 4'b1000;
														assign node7036 = (inp[7]) ? 4'b0001 : 4'b0000;
												assign node7040 = (inp[8]) ? node7046 : node7041;
													assign node7041 = (inp[2]) ? 4'b0000 : node7042;
														assign node7042 = (inp[14]) ? 4'b1001 : 4'b0001;
													assign node7046 = (inp[7]) ? 4'b1000 : 4'b1001;
											assign node7049 = (inp[7]) ? node7059 : node7050;
												assign node7050 = (inp[11]) ? node7054 : node7051;
													assign node7051 = (inp[13]) ? 4'b1000 : 4'b0000;
													assign node7054 = (inp[13]) ? node7056 : 4'b1000;
														assign node7056 = (inp[8]) ? 4'b0001 : 4'b0000;
												assign node7059 = (inp[11]) ? node7065 : node7060;
													assign node7060 = (inp[14]) ? 4'b1001 : node7061;
														assign node7061 = (inp[8]) ? 4'b1001 : 4'b0000;
													assign node7065 = (inp[2]) ? node7067 : 4'b0001;
														assign node7067 = (inp[8]) ? 4'b0000 : 4'b0001;
					assign node7070 = (inp[9]) ? node7808 : node7071;
						assign node7071 = (inp[12]) ? node7441 : node7072;
							assign node7072 = (inp[5]) ? node7248 : node7073;
								assign node7073 = (inp[10]) ? node7157 : node7074;
									assign node7074 = (inp[11]) ? node7110 : node7075;
										assign node7075 = (inp[6]) ? node7091 : node7076;
											assign node7076 = (inp[13]) ? node7084 : node7077;
												assign node7077 = (inp[7]) ? node7081 : node7078;
													assign node7078 = (inp[8]) ? 4'b1011 : 4'b1010;
													assign node7081 = (inp[8]) ? 4'b0010 : 4'b0011;
												assign node7084 = (inp[2]) ? 4'b0011 : node7085;
													assign node7085 = (inp[8]) ? 4'b0011 : node7086;
														assign node7086 = (inp[14]) ? 4'b0010 : 4'b0011;
											assign node7091 = (inp[13]) ? node7103 : node7092;
												assign node7092 = (inp[1]) ? node7098 : node7093;
													assign node7093 = (inp[8]) ? 4'b0011 : node7094;
														assign node7094 = (inp[14]) ? 4'b0010 : 4'b0010;
													assign node7098 = (inp[14]) ? 4'b1011 : node7099;
														assign node7099 = (inp[8]) ? 4'b0010 : 4'b1011;
												assign node7103 = (inp[8]) ? node7107 : node7104;
													assign node7104 = (inp[1]) ? 4'b1011 : 4'b0010;
													assign node7107 = (inp[7]) ? 4'b1010 : 4'b1011;
										assign node7110 = (inp[7]) ? node7132 : node7111;
											assign node7111 = (inp[8]) ? node7121 : node7112;
												assign node7112 = (inp[6]) ? node7116 : node7113;
													assign node7113 = (inp[13]) ? 4'b1010 : 4'b0010;
													assign node7116 = (inp[1]) ? node7118 : 4'b1010;
														assign node7118 = (inp[14]) ? 4'b0010 : 4'b1010;
												assign node7121 = (inp[14]) ? node7127 : node7122;
													assign node7122 = (inp[2]) ? 4'b1011 : node7123;
														assign node7123 = (inp[6]) ? 4'b1010 : 4'b0010;
													assign node7127 = (inp[2]) ? node7129 : 4'b0011;
														assign node7129 = (inp[6]) ? 4'b0011 : 4'b1011;
											assign node7132 = (inp[8]) ? node7144 : node7133;
												assign node7133 = (inp[2]) ? node7139 : node7134;
													assign node7134 = (inp[6]) ? node7136 : 4'b0010;
														assign node7136 = (inp[14]) ? 4'b1011 : 4'b1010;
													assign node7139 = (inp[6]) ? node7141 : 4'b0011;
														assign node7141 = (inp[1]) ? 4'b0011 : 4'b0011;
												assign node7144 = (inp[2]) ? node7152 : node7145;
													assign node7145 = (inp[14]) ? node7149 : node7146;
														assign node7146 = (inp[13]) ? 4'b0011 : 4'b1011;
														assign node7149 = (inp[1]) ? 4'b0010 : 4'b0010;
													assign node7152 = (inp[1]) ? node7154 : 4'b0010;
														assign node7154 = (inp[13]) ? 4'b0010 : 4'b1010;
									assign node7157 = (inp[6]) ? node7205 : node7158;
										assign node7158 = (inp[11]) ? node7180 : node7159;
											assign node7159 = (inp[1]) ? node7171 : node7160;
												assign node7160 = (inp[13]) ? node7166 : node7161;
													assign node7161 = (inp[8]) ? 4'b1010 : node7162;
														assign node7162 = (inp[2]) ? 4'b1011 : 4'b1010;
													assign node7166 = (inp[2]) ? node7168 : 4'b0011;
														assign node7168 = (inp[8]) ? 4'b0010 : 4'b1010;
												assign node7171 = (inp[13]) ? 4'b0011 : node7172;
													assign node7172 = (inp[8]) ? node7176 : node7173;
														assign node7173 = (inp[14]) ? 4'b0011 : 4'b1010;
														assign node7176 = (inp[7]) ? 4'b0010 : 4'b0011;
											assign node7180 = (inp[1]) ? node7192 : node7181;
												assign node7181 = (inp[7]) ? node7189 : node7182;
													assign node7182 = (inp[8]) ? node7186 : node7183;
														assign node7183 = (inp[13]) ? 4'b0010 : 4'b0010;
														assign node7186 = (inp[13]) ? 4'b0010 : 4'b0011;
													assign node7189 = (inp[13]) ? 4'b1101 : 4'b0011;
												assign node7192 = (inp[13]) ? node7200 : node7193;
													assign node7193 = (inp[2]) ? node7197 : node7194;
														assign node7194 = (inp[14]) ? 4'b1101 : 4'b0010;
														assign node7197 = (inp[14]) ? 4'b1100 : 4'b1101;
													assign node7200 = (inp[2]) ? node7202 : 4'b1100;
														assign node7202 = (inp[14]) ? 4'b1100 : 4'b1100;
										assign node7205 = (inp[11]) ? node7227 : node7206;
											assign node7206 = (inp[13]) ? node7222 : node7207;
												assign node7207 = (inp[1]) ? node7215 : node7208;
													assign node7208 = (inp[8]) ? node7212 : node7209;
														assign node7209 = (inp[7]) ? 4'b0010 : 4'b0010;
														assign node7212 = (inp[2]) ? 4'b0011 : 4'b0010;
													assign node7215 = (inp[8]) ? node7219 : node7216;
														assign node7216 = (inp[7]) ? 4'b1101 : 4'b0010;
														assign node7219 = (inp[7]) ? 4'b1100 : 4'b1101;
												assign node7222 = (inp[14]) ? 4'b1101 : node7223;
													assign node7223 = (inp[2]) ? 4'b1101 : 4'b0010;
											assign node7227 = (inp[13]) ? node7239 : node7228;
												assign node7228 = (inp[14]) ? node7236 : node7229;
													assign node7229 = (inp[7]) ? node7233 : node7230;
														assign node7230 = (inp[8]) ? 4'b1100 : 4'b1101;
														assign node7233 = (inp[1]) ? 4'b0101 : 4'b1101;
													assign node7236 = (inp[8]) ? 4'b0100 : 4'b1100;
												assign node7239 = (inp[8]) ? 4'b0101 : node7240;
													assign node7240 = (inp[1]) ? node7244 : node7241;
														assign node7241 = (inp[14]) ? 4'b1100 : 4'b0100;
														assign node7244 = (inp[2]) ? 4'b0100 : 4'b0101;
								assign node7248 = (inp[10]) ? node7344 : node7249;
									assign node7249 = (inp[8]) ? node7295 : node7250;
										assign node7250 = (inp[13]) ? node7278 : node7251;
											assign node7251 = (inp[1]) ? node7267 : node7252;
												assign node7252 = (inp[6]) ? node7260 : node7253;
													assign node7253 = (inp[11]) ? node7257 : node7254;
														assign node7254 = (inp[14]) ? 4'b1000 : 4'b1001;
														assign node7257 = (inp[14]) ? 4'b0001 : 4'b0000;
													assign node7260 = (inp[11]) ? node7264 : node7261;
														assign node7261 = (inp[2]) ? 4'b0000 : 4'b0001;
														assign node7264 = (inp[7]) ? 4'b1000 : 4'b1000;
												assign node7267 = (inp[14]) ? node7275 : node7268;
													assign node7268 = (inp[7]) ? node7272 : node7269;
														assign node7269 = (inp[6]) ? 4'b1000 : 4'b0001;
														assign node7272 = (inp[11]) ? 4'b0000 : 4'b1000;
													assign node7275 = (inp[7]) ? 4'b0001 : 4'b0000;
											assign node7278 = (inp[2]) ? node7290 : node7279;
												assign node7279 = (inp[7]) ? node7285 : node7280;
													assign node7280 = (inp[14]) ? 4'b0000 : node7281;
														assign node7281 = (inp[1]) ? 4'b0001 : 4'b1001;
													assign node7285 = (inp[14]) ? 4'b1001 : node7286;
														assign node7286 = (inp[1]) ? 4'b1000 : 4'b0000;
												assign node7290 = (inp[11]) ? node7292 : 4'b0001;
													assign node7292 = (inp[6]) ? 4'b0001 : 4'b1001;
										assign node7295 = (inp[7]) ? node7317 : node7296;
											assign node7296 = (inp[14]) ? node7306 : node7297;
												assign node7297 = (inp[2]) ? 4'b1001 : node7298;
													assign node7298 = (inp[1]) ? node7302 : node7299;
														assign node7299 = (inp[13]) ? 4'b0000 : 4'b1000;
														assign node7302 = (inp[11]) ? 4'b0000 : 4'b0000;
												assign node7306 = (inp[6]) ? node7312 : node7307;
													assign node7307 = (inp[11]) ? 4'b1001 : node7308;
														assign node7308 = (inp[1]) ? 4'b0001 : 4'b1001;
													assign node7312 = (inp[11]) ? 4'b0001 : node7313;
														assign node7313 = (inp[13]) ? 4'b1001 : 4'b0001;
											assign node7317 = (inp[14]) ? node7331 : node7318;
												assign node7318 = (inp[2]) ? node7326 : node7319;
													assign node7319 = (inp[1]) ? node7323 : node7320;
														assign node7320 = (inp[6]) ? 4'b0001 : 4'b1001;
														assign node7323 = (inp[11]) ? 4'b0001 : 4'b0001;
													assign node7326 = (inp[6]) ? node7328 : 4'b0000;
														assign node7328 = (inp[13]) ? 4'b0000 : 4'b1000;
												assign node7331 = (inp[1]) ? node7337 : node7332;
													assign node7332 = (inp[13]) ? node7334 : 4'b0000;
														assign node7334 = (inp[2]) ? 4'b0000 : 4'b1000;
													assign node7337 = (inp[6]) ? node7341 : node7338;
														assign node7338 = (inp[11]) ? 4'b1000 : 4'b0000;
														assign node7341 = (inp[11]) ? 4'b0000 : 4'b1000;
									assign node7344 = (inp[11]) ? node7390 : node7345;
										assign node7345 = (inp[6]) ? node7371 : node7346;
											assign node7346 = (inp[8]) ? node7358 : node7347;
												assign node7347 = (inp[7]) ? node7353 : node7348;
													assign node7348 = (inp[13]) ? node7350 : 4'b1000;
														assign node7350 = (inp[2]) ? 4'b1000 : 4'b1001;
													assign node7353 = (inp[14]) ? 4'b0001 : node7354;
														assign node7354 = (inp[1]) ? 4'b0000 : 4'b1000;
												assign node7358 = (inp[7]) ? node7364 : node7359;
													assign node7359 = (inp[1]) ? 4'b0001 : node7360;
														assign node7360 = (inp[13]) ? 4'b0001 : 4'b1001;
													assign node7364 = (inp[1]) ? node7368 : node7365;
														assign node7365 = (inp[13]) ? 4'b0000 : 4'b1000;
														assign node7368 = (inp[14]) ? 4'b0000 : 4'b0001;
											assign node7371 = (inp[13]) ? node7379 : node7372;
												assign node7372 = (inp[14]) ? node7376 : node7373;
													assign node7373 = (inp[7]) ? 4'b0001 : 4'b0000;
													assign node7376 = (inp[1]) ? 4'b1101 : 4'b0001;
												assign node7379 = (inp[8]) ? node7385 : node7380;
													assign node7380 = (inp[14]) ? node7382 : 4'b0000;
														assign node7382 = (inp[7]) ? 4'b1101 : 4'b0000;
													assign node7385 = (inp[7]) ? node7387 : 4'b1101;
														assign node7387 = (inp[14]) ? 4'b1100 : 4'b1101;
										assign node7390 = (inp[1]) ? node7416 : node7391;
											assign node7391 = (inp[6]) ? node7405 : node7392;
												assign node7392 = (inp[13]) ? node7400 : node7393;
													assign node7393 = (inp[7]) ? node7397 : node7394;
														assign node7394 = (inp[14]) ? 4'b0001 : 4'b0000;
														assign node7397 = (inp[8]) ? 4'b0000 : 4'b0000;
													assign node7400 = (inp[7]) ? node7402 : 4'b0000;
														assign node7402 = (inp[8]) ? 4'b1100 : 4'b1101;
												assign node7405 = (inp[13]) ? node7411 : node7406;
													assign node7406 = (inp[14]) ? 4'b1100 : node7407;
														assign node7407 = (inp[8]) ? 4'b1101 : 4'b1100;
													assign node7411 = (inp[7]) ? 4'b0101 : node7412;
														assign node7412 = (inp[2]) ? 4'b0101 : 4'b1100;
											assign node7416 = (inp[6]) ? node7430 : node7417;
												assign node7417 = (inp[13]) ? node7423 : node7418;
													assign node7418 = (inp[7]) ? 4'b1101 : node7419;
														assign node7419 = (inp[14]) ? 4'b1101 : 4'b0001;
													assign node7423 = (inp[2]) ? node7427 : node7424;
														assign node7424 = (inp[7]) ? 4'b1100 : 4'b1100;
														assign node7427 = (inp[8]) ? 4'b1100 : 4'b1101;
												assign node7430 = (inp[13]) ? node7438 : node7431;
													assign node7431 = (inp[7]) ? node7435 : node7432;
														assign node7432 = (inp[14]) ? 4'b1100 : 4'b1100;
														assign node7435 = (inp[14]) ? 4'b0100 : 4'b0101;
													assign node7438 = (inp[8]) ? 4'b0101 : 4'b0100;
							assign node7441 = (inp[10]) ? node7631 : node7442;
								assign node7442 = (inp[6]) ? node7538 : node7443;
									assign node7443 = (inp[5]) ? node7493 : node7444;
										assign node7444 = (inp[11]) ? node7470 : node7445;
											assign node7445 = (inp[13]) ? node7459 : node7446;
												assign node7446 = (inp[1]) ? node7454 : node7447;
													assign node7447 = (inp[2]) ? node7451 : node7448;
														assign node7448 = (inp[14]) ? 4'b1010 : 4'b1011;
														assign node7451 = (inp[14]) ? 4'b1010 : 4'b1010;
													assign node7454 = (inp[2]) ? 4'b0011 : node7455;
														assign node7455 = (inp[14]) ? 4'b1010 : 4'b1011;
												assign node7459 = (inp[2]) ? node7465 : node7460;
													assign node7460 = (inp[14]) ? node7462 : 4'b1010;
														assign node7462 = (inp[1]) ? 4'b0010 : 4'b0010;
													assign node7465 = (inp[14]) ? node7467 : 4'b0011;
														assign node7467 = (inp[8]) ? 4'b0011 : 4'b1010;
											assign node7470 = (inp[1]) ? node7484 : node7471;
												assign node7471 = (inp[8]) ? node7477 : node7472;
													assign node7472 = (inp[7]) ? node7474 : 4'b0010;
														assign node7474 = (inp[14]) ? 4'b0011 : 4'b0010;
													assign node7477 = (inp[13]) ? node7481 : node7478;
														assign node7478 = (inp[2]) ? 4'b0011 : 4'b0010;
														assign node7481 = (inp[7]) ? 4'b1100 : 4'b1101;
												assign node7484 = (inp[14]) ? node7490 : node7485;
													assign node7485 = (inp[13]) ? 4'b1100 : node7486;
														assign node7486 = (inp[7]) ? 4'b1100 : 4'b1101;
													assign node7490 = (inp[13]) ? 4'b1101 : 4'b1100;
										assign node7493 = (inp[11]) ? node7519 : node7494;
											assign node7494 = (inp[1]) ? node7504 : node7495;
												assign node7495 = (inp[7]) ? node7501 : node7496;
													assign node7496 = (inp[13]) ? node7498 : 4'b1000;
														assign node7498 = (inp[14]) ? 4'b0001 : 4'b1000;
													assign node7501 = (inp[8]) ? 4'b0001 : 4'b1001;
												assign node7504 = (inp[2]) ? node7512 : node7505;
													assign node7505 = (inp[14]) ? node7509 : node7506;
														assign node7506 = (inp[13]) ? 4'b0000 : 4'b1000;
														assign node7509 = (inp[8]) ? 4'b0000 : 4'b0000;
													assign node7512 = (inp[7]) ? node7516 : node7513;
														assign node7513 = (inp[8]) ? 4'b0001 : 4'b0000;
														assign node7516 = (inp[8]) ? 4'b0000 : 4'b0001;
											assign node7519 = (inp[1]) ? node7525 : node7520;
												assign node7520 = (inp[13]) ? node7522 : 4'b0001;
													assign node7522 = (inp[7]) ? 4'b1101 : 4'b0000;
												assign node7525 = (inp[7]) ? node7531 : node7526;
													assign node7526 = (inp[13]) ? 4'b1100 : node7527;
														assign node7527 = (inp[8]) ? 4'b1101 : 4'b0000;
													assign node7531 = (inp[8]) ? node7535 : node7532;
														assign node7532 = (inp[2]) ? 4'b1101 : 4'b1100;
														assign node7535 = (inp[14]) ? 4'b1100 : 4'b1101;
									assign node7538 = (inp[11]) ? node7590 : node7539;
										assign node7539 = (inp[13]) ? node7565 : node7540;
											assign node7540 = (inp[1]) ? node7552 : node7541;
												assign node7541 = (inp[5]) ? node7547 : node7542;
													assign node7542 = (inp[14]) ? node7544 : 4'b0011;
														assign node7544 = (inp[8]) ? 4'b0010 : 4'b0011;
													assign node7547 = (inp[2]) ? node7549 : 4'b0001;
														assign node7549 = (inp[7]) ? 4'b0000 : 4'b0001;
												assign node7552 = (inp[7]) ? node7560 : node7553;
													assign node7553 = (inp[5]) ? node7557 : node7554;
														assign node7554 = (inp[8]) ? 4'b1101 : 4'b0010;
														assign node7557 = (inp[8]) ? 4'b0000 : 4'b0000;
													assign node7560 = (inp[8]) ? node7562 : 4'b1101;
														assign node7562 = (inp[14]) ? 4'b1100 : 4'b1100;
											assign node7565 = (inp[14]) ? node7577 : node7566;
												assign node7566 = (inp[1]) ? node7572 : node7567;
													assign node7567 = (inp[8]) ? 4'b1101 : node7568;
														assign node7568 = (inp[5]) ? 4'b0000 : 4'b0010;
													assign node7572 = (inp[8]) ? node7574 : 4'b1101;
														assign node7574 = (inp[7]) ? 4'b1101 : 4'b1100;
												assign node7577 = (inp[5]) ? node7583 : node7578;
													assign node7578 = (inp[7]) ? node7580 : 4'b1101;
														assign node7580 = (inp[8]) ? 4'b1100 : 4'b1101;
													assign node7583 = (inp[8]) ? node7587 : node7584;
														assign node7584 = (inp[7]) ? 4'b1101 : 4'b1100;
														assign node7587 = (inp[7]) ? 4'b1100 : 4'b1101;
										assign node7590 = (inp[1]) ? node7614 : node7591;
											assign node7591 = (inp[13]) ? node7603 : node7592;
												assign node7592 = (inp[14]) ? node7598 : node7593;
													assign node7593 = (inp[2]) ? node7595 : 4'b1101;
														assign node7595 = (inp[8]) ? 4'b1101 : 4'b1100;
													assign node7598 = (inp[7]) ? 4'b1100 : node7599;
														assign node7599 = (inp[8]) ? 4'b1101 : 4'b1100;
												assign node7603 = (inp[8]) ? node7611 : node7604;
													assign node7604 = (inp[7]) ? node7608 : node7605;
														assign node7605 = (inp[14]) ? 4'b1100 : 4'b1100;
														assign node7608 = (inp[14]) ? 4'b0101 : 4'b1100;
													assign node7611 = (inp[7]) ? 4'b0100 : 4'b0101;
											assign node7614 = (inp[8]) ? node7622 : node7615;
												assign node7615 = (inp[13]) ? 4'b0100 : node7616;
													assign node7616 = (inp[7]) ? node7618 : 4'b1100;
														assign node7618 = (inp[14]) ? 4'b0101 : 4'b0100;
												assign node7622 = (inp[7]) ? node7626 : node7623;
													assign node7623 = (inp[14]) ? 4'b0101 : 4'b0100;
													assign node7626 = (inp[5]) ? 4'b0100 : node7627;
														assign node7627 = (inp[13]) ? 4'b0100 : 4'b0100;
								assign node7631 = (inp[1]) ? node7713 : node7632;
									assign node7632 = (inp[6]) ? node7676 : node7633;
										assign node7633 = (inp[7]) ? node7653 : node7634;
											assign node7634 = (inp[11]) ? node7644 : node7635;
												assign node7635 = (inp[13]) ? node7641 : node7636;
													assign node7636 = (inp[5]) ? node7638 : 4'b1100;
														assign node7638 = (inp[14]) ? 4'b1101 : 4'b1100;
													assign node7641 = (inp[2]) ? 4'b0101 : 4'b1100;
												assign node7644 = (inp[13]) ? 4'b0100 : node7645;
													assign node7645 = (inp[2]) ? node7649 : node7646;
														assign node7646 = (inp[8]) ? 4'b0100 : 4'b0101;
														assign node7649 = (inp[8]) ? 4'b0101 : 4'b0100;
											assign node7653 = (inp[8]) ? node7667 : node7654;
												assign node7654 = (inp[14]) ? node7660 : node7655;
													assign node7655 = (inp[13]) ? 4'b1101 : node7656;
														assign node7656 = (inp[5]) ? 4'b1100 : 4'b0100;
													assign node7660 = (inp[2]) ? node7664 : node7661;
														assign node7661 = (inp[13]) ? 4'b1101 : 4'b0101;
														assign node7664 = (inp[13]) ? 4'b0101 : 4'b1101;
												assign node7667 = (inp[2]) ? node7671 : node7668;
													assign node7668 = (inp[14]) ? 4'b1100 : 4'b1101;
													assign node7671 = (inp[14]) ? 4'b1100 : node7672;
														assign node7672 = (inp[13]) ? 4'b0100 : 4'b1100;
										assign node7676 = (inp[11]) ? node7696 : node7677;
											assign node7677 = (inp[13]) ? node7685 : node7678;
												assign node7678 = (inp[8]) ? node7680 : 4'b0101;
													assign node7680 = (inp[5]) ? node7682 : 4'b0100;
														assign node7682 = (inp[14]) ? 4'b0101 : 4'b0100;
												assign node7685 = (inp[8]) ? node7691 : node7686;
													assign node7686 = (inp[7]) ? node7688 : 4'b0100;
														assign node7688 = (inp[2]) ? 4'b1101 : 4'b0100;
													assign node7691 = (inp[7]) ? node7693 : 4'b1101;
														assign node7693 = (inp[14]) ? 4'b1100 : 4'b1101;
											assign node7696 = (inp[13]) ? node7706 : node7697;
												assign node7697 = (inp[2]) ? node7699 : 4'b1101;
													assign node7699 = (inp[14]) ? node7703 : node7700;
														assign node7700 = (inp[8]) ? 4'b1100 : 4'b1100;
														assign node7703 = (inp[5]) ? 4'b1100 : 4'b1101;
												assign node7706 = (inp[2]) ? 4'b0101 : node7707;
													assign node7707 = (inp[7]) ? node7709 : 4'b1100;
														assign node7709 = (inp[8]) ? 4'b0100 : 4'b0101;
									assign node7713 = (inp[11]) ? node7763 : node7714;
										assign node7714 = (inp[6]) ? node7738 : node7715;
											assign node7715 = (inp[7]) ? node7729 : node7716;
												assign node7716 = (inp[13]) ? node7724 : node7717;
													assign node7717 = (inp[8]) ? node7721 : node7718;
														assign node7718 = (inp[14]) ? 4'b1100 : 4'b1101;
														assign node7721 = (inp[14]) ? 4'b0101 : 4'b1100;
													assign node7724 = (inp[14]) ? 4'b0100 : node7725;
														assign node7725 = (inp[5]) ? 4'b0101 : 4'b0100;
												assign node7729 = (inp[8]) ? node7733 : node7730;
													assign node7730 = (inp[14]) ? 4'b0101 : 4'b0100;
													assign node7733 = (inp[2]) ? 4'b0100 : node7734;
														assign node7734 = (inp[14]) ? 4'b0100 : 4'b0101;
											assign node7738 = (inp[13]) ? node7750 : node7739;
												assign node7739 = (inp[8]) ? node7745 : node7740;
													assign node7740 = (inp[7]) ? node7742 : 4'b0100;
														assign node7742 = (inp[2]) ? 4'b1101 : 4'b0100;
													assign node7745 = (inp[7]) ? 4'b1100 : node7746;
														assign node7746 = (inp[5]) ? 4'b0100 : 4'b1101;
												assign node7750 = (inp[7]) ? node7756 : node7751;
													assign node7751 = (inp[14]) ? node7753 : 4'b1101;
														assign node7753 = (inp[2]) ? 4'b1101 : 4'b1100;
													assign node7756 = (inp[14]) ? node7760 : node7757;
														assign node7757 = (inp[5]) ? 4'b1100 : 4'b1100;
														assign node7760 = (inp[5]) ? 4'b1101 : 4'b1100;
										assign node7763 = (inp[6]) ? node7791 : node7764;
											assign node7764 = (inp[13]) ? node7778 : node7765;
												assign node7765 = (inp[7]) ? node7771 : node7766;
													assign node7766 = (inp[14]) ? node7768 : 4'b0100;
														assign node7768 = (inp[8]) ? 4'b1101 : 4'b0100;
													assign node7771 = (inp[8]) ? node7775 : node7772;
														assign node7772 = (inp[14]) ? 4'b1101 : 4'b0100;
														assign node7775 = (inp[14]) ? 4'b1100 : 4'b1101;
												assign node7778 = (inp[5]) ? node7786 : node7779;
													assign node7779 = (inp[7]) ? node7783 : node7780;
														assign node7780 = (inp[2]) ? 4'b1101 : 4'b1100;
														assign node7783 = (inp[8]) ? 4'b1100 : 4'b1101;
													assign node7786 = (inp[2]) ? 4'b1100 : node7787;
														assign node7787 = (inp[7]) ? 4'b1100 : 4'b1100;
											assign node7791 = (inp[8]) ? node7805 : node7792;
												assign node7792 = (inp[13]) ? node7800 : node7793;
													assign node7793 = (inp[5]) ? node7797 : node7794;
														assign node7794 = (inp[7]) ? 4'b0100 : 4'b1100;
														assign node7797 = (inp[7]) ? 4'b1100 : 4'b1100;
													assign node7800 = (inp[2]) ? 4'b0100 : node7801;
														assign node7801 = (inp[14]) ? 4'b0101 : 4'b0100;
												assign node7805 = (inp[7]) ? 4'b0100 : 4'b0101;
						assign node7808 = (inp[10]) ? node8150 : node7809;
							assign node7809 = (inp[12]) ? node7971 : node7810;
								assign node7810 = (inp[11]) ? node7896 : node7811;
									assign node7811 = (inp[8]) ? node7851 : node7812;
										assign node7812 = (inp[7]) ? node7830 : node7813;
											assign node7813 = (inp[6]) ? node7819 : node7814;
												assign node7814 = (inp[13]) ? 4'b1100 : node7815;
													assign node7815 = (inp[1]) ? 4'b1100 : 4'b1101;
												assign node7819 = (inp[14]) ? node7825 : node7820;
													assign node7820 = (inp[13]) ? 4'b1101 : node7821;
														assign node7821 = (inp[2]) ? 4'b0100 : 4'b0101;
													assign node7825 = (inp[5]) ? 4'b0100 : node7826;
														assign node7826 = (inp[2]) ? 4'b1100 : 4'b0100;
											assign node7830 = (inp[6]) ? node7842 : node7831;
												assign node7831 = (inp[1]) ? node7837 : node7832;
													assign node7832 = (inp[14]) ? 4'b0101 : node7833;
														assign node7833 = (inp[5]) ? 4'b1100 : 4'b1101;
													assign node7837 = (inp[14]) ? 4'b0101 : node7838;
														assign node7838 = (inp[2]) ? 4'b0101 : 4'b0100;
												assign node7842 = (inp[13]) ? node7846 : node7843;
													assign node7843 = (inp[1]) ? 4'b1101 : 4'b0101;
													assign node7846 = (inp[2]) ? 4'b1101 : node7847;
														assign node7847 = (inp[5]) ? 4'b1100 : 4'b1101;
										assign node7851 = (inp[7]) ? node7873 : node7852;
											assign node7852 = (inp[14]) ? node7864 : node7853;
												assign node7853 = (inp[2]) ? node7861 : node7854;
													assign node7854 = (inp[6]) ? node7858 : node7855;
														assign node7855 = (inp[13]) ? 4'b0100 : 4'b1100;
														assign node7858 = (inp[13]) ? 4'b0100 : 4'b0100;
													assign node7861 = (inp[6]) ? 4'b1101 : 4'b0101;
												assign node7864 = (inp[13]) ? node7870 : node7865;
													assign node7865 = (inp[2]) ? node7867 : 4'b1101;
														assign node7867 = (inp[6]) ? 4'b0101 : 4'b1101;
													assign node7870 = (inp[6]) ? 4'b1101 : 4'b0101;
											assign node7873 = (inp[6]) ? node7883 : node7874;
												assign node7874 = (inp[13]) ? node7878 : node7875;
													assign node7875 = (inp[1]) ? 4'b0100 : 4'b1100;
													assign node7878 = (inp[2]) ? 4'b0100 : node7879;
														assign node7879 = (inp[14]) ? 4'b0100 : 4'b0101;
												assign node7883 = (inp[13]) ? node7891 : node7884;
													assign node7884 = (inp[1]) ? node7888 : node7885;
														assign node7885 = (inp[14]) ? 4'b0100 : 4'b0101;
														assign node7888 = (inp[5]) ? 4'b1100 : 4'b1100;
													assign node7891 = (inp[14]) ? 4'b1100 : node7892;
														assign node7892 = (inp[2]) ? 4'b1100 : 4'b1101;
									assign node7896 = (inp[6]) ? node7940 : node7897;
										assign node7897 = (inp[1]) ? node7919 : node7898;
											assign node7898 = (inp[13]) ? node7906 : node7899;
												assign node7899 = (inp[7]) ? node7903 : node7900;
													assign node7900 = (inp[8]) ? 4'b0101 : 4'b0100;
													assign node7903 = (inp[8]) ? 4'b0100 : 4'b0101;
												assign node7906 = (inp[14]) ? node7914 : node7907;
													assign node7907 = (inp[2]) ? node7911 : node7908;
														assign node7908 = (inp[8]) ? 4'b0100 : 4'b0101;
														assign node7911 = (inp[8]) ? 4'b1101 : 4'b0100;
													assign node7914 = (inp[8]) ? node7916 : 4'b1101;
														assign node7916 = (inp[7]) ? 4'b1100 : 4'b1101;
											assign node7919 = (inp[7]) ? node7933 : node7920;
												assign node7920 = (inp[8]) ? node7928 : node7921;
													assign node7921 = (inp[13]) ? node7925 : node7922;
														assign node7922 = (inp[5]) ? 4'b0101 : 4'b0100;
														assign node7925 = (inp[2]) ? 4'b1100 : 4'b1100;
													assign node7928 = (inp[2]) ? 4'b1101 : node7929;
														assign node7929 = (inp[14]) ? 4'b1101 : 4'b0100;
												assign node7933 = (inp[8]) ? node7935 : 4'b1101;
													assign node7935 = (inp[14]) ? 4'b1100 : node7936;
														assign node7936 = (inp[2]) ? 4'b1100 : 4'b1101;
										assign node7940 = (inp[1]) ? node7956 : node7941;
											assign node7941 = (inp[13]) ? node7949 : node7942;
												assign node7942 = (inp[2]) ? 4'b1101 : node7943;
													assign node7943 = (inp[5]) ? 4'b1101 : node7944;
														assign node7944 = (inp[7]) ? 4'b1100 : 4'b1101;
												assign node7949 = (inp[8]) ? node7951 : 4'b1100;
													assign node7951 = (inp[7]) ? 4'b0100 : node7952;
														assign node7952 = (inp[2]) ? 4'b0101 : 4'b0100;
											assign node7956 = (inp[7]) ? node7966 : node7957;
												assign node7957 = (inp[8]) ? node7961 : node7958;
													assign node7958 = (inp[13]) ? 4'b0100 : 4'b1100;
													assign node7961 = (inp[14]) ? 4'b0101 : node7962;
														assign node7962 = (inp[2]) ? 4'b0101 : 4'b0100;
												assign node7966 = (inp[8]) ? node7968 : 4'b0101;
													assign node7968 = (inp[2]) ? 4'b0100 : 4'b0101;
								assign node7971 = (inp[11]) ? node8055 : node7972;
									assign node7972 = (inp[6]) ? node8014 : node7973;
										assign node7973 = (inp[1]) ? node7993 : node7974;
											assign node7974 = (inp[13]) ? node7982 : node7975;
												assign node7975 = (inp[8]) ? node7977 : 4'b1100;
													assign node7977 = (inp[2]) ? 4'b1101 : node7978;
														assign node7978 = (inp[5]) ? 4'b1101 : 4'b1100;
												assign node7982 = (inp[8]) ? node7990 : node7983;
													assign node7983 = (inp[7]) ? node7987 : node7984;
														assign node7984 = (inp[14]) ? 4'b1100 : 4'b1100;
														assign node7987 = (inp[2]) ? 4'b0101 : 4'b0100;
													assign node7990 = (inp[7]) ? 4'b0100 : 4'b0101;
											assign node7993 = (inp[13]) ? node8003 : node7994;
												assign node7994 = (inp[8]) ? node7998 : node7995;
													assign node7995 = (inp[7]) ? 4'b0101 : 4'b1100;
													assign node7998 = (inp[14]) ? node8000 : 4'b0101;
														assign node8000 = (inp[7]) ? 4'b0100 : 4'b0101;
												assign node8003 = (inp[5]) ? node8009 : node8004;
													assign node8004 = (inp[2]) ? node8006 : 4'b0101;
														assign node8006 = (inp[7]) ? 4'b0100 : 4'b0101;
													assign node8009 = (inp[8]) ? 4'b0100 : node8010;
														assign node8010 = (inp[2]) ? 4'b0100 : 4'b0100;
										assign node8014 = (inp[13]) ? node8034 : node8015;
											assign node8015 = (inp[5]) ? node8027 : node8016;
												assign node8016 = (inp[1]) ? node8022 : node8017;
													assign node8017 = (inp[8]) ? 4'b0101 : node8018;
														assign node8018 = (inp[7]) ? 4'b0101 : 4'b0100;
													assign node8022 = (inp[2]) ? 4'b1000 : node8023;
														assign node8023 = (inp[8]) ? 4'b0100 : 4'b0101;
												assign node8027 = (inp[7]) ? node8029 : 4'b0100;
													assign node8029 = (inp[14]) ? node8031 : 4'b0100;
														assign node8031 = (inp[2]) ? 4'b0100 : 4'b0101;
											assign node8034 = (inp[1]) ? node8046 : node8035;
												assign node8035 = (inp[7]) ? node8043 : node8036;
													assign node8036 = (inp[8]) ? node8040 : node8037;
														assign node8037 = (inp[2]) ? 4'b0100 : 4'b0101;
														assign node8040 = (inp[2]) ? 4'b1001 : 4'b0000;
													assign node8043 = (inp[8]) ? 4'b1000 : 4'b1001;
												assign node8046 = (inp[7]) ? node8050 : node8047;
													assign node8047 = (inp[8]) ? 4'b1001 : 4'b1000;
													assign node8050 = (inp[8]) ? 4'b1000 : node8051;
														assign node8051 = (inp[2]) ? 4'b1001 : 4'b1000;
									assign node8055 = (inp[6]) ? node8103 : node8056;
										assign node8056 = (inp[1]) ? node8078 : node8057;
											assign node8057 = (inp[13]) ? node8069 : node8058;
												assign node8058 = (inp[5]) ? node8066 : node8059;
													assign node8059 = (inp[2]) ? node8063 : node8060;
														assign node8060 = (inp[7]) ? 4'b0100 : 4'b0100;
														assign node8063 = (inp[14]) ? 4'b0101 : 4'b0100;
													assign node8066 = (inp[7]) ? 4'b0101 : 4'b0100;
												assign node8069 = (inp[8]) ? node8075 : node8070;
													assign node8070 = (inp[2]) ? 4'b0100 : node8071;
														assign node8071 = (inp[7]) ? 4'b0100 : 4'b0101;
													assign node8075 = (inp[7]) ? 4'b1000 : 4'b1001;
											assign node8078 = (inp[13]) ? node8090 : node8079;
												assign node8079 = (inp[8]) ? node8085 : node8080;
													assign node8080 = (inp[7]) ? node8082 : 4'b0100;
														assign node8082 = (inp[5]) ? 4'b0000 : 4'b1001;
													assign node8085 = (inp[7]) ? node8087 : 4'b1001;
														assign node8087 = (inp[14]) ? 4'b1000 : 4'b1000;
												assign node8090 = (inp[14]) ? node8096 : node8091;
													assign node8091 = (inp[8]) ? node8093 : 4'b1001;
														assign node8093 = (inp[5]) ? 4'b1001 : 4'b1000;
													assign node8096 = (inp[7]) ? node8100 : node8097;
														assign node8097 = (inp[8]) ? 4'b1001 : 4'b1000;
														assign node8100 = (inp[8]) ? 4'b1000 : 4'b1001;
										assign node8103 = (inp[1]) ? node8129 : node8104;
											assign node8104 = (inp[13]) ? node8118 : node8105;
												assign node8105 = (inp[8]) ? node8113 : node8106;
													assign node8106 = (inp[7]) ? node8110 : node8107;
														assign node8107 = (inp[2]) ? 4'b1000 : 4'b1001;
														assign node8110 = (inp[14]) ? 4'b1001 : 4'b1000;
													assign node8113 = (inp[7]) ? 4'b1000 : node8114;
														assign node8114 = (inp[2]) ? 4'b1001 : 4'b1000;
												assign node8118 = (inp[7]) ? node8124 : node8119;
													assign node8119 = (inp[8]) ? node8121 : 4'b1000;
														assign node8121 = (inp[14]) ? 4'b0001 : 4'b1000;
													assign node8124 = (inp[14]) ? 4'b0001 : node8125;
														assign node8125 = (inp[8]) ? 4'b0001 : 4'b1000;
											assign node8129 = (inp[2]) ? node8137 : node8130;
												assign node8130 = (inp[13]) ? 4'b0000 : node8131;
													assign node8131 = (inp[14]) ? 4'b0001 : node8132;
														assign node8132 = (inp[8]) ? 4'b1000 : 4'b1000;
												assign node8137 = (inp[13]) ? node8145 : node8138;
													assign node8138 = (inp[5]) ? node8142 : node8139;
														assign node8139 = (inp[14]) ? 4'b0000 : 4'b1000;
														assign node8142 = (inp[8]) ? 4'b0000 : 4'b0001;
													assign node8145 = (inp[5]) ? node8147 : 4'b0001;
														assign node8147 = (inp[7]) ? 4'b0001 : 4'b0000;
							assign node8150 = (inp[12]) ? node8322 : node8151;
								assign node8151 = (inp[6]) ? node8237 : node8152;
									assign node8152 = (inp[11]) ? node8194 : node8153;
										assign node8153 = (inp[13]) ? node8171 : node8154;
											assign node8154 = (inp[1]) ? node8162 : node8155;
												assign node8155 = (inp[2]) ? 4'b1100 : node8156;
													assign node8156 = (inp[5]) ? 4'b1101 : node8157;
														assign node8157 = (inp[7]) ? 4'b1101 : 4'b1100;
												assign node8162 = (inp[7]) ? node8168 : node8163;
													assign node8163 = (inp[8]) ? node8165 : 4'b1100;
														assign node8165 = (inp[2]) ? 4'b0101 : 4'b0100;
													assign node8168 = (inp[5]) ? 4'b0101 : 4'b0100;
											assign node8171 = (inp[5]) ? node8181 : node8172;
												assign node8172 = (inp[14]) ? node8176 : node8173;
													assign node8173 = (inp[7]) ? 4'b0101 : 4'b1101;
													assign node8176 = (inp[1]) ? 4'b0100 : node8177;
														assign node8177 = (inp[2]) ? 4'b0100 : 4'b0101;
												assign node8181 = (inp[7]) ? node8189 : node8182;
													assign node8182 = (inp[8]) ? node8186 : node8183;
														assign node8183 = (inp[1]) ? 4'b0100 : 4'b1100;
														assign node8186 = (inp[14]) ? 4'b0101 : 4'b0100;
													assign node8189 = (inp[14]) ? 4'b0100 : node8190;
														assign node8190 = (inp[1]) ? 4'b0100 : 4'b0101;
										assign node8194 = (inp[1]) ? node8214 : node8195;
											assign node8195 = (inp[13]) ? node8209 : node8196;
												assign node8196 = (inp[14]) ? node8204 : node8197;
													assign node8197 = (inp[2]) ? node8201 : node8198;
														assign node8198 = (inp[8]) ? 4'b0100 : 4'b0100;
														assign node8201 = (inp[7]) ? 4'b0101 : 4'b0100;
													assign node8204 = (inp[8]) ? 4'b0100 : node8205;
														assign node8205 = (inp[7]) ? 4'b0101 : 4'b0100;
												assign node8209 = (inp[14]) ? node8211 : 4'b0100;
													assign node8211 = (inp[8]) ? 4'b1000 : 4'b1001;
											assign node8214 = (inp[14]) ? node8228 : node8215;
												assign node8215 = (inp[13]) ? node8221 : node8216;
													assign node8216 = (inp[7]) ? 4'b1001 : node8217;
														assign node8217 = (inp[2]) ? 4'b0000 : 4'b0100;
													assign node8221 = (inp[5]) ? node8225 : node8222;
														assign node8222 = (inp[7]) ? 4'b1000 : 4'b1001;
														assign node8225 = (inp[2]) ? 4'b1000 : 4'b1001;
												assign node8228 = (inp[2]) ? node8230 : 4'b1001;
													assign node8230 = (inp[7]) ? node8234 : node8231;
														assign node8231 = (inp[8]) ? 4'b1001 : 4'b1000;
														assign node8234 = (inp[8]) ? 4'b1000 : 4'b1001;
									assign node8237 = (inp[11]) ? node8283 : node8238;
										assign node8238 = (inp[13]) ? node8264 : node8239;
											assign node8239 = (inp[1]) ? node8253 : node8240;
												assign node8240 = (inp[7]) ? node8248 : node8241;
													assign node8241 = (inp[14]) ? node8245 : node8242;
														assign node8242 = (inp[8]) ? 4'b0100 : 4'b0101;
														assign node8245 = (inp[8]) ? 4'b0101 : 4'b0100;
													assign node8248 = (inp[5]) ? node8250 : 4'b0100;
														assign node8250 = (inp[2]) ? 4'b0101 : 4'b0100;
												assign node8253 = (inp[7]) ? node8261 : node8254;
													assign node8254 = (inp[2]) ? node8258 : node8255;
														assign node8255 = (inp[14]) ? 4'b0100 : 4'b0100;
														assign node8258 = (inp[8]) ? 4'b1001 : 4'b0100;
													assign node8261 = (inp[8]) ? 4'b1000 : 4'b1001;
											assign node8264 = (inp[8]) ? node8274 : node8265;
												assign node8265 = (inp[7]) ? node8269 : node8266;
													assign node8266 = (inp[1]) ? 4'b1000 : 4'b0100;
													assign node8269 = (inp[2]) ? 4'b1001 : node8270;
														assign node8270 = (inp[14]) ? 4'b1001 : 4'b0000;
												assign node8274 = (inp[7]) ? node8280 : node8275;
													assign node8275 = (inp[14]) ? 4'b1001 : node8276;
														assign node8276 = (inp[2]) ? 4'b1001 : 4'b1000;
													assign node8280 = (inp[14]) ? 4'b1000 : 4'b1001;
										assign node8283 = (inp[1]) ? node8303 : node8284;
											assign node8284 = (inp[13]) ? node8296 : node8285;
												assign node8285 = (inp[14]) ? node8291 : node8286;
													assign node8286 = (inp[2]) ? node8288 : 4'b1001;
														assign node8288 = (inp[7]) ? 4'b1000 : 4'b1001;
													assign node8291 = (inp[2]) ? 4'b1000 : node8292;
														assign node8292 = (inp[7]) ? 4'b1001 : 4'b1000;
												assign node8296 = (inp[14]) ? node8298 : 4'b1000;
													assign node8298 = (inp[7]) ? node8300 : 4'b0001;
														assign node8300 = (inp[8]) ? 4'b0000 : 4'b0001;
											assign node8303 = (inp[8]) ? node8311 : node8304;
												assign node8304 = (inp[7]) ? node8306 : 4'b0000;
													assign node8306 = (inp[2]) ? 4'b0001 : node8307;
														assign node8307 = (inp[14]) ? 4'b0001 : 4'b0000;
												assign node8311 = (inp[7]) ? node8317 : node8312;
													assign node8312 = (inp[2]) ? 4'b0001 : node8313;
														assign node8313 = (inp[14]) ? 4'b0001 : 4'b1000;
													assign node8317 = (inp[2]) ? 4'b0000 : node8318;
														assign node8318 = (inp[14]) ? 4'b0000 : 4'b0001;
								assign node8322 = (inp[7]) ? node8406 : node8323;
									assign node8323 = (inp[8]) ? node8357 : node8324;
										assign node8324 = (inp[2]) ? node8346 : node8325;
											assign node8325 = (inp[14]) ? node8337 : node8326;
												assign node8326 = (inp[11]) ? node8332 : node8327;
													assign node8327 = (inp[6]) ? 4'b0001 : node8328;
														assign node8328 = (inp[13]) ? 4'b0001 : 4'b1001;
													assign node8332 = (inp[6]) ? node8334 : 4'b0001;
														assign node8334 = (inp[1]) ? 4'b0001 : 4'b1001;
												assign node8337 = (inp[5]) ? node8341 : node8338;
													assign node8338 = (inp[11]) ? 4'b0000 : 4'b1000;
													assign node8341 = (inp[11]) ? 4'b1000 : node8342;
														assign node8342 = (inp[6]) ? 4'b0000 : 4'b1000;
											assign node8346 = (inp[6]) ? node8352 : node8347;
												assign node8347 = (inp[11]) ? 4'b0000 : node8348;
													assign node8348 = (inp[13]) ? 4'b0000 : 4'b1000;
												assign node8352 = (inp[11]) ? 4'b1000 : node8353;
													assign node8353 = (inp[13]) ? 4'b1000 : 4'b0000;
										assign node8357 = (inp[14]) ? node8377 : node8358;
											assign node8358 = (inp[2]) ? node8366 : node8359;
												assign node8359 = (inp[5]) ? 4'b1000 : node8360;
													assign node8360 = (inp[11]) ? node8362 : 4'b0000;
														assign node8362 = (inp[13]) ? 4'b0000 : 4'b1000;
												assign node8366 = (inp[13]) ? node8372 : node8367;
													assign node8367 = (inp[1]) ? node8369 : 4'b0001;
														assign node8369 = (inp[5]) ? 4'b0001 : 4'b1001;
													assign node8372 = (inp[1]) ? node8374 : 4'b1001;
														assign node8374 = (inp[5]) ? 4'b1001 : 4'b0001;
											assign node8377 = (inp[2]) ? node8393 : node8378;
												assign node8378 = (inp[13]) ? node8386 : node8379;
													assign node8379 = (inp[6]) ? node8383 : node8380;
														assign node8380 = (inp[5]) ? 4'b1001 : 4'b0001;
														assign node8383 = (inp[11]) ? 4'b1001 : 4'b1001;
													assign node8386 = (inp[5]) ? node8390 : node8387;
														assign node8387 = (inp[6]) ? 4'b1001 : 4'b0001;
														assign node8390 = (inp[11]) ? 4'b0001 : 4'b0001;
												assign node8393 = (inp[5]) ? node8401 : node8394;
													assign node8394 = (inp[13]) ? node8398 : node8395;
														assign node8395 = (inp[6]) ? 4'b0001 : 4'b0001;
														assign node8398 = (inp[1]) ? 4'b1001 : 4'b0001;
													assign node8401 = (inp[13]) ? 4'b0001 : node8402;
														assign node8402 = (inp[1]) ? 4'b0001 : 4'b0001;
									assign node8406 = (inp[8]) ? node8434 : node8407;
										assign node8407 = (inp[14]) ? node8425 : node8408;
											assign node8408 = (inp[2]) ? node8420 : node8409;
												assign node8409 = (inp[13]) ? node8415 : node8410;
													assign node8410 = (inp[1]) ? node8412 : 4'b1000;
														assign node8412 = (inp[5]) ? 4'b0000 : 4'b1000;
													assign node8415 = (inp[6]) ? 4'b0000 : node8416;
														assign node8416 = (inp[5]) ? 4'b0000 : 4'b0000;
												assign node8420 = (inp[11]) ? 4'b1001 : node8421;
													assign node8421 = (inp[6]) ? 4'b1001 : 4'b0001;
											assign node8425 = (inp[1]) ? 4'b1001 : node8426;
												assign node8426 = (inp[11]) ? 4'b0001 : node8427;
													assign node8427 = (inp[6]) ? 4'b0001 : node8428;
														assign node8428 = (inp[13]) ? 4'b0001 : 4'b1001;
										assign node8434 = (inp[2]) ? node8454 : node8435;
											assign node8435 = (inp[14]) ? node8445 : node8436;
												assign node8436 = (inp[11]) ? node8442 : node8437;
													assign node8437 = (inp[6]) ? 4'b1001 : node8438;
														assign node8438 = (inp[5]) ? 4'b1001 : 4'b0001;
													assign node8442 = (inp[6]) ? 4'b0001 : 4'b1001;
												assign node8445 = (inp[1]) ? node8447 : 4'b1000;
													assign node8447 = (inp[6]) ? node8451 : node8448;
														assign node8448 = (inp[11]) ? 4'b1000 : 4'b0000;
														assign node8451 = (inp[13]) ? 4'b1000 : 4'b0000;
											assign node8454 = (inp[11]) ? node8464 : node8455;
												assign node8455 = (inp[6]) ? node8461 : node8456;
													assign node8456 = (inp[1]) ? 4'b0000 : node8457;
														assign node8457 = (inp[13]) ? 4'b0000 : 4'b1000;
													assign node8461 = (inp[1]) ? 4'b1000 : 4'b0000;
												assign node8464 = (inp[14]) ? node8470 : node8465;
													assign node8465 = (inp[5]) ? 4'b0000 : node8466;
														assign node8466 = (inp[13]) ? 4'b1000 : 4'b0000;
													assign node8470 = (inp[6]) ? node8474 : node8471;
														assign node8471 = (inp[13]) ? 4'b1000 : 4'b0000;
														assign node8474 = (inp[13]) ? 4'b0000 : 4'b1000;
				assign node8477 = (inp[3]) ? node9875 : node8478;
					assign node8478 = (inp[5]) ? node9160 : node8479;
						assign node8479 = (inp[9]) ? node8797 : node8480;
							assign node8480 = (inp[10]) ? node8640 : node8481;
								assign node8481 = (inp[12]) ? node8553 : node8482;
									assign node8482 = (inp[8]) ? node8524 : node8483;
										assign node8483 = (inp[7]) ? node8505 : node8484;
											assign node8484 = (inp[2]) ? node8496 : node8485;
												assign node8485 = (inp[14]) ? node8491 : node8486;
													assign node8486 = (inp[13]) ? 4'b0001 : node8487;
														assign node8487 = (inp[11]) ? 4'b0001 : 4'b1001;
													assign node8491 = (inp[11]) ? 4'b0000 : node8492;
														assign node8492 = (inp[13]) ? 4'b1000 : 4'b0000;
												assign node8496 = (inp[13]) ? 4'b1000 : node8497;
													assign node8497 = (inp[14]) ? node8501 : node8498;
														assign node8498 = (inp[1]) ? 4'b0000 : 4'b0000;
														assign node8501 = (inp[6]) ? 4'b1000 : 4'b0000;
											assign node8505 = (inp[14]) ? node8517 : node8506;
												assign node8506 = (inp[2]) ? node8512 : node8507;
													assign node8507 = (inp[6]) ? 4'b0000 : node8508;
														assign node8508 = (inp[13]) ? 4'b1000 : 4'b0000;
													assign node8512 = (inp[11]) ? 4'b0001 : node8513;
														assign node8513 = (inp[6]) ? 4'b1001 : 4'b0001;
												assign node8517 = (inp[2]) ? 4'b0001 : node8518;
													assign node8518 = (inp[1]) ? 4'b1001 : node8519;
														assign node8519 = (inp[13]) ? 4'b1001 : 4'b0001;
										assign node8524 = (inp[7]) ? node8542 : node8525;
											assign node8525 = (inp[2]) ? node8529 : node8526;
												assign node8526 = (inp[14]) ? 4'b1001 : 4'b1000;
												assign node8529 = (inp[14]) ? node8535 : node8530;
													assign node8530 = (inp[11]) ? 4'b1001 : node8531;
														assign node8531 = (inp[1]) ? 4'b1001 : 4'b0001;
													assign node8535 = (inp[1]) ? node8539 : node8536;
														assign node8536 = (inp[6]) ? 4'b0001 : 4'b0001;
														assign node8539 = (inp[13]) ? 4'b1001 : 4'b0001;
											assign node8542 = (inp[2]) ? node8548 : node8543;
												assign node8543 = (inp[14]) ? 4'b1000 : node8544;
													assign node8544 = (inp[1]) ? 4'b0001 : 4'b1001;
												assign node8548 = (inp[6]) ? node8550 : 4'b0000;
													assign node8550 = (inp[11]) ? 4'b0000 : 4'b1000;
									assign node8553 = (inp[11]) ? node8595 : node8554;
										assign node8554 = (inp[6]) ? node8578 : node8555;
											assign node8555 = (inp[13]) ? node8567 : node8556;
												assign node8556 = (inp[1]) ? node8562 : node8557;
													assign node8557 = (inp[7]) ? 4'b1000 : node8558;
														assign node8558 = (inp[14]) ? 4'b1001 : 4'b1000;
													assign node8562 = (inp[14]) ? node8564 : 4'b1000;
														assign node8564 = (inp[2]) ? 4'b0001 : 4'b0000;
												assign node8567 = (inp[1]) ? node8573 : node8568;
													assign node8568 = (inp[7]) ? 4'b0001 : node8569;
														assign node8569 = (inp[8]) ? 4'b0001 : 4'b1000;
													assign node8573 = (inp[8]) ? node8575 : 4'b0001;
														assign node8575 = (inp[7]) ? 4'b0000 : 4'b0001;
											assign node8578 = (inp[1]) ? node8588 : node8579;
												assign node8579 = (inp[13]) ? node8585 : node8580;
													assign node8580 = (inp[8]) ? 4'b0001 : node8581;
														assign node8581 = (inp[7]) ? 4'b0000 : 4'b0001;
													assign node8585 = (inp[7]) ? 4'b1101 : 4'b0000;
												assign node8588 = (inp[7]) ? node8590 : 4'b1101;
													assign node8590 = (inp[8]) ? 4'b1100 : node8591;
														assign node8591 = (inp[2]) ? 4'b1101 : 4'b0000;
										assign node8595 = (inp[6]) ? node8623 : node8596;
											assign node8596 = (inp[13]) ? node8612 : node8597;
												assign node8597 = (inp[1]) ? node8605 : node8598;
													assign node8598 = (inp[14]) ? node8602 : node8599;
														assign node8599 = (inp[8]) ? 4'b0001 : 4'b0000;
														assign node8602 = (inp[8]) ? 4'b0000 : 4'b0001;
													assign node8605 = (inp[7]) ? node8609 : node8606;
														assign node8606 = (inp[14]) ? 4'b1101 : 4'b0000;
														assign node8609 = (inp[8]) ? 4'b1100 : 4'b1101;
												assign node8612 = (inp[7]) ? node8618 : node8613;
													assign node8613 = (inp[14]) ? node8615 : 4'b1101;
														assign node8615 = (inp[8]) ? 4'b1101 : 4'b1100;
													assign node8618 = (inp[1]) ? 4'b1100 : node8619;
														assign node8619 = (inp[14]) ? 4'b1100 : 4'b1101;
											assign node8623 = (inp[13]) ? node8633 : node8624;
												assign node8624 = (inp[1]) ? node8630 : node8625;
													assign node8625 = (inp[2]) ? node8627 : 4'b1101;
														assign node8627 = (inp[8]) ? 4'b1100 : 4'b1101;
													assign node8630 = (inp[14]) ? 4'b0100 : 4'b1100;
												assign node8633 = (inp[8]) ? node8635 : 4'b0101;
													assign node8635 = (inp[7]) ? node8637 : 4'b0101;
														assign node8637 = (inp[2]) ? 4'b0100 : 4'b0101;
								assign node8640 = (inp[12]) ? node8714 : node8641;
									assign node8641 = (inp[6]) ? node8681 : node8642;
										assign node8642 = (inp[11]) ? node8658 : node8643;
											assign node8643 = (inp[1]) ? node8649 : node8644;
												assign node8644 = (inp[8]) ? node8646 : 4'b1000;
													assign node8646 = (inp[7]) ? 4'b1000 : 4'b1001;
												assign node8649 = (inp[2]) ? node8653 : node8650;
													assign node8650 = (inp[13]) ? 4'b0000 : 4'b1000;
													assign node8653 = (inp[8]) ? node8655 : 4'b0001;
														assign node8655 = (inp[7]) ? 4'b0000 : 4'b0001;
											assign node8658 = (inp[1]) ? node8672 : node8659;
												assign node8659 = (inp[13]) ? node8665 : node8660;
													assign node8660 = (inp[7]) ? 4'b0001 : node8661;
														assign node8661 = (inp[8]) ? 4'b0001 : 4'b0000;
													assign node8665 = (inp[8]) ? node8669 : node8666;
														assign node8666 = (inp[7]) ? 4'b1101 : 4'b0000;
														assign node8669 = (inp[7]) ? 4'b1100 : 4'b1101;
												assign node8672 = (inp[14]) ? node8678 : node8673;
													assign node8673 = (inp[2]) ? 4'b1101 : node8674;
														assign node8674 = (inp[8]) ? 4'b0000 : 4'b0001;
													assign node8678 = (inp[8]) ? 4'b1101 : 4'b1100;
										assign node8681 = (inp[11]) ? node8701 : node8682;
											assign node8682 = (inp[1]) ? node8692 : node8683;
												assign node8683 = (inp[7]) ? node8685 : 4'b0000;
													assign node8685 = (inp[13]) ? node8689 : node8686;
														assign node8686 = (inp[8]) ? 4'b0000 : 4'b0001;
														assign node8689 = (inp[8]) ? 4'b1100 : 4'b1101;
												assign node8692 = (inp[13]) ? node8696 : node8693;
													assign node8693 = (inp[8]) ? 4'b1100 : 4'b0000;
													assign node8696 = (inp[7]) ? node8698 : 4'b1101;
														assign node8698 = (inp[8]) ? 4'b1100 : 4'b1101;
											assign node8701 = (inp[1]) ? node8705 : node8702;
												assign node8702 = (inp[2]) ? 4'b0101 : 4'b1101;
												assign node8705 = (inp[13]) ? node8709 : node8706;
													assign node8706 = (inp[8]) ? 4'b0100 : 4'b1100;
													assign node8709 = (inp[8]) ? 4'b0100 : node8710;
														assign node8710 = (inp[7]) ? 4'b0100 : 4'b0100;
									assign node8714 = (inp[7]) ? node8754 : node8715;
										assign node8715 = (inp[8]) ? node8729 : node8716;
											assign node8716 = (inp[14]) ? node8724 : node8717;
												assign node8717 = (inp[2]) ? 4'b1100 : node8718;
													assign node8718 = (inp[13]) ? 4'b0101 : node8719;
														assign node8719 = (inp[11]) ? 4'b0101 : 4'b1101;
												assign node8724 = (inp[6]) ? node8726 : 4'b0100;
													assign node8726 = (inp[13]) ? 4'b1100 : 4'b0100;
											assign node8729 = (inp[11]) ? node8743 : node8730;
												assign node8730 = (inp[14]) ? node8738 : node8731;
													assign node8731 = (inp[2]) ? node8735 : node8732;
														assign node8732 = (inp[1]) ? 4'b0100 : 4'b1100;
														assign node8735 = (inp[1]) ? 4'b0101 : 4'b0101;
													assign node8738 = (inp[6]) ? node8740 : 4'b0101;
														assign node8740 = (inp[2]) ? 4'b0101 : 4'b1101;
												assign node8743 = (inp[6]) ? node8749 : node8744;
													assign node8744 = (inp[14]) ? 4'b1101 : node8745;
														assign node8745 = (inp[2]) ? 4'b1101 : 4'b1100;
													assign node8749 = (inp[1]) ? node8751 : 4'b1101;
														assign node8751 = (inp[14]) ? 4'b0101 : 4'b0100;
										assign node8754 = (inp[8]) ? node8778 : node8755;
											assign node8755 = (inp[14]) ? node8767 : node8756;
												assign node8756 = (inp[2]) ? node8762 : node8757;
													assign node8757 = (inp[13]) ? node8759 : 4'b1100;
														assign node8759 = (inp[6]) ? 4'b0100 : 4'b1100;
													assign node8762 = (inp[1]) ? 4'b1101 : node8763;
														assign node8763 = (inp[6]) ? 4'b1101 : 4'b0101;
												assign node8767 = (inp[2]) ? node8773 : node8768;
													assign node8768 = (inp[11]) ? node8770 : 4'b0101;
														assign node8770 = (inp[1]) ? 4'b0101 : 4'b0101;
													assign node8773 = (inp[13]) ? node8775 : 4'b1101;
														assign node8775 = (inp[1]) ? 4'b1101 : 4'b0101;
											assign node8778 = (inp[2]) ? node8790 : node8779;
												assign node8779 = (inp[14]) ? node8785 : node8780;
													assign node8780 = (inp[13]) ? node8782 : 4'b0101;
														assign node8782 = (inp[11]) ? 4'b0101 : 4'b1101;
													assign node8785 = (inp[6]) ? 4'b1100 : node8786;
														assign node8786 = (inp[13]) ? 4'b0100 : 4'b0100;
												assign node8790 = (inp[1]) ? 4'b0100 : node8791;
													assign node8791 = (inp[11]) ? node8793 : 4'b0100;
														assign node8793 = (inp[6]) ? 4'b1100 : 4'b0100;
							assign node8797 = (inp[10]) ? node8967 : node8798;
								assign node8798 = (inp[12]) ? node8878 : node8799;
									assign node8799 = (inp[8]) ? node8839 : node8800;
										assign node8800 = (inp[7]) ? node8816 : node8801;
											assign node8801 = (inp[2]) ? node8809 : node8802;
												assign node8802 = (inp[14]) ? 4'b1100 : node8803;
													assign node8803 = (inp[6]) ? node8805 : 4'b1101;
														assign node8805 = (inp[1]) ? 4'b0101 : 4'b1101;
												assign node8809 = (inp[13]) ? 4'b1100 : node8810;
													assign node8810 = (inp[6]) ? 4'b1100 : node8811;
														assign node8811 = (inp[11]) ? 4'b0100 : 4'b1100;
											assign node8816 = (inp[14]) ? node8828 : node8817;
												assign node8817 = (inp[2]) ? node8823 : node8818;
													assign node8818 = (inp[1]) ? node8820 : 4'b1100;
														assign node8820 = (inp[11]) ? 4'b1100 : 4'b0100;
													assign node8823 = (inp[1]) ? 4'b1101 : node8824;
														assign node8824 = (inp[6]) ? 4'b0101 : 4'b1101;
												assign node8828 = (inp[11]) ? node8836 : node8829;
													assign node8829 = (inp[6]) ? node8833 : node8830;
														assign node8830 = (inp[1]) ? 4'b0101 : 4'b1101;
														assign node8833 = (inp[2]) ? 4'b1101 : 4'b1101;
													assign node8836 = (inp[6]) ? 4'b0101 : 4'b1101;
										assign node8839 = (inp[7]) ? node8859 : node8840;
											assign node8840 = (inp[2]) ? node8848 : node8841;
												assign node8841 = (inp[14]) ? node8845 : node8842;
													assign node8842 = (inp[6]) ? 4'b1100 : 4'b0100;
													assign node8845 = (inp[13]) ? 4'b1101 : 4'b0101;
												assign node8848 = (inp[6]) ? node8854 : node8849;
													assign node8849 = (inp[1]) ? node8851 : 4'b0101;
														assign node8851 = (inp[11]) ? 4'b1101 : 4'b0101;
													assign node8854 = (inp[13]) ? 4'b1101 : node8855;
														assign node8855 = (inp[14]) ? 4'b0101 : 4'b0101;
											assign node8859 = (inp[14]) ? node8871 : node8860;
												assign node8860 = (inp[2]) ? node8866 : node8861;
													assign node8861 = (inp[13]) ? node8863 : 4'b0101;
														assign node8863 = (inp[11]) ? 4'b0101 : 4'b0101;
													assign node8866 = (inp[13]) ? 4'b0100 : node8867;
														assign node8867 = (inp[6]) ? 4'b1100 : 4'b0100;
												assign node8871 = (inp[13]) ? 4'b1100 : node8872;
													assign node8872 = (inp[2]) ? 4'b0100 : node8873;
														assign node8873 = (inp[6]) ? 4'b0100 : 4'b1100;
									assign node8878 = (inp[6]) ? node8920 : node8879;
										assign node8879 = (inp[11]) ? node8901 : node8880;
											assign node8880 = (inp[13]) ? node8892 : node8881;
												assign node8881 = (inp[1]) ? node8887 : node8882;
													assign node8882 = (inp[7]) ? node8884 : 4'b1101;
														assign node8884 = (inp[2]) ? 4'b1101 : 4'b1100;
													assign node8887 = (inp[7]) ? node8889 : 4'b1100;
														assign node8889 = (inp[8]) ? 4'b0100 : 4'b0101;
												assign node8892 = (inp[1]) ? node8898 : node8893;
													assign node8893 = (inp[7]) ? node8895 : 4'b1100;
														assign node8895 = (inp[8]) ? 4'b0100 : 4'b0100;
													assign node8898 = (inp[8]) ? 4'b0101 : 4'b0100;
											assign node8901 = (inp[1]) ? node8911 : node8902;
												assign node8902 = (inp[8]) ? node8906 : node8903;
													assign node8903 = (inp[2]) ? 4'b0100 : 4'b0101;
													assign node8906 = (inp[13]) ? node8908 : 4'b0100;
														assign node8908 = (inp[7]) ? 4'b1000 : 4'b1001;
												assign node8911 = (inp[14]) ? 4'b1001 : node8912;
													assign node8912 = (inp[2]) ? node8916 : node8913;
														assign node8913 = (inp[13]) ? 4'b1000 : 4'b0100;
														assign node8916 = (inp[8]) ? 4'b1000 : 4'b1001;
										assign node8920 = (inp[11]) ? node8946 : node8921;
											assign node8921 = (inp[13]) ? node8933 : node8922;
												assign node8922 = (inp[1]) ? node8928 : node8923;
													assign node8923 = (inp[8]) ? 4'b0101 : node8924;
														assign node8924 = (inp[7]) ? 4'b0100 : 4'b0100;
													assign node8928 = (inp[7]) ? node8930 : 4'b0100;
														assign node8930 = (inp[8]) ? 4'b1000 : 4'b1001;
												assign node8933 = (inp[14]) ? node8941 : node8934;
													assign node8934 = (inp[2]) ? node8938 : node8935;
														assign node8935 = (inp[8]) ? 4'b1001 : 4'b1000;
														assign node8938 = (inp[8]) ? 4'b1000 : 4'b1001;
													assign node8941 = (inp[1]) ? node8943 : 4'b1000;
														assign node8943 = (inp[8]) ? 4'b1001 : 4'b1000;
											assign node8946 = (inp[7]) ? node8960 : node8947;
												assign node8947 = (inp[8]) ? node8955 : node8948;
													assign node8948 = (inp[13]) ? node8952 : node8949;
														assign node8949 = (inp[14]) ? 4'b1000 : 4'b1000;
														assign node8952 = (inp[1]) ? 4'b0000 : 4'b1000;
													assign node8955 = (inp[1]) ? 4'b0001 : node8956;
														assign node8956 = (inp[13]) ? 4'b0000 : 4'b1001;
												assign node8960 = (inp[8]) ? node8962 : 4'b0001;
													assign node8962 = (inp[14]) ? node8964 : 4'b0001;
														assign node8964 = (inp[13]) ? 4'b0000 : 4'b1000;
								assign node8967 = (inp[12]) ? node9065 : node8968;
									assign node8968 = (inp[6]) ? node9022 : node8969;
										assign node8969 = (inp[11]) ? node8997 : node8970;
											assign node8970 = (inp[7]) ? node8984 : node8971;
												assign node8971 = (inp[14]) ? node8977 : node8972;
													assign node8972 = (inp[2]) ? node8974 : 4'b1100;
														assign node8974 = (inp[13]) ? 4'b1100 : 4'b1101;
													assign node8977 = (inp[8]) ? node8981 : node8978;
														assign node8978 = (inp[13]) ? 4'b0100 : 4'b1100;
														assign node8981 = (inp[1]) ? 4'b0101 : 4'b0101;
												assign node8984 = (inp[2]) ? node8992 : node8985;
													assign node8985 = (inp[1]) ? node8989 : node8986;
														assign node8986 = (inp[13]) ? 4'b0101 : 4'b1101;
														assign node8989 = (inp[8]) ? 4'b0100 : 4'b0101;
													assign node8992 = (inp[1]) ? 4'b0100 : node8993;
														assign node8993 = (inp[13]) ? 4'b0100 : 4'b1100;
											assign node8997 = (inp[1]) ? node9009 : node8998;
												assign node8998 = (inp[7]) ? node9006 : node8999;
													assign node8999 = (inp[14]) ? node9003 : node9000;
														assign node9000 = (inp[2]) ? 4'b0101 : 4'b0100;
														assign node9003 = (inp[8]) ? 4'b1001 : 4'b0100;
													assign node9006 = (inp[2]) ? 4'b0101 : 4'b1001;
												assign node9009 = (inp[13]) ? node9015 : node9010;
													assign node9010 = (inp[7]) ? 4'b1001 : node9011;
														assign node9011 = (inp[8]) ? 4'b1001 : 4'b0100;
													assign node9015 = (inp[7]) ? node9019 : node9016;
														assign node9016 = (inp[8]) ? 4'b1001 : 4'b1000;
														assign node9019 = (inp[8]) ? 4'b1000 : 4'b1001;
										assign node9022 = (inp[11]) ? node9040 : node9023;
											assign node9023 = (inp[1]) ? node9031 : node9024;
												assign node9024 = (inp[13]) ? node9026 : 4'b0101;
													assign node9026 = (inp[8]) ? node9028 : 4'b0100;
														assign node9028 = (inp[2]) ? 4'b1000 : 4'b1001;
												assign node9031 = (inp[7]) ? node9033 : 4'b1001;
													assign node9033 = (inp[2]) ? node9037 : node9034;
														assign node9034 = (inp[8]) ? 4'b1001 : 4'b1000;
														assign node9037 = (inp[8]) ? 4'b1000 : 4'b1001;
											assign node9040 = (inp[13]) ? node9054 : node9041;
												assign node9041 = (inp[8]) ? node9049 : node9042;
													assign node9042 = (inp[2]) ? node9046 : node9043;
														assign node9043 = (inp[7]) ? 4'b1000 : 4'b1001;
														assign node9046 = (inp[7]) ? 4'b0001 : 4'b1000;
													assign node9049 = (inp[7]) ? node9051 : 4'b0001;
														assign node9051 = (inp[14]) ? 4'b0000 : 4'b0001;
												assign node9054 = (inp[8]) ? node9060 : node9055;
													assign node9055 = (inp[14]) ? 4'b0001 : node9056;
														assign node9056 = (inp[7]) ? 4'b0000 : 4'b0001;
													assign node9060 = (inp[2]) ? 4'b0000 : node9061;
														assign node9061 = (inp[1]) ? 4'b0000 : 4'b0000;
									assign node9065 = (inp[2]) ? node9107 : node9066;
										assign node9066 = (inp[7]) ? node9092 : node9067;
											assign node9067 = (inp[13]) ? node9081 : node9068;
												assign node9068 = (inp[11]) ? node9074 : node9069;
													assign node9069 = (inp[8]) ? 4'b1000 : node9070;
														assign node9070 = (inp[14]) ? 4'b0000 : 4'b0001;
													assign node9074 = (inp[14]) ? node9078 : node9075;
														assign node9075 = (inp[6]) ? 4'b1001 : 4'b0000;
														assign node9078 = (inp[8]) ? 4'b1001 : 4'b1000;
												assign node9081 = (inp[8]) ? node9087 : node9082;
													assign node9082 = (inp[14]) ? 4'b1000 : node9083;
														assign node9083 = (inp[11]) ? 4'b1001 : 4'b1001;
													assign node9087 = (inp[14]) ? 4'b1001 : node9088;
														assign node9088 = (inp[11]) ? 4'b0000 : 4'b1000;
											assign node9092 = (inp[14]) ? node9098 : node9093;
												assign node9093 = (inp[8]) ? node9095 : 4'b1000;
													assign node9095 = (inp[13]) ? 4'b0001 : 4'b1001;
												assign node9098 = (inp[8]) ? node9100 : 4'b0001;
													assign node9100 = (inp[1]) ? node9104 : node9101;
														assign node9101 = (inp[6]) ? 4'b1000 : 4'b0000;
														assign node9104 = (inp[11]) ? 4'b1000 : 4'b0000;
										assign node9107 = (inp[6]) ? node9133 : node9108;
											assign node9108 = (inp[11]) ? node9120 : node9109;
												assign node9109 = (inp[1]) ? node9113 : node9110;
													assign node9110 = (inp[13]) ? 4'b0000 : 4'b1000;
													assign node9113 = (inp[7]) ? node9117 : node9114;
														assign node9114 = (inp[8]) ? 4'b0001 : 4'b0000;
														assign node9117 = (inp[8]) ? 4'b0000 : 4'b0001;
												assign node9120 = (inp[1]) ? node9128 : node9121;
													assign node9121 = (inp[13]) ? node9125 : node9122;
														assign node9122 = (inp[8]) ? 4'b0000 : 4'b0000;
														assign node9125 = (inp[8]) ? 4'b1000 : 4'b0000;
													assign node9128 = (inp[14]) ? node9130 : 4'b1000;
														assign node9130 = (inp[7]) ? 4'b1000 : 4'b1001;
											assign node9133 = (inp[1]) ? node9149 : node9134;
												assign node9134 = (inp[11]) ? node9142 : node9135;
													assign node9135 = (inp[13]) ? node9139 : node9136;
														assign node9136 = (inp[7]) ? 4'b0001 : 4'b0000;
														assign node9139 = (inp[14]) ? 4'b1001 : 4'b1000;
													assign node9142 = (inp[13]) ? node9146 : node9143;
														assign node9143 = (inp[7]) ? 4'b1000 : 4'b1000;
														assign node9146 = (inp[7]) ? 4'b0001 : 4'b1000;
												assign node9149 = (inp[11]) ? node9155 : node9150;
													assign node9150 = (inp[14]) ? node9152 : 4'b1001;
														assign node9152 = (inp[7]) ? 4'b1001 : 4'b0000;
													assign node9155 = (inp[13]) ? node9157 : 4'b0001;
														assign node9157 = (inp[14]) ? 4'b0000 : 4'b0000;
						assign node9160 = (inp[9]) ? node9522 : node9161;
							assign node9161 = (inp[12]) ? node9345 : node9162;
								assign node9162 = (inp[10]) ? node9262 : node9163;
									assign node9163 = (inp[2]) ? node9217 : node9164;
										assign node9164 = (inp[6]) ? node9190 : node9165;
											assign node9165 = (inp[8]) ? node9177 : node9166;
												assign node9166 = (inp[13]) ? node9170 : node9167;
													assign node9167 = (inp[11]) ? 4'b0000 : 4'b0001;
													assign node9170 = (inp[11]) ? node9174 : node9171;
														assign node9171 = (inp[1]) ? 4'b0000 : 4'b1000;
														assign node9174 = (inp[1]) ? 4'b1000 : 4'b0000;
												assign node9177 = (inp[7]) ? node9185 : node9178;
													assign node9178 = (inp[14]) ? node9182 : node9179;
														assign node9179 = (inp[13]) ? 4'b0000 : 4'b1000;
														assign node9182 = (inp[1]) ? 4'b1001 : 4'b0001;
													assign node9185 = (inp[14]) ? 4'b0000 : node9186;
														assign node9186 = (inp[11]) ? 4'b1001 : 4'b0001;
											assign node9190 = (inp[14]) ? node9202 : node9191;
												assign node9191 = (inp[8]) ? node9199 : node9192;
													assign node9192 = (inp[7]) ? node9196 : node9193;
														assign node9193 = (inp[1]) ? 4'b1001 : 4'b0001;
														assign node9196 = (inp[13]) ? 4'b1000 : 4'b0000;
													assign node9199 = (inp[7]) ? 4'b0001 : 4'b0000;
												assign node9202 = (inp[11]) ? node9210 : node9203;
													assign node9203 = (inp[13]) ? node9207 : node9204;
														assign node9204 = (inp[8]) ? 4'b0001 : 4'b0000;
														assign node9207 = (inp[1]) ? 4'b1001 : 4'b0000;
													assign node9210 = (inp[13]) ? node9214 : node9211;
														assign node9211 = (inp[1]) ? 4'b1000 : 4'b1000;
														assign node9214 = (inp[8]) ? 4'b0000 : 4'b0001;
										assign node9217 = (inp[11]) ? node9239 : node9218;
											assign node9218 = (inp[6]) ? node9230 : node9219;
												assign node9219 = (inp[13]) ? node9225 : node9220;
													assign node9220 = (inp[8]) ? 4'b0000 : node9221;
														assign node9221 = (inp[7]) ? 4'b1001 : 4'b1000;
													assign node9225 = (inp[8]) ? node9227 : 4'b0001;
														assign node9227 = (inp[7]) ? 4'b0000 : 4'b0001;
												assign node9230 = (inp[7]) ? node9236 : node9231;
													assign node9231 = (inp[8]) ? 4'b1001 : node9232;
														assign node9232 = (inp[13]) ? 4'b1000 : 4'b0000;
													assign node9236 = (inp[8]) ? 4'b1000 : 4'b1001;
											assign node9239 = (inp[8]) ? node9251 : node9240;
												assign node9240 = (inp[7]) ? node9246 : node9241;
													assign node9241 = (inp[1]) ? node9243 : 4'b1000;
														assign node9243 = (inp[14]) ? 4'b0000 : 4'b1000;
													assign node9246 = (inp[6]) ? 4'b0001 : node9247;
														assign node9247 = (inp[1]) ? 4'b1001 : 4'b0001;
												assign node9251 = (inp[7]) ? node9257 : node9252;
													assign node9252 = (inp[1]) ? 4'b1001 : node9253;
														assign node9253 = (inp[6]) ? 4'b1001 : 4'b0001;
													assign node9257 = (inp[13]) ? 4'b1000 : node9258;
														assign node9258 = (inp[14]) ? 4'b0000 : 4'b1000;
									assign node9262 = (inp[6]) ? node9306 : node9263;
										assign node9263 = (inp[11]) ? node9285 : node9264;
											assign node9264 = (inp[1]) ? node9278 : node9265;
												assign node9265 = (inp[13]) ? node9273 : node9266;
													assign node9266 = (inp[7]) ? node9270 : node9267;
														assign node9267 = (inp[8]) ? 4'b1001 : 4'b1000;
														assign node9270 = (inp[8]) ? 4'b1000 : 4'b1000;
													assign node9273 = (inp[8]) ? 4'b0000 : node9274;
														assign node9274 = (inp[7]) ? 4'b0001 : 4'b1001;
												assign node9278 = (inp[13]) ? 4'b0000 : node9279;
													assign node9279 = (inp[8]) ? 4'b0001 : node9280;
														assign node9280 = (inp[14]) ? 4'b1000 : 4'b0001;
											assign node9285 = (inp[13]) ? node9297 : node9286;
												assign node9286 = (inp[1]) ? node9292 : node9287;
													assign node9287 = (inp[7]) ? node9289 : 4'b0001;
														assign node9289 = (inp[14]) ? 4'b0000 : 4'b0000;
													assign node9292 = (inp[8]) ? 4'b1111 : node9293;
														assign node9293 = (inp[14]) ? 4'b0000 : 4'b0001;
												assign node9297 = (inp[8]) ? node9303 : node9298;
													assign node9298 = (inp[7]) ? node9300 : 4'b0000;
														assign node9300 = (inp[2]) ? 4'b1111 : 4'b0000;
													assign node9303 = (inp[7]) ? 4'b1110 : 4'b1111;
										assign node9306 = (inp[11]) ? node9330 : node9307;
											assign node9307 = (inp[13]) ? node9321 : node9308;
												assign node9308 = (inp[1]) ? node9316 : node9309;
													assign node9309 = (inp[8]) ? node9313 : node9310;
														assign node9310 = (inp[7]) ? 4'b0000 : 4'b0000;
														assign node9313 = (inp[7]) ? 4'b0000 : 4'b0001;
													assign node9316 = (inp[8]) ? node9318 : 4'b0000;
														assign node9318 = (inp[2]) ? 4'b1110 : 4'b1111;
												assign node9321 = (inp[7]) ? node9325 : node9322;
													assign node9322 = (inp[2]) ? 4'b1111 : 4'b0000;
													assign node9325 = (inp[1]) ? node9327 : 4'b1111;
														assign node9327 = (inp[14]) ? 4'b1111 : 4'b1110;
											assign node9330 = (inp[13]) ? node9338 : node9331;
												assign node9331 = (inp[1]) ? 4'b0111 : node9332;
													assign node9332 = (inp[7]) ? 4'b1111 : node9333;
														assign node9333 = (inp[2]) ? 4'b1111 : 4'b1110;
												assign node9338 = (inp[8]) ? node9342 : node9339;
													assign node9339 = (inp[7]) ? 4'b0111 : 4'b0110;
													assign node9342 = (inp[7]) ? 4'b0110 : 4'b0111;
								assign node9345 = (inp[10]) ? node9443 : node9346;
									assign node9346 = (inp[11]) ? node9398 : node9347;
										assign node9347 = (inp[6]) ? node9375 : node9348;
											assign node9348 = (inp[13]) ? node9364 : node9349;
												assign node9349 = (inp[1]) ? node9357 : node9350;
													assign node9350 = (inp[7]) ? node9354 : node9351;
														assign node9351 = (inp[14]) ? 4'b1000 : 4'b1000;
														assign node9354 = (inp[14]) ? 4'b1000 : 4'b1001;
													assign node9357 = (inp[8]) ? node9361 : node9358;
														assign node9358 = (inp[14]) ? 4'b0000 : 4'b1000;
														assign node9361 = (inp[14]) ? 4'b0000 : 4'b0001;
												assign node9364 = (inp[1]) ? node9370 : node9365;
													assign node9365 = (inp[7]) ? node9367 : 4'b0001;
														assign node9367 = (inp[14]) ? 4'b0001 : 4'b0000;
													assign node9370 = (inp[14]) ? node9372 : 4'b0000;
														assign node9372 = (inp[8]) ? 4'b0000 : 4'b0001;
											assign node9375 = (inp[8]) ? node9387 : node9376;
												assign node9376 = (inp[1]) ? node9382 : node9377;
													assign node9377 = (inp[13]) ? 4'b0000 : node9378;
														assign node9378 = (inp[2]) ? 4'b0001 : 4'b0000;
													assign node9382 = (inp[13]) ? node9384 : 4'b0000;
														assign node9384 = (inp[7]) ? 4'b1111 : 4'b1110;
												assign node9387 = (inp[13]) ? node9391 : node9388;
													assign node9388 = (inp[1]) ? 4'b1111 : 4'b0001;
													assign node9391 = (inp[7]) ? node9395 : node9392;
														assign node9392 = (inp[2]) ? 4'b1111 : 4'b1110;
														assign node9395 = (inp[1]) ? 4'b1110 : 4'b1110;
										assign node9398 = (inp[6]) ? node9418 : node9399;
											assign node9399 = (inp[13]) ? node9409 : node9400;
												assign node9400 = (inp[8]) ? node9406 : node9401;
													assign node9401 = (inp[7]) ? 4'b0001 : node9402;
														assign node9402 = (inp[14]) ? 4'b0000 : 4'b0000;
													assign node9406 = (inp[7]) ? 4'b0000 : 4'b1111;
												assign node9409 = (inp[8]) ? node9415 : node9410;
													assign node9410 = (inp[14]) ? 4'b1111 : node9411;
														assign node9411 = (inp[2]) ? 4'b1110 : 4'b1111;
													assign node9415 = (inp[7]) ? 4'b1110 : 4'b1111;
											assign node9418 = (inp[1]) ? node9430 : node9419;
												assign node9419 = (inp[13]) ? node9427 : node9420;
													assign node9420 = (inp[2]) ? node9424 : node9421;
														assign node9421 = (inp[8]) ? 4'b1111 : 4'b1111;
														assign node9424 = (inp[8]) ? 4'b1110 : 4'b1110;
													assign node9427 = (inp[2]) ? 4'b0111 : 4'b1110;
												assign node9430 = (inp[13]) ? node9438 : node9431;
													assign node9431 = (inp[8]) ? node9435 : node9432;
														assign node9432 = (inp[7]) ? 4'b0111 : 4'b1110;
														assign node9435 = (inp[14]) ? 4'b0110 : 4'b0111;
													assign node9438 = (inp[7]) ? 4'b0110 : node9439;
														assign node9439 = (inp[2]) ? 4'b0110 : 4'b0110;
									assign node9443 = (inp[7]) ? node9483 : node9444;
										assign node9444 = (inp[8]) ? node9466 : node9445;
											assign node9445 = (inp[2]) ? node9455 : node9446;
												assign node9446 = (inp[14]) ? node9452 : node9447;
													assign node9447 = (inp[13]) ? 4'b1111 : node9448;
														assign node9448 = (inp[11]) ? 4'b0111 : 4'b0111;
													assign node9452 = (inp[6]) ? 4'b1110 : 4'b0110;
												assign node9455 = (inp[14]) ? node9461 : node9456;
													assign node9456 = (inp[1]) ? 4'b0110 : node9457;
														assign node9457 = (inp[6]) ? 4'b1110 : 4'b0110;
													assign node9461 = (inp[6]) ? node9463 : 4'b1110;
														assign node9463 = (inp[13]) ? 4'b1110 : 4'b0110;
											assign node9466 = (inp[2]) ? node9474 : node9467;
												assign node9467 = (inp[14]) ? node9471 : node9468;
													assign node9468 = (inp[6]) ? 4'b1110 : 4'b0110;
													assign node9471 = (inp[11]) ? 4'b0111 : 4'b1111;
												assign node9474 = (inp[6]) ? node9480 : node9475;
													assign node9475 = (inp[11]) ? 4'b1111 : node9476;
														assign node9476 = (inp[1]) ? 4'b0111 : 4'b1111;
													assign node9480 = (inp[13]) ? 4'b0111 : 4'b1111;
										assign node9483 = (inp[8]) ? node9503 : node9484;
											assign node9484 = (inp[14]) ? node9496 : node9485;
												assign node9485 = (inp[2]) ? node9491 : node9486;
													assign node9486 = (inp[13]) ? node9488 : 4'b0110;
														assign node9488 = (inp[11]) ? 4'b1110 : 4'b0110;
													assign node9491 = (inp[1]) ? node9493 : 4'b0111;
														assign node9493 = (inp[6]) ? 4'b0111 : 4'b1111;
												assign node9496 = (inp[13]) ? node9498 : 4'b0111;
													assign node9498 = (inp[1]) ? node9500 : 4'b1111;
														assign node9500 = (inp[2]) ? 4'b0111 : 4'b0111;
											assign node9503 = (inp[2]) ? node9513 : node9504;
												assign node9504 = (inp[14]) ? node9510 : node9505;
													assign node9505 = (inp[11]) ? 4'b1111 : node9506;
														assign node9506 = (inp[13]) ? 4'b0111 : 4'b0111;
													assign node9510 = (inp[6]) ? 4'b1110 : 4'b0110;
												assign node9513 = (inp[14]) ? 4'b0110 : node9514;
													assign node9514 = (inp[1]) ? node9518 : node9515;
														assign node9515 = (inp[13]) ? 4'b0110 : 4'b0110;
														assign node9518 = (inp[11]) ? 4'b1110 : 4'b0110;
							assign node9522 = (inp[12]) ? node9688 : node9523;
								assign node9523 = (inp[10]) ? node9603 : node9524;
									assign node9524 = (inp[11]) ? node9568 : node9525;
										assign node9525 = (inp[8]) ? node9547 : node9526;
											assign node9526 = (inp[7]) ? node9536 : node9527;
												assign node9527 = (inp[6]) ? node9533 : node9528;
													assign node9528 = (inp[2]) ? node9530 : 4'b1111;
														assign node9530 = (inp[1]) ? 4'b0110 : 4'b1110;
													assign node9533 = (inp[13]) ? 4'b0111 : 4'b0110;
												assign node9536 = (inp[14]) ? node9542 : node9537;
													assign node9537 = (inp[2]) ? 4'b0111 : node9538;
														assign node9538 = (inp[6]) ? 4'b0110 : 4'b1110;
													assign node9542 = (inp[6]) ? 4'b1111 : node9543;
														assign node9543 = (inp[2]) ? 4'b0111 : 4'b0111;
											assign node9547 = (inp[7]) ? node9557 : node9548;
												assign node9548 = (inp[2]) ? node9552 : node9549;
													assign node9549 = (inp[14]) ? 4'b0111 : 4'b0110;
													assign node9552 = (inp[13]) ? 4'b1111 : node9553;
														assign node9553 = (inp[1]) ? 4'b0111 : 4'b0111;
												assign node9557 = (inp[6]) ? node9563 : node9558;
													assign node9558 = (inp[13]) ? 4'b0110 : node9559;
														assign node9559 = (inp[1]) ? 4'b0110 : 4'b1110;
													assign node9563 = (inp[14]) ? 4'b1110 : node9564;
														assign node9564 = (inp[2]) ? 4'b1110 : 4'b0111;
										assign node9568 = (inp[14]) ? node9588 : node9569;
											assign node9569 = (inp[8]) ? node9577 : node9570;
												assign node9570 = (inp[2]) ? 4'b1110 : node9571;
													assign node9571 = (inp[7]) ? node9573 : 4'b0111;
														assign node9573 = (inp[1]) ? 4'b1110 : 4'b0110;
												assign node9577 = (inp[2]) ? node9583 : node9578;
													assign node9578 = (inp[7]) ? 4'b0111 : node9579;
														assign node9579 = (inp[6]) ? 4'b1110 : 4'b0110;
													assign node9583 = (inp[7]) ? 4'b0110 : node9584;
														assign node9584 = (inp[13]) ? 4'b0111 : 4'b0111;
											assign node9588 = (inp[6]) ? node9596 : node9589;
												assign node9589 = (inp[2]) ? 4'b1110 : node9590;
													assign node9590 = (inp[13]) ? node9592 : 4'b0110;
														assign node9592 = (inp[8]) ? 4'b1110 : 4'b1111;
												assign node9596 = (inp[8]) ? node9598 : 4'b1110;
													assign node9598 = (inp[7]) ? node9600 : 4'b0111;
														assign node9600 = (inp[1]) ? 4'b0110 : 4'b0110;
									assign node9603 = (inp[11]) ? node9655 : node9604;
										assign node9604 = (inp[6]) ? node9628 : node9605;
											assign node9605 = (inp[1]) ? node9617 : node9606;
												assign node9606 = (inp[2]) ? node9612 : node9607;
													assign node9607 = (inp[7]) ? node9609 : 4'b1110;
														assign node9609 = (inp[13]) ? 4'b0110 : 4'b1110;
													assign node9612 = (inp[13]) ? node9614 : 4'b1111;
														assign node9614 = (inp[14]) ? 4'b0111 : 4'b0111;
												assign node9617 = (inp[8]) ? node9623 : node9618;
													assign node9618 = (inp[13]) ? node9620 : 4'b1110;
														assign node9620 = (inp[7]) ? 4'b0111 : 4'b0110;
													assign node9623 = (inp[7]) ? node9625 : 4'b0111;
														assign node9625 = (inp[14]) ? 4'b0110 : 4'b0111;
											assign node9628 = (inp[1]) ? node9640 : node9629;
												assign node9629 = (inp[13]) ? node9635 : node9630;
													assign node9630 = (inp[8]) ? 4'b0110 : node9631;
														assign node9631 = (inp[7]) ? 4'b0111 : 4'b0110;
													assign node9635 = (inp[14]) ? 4'b1011 : node9636;
														assign node9636 = (inp[8]) ? 4'b1011 : 4'b0110;
												assign node9640 = (inp[13]) ? node9648 : node9641;
													assign node9641 = (inp[8]) ? node9645 : node9642;
														assign node9642 = (inp[7]) ? 4'b1011 : 4'b0110;
														assign node9645 = (inp[7]) ? 4'b1010 : 4'b1011;
													assign node9648 = (inp[14]) ? node9652 : node9649;
														assign node9649 = (inp[7]) ? 4'b1010 : 4'b1011;
														assign node9652 = (inp[7]) ? 4'b1010 : 4'b1010;
										assign node9655 = (inp[6]) ? node9673 : node9656;
											assign node9656 = (inp[1]) ? node9664 : node9657;
												assign node9657 = (inp[13]) ? node9661 : node9658;
													assign node9658 = (inp[8]) ? 4'b0110 : 4'b0111;
													assign node9661 = (inp[14]) ? 4'b1011 : 4'b0110;
												assign node9664 = (inp[7]) ? node9668 : node9665;
													assign node9665 = (inp[14]) ? 4'b0110 : 4'b1011;
													assign node9668 = (inp[8]) ? 4'b1010 : node9669;
														assign node9669 = (inp[14]) ? 4'b1011 : 4'b1010;
											assign node9673 = (inp[1]) ? node9681 : node9674;
												assign node9674 = (inp[8]) ? node9676 : 4'b1010;
													assign node9676 = (inp[7]) ? 4'b1010 : node9677;
														assign node9677 = (inp[13]) ? 4'b0011 : 4'b1011;
												assign node9681 = (inp[8]) ? node9685 : node9682;
													assign node9682 = (inp[7]) ? 4'b0011 : 4'b1010;
													assign node9685 = (inp[7]) ? 4'b0010 : 4'b0011;
								assign node9688 = (inp[10]) ? node9780 : node9689;
									assign node9689 = (inp[11]) ? node9735 : node9690;
										assign node9690 = (inp[6]) ? node9710 : node9691;
											assign node9691 = (inp[1]) ? node9701 : node9692;
												assign node9692 = (inp[8]) ? node9696 : node9693;
													assign node9693 = (inp[2]) ? 4'b1110 : 4'b1111;
													assign node9696 = (inp[13]) ? node9698 : 4'b1111;
														assign node9698 = (inp[7]) ? 4'b0110 : 4'b0111;
												assign node9701 = (inp[14]) ? node9705 : node9702;
													assign node9702 = (inp[8]) ? 4'b0110 : 4'b1110;
													assign node9705 = (inp[2]) ? node9707 : 4'b0111;
														assign node9707 = (inp[13]) ? 4'b0110 : 4'b0111;
											assign node9710 = (inp[13]) ? node9724 : node9711;
												assign node9711 = (inp[14]) ? node9719 : node9712;
													assign node9712 = (inp[2]) ? node9716 : node9713;
														assign node9713 = (inp[1]) ? 4'b0111 : 4'b0110;
														assign node9716 = (inp[1]) ? 4'b1011 : 4'b0111;
													assign node9719 = (inp[1]) ? 4'b0110 : node9720;
														assign node9720 = (inp[2]) ? 4'b0110 : 4'b0110;
												assign node9724 = (inp[2]) ? node9730 : node9725;
													assign node9725 = (inp[7]) ? node9727 : 4'b1011;
														assign node9727 = (inp[1]) ? 4'b1010 : 4'b1011;
													assign node9730 = (inp[7]) ? node9732 : 4'b0110;
														assign node9732 = (inp[8]) ? 4'b1010 : 4'b1011;
										assign node9735 = (inp[6]) ? node9761 : node9736;
											assign node9736 = (inp[1]) ? node9748 : node9737;
												assign node9737 = (inp[13]) ? node9743 : node9738;
													assign node9738 = (inp[8]) ? 4'b0110 : node9739;
														assign node9739 = (inp[7]) ? 4'b0110 : 4'b0111;
													assign node9743 = (inp[8]) ? 4'b1011 : node9744;
														assign node9744 = (inp[7]) ? 4'b1011 : 4'b0110;
												assign node9748 = (inp[13]) ? node9756 : node9749;
													assign node9749 = (inp[7]) ? node9753 : node9750;
														assign node9750 = (inp[8]) ? 4'b1011 : 4'b0110;
														assign node9753 = (inp[8]) ? 4'b1010 : 4'b1011;
													assign node9756 = (inp[7]) ? 4'b1010 : node9757;
														assign node9757 = (inp[8]) ? 4'b1011 : 4'b1010;
											assign node9761 = (inp[1]) ? node9775 : node9762;
												assign node9762 = (inp[13]) ? node9770 : node9763;
													assign node9763 = (inp[8]) ? node9767 : node9764;
														assign node9764 = (inp[7]) ? 4'b1011 : 4'b1010;
														assign node9767 = (inp[7]) ? 4'b1010 : 4'b1011;
													assign node9770 = (inp[14]) ? node9772 : 4'b1010;
														assign node9772 = (inp[2]) ? 4'b0010 : 4'b0011;
												assign node9775 = (inp[8]) ? node9777 : 4'b1010;
													assign node9777 = (inp[7]) ? 4'b0010 : 4'b0011;
									assign node9780 = (inp[13]) ? node9824 : node9781;
										assign node9781 = (inp[1]) ? node9799 : node9782;
											assign node9782 = (inp[11]) ? node9790 : node9783;
												assign node9783 = (inp[6]) ? 4'b0010 : node9784;
													assign node9784 = (inp[2]) ? 4'b1010 : node9785;
														assign node9785 = (inp[14]) ? 4'b1010 : 4'b1011;
												assign node9790 = (inp[7]) ? node9792 : 4'b1011;
													assign node9792 = (inp[8]) ? node9796 : node9793;
														assign node9793 = (inp[2]) ? 4'b1011 : 4'b1010;
														assign node9796 = (inp[2]) ? 4'b1010 : 4'b1010;
											assign node9799 = (inp[2]) ? node9813 : node9800;
												assign node9800 = (inp[14]) ? node9806 : node9801;
													assign node9801 = (inp[6]) ? node9803 : 4'b1010;
														assign node9803 = (inp[7]) ? 4'b1010 : 4'b1011;
													assign node9806 = (inp[11]) ? node9810 : node9807;
														assign node9807 = (inp[6]) ? 4'b1011 : 4'b0010;
														assign node9810 = (inp[6]) ? 4'b0011 : 4'b1011;
												assign node9813 = (inp[6]) ? node9817 : node9814;
													assign node9814 = (inp[11]) ? 4'b0010 : 4'b0011;
													assign node9817 = (inp[11]) ? node9821 : node9818;
														assign node9818 = (inp[14]) ? 4'b1010 : 4'b1011;
														assign node9821 = (inp[7]) ? 4'b0011 : 4'b1010;
										assign node9824 = (inp[8]) ? node9850 : node9825;
											assign node9825 = (inp[7]) ? node9837 : node9826;
												assign node9826 = (inp[2]) ? node9832 : node9827;
													assign node9827 = (inp[14]) ? node9829 : 4'b0011;
														assign node9829 = (inp[1]) ? 4'b1010 : 4'b0010;
													assign node9832 = (inp[11]) ? node9834 : 4'b1010;
														assign node9834 = (inp[1]) ? 4'b1010 : 4'b0010;
												assign node9837 = (inp[14]) ? node9843 : node9838;
													assign node9838 = (inp[2]) ? 4'b0011 : node9839;
														assign node9839 = (inp[6]) ? 4'b1010 : 4'b0010;
													assign node9843 = (inp[11]) ? node9847 : node9844;
														assign node9844 = (inp[1]) ? 4'b1011 : 4'b0011;
														assign node9847 = (inp[2]) ? 4'b1011 : 4'b0011;
											assign node9850 = (inp[7]) ? node9866 : node9851;
												assign node9851 = (inp[14]) ? node9859 : node9852;
													assign node9852 = (inp[2]) ? node9856 : node9853;
														assign node9853 = (inp[11]) ? 4'b0010 : 4'b0010;
														assign node9856 = (inp[6]) ? 4'b1011 : 4'b0011;
													assign node9859 = (inp[6]) ? node9863 : node9860;
														assign node9860 = (inp[11]) ? 4'b1011 : 4'b0011;
														assign node9863 = (inp[11]) ? 4'b0011 : 4'b1011;
												assign node9866 = (inp[2]) ? node9872 : node9867;
													assign node9867 = (inp[14]) ? 4'b1010 : node9868;
														assign node9868 = (inp[11]) ? 4'b0011 : 4'b1011;
													assign node9872 = (inp[6]) ? 4'b0010 : 4'b1010;
					assign node9875 = (inp[9]) ? node10603 : node9876;
						assign node9876 = (inp[10]) ? node10252 : node9877;
							assign node9877 = (inp[5]) ? node10067 : node9878;
								assign node9878 = (inp[12]) ? node9974 : node9879;
									assign node9879 = (inp[14]) ? node9933 : node9880;
										assign node9880 = (inp[1]) ? node9906 : node9881;
											assign node9881 = (inp[2]) ? node9893 : node9882;
												assign node9882 = (inp[11]) ? node9888 : node9883;
													assign node9883 = (inp[6]) ? node9885 : 4'b1001;
														assign node9885 = (inp[13]) ? 4'b0000 : 4'b0001;
													assign node9888 = (inp[7]) ? 4'b1000 : node9889;
														assign node9889 = (inp[8]) ? 4'b0000 : 4'b0001;
												assign node9893 = (inp[11]) ? node9901 : node9894;
													assign node9894 = (inp[13]) ? node9898 : node9895;
														assign node9895 = (inp[6]) ? 4'b0000 : 4'b1000;
														assign node9898 = (inp[6]) ? 4'b1001 : 4'b0001;
													assign node9901 = (inp[8]) ? 4'b0001 : node9902;
														assign node9902 = (inp[6]) ? 4'b1001 : 4'b0001;
											assign node9906 = (inp[7]) ? node9918 : node9907;
												assign node9907 = (inp[8]) ? node9913 : node9908;
													assign node9908 = (inp[2]) ? node9910 : 4'b0001;
														assign node9910 = (inp[11]) ? 4'b1000 : 4'b0000;
													assign node9913 = (inp[2]) ? node9915 : 4'b0000;
														assign node9915 = (inp[6]) ? 4'b0001 : 4'b0001;
												assign node9918 = (inp[6]) ? node9926 : node9919;
													assign node9919 = (inp[11]) ? node9923 : node9920;
														assign node9920 = (inp[8]) ? 4'b0000 : 4'b0000;
														assign node9923 = (inp[13]) ? 4'b1001 : 4'b0000;
													assign node9926 = (inp[11]) ? node9930 : node9927;
														assign node9927 = (inp[8]) ? 4'b1000 : 4'b1000;
														assign node9930 = (inp[13]) ? 4'b0000 : 4'b0001;
										assign node9933 = (inp[1]) ? node9955 : node9934;
											assign node9934 = (inp[7]) ? node9946 : node9935;
												assign node9935 = (inp[8]) ? node9941 : node9936;
													assign node9936 = (inp[13]) ? 4'b0000 : node9937;
														assign node9937 = (inp[6]) ? 4'b1000 : 4'b0000;
													assign node9941 = (inp[2]) ? 4'b1001 : node9942;
														assign node9942 = (inp[13]) ? 4'b1001 : 4'b0001;
												assign node9946 = (inp[8]) ? node9950 : node9947;
													assign node9947 = (inp[6]) ? 4'b0001 : 4'b1001;
													assign node9950 = (inp[2]) ? node9952 : 4'b0000;
														assign node9952 = (inp[13]) ? 4'b1000 : 4'b0000;
											assign node9955 = (inp[8]) ? node9965 : node9956;
												assign node9956 = (inp[7]) ? node9960 : node9957;
													assign node9957 = (inp[2]) ? 4'b1000 : 4'b0000;
													assign node9960 = (inp[2]) ? node9962 : 4'b0001;
														assign node9962 = (inp[13]) ? 4'b0001 : 4'b1001;
												assign node9965 = (inp[2]) ? node9969 : node9966;
													assign node9966 = (inp[7]) ? 4'b1000 : 4'b1001;
													assign node9969 = (inp[13]) ? node9971 : 4'b0001;
														assign node9971 = (inp[6]) ? 4'b0001 : 4'b1001;
									assign node9974 = (inp[6]) ? node10018 : node9975;
										assign node9975 = (inp[11]) ? node9997 : node9976;
											assign node9976 = (inp[1]) ? node9986 : node9977;
												assign node9977 = (inp[13]) ? node9981 : node9978;
													assign node9978 = (inp[14]) ? 4'b1001 : 4'b1000;
													assign node9981 = (inp[7]) ? node9983 : 4'b1000;
														assign node9983 = (inp[8]) ? 4'b0000 : 4'b0001;
												assign node9986 = (inp[2]) ? node9992 : node9987;
													assign node9987 = (inp[7]) ? node9989 : 4'b0001;
														assign node9989 = (inp[13]) ? 4'b0000 : 4'b0001;
													assign node9992 = (inp[7]) ? 4'b0000 : node9993;
														assign node9993 = (inp[8]) ? 4'b0001 : 4'b0000;
											assign node9997 = (inp[1]) ? node10007 : node9998;
												assign node9998 = (inp[13]) ? node10004 : node9999;
													assign node9999 = (inp[7]) ? 4'b0000 : node10000;
														assign node10000 = (inp[2]) ? 4'b0000 : 4'b0000;
													assign node10004 = (inp[7]) ? 4'b1110 : 4'b0000;
												assign node10007 = (inp[8]) ? node10011 : node10008;
													assign node10008 = (inp[2]) ? 4'b0000 : 4'b1110;
													assign node10011 = (inp[7]) ? node10015 : node10012;
														assign node10012 = (inp[14]) ? 4'b1111 : 4'b1110;
														assign node10015 = (inp[2]) ? 4'b1110 : 4'b1111;
										assign node10018 = (inp[11]) ? node10046 : node10019;
											assign node10019 = (inp[1]) ? node10033 : node10020;
												assign node10020 = (inp[13]) ? node10028 : node10021;
													assign node10021 = (inp[7]) ? node10025 : node10022;
														assign node10022 = (inp[8]) ? 4'b0000 : 4'b0000;
														assign node10025 = (inp[8]) ? 4'b0000 : 4'b0001;
													assign node10028 = (inp[8]) ? node10030 : 4'b0000;
														assign node10030 = (inp[7]) ? 4'b1110 : 4'b1111;
												assign node10033 = (inp[7]) ? node10041 : node10034;
													assign node10034 = (inp[8]) ? node10038 : node10035;
														assign node10035 = (inp[13]) ? 4'b1110 : 4'b0000;
														assign node10038 = (inp[13]) ? 4'b1110 : 4'b1111;
													assign node10041 = (inp[8]) ? node10043 : 4'b1111;
														assign node10043 = (inp[14]) ? 4'b1110 : 4'b1111;
											assign node10046 = (inp[8]) ? node10058 : node10047;
												assign node10047 = (inp[13]) ? node10053 : node10048;
													assign node10048 = (inp[2]) ? 4'b1110 : node10049;
														assign node10049 = (inp[14]) ? 4'b0111 : 4'b1110;
													assign node10053 = (inp[7]) ? 4'b0111 : node10054;
														assign node10054 = (inp[1]) ? 4'b0110 : 4'b1110;
												assign node10058 = (inp[1]) ? node10062 : node10059;
													assign node10059 = (inp[13]) ? 4'b0110 : 4'b1110;
													assign node10062 = (inp[2]) ? node10064 : 4'b0110;
														assign node10064 = (inp[7]) ? 4'b0110 : 4'b0111;
								assign node10067 = (inp[12]) ? node10157 : node10068;
									assign node10068 = (inp[11]) ? node10108 : node10069;
										assign node10069 = (inp[7]) ? node10085 : node10070;
											assign node10070 = (inp[8]) ? node10078 : node10071;
												assign node10071 = (inp[2]) ? 4'b0010 : node10072;
													assign node10072 = (inp[14]) ? 4'b1010 : node10073;
														assign node10073 = (inp[6]) ? 4'b1011 : 4'b1011;
												assign node10078 = (inp[14]) ? node10080 : 4'b0011;
													assign node10080 = (inp[2]) ? 4'b1011 : node10081;
														assign node10081 = (inp[6]) ? 4'b0011 : 4'b0011;
											assign node10085 = (inp[6]) ? node10099 : node10086;
												assign node10086 = (inp[1]) ? node10092 : node10087;
													assign node10087 = (inp[13]) ? node10089 : 4'b1010;
														assign node10089 = (inp[8]) ? 4'b0011 : 4'b0010;
													assign node10092 = (inp[8]) ? node10096 : node10093;
														assign node10093 = (inp[13]) ? 4'b0010 : 4'b0011;
														assign node10096 = (inp[2]) ? 4'b0010 : 4'b0010;
												assign node10099 = (inp[13]) ? node10105 : node10100;
													assign node10100 = (inp[1]) ? 4'b1010 : node10101;
														assign node10101 = (inp[2]) ? 4'b0010 : 4'b0010;
													assign node10105 = (inp[14]) ? 4'b1010 : 4'b1011;
										assign node10108 = (inp[1]) ? node10134 : node10109;
											assign node10109 = (inp[8]) ? node10123 : node10110;
												assign node10110 = (inp[7]) ? node10116 : node10111;
													assign node10111 = (inp[14]) ? 4'b1010 : node10112;
														assign node10112 = (inp[2]) ? 4'b1010 : 4'b1011;
													assign node10116 = (inp[13]) ? node10120 : node10117;
														assign node10117 = (inp[6]) ? 4'b1011 : 4'b0011;
														assign node10120 = (inp[2]) ? 4'b0011 : 4'b1010;
												assign node10123 = (inp[7]) ? node10127 : node10124;
													assign node10124 = (inp[13]) ? 4'b1011 : 4'b0011;
													assign node10127 = (inp[14]) ? node10131 : node10128;
														assign node10128 = (inp[2]) ? 4'b0010 : 4'b0011;
														assign node10131 = (inp[13]) ? 4'b0010 : 4'b1010;
											assign node10134 = (inp[6]) ? node10146 : node10135;
												assign node10135 = (inp[7]) ? node10143 : node10136;
													assign node10136 = (inp[2]) ? node10140 : node10137;
														assign node10137 = (inp[13]) ? 4'b1010 : 4'b0010;
														assign node10140 = (inp[8]) ? 4'b1011 : 4'b1010;
													assign node10143 = (inp[14]) ? 4'b1010 : 4'b1011;
												assign node10146 = (inp[7]) ? node10154 : node10147;
													assign node10147 = (inp[8]) ? node10151 : node10148;
														assign node10148 = (inp[13]) ? 4'b0010 : 4'b1010;
														assign node10151 = (inp[2]) ? 4'b0011 : 4'b0010;
													assign node10154 = (inp[8]) ? 4'b0010 : 4'b0011;
									assign node10157 = (inp[6]) ? node10203 : node10158;
										assign node10158 = (inp[13]) ? node10182 : node10159;
											assign node10159 = (inp[7]) ? node10171 : node10160;
												assign node10160 = (inp[8]) ? node10166 : node10161;
													assign node10161 = (inp[11]) ? node10163 : 4'b1010;
														assign node10163 = (inp[2]) ? 4'b0010 : 4'b0010;
													assign node10166 = (inp[14]) ? 4'b0011 : node10167;
														assign node10167 = (inp[1]) ? 4'b0010 : 4'b0011;
												assign node10171 = (inp[1]) ? node10175 : node10172;
													assign node10172 = (inp[14]) ? 4'b0011 : 4'b0010;
													assign node10175 = (inp[11]) ? node10179 : node10176;
														assign node10176 = (inp[14]) ? 4'b0010 : 4'b1010;
														assign node10179 = (inp[14]) ? 4'b1110 : 4'b1111;
											assign node10182 = (inp[11]) ? node10192 : node10183;
												assign node10183 = (inp[8]) ? 4'b0011 : node10184;
													assign node10184 = (inp[1]) ? node10188 : node10185;
														assign node10185 = (inp[2]) ? 4'b1010 : 4'b1011;
														assign node10188 = (inp[7]) ? 4'b0010 : 4'b0011;
												assign node10192 = (inp[1]) ? node10198 : node10193;
													assign node10193 = (inp[7]) ? 4'b1111 : node10194;
														assign node10194 = (inp[8]) ? 4'b1111 : 4'b0010;
													assign node10198 = (inp[8]) ? 4'b1111 : node10199;
														assign node10199 = (inp[7]) ? 4'b1111 : 4'b1110;
										assign node10203 = (inp[11]) ? node10231 : node10204;
											assign node10204 = (inp[13]) ? node10220 : node10205;
												assign node10205 = (inp[1]) ? node10213 : node10206;
													assign node10206 = (inp[7]) ? node10210 : node10207;
														assign node10207 = (inp[14]) ? 4'b0010 : 4'b0011;
														assign node10210 = (inp[2]) ? 4'b0010 : 4'b0010;
													assign node10213 = (inp[7]) ? node10217 : node10214;
														assign node10214 = (inp[8]) ? 4'b1111 : 4'b0010;
														assign node10217 = (inp[14]) ? 4'b1110 : 4'b0010;
												assign node10220 = (inp[8]) ? node10226 : node10221;
													assign node10221 = (inp[7]) ? 4'b1111 : node10222;
														assign node10222 = (inp[1]) ? 4'b1111 : 4'b0010;
													assign node10226 = (inp[7]) ? 4'b1110 : node10227;
														assign node10227 = (inp[2]) ? 4'b1111 : 4'b1110;
											assign node10231 = (inp[13]) ? node10245 : node10232;
												assign node10232 = (inp[2]) ? node10238 : node10233;
													assign node10233 = (inp[14]) ? node10235 : 4'b1111;
														assign node10235 = (inp[7]) ? 4'b1110 : 4'b1110;
													assign node10238 = (inp[14]) ? node10242 : node10239;
														assign node10239 = (inp[8]) ? 4'b0110 : 4'b0111;
														assign node10242 = (inp[8]) ? 4'b0110 : 4'b1110;
												assign node10245 = (inp[7]) ? 4'b0110 : node10246;
													assign node10246 = (inp[1]) ? node10248 : 4'b1110;
														assign node10248 = (inp[14]) ? 4'b0110 : 4'b0111;
							assign node10252 = (inp[12]) ? node10444 : node10253;
								assign node10253 = (inp[11]) ? node10355 : node10254;
									assign node10254 = (inp[5]) ? node10304 : node10255;
										assign node10255 = (inp[6]) ? node10281 : node10256;
											assign node10256 = (inp[13]) ? node10270 : node10257;
												assign node10257 = (inp[1]) ? node10263 : node10258;
													assign node10258 = (inp[8]) ? 4'b1001 : node10259;
														assign node10259 = (inp[2]) ? 4'b1000 : 4'b1001;
													assign node10263 = (inp[2]) ? node10267 : node10264;
														assign node10264 = (inp[14]) ? 4'b0001 : 4'b0001;
														assign node10267 = (inp[14]) ? 4'b0000 : 4'b1000;
												assign node10270 = (inp[14]) ? node10276 : node10271;
													assign node10271 = (inp[8]) ? node10273 : 4'b0001;
														assign node10273 = (inp[2]) ? 4'b0000 : 4'b0001;
													assign node10276 = (inp[8]) ? 4'b0000 : node10277;
														assign node10277 = (inp[2]) ? 4'b1000 : 4'b0000;
											assign node10281 = (inp[13]) ? node10297 : node10282;
												assign node10282 = (inp[1]) ? node10290 : node10283;
													assign node10283 = (inp[7]) ? node10287 : node10284;
														assign node10284 = (inp[8]) ? 4'b0001 : 4'b0000;
														assign node10287 = (inp[8]) ? 4'b0000 : 4'b0001;
													assign node10290 = (inp[14]) ? node10294 : node10291;
														assign node10291 = (inp[2]) ? 4'b0000 : 4'b0000;
														assign node10294 = (inp[2]) ? 4'b1111 : 4'b1110;
												assign node10297 = (inp[14]) ? node10299 : 4'b1111;
													assign node10299 = (inp[1]) ? 4'b1110 : node10300;
														assign node10300 = (inp[7]) ? 4'b1110 : 4'b1111;
										assign node10304 = (inp[6]) ? node10328 : node10305;
											assign node10305 = (inp[1]) ? node10319 : node10306;
												assign node10306 = (inp[13]) ? node10312 : node10307;
													assign node10307 = (inp[2]) ? 4'b1010 : node10308;
														assign node10308 = (inp[7]) ? 4'b1010 : 4'b1010;
													assign node10312 = (inp[7]) ? node10316 : node10313;
														assign node10313 = (inp[8]) ? 4'b0010 : 4'b1010;
														assign node10316 = (inp[2]) ? 4'b0011 : 4'b0010;
												assign node10319 = (inp[8]) ? node10323 : node10320;
													assign node10320 = (inp[14]) ? 4'b1010 : 4'b0010;
													assign node10323 = (inp[14]) ? 4'b0011 : node10324;
														assign node10324 = (inp[13]) ? 4'b0010 : 4'b0010;
											assign node10328 = (inp[13]) ? node10342 : node10329;
												assign node10329 = (inp[7]) ? node10335 : node10330;
													assign node10330 = (inp[14]) ? node10332 : 4'b0011;
														assign node10332 = (inp[8]) ? 4'b0011 : 4'b0010;
													assign node10335 = (inp[14]) ? node10339 : node10336;
														assign node10336 = (inp[8]) ? 4'b1110 : 4'b0010;
														assign node10339 = (inp[1]) ? 4'b1111 : 4'b0011;
												assign node10342 = (inp[8]) ? node10350 : node10343;
													assign node10343 = (inp[1]) ? node10347 : node10344;
														assign node10344 = (inp[2]) ? 4'b0010 : 4'b0011;
														assign node10347 = (inp[7]) ? 4'b1111 : 4'b1110;
													assign node10350 = (inp[7]) ? node10352 : 4'b1111;
														assign node10352 = (inp[2]) ? 4'b1110 : 4'b1111;
									assign node10355 = (inp[6]) ? node10401 : node10356;
										assign node10356 = (inp[13]) ? node10376 : node10357;
											assign node10357 = (inp[1]) ? node10365 : node10358;
												assign node10358 = (inp[5]) ? node10360 : 4'b0000;
													assign node10360 = (inp[14]) ? node10362 : 4'b0011;
														assign node10362 = (inp[7]) ? 4'b0010 : 4'b0010;
												assign node10365 = (inp[5]) ? node10373 : node10366;
													assign node10366 = (inp[7]) ? node10370 : node10367;
														assign node10367 = (inp[8]) ? 4'b0000 : 4'b0001;
														assign node10370 = (inp[14]) ? 4'b1111 : 4'b0000;
													assign node10373 = (inp[2]) ? 4'b1110 : 4'b1111;
											assign node10376 = (inp[1]) ? node10388 : node10377;
												assign node10377 = (inp[7]) ? node10385 : node10378;
													assign node10378 = (inp[14]) ? node10382 : node10379;
														assign node10379 = (inp[5]) ? 4'b0010 : 4'b0000;
														assign node10382 = (inp[8]) ? 4'b1111 : 4'b0000;
													assign node10385 = (inp[8]) ? 4'b1110 : 4'b1111;
												assign node10388 = (inp[5]) ? node10394 : node10389;
													assign node10389 = (inp[7]) ? node10391 : 4'b1111;
														assign node10391 = (inp[8]) ? 4'b1110 : 4'b1111;
													assign node10394 = (inp[2]) ? node10398 : node10395;
														assign node10395 = (inp[8]) ? 4'b1111 : 4'b1110;
														assign node10398 = (inp[14]) ? 4'b1110 : 4'b1110;
										assign node10401 = (inp[13]) ? node10419 : node10402;
											assign node10402 = (inp[1]) ? node10408 : node10403;
												assign node10403 = (inp[7]) ? node10405 : 4'b1110;
													assign node10405 = (inp[8]) ? 4'b1110 : 4'b1111;
												assign node10408 = (inp[7]) ? node10414 : node10409;
													assign node10409 = (inp[8]) ? node10411 : 4'b1110;
														assign node10411 = (inp[14]) ? 4'b0111 : 4'b1110;
													assign node10414 = (inp[8]) ? node10416 : 4'b0111;
														assign node10416 = (inp[2]) ? 4'b0110 : 4'b0111;
											assign node10419 = (inp[14]) ? node10433 : node10420;
												assign node10420 = (inp[1]) ? node10426 : node10421;
													assign node10421 = (inp[8]) ? node10423 : 4'b1110;
														assign node10423 = (inp[5]) ? 4'b0110 : 4'b0111;
													assign node10426 = (inp[7]) ? node10430 : node10427;
														assign node10427 = (inp[2]) ? 4'b0110 : 4'b0111;
														assign node10430 = (inp[8]) ? 4'b0110 : 4'b0110;
												assign node10433 = (inp[5]) ? node10439 : node10434;
													assign node10434 = (inp[7]) ? node10436 : 4'b0111;
														assign node10436 = (inp[1]) ? 4'b0110 : 4'b0111;
													assign node10439 = (inp[2]) ? 4'b0110 : node10440;
														assign node10440 = (inp[1]) ? 4'b0110 : 4'b0111;
								assign node10444 = (inp[14]) ? node10528 : node10445;
									assign node10445 = (inp[8]) ? node10481 : node10446;
										assign node10446 = (inp[2]) ? node10462 : node10447;
											assign node10447 = (inp[7]) ? node10455 : node10448;
												assign node10448 = (inp[6]) ? node10450 : 4'b0111;
													assign node10450 = (inp[13]) ? 4'b0111 : node10451;
														assign node10451 = (inp[5]) ? 4'b0111 : 4'b1111;
												assign node10455 = (inp[5]) ? 4'b0110 : node10456;
													assign node10456 = (inp[6]) ? 4'b0110 : node10457;
														assign node10457 = (inp[13]) ? 4'b1110 : 4'b0110;
											assign node10462 = (inp[7]) ? node10474 : node10463;
												assign node10463 = (inp[11]) ? node10469 : node10464;
													assign node10464 = (inp[1]) ? node10466 : 4'b1110;
														assign node10466 = (inp[13]) ? 4'b0110 : 4'b0110;
													assign node10469 = (inp[1]) ? node10471 : 4'b0110;
														assign node10471 = (inp[6]) ? 4'b0110 : 4'b0110;
												assign node10474 = (inp[5]) ? node10476 : 4'b0111;
													assign node10476 = (inp[11]) ? 4'b1111 : node10477;
														assign node10477 = (inp[1]) ? 4'b0111 : 4'b0111;
										assign node10481 = (inp[6]) ? node10501 : node10482;
											assign node10482 = (inp[11]) ? node10494 : node10483;
												assign node10483 = (inp[1]) ? node10489 : node10484;
													assign node10484 = (inp[2]) ? 4'b0111 : node10485;
														assign node10485 = (inp[7]) ? 4'b0111 : 4'b1110;
													assign node10489 = (inp[13]) ? 4'b0111 : node10490;
														assign node10490 = (inp[7]) ? 4'b0110 : 4'b0111;
												assign node10494 = (inp[2]) ? 4'b1111 : node10495;
													assign node10495 = (inp[7]) ? 4'b0111 : node10496;
														assign node10496 = (inp[13]) ? 4'b0110 : 4'b0110;
											assign node10501 = (inp[13]) ? node10513 : node10502;
												assign node10502 = (inp[11]) ? node10508 : node10503;
													assign node10503 = (inp[5]) ? node10505 : 4'b0110;
														assign node10505 = (inp[2]) ? 4'b0111 : 4'b0110;
													assign node10508 = (inp[1]) ? 4'b0111 : node10509;
														assign node10509 = (inp[2]) ? 4'b1110 : 4'b1110;
												assign node10513 = (inp[11]) ? node10521 : node10514;
													assign node10514 = (inp[2]) ? node10518 : node10515;
														assign node10515 = (inp[7]) ? 4'b1111 : 4'b1110;
														assign node10518 = (inp[7]) ? 4'b1110 : 4'b1111;
													assign node10521 = (inp[1]) ? node10525 : node10522;
														assign node10522 = (inp[2]) ? 4'b0110 : 4'b1110;
														assign node10525 = (inp[7]) ? 4'b0110 : 4'b0110;
									assign node10528 = (inp[8]) ? node10564 : node10529;
										assign node10529 = (inp[7]) ? node10545 : node10530;
											assign node10530 = (inp[2]) ? node10540 : node10531;
												assign node10531 = (inp[6]) ? node10537 : node10532;
													assign node10532 = (inp[5]) ? 4'b1110 : node10533;
														assign node10533 = (inp[1]) ? 4'b0110 : 4'b1110;
													assign node10537 = (inp[11]) ? 4'b1110 : 4'b0110;
												assign node10540 = (inp[13]) ? 4'b1110 : node10541;
													assign node10541 = (inp[5]) ? 4'b0110 : 4'b1110;
											assign node10545 = (inp[6]) ? node10557 : node10546;
												assign node10546 = (inp[11]) ? node10552 : node10547;
													assign node10547 = (inp[13]) ? 4'b0111 : node10548;
														assign node10548 = (inp[1]) ? 4'b0111 : 4'b1111;
													assign node10552 = (inp[13]) ? 4'b1111 : node10553;
														assign node10553 = (inp[1]) ? 4'b1111 : 4'b0111;
												assign node10557 = (inp[11]) ? node10559 : 4'b1111;
													assign node10559 = (inp[13]) ? 4'b0111 : node10560;
														assign node10560 = (inp[1]) ? 4'b0111 : 4'b1111;
										assign node10564 = (inp[7]) ? node10586 : node10565;
											assign node10565 = (inp[6]) ? node10575 : node10566;
												assign node10566 = (inp[11]) ? node10572 : node10567;
													assign node10567 = (inp[1]) ? 4'b0111 : node10568;
														assign node10568 = (inp[13]) ? 4'b0111 : 4'b1111;
													assign node10572 = (inp[1]) ? 4'b1111 : 4'b0111;
												assign node10575 = (inp[11]) ? node10581 : node10576;
													assign node10576 = (inp[1]) ? 4'b1111 : node10577;
														assign node10577 = (inp[13]) ? 4'b1111 : 4'b0111;
													assign node10581 = (inp[1]) ? 4'b0111 : node10582;
														assign node10582 = (inp[13]) ? 4'b0111 : 4'b1111;
											assign node10586 = (inp[11]) ? node10598 : node10587;
												assign node10587 = (inp[6]) ? node10593 : node10588;
													assign node10588 = (inp[1]) ? 4'b0110 : node10589;
														assign node10589 = (inp[13]) ? 4'b0110 : 4'b1110;
													assign node10593 = (inp[13]) ? 4'b1110 : node10594;
														assign node10594 = (inp[1]) ? 4'b1110 : 4'b0110;
												assign node10598 = (inp[6]) ? 4'b0110 : node10599;
													assign node10599 = (inp[13]) ? 4'b1110 : 4'b0110;
						assign node10603 = (inp[10]) ? node10957 : node10604;
							assign node10604 = (inp[12]) ? node10790 : node10605;
								assign node10605 = (inp[5]) ? node10693 : node10606;
									assign node10606 = (inp[2]) ? node10646 : node10607;
										assign node10607 = (inp[6]) ? node10631 : node10608;
											assign node10608 = (inp[7]) ? node10620 : node10609;
												assign node10609 = (inp[8]) ? node10617 : node10610;
													assign node10610 = (inp[14]) ? node10614 : node10611;
														assign node10611 = (inp[1]) ? 4'b0111 : 4'b0111;
														assign node10614 = (inp[1]) ? 4'b1110 : 4'b0110;
													assign node10617 = (inp[14]) ? 4'b0111 : 4'b0110;
												assign node10620 = (inp[8]) ? node10626 : node10621;
													assign node10621 = (inp[14]) ? node10623 : 4'b0110;
														assign node10623 = (inp[1]) ? 4'b0111 : 4'b1111;
													assign node10626 = (inp[14]) ? node10628 : 4'b1111;
														assign node10628 = (inp[1]) ? 4'b0110 : 4'b1110;
											assign node10631 = (inp[11]) ? node10635 : node10632;
												assign node10632 = (inp[13]) ? 4'b1110 : 4'b0110;
												assign node10635 = (inp[1]) ? node10641 : node10636;
													assign node10636 = (inp[8]) ? node10638 : 4'b1110;
														assign node10638 = (inp[7]) ? 4'b1111 : 4'b1110;
													assign node10641 = (inp[7]) ? node10643 : 4'b1111;
														assign node10643 = (inp[14]) ? 4'b0110 : 4'b0110;
										assign node10646 = (inp[11]) ? node10670 : node10647;
											assign node10647 = (inp[6]) ? node10659 : node10648;
												assign node10648 = (inp[13]) ? node10654 : node10649;
													assign node10649 = (inp[7]) ? node10651 : 4'b1110;
														assign node10651 = (inp[1]) ? 4'b0111 : 4'b1111;
													assign node10654 = (inp[14]) ? 4'b0111 : node10655;
														assign node10655 = (inp[7]) ? 4'b0110 : 4'b0110;
												assign node10659 = (inp[8]) ? node10665 : node10660;
													assign node10660 = (inp[7]) ? 4'b1111 : node10661;
														assign node10661 = (inp[13]) ? 4'b1110 : 4'b0110;
													assign node10665 = (inp[7]) ? node10667 : 4'b1111;
														assign node10667 = (inp[1]) ? 4'b1110 : 4'b1110;
											assign node10670 = (inp[6]) ? node10682 : node10671;
												assign node10671 = (inp[1]) ? node10677 : node10672;
													assign node10672 = (inp[8]) ? node10674 : 4'b0110;
														assign node10674 = (inp[7]) ? 4'b1110 : 4'b0111;
													assign node10677 = (inp[7]) ? node10679 : 4'b1111;
														assign node10679 = (inp[8]) ? 4'b1110 : 4'b1111;
												assign node10682 = (inp[13]) ? node10686 : node10683;
													assign node10683 = (inp[1]) ? 4'b0110 : 4'b1110;
													assign node10686 = (inp[7]) ? node10690 : node10687;
														assign node10687 = (inp[8]) ? 4'b0111 : 4'b1110;
														assign node10690 = (inp[8]) ? 4'b0110 : 4'b0111;
									assign node10693 = (inp[11]) ? node10743 : node10694;
										assign node10694 = (inp[1]) ? node10720 : node10695;
											assign node10695 = (inp[7]) ? node10705 : node10696;
												assign node10696 = (inp[8]) ? node10700 : node10697;
													assign node10697 = (inp[2]) ? 4'b1110 : 4'b1111;
													assign node10700 = (inp[14]) ? 4'b1111 : node10701;
														assign node10701 = (inp[2]) ? 4'b0111 : 4'b0110;
												assign node10705 = (inp[8]) ? node10713 : node10706;
													assign node10706 = (inp[14]) ? node10710 : node10707;
														assign node10707 = (inp[13]) ? 4'b1111 : 4'b0110;
														assign node10710 = (inp[2]) ? 4'b0111 : 4'b1111;
													assign node10713 = (inp[2]) ? node10717 : node10714;
														assign node10714 = (inp[14]) ? 4'b0110 : 4'b1111;
														assign node10717 = (inp[6]) ? 4'b1110 : 4'b0110;
											assign node10720 = (inp[6]) ? node10732 : node10721;
												assign node10721 = (inp[8]) ? node10727 : node10722;
													assign node10722 = (inp[13]) ? 4'b0111 : node10723;
														assign node10723 = (inp[14]) ? 4'b1110 : 4'b0110;
													assign node10727 = (inp[14]) ? node10729 : 4'b0110;
														assign node10729 = (inp[7]) ? 4'b0110 : 4'b0111;
												assign node10732 = (inp[14]) ? node10738 : node10733;
													assign node10733 = (inp[8]) ? 4'b1111 : node10734;
														assign node10734 = (inp[7]) ? 4'b1111 : 4'b0110;
													assign node10738 = (inp[8]) ? node10740 : 4'b1111;
														assign node10740 = (inp[2]) ? 4'b1110 : 4'b1111;
										assign node10743 = (inp[8]) ? node10767 : node10744;
											assign node10744 = (inp[7]) ? node10756 : node10745;
												assign node10745 = (inp[6]) ? node10751 : node10746;
													assign node10746 = (inp[14]) ? 4'b0110 : node10747;
														assign node10747 = (inp[2]) ? 4'b1110 : 4'b0111;
													assign node10751 = (inp[14]) ? 4'b1110 : node10752;
														assign node10752 = (inp[2]) ? 4'b1110 : 4'b0111;
												assign node10756 = (inp[14]) ? node10762 : node10757;
													assign node10757 = (inp[2]) ? 4'b1111 : node10758;
														assign node10758 = (inp[6]) ? 4'b0110 : 4'b0110;
													assign node10762 = (inp[13]) ? 4'b0111 : node10763;
														assign node10763 = (inp[6]) ? 4'b0111 : 4'b1111;
											assign node10767 = (inp[7]) ? node10777 : node10768;
												assign node10768 = (inp[6]) ? node10772 : node10769;
													assign node10769 = (inp[14]) ? 4'b0111 : 4'b1111;
													assign node10772 = (inp[2]) ? 4'b0111 : node10773;
														assign node10773 = (inp[13]) ? 4'b0110 : 4'b0111;
												assign node10777 = (inp[14]) ? node10785 : node10778;
													assign node10778 = (inp[2]) ? node10782 : node10779;
														assign node10779 = (inp[6]) ? 4'b0111 : 4'b1111;
														assign node10782 = (inp[6]) ? 4'b0110 : 4'b1110;
													assign node10785 = (inp[1]) ? 4'b1110 : node10786;
														assign node10786 = (inp[13]) ? 4'b0110 : 4'b0110;
								assign node10790 = (inp[6]) ? node10880 : node10791;
									assign node10791 = (inp[11]) ? node10843 : node10792;
										assign node10792 = (inp[1]) ? node10816 : node10793;
											assign node10793 = (inp[13]) ? node10807 : node10794;
												assign node10794 = (inp[7]) ? node10802 : node10795;
													assign node10795 = (inp[8]) ? node10799 : node10796;
														assign node10796 = (inp[14]) ? 4'b1110 : 4'b1111;
														assign node10799 = (inp[5]) ? 4'b1110 : 4'b1111;
													assign node10802 = (inp[5]) ? 4'b1111 : node10803;
														assign node10803 = (inp[8]) ? 4'b1110 : 4'b1111;
												assign node10807 = (inp[7]) ? node10813 : node10808;
													assign node10808 = (inp[2]) ? 4'b0111 : node10809;
														assign node10809 = (inp[14]) ? 4'b1110 : 4'b1111;
													assign node10813 = (inp[2]) ? 4'b0110 : 4'b0111;
											assign node10816 = (inp[13]) ? node10828 : node10817;
												assign node10817 = (inp[7]) ? node10825 : node10818;
													assign node10818 = (inp[8]) ? node10822 : node10819;
														assign node10819 = (inp[2]) ? 4'b1110 : 4'b1111;
														assign node10822 = (inp[14]) ? 4'b0111 : 4'b0110;
													assign node10825 = (inp[8]) ? 4'b0110 : 4'b0111;
												assign node10828 = (inp[5]) ? node10836 : node10829;
													assign node10829 = (inp[8]) ? node10833 : node10830;
														assign node10830 = (inp[2]) ? 4'b0110 : 4'b0111;
														assign node10833 = (inp[7]) ? 4'b0110 : 4'b0111;
													assign node10836 = (inp[14]) ? node10840 : node10837;
														assign node10837 = (inp[2]) ? 4'b0110 : 4'b0110;
														assign node10840 = (inp[8]) ? 4'b0111 : 4'b0110;
										assign node10843 = (inp[13]) ? node10863 : node10844;
											assign node10844 = (inp[1]) ? node10856 : node10845;
												assign node10845 = (inp[2]) ? node10849 : node10846;
													assign node10846 = (inp[14]) ? 4'b0110 : 4'b0111;
													assign node10849 = (inp[7]) ? node10853 : node10850;
														assign node10850 = (inp[8]) ? 4'b0111 : 4'b0110;
														assign node10853 = (inp[8]) ? 4'b0110 : 4'b0111;
												assign node10856 = (inp[7]) ? 4'b1010 : node10857;
													assign node10857 = (inp[5]) ? 4'b0110 : node10858;
														assign node10858 = (inp[8]) ? 4'b0010 : 4'b0110;
											assign node10863 = (inp[2]) ? node10871 : node10864;
												assign node10864 = (inp[1]) ? node10866 : 4'b0110;
													assign node10866 = (inp[8]) ? 4'b1010 : node10867;
														assign node10867 = (inp[5]) ? 4'b1010 : 4'b1010;
												assign node10871 = (inp[14]) ? node10873 : 4'b1011;
													assign node10873 = (inp[5]) ? node10877 : node10874;
														assign node10874 = (inp[8]) ? 4'b1011 : 4'b1010;
														assign node10877 = (inp[8]) ? 4'b1010 : 4'b1010;
									assign node10880 = (inp[11]) ? node10918 : node10881;
										assign node10881 = (inp[1]) ? node10903 : node10882;
											assign node10882 = (inp[13]) ? node10894 : node10883;
												assign node10883 = (inp[7]) ? node10889 : node10884;
													assign node10884 = (inp[8]) ? 4'b0111 : node10885;
														assign node10885 = (inp[2]) ? 4'b0110 : 4'b0111;
													assign node10889 = (inp[8]) ? 4'b0110 : node10890;
														assign node10890 = (inp[14]) ? 4'b0111 : 4'b0110;
												assign node10894 = (inp[14]) ? node10900 : node10895;
													assign node10895 = (inp[8]) ? node10897 : 4'b0110;
														assign node10897 = (inp[7]) ? 4'b1010 : 4'b0010;
													assign node10900 = (inp[8]) ? 4'b1010 : 4'b1011;
											assign node10903 = (inp[8]) ? node10915 : node10904;
												assign node10904 = (inp[13]) ? node10912 : node10905;
													assign node10905 = (inp[7]) ? node10909 : node10906;
														assign node10906 = (inp[2]) ? 4'b0110 : 4'b0110;
														assign node10909 = (inp[2]) ? 4'b1011 : 4'b0110;
													assign node10912 = (inp[7]) ? 4'b1011 : 4'b1010;
												assign node10915 = (inp[7]) ? 4'b1010 : 4'b1011;
										assign node10918 = (inp[1]) ? node10934 : node10919;
											assign node10919 = (inp[7]) ? node10927 : node10920;
												assign node10920 = (inp[13]) ? 4'b1010 : node10921;
													assign node10921 = (inp[5]) ? 4'b1011 : node10922;
														assign node10922 = (inp[8]) ? 4'b1010 : 4'b1010;
												assign node10927 = (inp[13]) ? 4'b0011 : node10928;
													assign node10928 = (inp[8]) ? 4'b1010 : node10929;
														assign node10929 = (inp[14]) ? 4'b1011 : 4'b1010;
											assign node10934 = (inp[8]) ? node10946 : node10935;
												assign node10935 = (inp[7]) ? node10943 : node10936;
													assign node10936 = (inp[13]) ? node10940 : node10937;
														assign node10937 = (inp[14]) ? 4'b1010 : 4'b1011;
														assign node10940 = (inp[2]) ? 4'b0010 : 4'b0010;
													assign node10943 = (inp[14]) ? 4'b0011 : 4'b0010;
												assign node10946 = (inp[7]) ? node10952 : node10947;
													assign node10947 = (inp[2]) ? 4'b0011 : node10948;
														assign node10948 = (inp[13]) ? 4'b0010 : 4'b0011;
													assign node10952 = (inp[2]) ? 4'b0010 : node10953;
														assign node10953 = (inp[14]) ? 4'b0010 : 4'b0011;
							assign node10957 = (inp[12]) ? node11121 : node10958;
								assign node10958 = (inp[6]) ? node11044 : node10959;
									assign node10959 = (inp[11]) ? node10999 : node10960;
										assign node10960 = (inp[1]) ? node10978 : node10961;
											assign node10961 = (inp[13]) ? node10971 : node10962;
												assign node10962 = (inp[8]) ? node10968 : node10963;
													assign node10963 = (inp[7]) ? 4'b1111 : node10964;
														assign node10964 = (inp[5]) ? 4'b1110 : 4'b1110;
													assign node10968 = (inp[7]) ? 4'b1110 : 4'b1111;
												assign node10971 = (inp[14]) ? 4'b0111 : node10972;
													assign node10972 = (inp[8]) ? node10974 : 4'b1110;
														assign node10974 = (inp[7]) ? 4'b0110 : 4'b0111;
											assign node10978 = (inp[2]) ? node10988 : node10979;
												assign node10979 = (inp[13]) ? node10983 : node10980;
													assign node10980 = (inp[14]) ? 4'b1110 : 4'b0111;
													assign node10983 = (inp[5]) ? 4'b0111 : node10984;
														assign node10984 = (inp[7]) ? 4'b0110 : 4'b0111;
												assign node10988 = (inp[13]) ? node10994 : node10989;
													assign node10989 = (inp[8]) ? node10991 : 4'b0111;
														assign node10991 = (inp[7]) ? 4'b0110 : 4'b0111;
													assign node10994 = (inp[14]) ? 4'b0110 : node10995;
														assign node10995 = (inp[8]) ? 4'b0111 : 4'b0110;
										assign node10999 = (inp[1]) ? node11021 : node11000;
											assign node11000 = (inp[13]) ? node11012 : node11001;
												assign node11001 = (inp[14]) ? node11007 : node11002;
													assign node11002 = (inp[7]) ? node11004 : 4'b0111;
														assign node11004 = (inp[2]) ? 4'b0110 : 4'b0111;
													assign node11007 = (inp[8]) ? 4'b0110 : node11008;
														assign node11008 = (inp[2]) ? 4'b0111 : 4'b0110;
												assign node11012 = (inp[2]) ? node11018 : node11013;
													assign node11013 = (inp[14]) ? node11015 : 4'b0110;
														assign node11015 = (inp[5]) ? 4'b1011 : 4'b0110;
													assign node11018 = (inp[5]) ? 4'b1010 : 4'b1011;
											assign node11021 = (inp[8]) ? node11033 : node11022;
												assign node11022 = (inp[7]) ? node11028 : node11023;
													assign node11023 = (inp[2]) ? 4'b0110 : node11024;
														assign node11024 = (inp[5]) ? 4'b1010 : 4'b1011;
													assign node11028 = (inp[14]) ? 4'b1011 : node11029;
														assign node11029 = (inp[2]) ? 4'b1011 : 4'b0110;
												assign node11033 = (inp[7]) ? node11039 : node11034;
													assign node11034 = (inp[14]) ? 4'b1011 : node11035;
														assign node11035 = (inp[2]) ? 4'b1011 : 4'b1010;
													assign node11039 = (inp[14]) ? 4'b1010 : node11040;
														assign node11040 = (inp[2]) ? 4'b1010 : 4'b1011;
									assign node11044 = (inp[11]) ? node11076 : node11045;
										assign node11045 = (inp[1]) ? node11063 : node11046;
											assign node11046 = (inp[13]) ? node11052 : node11047;
												assign node11047 = (inp[2]) ? node11049 : 4'b0110;
													assign node11049 = (inp[7]) ? 4'b0111 : 4'b0110;
												assign node11052 = (inp[8]) ? node11058 : node11053;
													assign node11053 = (inp[7]) ? 4'b1011 : node11054;
														assign node11054 = (inp[2]) ? 4'b0110 : 4'b0111;
													assign node11058 = (inp[14]) ? 4'b1010 : node11059;
														assign node11059 = (inp[7]) ? 4'b1010 : 4'b1011;
											assign node11063 = (inp[8]) ? node11071 : node11064;
												assign node11064 = (inp[7]) ? 4'b1011 : node11065;
													assign node11065 = (inp[13]) ? node11067 : 4'b0111;
														assign node11067 = (inp[2]) ? 4'b1010 : 4'b1011;
												assign node11071 = (inp[7]) ? 4'b1010 : node11072;
													assign node11072 = (inp[14]) ? 4'b1011 : 4'b1010;
										assign node11076 = (inp[1]) ? node11104 : node11077;
											assign node11077 = (inp[13]) ? node11091 : node11078;
												assign node11078 = (inp[5]) ? node11086 : node11079;
													assign node11079 = (inp[8]) ? node11083 : node11080;
														assign node11080 = (inp[2]) ? 4'b1010 : 4'b1011;
														assign node11083 = (inp[2]) ? 4'b1010 : 4'b1010;
													assign node11086 = (inp[8]) ? 4'b1011 : node11087;
														assign node11087 = (inp[7]) ? 4'b1011 : 4'b1010;
												assign node11091 = (inp[2]) ? node11097 : node11092;
													assign node11092 = (inp[14]) ? 4'b0011 : node11093;
														assign node11093 = (inp[8]) ? 4'b1010 : 4'b1010;
													assign node11097 = (inp[8]) ? node11101 : node11098;
														assign node11098 = (inp[7]) ? 4'b0011 : 4'b1010;
														assign node11101 = (inp[7]) ? 4'b0010 : 4'b0011;
											assign node11104 = (inp[13]) ? node11114 : node11105;
												assign node11105 = (inp[8]) ? node11107 : 4'b0011;
													assign node11107 = (inp[14]) ? node11111 : node11108;
														assign node11108 = (inp[5]) ? 4'b1010 : 4'b0011;
														assign node11111 = (inp[5]) ? 4'b0011 : 4'b0010;
												assign node11114 = (inp[7]) ? 4'b0010 : node11115;
													assign node11115 = (inp[2]) ? 4'b0010 : node11116;
														assign node11116 = (inp[14]) ? 4'b0010 : 4'b0010;
								assign node11121 = (inp[7]) ? node11199 : node11122;
									assign node11122 = (inp[8]) ? node11156 : node11123;
										assign node11123 = (inp[2]) ? node11139 : node11124;
											assign node11124 = (inp[14]) ? node11132 : node11125;
												assign node11125 = (inp[11]) ? 4'b0011 : node11126;
													assign node11126 = (inp[5]) ? node11128 : 4'b1011;
														assign node11128 = (inp[6]) ? 4'b0011 : 4'b1011;
												assign node11132 = (inp[1]) ? node11134 : 4'b1010;
													assign node11134 = (inp[13]) ? 4'b0010 : node11135;
														assign node11135 = (inp[5]) ? 4'b0010 : 4'b1010;
											assign node11139 = (inp[6]) ? node11147 : node11140;
												assign node11140 = (inp[13]) ? node11142 : 4'b0010;
													assign node11142 = (inp[5]) ? 4'b0010 : node11143;
														assign node11143 = (inp[14]) ? 4'b1010 : 4'b0010;
												assign node11147 = (inp[11]) ? node11151 : node11148;
													assign node11148 = (inp[5]) ? 4'b1010 : 4'b0010;
													assign node11151 = (inp[1]) ? node11153 : 4'b1010;
														assign node11153 = (inp[13]) ? 4'b0010 : 4'b1010;
										assign node11156 = (inp[2]) ? node11178 : node11157;
											assign node11157 = (inp[14]) ? node11165 : node11158;
												assign node11158 = (inp[5]) ? node11160 : 4'b0010;
													assign node11160 = (inp[11]) ? 4'b1010 : node11161;
														assign node11161 = (inp[13]) ? 4'b1010 : 4'b0010;
												assign node11165 = (inp[13]) ? node11173 : node11166;
													assign node11166 = (inp[5]) ? node11170 : node11167;
														assign node11167 = (inp[11]) ? 4'b0011 : 4'b0011;
														assign node11170 = (inp[11]) ? 4'b1011 : 4'b0011;
													assign node11173 = (inp[1]) ? 4'b1011 : node11174;
														assign node11174 = (inp[11]) ? 4'b0011 : 4'b1011;
											assign node11178 = (inp[1]) ? node11192 : node11179;
												assign node11179 = (inp[11]) ? node11187 : node11180;
													assign node11180 = (inp[13]) ? node11184 : node11181;
														assign node11181 = (inp[6]) ? 4'b0011 : 4'b1011;
														assign node11184 = (inp[6]) ? 4'b1011 : 4'b0011;
													assign node11187 = (inp[5]) ? 4'b1011 : node11188;
														assign node11188 = (inp[6]) ? 4'b0011 : 4'b1011;
												assign node11192 = (inp[6]) ? node11196 : node11193;
													assign node11193 = (inp[11]) ? 4'b1011 : 4'b0011;
													assign node11196 = (inp[11]) ? 4'b0011 : 4'b1011;
									assign node11199 = (inp[8]) ? node11239 : node11200;
										assign node11200 = (inp[14]) ? node11224 : node11201;
											assign node11201 = (inp[2]) ? node11215 : node11202;
												assign node11202 = (inp[5]) ? node11208 : node11203;
													assign node11203 = (inp[6]) ? node11205 : 4'b0010;
														assign node11205 = (inp[11]) ? 4'b1010 : 4'b0010;
													assign node11208 = (inp[13]) ? node11212 : node11209;
														assign node11209 = (inp[1]) ? 4'b0010 : 4'b1010;
														assign node11212 = (inp[6]) ? 4'b0010 : 4'b0010;
												assign node11215 = (inp[11]) ? node11219 : node11216;
													assign node11216 = (inp[6]) ? 4'b1011 : 4'b0011;
													assign node11219 = (inp[6]) ? 4'b0011 : node11220;
														assign node11220 = (inp[5]) ? 4'b0011 : 4'b1011;
											assign node11224 = (inp[6]) ? node11232 : node11225;
												assign node11225 = (inp[11]) ? node11229 : node11226;
													assign node11226 = (inp[1]) ? 4'b0011 : 4'b1011;
													assign node11229 = (inp[1]) ? 4'b1011 : 4'b0011;
												assign node11232 = (inp[11]) ? node11234 : 4'b1011;
													assign node11234 = (inp[13]) ? 4'b0011 : node11235;
														assign node11235 = (inp[1]) ? 4'b0011 : 4'b1011;
										assign node11239 = (inp[2]) ? node11255 : node11240;
											assign node11240 = (inp[14]) ? node11246 : node11241;
												assign node11241 = (inp[11]) ? 4'b0011 : node11242;
													assign node11242 = (inp[1]) ? 4'b1011 : 4'b0011;
												assign node11246 = (inp[5]) ? 4'b0010 : node11247;
													assign node11247 = (inp[11]) ? node11251 : node11248;
														assign node11248 = (inp[6]) ? 4'b0010 : 4'b0010;
														assign node11251 = (inp[6]) ? 4'b0010 : 4'b1010;
											assign node11255 = (inp[11]) ? node11261 : node11256;
												assign node11256 = (inp[6]) ? node11258 : 4'b0010;
													assign node11258 = (inp[14]) ? 4'b0010 : 4'b1010;
												assign node11261 = (inp[6]) ? node11267 : node11262;
													assign node11262 = (inp[1]) ? 4'b1010 : node11263;
														assign node11263 = (inp[13]) ? 4'b1010 : 4'b0010;
													assign node11267 = (inp[1]) ? 4'b0010 : 4'b1010;
		assign node11270 = (inp[6]) ? node16998 : node11271;
			assign node11271 = (inp[11]) ? node14091 : node11272;
				assign node11272 = (inp[13]) ? node12692 : node11273;
					assign node11273 = (inp[1]) ? node12001 : node11274;
						assign node11274 = (inp[15]) ? node11624 : node11275;
							assign node11275 = (inp[5]) ? node11449 : node11276;
								assign node11276 = (inp[3]) ? node11362 : node11277;
									assign node11277 = (inp[8]) ? node11323 : node11278;
										assign node11278 = (inp[7]) ? node11304 : node11279;
											assign node11279 = (inp[14]) ? node11291 : node11280;
												assign node11280 = (inp[2]) ? node11286 : node11281;
													assign node11281 = (inp[10]) ? 4'b1101 : node11282;
														assign node11282 = (inp[9]) ? 4'b1001 : 4'b1001;
													assign node11286 = (inp[12]) ? node11288 : 4'b1000;
														assign node11288 = (inp[10]) ? 4'b1100 : 4'b1000;
												assign node11291 = (inp[9]) ? node11297 : node11292;
													assign node11292 = (inp[4]) ? 4'b1000 : node11293;
														assign node11293 = (inp[10]) ? 4'b1000 : 4'b1100;
													assign node11297 = (inp[4]) ? node11301 : node11298;
														assign node11298 = (inp[10]) ? 4'b1000 : 4'b1000;
														assign node11301 = (inp[2]) ? 4'b1100 : 4'b1000;
											assign node11304 = (inp[14]) ? node11316 : node11305;
												assign node11305 = (inp[2]) ? node11311 : node11306;
													assign node11306 = (inp[10]) ? 4'b1100 : node11307;
														assign node11307 = (inp[12]) ? 4'b1100 : 4'b1000;
													assign node11311 = (inp[12]) ? node11313 : 4'b1001;
														assign node11313 = (inp[10]) ? 4'b1101 : 4'b1001;
												assign node11316 = (inp[12]) ? 4'b1101 : node11317;
													assign node11317 = (inp[10]) ? 4'b1001 : node11318;
														assign node11318 = (inp[9]) ? 4'b1101 : 4'b1001;
										assign node11323 = (inp[7]) ? node11345 : node11324;
											assign node11324 = (inp[2]) ? node11336 : node11325;
												assign node11325 = (inp[14]) ? node11331 : node11326;
													assign node11326 = (inp[10]) ? 4'b1000 : node11327;
														assign node11327 = (inp[12]) ? 4'b1000 : 4'b1100;
													assign node11331 = (inp[10]) ? node11333 : 4'b1101;
														assign node11333 = (inp[4]) ? 4'b1001 : 4'b1101;
												assign node11336 = (inp[4]) ? node11342 : node11337;
													assign node11337 = (inp[9]) ? node11339 : 4'b1101;
														assign node11339 = (inp[10]) ? 4'b1101 : 4'b1001;
													assign node11342 = (inp[9]) ? 4'b1101 : 4'b1001;
											assign node11345 = (inp[14]) ? node11355 : node11346;
												assign node11346 = (inp[2]) ? node11352 : node11347;
													assign node11347 = (inp[4]) ? 4'b1101 : node11348;
														assign node11348 = (inp[10]) ? 4'b1101 : 4'b1001;
													assign node11352 = (inp[12]) ? 4'b1000 : 4'b1100;
												assign node11355 = (inp[10]) ? 4'b1100 : node11356;
													assign node11356 = (inp[12]) ? node11358 : 4'b1000;
														assign node11358 = (inp[9]) ? 4'b1100 : 4'b1000;
									assign node11362 = (inp[4]) ? node11408 : node11363;
										assign node11363 = (inp[9]) ? node11387 : node11364;
											assign node11364 = (inp[10]) ? node11374 : node11365;
												assign node11365 = (inp[2]) ? node11369 : node11366;
													assign node11366 = (inp[8]) ? 4'b1101 : 4'b1100;
													assign node11369 = (inp[8]) ? node11371 : 4'b1101;
														assign node11371 = (inp[7]) ? 4'b1100 : 4'b1101;
												assign node11374 = (inp[12]) ? node11380 : node11375;
													assign node11375 = (inp[14]) ? 4'b1101 : node11376;
														assign node11376 = (inp[7]) ? 4'b1100 : 4'b1101;
													assign node11380 = (inp[8]) ? node11384 : node11381;
														assign node11381 = (inp[2]) ? 4'b1000 : 4'b1001;
														assign node11384 = (inp[2]) ? 4'b1001 : 4'b1000;
											assign node11387 = (inp[12]) ? node11399 : node11388;
												assign node11388 = (inp[7]) ? node11394 : node11389;
													assign node11389 = (inp[2]) ? node11391 : 4'b1000;
														assign node11391 = (inp[14]) ? 4'b1001 : 4'b1000;
													assign node11394 = (inp[8]) ? node11396 : 4'b1001;
														assign node11396 = (inp[14]) ? 4'b1000 : 4'b1001;
												assign node11399 = (inp[10]) ? node11405 : node11400;
													assign node11400 = (inp[14]) ? node11402 : 4'b1001;
														assign node11402 = (inp[7]) ? 4'b1000 : 4'b1000;
													assign node11405 = (inp[14]) ? 4'b1110 : 4'b1111;
										assign node11408 = (inp[9]) ? node11424 : node11409;
											assign node11409 = (inp[12]) ? node11419 : node11410;
												assign node11410 = (inp[7]) ? node11414 : node11411;
													assign node11411 = (inp[8]) ? 4'b1001 : 4'b1000;
													assign node11414 = (inp[14]) ? 4'b1001 : node11415;
														assign node11415 = (inp[2]) ? 4'b1001 : 4'b1000;
												assign node11419 = (inp[10]) ? node11421 : 4'b1000;
													assign node11421 = (inp[2]) ? 4'b1110 : 4'b1111;
											assign node11424 = (inp[12]) ? node11436 : node11425;
												assign node11425 = (inp[2]) ? node11431 : node11426;
													assign node11426 = (inp[7]) ? 4'b1111 : node11427;
														assign node11427 = (inp[10]) ? 4'b1110 : 4'b1110;
													assign node11431 = (inp[14]) ? 4'b1111 : node11432;
														assign node11432 = (inp[8]) ? 4'b1110 : 4'b1111;
												assign node11436 = (inp[10]) ? node11444 : node11437;
													assign node11437 = (inp[2]) ? node11441 : node11438;
														assign node11438 = (inp[7]) ? 4'b1111 : 4'b1110;
														assign node11441 = (inp[14]) ? 4'b1111 : 4'b1110;
													assign node11444 = (inp[14]) ? 4'b1011 : node11445;
														assign node11445 = (inp[2]) ? 4'b1010 : 4'b1010;
								assign node11449 = (inp[3]) ? node11539 : node11450;
									assign node11450 = (inp[9]) ? node11496 : node11451;
										assign node11451 = (inp[4]) ? node11477 : node11452;
											assign node11452 = (inp[12]) ? node11464 : node11453;
												assign node11453 = (inp[10]) ? node11459 : node11454;
													assign node11454 = (inp[8]) ? 4'b1100 : node11455;
														assign node11455 = (inp[2]) ? 4'b1101 : 4'b1100;
													assign node11459 = (inp[7]) ? 4'b1100 : node11460;
														assign node11460 = (inp[14]) ? 4'b1100 : 4'b1100;
												assign node11464 = (inp[10]) ? node11470 : node11465;
													assign node11465 = (inp[14]) ? node11467 : 4'b1101;
														assign node11467 = (inp[2]) ? 4'b1100 : 4'b1101;
													assign node11470 = (inp[2]) ? node11474 : node11471;
														assign node11471 = (inp[8]) ? 4'b1000 : 4'b1000;
														assign node11474 = (inp[7]) ? 4'b1000 : 4'b1001;
											assign node11477 = (inp[10]) ? node11489 : node11478;
												assign node11478 = (inp[12]) ? node11484 : node11479;
													assign node11479 = (inp[2]) ? node11481 : 4'b1000;
														assign node11481 = (inp[8]) ? 4'b1000 : 4'b1001;
													assign node11484 = (inp[2]) ? 4'b1001 : node11485;
														assign node11485 = (inp[7]) ? 4'b1001 : 4'b1000;
												assign node11489 = (inp[12]) ? node11491 : 4'b1001;
													assign node11491 = (inp[7]) ? node11493 : 4'b1110;
														assign node11493 = (inp[2]) ? 4'b1111 : 4'b1111;
										assign node11496 = (inp[4]) ? node11518 : node11497;
											assign node11497 = (inp[10]) ? node11511 : node11498;
												assign node11498 = (inp[14]) ? node11506 : node11499;
													assign node11499 = (inp[7]) ? node11503 : node11500;
														assign node11500 = (inp[2]) ? 4'b1001 : 4'b1000;
														assign node11503 = (inp[12]) ? 4'b1001 : 4'b1001;
													assign node11506 = (inp[12]) ? node11508 : 4'b1000;
														assign node11508 = (inp[7]) ? 4'b1000 : 4'b1000;
												assign node11511 = (inp[7]) ? 4'b1111 : node11512;
													assign node11512 = (inp[14]) ? 4'b1110 : node11513;
														assign node11513 = (inp[2]) ? 4'b1110 : 4'b1111;
											assign node11518 = (inp[10]) ? node11528 : node11519;
												assign node11519 = (inp[7]) ? node11525 : node11520;
													assign node11520 = (inp[8]) ? 4'b1111 : node11521;
														assign node11521 = (inp[14]) ? 4'b1110 : 4'b1111;
													assign node11525 = (inp[8]) ? 4'b1110 : 4'b1111;
												assign node11528 = (inp[12]) ? node11534 : node11529;
													assign node11529 = (inp[8]) ? node11531 : 4'b1111;
														assign node11531 = (inp[7]) ? 4'b1110 : 4'b1111;
													assign node11534 = (inp[8]) ? 4'b1010 : node11535;
														assign node11535 = (inp[2]) ? 4'b1010 : 4'b1010;
									assign node11539 = (inp[4]) ? node11581 : node11540;
										assign node11540 = (inp[9]) ? node11564 : node11541;
											assign node11541 = (inp[10]) ? node11553 : node11542;
												assign node11542 = (inp[8]) ? node11550 : node11543;
													assign node11543 = (inp[2]) ? node11547 : node11544;
														assign node11544 = (inp[12]) ? 4'b1110 : 4'b1111;
														assign node11547 = (inp[7]) ? 4'b1111 : 4'b1110;
													assign node11550 = (inp[7]) ? 4'b1110 : 4'b1111;
												assign node11553 = (inp[12]) ? node11559 : node11554;
													assign node11554 = (inp[7]) ? node11556 : 4'b1110;
														assign node11556 = (inp[8]) ? 4'b1110 : 4'b1110;
													assign node11559 = (inp[14]) ? 4'b1010 : node11560;
														assign node11560 = (inp[8]) ? 4'b1010 : 4'b1010;
											assign node11564 = (inp[10]) ? node11572 : node11565;
												assign node11565 = (inp[2]) ? node11567 : 4'b1010;
													assign node11567 = (inp[8]) ? node11569 : 4'b1011;
														assign node11569 = (inp[7]) ? 4'b1010 : 4'b1011;
												assign node11572 = (inp[12]) ? node11576 : node11573;
													assign node11573 = (inp[7]) ? 4'b1010 : 4'b1011;
													assign node11576 = (inp[14]) ? node11578 : 4'b1111;
														assign node11578 = (inp[7]) ? 4'b1110 : 4'b1111;
										assign node11581 = (inp[9]) ? node11605 : node11582;
											assign node11582 = (inp[10]) ? node11594 : node11583;
												assign node11583 = (inp[8]) ? node11589 : node11584;
													assign node11584 = (inp[7]) ? 4'b1011 : node11585;
														assign node11585 = (inp[12]) ? 4'b1010 : 4'b1011;
													assign node11589 = (inp[7]) ? node11591 : 4'b1011;
														assign node11591 = (inp[12]) ? 4'b1011 : 4'b1010;
												assign node11594 = (inp[12]) ? node11600 : node11595;
													assign node11595 = (inp[7]) ? node11597 : 4'b1011;
														assign node11597 = (inp[14]) ? 4'b1010 : 4'b1011;
													assign node11600 = (inp[14]) ? 4'b1111 : node11601;
														assign node11601 = (inp[7]) ? 4'b1110 : 4'b1111;
											assign node11605 = (inp[10]) ? node11617 : node11606;
												assign node11606 = (inp[12]) ? node11612 : node11607;
													assign node11607 = (inp[7]) ? 4'b1111 : node11608;
														assign node11608 = (inp[8]) ? 4'b1111 : 4'b1110;
													assign node11612 = (inp[14]) ? 4'b1110 : node11613;
														assign node11613 = (inp[7]) ? 4'b1110 : 4'b1111;
												assign node11617 = (inp[12]) ? 4'b1011 : node11618;
													assign node11618 = (inp[7]) ? 4'b1111 : node11619;
														assign node11619 = (inp[14]) ? 4'b1110 : 4'b1111;
							assign node11624 = (inp[3]) ? node11828 : node11625;
								assign node11625 = (inp[5]) ? node11729 : node11626;
									assign node11626 = (inp[12]) ? node11676 : node11627;
										assign node11627 = (inp[8]) ? node11653 : node11628;
											assign node11628 = (inp[7]) ? node11644 : node11629;
												assign node11629 = (inp[2]) ? node11637 : node11630;
													assign node11630 = (inp[14]) ? node11634 : node11631;
														assign node11631 = (inp[10]) ? 4'b1011 : 4'b1111;
														assign node11634 = (inp[10]) ? 4'b1010 : 4'b1110;
													assign node11637 = (inp[9]) ? node11641 : node11638;
														assign node11638 = (inp[4]) ? 4'b1010 : 4'b1110;
														assign node11641 = (inp[4]) ? 4'b1110 : 4'b1010;
												assign node11644 = (inp[2]) ? node11648 : node11645;
													assign node11645 = (inp[9]) ? 4'b1110 : 4'b1010;
													assign node11648 = (inp[9]) ? node11650 : 4'b1111;
														assign node11650 = (inp[4]) ? 4'b1111 : 4'b1011;
											assign node11653 = (inp[4]) ? node11667 : node11654;
												assign node11654 = (inp[9]) ? node11662 : node11655;
													assign node11655 = (inp[2]) ? node11659 : node11656;
														assign node11656 = (inp[7]) ? 4'b1111 : 4'b1110;
														assign node11659 = (inp[7]) ? 4'b1110 : 4'b1111;
													assign node11662 = (inp[7]) ? 4'b1010 : node11663;
														assign node11663 = (inp[14]) ? 4'b1011 : 4'b1010;
												assign node11667 = (inp[9]) ? node11671 : node11668;
													assign node11668 = (inp[14]) ? 4'b1010 : 4'b1011;
													assign node11671 = (inp[7]) ? node11673 : 4'b1111;
														assign node11673 = (inp[14]) ? 4'b1110 : 4'b1111;
										assign node11676 = (inp[2]) ? node11702 : node11677;
											assign node11677 = (inp[4]) ? node11687 : node11678;
												assign node11678 = (inp[10]) ? node11682 : node11679;
													assign node11679 = (inp[9]) ? 4'b1011 : 4'b1111;
													assign node11682 = (inp[9]) ? node11684 : 4'b1011;
														assign node11684 = (inp[7]) ? 4'b1111 : 4'b1110;
												assign node11687 = (inp[14]) ? node11695 : node11688;
													assign node11688 = (inp[10]) ? node11692 : node11689;
														assign node11689 = (inp[9]) ? 4'b1111 : 4'b1010;
														assign node11692 = (inp[9]) ? 4'b1011 : 4'b1111;
													assign node11695 = (inp[8]) ? node11699 : node11696;
														assign node11696 = (inp[7]) ? 4'b1011 : 4'b1010;
														assign node11699 = (inp[7]) ? 4'b1010 : 4'b1011;
											assign node11702 = (inp[9]) ? node11714 : node11703;
												assign node11703 = (inp[8]) ? node11709 : node11704;
													assign node11704 = (inp[7]) ? node11706 : 4'b1110;
														assign node11706 = (inp[10]) ? 4'b1111 : 4'b1011;
													assign node11709 = (inp[7]) ? node11711 : 4'b1011;
														assign node11711 = (inp[4]) ? 4'b1010 : 4'b1110;
												assign node11714 = (inp[14]) ? node11722 : node11715;
													assign node11715 = (inp[4]) ? node11719 : node11716;
														assign node11716 = (inp[10]) ? 4'b1110 : 4'b1010;
														assign node11719 = (inp[10]) ? 4'b1010 : 4'b1110;
													assign node11722 = (inp[7]) ? node11726 : node11723;
														assign node11723 = (inp[8]) ? 4'b1011 : 4'b1010;
														assign node11726 = (inp[10]) ? 4'b1010 : 4'b1011;
									assign node11729 = (inp[4]) ? node11783 : node11730;
										assign node11730 = (inp[9]) ? node11754 : node11731;
											assign node11731 = (inp[12]) ? node11743 : node11732;
												assign node11732 = (inp[10]) ? node11738 : node11733;
													assign node11733 = (inp[8]) ? 4'b1110 : node11734;
														assign node11734 = (inp[7]) ? 4'b1111 : 4'b1110;
													assign node11738 = (inp[2]) ? node11740 : 4'b1111;
														assign node11740 = (inp[8]) ? 4'b1110 : 4'b1110;
												assign node11743 = (inp[10]) ? node11749 : node11744;
													assign node11744 = (inp[14]) ? node11746 : 4'b1111;
														assign node11746 = (inp[8]) ? 4'b1111 : 4'b1110;
													assign node11749 = (inp[2]) ? node11751 : 4'b1011;
														assign node11751 = (inp[14]) ? 4'b1011 : 4'b1010;
											assign node11754 = (inp[12]) ? node11770 : node11755;
												assign node11755 = (inp[10]) ? node11763 : node11756;
													assign node11756 = (inp[2]) ? node11760 : node11757;
														assign node11757 = (inp[7]) ? 4'b1010 : 4'b1010;
														assign node11760 = (inp[7]) ? 4'b1010 : 4'b1010;
													assign node11763 = (inp[14]) ? node11767 : node11764;
														assign node11764 = (inp[7]) ? 4'b1011 : 4'b1010;
														assign node11767 = (inp[2]) ? 4'b1010 : 4'b1011;
												assign node11770 = (inp[10]) ? node11776 : node11771;
													assign node11771 = (inp[2]) ? 4'b1010 : node11772;
														assign node11772 = (inp[8]) ? 4'b1010 : 4'b1011;
													assign node11776 = (inp[14]) ? node11780 : node11777;
														assign node11777 = (inp[7]) ? 4'b1100 : 4'b1101;
														assign node11780 = (inp[2]) ? 4'b1101 : 4'b1100;
										assign node11783 = (inp[9]) ? node11807 : node11784;
											assign node11784 = (inp[10]) ? node11796 : node11785;
												assign node11785 = (inp[8]) ? node11791 : node11786;
													assign node11786 = (inp[12]) ? 4'b1010 : node11787;
														assign node11787 = (inp[7]) ? 4'b1011 : 4'b1010;
													assign node11791 = (inp[7]) ? node11793 : 4'b1011;
														assign node11793 = (inp[14]) ? 4'b1010 : 4'b1010;
												assign node11796 = (inp[12]) ? node11802 : node11797;
													assign node11797 = (inp[2]) ? 4'b1010 : node11798;
														assign node11798 = (inp[7]) ? 4'b1010 : 4'b1011;
													assign node11802 = (inp[8]) ? 4'b1100 : node11803;
														assign node11803 = (inp[7]) ? 4'b1101 : 4'b1100;
											assign node11807 = (inp[12]) ? node11819 : node11808;
												assign node11808 = (inp[8]) ? node11814 : node11809;
													assign node11809 = (inp[7]) ? 4'b1101 : node11810;
														assign node11810 = (inp[2]) ? 4'b1100 : 4'b1101;
													assign node11814 = (inp[7]) ? 4'b1100 : node11815;
														assign node11815 = (inp[14]) ? 4'b1101 : 4'b1100;
												assign node11819 = (inp[10]) ? node11825 : node11820;
													assign node11820 = (inp[7]) ? 4'b1101 : node11821;
														assign node11821 = (inp[14]) ? 4'b1100 : 4'b1101;
													assign node11825 = (inp[8]) ? 4'b1000 : 4'b1001;
								assign node11828 = (inp[5]) ? node11918 : node11829;
									assign node11829 = (inp[4]) ? node11869 : node11830;
										assign node11830 = (inp[9]) ? node11852 : node11831;
											assign node11831 = (inp[10]) ? node11843 : node11832;
												assign node11832 = (inp[12]) ? node11838 : node11833;
													assign node11833 = (inp[7]) ? node11835 : 4'b1110;
														assign node11835 = (inp[8]) ? 4'b1110 : 4'b1111;
													assign node11838 = (inp[14]) ? node11840 : 4'b1111;
														assign node11840 = (inp[8]) ? 4'b1110 : 4'b1111;
												assign node11843 = (inp[12]) ? node11847 : node11844;
													assign node11844 = (inp[14]) ? 4'b1110 : 4'b1111;
													assign node11847 = (inp[14]) ? node11849 : 4'b1010;
														assign node11849 = (inp[2]) ? 4'b1010 : 4'b1011;
											assign node11852 = (inp[10]) ? node11864 : node11853;
												assign node11853 = (inp[7]) ? node11859 : node11854;
													assign node11854 = (inp[8]) ? 4'b1011 : node11855;
														assign node11855 = (inp[2]) ? 4'b1010 : 4'b1010;
													assign node11859 = (inp[8]) ? 4'b1010 : node11860;
														assign node11860 = (inp[12]) ? 4'b1011 : 4'b1010;
												assign node11864 = (inp[12]) ? 4'b1101 : node11865;
													assign node11865 = (inp[14]) ? 4'b1011 : 4'b1010;
										assign node11869 = (inp[9]) ? node11893 : node11870;
											assign node11870 = (inp[12]) ? node11882 : node11871;
												assign node11871 = (inp[7]) ? node11877 : node11872;
													assign node11872 = (inp[14]) ? node11874 : 4'b1011;
														assign node11874 = (inp[8]) ? 4'b1011 : 4'b1010;
													assign node11877 = (inp[8]) ? 4'b1010 : node11878;
														assign node11878 = (inp[2]) ? 4'b1011 : 4'b1010;
												assign node11882 = (inp[10]) ? node11886 : node11883;
													assign node11883 = (inp[2]) ? 4'b1010 : 4'b1011;
													assign node11886 = (inp[7]) ? node11890 : node11887;
														assign node11887 = (inp[8]) ? 4'b1100 : 4'b1100;
														assign node11890 = (inp[8]) ? 4'b1101 : 4'b1101;
											assign node11893 = (inp[10]) ? node11907 : node11894;
												assign node11894 = (inp[2]) ? node11900 : node11895;
													assign node11895 = (inp[8]) ? node11897 : 4'b1101;
														assign node11897 = (inp[12]) ? 4'b1100 : 4'b1101;
													assign node11900 = (inp[8]) ? node11904 : node11901;
														assign node11901 = (inp[7]) ? 4'b1101 : 4'b1100;
														assign node11904 = (inp[7]) ? 4'b1100 : 4'b1101;
												assign node11907 = (inp[12]) ? node11913 : node11908;
													assign node11908 = (inp[7]) ? 4'b1101 : node11909;
														assign node11909 = (inp[2]) ? 4'b1101 : 4'b1100;
													assign node11913 = (inp[14]) ? 4'b1001 : node11914;
														assign node11914 = (inp[7]) ? 4'b1000 : 4'b1001;
									assign node11918 = (inp[7]) ? node11960 : node11919;
										assign node11919 = (inp[8]) ? node11939 : node11920;
											assign node11920 = (inp[14]) ? node11932 : node11921;
												assign node11921 = (inp[2]) ? node11927 : node11922;
													assign node11922 = (inp[4]) ? node11924 : 4'b1101;
														assign node11924 = (inp[12]) ? 4'b1001 : 4'b1101;
													assign node11927 = (inp[12]) ? 4'b1100 : node11928;
														assign node11928 = (inp[10]) ? 4'b1000 : 4'b1000;
												assign node11932 = (inp[4]) ? node11936 : node11933;
													assign node11933 = (inp[9]) ? 4'b1000 : 4'b1100;
													assign node11936 = (inp[9]) ? 4'b1100 : 4'b1000;
											assign node11939 = (inp[14]) ? node11947 : node11940;
												assign node11940 = (inp[2]) ? node11944 : node11941;
													assign node11941 = (inp[4]) ? 4'b1000 : 4'b1100;
													assign node11944 = (inp[12]) ? 4'b1101 : 4'b1001;
												assign node11947 = (inp[12]) ? node11955 : node11948;
													assign node11948 = (inp[10]) ? node11952 : node11949;
														assign node11949 = (inp[9]) ? 4'b1101 : 4'b1101;
														assign node11952 = (inp[9]) ? 4'b1001 : 4'b1101;
													assign node11955 = (inp[9]) ? 4'b1001 : node11956;
														assign node11956 = (inp[10]) ? 4'b1001 : 4'b1001;
										assign node11960 = (inp[8]) ? node11980 : node11961;
											assign node11961 = (inp[14]) ? node11971 : node11962;
												assign node11962 = (inp[2]) ? node11968 : node11963;
													assign node11963 = (inp[10]) ? 4'b1000 : node11964;
														assign node11964 = (inp[9]) ? 4'b1000 : 4'b1100;
													assign node11968 = (inp[12]) ? 4'b1001 : 4'b1101;
												assign node11971 = (inp[9]) ? node11975 : node11972;
													assign node11972 = (inp[4]) ? 4'b1001 : 4'b1101;
													assign node11975 = (inp[10]) ? 4'b1001 : node11976;
														assign node11976 = (inp[4]) ? 4'b1101 : 4'b1001;
											assign node11980 = (inp[14]) ? node11992 : node11981;
												assign node11981 = (inp[2]) ? node11987 : node11982;
													assign node11982 = (inp[9]) ? 4'b1001 : node11983;
														assign node11983 = (inp[10]) ? 4'b1101 : 4'b1001;
													assign node11987 = (inp[10]) ? 4'b1000 : node11988;
														assign node11988 = (inp[12]) ? 4'b1000 : 4'b1100;
												assign node11992 = (inp[12]) ? node11998 : node11993;
													assign node11993 = (inp[4]) ? 4'b1000 : node11994;
														assign node11994 = (inp[9]) ? 4'b1000 : 4'b1100;
													assign node11998 = (inp[9]) ? 4'b1100 : 4'b1000;
						assign node12001 = (inp[8]) ? node12361 : node12002;
							assign node12002 = (inp[7]) ? node12182 : node12003;
								assign node12003 = (inp[2]) ? node12085 : node12004;
									assign node12004 = (inp[14]) ? node12050 : node12005;
										assign node12005 = (inp[10]) ? node12023 : node12006;
											assign node12006 = (inp[4]) ? node12016 : node12007;
												assign node12007 = (inp[9]) ? node12011 : node12008;
													assign node12008 = (inp[15]) ? 4'b1111 : 4'b1101;
													assign node12011 = (inp[5]) ? node12013 : 4'b1001;
														assign node12013 = (inp[15]) ? 4'b1001 : 4'b1001;
												assign node12016 = (inp[9]) ? 4'b1111 : node12017;
													assign node12017 = (inp[12]) ? node12019 : 4'b1011;
														assign node12019 = (inp[3]) ? 4'b1001 : 4'b1011;
											assign node12023 = (inp[3]) ? node12039 : node12024;
												assign node12024 = (inp[4]) ? node12032 : node12025;
													assign node12025 = (inp[15]) ? node12029 : node12026;
														assign node12026 = (inp[9]) ? 4'b1111 : 4'b1101;
														assign node12029 = (inp[12]) ? 4'b1101 : 4'b1111;
													assign node12032 = (inp[15]) ? node12036 : node12033;
														assign node12033 = (inp[9]) ? 4'b1011 : 4'b1101;
														assign node12036 = (inp[9]) ? 4'b1011 : 4'b1011;
												assign node12039 = (inp[4]) ? node12047 : node12040;
													assign node12040 = (inp[9]) ? node12044 : node12041;
														assign node12041 = (inp[12]) ? 4'b1001 : 4'b1101;
														assign node12044 = (inp[5]) ? 4'b1101 : 4'b1001;
													assign node12047 = (inp[15]) ? 4'b1101 : 4'b1111;
										assign node12050 = (inp[15]) ? node12072 : node12051;
											assign node12051 = (inp[5]) ? node12061 : node12052;
												assign node12052 = (inp[9]) ? node12054 : 4'b1000;
													assign node12054 = (inp[3]) ? node12058 : node12055;
														assign node12055 = (inp[4]) ? 4'b1100 : 4'b1000;
														assign node12058 = (inp[10]) ? 4'b1010 : 4'b1000;
												assign node12061 = (inp[3]) ? node12067 : node12062;
													assign node12062 = (inp[12]) ? node12064 : 4'b1000;
														assign node12064 = (inp[4]) ? 4'b1110 : 4'b1000;
													assign node12067 = (inp[9]) ? node12069 : 4'b1110;
														assign node12069 = (inp[4]) ? 4'b1110 : 4'b1010;
											assign node12072 = (inp[5]) ? node12078 : node12073;
												assign node12073 = (inp[10]) ? node12075 : 4'b1110;
													assign node12075 = (inp[12]) ? 4'b1110 : 4'b1010;
												assign node12078 = (inp[4]) ? 4'b1100 : node12079;
													assign node12079 = (inp[9]) ? node12081 : 4'b1100;
														assign node12081 = (inp[3]) ? 4'b1000 : 4'b1010;
									assign node12085 = (inp[14]) ? node12135 : node12086;
										assign node12086 = (inp[9]) ? node12110 : node12087;
											assign node12087 = (inp[4]) ? node12097 : node12088;
												assign node12088 = (inp[12]) ? node12094 : node12089;
													assign node12089 = (inp[15]) ? 4'b1110 : node12090;
														assign node12090 = (inp[3]) ? 4'b1100 : 4'b1100;
													assign node12094 = (inp[5]) ? 4'b1010 : 4'b1000;
												assign node12097 = (inp[10]) ? node12105 : node12098;
													assign node12098 = (inp[15]) ? node12102 : node12099;
														assign node12099 = (inp[5]) ? 4'b1000 : 4'b1000;
														assign node12102 = (inp[3]) ? 4'b1000 : 4'b1010;
													assign node12105 = (inp[12]) ? node12107 : 4'b1010;
														assign node12107 = (inp[5]) ? 4'b1100 : 4'b1110;
											assign node12110 = (inp[4]) ? node12122 : node12111;
												assign node12111 = (inp[12]) ? node12119 : node12112;
													assign node12112 = (inp[15]) ? node12116 : node12113;
														assign node12113 = (inp[3]) ? 4'b1010 : 4'b1000;
														assign node12116 = (inp[5]) ? 4'b1000 : 4'b1010;
													assign node12119 = (inp[10]) ? 4'b1110 : 4'b1010;
												assign node12122 = (inp[12]) ? node12128 : node12123;
													assign node12123 = (inp[15]) ? node12125 : 4'b1110;
														assign node12125 = (inp[3]) ? 4'b1100 : 4'b1110;
													assign node12128 = (inp[10]) ? node12132 : node12129;
														assign node12129 = (inp[5]) ? 4'b1100 : 4'b1110;
														assign node12132 = (inp[15]) ? 4'b1000 : 4'b1010;
										assign node12135 = (inp[10]) ? node12159 : node12136;
											assign node12136 = (inp[12]) ? node12148 : node12137;
												assign node12137 = (inp[15]) ? node12143 : node12138;
													assign node12138 = (inp[5]) ? 4'b1110 : node12139;
														assign node12139 = (inp[3]) ? 4'b1000 : 4'b1100;
													assign node12143 = (inp[5]) ? 4'b1100 : node12144;
														assign node12144 = (inp[9]) ? 4'b1100 : 4'b1110;
												assign node12148 = (inp[9]) ? node12154 : node12149;
													assign node12149 = (inp[4]) ? 4'b1000 : node12150;
														assign node12150 = (inp[15]) ? 4'b1100 : 4'b1100;
													assign node12154 = (inp[15]) ? node12156 : 4'b1110;
														assign node12156 = (inp[5]) ? 4'b1000 : 4'b1010;
											assign node12159 = (inp[12]) ? node12173 : node12160;
												assign node12160 = (inp[3]) ? node12166 : node12161;
													assign node12161 = (inp[4]) ? node12163 : 4'b1110;
														assign node12163 = (inp[9]) ? 4'b1100 : 4'b1000;
													assign node12166 = (inp[9]) ? node12170 : node12167;
														assign node12167 = (inp[4]) ? 4'b1010 : 4'b1110;
														assign node12170 = (inp[4]) ? 4'b1110 : 4'b1010;
												assign node12173 = (inp[4]) ? node12179 : node12174;
													assign node12174 = (inp[9]) ? 4'b1110 : node12175;
														assign node12175 = (inp[15]) ? 4'b1010 : 4'b1000;
													assign node12179 = (inp[9]) ? 4'b1000 : 4'b1100;
								assign node12182 = (inp[14]) ? node12278 : node12183;
									assign node12183 = (inp[2]) ? node12239 : node12184;
										assign node12184 = (inp[15]) ? node12212 : node12185;
											assign node12185 = (inp[3]) ? node12199 : node12186;
												assign node12186 = (inp[5]) ? node12194 : node12187;
													assign node12187 = (inp[4]) ? node12191 : node12188;
														assign node12188 = (inp[12]) ? 4'b1000 : 4'b1000;
														assign node12191 = (inp[12]) ? 4'b1000 : 4'b1100;
													assign node12194 = (inp[12]) ? 4'b1110 : node12195;
														assign node12195 = (inp[10]) ? 4'b1000 : 4'b1100;
												assign node12199 = (inp[5]) ? node12207 : node12200;
													assign node12200 = (inp[4]) ? node12204 : node12201;
														assign node12201 = (inp[12]) ? 4'b1000 : 4'b1000;
														assign node12204 = (inp[12]) ? 4'b1010 : 4'b1110;
													assign node12207 = (inp[9]) ? node12209 : 4'b1110;
														assign node12209 = (inp[4]) ? 4'b1110 : 4'b1010;
											assign node12212 = (inp[3]) ? node12226 : node12213;
												assign node12213 = (inp[4]) ? node12221 : node12214;
													assign node12214 = (inp[5]) ? node12218 : node12215;
														assign node12215 = (inp[10]) ? 4'b1110 : 4'b1010;
														assign node12218 = (inp[9]) ? 4'b1010 : 4'b1010;
													assign node12221 = (inp[9]) ? node12223 : 4'b1010;
														assign node12223 = (inp[12]) ? 4'b1000 : 4'b1100;
												assign node12226 = (inp[5]) ? node12234 : node12227;
													assign node12227 = (inp[9]) ? node12231 : node12228;
														assign node12228 = (inp[10]) ? 4'b1010 : 4'b1010;
														assign node12231 = (inp[4]) ? 4'b1000 : 4'b1010;
													assign node12234 = (inp[4]) ? node12236 : 4'b1000;
														assign node12236 = (inp[9]) ? 4'b1100 : 4'b1000;
										assign node12239 = (inp[4]) ? node12259 : node12240;
											assign node12240 = (inp[12]) ? node12250 : node12241;
												assign node12241 = (inp[9]) ? node12245 : node12242;
													assign node12242 = (inp[15]) ? 4'b0101 : 4'b0111;
													assign node12245 = (inp[15]) ? 4'b0011 : node12246;
														assign node12246 = (inp[5]) ? 4'b0011 : 4'b0001;
												assign node12250 = (inp[10]) ? node12254 : node12251;
													assign node12251 = (inp[9]) ? 4'b0011 : 4'b0111;
													assign node12254 = (inp[15]) ? node12256 : 4'b0111;
														assign node12256 = (inp[3]) ? 4'b0101 : 4'b0111;
											assign node12259 = (inp[9]) ? node12273 : node12260;
												assign node12260 = (inp[5]) ? node12266 : node12261;
													assign node12261 = (inp[15]) ? node12263 : 4'b0001;
														assign node12263 = (inp[3]) ? 4'b0011 : 4'b0011;
													assign node12266 = (inp[10]) ? node12270 : node12267;
														assign node12267 = (inp[12]) ? 4'b0001 : 4'b0001;
														assign node12270 = (inp[12]) ? 4'b0101 : 4'b0001;
												assign node12273 = (inp[10]) ? node12275 : 4'b0101;
													assign node12275 = (inp[12]) ? 4'b0001 : 4'b0101;
									assign node12278 = (inp[10]) ? node12320 : node12279;
										assign node12279 = (inp[15]) ? node12297 : node12280;
											assign node12280 = (inp[12]) ? node12288 : node12281;
												assign node12281 = (inp[3]) ? node12283 : 4'b0001;
													assign node12283 = (inp[9]) ? node12285 : 4'b0001;
														assign node12285 = (inp[4]) ? 4'b0111 : 4'b0011;
												assign node12288 = (inp[5]) ? node12290 : 4'b0101;
													assign node12290 = (inp[3]) ? node12294 : node12291;
														assign node12291 = (inp[4]) ? 4'b0111 : 4'b0101;
														assign node12294 = (inp[9]) ? 4'b0011 : 4'b0011;
											assign node12297 = (inp[5]) ? node12311 : node12298;
												assign node12298 = (inp[2]) ? node12304 : node12299;
													assign node12299 = (inp[12]) ? node12301 : 4'b0011;
														assign node12301 = (inp[9]) ? 4'b0011 : 4'b0111;
													assign node12304 = (inp[9]) ? node12308 : node12305;
														assign node12305 = (inp[4]) ? 4'b0011 : 4'b0111;
														assign node12308 = (inp[4]) ? 4'b0111 : 4'b0011;
												assign node12311 = (inp[9]) ? node12315 : node12312;
													assign node12312 = (inp[4]) ? 4'b0011 : 4'b0111;
													assign node12315 = (inp[4]) ? 4'b0101 : node12316;
														assign node12316 = (inp[12]) ? 4'b0001 : 4'b0011;
										assign node12320 = (inp[12]) ? node12340 : node12321;
											assign node12321 = (inp[15]) ? node12329 : node12322;
												assign node12322 = (inp[4]) ? node12324 : 4'b0101;
													assign node12324 = (inp[2]) ? node12326 : 4'b0001;
														assign node12326 = (inp[3]) ? 4'b0111 : 4'b0101;
												assign node12329 = (inp[4]) ? node12333 : node12330;
													assign node12330 = (inp[9]) ? 4'b0011 : 4'b0111;
													assign node12333 = (inp[9]) ? node12337 : node12334;
														assign node12334 = (inp[3]) ? 4'b0001 : 4'b0011;
														assign node12337 = (inp[3]) ? 4'b0101 : 4'b0111;
											assign node12340 = (inp[15]) ? node12352 : node12341;
												assign node12341 = (inp[5]) ? node12347 : node12342;
													assign node12342 = (inp[4]) ? node12344 : 4'b0001;
														assign node12344 = (inp[9]) ? 4'b0001 : 4'b0101;
													assign node12347 = (inp[3]) ? 4'b0011 : node12348;
														assign node12348 = (inp[2]) ? 4'b0111 : 4'b0011;
												assign node12352 = (inp[9]) ? node12358 : node12353;
													assign node12353 = (inp[4]) ? node12355 : 4'b0011;
														assign node12355 = (inp[3]) ? 4'b0101 : 4'b0111;
													assign node12358 = (inp[4]) ? 4'b0001 : 4'b0101;
							assign node12361 = (inp[7]) ? node12521 : node12362;
								assign node12362 = (inp[14]) ? node12450 : node12363;
									assign node12363 = (inp[2]) ? node12403 : node12364;
										assign node12364 = (inp[3]) ? node12384 : node12365;
											assign node12365 = (inp[15]) ? node12377 : node12366;
												assign node12366 = (inp[9]) ? node12372 : node12367;
													assign node12367 = (inp[5]) ? 4'b1000 : node12368;
														assign node12368 = (inp[10]) ? 4'b1000 : 4'b1100;
													assign node12372 = (inp[5]) ? 4'b1110 : node12373;
														assign node12373 = (inp[10]) ? 4'b1000 : 4'b1000;
												assign node12377 = (inp[12]) ? 4'b1110 : node12378;
													assign node12378 = (inp[9]) ? node12380 : 4'b1010;
														assign node12380 = (inp[4]) ? 4'b1110 : 4'b1010;
											assign node12384 = (inp[15]) ? node12394 : node12385;
												assign node12385 = (inp[12]) ? node12389 : node12386;
													assign node12386 = (inp[9]) ? 4'b1110 : 4'b1100;
													assign node12389 = (inp[9]) ? 4'b1010 : node12390;
														assign node12390 = (inp[4]) ? 4'b1110 : 4'b1010;
												assign node12394 = (inp[9]) ? node12396 : 4'b1100;
													assign node12396 = (inp[5]) ? node12400 : node12397;
														assign node12397 = (inp[12]) ? 4'b1000 : 4'b1100;
														assign node12400 = (inp[12]) ? 4'b1000 : 4'b1000;
										assign node12403 = (inp[3]) ? node12427 : node12404;
											assign node12404 = (inp[15]) ? node12414 : node12405;
												assign node12405 = (inp[5]) ? node12407 : 4'b0001;
													assign node12407 = (inp[4]) ? node12411 : node12408;
														assign node12408 = (inp[10]) ? 4'b0001 : 4'b0101;
														assign node12411 = (inp[10]) ? 4'b0011 : 4'b0111;
												assign node12414 = (inp[4]) ? node12420 : node12415;
													assign node12415 = (inp[9]) ? 4'b0011 : node12416;
														assign node12416 = (inp[12]) ? 4'b0011 : 4'b0111;
													assign node12420 = (inp[5]) ? node12424 : node12421;
														assign node12421 = (inp[9]) ? 4'b0011 : 4'b0111;
														assign node12424 = (inp[10]) ? 4'b0001 : 4'b0101;
											assign node12427 = (inp[15]) ? node12439 : node12428;
												assign node12428 = (inp[4]) ? node12434 : node12429;
													assign node12429 = (inp[10]) ? 4'b0111 : node12430;
														assign node12430 = (inp[5]) ? 4'b0011 : 4'b0001;
													assign node12434 = (inp[12]) ? node12436 : 4'b0111;
														assign node12436 = (inp[9]) ? 4'b0011 : 4'b0111;
												assign node12439 = (inp[5]) ? node12445 : node12440;
													assign node12440 = (inp[9]) ? 4'b0101 : node12441;
														assign node12441 = (inp[12]) ? 4'b0101 : 4'b0011;
													assign node12445 = (inp[12]) ? node12447 : 4'b0101;
														assign node12447 = (inp[10]) ? 4'b0001 : 4'b0001;
									assign node12450 = (inp[15]) ? node12484 : node12451;
										assign node12451 = (inp[3]) ? node12467 : node12452;
											assign node12452 = (inp[4]) ? node12462 : node12453;
												assign node12453 = (inp[12]) ? node12457 : node12454;
													assign node12454 = (inp[9]) ? 4'b0001 : 4'b0101;
													assign node12457 = (inp[5]) ? 4'b0001 : node12458;
														assign node12458 = (inp[9]) ? 4'b0101 : 4'b0001;
												assign node12462 = (inp[9]) ? node12464 : 4'b0001;
													assign node12464 = (inp[12]) ? 4'b0011 : 4'b0111;
											assign node12467 = (inp[12]) ? node12479 : node12468;
												assign node12468 = (inp[5]) ? node12474 : node12469;
													assign node12469 = (inp[9]) ? 4'b0001 : node12470;
														assign node12470 = (inp[4]) ? 4'b0001 : 4'b0101;
													assign node12474 = (inp[9]) ? 4'b0011 : node12475;
														assign node12475 = (inp[4]) ? 4'b0011 : 4'b0111;
												assign node12479 = (inp[4]) ? node12481 : 4'b0111;
													assign node12481 = (inp[10]) ? 4'b0011 : 4'b0111;
										assign node12484 = (inp[5]) ? node12502 : node12485;
											assign node12485 = (inp[4]) ? node12493 : node12486;
												assign node12486 = (inp[9]) ? node12488 : 4'b0111;
													assign node12488 = (inp[12]) ? node12490 : 4'b0011;
														assign node12490 = (inp[10]) ? 4'b0111 : 4'b0011;
												assign node12493 = (inp[9]) ? node12499 : node12494;
													assign node12494 = (inp[12]) ? node12496 : 4'b0011;
														assign node12496 = (inp[10]) ? 4'b0101 : 4'b0011;
													assign node12499 = (inp[2]) ? 4'b0101 : 4'b0111;
											assign node12502 = (inp[3]) ? node12514 : node12503;
												assign node12503 = (inp[9]) ? node12509 : node12504;
													assign node12504 = (inp[4]) ? 4'b0011 : node12505;
														assign node12505 = (inp[10]) ? 4'b0011 : 4'b0111;
													assign node12509 = (inp[4]) ? 4'b0101 : node12510;
														assign node12510 = (inp[2]) ? 4'b0011 : 4'b0001;
												assign node12514 = (inp[10]) ? node12516 : 4'b0101;
													assign node12516 = (inp[2]) ? 4'b0101 : node12517;
														assign node12517 = (inp[4]) ? 4'b0101 : 4'b0001;
								assign node12521 = (inp[2]) ? node12609 : node12522;
									assign node12522 = (inp[14]) ? node12570 : node12523;
										assign node12523 = (inp[10]) ? node12547 : node12524;
											assign node12524 = (inp[15]) ? node12536 : node12525;
												assign node12525 = (inp[3]) ? node12533 : node12526;
													assign node12526 = (inp[4]) ? node12530 : node12527;
														assign node12527 = (inp[9]) ? 4'b0001 : 4'b0101;
														assign node12530 = (inp[9]) ? 4'b0101 : 4'b0001;
													assign node12533 = (inp[12]) ? 4'b0111 : 4'b0011;
												assign node12536 = (inp[5]) ? node12542 : node12537;
													assign node12537 = (inp[4]) ? 4'b0011 : node12538;
														assign node12538 = (inp[9]) ? 4'b0011 : 4'b0111;
													assign node12542 = (inp[3]) ? node12544 : 4'b0111;
														assign node12544 = (inp[12]) ? 4'b0001 : 4'b0001;
											assign node12547 = (inp[15]) ? node12561 : node12548;
												assign node12548 = (inp[5]) ? node12556 : node12549;
													assign node12549 = (inp[3]) ? node12553 : node12550;
														assign node12550 = (inp[9]) ? 4'b0001 : 4'b0001;
														assign node12553 = (inp[9]) ? 4'b0111 : 4'b0001;
													assign node12556 = (inp[3]) ? node12558 : 4'b0111;
														assign node12558 = (inp[9]) ? 4'b0011 : 4'b0111;
												assign node12561 = (inp[5]) ? node12565 : node12562;
													assign node12562 = (inp[12]) ? 4'b0101 : 4'b0011;
													assign node12565 = (inp[4]) ? 4'b0101 : node12566;
														assign node12566 = (inp[12]) ? 4'b0001 : 4'b0001;
										assign node12570 = (inp[12]) ? node12590 : node12571;
											assign node12571 = (inp[9]) ? node12579 : node12572;
												assign node12572 = (inp[4]) ? 4'b0010 : node12573;
													assign node12573 = (inp[10]) ? node12575 : 4'b0110;
														assign node12575 = (inp[5]) ? 4'b0100 : 4'b0110;
												assign node12579 = (inp[4]) ? node12583 : node12580;
													assign node12580 = (inp[15]) ? 4'b0010 : 4'b0000;
													assign node12583 = (inp[10]) ? node12587 : node12584;
														assign node12584 = (inp[15]) ? 4'b0100 : 4'b0110;
														assign node12587 = (inp[5]) ? 4'b0100 : 4'b0100;
											assign node12590 = (inp[4]) ? node12600 : node12591;
												assign node12591 = (inp[9]) ? node12595 : node12592;
													assign node12592 = (inp[10]) ? 4'b0010 : 4'b0110;
													assign node12595 = (inp[5]) ? node12597 : 4'b0000;
														assign node12597 = (inp[15]) ? 4'b0000 : 4'b0010;
												assign node12600 = (inp[5]) ? 4'b0110 : node12601;
													assign node12601 = (inp[15]) ? node12605 : node12602;
														assign node12602 = (inp[10]) ? 4'b0010 : 4'b0000;
														assign node12605 = (inp[9]) ? 4'b0100 : 4'b0000;
									assign node12609 = (inp[3]) ? node12651 : node12610;
										assign node12610 = (inp[15]) ? node12634 : node12611;
											assign node12611 = (inp[5]) ? node12623 : node12612;
												assign node12612 = (inp[14]) ? node12618 : node12613;
													assign node12613 = (inp[9]) ? 4'b0100 : node12614;
														assign node12614 = (inp[4]) ? 4'b0000 : 4'b0100;
													assign node12618 = (inp[4]) ? node12620 : 4'b0000;
														assign node12620 = (inp[12]) ? 4'b0000 : 4'b0000;
												assign node12623 = (inp[10]) ? node12629 : node12624;
													assign node12624 = (inp[14]) ? node12626 : 4'b0000;
														assign node12626 = (inp[9]) ? 4'b0000 : 4'b0100;
													assign node12629 = (inp[4]) ? node12631 : 4'b0000;
														assign node12631 = (inp[14]) ? 4'b0110 : 4'b0010;
											assign node12634 = (inp[5]) ? node12642 : node12635;
												assign node12635 = (inp[4]) ? node12639 : node12636;
													assign node12636 = (inp[9]) ? 4'b0010 : 4'b0110;
													assign node12639 = (inp[9]) ? 4'b0110 : 4'b0010;
												assign node12642 = (inp[9]) ? node12646 : node12643;
													assign node12643 = (inp[4]) ? 4'b0010 : 4'b0110;
													assign node12646 = (inp[10]) ? node12648 : 4'b0100;
														assign node12648 = (inp[12]) ? 4'b0100 : 4'b0010;
										assign node12651 = (inp[15]) ? node12677 : node12652;
											assign node12652 = (inp[5]) ? node12664 : node12653;
												assign node12653 = (inp[4]) ? node12659 : node12654;
													assign node12654 = (inp[14]) ? 4'b0000 : node12655;
														assign node12655 = (inp[10]) ? 4'b0100 : 4'b0000;
													assign node12659 = (inp[9]) ? node12661 : 4'b0000;
														assign node12661 = (inp[10]) ? 4'b0010 : 4'b0110;
												assign node12664 = (inp[9]) ? node12672 : node12665;
													assign node12665 = (inp[4]) ? node12669 : node12666;
														assign node12666 = (inp[12]) ? 4'b0010 : 4'b0110;
														assign node12669 = (inp[12]) ? 4'b0010 : 4'b0010;
													assign node12672 = (inp[4]) ? node12674 : 4'b0010;
														assign node12674 = (inp[10]) ? 4'b0010 : 4'b0110;
											assign node12677 = (inp[5]) ? node12685 : node12678;
												assign node12678 = (inp[14]) ? 4'b0010 : node12679;
													assign node12679 = (inp[9]) ? 4'b0100 : node12680;
														assign node12680 = (inp[12]) ? 4'b0110 : 4'b0010;
												assign node12685 = (inp[12]) ? 4'b0000 : node12686;
													assign node12686 = (inp[4]) ? node12688 : 4'b0100;
														assign node12688 = (inp[9]) ? 4'b0100 : 4'b0000;
					assign node12692 = (inp[1]) ? node13390 : node12693;
						assign node12693 = (inp[7]) ? node13037 : node12694;
							assign node12694 = (inp[8]) ? node12868 : node12695;
								assign node12695 = (inp[2]) ? node12793 : node12696;
									assign node12696 = (inp[14]) ? node12752 : node12697;
										assign node12697 = (inp[10]) ? node12725 : node12698;
											assign node12698 = (inp[5]) ? node12712 : node12699;
												assign node12699 = (inp[15]) ? node12707 : node12700;
													assign node12700 = (inp[9]) ? node12704 : node12701;
														assign node12701 = (inp[4]) ? 4'b1001 : 4'b1101;
														assign node12704 = (inp[12]) ? 4'b1111 : 4'b1001;
													assign node12707 = (inp[3]) ? node12709 : 4'b1111;
														assign node12709 = (inp[4]) ? 4'b1011 : 4'b1111;
												assign node12712 = (inp[12]) ? node12720 : node12713;
													assign node12713 = (inp[4]) ? node12717 : node12714;
														assign node12714 = (inp[15]) ? 4'b1001 : 4'b1111;
														assign node12717 = (inp[9]) ? 4'b1101 : 4'b1001;
													assign node12720 = (inp[15]) ? 4'b1011 : node12721;
														assign node12721 = (inp[3]) ? 4'b1111 : 4'b1101;
											assign node12725 = (inp[12]) ? node12739 : node12726;
												assign node12726 = (inp[15]) ? node12734 : node12727;
													assign node12727 = (inp[9]) ? node12731 : node12728;
														assign node12728 = (inp[4]) ? 4'b1001 : 4'b1101;
														assign node12731 = (inp[3]) ? 4'b1001 : 4'b1001;
													assign node12734 = (inp[9]) ? 4'b1101 : node12735;
														assign node12735 = (inp[5]) ? 4'b1001 : 4'b1011;
												assign node12739 = (inp[15]) ? node12747 : node12740;
													assign node12740 = (inp[3]) ? node12744 : node12741;
														assign node12741 = (inp[4]) ? 4'b1101 : 4'b1001;
														assign node12744 = (inp[9]) ? 4'b1111 : 4'b1011;
													assign node12747 = (inp[5]) ? node12749 : 4'b1111;
														assign node12749 = (inp[3]) ? 4'b1001 : 4'b1101;
										assign node12752 = (inp[4]) ? node12776 : node12753;
											assign node12753 = (inp[9]) ? node12767 : node12754;
												assign node12754 = (inp[15]) ? node12762 : node12755;
													assign node12755 = (inp[5]) ? node12759 : node12756;
														assign node12756 = (inp[10]) ? 4'b1000 : 4'b1100;
														assign node12759 = (inp[12]) ? 4'b1010 : 4'b1110;
													assign node12762 = (inp[12]) ? node12764 : 4'b1110;
														assign node12764 = (inp[10]) ? 4'b1010 : 4'b1110;
												assign node12767 = (inp[12]) ? node12773 : node12768;
													assign node12768 = (inp[5]) ? node12770 : 4'b1010;
														assign node12770 = (inp[3]) ? 4'b1010 : 4'b1000;
													assign node12773 = (inp[15]) ? 4'b1010 : 4'b1110;
											assign node12776 = (inp[15]) ? node12784 : node12777;
												assign node12777 = (inp[9]) ? node12781 : node12778;
													assign node12778 = (inp[12]) ? 4'b1110 : 4'b1000;
													assign node12781 = (inp[12]) ? 4'b1010 : 4'b1110;
												assign node12784 = (inp[3]) ? node12788 : node12785;
													assign node12785 = (inp[10]) ? 4'b1110 : 4'b1100;
													assign node12788 = (inp[10]) ? node12790 : 4'b1100;
														assign node12790 = (inp[5]) ? 4'b1000 : 4'b1100;
									assign node12793 = (inp[15]) ? node12837 : node12794;
										assign node12794 = (inp[5]) ? node12820 : node12795;
											assign node12795 = (inp[3]) ? node12807 : node12796;
												assign node12796 = (inp[14]) ? node12802 : node12797;
													assign node12797 = (inp[9]) ? node12799 : 4'b1000;
														assign node12799 = (inp[12]) ? 4'b1000 : 4'b1000;
													assign node12802 = (inp[12]) ? node12804 : 4'b1100;
														assign node12804 = (inp[10]) ? 4'b1000 : 4'b1100;
												assign node12807 = (inp[12]) ? node12815 : node12808;
													assign node12808 = (inp[4]) ? node12812 : node12809;
														assign node12809 = (inp[9]) ? 4'b1000 : 4'b1100;
														assign node12812 = (inp[14]) ? 4'b1000 : 4'b1110;
													assign node12815 = (inp[10]) ? node12817 : 4'b1000;
														assign node12817 = (inp[4]) ? 4'b1010 : 4'b1110;
											assign node12820 = (inp[4]) ? node12832 : node12821;
												assign node12821 = (inp[3]) ? node12827 : node12822;
													assign node12822 = (inp[9]) ? 4'b1000 : node12823;
														assign node12823 = (inp[10]) ? 4'b1000 : 4'b1100;
													assign node12827 = (inp[9]) ? 4'b1010 : node12828;
														assign node12828 = (inp[10]) ? 4'b1010 : 4'b1110;
												assign node12832 = (inp[10]) ? node12834 : 4'b1110;
													assign node12834 = (inp[9]) ? 4'b1010 : 4'b1110;
										assign node12837 = (inp[3]) ? node12855 : node12838;
											assign node12838 = (inp[9]) ? node12846 : node12839;
												assign node12839 = (inp[10]) ? node12841 : 4'b1110;
													assign node12841 = (inp[5]) ? node12843 : 4'b1110;
														assign node12843 = (inp[14]) ? 4'b1010 : 4'b1110;
												assign node12846 = (inp[10]) ? node12848 : 4'b1010;
													assign node12848 = (inp[5]) ? node12852 : node12849;
														assign node12849 = (inp[14]) ? 4'b1010 : 4'b1110;
														assign node12852 = (inp[4]) ? 4'b1000 : 4'b1000;
											assign node12855 = (inp[5]) ? node12863 : node12856;
												assign node12856 = (inp[9]) ? node12860 : node12857;
													assign node12857 = (inp[4]) ? 4'b1010 : 4'b1110;
													assign node12860 = (inp[4]) ? 4'b1100 : 4'b1010;
												assign node12863 = (inp[4]) ? 4'b1000 : node12864;
													assign node12864 = (inp[9]) ? 4'b1000 : 4'b1100;
								assign node12868 = (inp[2]) ? node12956 : node12869;
									assign node12869 = (inp[14]) ? node12911 : node12870;
										assign node12870 = (inp[9]) ? node12890 : node12871;
											assign node12871 = (inp[4]) ? node12881 : node12872;
												assign node12872 = (inp[10]) ? node12878 : node12873;
													assign node12873 = (inp[15]) ? 4'b1110 : node12874;
														assign node12874 = (inp[5]) ? 4'b1110 : 4'b1100;
													assign node12878 = (inp[12]) ? 4'b1010 : 4'b1110;
												assign node12881 = (inp[3]) ? node12885 : node12882;
													assign node12882 = (inp[15]) ? 4'b1010 : 4'b1000;
													assign node12885 = (inp[10]) ? node12887 : 4'b1010;
														assign node12887 = (inp[12]) ? 4'b1100 : 4'b1000;
											assign node12890 = (inp[4]) ? node12904 : node12891;
												assign node12891 = (inp[10]) ? node12897 : node12892;
													assign node12892 = (inp[5]) ? node12894 : 4'b1000;
														assign node12894 = (inp[3]) ? 4'b1010 : 4'b1000;
													assign node12897 = (inp[12]) ? node12901 : node12898;
														assign node12898 = (inp[3]) ? 4'b1000 : 4'b1010;
														assign node12901 = (inp[5]) ? 4'b1100 : 4'b1110;
												assign node12904 = (inp[10]) ? node12906 : 4'b1100;
													assign node12906 = (inp[12]) ? node12908 : 4'b1100;
														assign node12908 = (inp[15]) ? 4'b1000 : 4'b1010;
										assign node12911 = (inp[5]) ? node12935 : node12912;
											assign node12912 = (inp[15]) ? node12924 : node12913;
												assign node12913 = (inp[9]) ? node12919 : node12914;
													assign node12914 = (inp[4]) ? node12916 : 4'b0101;
														assign node12916 = (inp[10]) ? 4'b0001 : 4'b0001;
													assign node12919 = (inp[4]) ? node12921 : 4'b0001;
														assign node12921 = (inp[12]) ? 4'b0011 : 4'b0111;
												assign node12924 = (inp[12]) ? node12930 : node12925;
													assign node12925 = (inp[10]) ? node12927 : 4'b0011;
														assign node12927 = (inp[9]) ? 4'b0011 : 4'b0111;
													assign node12930 = (inp[3]) ? node12932 : 4'b0011;
														assign node12932 = (inp[10]) ? 4'b0101 : 4'b0111;
											assign node12935 = (inp[15]) ? node12945 : node12936;
												assign node12936 = (inp[3]) ? node12940 : node12937;
													assign node12937 = (inp[10]) ? 4'b0111 : 4'b0001;
													assign node12940 = (inp[10]) ? 4'b0111 : node12941;
														assign node12941 = (inp[4]) ? 4'b0111 : 4'b0011;
												assign node12945 = (inp[3]) ? node12953 : node12946;
													assign node12946 = (inp[10]) ? node12950 : node12947;
														assign node12947 = (inp[4]) ? 4'b0011 : 4'b0111;
														assign node12950 = (inp[12]) ? 4'b0101 : 4'b0111;
													assign node12953 = (inp[9]) ? 4'b0001 : 4'b0101;
									assign node12956 = (inp[4]) ? node12998 : node12957;
										assign node12957 = (inp[9]) ? node12981 : node12958;
											assign node12958 = (inp[10]) ? node12968 : node12959;
												assign node12959 = (inp[15]) ? node12965 : node12960;
													assign node12960 = (inp[14]) ? node12962 : 4'b0101;
														assign node12962 = (inp[5]) ? 4'b0111 : 4'b0101;
													assign node12965 = (inp[5]) ? 4'b0101 : 4'b0111;
												assign node12968 = (inp[12]) ? node12974 : node12969;
													assign node12969 = (inp[5]) ? 4'b0101 : node12970;
														assign node12970 = (inp[15]) ? 4'b0111 : 4'b0101;
													assign node12974 = (inp[3]) ? node12978 : node12975;
														assign node12975 = (inp[5]) ? 4'b0001 : 4'b0011;
														assign node12978 = (inp[15]) ? 4'b0001 : 4'b0011;
											assign node12981 = (inp[12]) ? node12989 : node12982;
												assign node12982 = (inp[15]) ? node12986 : node12983;
													assign node12983 = (inp[3]) ? 4'b0011 : 4'b0001;
													assign node12986 = (inp[3]) ? 4'b0001 : 4'b0011;
												assign node12989 = (inp[10]) ? node12993 : node12990;
													assign node12990 = (inp[14]) ? 4'b0011 : 4'b0001;
													assign node12993 = (inp[15]) ? node12995 : 4'b0111;
														assign node12995 = (inp[3]) ? 4'b0101 : 4'b0111;
										assign node12998 = (inp[9]) ? node13022 : node12999;
											assign node12999 = (inp[10]) ? node13011 : node13000;
												assign node13000 = (inp[15]) ? node13006 : node13001;
													assign node13001 = (inp[3]) ? node13003 : 4'b0001;
														assign node13003 = (inp[14]) ? 4'b0011 : 4'b0001;
													assign node13006 = (inp[14]) ? node13008 : 4'b0011;
														assign node13008 = (inp[12]) ? 4'b0001 : 4'b0011;
												assign node13011 = (inp[12]) ? node13015 : node13012;
													assign node13012 = (inp[15]) ? 4'b0011 : 4'b0001;
													assign node13015 = (inp[14]) ? node13019 : node13016;
														assign node13016 = (inp[15]) ? 4'b0101 : 4'b0111;
														assign node13019 = (inp[5]) ? 4'b0101 : 4'b0101;
											assign node13022 = (inp[15]) ? node13032 : node13023;
												assign node13023 = (inp[5]) ? 4'b0111 : node13024;
													assign node13024 = (inp[10]) ? node13028 : node13025;
														assign node13025 = (inp[14]) ? 4'b0101 : 4'b0111;
														assign node13028 = (inp[3]) ? 4'b0011 : 4'b0001;
												assign node13032 = (inp[12]) ? node13034 : 4'b0101;
													assign node13034 = (inp[10]) ? 4'b0001 : 4'b0111;
							assign node13037 = (inp[8]) ? node13223 : node13038;
								assign node13038 = (inp[2]) ? node13132 : node13039;
									assign node13039 = (inp[14]) ? node13089 : node13040;
										assign node13040 = (inp[15]) ? node13060 : node13041;
											assign node13041 = (inp[5]) ? node13053 : node13042;
												assign node13042 = (inp[9]) ? node13048 : node13043;
													assign node13043 = (inp[3]) ? node13045 : 4'b1000;
														assign node13045 = (inp[4]) ? 4'b1000 : 4'b1100;
													assign node13048 = (inp[4]) ? node13050 : 4'b1000;
														assign node13050 = (inp[3]) ? 4'b1110 : 4'b1100;
												assign node13053 = (inp[4]) ? node13057 : node13054;
													assign node13054 = (inp[3]) ? 4'b1010 : 4'b1000;
													assign node13057 = (inp[10]) ? 4'b1010 : 4'b1110;
											assign node13060 = (inp[3]) ? node13074 : node13061;
												assign node13061 = (inp[12]) ? node13069 : node13062;
													assign node13062 = (inp[5]) ? node13066 : node13063;
														assign node13063 = (inp[10]) ? 4'b1110 : 4'b1010;
														assign node13066 = (inp[9]) ? 4'b1100 : 4'b1110;
													assign node13069 = (inp[10]) ? 4'b1010 : node13070;
														assign node13070 = (inp[9]) ? 4'b1010 : 4'b1110;
												assign node13074 = (inp[5]) ? node13082 : node13075;
													assign node13075 = (inp[9]) ? node13079 : node13076;
														assign node13076 = (inp[10]) ? 4'b1010 : 4'b1010;
														assign node13079 = (inp[10]) ? 4'b1100 : 4'b1000;
													assign node13082 = (inp[10]) ? node13086 : node13083;
														assign node13083 = (inp[4]) ? 4'b1000 : 4'b1100;
														assign node13086 = (inp[4]) ? 4'b1100 : 4'b1000;
										assign node13089 = (inp[9]) ? node13109 : node13090;
											assign node13090 = (inp[4]) ? node13098 : node13091;
												assign node13091 = (inp[15]) ? node13093 : 4'b0101;
													assign node13093 = (inp[3]) ? node13095 : 4'b0111;
														assign node13095 = (inp[10]) ? 4'b0001 : 4'b0101;
												assign node13098 = (inp[12]) ? node13102 : node13099;
													assign node13099 = (inp[5]) ? 4'b0011 : 4'b0001;
													assign node13102 = (inp[10]) ? node13106 : node13103;
														assign node13103 = (inp[15]) ? 4'b0011 : 4'b0001;
														assign node13106 = (inp[15]) ? 4'b0101 : 4'b0111;
											assign node13109 = (inp[4]) ? node13121 : node13110;
												assign node13110 = (inp[12]) ? node13116 : node13111;
													assign node13111 = (inp[15]) ? node13113 : 4'b0001;
														assign node13113 = (inp[3]) ? 4'b0001 : 4'b0011;
													assign node13116 = (inp[10]) ? 4'b0101 : node13117;
														assign node13117 = (inp[5]) ? 4'b0001 : 4'b0001;
												assign node13121 = (inp[12]) ? node13127 : node13122;
													assign node13122 = (inp[15]) ? 4'b0101 : node13123;
														assign node13123 = (inp[10]) ? 4'b0111 : 4'b0101;
													assign node13127 = (inp[10]) ? node13129 : 4'b0101;
														assign node13129 = (inp[15]) ? 4'b0001 : 4'b0011;
									assign node13132 = (inp[10]) ? node13174 : node13133;
										assign node13133 = (inp[15]) ? node13155 : node13134;
											assign node13134 = (inp[3]) ? node13144 : node13135;
												assign node13135 = (inp[4]) ? node13139 : node13136;
													assign node13136 = (inp[9]) ? 4'b0001 : 4'b0101;
													assign node13139 = (inp[9]) ? node13141 : 4'b0001;
														assign node13141 = (inp[12]) ? 4'b0111 : 4'b0101;
												assign node13144 = (inp[5]) ? node13150 : node13145;
													assign node13145 = (inp[9]) ? 4'b0111 : node13146;
														assign node13146 = (inp[12]) ? 4'b0101 : 4'b0001;
													assign node13150 = (inp[12]) ? node13152 : 4'b0111;
														assign node13152 = (inp[14]) ? 4'b0011 : 4'b0011;
											assign node13155 = (inp[3]) ? node13167 : node13156;
												assign node13156 = (inp[14]) ? node13162 : node13157;
													assign node13157 = (inp[9]) ? node13159 : 4'b0011;
														assign node13159 = (inp[4]) ? 4'b0101 : 4'b0011;
													assign node13162 = (inp[12]) ? 4'b0111 : node13163;
														assign node13163 = (inp[9]) ? 4'b0011 : 4'b0011;
												assign node13167 = (inp[5]) ? 4'b0001 : node13168;
													assign node13168 = (inp[9]) ? 4'b0101 : node13169;
														assign node13169 = (inp[4]) ? 4'b0011 : 4'b0111;
										assign node13174 = (inp[14]) ? node13196 : node13175;
											assign node13175 = (inp[15]) ? node13187 : node13176;
												assign node13176 = (inp[4]) ? node13182 : node13177;
													assign node13177 = (inp[12]) ? 4'b0001 : node13178;
														assign node13178 = (inp[9]) ? 4'b0001 : 4'b0101;
													assign node13182 = (inp[3]) ? node13184 : 4'b0001;
														assign node13184 = (inp[5]) ? 4'b0011 : 4'b0001;
												assign node13187 = (inp[5]) ? node13191 : node13188;
													assign node13188 = (inp[12]) ? 4'b0101 : 4'b0011;
													assign node13191 = (inp[3]) ? 4'b0001 : node13192;
														assign node13192 = (inp[4]) ? 4'b0001 : 4'b0011;
											assign node13196 = (inp[12]) ? node13212 : node13197;
												assign node13197 = (inp[5]) ? node13205 : node13198;
													assign node13198 = (inp[15]) ? node13202 : node13199;
														assign node13199 = (inp[9]) ? 4'b0001 : 4'b0101;
														assign node13202 = (inp[3]) ? 4'b0101 : 4'b0111;
													assign node13205 = (inp[3]) ? node13209 : node13206;
														assign node13206 = (inp[15]) ? 4'b0011 : 4'b0001;
														assign node13209 = (inp[15]) ? 4'b0001 : 4'b0111;
												assign node13212 = (inp[9]) ? node13218 : node13213;
													assign node13213 = (inp[4]) ? 4'b0101 : node13214;
														assign node13214 = (inp[15]) ? 4'b0001 : 4'b0001;
													assign node13218 = (inp[4]) ? node13220 : 4'b0111;
														assign node13220 = (inp[3]) ? 4'b0001 : 4'b0011;
								assign node13223 = (inp[14]) ? node13303 : node13224;
									assign node13224 = (inp[2]) ? node13260 : node13225;
										assign node13225 = (inp[10]) ? node13237 : node13226;
											assign node13226 = (inp[4]) ? node13234 : node13227;
												assign node13227 = (inp[9]) ? node13231 : node13228;
													assign node13228 = (inp[12]) ? 4'b0111 : 4'b0101;
													assign node13231 = (inp[5]) ? 4'b0001 : 4'b0011;
												assign node13234 = (inp[9]) ? 4'b0111 : 4'b0011;
											assign node13237 = (inp[9]) ? node13249 : node13238;
												assign node13238 = (inp[4]) ? node13244 : node13239;
													assign node13239 = (inp[12]) ? 4'b0011 : node13240;
														assign node13240 = (inp[5]) ? 4'b0101 : 4'b0111;
													assign node13244 = (inp[12]) ? node13246 : 4'b0001;
														assign node13246 = (inp[5]) ? 4'b0101 : 4'b0101;
												assign node13249 = (inp[12]) ? node13255 : node13250;
													assign node13250 = (inp[3]) ? node13252 : 4'b0011;
														assign node13252 = (inp[15]) ? 4'b0001 : 4'b0001;
													assign node13255 = (inp[4]) ? 4'b0001 : node13256;
														assign node13256 = (inp[3]) ? 4'b0111 : 4'b0101;
										assign node13260 = (inp[12]) ? node13280 : node13261;
											assign node13261 = (inp[4]) ? node13271 : node13262;
												assign node13262 = (inp[15]) ? node13266 : node13263;
													assign node13263 = (inp[9]) ? 4'b0000 : 4'b0100;
													assign node13266 = (inp[3]) ? node13268 : 4'b0010;
														assign node13268 = (inp[5]) ? 4'b0000 : 4'b0010;
												assign node13271 = (inp[9]) ? node13275 : node13272;
													assign node13272 = (inp[10]) ? 4'b0010 : 4'b0000;
													assign node13275 = (inp[3]) ? node13277 : 4'b0110;
														assign node13277 = (inp[10]) ? 4'b0110 : 4'b0100;
											assign node13280 = (inp[5]) ? node13292 : node13281;
												assign node13281 = (inp[10]) ? node13289 : node13282;
													assign node13282 = (inp[15]) ? node13286 : node13283;
														assign node13283 = (inp[3]) ? 4'b0100 : 4'b0000;
														assign node13286 = (inp[9]) ? 4'b0010 : 4'b0110;
													assign node13289 = (inp[4]) ? 4'b0000 : 4'b0100;
												assign node13292 = (inp[15]) ? node13298 : node13293;
													assign node13293 = (inp[10]) ? 4'b0110 : node13294;
														assign node13294 = (inp[9]) ? 4'b0110 : 4'b0000;
													assign node13298 = (inp[10]) ? node13300 : 4'b0100;
														assign node13300 = (inp[3]) ? 4'b0000 : 4'b0000;
									assign node13303 = (inp[15]) ? node13349 : node13304;
										assign node13304 = (inp[3]) ? node13322 : node13305;
											assign node13305 = (inp[4]) ? node13317 : node13306;
												assign node13306 = (inp[9]) ? node13312 : node13307;
													assign node13307 = (inp[12]) ? node13309 : 4'b0100;
														assign node13309 = (inp[10]) ? 4'b0000 : 4'b0100;
													assign node13312 = (inp[12]) ? node13314 : 4'b0000;
														assign node13314 = (inp[2]) ? 4'b0000 : 4'b0100;
												assign node13317 = (inp[9]) ? node13319 : 4'b0000;
													assign node13319 = (inp[5]) ? 4'b0110 : 4'b0100;
											assign node13322 = (inp[5]) ? node13338 : node13323;
												assign node13323 = (inp[4]) ? node13331 : node13324;
													assign node13324 = (inp[9]) ? node13328 : node13325;
														assign node13325 = (inp[10]) ? 4'b0000 : 4'b0100;
														assign node13328 = (inp[10]) ? 4'b0000 : 4'b0000;
													assign node13331 = (inp[9]) ? node13335 : node13332;
														assign node13332 = (inp[12]) ? 4'b0110 : 4'b0000;
														assign node13335 = (inp[12]) ? 4'b0010 : 4'b0110;
												assign node13338 = (inp[12]) ? node13344 : node13339;
													assign node13339 = (inp[10]) ? 4'b0110 : node13340;
														assign node13340 = (inp[4]) ? 4'b0110 : 4'b0010;
													assign node13344 = (inp[10]) ? 4'b0010 : node13345;
														assign node13345 = (inp[9]) ? 4'b0110 : 4'b0010;
										assign node13349 = (inp[5]) ? node13367 : node13350;
											assign node13350 = (inp[4]) ? node13360 : node13351;
												assign node13351 = (inp[12]) ? node13353 : 4'b0010;
													assign node13353 = (inp[10]) ? node13357 : node13354;
														assign node13354 = (inp[9]) ? 4'b0010 : 4'b0110;
														assign node13357 = (inp[3]) ? 4'b0010 : 4'b0110;
												assign node13360 = (inp[9]) ? node13362 : 4'b0010;
													assign node13362 = (inp[10]) ? node13364 : 4'b0100;
														assign node13364 = (inp[12]) ? 4'b0010 : 4'b0110;
											assign node13367 = (inp[3]) ? node13381 : node13368;
												assign node13368 = (inp[9]) ? node13374 : node13369;
													assign node13369 = (inp[4]) ? 4'b0010 : node13370;
														assign node13370 = (inp[12]) ? 4'b0010 : 4'b0110;
													assign node13374 = (inp[4]) ? node13378 : node13375;
														assign node13375 = (inp[12]) ? 4'b0100 : 4'b0010;
														assign node13378 = (inp[12]) ? 4'b0000 : 4'b0100;
												assign node13381 = (inp[12]) ? node13383 : 4'b0000;
													assign node13383 = (inp[9]) ? node13387 : node13384;
														assign node13384 = (inp[10]) ? 4'b0100 : 4'b0000;
														assign node13387 = (inp[2]) ? 4'b0000 : 4'b0000;
						assign node13390 = (inp[15]) ? node13754 : node13391;
							assign node13391 = (inp[5]) ? node13575 : node13392;
								assign node13392 = (inp[3]) ? node13484 : node13393;
									assign node13393 = (inp[4]) ? node13435 : node13394;
										assign node13394 = (inp[9]) ? node13412 : node13395;
											assign node13395 = (inp[10]) ? node13403 : node13396;
												assign node13396 = (inp[2]) ? node13398 : 4'b0101;
													assign node13398 = (inp[8]) ? 4'b0101 : node13399;
														assign node13399 = (inp[7]) ? 4'b0101 : 4'b0100;
												assign node13403 = (inp[12]) ? node13407 : node13404;
													assign node13404 = (inp[8]) ? 4'b0101 : 4'b0100;
													assign node13407 = (inp[7]) ? node13409 : 4'b0001;
														assign node13409 = (inp[2]) ? 4'b0000 : 4'b0000;
											assign node13412 = (inp[14]) ? node13424 : node13413;
												assign node13413 = (inp[10]) ? node13419 : node13414;
													assign node13414 = (inp[12]) ? node13416 : 4'b0000;
														assign node13416 = (inp[8]) ? 4'b0000 : 4'b0001;
													assign node13419 = (inp[2]) ? node13421 : 4'b0000;
														assign node13421 = (inp[12]) ? 4'b0101 : 4'b0001;
												assign node13424 = (inp[12]) ? node13430 : node13425;
													assign node13425 = (inp[8]) ? node13427 : 4'b0001;
														assign node13427 = (inp[7]) ? 4'b0000 : 4'b0001;
													assign node13430 = (inp[10]) ? 4'b0101 : node13431;
														assign node13431 = (inp[8]) ? 4'b0001 : 4'b0000;
										assign node13435 = (inp[9]) ? node13459 : node13436;
											assign node13436 = (inp[12]) ? node13448 : node13437;
												assign node13437 = (inp[8]) ? node13443 : node13438;
													assign node13438 = (inp[7]) ? 4'b0001 : node13439;
														assign node13439 = (inp[14]) ? 4'b0000 : 4'b0001;
													assign node13443 = (inp[10]) ? node13445 : 4'b0000;
														assign node13445 = (inp[2]) ? 4'b0000 : 4'b0001;
												assign node13448 = (inp[10]) ? node13454 : node13449;
													assign node13449 = (inp[2]) ? 4'b0001 : node13450;
														assign node13450 = (inp[7]) ? 4'b0000 : 4'b0000;
													assign node13454 = (inp[8]) ? node13456 : 4'b0101;
														assign node13456 = (inp[7]) ? 4'b0100 : 4'b0100;
											assign node13459 = (inp[10]) ? node13473 : node13460;
												assign node13460 = (inp[7]) ? node13468 : node13461;
													assign node13461 = (inp[8]) ? node13465 : node13462;
														assign node13462 = (inp[12]) ? 4'b0100 : 4'b0101;
														assign node13465 = (inp[14]) ? 4'b0101 : 4'b0100;
													assign node13468 = (inp[14]) ? node13470 : 4'b0101;
														assign node13470 = (inp[8]) ? 4'b0100 : 4'b0101;
												assign node13473 = (inp[12]) ? node13479 : node13474;
													assign node13474 = (inp[2]) ? 4'b0100 : node13475;
														assign node13475 = (inp[14]) ? 4'b0100 : 4'b0101;
													assign node13479 = (inp[7]) ? node13481 : 4'b0000;
														assign node13481 = (inp[14]) ? 4'b0000 : 4'b0001;
									assign node13484 = (inp[9]) ? node13526 : node13485;
										assign node13485 = (inp[4]) ? node13503 : node13486;
											assign node13486 = (inp[12]) ? node13492 : node13487;
												assign node13487 = (inp[10]) ? 4'b0101 : node13488;
													assign node13488 = (inp[7]) ? 4'b0101 : 4'b0100;
												assign node13492 = (inp[10]) ? node13498 : node13493;
													assign node13493 = (inp[7]) ? 4'b0101 : node13494;
														assign node13494 = (inp[14]) ? 4'b0100 : 4'b0101;
													assign node13498 = (inp[8]) ? 4'b0000 : node13499;
														assign node13499 = (inp[14]) ? 4'b0001 : 4'b0000;
											assign node13503 = (inp[10]) ? node13517 : node13504;
												assign node13504 = (inp[14]) ? node13512 : node13505;
													assign node13505 = (inp[7]) ? node13509 : node13506;
														assign node13506 = (inp[12]) ? 4'b0001 : 4'b0000;
														assign node13509 = (inp[12]) ? 4'b0000 : 4'b0001;
													assign node13512 = (inp[7]) ? 4'b0001 : node13513;
														assign node13513 = (inp[8]) ? 4'b0001 : 4'b0000;
												assign node13517 = (inp[12]) ? node13521 : node13518;
													assign node13518 = (inp[14]) ? 4'b0001 : 4'b0000;
													assign node13521 = (inp[14]) ? 4'b0110 : node13522;
														assign node13522 = (inp[2]) ? 4'b0111 : 4'b0110;
										assign node13526 = (inp[4]) ? node13554 : node13527;
											assign node13527 = (inp[12]) ? node13541 : node13528;
												assign node13528 = (inp[2]) ? node13534 : node13529;
													assign node13529 = (inp[7]) ? 4'b0000 : node13530;
														assign node13530 = (inp[14]) ? 4'b0000 : 4'b0000;
													assign node13534 = (inp[8]) ? node13538 : node13535;
														assign node13535 = (inp[7]) ? 4'b0001 : 4'b0000;
														assign node13538 = (inp[7]) ? 4'b0000 : 4'b0001;
												assign node13541 = (inp[10]) ? node13547 : node13542;
													assign node13542 = (inp[8]) ? 4'b0001 : node13543;
														assign node13543 = (inp[2]) ? 4'b0000 : 4'b0000;
													assign node13547 = (inp[8]) ? node13551 : node13548;
														assign node13548 = (inp[7]) ? 4'b0111 : 4'b0110;
														assign node13551 = (inp[7]) ? 4'b0110 : 4'b0111;
											assign node13554 = (inp[10]) ? node13564 : node13555;
												assign node13555 = (inp[14]) ? node13557 : 4'b0110;
													assign node13557 = (inp[8]) ? node13561 : node13558;
														assign node13558 = (inp[7]) ? 4'b0111 : 4'b0110;
														assign node13561 = (inp[7]) ? 4'b0110 : 4'b0111;
												assign node13564 = (inp[12]) ? node13570 : node13565;
													assign node13565 = (inp[2]) ? 4'b0111 : node13566;
														assign node13566 = (inp[7]) ? 4'b0110 : 4'b0110;
													assign node13570 = (inp[14]) ? node13572 : 4'b0011;
														assign node13572 = (inp[7]) ? 4'b0011 : 4'b0010;
								assign node13575 = (inp[3]) ? node13671 : node13576;
									assign node13576 = (inp[9]) ? node13622 : node13577;
										assign node13577 = (inp[4]) ? node13599 : node13578;
											assign node13578 = (inp[10]) ? node13590 : node13579;
												assign node13579 = (inp[7]) ? node13585 : node13580;
													assign node13580 = (inp[12]) ? 4'b0100 : node13581;
														assign node13581 = (inp[14]) ? 4'b0100 : 4'b0101;
													assign node13585 = (inp[12]) ? 4'b0101 : node13586;
														assign node13586 = (inp[14]) ? 4'b0100 : 4'b0100;
												assign node13590 = (inp[12]) ? node13594 : node13591;
													assign node13591 = (inp[2]) ? 4'b0101 : 4'b0100;
													assign node13594 = (inp[7]) ? 4'b0001 : node13595;
														assign node13595 = (inp[14]) ? 4'b0000 : 4'b0000;
											assign node13599 = (inp[12]) ? node13611 : node13600;
												assign node13600 = (inp[14]) ? node13606 : node13601;
													assign node13601 = (inp[10]) ? 4'b0001 : node13602;
														assign node13602 = (inp[8]) ? 4'b0000 : 4'b0001;
													assign node13606 = (inp[7]) ? 4'b0000 : node13607;
														assign node13607 = (inp[8]) ? 4'b0001 : 4'b0000;
												assign node13611 = (inp[10]) ? node13617 : node13612;
													assign node13612 = (inp[8]) ? 4'b0000 : node13613;
														assign node13613 = (inp[7]) ? 4'b0001 : 4'b0000;
													assign node13617 = (inp[7]) ? 4'b0111 : node13618;
														assign node13618 = (inp[8]) ? 4'b0111 : 4'b0110;
										assign node13622 = (inp[4]) ? node13648 : node13623;
											assign node13623 = (inp[12]) ? node13635 : node13624;
												assign node13624 = (inp[7]) ? node13630 : node13625;
													assign node13625 = (inp[8]) ? node13627 : 4'b0000;
														assign node13627 = (inp[2]) ? 4'b0001 : 4'b0000;
													assign node13630 = (inp[10]) ? 4'b0001 : node13631;
														assign node13631 = (inp[14]) ? 4'b0001 : 4'b0000;
												assign node13635 = (inp[10]) ? node13641 : node13636;
													assign node13636 = (inp[8]) ? node13638 : 4'b0001;
														assign node13638 = (inp[7]) ? 4'b0000 : 4'b0001;
													assign node13641 = (inp[7]) ? node13645 : node13642;
														assign node13642 = (inp[2]) ? 4'b0110 : 4'b0110;
														assign node13645 = (inp[14]) ? 4'b0111 : 4'b0110;
											assign node13648 = (inp[10]) ? node13660 : node13649;
												assign node13649 = (inp[2]) ? node13655 : node13650;
													assign node13650 = (inp[8]) ? node13652 : 4'b0110;
														assign node13652 = (inp[14]) ? 4'b0111 : 4'b0110;
													assign node13655 = (inp[14]) ? 4'b0110 : node13656;
														assign node13656 = (inp[8]) ? 4'b0110 : 4'b0111;
												assign node13660 = (inp[12]) ? node13666 : node13661;
													assign node13661 = (inp[14]) ? node13663 : 4'b0110;
														assign node13663 = (inp[8]) ? 4'b0110 : 4'b0111;
													assign node13666 = (inp[7]) ? 4'b0011 : node13667;
														assign node13667 = (inp[8]) ? 4'b0010 : 4'b0010;
									assign node13671 = (inp[9]) ? node13713 : node13672;
										assign node13672 = (inp[4]) ? node13696 : node13673;
											assign node13673 = (inp[12]) ? node13685 : node13674;
												assign node13674 = (inp[2]) ? node13680 : node13675;
													assign node13675 = (inp[7]) ? node13677 : 4'b0111;
														assign node13677 = (inp[14]) ? 4'b0110 : 4'b0111;
													assign node13680 = (inp[14]) ? node13682 : 4'b0110;
														assign node13682 = (inp[8]) ? 4'b0111 : 4'b0110;
												assign node13685 = (inp[10]) ? node13691 : node13686;
													assign node13686 = (inp[8]) ? node13688 : 4'b0111;
														assign node13688 = (inp[7]) ? 4'b0110 : 4'b0110;
													assign node13691 = (inp[14]) ? 4'b0010 : node13692;
														assign node13692 = (inp[2]) ? 4'b0011 : 4'b0010;
											assign node13696 = (inp[12]) ? node13706 : node13697;
												assign node13697 = (inp[14]) ? node13701 : node13698;
													assign node13698 = (inp[2]) ? 4'b0010 : 4'b0011;
													assign node13701 = (inp[2]) ? 4'b0011 : node13702;
														assign node13702 = (inp[10]) ? 4'b0011 : 4'b0010;
												assign node13706 = (inp[10]) ? 4'b0110 : node13707;
													assign node13707 = (inp[2]) ? 4'b0010 : node13708;
														assign node13708 = (inp[8]) ? 4'b0010 : 4'b0010;
										assign node13713 = (inp[4]) ? node13731 : node13714;
											assign node13714 = (inp[12]) ? node13726 : node13715;
												assign node13715 = (inp[7]) ? node13721 : node13716;
													assign node13716 = (inp[2]) ? 4'b0011 : node13717;
														assign node13717 = (inp[8]) ? 4'b0010 : 4'b0010;
													assign node13721 = (inp[14]) ? 4'b0010 : node13722;
														assign node13722 = (inp[2]) ? 4'b0010 : 4'b0011;
												assign node13726 = (inp[10]) ? node13728 : 4'b0011;
													assign node13728 = (inp[7]) ? 4'b0110 : 4'b0111;
											assign node13731 = (inp[12]) ? node13745 : node13732;
												assign node13732 = (inp[14]) ? node13740 : node13733;
													assign node13733 = (inp[10]) ? node13737 : node13734;
														assign node13734 = (inp[7]) ? 4'b0110 : 4'b0111;
														assign node13737 = (inp[7]) ? 4'b0111 : 4'b0110;
													assign node13740 = (inp[8]) ? 4'b0110 : node13741;
														assign node13741 = (inp[7]) ? 4'b0111 : 4'b0110;
												assign node13745 = (inp[10]) ? node13751 : node13746;
													assign node13746 = (inp[7]) ? 4'b0110 : node13747;
														assign node13747 = (inp[8]) ? 4'b0111 : 4'b0110;
													assign node13751 = (inp[7]) ? 4'b0011 : 4'b0010;
							assign node13754 = (inp[3]) ? node13924 : node13755;
								assign node13755 = (inp[5]) ? node13831 : node13756;
									assign node13756 = (inp[4]) ? node13792 : node13757;
										assign node13757 = (inp[9]) ? node13773 : node13758;
											assign node13758 = (inp[10]) ? node13766 : node13759;
												assign node13759 = (inp[14]) ? 4'b0111 : node13760;
													assign node13760 = (inp[7]) ? node13762 : 4'b0110;
														assign node13762 = (inp[12]) ? 4'b0111 : 4'b0110;
												assign node13766 = (inp[12]) ? node13768 : 4'b0111;
													assign node13768 = (inp[2]) ? 4'b0011 : node13769;
														assign node13769 = (inp[14]) ? 4'b0010 : 4'b0011;
											assign node13773 = (inp[12]) ? node13783 : node13774;
												assign node13774 = (inp[7]) ? node13780 : node13775;
													assign node13775 = (inp[8]) ? 4'b0011 : node13776;
														assign node13776 = (inp[14]) ? 4'b0010 : 4'b0011;
													assign node13780 = (inp[8]) ? 4'b0010 : 4'b0011;
												assign node13783 = (inp[10]) ? node13785 : 4'b0011;
													assign node13785 = (inp[14]) ? node13789 : node13786;
														assign node13786 = (inp[8]) ? 4'b0111 : 4'b0110;
														assign node13789 = (inp[8]) ? 4'b0110 : 4'b0111;
										assign node13792 = (inp[9]) ? node13810 : node13793;
											assign node13793 = (inp[10]) ? node13807 : node13794;
												assign node13794 = (inp[14]) ? node13800 : node13795;
													assign node13795 = (inp[2]) ? 4'b0011 : node13796;
														assign node13796 = (inp[8]) ? 4'b0010 : 4'b0010;
													assign node13800 = (inp[8]) ? node13804 : node13801;
														assign node13801 = (inp[7]) ? 4'b0011 : 4'b0010;
														assign node13804 = (inp[7]) ? 4'b0010 : 4'b0011;
												assign node13807 = (inp[12]) ? 4'b0111 : 4'b0011;
											assign node13810 = (inp[10]) ? node13824 : node13811;
												assign node13811 = (inp[12]) ? node13817 : node13812;
													assign node13812 = (inp[14]) ? node13814 : 4'b0111;
														assign node13814 = (inp[7]) ? 4'b0110 : 4'b0110;
													assign node13817 = (inp[2]) ? node13821 : node13818;
														assign node13818 = (inp[8]) ? 4'b0110 : 4'b0110;
														assign node13821 = (inp[14]) ? 4'b0111 : 4'b0110;
												assign node13824 = (inp[12]) ? node13828 : node13825;
													assign node13825 = (inp[7]) ? 4'b0111 : 4'b0110;
													assign node13828 = (inp[7]) ? 4'b0010 : 4'b0011;
									assign node13831 = (inp[4]) ? node13875 : node13832;
										assign node13832 = (inp[9]) ? node13854 : node13833;
											assign node13833 = (inp[10]) ? node13845 : node13834;
												assign node13834 = (inp[8]) ? node13838 : node13835;
													assign node13835 = (inp[7]) ? 4'b0111 : 4'b0110;
													assign node13838 = (inp[7]) ? node13842 : node13839;
														assign node13839 = (inp[12]) ? 4'b0111 : 4'b0110;
														assign node13842 = (inp[14]) ? 4'b0110 : 4'b0110;
												assign node13845 = (inp[12]) ? node13847 : 4'b0111;
													assign node13847 = (inp[14]) ? node13851 : node13848;
														assign node13848 = (inp[7]) ? 4'b0010 : 4'b0010;
														assign node13851 = (inp[2]) ? 4'b0011 : 4'b0011;
											assign node13854 = (inp[10]) ? node13866 : node13855;
												assign node13855 = (inp[12]) ? node13861 : node13856;
													assign node13856 = (inp[14]) ? 4'b0010 : node13857;
														assign node13857 = (inp[7]) ? 4'b0010 : 4'b0011;
													assign node13861 = (inp[8]) ? 4'b0011 : node13862;
														assign node13862 = (inp[7]) ? 4'b0011 : 4'b0010;
												assign node13866 = (inp[12]) ? node13870 : node13867;
													assign node13867 = (inp[2]) ? 4'b0011 : 4'b0010;
													assign node13870 = (inp[2]) ? 4'b0100 : node13871;
														assign node13871 = (inp[8]) ? 4'b0100 : 4'b0101;
										assign node13875 = (inp[9]) ? node13899 : node13876;
											assign node13876 = (inp[12]) ? node13888 : node13877;
												assign node13877 = (inp[2]) ? node13885 : node13878;
													assign node13878 = (inp[7]) ? node13882 : node13879;
														assign node13879 = (inp[8]) ? 4'b0010 : 4'b0011;
														assign node13882 = (inp[10]) ? 4'b0011 : 4'b0010;
													assign node13885 = (inp[10]) ? 4'b0010 : 4'b0011;
												assign node13888 = (inp[10]) ? node13894 : node13889;
													assign node13889 = (inp[8]) ? node13891 : 4'b0011;
														assign node13891 = (inp[7]) ? 4'b0010 : 4'b0011;
													assign node13894 = (inp[2]) ? node13896 : 4'b0101;
														assign node13896 = (inp[8]) ? 4'b0100 : 4'b0100;
											assign node13899 = (inp[10]) ? node13911 : node13900;
												assign node13900 = (inp[7]) ? node13906 : node13901;
													assign node13901 = (inp[8]) ? node13903 : 4'b0100;
														assign node13903 = (inp[12]) ? 4'b0101 : 4'b0100;
													assign node13906 = (inp[8]) ? node13908 : 4'b0101;
														assign node13908 = (inp[2]) ? 4'b0100 : 4'b0101;
												assign node13911 = (inp[12]) ? node13919 : node13912;
													assign node13912 = (inp[7]) ? node13916 : node13913;
														assign node13913 = (inp[8]) ? 4'b0101 : 4'b0100;
														assign node13916 = (inp[8]) ? 4'b0100 : 4'b0101;
													assign node13919 = (inp[14]) ? node13921 : 4'b0000;
														assign node13921 = (inp[2]) ? 4'b0001 : 4'b0001;
								assign node13924 = (inp[5]) ? node14016 : node13925;
									assign node13925 = (inp[9]) ? node13967 : node13926;
										assign node13926 = (inp[4]) ? node13950 : node13927;
											assign node13927 = (inp[10]) ? node13939 : node13928;
												assign node13928 = (inp[12]) ? node13934 : node13929;
													assign node13929 = (inp[14]) ? 4'b0110 : node13930;
														assign node13930 = (inp[8]) ? 4'b0110 : 4'b0110;
													assign node13934 = (inp[7]) ? node13936 : 4'b0111;
														assign node13936 = (inp[8]) ? 4'b0110 : 4'b0110;
												assign node13939 = (inp[12]) ? node13945 : node13940;
													assign node13940 = (inp[2]) ? node13942 : 4'b0110;
														assign node13942 = (inp[8]) ? 4'b0110 : 4'b0111;
													assign node13945 = (inp[8]) ? node13947 : 4'b0011;
														assign node13947 = (inp[7]) ? 4'b0010 : 4'b0011;
											assign node13950 = (inp[12]) ? node13962 : node13951;
												assign node13951 = (inp[2]) ? node13955 : node13952;
													assign node13952 = (inp[7]) ? 4'b0011 : 4'b0010;
													assign node13955 = (inp[8]) ? node13959 : node13956;
														assign node13956 = (inp[7]) ? 4'b0011 : 4'b0010;
														assign node13959 = (inp[7]) ? 4'b0010 : 4'b0011;
												assign node13962 = (inp[10]) ? 4'b0100 : node13963;
													assign node13963 = (inp[7]) ? 4'b0011 : 4'b0010;
										assign node13967 = (inp[4]) ? node13993 : node13968;
											assign node13968 = (inp[10]) ? node13982 : node13969;
												assign node13969 = (inp[14]) ? node13975 : node13970;
													assign node13970 = (inp[8]) ? 4'b0011 : node13971;
														assign node13971 = (inp[2]) ? 4'b0011 : 4'b0010;
													assign node13975 = (inp[7]) ? node13979 : node13976;
														assign node13976 = (inp[8]) ? 4'b0011 : 4'b0010;
														assign node13979 = (inp[8]) ? 4'b0010 : 4'b0011;
												assign node13982 = (inp[12]) ? node13988 : node13983;
													assign node13983 = (inp[2]) ? 4'b0010 : node13984;
														assign node13984 = (inp[8]) ? 4'b0010 : 4'b0011;
													assign node13988 = (inp[8]) ? 4'b0101 : node13989;
														assign node13989 = (inp[2]) ? 4'b0100 : 4'b0100;
											assign node13993 = (inp[10]) ? node14001 : node13994;
												assign node13994 = (inp[8]) ? node13996 : 4'b0101;
													assign node13996 = (inp[7]) ? 4'b0100 : node13997;
														assign node13997 = (inp[14]) ? 4'b0101 : 4'b0101;
												assign node14001 = (inp[12]) ? node14009 : node14002;
													assign node14002 = (inp[2]) ? node14006 : node14003;
														assign node14003 = (inp[8]) ? 4'b0100 : 4'b0101;
														assign node14006 = (inp[8]) ? 4'b0101 : 4'b0100;
													assign node14009 = (inp[14]) ? node14013 : node14010;
														assign node14010 = (inp[8]) ? 4'b0000 : 4'b0000;
														assign node14013 = (inp[8]) ? 4'b0001 : 4'b0000;
									assign node14016 = (inp[9]) ? node14054 : node14017;
										assign node14017 = (inp[4]) ? node14031 : node14018;
											assign node14018 = (inp[10]) ? node14026 : node14019;
												assign node14019 = (inp[12]) ? node14021 : 4'b0101;
													assign node14021 = (inp[7]) ? 4'b0101 : node14022;
														assign node14022 = (inp[8]) ? 4'b0101 : 4'b0100;
												assign node14026 = (inp[12]) ? 4'b0000 : node14027;
													assign node14027 = (inp[2]) ? 4'b0100 : 4'b0101;
											assign node14031 = (inp[12]) ? node14045 : node14032;
												assign node14032 = (inp[10]) ? node14040 : node14033;
													assign node14033 = (inp[2]) ? node14037 : node14034;
														assign node14034 = (inp[8]) ? 4'b0000 : 4'b0001;
														assign node14037 = (inp[8]) ? 4'b0001 : 4'b0000;
													assign node14040 = (inp[7]) ? node14042 : 4'b0001;
														assign node14042 = (inp[2]) ? 4'b0001 : 4'b0000;
												assign node14045 = (inp[10]) ? node14051 : node14046;
													assign node14046 = (inp[8]) ? 4'b0001 : node14047;
														assign node14047 = (inp[7]) ? 4'b0001 : 4'b0000;
													assign node14051 = (inp[2]) ? 4'b0101 : 4'b0100;
										assign node14054 = (inp[4]) ? node14074 : node14055;
											assign node14055 = (inp[12]) ? node14063 : node14056;
												assign node14056 = (inp[7]) ? node14058 : 4'b0001;
													assign node14058 = (inp[8]) ? 4'b0000 : node14059;
														assign node14059 = (inp[14]) ? 4'b0001 : 4'b0000;
												assign node14063 = (inp[10]) ? node14069 : node14064;
													assign node14064 = (inp[8]) ? 4'b0001 : node14065;
														assign node14065 = (inp[14]) ? 4'b0000 : 4'b0001;
													assign node14069 = (inp[14]) ? node14071 : 4'b0100;
														assign node14071 = (inp[8]) ? 4'b0100 : 4'b0101;
											assign node14074 = (inp[12]) ? node14082 : node14075;
												assign node14075 = (inp[8]) ? node14077 : 4'b0100;
													assign node14077 = (inp[7]) ? node14079 : 4'b0101;
														assign node14079 = (inp[2]) ? 4'b0100 : 4'b0101;
												assign node14082 = (inp[10]) ? node14086 : node14083;
													assign node14083 = (inp[2]) ? 4'b0101 : 4'b0100;
													assign node14086 = (inp[14]) ? 4'b0000 : node14087;
														assign node14087 = (inp[8]) ? 4'b0000 : 4'b0001;
				assign node14091 = (inp[1]) ? node15517 : node14092;
					assign node14092 = (inp[13]) ? node14792 : node14093;
						assign node14093 = (inp[15]) ? node14427 : node14094;
							assign node14094 = (inp[5]) ? node14256 : node14095;
								assign node14095 = (inp[3]) ? node14181 : node14096;
									assign node14096 = (inp[10]) ? node14140 : node14097;
										assign node14097 = (inp[8]) ? node14125 : node14098;
											assign node14098 = (inp[14]) ? node14112 : node14099;
												assign node14099 = (inp[7]) ? node14107 : node14100;
													assign node14100 = (inp[2]) ? node14104 : node14101;
														assign node14101 = (inp[4]) ? 4'b0101 : 4'b0101;
														assign node14104 = (inp[9]) ? 4'b0100 : 4'b0000;
													assign node14107 = (inp[9]) ? node14109 : 4'b0100;
														assign node14109 = (inp[4]) ? 4'b0100 : 4'b0000;
												assign node14112 = (inp[7]) ? node14118 : node14113;
													assign node14113 = (inp[12]) ? 4'b0000 : node14114;
														assign node14114 = (inp[9]) ? 4'b0000 : 4'b0100;
													assign node14118 = (inp[2]) ? node14122 : node14119;
														assign node14119 = (inp[4]) ? 4'b0001 : 4'b0001;
														assign node14122 = (inp[12]) ? 4'b0001 : 4'b0101;
											assign node14125 = (inp[2]) ? node14133 : node14126;
												assign node14126 = (inp[12]) ? node14128 : 4'b0000;
													assign node14128 = (inp[4]) ? node14130 : 4'b0001;
														assign node14130 = (inp[14]) ? 4'b0000 : 4'b0000;
												assign node14133 = (inp[7]) ? node14137 : node14134;
													assign node14134 = (inp[12]) ? 4'b0101 : 4'b0001;
													assign node14137 = (inp[12]) ? 4'b0000 : 4'b0100;
										assign node14140 = (inp[4]) ? node14160 : node14141;
											assign node14141 = (inp[9]) ? node14153 : node14142;
												assign node14142 = (inp[12]) ? node14148 : node14143;
													assign node14143 = (inp[14]) ? 4'b0101 : node14144;
														assign node14144 = (inp[2]) ? 4'b0101 : 4'b0100;
													assign node14148 = (inp[7]) ? 4'b0001 : node14149;
														assign node14149 = (inp[8]) ? 4'b0001 : 4'b0000;
												assign node14153 = (inp[12]) ? node14157 : node14154;
													assign node14154 = (inp[8]) ? 4'b0000 : 4'b0001;
													assign node14157 = (inp[2]) ? 4'b0100 : 4'b0101;
											assign node14160 = (inp[9]) ? node14170 : node14161;
												assign node14161 = (inp[12]) ? node14167 : node14162;
													assign node14162 = (inp[14]) ? 4'b0000 : node14163;
														assign node14163 = (inp[7]) ? 4'b0000 : 4'b0001;
													assign node14167 = (inp[2]) ? 4'b0101 : 4'b0100;
												assign node14170 = (inp[12]) ? node14176 : node14171;
													assign node14171 = (inp[2]) ? node14173 : 4'b0100;
														assign node14173 = (inp[7]) ? 4'b0100 : 4'b0101;
													assign node14176 = (inp[2]) ? node14178 : 4'b0000;
														assign node14178 = (inp[7]) ? 4'b0001 : 4'b0000;
									assign node14181 = (inp[9]) ? node14219 : node14182;
										assign node14182 = (inp[4]) ? node14202 : node14183;
											assign node14183 = (inp[12]) ? node14193 : node14184;
												assign node14184 = (inp[2]) ? node14186 : 4'b0101;
													assign node14186 = (inp[14]) ? node14190 : node14187;
														assign node14187 = (inp[7]) ? 4'b0101 : 4'b0100;
														assign node14190 = (inp[8]) ? 4'b0100 : 4'b0101;
												assign node14193 = (inp[10]) ? node14197 : node14194;
													assign node14194 = (inp[2]) ? 4'b0100 : 4'b0101;
													assign node14197 = (inp[8]) ? node14199 : 4'b0000;
														assign node14199 = (inp[14]) ? 4'b0001 : 4'b0000;
											assign node14202 = (inp[10]) ? node14214 : node14203;
												assign node14203 = (inp[14]) ? node14209 : node14204;
													assign node14204 = (inp[8]) ? 4'b0001 : node14205;
														assign node14205 = (inp[2]) ? 4'b0000 : 4'b0001;
													assign node14209 = (inp[2]) ? 4'b0000 : node14210;
														assign node14210 = (inp[7]) ? 4'b0000 : 4'b0000;
												assign node14214 = (inp[12]) ? 4'b0110 : node14215;
													assign node14215 = (inp[7]) ? 4'b0000 : 4'b0001;
										assign node14219 = (inp[4]) ? node14241 : node14220;
											assign node14220 = (inp[10]) ? node14232 : node14221;
												assign node14221 = (inp[7]) ? node14227 : node14222;
													assign node14222 = (inp[8]) ? node14224 : 4'b0000;
														assign node14224 = (inp[2]) ? 4'b0001 : 4'b0000;
													assign node14227 = (inp[8]) ? 4'b0000 : node14228;
														assign node14228 = (inp[2]) ? 4'b0001 : 4'b0000;
												assign node14232 = (inp[12]) ? node14238 : node14233;
													assign node14233 = (inp[8]) ? 4'b0001 : node14234;
														assign node14234 = (inp[7]) ? 4'b0000 : 4'b0000;
													assign node14238 = (inp[7]) ? 4'b0110 : 4'b0111;
											assign node14241 = (inp[10]) ? node14249 : node14242;
												assign node14242 = (inp[8]) ? node14244 : 4'b0110;
													assign node14244 = (inp[12]) ? 4'b0110 : node14245;
														assign node14245 = (inp[2]) ? 4'b0111 : 4'b0110;
												assign node14249 = (inp[12]) ? node14253 : node14250;
													assign node14250 = (inp[7]) ? 4'b0110 : 4'b0111;
													assign node14253 = (inp[7]) ? 4'b0011 : 4'b0010;
								assign node14256 = (inp[3]) ? node14334 : node14257;
									assign node14257 = (inp[9]) ? node14295 : node14258;
										assign node14258 = (inp[4]) ? node14276 : node14259;
											assign node14259 = (inp[10]) ? node14267 : node14260;
												assign node14260 = (inp[2]) ? node14262 : 4'b0101;
													assign node14262 = (inp[8]) ? node14264 : 4'b0100;
														assign node14264 = (inp[14]) ? 4'b0101 : 4'b0100;
												assign node14267 = (inp[12]) ? node14271 : node14268;
													assign node14268 = (inp[8]) ? 4'b0100 : 4'b0101;
													assign node14271 = (inp[14]) ? node14273 : 4'b0001;
														assign node14273 = (inp[7]) ? 4'b0000 : 4'b0001;
											assign node14276 = (inp[10]) ? node14286 : node14277;
												assign node14277 = (inp[7]) ? node14283 : node14278;
													assign node14278 = (inp[8]) ? node14280 : 4'b0000;
														assign node14280 = (inp[14]) ? 4'b0001 : 4'b0000;
													assign node14283 = (inp[8]) ? 4'b0000 : 4'b0001;
												assign node14286 = (inp[12]) ? node14292 : node14287;
													assign node14287 = (inp[7]) ? node14289 : 4'b0000;
														assign node14289 = (inp[2]) ? 4'b0000 : 4'b0001;
													assign node14292 = (inp[7]) ? 4'b0111 : 4'b0110;
										assign node14295 = (inp[4]) ? node14319 : node14296;
											assign node14296 = (inp[12]) ? node14308 : node14297;
												assign node14297 = (inp[7]) ? node14303 : node14298;
													assign node14298 = (inp[14]) ? 4'b0000 : node14299;
														assign node14299 = (inp[8]) ? 4'b0000 : 4'b0001;
													assign node14303 = (inp[10]) ? node14305 : 4'b0001;
														assign node14305 = (inp[8]) ? 4'b0001 : 4'b0000;
												assign node14308 = (inp[10]) ? node14314 : node14309;
													assign node14309 = (inp[8]) ? node14311 : 4'b0001;
														assign node14311 = (inp[2]) ? 4'b0001 : 4'b0000;
													assign node14314 = (inp[8]) ? node14316 : 4'b0110;
														assign node14316 = (inp[14]) ? 4'b0111 : 4'b0110;
											assign node14319 = (inp[12]) ? node14325 : node14320;
												assign node14320 = (inp[7]) ? node14322 : 4'b0111;
													assign node14322 = (inp[10]) ? 4'b0110 : 4'b0111;
												assign node14325 = (inp[10]) ? node14331 : node14326;
													assign node14326 = (inp[2]) ? node14328 : 4'b0110;
														assign node14328 = (inp[14]) ? 4'b0110 : 4'b0111;
													assign node14331 = (inp[8]) ? 4'b0011 : 4'b0010;
									assign node14334 = (inp[10]) ? node14376 : node14335;
										assign node14335 = (inp[7]) ? node14359 : node14336;
											assign node14336 = (inp[8]) ? node14344 : node14337;
												assign node14337 = (inp[14]) ? 4'b0110 : node14338;
													assign node14338 = (inp[2]) ? 4'b0110 : node14339;
														assign node14339 = (inp[4]) ? 4'b0011 : 4'b0111;
												assign node14344 = (inp[12]) ? node14352 : node14345;
													assign node14345 = (inp[14]) ? node14349 : node14346;
														assign node14346 = (inp[2]) ? 4'b0011 : 4'b0110;
														assign node14349 = (inp[9]) ? 4'b0011 : 4'b0011;
													assign node14352 = (inp[2]) ? node14356 : node14353;
														assign node14353 = (inp[4]) ? 4'b0011 : 4'b0111;
														assign node14356 = (inp[4]) ? 4'b0111 : 4'b0011;
											assign node14359 = (inp[8]) ? node14369 : node14360;
												assign node14360 = (inp[9]) ? node14364 : node14361;
													assign node14361 = (inp[4]) ? 4'b0011 : 4'b0111;
													assign node14364 = (inp[4]) ? 4'b0111 : node14365;
														assign node14365 = (inp[2]) ? 4'b0011 : 4'b0010;
												assign node14369 = (inp[2]) ? 4'b0110 : node14370;
													assign node14370 = (inp[9]) ? node14372 : 4'b0110;
														assign node14372 = (inp[4]) ? 4'b0110 : 4'b0010;
										assign node14376 = (inp[9]) ? node14404 : node14377;
											assign node14377 = (inp[7]) ? node14391 : node14378;
												assign node14378 = (inp[8]) ? node14386 : node14379;
													assign node14379 = (inp[12]) ? node14383 : node14380;
														assign node14380 = (inp[4]) ? 4'b0010 : 4'b0110;
														assign node14383 = (inp[4]) ? 4'b0110 : 4'b0010;
													assign node14386 = (inp[4]) ? node14388 : 4'b0111;
														assign node14388 = (inp[14]) ? 4'b0111 : 4'b0110;
												assign node14391 = (inp[8]) ? node14399 : node14392;
													assign node14392 = (inp[14]) ? node14396 : node14393;
														assign node14393 = (inp[4]) ? 4'b0111 : 4'b0010;
														assign node14396 = (inp[2]) ? 4'b0011 : 4'b0111;
													assign node14399 = (inp[2]) ? 4'b0110 : node14400;
														assign node14400 = (inp[14]) ? 4'b0010 : 4'b0011;
											assign node14404 = (inp[2]) ? node14418 : node14405;
												assign node14405 = (inp[12]) ? node14413 : node14406;
													assign node14406 = (inp[4]) ? node14410 : node14407;
														assign node14407 = (inp[7]) ? 4'b0011 : 4'b0010;
														assign node14410 = (inp[8]) ? 4'b0110 : 4'b0110;
													assign node14413 = (inp[4]) ? node14415 : 4'b0111;
														assign node14415 = (inp[7]) ? 4'b0011 : 4'b0011;
												assign node14418 = (inp[8]) ? node14424 : node14419;
													assign node14419 = (inp[14]) ? 4'b0010 : node14420;
														assign node14420 = (inp[4]) ? 4'b0010 : 4'b0110;
													assign node14424 = (inp[7]) ? 4'b0010 : 4'b0011;
							assign node14427 = (inp[3]) ? node14605 : node14428;
								assign node14428 = (inp[5]) ? node14520 : node14429;
									assign node14429 = (inp[7]) ? node14471 : node14430;
										assign node14430 = (inp[8]) ? node14456 : node14431;
											assign node14431 = (inp[14]) ? node14443 : node14432;
												assign node14432 = (inp[2]) ? node14438 : node14433;
													assign node14433 = (inp[9]) ? node14435 : 4'b0011;
														assign node14435 = (inp[10]) ? 4'b0111 : 4'b0011;
													assign node14438 = (inp[12]) ? 4'b0110 : node14439;
														assign node14439 = (inp[9]) ? 4'b0010 : 4'b0110;
												assign node14443 = (inp[12]) ? node14451 : node14444;
													assign node14444 = (inp[10]) ? node14448 : node14445;
														assign node14445 = (inp[9]) ? 4'b0010 : 4'b0110;
														assign node14448 = (inp[9]) ? 4'b0110 : 4'b0010;
													assign node14451 = (inp[9]) ? node14453 : 4'b0010;
														assign node14453 = (inp[10]) ? 4'b0110 : 4'b0010;
											assign node14456 = (inp[2]) ? node14462 : node14457;
												assign node14457 = (inp[14]) ? 4'b0111 : node14458;
													assign node14458 = (inp[9]) ? 4'b0110 : 4'b0010;
												assign node14462 = (inp[14]) ? node14468 : node14463;
													assign node14463 = (inp[9]) ? node14465 : 4'b0011;
														assign node14465 = (inp[12]) ? 4'b0111 : 4'b0011;
													assign node14468 = (inp[12]) ? 4'b0011 : 4'b0111;
										assign node14471 = (inp[8]) ? node14499 : node14472;
											assign node14472 = (inp[2]) ? node14486 : node14473;
												assign node14473 = (inp[14]) ? node14479 : node14474;
													assign node14474 = (inp[4]) ? 4'b0110 : node14475;
														assign node14475 = (inp[9]) ? 4'b0010 : 4'b0110;
													assign node14479 = (inp[9]) ? node14483 : node14480;
														assign node14480 = (inp[4]) ? 4'b0011 : 4'b0111;
														assign node14483 = (inp[10]) ? 4'b0011 : 4'b0011;
												assign node14486 = (inp[9]) ? node14494 : node14487;
													assign node14487 = (inp[4]) ? node14491 : node14488;
														assign node14488 = (inp[12]) ? 4'b0011 : 4'b0111;
														assign node14491 = (inp[12]) ? 4'b0011 : 4'b0011;
													assign node14494 = (inp[4]) ? 4'b0111 : node14495;
														assign node14495 = (inp[12]) ? 4'b0011 : 4'b0011;
											assign node14499 = (inp[2]) ? node14509 : node14500;
												assign node14500 = (inp[14]) ? node14506 : node14501;
													assign node14501 = (inp[12]) ? node14503 : 4'b0011;
														assign node14503 = (inp[10]) ? 4'b0111 : 4'b0011;
													assign node14506 = (inp[4]) ? 4'b0110 : 4'b0010;
												assign node14509 = (inp[10]) ? node14515 : node14510;
													assign node14510 = (inp[12]) ? 4'b0010 : node14511;
														assign node14511 = (inp[4]) ? 4'b0010 : 4'b0110;
													assign node14515 = (inp[12]) ? 4'b0110 : node14516;
														assign node14516 = (inp[9]) ? 4'b0010 : 4'b0110;
									assign node14520 = (inp[4]) ? node14564 : node14521;
										assign node14521 = (inp[9]) ? node14547 : node14522;
											assign node14522 = (inp[10]) ? node14536 : node14523;
												assign node14523 = (inp[12]) ? node14529 : node14524;
													assign node14524 = (inp[7]) ? 4'b0111 : node14525;
														assign node14525 = (inp[14]) ? 4'b0110 : 4'b0111;
													assign node14529 = (inp[7]) ? node14533 : node14530;
														assign node14530 = (inp[2]) ? 4'b0110 : 4'b0111;
														assign node14533 = (inp[8]) ? 4'b0110 : 4'b0111;
												assign node14536 = (inp[12]) ? node14542 : node14537;
													assign node14537 = (inp[8]) ? 4'b0111 : node14538;
														assign node14538 = (inp[14]) ? 4'b0111 : 4'b0110;
													assign node14542 = (inp[14]) ? node14544 : 4'b0011;
														assign node14544 = (inp[7]) ? 4'b0011 : 4'b0010;
											assign node14547 = (inp[10]) ? node14557 : node14548;
												assign node14548 = (inp[8]) ? node14552 : node14549;
													assign node14549 = (inp[14]) ? 4'b0011 : 4'b0010;
													assign node14552 = (inp[2]) ? 4'b0011 : node14553;
														assign node14553 = (inp[12]) ? 4'b0010 : 4'b0011;
												assign node14557 = (inp[12]) ? 4'b0100 : node14558;
													assign node14558 = (inp[8]) ? 4'b0011 : node14559;
														assign node14559 = (inp[7]) ? 4'b0010 : 4'b0010;
										assign node14564 = (inp[9]) ? node14584 : node14565;
											assign node14565 = (inp[10]) ? node14577 : node14566;
												assign node14566 = (inp[14]) ? node14572 : node14567;
													assign node14567 = (inp[2]) ? node14569 : 4'b0010;
														assign node14569 = (inp[7]) ? 4'b0010 : 4'b0010;
													assign node14572 = (inp[7]) ? 4'b0011 : node14573;
														assign node14573 = (inp[8]) ? 4'b0011 : 4'b0010;
												assign node14577 = (inp[12]) ? node14579 : 4'b0011;
													assign node14579 = (inp[2]) ? 4'b0100 : node14580;
														assign node14580 = (inp[7]) ? 4'b0100 : 4'b0101;
											assign node14584 = (inp[12]) ? node14592 : node14585;
												assign node14585 = (inp[8]) ? 4'b0100 : node14586;
													assign node14586 = (inp[14]) ? node14588 : 4'b0101;
														assign node14588 = (inp[7]) ? 4'b0101 : 4'b0100;
												assign node14592 = (inp[10]) ? node14598 : node14593;
													assign node14593 = (inp[2]) ? 4'b0101 : node14594;
														assign node14594 = (inp[8]) ? 4'b0101 : 4'b0100;
													assign node14598 = (inp[14]) ? node14602 : node14599;
														assign node14599 = (inp[7]) ? 4'b0000 : 4'b0001;
														assign node14602 = (inp[8]) ? 4'b0000 : 4'b0000;
								assign node14605 = (inp[5]) ? node14695 : node14606;
									assign node14606 = (inp[4]) ? node14654 : node14607;
										assign node14607 = (inp[9]) ? node14633 : node14608;
											assign node14608 = (inp[12]) ? node14622 : node14609;
												assign node14609 = (inp[14]) ? node14617 : node14610;
													assign node14610 = (inp[7]) ? node14614 : node14611;
														assign node14611 = (inp[10]) ? 4'b0110 : 4'b0110;
														assign node14614 = (inp[2]) ? 4'b0111 : 4'b0110;
													assign node14617 = (inp[10]) ? 4'b0110 : node14618;
														assign node14618 = (inp[2]) ? 4'b0110 : 4'b0110;
												assign node14622 = (inp[10]) ? node14628 : node14623;
													assign node14623 = (inp[7]) ? 4'b0111 : node14624;
														assign node14624 = (inp[8]) ? 4'b0111 : 4'b0110;
													assign node14628 = (inp[14]) ? 4'b0011 : node14629;
														assign node14629 = (inp[7]) ? 4'b0010 : 4'b0011;
											assign node14633 = (inp[10]) ? node14645 : node14634;
												assign node14634 = (inp[2]) ? node14640 : node14635;
													assign node14635 = (inp[12]) ? node14637 : 4'b0010;
														assign node14637 = (inp[14]) ? 4'b0011 : 4'b0010;
													assign node14640 = (inp[14]) ? 4'b0011 : node14641;
														assign node14641 = (inp[12]) ? 4'b0010 : 4'b0011;
												assign node14645 = (inp[12]) ? node14651 : node14646;
													assign node14646 = (inp[8]) ? 4'b0010 : node14647;
														assign node14647 = (inp[2]) ? 4'b0010 : 4'b0010;
													assign node14651 = (inp[14]) ? 4'b0100 : 4'b0101;
										assign node14654 = (inp[9]) ? node14672 : node14655;
											assign node14655 = (inp[10]) ? node14663 : node14656;
												assign node14656 = (inp[8]) ? 4'b0010 : node14657;
													assign node14657 = (inp[7]) ? node14659 : 4'b0010;
														assign node14659 = (inp[2]) ? 4'b0011 : 4'b0010;
												assign node14663 = (inp[12]) ? node14669 : node14664;
													assign node14664 = (inp[8]) ? node14666 : 4'b0011;
														assign node14666 = (inp[2]) ? 4'b0010 : 4'b0011;
													assign node14669 = (inp[14]) ? 4'b0101 : 4'b0100;
											assign node14672 = (inp[10]) ? node14686 : node14673;
												assign node14673 = (inp[2]) ? node14681 : node14674;
													assign node14674 = (inp[12]) ? node14678 : node14675;
														assign node14675 = (inp[14]) ? 4'b0100 : 4'b0100;
														assign node14678 = (inp[14]) ? 4'b0101 : 4'b0100;
													assign node14681 = (inp[12]) ? 4'b0100 : node14682;
														assign node14682 = (inp[8]) ? 4'b0101 : 4'b0100;
												assign node14686 = (inp[12]) ? node14690 : node14687;
													assign node14687 = (inp[8]) ? 4'b0100 : 4'b0101;
													assign node14690 = (inp[2]) ? 4'b0000 : node14691;
														assign node14691 = (inp[7]) ? 4'b0000 : 4'b0001;
									assign node14695 = (inp[2]) ? node14749 : node14696;
										assign node14696 = (inp[14]) ? node14724 : node14697;
											assign node14697 = (inp[9]) ? node14711 : node14698;
												assign node14698 = (inp[4]) ? node14704 : node14699;
													assign node14699 = (inp[12]) ? 4'b0001 : node14700;
														assign node14700 = (inp[10]) ? 4'b0100 : 4'b0100;
													assign node14704 = (inp[7]) ? node14708 : node14705;
														assign node14705 = (inp[8]) ? 4'b0000 : 4'b0001;
														assign node14708 = (inp[12]) ? 4'b0101 : 4'b0001;
												assign node14711 = (inp[4]) ? node14717 : node14712;
													assign node14712 = (inp[10]) ? node14714 : 4'b0000;
														assign node14714 = (inp[12]) ? 4'b0101 : 4'b0000;
													assign node14717 = (inp[10]) ? node14721 : node14718;
														assign node14718 = (inp[7]) ? 4'b0101 : 4'b0101;
														assign node14721 = (inp[12]) ? 4'b0000 : 4'b0100;
											assign node14724 = (inp[8]) ? node14736 : node14725;
												assign node14725 = (inp[7]) ? node14731 : node14726;
													assign node14726 = (inp[10]) ? node14728 : 4'b0000;
														assign node14728 = (inp[9]) ? 4'b0000 : 4'b0100;
													assign node14731 = (inp[9]) ? node14733 : 4'b0001;
														assign node14733 = (inp[4]) ? 4'b0101 : 4'b0001;
												assign node14736 = (inp[7]) ? node14742 : node14737;
													assign node14737 = (inp[10]) ? 4'b0001 : node14738;
														assign node14738 = (inp[12]) ? 4'b0101 : 4'b0001;
													assign node14742 = (inp[10]) ? node14746 : node14743;
														assign node14743 = (inp[9]) ? 4'b0000 : 4'b0100;
														assign node14746 = (inp[4]) ? 4'b0100 : 4'b0000;
										assign node14749 = (inp[12]) ? node14771 : node14750;
											assign node14750 = (inp[14]) ? node14758 : node14751;
												assign node14751 = (inp[10]) ? node14753 : 4'b0100;
													assign node14753 = (inp[4]) ? 4'b0100 : node14754;
														assign node14754 = (inp[9]) ? 4'b0000 : 4'b0100;
												assign node14758 = (inp[8]) ? node14766 : node14759;
													assign node14759 = (inp[7]) ? node14763 : node14760;
														assign node14760 = (inp[10]) ? 4'b0100 : 4'b0000;
														assign node14763 = (inp[9]) ? 4'b0101 : 4'b0001;
													assign node14766 = (inp[7]) ? node14768 : 4'b0001;
														assign node14768 = (inp[9]) ? 4'b0000 : 4'b0000;
											assign node14771 = (inp[7]) ? node14785 : node14772;
												assign node14772 = (inp[8]) ? node14780 : node14773;
													assign node14773 = (inp[10]) ? node14777 : node14774;
														assign node14774 = (inp[9]) ? 4'b0100 : 4'b0000;
														assign node14777 = (inp[9]) ? 4'b0000 : 4'b0100;
													assign node14780 = (inp[9]) ? node14782 : 4'b0001;
														assign node14782 = (inp[14]) ? 4'b0101 : 4'b0001;
												assign node14785 = (inp[8]) ? 4'b0100 : node14786;
													assign node14786 = (inp[10]) ? node14788 : 4'b0101;
														assign node14788 = (inp[9]) ? 4'b0001 : 4'b0101;
						assign node14792 = (inp[8]) ? node15184 : node14793;
							assign node14793 = (inp[7]) ? node14991 : node14794;
								assign node14794 = (inp[14]) ? node14890 : node14795;
									assign node14795 = (inp[2]) ? node14841 : node14796;
										assign node14796 = (inp[10]) ? node14820 : node14797;
											assign node14797 = (inp[12]) ? node14807 : node14798;
												assign node14798 = (inp[4]) ? node14804 : node14799;
													assign node14799 = (inp[9]) ? node14801 : 4'b0101;
														assign node14801 = (inp[15]) ? 4'b0001 : 4'b0001;
													assign node14804 = (inp[9]) ? 4'b0101 : 4'b0011;
												assign node14807 = (inp[4]) ? node14815 : node14808;
													assign node14808 = (inp[15]) ? node14812 : node14809;
														assign node14809 = (inp[5]) ? 4'b0111 : 4'b0101;
														assign node14812 = (inp[5]) ? 4'b0101 : 4'b0111;
													assign node14815 = (inp[9]) ? node14817 : 4'b0001;
														assign node14817 = (inp[15]) ? 4'b0101 : 4'b0111;
											assign node14820 = (inp[5]) ? node14828 : node14821;
												assign node14821 = (inp[15]) ? node14823 : 4'b0001;
													assign node14823 = (inp[9]) ? 4'b0011 : node14824;
														assign node14824 = (inp[12]) ? 4'b0111 : 4'b0011;
												assign node14828 = (inp[15]) ? node14834 : node14829;
													assign node14829 = (inp[12]) ? node14831 : 4'b0001;
														assign node14831 = (inp[9]) ? 4'b0011 : 4'b0111;
													assign node14834 = (inp[12]) ? node14838 : node14835;
														assign node14835 = (inp[3]) ? 4'b0101 : 4'b0111;
														assign node14838 = (inp[9]) ? 4'b0101 : 4'b0001;
										assign node14841 = (inp[9]) ? node14861 : node14842;
											assign node14842 = (inp[10]) ? node14850 : node14843;
												assign node14843 = (inp[4]) ? 4'b0010 : node14844;
													assign node14844 = (inp[15]) ? node14846 : 4'b0100;
														assign node14846 = (inp[5]) ? 4'b0100 : 4'b0110;
												assign node14850 = (inp[15]) ? node14856 : node14851;
													assign node14851 = (inp[5]) ? node14853 : 4'b0110;
														assign node14853 = (inp[12]) ? 4'b0010 : 4'b0110;
													assign node14856 = (inp[5]) ? node14858 : 4'b0010;
														assign node14858 = (inp[12]) ? 4'b0000 : 4'b0010;
											assign node14861 = (inp[4]) ? node14875 : node14862;
												assign node14862 = (inp[10]) ? node14870 : node14863;
													assign node14863 = (inp[5]) ? node14867 : node14864;
														assign node14864 = (inp[15]) ? 4'b0010 : 4'b0000;
														assign node14867 = (inp[3]) ? 4'b0000 : 4'b0000;
													assign node14870 = (inp[12]) ? node14872 : 4'b0000;
														assign node14872 = (inp[15]) ? 4'b0100 : 4'b0100;
												assign node14875 = (inp[10]) ? node14883 : node14876;
													assign node14876 = (inp[5]) ? node14880 : node14877;
														assign node14877 = (inp[12]) ? 4'b0100 : 4'b0100;
														assign node14880 = (inp[12]) ? 4'b0110 : 4'b0100;
													assign node14883 = (inp[12]) ? node14887 : node14884;
														assign node14884 = (inp[15]) ? 4'b0110 : 4'b0100;
														assign node14887 = (inp[5]) ? 4'b0010 : 4'b0000;
									assign node14890 = (inp[2]) ? node14936 : node14891;
										assign node14891 = (inp[15]) ? node14913 : node14892;
											assign node14892 = (inp[5]) ? node14906 : node14893;
												assign node14893 = (inp[10]) ? node14901 : node14894;
													assign node14894 = (inp[9]) ? node14898 : node14895;
														assign node14895 = (inp[4]) ? 4'b0000 : 4'b0100;
														assign node14898 = (inp[4]) ? 4'b0100 : 4'b0000;
													assign node14901 = (inp[9]) ? node14903 : 4'b0000;
														assign node14903 = (inp[12]) ? 4'b0100 : 4'b0000;
												assign node14906 = (inp[9]) ? node14910 : node14907;
													assign node14907 = (inp[3]) ? 4'b0010 : 4'b0110;
													assign node14910 = (inp[3]) ? 4'b0110 : 4'b0000;
											assign node14913 = (inp[3]) ? node14927 : node14914;
												assign node14914 = (inp[4]) ? node14922 : node14915;
													assign node14915 = (inp[9]) ? node14919 : node14916;
														assign node14916 = (inp[5]) ? 4'b0110 : 4'b0010;
														assign node14919 = (inp[12]) ? 4'b0010 : 4'b0010;
													assign node14922 = (inp[5]) ? 4'b0100 : node14923;
														assign node14923 = (inp[9]) ? 4'b0110 : 4'b0010;
												assign node14927 = (inp[10]) ? node14931 : node14928;
													assign node14928 = (inp[12]) ? 4'b0110 : 4'b0100;
													assign node14931 = (inp[12]) ? node14933 : 4'b0010;
														assign node14933 = (inp[9]) ? 4'b0000 : 4'b0000;
										assign node14936 = (inp[10]) ? node14966 : node14937;
											assign node14937 = (inp[12]) ? node14953 : node14938;
												assign node14938 = (inp[9]) ? node14946 : node14939;
													assign node14939 = (inp[4]) ? node14943 : node14940;
														assign node14940 = (inp[5]) ? 4'b0100 : 4'b0110;
														assign node14943 = (inp[15]) ? 4'b0010 : 4'b0000;
													assign node14946 = (inp[4]) ? node14950 : node14947;
														assign node14947 = (inp[5]) ? 4'b0010 : 4'b0000;
														assign node14950 = (inp[15]) ? 4'b0100 : 4'b0110;
												assign node14953 = (inp[4]) ? node14961 : node14954;
													assign node14954 = (inp[9]) ? node14958 : node14955;
														assign node14955 = (inp[15]) ? 4'b0110 : 4'b0100;
														assign node14958 = (inp[5]) ? 4'b0010 : 4'b0000;
													assign node14961 = (inp[9]) ? 4'b0110 : node14962;
														assign node14962 = (inp[3]) ? 4'b0000 : 4'b0010;
											assign node14966 = (inp[12]) ? node14980 : node14967;
												assign node14967 = (inp[3]) ? node14975 : node14968;
													assign node14968 = (inp[15]) ? node14972 : node14969;
														assign node14969 = (inp[4]) ? 4'b0110 : 4'b0100;
														assign node14972 = (inp[5]) ? 4'b0010 : 4'b0110;
													assign node14975 = (inp[5]) ? node14977 : 4'b0010;
														assign node14977 = (inp[9]) ? 4'b0010 : 4'b0010;
												assign node14980 = (inp[5]) ? node14988 : node14981;
													assign node14981 = (inp[9]) ? node14985 : node14982;
														assign node14982 = (inp[4]) ? 4'b0110 : 4'b0010;
														assign node14985 = (inp[4]) ? 4'b0010 : 4'b0100;
													assign node14988 = (inp[15]) ? 4'b0100 : 4'b0110;
								assign node14991 = (inp[14]) ? node15089 : node14992;
									assign node14992 = (inp[2]) ? node15048 : node14993;
										assign node14993 = (inp[4]) ? node15021 : node14994;
											assign node14994 = (inp[9]) ? node15008 : node14995;
												assign node14995 = (inp[12]) ? node15001 : node14996;
													assign node14996 = (inp[10]) ? 4'b0100 : node14997;
														assign node14997 = (inp[15]) ? 4'b0100 : 4'b0100;
													assign node15001 = (inp[10]) ? node15005 : node15002;
														assign node15002 = (inp[5]) ? 4'b0110 : 4'b0100;
														assign node15005 = (inp[15]) ? 4'b0010 : 4'b0000;
												assign node15008 = (inp[10]) ? node15016 : node15009;
													assign node15009 = (inp[15]) ? node15013 : node15010;
														assign node15010 = (inp[3]) ? 4'b0000 : 4'b0000;
														assign node15013 = (inp[3]) ? 4'b0000 : 4'b0010;
													assign node15016 = (inp[12]) ? node15018 : 4'b0000;
														assign node15018 = (inp[15]) ? 4'b0100 : 4'b0110;
											assign node15021 = (inp[9]) ? node15037 : node15022;
												assign node15022 = (inp[12]) ? node15030 : node15023;
													assign node15023 = (inp[15]) ? node15027 : node15024;
														assign node15024 = (inp[5]) ? 4'b0000 : 4'b0000;
														assign node15027 = (inp[3]) ? 4'b0000 : 4'b0010;
													assign node15030 = (inp[10]) ? node15034 : node15031;
														assign node15031 = (inp[5]) ? 4'b0000 : 4'b0010;
														assign node15034 = (inp[15]) ? 4'b0100 : 4'b0110;
												assign node15037 = (inp[12]) ? node15043 : node15038;
													assign node15038 = (inp[10]) ? 4'b0100 : node15039;
														assign node15039 = (inp[5]) ? 4'b0100 : 4'b0110;
													assign node15043 = (inp[10]) ? 4'b0010 : node15044;
														assign node15044 = (inp[15]) ? 4'b0110 : 4'b0100;
										assign node15048 = (inp[10]) ? node15072 : node15049;
											assign node15049 = (inp[15]) ? node15059 : node15050;
												assign node15050 = (inp[3]) ? node15054 : node15051;
													assign node15051 = (inp[12]) ? 4'b1001 : 4'b1101;
													assign node15054 = (inp[5]) ? node15056 : 4'b1111;
														assign node15056 = (inp[12]) ? 4'b1111 : 4'b1011;
												assign node15059 = (inp[3]) ? node15065 : node15060;
													assign node15060 = (inp[12]) ? node15062 : 4'b1111;
														assign node15062 = (inp[9]) ? 4'b1011 : 4'b1011;
													assign node15065 = (inp[12]) ? node15069 : node15066;
														assign node15066 = (inp[4]) ? 4'b1101 : 4'b1001;
														assign node15069 = (inp[5]) ? 4'b1101 : 4'b1001;
											assign node15072 = (inp[9]) ? node15082 : node15073;
												assign node15073 = (inp[4]) ? node15077 : node15074;
													assign node15074 = (inp[15]) ? 4'b1011 : 4'b1001;
													assign node15077 = (inp[5]) ? node15079 : 4'b1111;
														assign node15079 = (inp[15]) ? 4'b1101 : 4'b1111;
												assign node15082 = (inp[4]) ? node15084 : 4'b1101;
													assign node15084 = (inp[15]) ? 4'b1001 : node15085;
														assign node15085 = (inp[5]) ? 4'b1011 : 4'b1001;
									assign node15089 = (inp[10]) ? node15145 : node15090;
										assign node15090 = (inp[9]) ? node15122 : node15091;
											assign node15091 = (inp[15]) ? node15107 : node15092;
												assign node15092 = (inp[3]) ? node15100 : node15093;
													assign node15093 = (inp[4]) ? node15097 : node15094;
														assign node15094 = (inp[12]) ? 4'b1001 : 4'b1101;
														assign node15097 = (inp[12]) ? 4'b1101 : 4'b1001;
													assign node15100 = (inp[5]) ? node15104 : node15101;
														assign node15101 = (inp[12]) ? 4'b1001 : 4'b1001;
														assign node15104 = (inp[2]) ? 4'b1111 : 4'b1011;
												assign node15107 = (inp[3]) ? node15115 : node15108;
													assign node15108 = (inp[4]) ? node15112 : node15109;
														assign node15109 = (inp[12]) ? 4'b1011 : 4'b1111;
														assign node15112 = (inp[12]) ? 4'b1101 : 4'b1011;
													assign node15115 = (inp[5]) ? node15119 : node15116;
														assign node15116 = (inp[12]) ? 4'b1011 : 4'b1111;
														assign node15119 = (inp[2]) ? 4'b1001 : 4'b1001;
											assign node15122 = (inp[4]) ? node15132 : node15123;
												assign node15123 = (inp[12]) ? node15125 : 4'b1011;
													assign node15125 = (inp[15]) ? node15129 : node15126;
														assign node15126 = (inp[3]) ? 4'b1111 : 4'b1101;
														assign node15129 = (inp[5]) ? 4'b1101 : 4'b1111;
												assign node15132 = (inp[12]) ? node15138 : node15133;
													assign node15133 = (inp[15]) ? 4'b1101 : node15134;
														assign node15134 = (inp[3]) ? 4'b1111 : 4'b1101;
													assign node15138 = (inp[15]) ? node15142 : node15139;
														assign node15139 = (inp[3]) ? 4'b1011 : 4'b1001;
														assign node15142 = (inp[5]) ? 4'b1001 : 4'b1011;
										assign node15145 = (inp[12]) ? node15167 : node15146;
											assign node15146 = (inp[15]) ? node15158 : node15147;
												assign node15147 = (inp[3]) ? node15155 : node15148;
													assign node15148 = (inp[5]) ? node15152 : node15149;
														assign node15149 = (inp[4]) ? 4'b1101 : 4'b1101;
														assign node15152 = (inp[9]) ? 4'b1111 : 4'b1001;
													assign node15155 = (inp[4]) ? 4'b1011 : 4'b1111;
												assign node15158 = (inp[3]) ? node15162 : node15159;
													assign node15159 = (inp[5]) ? 4'b1001 : 4'b1011;
													assign node15162 = (inp[2]) ? node15164 : 4'b1101;
														assign node15164 = (inp[4]) ? 4'b1001 : 4'b1011;
											assign node15167 = (inp[4]) ? node15175 : node15168;
												assign node15168 = (inp[9]) ? 4'b1101 : node15169;
													assign node15169 = (inp[3]) ? 4'b1001 : node15170;
														assign node15170 = (inp[15]) ? 4'b1011 : 4'b1001;
												assign node15175 = (inp[9]) ? node15179 : node15176;
													assign node15176 = (inp[5]) ? 4'b1111 : 4'b1101;
													assign node15179 = (inp[5]) ? 4'b1001 : node15180;
														assign node15180 = (inp[3]) ? 4'b1001 : 4'b1001;
							assign node15184 = (inp[7]) ? node15356 : node15185;
								assign node15185 = (inp[2]) ? node15271 : node15186;
									assign node15186 = (inp[14]) ? node15226 : node15187;
										assign node15187 = (inp[4]) ? node15205 : node15188;
											assign node15188 = (inp[15]) ? node15196 : node15189;
												assign node15189 = (inp[9]) ? 4'b0000 : node15190;
													assign node15190 = (inp[12]) ? 4'b0000 : node15191;
														assign node15191 = (inp[5]) ? 4'b0110 : 4'b0100;
												assign node15196 = (inp[5]) ? node15202 : node15197;
													assign node15197 = (inp[9]) ? node15199 : 4'b0110;
														assign node15199 = (inp[12]) ? 4'b0000 : 4'b0010;
													assign node15202 = (inp[3]) ? 4'b0000 : 4'b0010;
											assign node15205 = (inp[9]) ? node15217 : node15206;
												assign node15206 = (inp[10]) ? node15212 : node15207;
													assign node15207 = (inp[12]) ? 4'b0000 : node15208;
														assign node15208 = (inp[3]) ? 4'b0010 : 4'b0000;
													assign node15212 = (inp[12]) ? node15214 : 4'b0000;
														assign node15214 = (inp[3]) ? 4'b0100 : 4'b0110;
												assign node15217 = (inp[12]) ? 4'b0000 : node15218;
													assign node15218 = (inp[10]) ? node15222 : node15219;
														assign node15219 = (inp[5]) ? 4'b0100 : 4'b0100;
														assign node15222 = (inp[5]) ? 4'b0100 : 4'b0110;
										assign node15226 = (inp[12]) ? node15244 : node15227;
											assign node15227 = (inp[15]) ? node15237 : node15228;
												assign node15228 = (inp[3]) ? node15232 : node15229;
													assign node15229 = (inp[10]) ? 4'b1001 : 4'b1101;
													assign node15232 = (inp[10]) ? node15234 : 4'b1001;
														assign node15234 = (inp[9]) ? 4'b1111 : 4'b1011;
												assign node15237 = (inp[3]) ? 4'b1011 : node15238;
													assign node15238 = (inp[9]) ? 4'b1111 : node15239;
														assign node15239 = (inp[10]) ? 4'b1011 : 4'b1111;
											assign node15244 = (inp[5]) ? node15258 : node15245;
												assign node15245 = (inp[15]) ? node15251 : node15246;
													assign node15246 = (inp[9]) ? 4'b1011 : node15247;
														assign node15247 = (inp[4]) ? 4'b1101 : 4'b1001;
													assign node15251 = (inp[3]) ? node15255 : node15252;
														assign node15252 = (inp[10]) ? 4'b1111 : 4'b1011;
														assign node15255 = (inp[4]) ? 4'b1001 : 4'b1011;
												assign node15258 = (inp[15]) ? node15266 : node15259;
													assign node15259 = (inp[9]) ? node15263 : node15260;
														assign node15260 = (inp[4]) ? 4'b1111 : 4'b1001;
														assign node15263 = (inp[4]) ? 4'b1011 : 4'b1111;
													assign node15266 = (inp[3]) ? 4'b1101 : node15267;
														assign node15267 = (inp[9]) ? 4'b1001 : 4'b1011;
									assign node15271 = (inp[15]) ? node15319 : node15272;
										assign node15272 = (inp[3]) ? node15296 : node15273;
											assign node15273 = (inp[5]) ? node15285 : node15274;
												assign node15274 = (inp[9]) ? node15280 : node15275;
													assign node15275 = (inp[12]) ? 4'b1001 : node15276;
														assign node15276 = (inp[4]) ? 4'b1001 : 4'b1101;
													assign node15280 = (inp[4]) ? node15282 : 4'b1101;
														assign node15282 = (inp[10]) ? 4'b1001 : 4'b1101;
												assign node15285 = (inp[14]) ? node15291 : node15286;
													assign node15286 = (inp[4]) ? node15288 : 4'b1111;
														assign node15288 = (inp[9]) ? 4'b1011 : 4'b1001;
													assign node15291 = (inp[12]) ? node15293 : 4'b1001;
														assign node15293 = (inp[10]) ? 4'b1001 : 4'b1111;
											assign node15296 = (inp[5]) ? node15308 : node15297;
												assign node15297 = (inp[4]) ? node15303 : node15298;
													assign node15298 = (inp[9]) ? 4'b1111 : node15299;
														assign node15299 = (inp[10]) ? 4'b1001 : 4'b1101;
													assign node15303 = (inp[9]) ? node15305 : 4'b1111;
														assign node15305 = (inp[12]) ? 4'b1011 : 4'b1111;
												assign node15308 = (inp[4]) ? node15316 : node15309;
													assign node15309 = (inp[9]) ? node15313 : node15310;
														assign node15310 = (inp[10]) ? 4'b1011 : 4'b1111;
														assign node15313 = (inp[12]) ? 4'b1111 : 4'b1011;
													assign node15316 = (inp[9]) ? 4'b1011 : 4'b1111;
										assign node15319 = (inp[4]) ? node15341 : node15320;
											assign node15320 = (inp[9]) ? node15330 : node15321;
												assign node15321 = (inp[12]) ? node15325 : node15322;
													assign node15322 = (inp[10]) ? 4'b1011 : 4'b1111;
													assign node15325 = (inp[14]) ? 4'b1011 : node15326;
														assign node15326 = (inp[3]) ? 4'b1001 : 4'b1011;
												assign node15330 = (inp[12]) ? node15336 : node15331;
													assign node15331 = (inp[10]) ? 4'b1101 : node15332;
														assign node15332 = (inp[14]) ? 4'b1001 : 4'b1011;
													assign node15336 = (inp[5]) ? 4'b1101 : node15337;
														assign node15337 = (inp[3]) ? 4'b1101 : 4'b1111;
											assign node15341 = (inp[9]) ? node15347 : node15342;
												assign node15342 = (inp[3]) ? 4'b1101 : node15343;
													assign node15343 = (inp[5]) ? 4'b1101 : 4'b1111;
												assign node15347 = (inp[10]) ? node15351 : node15348;
													assign node15348 = (inp[12]) ? 4'b1001 : 4'b1101;
													assign node15351 = (inp[14]) ? 4'b1001 : node15352;
														assign node15352 = (inp[5]) ? 4'b1001 : 4'b1011;
								assign node15356 = (inp[2]) ? node15440 : node15357;
									assign node15357 = (inp[14]) ? node15403 : node15358;
										assign node15358 = (inp[15]) ? node15382 : node15359;
											assign node15359 = (inp[3]) ? node15371 : node15360;
												assign node15360 = (inp[5]) ? node15366 : node15361;
													assign node15361 = (inp[10]) ? node15363 : 4'b1101;
														assign node15363 = (inp[12]) ? 4'b1001 : 4'b1001;
													assign node15366 = (inp[12]) ? 4'b1011 : node15367;
														assign node15367 = (inp[10]) ? 4'b1111 : 4'b1001;
												assign node15371 = (inp[4]) ? node15377 : node15372;
													assign node15372 = (inp[12]) ? 4'b1111 : node15373;
														assign node15373 = (inp[5]) ? 4'b1011 : 4'b1001;
													assign node15377 = (inp[9]) ? node15379 : 4'b1111;
														assign node15379 = (inp[12]) ? 4'b1011 : 4'b1111;
											assign node15382 = (inp[5]) ? node15394 : node15383;
												assign node15383 = (inp[3]) ? node15389 : node15384;
													assign node15384 = (inp[10]) ? 4'b1111 : node15385;
														assign node15385 = (inp[12]) ? 4'b1011 : 4'b1011;
													assign node15389 = (inp[9]) ? node15391 : 4'b1011;
														assign node15391 = (inp[4]) ? 4'b1001 : 4'b1101;
												assign node15394 = (inp[12]) ? node15400 : node15395;
													assign node15395 = (inp[10]) ? node15397 : 4'b1001;
														assign node15397 = (inp[4]) ? 4'b1101 : 4'b1001;
													assign node15400 = (inp[10]) ? 4'b1001 : 4'b1101;
										assign node15403 = (inp[4]) ? node15429 : node15404;
											assign node15404 = (inp[9]) ? node15418 : node15405;
												assign node15405 = (inp[15]) ? node15411 : node15406;
													assign node15406 = (inp[10]) ? 4'b1000 : node15407;
														assign node15407 = (inp[5]) ? 4'b1010 : 4'b1000;
													assign node15411 = (inp[12]) ? node15415 : node15412;
														assign node15412 = (inp[3]) ? 4'b1010 : 4'b1110;
														assign node15415 = (inp[5]) ? 4'b1000 : 4'b1010;
												assign node15418 = (inp[15]) ? node15424 : node15419;
													assign node15419 = (inp[3]) ? 4'b1110 : node15420;
														assign node15420 = (inp[5]) ? 4'b1110 : 4'b1100;
													assign node15424 = (inp[3]) ? node15426 : 4'b1110;
														assign node15426 = (inp[10]) ? 4'b1100 : 4'b1000;
											assign node15429 = (inp[9]) ? node15437 : node15430;
												assign node15430 = (inp[15]) ? node15432 : 4'b1110;
													assign node15432 = (inp[3]) ? 4'b1100 : node15433;
														assign node15433 = (inp[12]) ? 4'b1110 : 4'b1100;
												assign node15437 = (inp[10]) ? 4'b1010 : 4'b1100;
									assign node15440 = (inp[15]) ? node15476 : node15441;
										assign node15441 = (inp[3]) ? node15459 : node15442;
											assign node15442 = (inp[9]) ? node15450 : node15443;
												assign node15443 = (inp[4]) ? node15447 : node15444;
													assign node15444 = (inp[10]) ? 4'b1000 : 4'b1100;
													assign node15447 = (inp[5]) ? 4'b1000 : 4'b1100;
												assign node15450 = (inp[5]) ? node15456 : node15451;
													assign node15451 = (inp[4]) ? 4'b1000 : node15452;
														assign node15452 = (inp[12]) ? 4'b1100 : 4'b1000;
													assign node15456 = (inp[4]) ? 4'b1010 : 4'b1110;
											assign node15459 = (inp[4]) ? node15467 : node15460;
												assign node15460 = (inp[9]) ? 4'b1110 : node15461;
													assign node15461 = (inp[14]) ? 4'b1110 : node15462;
														assign node15462 = (inp[5]) ? 4'b1010 : 4'b1000;
												assign node15467 = (inp[9]) ? node15471 : node15468;
													assign node15468 = (inp[10]) ? 4'b1110 : 4'b1000;
													assign node15471 = (inp[10]) ? 4'b1010 : node15472;
														assign node15472 = (inp[12]) ? 4'b1010 : 4'b1110;
										assign node15476 = (inp[3]) ? node15500 : node15477;
											assign node15477 = (inp[5]) ? node15487 : node15478;
												assign node15478 = (inp[9]) ? node15482 : node15479;
													assign node15479 = (inp[4]) ? 4'b1110 : 4'b1010;
													assign node15482 = (inp[14]) ? 4'b1110 : node15483;
														assign node15483 = (inp[4]) ? 4'b1010 : 4'b1010;
												assign node15487 = (inp[9]) ? node15493 : node15488;
													assign node15488 = (inp[4]) ? 4'b1100 : node15489;
														assign node15489 = (inp[10]) ? 4'b1010 : 4'b1110;
													assign node15493 = (inp[12]) ? node15497 : node15494;
														assign node15494 = (inp[4]) ? 4'b1100 : 4'b1010;
														assign node15497 = (inp[4]) ? 4'b1000 : 4'b1100;
											assign node15500 = (inp[5]) ? node15506 : node15501;
												assign node15501 = (inp[14]) ? node15503 : 4'b1100;
													assign node15503 = (inp[4]) ? 4'b1000 : 4'b1010;
												assign node15506 = (inp[12]) ? node15512 : node15507;
													assign node15507 = (inp[4]) ? 4'b1100 : node15508;
														assign node15508 = (inp[9]) ? 4'b1000 : 4'b1100;
													assign node15512 = (inp[14]) ? node15514 : 4'b1000;
														assign node15514 = (inp[10]) ? 4'b1100 : 4'b1000;
					assign node15517 = (inp[13]) ? node16253 : node15518;
						assign node15518 = (inp[7]) ? node15882 : node15519;
							assign node15519 = (inp[8]) ? node15697 : node15520;
								assign node15520 = (inp[14]) ? node15596 : node15521;
									assign node15521 = (inp[2]) ? node15561 : node15522;
										assign node15522 = (inp[15]) ? node15540 : node15523;
											assign node15523 = (inp[5]) ? node15535 : node15524;
												assign node15524 = (inp[9]) ? node15530 : node15525;
													assign node15525 = (inp[4]) ? 4'b0001 : node15526;
														assign node15526 = (inp[12]) ? 4'b0001 : 4'b0101;
													assign node15530 = (inp[3]) ? 4'b0111 : node15531;
														assign node15531 = (inp[10]) ? 4'b0101 : 4'b0001;
												assign node15535 = (inp[3]) ? 4'b0111 : node15536;
													assign node15536 = (inp[9]) ? 4'b0111 : 4'b0001;
											assign node15540 = (inp[3]) ? node15548 : node15541;
												assign node15541 = (inp[12]) ? node15543 : 4'b0011;
													assign node15543 = (inp[9]) ? 4'b0001 : node15544;
														assign node15544 = (inp[5]) ? 4'b0101 : 4'b0111;
												assign node15548 = (inp[9]) ? node15554 : node15549;
													assign node15549 = (inp[5]) ? node15551 : 4'b0011;
														assign node15551 = (inp[4]) ? 4'b0001 : 4'b0101;
													assign node15554 = (inp[5]) ? node15558 : node15555;
														assign node15555 = (inp[10]) ? 4'b0101 : 4'b0101;
														assign node15558 = (inp[4]) ? 4'b0101 : 4'b0001;
										assign node15561 = (inp[4]) ? node15573 : node15562;
											assign node15562 = (inp[9]) ? node15568 : node15563;
												assign node15563 = (inp[15]) ? node15565 : 4'b0100;
													assign node15565 = (inp[5]) ? 4'b0100 : 4'b0110;
												assign node15568 = (inp[12]) ? node15570 : 4'b0010;
													assign node15570 = (inp[10]) ? 4'b0100 : 4'b0000;
											assign node15573 = (inp[9]) ? node15585 : node15574;
												assign node15574 = (inp[10]) ? node15582 : node15575;
													assign node15575 = (inp[15]) ? node15579 : node15576;
														assign node15576 = (inp[3]) ? 4'b0010 : 4'b0000;
														assign node15579 = (inp[5]) ? 4'b0000 : 4'b0010;
													assign node15582 = (inp[12]) ? 4'b0110 : 4'b0010;
												assign node15585 = (inp[10]) ? node15591 : node15586;
													assign node15586 = (inp[15]) ? node15588 : 4'b0110;
														assign node15588 = (inp[3]) ? 4'b0100 : 4'b0110;
													assign node15591 = (inp[15]) ? 4'b0100 : node15592;
														assign node15592 = (inp[5]) ? 4'b0010 : 4'b0000;
									assign node15596 = (inp[12]) ? node15644 : node15597;
										assign node15597 = (inp[10]) ? node15619 : node15598;
											assign node15598 = (inp[15]) ? node15610 : node15599;
												assign node15599 = (inp[4]) ? node15603 : node15600;
													assign node15600 = (inp[9]) ? 4'b0000 : 4'b0100;
													assign node15603 = (inp[9]) ? node15607 : node15604;
														assign node15604 = (inp[2]) ? 4'b0000 : 4'b0000;
														assign node15607 = (inp[3]) ? 4'b0110 : 4'b0100;
												assign node15610 = (inp[4]) ? node15616 : node15611;
													assign node15611 = (inp[9]) ? node15613 : 4'b0110;
														assign node15613 = (inp[3]) ? 4'b0000 : 4'b0010;
													assign node15616 = (inp[9]) ? 4'b0100 : 4'b0000;
											assign node15619 = (inp[2]) ? node15629 : node15620;
												assign node15620 = (inp[5]) ? node15624 : node15621;
													assign node15621 = (inp[9]) ? 4'b0100 : 4'b0000;
													assign node15624 = (inp[9]) ? 4'b0110 : node15625;
														assign node15625 = (inp[3]) ? 4'b0100 : 4'b0100;
												assign node15629 = (inp[3]) ? node15637 : node15630;
													assign node15630 = (inp[5]) ? node15634 : node15631;
														assign node15631 = (inp[9]) ? 4'b0110 : 4'b0010;
														assign node15634 = (inp[9]) ? 4'b0010 : 4'b0110;
													assign node15637 = (inp[15]) ? node15641 : node15638;
														assign node15638 = (inp[4]) ? 4'b0110 : 4'b0010;
														assign node15641 = (inp[5]) ? 4'b0000 : 4'b0010;
										assign node15644 = (inp[15]) ? node15670 : node15645;
											assign node15645 = (inp[5]) ? node15657 : node15646;
												assign node15646 = (inp[9]) ? node15652 : node15647;
													assign node15647 = (inp[2]) ? node15649 : 4'b0100;
														assign node15649 = (inp[10]) ? 4'b0100 : 4'b0000;
													assign node15652 = (inp[3]) ? node15654 : 4'b0000;
														assign node15654 = (inp[4]) ? 4'b0110 : 4'b0000;
												assign node15657 = (inp[9]) ? node15663 : node15658;
													assign node15658 = (inp[3]) ? node15660 : 4'b0000;
														assign node15660 = (inp[2]) ? 4'b0010 : 4'b0010;
													assign node15663 = (inp[10]) ? node15667 : node15664;
														assign node15664 = (inp[4]) ? 4'b0110 : 4'b0010;
														assign node15667 = (inp[4]) ? 4'b0010 : 4'b0110;
											assign node15670 = (inp[9]) ? node15684 : node15671;
												assign node15671 = (inp[5]) ? node15677 : node15672;
													assign node15672 = (inp[3]) ? 4'b0010 : node15673;
														assign node15673 = (inp[4]) ? 4'b0010 : 4'b0110;
													assign node15677 = (inp[4]) ? node15681 : node15678;
														assign node15678 = (inp[10]) ? 4'b0010 : 4'b0110;
														assign node15681 = (inp[10]) ? 4'b0100 : 4'b0000;
												assign node15684 = (inp[3]) ? node15690 : node15685;
													assign node15685 = (inp[4]) ? 4'b0100 : node15686;
														assign node15686 = (inp[5]) ? 4'b0010 : 4'b0110;
													assign node15690 = (inp[5]) ? node15694 : node15691;
														assign node15691 = (inp[4]) ? 4'b0000 : 4'b0100;
														assign node15694 = (inp[2]) ? 4'b0000 : 4'b0000;
								assign node15697 = (inp[14]) ? node15781 : node15698;
									assign node15698 = (inp[2]) ? node15742 : node15699;
										assign node15699 = (inp[15]) ? node15719 : node15700;
											assign node15700 = (inp[5]) ? node15710 : node15701;
												assign node15701 = (inp[9]) ? node15707 : node15702;
													assign node15702 = (inp[4]) ? 4'b0000 : node15703;
														assign node15703 = (inp[10]) ? 4'b0000 : 4'b0100;
													assign node15707 = (inp[4]) ? 4'b0100 : 4'b0000;
												assign node15710 = (inp[12]) ? node15712 : 4'b0000;
													assign node15712 = (inp[4]) ? node15716 : node15713;
														assign node15713 = (inp[3]) ? 4'b0010 : 4'b0110;
														assign node15716 = (inp[10]) ? 4'b0010 : 4'b0000;
											assign node15719 = (inp[3]) ? node15731 : node15720;
												assign node15720 = (inp[9]) ? node15726 : node15721;
													assign node15721 = (inp[4]) ? 4'b0010 : node15722;
														assign node15722 = (inp[10]) ? 4'b0110 : 4'b0110;
													assign node15726 = (inp[4]) ? node15728 : 4'b0010;
														assign node15728 = (inp[5]) ? 4'b0100 : 4'b0110;
												assign node15731 = (inp[12]) ? node15737 : node15732;
													assign node15732 = (inp[9]) ? 4'b0010 : node15733;
														assign node15733 = (inp[4]) ? 4'b0010 : 4'b0110;
													assign node15737 = (inp[9]) ? node15739 : 4'b0000;
														assign node15739 = (inp[10]) ? 4'b0100 : 4'b0000;
										assign node15742 = (inp[15]) ? node15764 : node15743;
											assign node15743 = (inp[3]) ? node15755 : node15744;
												assign node15744 = (inp[5]) ? node15750 : node15745;
													assign node15745 = (inp[4]) ? node15747 : 4'b1101;
														assign node15747 = (inp[10]) ? 4'b1001 : 4'b1101;
													assign node15750 = (inp[9]) ? node15752 : 4'b1001;
														assign node15752 = (inp[4]) ? 4'b1011 : 4'b1111;
												assign node15755 = (inp[5]) ? node15757 : 4'b1111;
													assign node15757 = (inp[12]) ? node15761 : node15758;
														assign node15758 = (inp[9]) ? 4'b1111 : 4'b1011;
														assign node15761 = (inp[9]) ? 4'b1011 : 4'b1111;
											assign node15764 = (inp[5]) ? node15774 : node15765;
												assign node15765 = (inp[9]) ? node15769 : node15766;
													assign node15766 = (inp[4]) ? 4'b1111 : 4'b1011;
													assign node15769 = (inp[3]) ? node15771 : 4'b1011;
														assign node15771 = (inp[12]) ? 4'b1001 : 4'b1101;
												assign node15774 = (inp[4]) ? 4'b1101 : node15775;
													assign node15775 = (inp[3]) ? node15777 : 4'b1011;
														assign node15777 = (inp[9]) ? 4'b1101 : 4'b1001;
									assign node15781 = (inp[10]) ? node15835 : node15782;
										assign node15782 = (inp[15]) ? node15810 : node15783;
											assign node15783 = (inp[3]) ? node15795 : node15784;
												assign node15784 = (inp[4]) ? node15790 : node15785;
													assign node15785 = (inp[9]) ? 4'b1001 : node15786;
														assign node15786 = (inp[2]) ? 4'b1101 : 4'b1001;
													assign node15790 = (inp[5]) ? 4'b1111 : node15791;
														assign node15791 = (inp[9]) ? 4'b1001 : 4'b1101;
												assign node15795 = (inp[5]) ? node15803 : node15796;
													assign node15796 = (inp[12]) ? node15800 : node15797;
														assign node15797 = (inp[9]) ? 4'b1111 : 4'b1001;
														assign node15800 = (inp[9]) ? 4'b1011 : 4'b1111;
													assign node15803 = (inp[2]) ? node15807 : node15804;
														assign node15804 = (inp[12]) ? 4'b1011 : 4'b1111;
														assign node15807 = (inp[9]) ? 4'b1011 : 4'b1011;
											assign node15810 = (inp[3]) ? node15824 : node15811;
												assign node15811 = (inp[5]) ? node15817 : node15812;
													assign node15812 = (inp[9]) ? 4'b1111 : node15813;
														assign node15813 = (inp[2]) ? 4'b1011 : 4'b1111;
													assign node15817 = (inp[12]) ? node15821 : node15818;
														assign node15818 = (inp[2]) ? 4'b1011 : 4'b1011;
														assign node15821 = (inp[9]) ? 4'b1001 : 4'b1011;
												assign node15824 = (inp[5]) ? node15830 : node15825;
													assign node15825 = (inp[9]) ? node15827 : 4'b1011;
														assign node15827 = (inp[12]) ? 4'b1001 : 4'b1101;
													assign node15830 = (inp[9]) ? 4'b1101 : node15831;
														assign node15831 = (inp[12]) ? 4'b1001 : 4'b1001;
										assign node15835 = (inp[15]) ? node15865 : node15836;
											assign node15836 = (inp[5]) ? node15852 : node15837;
												assign node15837 = (inp[3]) ? node15845 : node15838;
													assign node15838 = (inp[4]) ? node15842 : node15839;
														assign node15839 = (inp[9]) ? 4'b1101 : 4'b1001;
														assign node15842 = (inp[9]) ? 4'b1001 : 4'b1101;
													assign node15845 = (inp[4]) ? node15849 : node15846;
														assign node15846 = (inp[9]) ? 4'b1111 : 4'b1001;
														assign node15849 = (inp[9]) ? 4'b1011 : 4'b1111;
												assign node15852 = (inp[2]) ? node15860 : node15853;
													assign node15853 = (inp[4]) ? node15857 : node15854;
														assign node15854 = (inp[9]) ? 4'b1111 : 4'b1001;
														assign node15857 = (inp[9]) ? 4'b1011 : 4'b1111;
													assign node15860 = (inp[3]) ? node15862 : 4'b1111;
														assign node15862 = (inp[4]) ? 4'b1111 : 4'b1011;
											assign node15865 = (inp[2]) ? node15873 : node15866;
												assign node15866 = (inp[5]) ? node15868 : 4'b1101;
													assign node15868 = (inp[3]) ? node15870 : 4'b1101;
														assign node15870 = (inp[12]) ? 4'b1001 : 4'b1001;
												assign node15873 = (inp[9]) ? node15879 : node15874;
													assign node15874 = (inp[4]) ? 4'b1101 : node15875;
														assign node15875 = (inp[3]) ? 4'b1001 : 4'b1011;
													assign node15879 = (inp[4]) ? 4'b1001 : 4'b1101;
							assign node15882 = (inp[8]) ? node16066 : node15883;
								assign node15883 = (inp[2]) ? node15981 : node15884;
									assign node15884 = (inp[14]) ? node15930 : node15885;
										assign node15885 = (inp[12]) ? node15909 : node15886;
											assign node15886 = (inp[3]) ? node15898 : node15887;
												assign node15887 = (inp[15]) ? node15893 : node15888;
													assign node15888 = (inp[10]) ? 4'b0000 : node15889;
														assign node15889 = (inp[4]) ? 4'b0000 : 4'b0100;
													assign node15893 = (inp[5]) ? node15895 : 4'b0010;
														assign node15895 = (inp[10]) ? 4'b0010 : 4'b0110;
												assign node15898 = (inp[4]) ? node15902 : node15899;
													assign node15899 = (inp[9]) ? 4'b0000 : 4'b0100;
													assign node15902 = (inp[9]) ? node15906 : node15903;
														assign node15903 = (inp[15]) ? 4'b0010 : 4'b0000;
														assign node15906 = (inp[15]) ? 4'b0100 : 4'b0110;
											assign node15909 = (inp[15]) ? node15921 : node15910;
												assign node15910 = (inp[5]) ? node15916 : node15911;
													assign node15911 = (inp[9]) ? node15913 : 4'b0100;
														assign node15913 = (inp[10]) ? 4'b0000 : 4'b0110;
													assign node15916 = (inp[10]) ? 4'b0110 : node15917;
														assign node15917 = (inp[4]) ? 4'b0010 : 4'b0010;
												assign node15921 = (inp[10]) ? node15927 : node15922;
													assign node15922 = (inp[5]) ? 4'b0100 : node15923;
														assign node15923 = (inp[9]) ? 4'b0110 : 4'b0010;
													assign node15927 = (inp[9]) ? 4'b0000 : 4'b0100;
										assign node15930 = (inp[15]) ? node15956 : node15931;
											assign node15931 = (inp[3]) ? node15943 : node15932;
												assign node15932 = (inp[4]) ? node15940 : node15933;
													assign node15933 = (inp[9]) ? node15937 : node15934;
														assign node15934 = (inp[10]) ? 4'b1001 : 4'b1101;
														assign node15937 = (inp[10]) ? 4'b1111 : 4'b1101;
													assign node15940 = (inp[5]) ? 4'b1111 : 4'b1101;
												assign node15943 = (inp[4]) ? node15949 : node15944;
													assign node15944 = (inp[12]) ? 4'b1111 : node15945;
														assign node15945 = (inp[9]) ? 4'b1011 : 4'b1011;
													assign node15949 = (inp[9]) ? node15953 : node15950;
														assign node15950 = (inp[12]) ? 4'b1111 : 4'b1011;
														assign node15953 = (inp[10]) ? 4'b1011 : 4'b1011;
											assign node15956 = (inp[3]) ? node15970 : node15957;
												assign node15957 = (inp[5]) ? node15963 : node15958;
													assign node15958 = (inp[12]) ? 4'b1011 : node15959;
														assign node15959 = (inp[10]) ? 4'b1011 : 4'b1111;
													assign node15963 = (inp[4]) ? node15967 : node15964;
														assign node15964 = (inp[9]) ? 4'b1001 : 4'b1011;
														assign node15967 = (inp[9]) ? 4'b1001 : 4'b1101;
												assign node15970 = (inp[10]) ? node15976 : node15971;
													assign node15971 = (inp[5]) ? node15973 : 4'b1101;
														assign node15973 = (inp[12]) ? 4'b1001 : 4'b1001;
													assign node15976 = (inp[9]) ? 4'b1001 : node15977;
														assign node15977 = (inp[5]) ? 4'b1001 : 4'b1101;
									assign node15981 = (inp[15]) ? node16027 : node15982;
										assign node15982 = (inp[5]) ? node16004 : node15983;
											assign node15983 = (inp[3]) ? node15993 : node15984;
												assign node15984 = (inp[12]) ? node15988 : node15985;
													assign node15985 = (inp[9]) ? 4'b1001 : 4'b1101;
													assign node15988 = (inp[4]) ? 4'b1101 : node15989;
														assign node15989 = (inp[10]) ? 4'b1101 : 4'b1001;
												assign node15993 = (inp[4]) ? node16001 : node15994;
													assign node15994 = (inp[9]) ? node15998 : node15995;
														assign node15995 = (inp[12]) ? 4'b1001 : 4'b1001;
														assign node15998 = (inp[10]) ? 4'b1111 : 4'b1001;
													assign node16001 = (inp[9]) ? 4'b1011 : 4'b1111;
											assign node16004 = (inp[3]) ? node16016 : node16005;
												assign node16005 = (inp[4]) ? node16011 : node16006;
													assign node16006 = (inp[14]) ? 4'b1001 : node16007;
														assign node16007 = (inp[10]) ? 4'b1111 : 4'b1001;
													assign node16011 = (inp[10]) ? 4'b1011 : node16012;
														assign node16012 = (inp[14]) ? 4'b1111 : 4'b1011;
												assign node16016 = (inp[10]) ? node16022 : node16017;
													assign node16017 = (inp[4]) ? 4'b1111 : node16018;
														assign node16018 = (inp[14]) ? 4'b1111 : 4'b1011;
													assign node16022 = (inp[4]) ? node16024 : 4'b1011;
														assign node16024 = (inp[9]) ? 4'b1011 : 4'b1111;
										assign node16027 = (inp[3]) ? node16045 : node16028;
											assign node16028 = (inp[5]) ? node16036 : node16029;
												assign node16029 = (inp[12]) ? node16031 : 4'b1111;
													assign node16031 = (inp[14]) ? node16033 : 4'b1011;
														assign node16033 = (inp[10]) ? 4'b1011 : 4'b1111;
												assign node16036 = (inp[9]) ? node16042 : node16037;
													assign node16037 = (inp[4]) ? 4'b1101 : node16038;
														assign node16038 = (inp[12]) ? 4'b1011 : 4'b1111;
													assign node16042 = (inp[12]) ? 4'b1001 : 4'b1101;
											assign node16045 = (inp[4]) ? node16059 : node16046;
												assign node16046 = (inp[5]) ? node16054 : node16047;
													assign node16047 = (inp[9]) ? node16051 : node16048;
														assign node16048 = (inp[10]) ? 4'b1011 : 4'b1111;
														assign node16051 = (inp[14]) ? 4'b1101 : 4'b1001;
													assign node16054 = (inp[14]) ? 4'b1101 : node16055;
														assign node16055 = (inp[12]) ? 4'b1101 : 4'b1001;
												assign node16059 = (inp[9]) ? 4'b1001 : node16060;
													assign node16060 = (inp[14]) ? 4'b1101 : node16061;
														assign node16061 = (inp[12]) ? 4'b1101 : 4'b1001;
								assign node16066 = (inp[2]) ? node16166 : node16067;
									assign node16067 = (inp[14]) ? node16121 : node16068;
										assign node16068 = (inp[3]) ? node16096 : node16069;
											assign node16069 = (inp[10]) ? node16083 : node16070;
												assign node16070 = (inp[15]) ? node16078 : node16071;
													assign node16071 = (inp[12]) ? node16075 : node16072;
														assign node16072 = (inp[4]) ? 4'b1001 : 4'b1001;
														assign node16075 = (inp[9]) ? 4'b1011 : 4'b1001;
													assign node16078 = (inp[9]) ? node16080 : 4'b1011;
														assign node16080 = (inp[4]) ? 4'b1001 : 4'b1111;
												assign node16083 = (inp[5]) ? node16089 : node16084;
													assign node16084 = (inp[9]) ? 4'b1011 : node16085;
														assign node16085 = (inp[4]) ? 4'b1111 : 4'b1011;
													assign node16089 = (inp[15]) ? node16093 : node16090;
														assign node16090 = (inp[4]) ? 4'b1011 : 4'b1001;
														assign node16093 = (inp[9]) ? 4'b1001 : 4'b1011;
											assign node16096 = (inp[15]) ? node16108 : node16097;
												assign node16097 = (inp[12]) ? node16103 : node16098;
													assign node16098 = (inp[5]) ? node16100 : 4'b1111;
														assign node16100 = (inp[4]) ? 4'b1011 : 4'b1111;
													assign node16103 = (inp[4]) ? node16105 : 4'b1001;
														assign node16105 = (inp[9]) ? 4'b1011 : 4'b1111;
												assign node16108 = (inp[12]) ? node16116 : node16109;
													assign node16109 = (inp[9]) ? node16113 : node16110;
														assign node16110 = (inp[4]) ? 4'b1001 : 4'b1011;
														assign node16113 = (inp[4]) ? 4'b1001 : 4'b1101;
													assign node16116 = (inp[9]) ? 4'b1101 : node16117;
														assign node16117 = (inp[4]) ? 4'b1101 : 4'b1011;
										assign node16121 = (inp[5]) ? node16145 : node16122;
											assign node16122 = (inp[9]) ? node16130 : node16123;
												assign node16123 = (inp[4]) ? node16127 : node16124;
													assign node16124 = (inp[15]) ? 4'b1010 : 4'b1000;
													assign node16127 = (inp[10]) ? 4'b1110 : 4'b1010;
												assign node16130 = (inp[4]) ? node16138 : node16131;
													assign node16131 = (inp[10]) ? node16135 : node16132;
														assign node16132 = (inp[12]) ? 4'b1100 : 4'b1010;
														assign node16135 = (inp[15]) ? 4'b1100 : 4'b1100;
													assign node16138 = (inp[10]) ? node16142 : node16139;
														assign node16139 = (inp[12]) ? 4'b1010 : 4'b1110;
														assign node16142 = (inp[12]) ? 4'b1010 : 4'b1000;
											assign node16145 = (inp[15]) ? node16155 : node16146;
												assign node16146 = (inp[4]) ? node16152 : node16147;
													assign node16147 = (inp[3]) ? 4'b1010 : node16148;
														assign node16148 = (inp[10]) ? 4'b1000 : 4'b1000;
													assign node16152 = (inp[9]) ? 4'b1010 : 4'b1110;
												assign node16155 = (inp[3]) ? node16159 : node16156;
													assign node16156 = (inp[12]) ? 4'b1000 : 4'b1100;
													assign node16159 = (inp[9]) ? node16163 : node16160;
														assign node16160 = (inp[12]) ? 4'b1100 : 4'b1000;
														assign node16163 = (inp[4]) ? 4'b1000 : 4'b1100;
									assign node16166 = (inp[15]) ? node16210 : node16167;
										assign node16167 = (inp[3]) ? node16191 : node16168;
											assign node16168 = (inp[5]) ? node16180 : node16169;
												assign node16169 = (inp[12]) ? node16175 : node16170;
													assign node16170 = (inp[9]) ? 4'b1000 : node16171;
														assign node16171 = (inp[4]) ? 4'b1000 : 4'b1000;
													assign node16175 = (inp[14]) ? node16177 : 4'b1100;
														assign node16177 = (inp[10]) ? 4'b1100 : 4'b1000;
												assign node16180 = (inp[4]) ? node16188 : node16181;
													assign node16181 = (inp[9]) ? node16185 : node16182;
														assign node16182 = (inp[12]) ? 4'b1000 : 4'b1100;
														assign node16185 = (inp[14]) ? 4'b1000 : 4'b1110;
													assign node16188 = (inp[12]) ? 4'b1110 : 4'b1010;
											assign node16191 = (inp[9]) ? node16201 : node16192;
												assign node16192 = (inp[4]) ? node16196 : node16193;
													assign node16193 = (inp[5]) ? 4'b1010 : 4'b1000;
													assign node16196 = (inp[10]) ? 4'b1110 : node16197;
														assign node16197 = (inp[12]) ? 4'b1110 : 4'b1010;
												assign node16201 = (inp[4]) ? node16207 : node16202;
													assign node16202 = (inp[12]) ? 4'b1110 : node16203;
														assign node16203 = (inp[10]) ? 4'b1110 : 4'b1010;
													assign node16207 = (inp[10]) ? 4'b1010 : 4'b1110;
										assign node16210 = (inp[3]) ? node16232 : node16211;
											assign node16211 = (inp[5]) ? node16223 : node16212;
												assign node16212 = (inp[10]) ? node16218 : node16213;
													assign node16213 = (inp[4]) ? 4'b1110 : node16214;
														assign node16214 = (inp[9]) ? 4'b1010 : 4'b1110;
													assign node16218 = (inp[14]) ? node16220 : 4'b1010;
														assign node16220 = (inp[9]) ? 4'b1010 : 4'b1110;
												assign node16223 = (inp[4]) ? node16229 : node16224;
													assign node16224 = (inp[9]) ? node16226 : 4'b1010;
														assign node16226 = (inp[10]) ? 4'b1100 : 4'b1010;
													assign node16229 = (inp[9]) ? 4'b1000 : 4'b1100;
											assign node16232 = (inp[4]) ? node16242 : node16233;
												assign node16233 = (inp[9]) ? node16237 : node16234;
													assign node16234 = (inp[5]) ? 4'b1000 : 4'b1010;
													assign node16237 = (inp[12]) ? 4'b1100 : node16238;
														assign node16238 = (inp[10]) ? 4'b1100 : 4'b1000;
												assign node16242 = (inp[9]) ? node16248 : node16243;
													assign node16243 = (inp[12]) ? 4'b1100 : node16244;
														assign node16244 = (inp[10]) ? 4'b1100 : 4'b1000;
													assign node16248 = (inp[12]) ? 4'b1000 : node16249;
														assign node16249 = (inp[14]) ? 4'b1000 : 4'b1100;
						assign node16253 = (inp[15]) ? node16623 : node16254;
							assign node16254 = (inp[5]) ? node16432 : node16255;
								assign node16255 = (inp[3]) ? node16353 : node16256;
									assign node16256 = (inp[12]) ? node16302 : node16257;
										assign node16257 = (inp[7]) ? node16279 : node16258;
											assign node16258 = (inp[8]) ? node16268 : node16259;
												assign node16259 = (inp[14]) ? node16265 : node16260;
													assign node16260 = (inp[2]) ? 4'b1100 : node16261;
														assign node16261 = (inp[10]) ? 4'b1101 : 4'b1001;
													assign node16265 = (inp[4]) ? 4'b1000 : 4'b1100;
												assign node16268 = (inp[2]) ? node16272 : node16269;
													assign node16269 = (inp[14]) ? 4'b1101 : 4'b1100;
													assign node16272 = (inp[9]) ? node16276 : node16273;
														assign node16273 = (inp[4]) ? 4'b1001 : 4'b1001;
														assign node16276 = (inp[4]) ? 4'b1001 : 4'b1101;
											assign node16279 = (inp[8]) ? node16295 : node16280;
												assign node16280 = (inp[10]) ? node16288 : node16281;
													assign node16281 = (inp[14]) ? node16285 : node16282;
														assign node16282 = (inp[9]) ? 4'b1001 : 4'b1001;
														assign node16285 = (inp[9]) ? 4'b1101 : 4'b1001;
													assign node16288 = (inp[2]) ? node16292 : node16289;
														assign node16289 = (inp[4]) ? 4'b1000 : 4'b1001;
														assign node16292 = (inp[4]) ? 4'b1001 : 4'b1001;
												assign node16295 = (inp[2]) ? 4'b1000 : node16296;
													assign node16296 = (inp[14]) ? node16298 : 4'b1101;
														assign node16298 = (inp[9]) ? 4'b1000 : 4'b1000;
										assign node16302 = (inp[10]) ? node16328 : node16303;
											assign node16303 = (inp[2]) ? node16319 : node16304;
												assign node16304 = (inp[7]) ? node16312 : node16305;
													assign node16305 = (inp[9]) ? node16309 : node16306;
														assign node16306 = (inp[4]) ? 4'b1101 : 4'b1000;
														assign node16309 = (inp[4]) ? 4'b1000 : 4'b1100;
													assign node16312 = (inp[8]) ? node16316 : node16313;
														assign node16313 = (inp[9]) ? 4'b1000 : 4'b1000;
														assign node16316 = (inp[9]) ? 4'b1101 : 4'b1100;
												assign node16319 = (inp[9]) ? node16325 : node16320;
													assign node16320 = (inp[14]) ? 4'b1000 : node16321;
														assign node16321 = (inp[8]) ? 4'b1000 : 4'b1000;
													assign node16325 = (inp[4]) ? 4'b1000 : 4'b1100;
											assign node16328 = (inp[7]) ? node16344 : node16329;
												assign node16329 = (inp[8]) ? node16337 : node16330;
													assign node16330 = (inp[14]) ? node16334 : node16331;
														assign node16331 = (inp[2]) ? 4'b1000 : 4'b1001;
														assign node16334 = (inp[4]) ? 4'b1000 : 4'b1000;
													assign node16337 = (inp[2]) ? node16341 : node16338;
														assign node16338 = (inp[14]) ? 4'b1101 : 4'b1000;
														assign node16341 = (inp[4]) ? 4'b1101 : 4'b1001;
												assign node16344 = (inp[8]) ? node16348 : node16345;
													assign node16345 = (inp[14]) ? 4'b1101 : 4'b1001;
													assign node16348 = (inp[14]) ? node16350 : 4'b1101;
														assign node16350 = (inp[9]) ? 4'b1100 : 4'b1000;
									assign node16353 = (inp[9]) ? node16395 : node16354;
										assign node16354 = (inp[4]) ? node16376 : node16355;
											assign node16355 = (inp[10]) ? node16365 : node16356;
												assign node16356 = (inp[12]) ? 4'b1001 : node16357;
													assign node16357 = (inp[2]) ? node16361 : node16358;
														assign node16358 = (inp[14]) ? 4'b1101 : 4'b1100;
														assign node16361 = (inp[14]) ? 4'b1100 : 4'b1101;
												assign node16365 = (inp[8]) ? node16371 : node16366;
													assign node16366 = (inp[12]) ? node16368 : 4'b1001;
														assign node16368 = (inp[14]) ? 4'b1001 : 4'b1000;
													assign node16371 = (inp[14]) ? 4'b1000 : node16372;
														assign node16372 = (inp[12]) ? 4'b1000 : 4'b1000;
											assign node16376 = (inp[12]) ? node16388 : node16377;
												assign node16377 = (inp[10]) ? node16383 : node16378;
													assign node16378 = (inp[8]) ? node16380 : 4'b1001;
														assign node16380 = (inp[2]) ? 4'b1000 : 4'b1000;
													assign node16383 = (inp[14]) ? 4'b1110 : node16384;
														assign node16384 = (inp[2]) ? 4'b1110 : 4'b1111;
												assign node16388 = (inp[2]) ? node16390 : 4'b1111;
													assign node16390 = (inp[14]) ? node16392 : 4'b1111;
														assign node16392 = (inp[7]) ? 4'b1111 : 4'b1110;
										assign node16395 = (inp[4]) ? node16413 : node16396;
											assign node16396 = (inp[12]) ? node16404 : node16397;
												assign node16397 = (inp[10]) ? node16399 : 4'b1001;
													assign node16399 = (inp[8]) ? node16401 : 4'b1111;
														assign node16401 = (inp[7]) ? 4'b1110 : 4'b1111;
												assign node16404 = (inp[2]) ? node16408 : node16405;
													assign node16405 = (inp[10]) ? 4'b1110 : 4'b1111;
													assign node16408 = (inp[7]) ? 4'b1110 : node16409;
														assign node16409 = (inp[8]) ? 4'b1111 : 4'b1110;
											assign node16413 = (inp[12]) ? node16425 : node16414;
												assign node16414 = (inp[10]) ? node16420 : node16415;
													assign node16415 = (inp[2]) ? 4'b1110 : node16416;
														assign node16416 = (inp[7]) ? 4'b1110 : 4'b1111;
													assign node16420 = (inp[8]) ? 4'b1011 : node16421;
														assign node16421 = (inp[14]) ? 4'b1010 : 4'b1010;
												assign node16425 = (inp[7]) ? node16427 : 4'b1010;
													assign node16427 = (inp[8]) ? node16429 : 4'b1011;
														assign node16429 = (inp[2]) ? 4'b1010 : 4'b1011;
								assign node16432 = (inp[3]) ? node16528 : node16433;
									assign node16433 = (inp[4]) ? node16477 : node16434;
										assign node16434 = (inp[9]) ? node16456 : node16435;
											assign node16435 = (inp[12]) ? node16449 : node16436;
												assign node16436 = (inp[10]) ? node16444 : node16437;
													assign node16437 = (inp[14]) ? node16441 : node16438;
														assign node16438 = (inp[7]) ? 4'b1100 : 4'b1100;
														assign node16441 = (inp[8]) ? 4'b1101 : 4'b1100;
													assign node16444 = (inp[8]) ? 4'b1000 : node16445;
														assign node16445 = (inp[14]) ? 4'b1000 : 4'b1000;
												assign node16449 = (inp[14]) ? 4'b1000 : node16450;
													assign node16450 = (inp[7]) ? node16452 : 4'b1000;
														assign node16452 = (inp[2]) ? 4'b1001 : 4'b1000;
											assign node16456 = (inp[12]) ? node16466 : node16457;
												assign node16457 = (inp[10]) ? node16463 : node16458;
													assign node16458 = (inp[2]) ? node16460 : 4'b1001;
														assign node16460 = (inp[7]) ? 4'b1000 : 4'b1000;
													assign node16463 = (inp[8]) ? 4'b1110 : 4'b1111;
												assign node16466 = (inp[7]) ? node16472 : node16467;
													assign node16467 = (inp[2]) ? node16469 : 4'b1111;
														assign node16469 = (inp[8]) ? 4'b1111 : 4'b1110;
													assign node16472 = (inp[10]) ? 4'b1110 : node16473;
														assign node16473 = (inp[8]) ? 4'b1110 : 4'b1111;
										assign node16477 = (inp[9]) ? node16503 : node16478;
											assign node16478 = (inp[10]) ? node16490 : node16479;
												assign node16479 = (inp[12]) ? node16485 : node16480;
													assign node16480 = (inp[14]) ? 4'b1001 : node16481;
														assign node16481 = (inp[8]) ? 4'b1000 : 4'b1001;
													assign node16485 = (inp[2]) ? 4'b1110 : node16486;
														assign node16486 = (inp[7]) ? 4'b1111 : 4'b1110;
												assign node16490 = (inp[8]) ? node16496 : node16491;
													assign node16491 = (inp[14]) ? 4'b1111 : node16492;
														assign node16492 = (inp[2]) ? 4'b1110 : 4'b1110;
													assign node16496 = (inp[2]) ? node16500 : node16497;
														assign node16497 = (inp[7]) ? 4'b1110 : 4'b1110;
														assign node16500 = (inp[7]) ? 4'b1110 : 4'b1111;
											assign node16503 = (inp[10]) ? node16517 : node16504;
												assign node16504 = (inp[12]) ? node16510 : node16505;
													assign node16505 = (inp[14]) ? 4'b1110 : node16506;
														assign node16506 = (inp[8]) ? 4'b1110 : 4'b1111;
													assign node16510 = (inp[8]) ? node16514 : node16511;
														assign node16511 = (inp[2]) ? 4'b1010 : 4'b1011;
														assign node16514 = (inp[2]) ? 4'b1011 : 4'b1010;
												assign node16517 = (inp[14]) ? node16523 : node16518;
													assign node16518 = (inp[2]) ? 4'b1011 : node16519;
														assign node16519 = (inp[7]) ? 4'b1010 : 4'b1010;
													assign node16523 = (inp[12]) ? node16525 : 4'b1011;
														assign node16525 = (inp[7]) ? 4'b1010 : 4'b1011;
									assign node16528 = (inp[12]) ? node16576 : node16529;
										assign node16529 = (inp[7]) ? node16555 : node16530;
											assign node16530 = (inp[8]) ? node16542 : node16531;
												assign node16531 = (inp[14]) ? node16537 : node16532;
													assign node16532 = (inp[2]) ? node16534 : 4'b1011;
														assign node16534 = (inp[9]) ? 4'b1010 : 4'b1010;
													assign node16537 = (inp[9]) ? 4'b1110 : node16538;
														assign node16538 = (inp[2]) ? 4'b1110 : 4'b1010;
												assign node16542 = (inp[2]) ? node16550 : node16543;
													assign node16543 = (inp[14]) ? node16547 : node16544;
														assign node16544 = (inp[9]) ? 4'b1010 : 4'b1110;
														assign node16547 = (inp[10]) ? 4'b1011 : 4'b1111;
													assign node16550 = (inp[10]) ? 4'b1111 : node16551;
														assign node16551 = (inp[4]) ? 4'b1111 : 4'b1011;
											assign node16555 = (inp[8]) ? node16567 : node16556;
												assign node16556 = (inp[9]) ? node16562 : node16557;
													assign node16557 = (inp[10]) ? 4'b1111 : node16558;
														assign node16558 = (inp[4]) ? 4'b1011 : 4'b1111;
													assign node16562 = (inp[14]) ? node16564 : 4'b1111;
														assign node16564 = (inp[10]) ? 4'b1011 : 4'b1011;
												assign node16567 = (inp[2]) ? node16571 : node16568;
													assign node16568 = (inp[14]) ? 4'b1010 : 4'b1111;
													assign node16571 = (inp[9]) ? node16573 : 4'b1110;
														assign node16573 = (inp[10]) ? 4'b1010 : 4'b1110;
										assign node16576 = (inp[9]) ? node16598 : node16577;
											assign node16577 = (inp[4]) ? node16591 : node16578;
												assign node16578 = (inp[14]) ? node16584 : node16579;
													assign node16579 = (inp[10]) ? node16581 : 4'b1011;
														assign node16581 = (inp[8]) ? 4'b1010 : 4'b1010;
													assign node16584 = (inp[10]) ? node16588 : node16585;
														assign node16585 = (inp[7]) ? 4'b1010 : 4'b1010;
														assign node16588 = (inp[8]) ? 4'b1010 : 4'b1010;
												assign node16591 = (inp[7]) ? 4'b1110 : node16592;
													assign node16592 = (inp[8]) ? node16594 : 4'b1110;
														assign node16594 = (inp[14]) ? 4'b1111 : 4'b1110;
											assign node16598 = (inp[4]) ? node16610 : node16599;
												assign node16599 = (inp[10]) ? node16605 : node16600;
													assign node16600 = (inp[14]) ? 4'b1111 : node16601;
														assign node16601 = (inp[8]) ? 4'b1110 : 4'b1111;
													assign node16605 = (inp[2]) ? 4'b1110 : node16606;
														assign node16606 = (inp[7]) ? 4'b1110 : 4'b1111;
												assign node16610 = (inp[14]) ? node16618 : node16611;
													assign node16611 = (inp[8]) ? node16615 : node16612;
														assign node16612 = (inp[7]) ? 4'b1010 : 4'b1010;
														assign node16615 = (inp[7]) ? 4'b1010 : 4'b1010;
													assign node16618 = (inp[7]) ? node16620 : 4'b1011;
														assign node16620 = (inp[8]) ? 4'b1010 : 4'b1011;
							assign node16623 = (inp[5]) ? node16807 : node16624;
								assign node16624 = (inp[3]) ? node16726 : node16625;
									assign node16625 = (inp[12]) ? node16681 : node16626;
										assign node16626 = (inp[2]) ? node16652 : node16627;
											assign node16627 = (inp[9]) ? node16639 : node16628;
												assign node16628 = (inp[10]) ? node16634 : node16629;
													assign node16629 = (inp[8]) ? node16631 : 4'b1010;
														assign node16631 = (inp[7]) ? 4'b1010 : 4'b1011;
													assign node16634 = (inp[4]) ? 4'b1111 : node16635;
														assign node16635 = (inp[7]) ? 4'b1011 : 4'b1010;
												assign node16639 = (inp[8]) ? node16645 : node16640;
													assign node16640 = (inp[14]) ? 4'b1110 : node16641;
														assign node16641 = (inp[7]) ? 4'b1010 : 4'b1011;
													assign node16645 = (inp[4]) ? node16649 : node16646;
														assign node16646 = (inp[10]) ? 4'b1111 : 4'b1011;
														assign node16649 = (inp[10]) ? 4'b1010 : 4'b1110;
											assign node16652 = (inp[14]) ? node16668 : node16653;
												assign node16653 = (inp[9]) ? node16661 : node16654;
													assign node16654 = (inp[8]) ? node16658 : node16655;
														assign node16655 = (inp[7]) ? 4'b1011 : 4'b1010;
														assign node16658 = (inp[4]) ? 4'b1010 : 4'b1111;
													assign node16661 = (inp[7]) ? node16665 : node16662;
														assign node16662 = (inp[10]) ? 4'b1111 : 4'b1010;
														assign node16665 = (inp[10]) ? 4'b1010 : 4'b1010;
												assign node16668 = (inp[10]) ? node16676 : node16669;
													assign node16669 = (inp[7]) ? node16673 : node16670;
														assign node16670 = (inp[8]) ? 4'b1111 : 4'b1010;
														assign node16673 = (inp[8]) ? 4'b1010 : 4'b1011;
													assign node16676 = (inp[8]) ? 4'b1011 : node16677;
														assign node16677 = (inp[4]) ? 4'b1011 : 4'b1111;
										assign node16681 = (inp[4]) ? node16703 : node16682;
											assign node16682 = (inp[9]) ? node16690 : node16683;
												assign node16683 = (inp[2]) ? 4'b1011 : node16684;
													assign node16684 = (inp[7]) ? node16686 : 4'b1011;
														assign node16686 = (inp[10]) ? 4'b1010 : 4'b1010;
												assign node16690 = (inp[14]) ? node16698 : node16691;
													assign node16691 = (inp[2]) ? node16695 : node16692;
														assign node16692 = (inp[8]) ? 4'b1110 : 4'b1110;
														assign node16695 = (inp[8]) ? 4'b1110 : 4'b1110;
													assign node16698 = (inp[2]) ? 4'b1111 : node16699;
														assign node16699 = (inp[8]) ? 4'b1110 : 4'b1110;
											assign node16703 = (inp[9]) ? node16711 : node16704;
												assign node16704 = (inp[2]) ? 4'b1111 : node16705;
													assign node16705 = (inp[7]) ? node16707 : 4'b1111;
														assign node16707 = (inp[8]) ? 4'b1110 : 4'b1111;
												assign node16711 = (inp[2]) ? node16719 : node16712;
													assign node16712 = (inp[8]) ? node16716 : node16713;
														assign node16713 = (inp[14]) ? 4'b1010 : 4'b1011;
														assign node16716 = (inp[14]) ? 4'b1011 : 4'b1010;
													assign node16719 = (inp[14]) ? node16723 : node16720;
														assign node16720 = (inp[10]) ? 4'b1010 : 4'b1011;
														assign node16723 = (inp[8]) ? 4'b1010 : 4'b1010;
									assign node16726 = (inp[4]) ? node16766 : node16727;
										assign node16727 = (inp[9]) ? node16751 : node16728;
											assign node16728 = (inp[8]) ? node16742 : node16729;
												assign node16729 = (inp[12]) ? node16737 : node16730;
													assign node16730 = (inp[10]) ? node16734 : node16731;
														assign node16731 = (inp[14]) ? 4'b1110 : 4'b1111;
														assign node16734 = (inp[2]) ? 4'b1010 : 4'b1010;
													assign node16737 = (inp[10]) ? node16739 : 4'b1010;
														assign node16739 = (inp[2]) ? 4'b1011 : 4'b1010;
												assign node16742 = (inp[14]) ? node16748 : node16743;
													assign node16743 = (inp[7]) ? 4'b1011 : node16744;
														assign node16744 = (inp[2]) ? 4'b1011 : 4'b1010;
													assign node16748 = (inp[7]) ? 4'b1010 : 4'b1011;
											assign node16751 = (inp[12]) ? node16757 : node16752;
												assign node16752 = (inp[10]) ? node16754 : 4'b1011;
													assign node16754 = (inp[2]) ? 4'b1101 : 4'b1100;
												assign node16757 = (inp[2]) ? node16759 : 4'b1100;
													assign node16759 = (inp[7]) ? node16763 : node16760;
														assign node16760 = (inp[8]) ? 4'b1101 : 4'b1100;
														assign node16763 = (inp[8]) ? 4'b1100 : 4'b1101;
										assign node16766 = (inp[9]) ? node16788 : node16767;
											assign node16767 = (inp[12]) ? node16777 : node16768;
												assign node16768 = (inp[10]) ? node16774 : node16769;
													assign node16769 = (inp[7]) ? 4'b1010 : node16770;
														assign node16770 = (inp[2]) ? 4'b1011 : 4'b1010;
													assign node16774 = (inp[7]) ? 4'b1101 : 4'b1100;
												assign node16777 = (inp[14]) ? node16783 : node16778;
													assign node16778 = (inp[7]) ? node16780 : 4'b1100;
														assign node16780 = (inp[8]) ? 4'b1100 : 4'b1100;
													assign node16783 = (inp[2]) ? 4'b1101 : node16784;
														assign node16784 = (inp[7]) ? 4'b1100 : 4'b1101;
											assign node16788 = (inp[7]) ? node16800 : node16789;
												assign node16789 = (inp[14]) ? node16797 : node16790;
													assign node16790 = (inp[8]) ? node16794 : node16791;
														assign node16791 = (inp[2]) ? 4'b1000 : 4'b1001;
														assign node16794 = (inp[2]) ? 4'b1001 : 4'b1000;
													assign node16797 = (inp[10]) ? 4'b1000 : 4'b1100;
												assign node16800 = (inp[8]) ? node16804 : node16801;
													assign node16801 = (inp[2]) ? 4'b1001 : 4'b1101;
													assign node16804 = (inp[2]) ? 4'b1000 : 4'b1001;
								assign node16807 = (inp[3]) ? node16901 : node16808;
									assign node16808 = (inp[9]) ? node16854 : node16809;
										assign node16809 = (inp[4]) ? node16833 : node16810;
											assign node16810 = (inp[10]) ? node16822 : node16811;
												assign node16811 = (inp[12]) ? node16817 : node16812;
													assign node16812 = (inp[8]) ? 4'b1111 : node16813;
														assign node16813 = (inp[2]) ? 4'b1110 : 4'b1111;
													assign node16817 = (inp[7]) ? 4'b1011 : node16818;
														assign node16818 = (inp[14]) ? 4'b1011 : 4'b1010;
												assign node16822 = (inp[7]) ? node16828 : node16823;
													assign node16823 = (inp[8]) ? node16825 : 4'b1010;
														assign node16825 = (inp[2]) ? 4'b1011 : 4'b1010;
													assign node16828 = (inp[14]) ? 4'b1011 : node16829;
														assign node16829 = (inp[8]) ? 4'b1011 : 4'b1010;
											assign node16833 = (inp[12]) ? node16845 : node16834;
												assign node16834 = (inp[10]) ? node16840 : node16835;
													assign node16835 = (inp[2]) ? 4'b1011 : node16836;
														assign node16836 = (inp[14]) ? 4'b1011 : 4'b1010;
													assign node16840 = (inp[8]) ? node16842 : 4'b1101;
														assign node16842 = (inp[7]) ? 4'b1100 : 4'b1100;
												assign node16845 = (inp[8]) ? node16849 : node16846;
													assign node16846 = (inp[7]) ? 4'b1101 : 4'b1100;
													assign node16849 = (inp[7]) ? 4'b1100 : node16850;
														assign node16850 = (inp[14]) ? 4'b1101 : 4'b1100;
										assign node16854 = (inp[4]) ? node16878 : node16855;
											assign node16855 = (inp[10]) ? node16867 : node16856;
												assign node16856 = (inp[12]) ? node16860 : node16857;
													assign node16857 = (inp[14]) ? 4'b1010 : 4'b1011;
													assign node16860 = (inp[14]) ? node16864 : node16861;
														assign node16861 = (inp[2]) ? 4'b1100 : 4'b1101;
														assign node16864 = (inp[8]) ? 4'b1100 : 4'b1100;
												assign node16867 = (inp[7]) ? node16873 : node16868;
													assign node16868 = (inp[8]) ? 4'b1101 : node16869;
														assign node16869 = (inp[14]) ? 4'b1100 : 4'b1101;
													assign node16873 = (inp[14]) ? node16875 : 4'b1100;
														assign node16875 = (inp[8]) ? 4'b1100 : 4'b1101;
											assign node16878 = (inp[12]) ? node16890 : node16879;
												assign node16879 = (inp[10]) ? node16885 : node16880;
													assign node16880 = (inp[8]) ? node16882 : 4'b1101;
														assign node16882 = (inp[2]) ? 4'b1100 : 4'b1100;
													assign node16885 = (inp[7]) ? 4'b1001 : node16886;
														assign node16886 = (inp[8]) ? 4'b1001 : 4'b1000;
												assign node16890 = (inp[14]) ? node16896 : node16891;
													assign node16891 = (inp[8]) ? node16893 : 4'b1000;
														assign node16893 = (inp[10]) ? 4'b1000 : 4'b1001;
													assign node16896 = (inp[2]) ? 4'b1001 : node16897;
														assign node16897 = (inp[7]) ? 4'b1000 : 4'b1001;
									assign node16901 = (inp[9]) ? node16945 : node16902;
										assign node16902 = (inp[4]) ? node16922 : node16903;
											assign node16903 = (inp[12]) ? node16909 : node16904;
												assign node16904 = (inp[10]) ? node16906 : 4'b1101;
													assign node16906 = (inp[8]) ? 4'b1000 : 4'b1001;
												assign node16909 = (inp[14]) ? node16915 : node16910;
													assign node16910 = (inp[10]) ? 4'b1001 : node16911;
														assign node16911 = (inp[8]) ? 4'b1001 : 4'b1000;
													assign node16915 = (inp[10]) ? node16919 : node16916;
														assign node16916 = (inp[8]) ? 4'b1001 : 4'b1000;
														assign node16919 = (inp[8]) ? 4'b1000 : 4'b1001;
											assign node16922 = (inp[12]) ? node16934 : node16923;
												assign node16923 = (inp[10]) ? node16929 : node16924;
													assign node16924 = (inp[14]) ? node16926 : 4'b1001;
														assign node16926 = (inp[7]) ? 4'b1000 : 4'b1000;
													assign node16929 = (inp[2]) ? node16931 : 4'b1101;
														assign node16931 = (inp[7]) ? 4'b1100 : 4'b1101;
												assign node16934 = (inp[7]) ? node16940 : node16935;
													assign node16935 = (inp[8]) ? node16937 : 4'b1100;
														assign node16937 = (inp[14]) ? 4'b1101 : 4'b1100;
													assign node16940 = (inp[2]) ? node16942 : 4'b1101;
														assign node16942 = (inp[8]) ? 4'b1100 : 4'b1101;
										assign node16945 = (inp[4]) ? node16975 : node16946;
											assign node16946 = (inp[10]) ? node16962 : node16947;
												assign node16947 = (inp[12]) ? node16955 : node16948;
													assign node16948 = (inp[2]) ? node16952 : node16949;
														assign node16949 = (inp[8]) ? 4'b1000 : 4'b1001;
														assign node16952 = (inp[8]) ? 4'b1001 : 4'b1000;
													assign node16955 = (inp[2]) ? node16959 : node16956;
														assign node16956 = (inp[14]) ? 4'b1100 : 4'b1101;
														assign node16959 = (inp[8]) ? 4'b1101 : 4'b1100;
												assign node16962 = (inp[2]) ? node16970 : node16963;
													assign node16963 = (inp[8]) ? node16967 : node16964;
														assign node16964 = (inp[12]) ? 4'b1100 : 4'b1100;
														assign node16967 = (inp[12]) ? 4'b1101 : 4'b1100;
													assign node16970 = (inp[12]) ? 4'b1101 : node16971;
														assign node16971 = (inp[7]) ? 4'b1100 : 4'b1101;
											assign node16975 = (inp[10]) ? node16987 : node16976;
												assign node16976 = (inp[12]) ? node16982 : node16977;
													assign node16977 = (inp[14]) ? node16979 : 4'b1100;
														assign node16979 = (inp[7]) ? 4'b1101 : 4'b1100;
													assign node16982 = (inp[8]) ? node16984 : 4'b1000;
														assign node16984 = (inp[7]) ? 4'b1001 : 4'b1000;
												assign node16987 = (inp[7]) ? node16993 : node16988;
													assign node16988 = (inp[14]) ? 4'b1001 : node16989;
														assign node16989 = (inp[12]) ? 4'b1000 : 4'b1000;
													assign node16993 = (inp[8]) ? 4'b1000 : node16994;
														assign node16994 = (inp[14]) ? 4'b1001 : 4'b1000;
			assign node16998 = (inp[11]) ? node19874 : node16999;
				assign node16999 = (inp[1]) ? node18443 : node17000;
					assign node17000 = (inp[13]) ? node17742 : node17001;
						assign node17001 = (inp[15]) ? node17373 : node17002;
							assign node17002 = (inp[3]) ? node17192 : node17003;
								assign node17003 = (inp[5]) ? node17101 : node17004;
									assign node17004 = (inp[9]) ? node17050 : node17005;
										assign node17005 = (inp[4]) ? node17025 : node17006;
											assign node17006 = (inp[10]) ? node17016 : node17007;
												assign node17007 = (inp[2]) ? 4'b0100 : node17008;
													assign node17008 = (inp[14]) ? node17012 : node17009;
														assign node17009 = (inp[8]) ? 4'b0100 : 4'b0100;
														assign node17012 = (inp[7]) ? 4'b0100 : 4'b0101;
												assign node17016 = (inp[12]) ? node17020 : node17017;
													assign node17017 = (inp[7]) ? 4'b0100 : 4'b0101;
													assign node17020 = (inp[14]) ? node17022 : 4'b0000;
														assign node17022 = (inp[7]) ? 4'b0000 : 4'b0000;
											assign node17025 = (inp[12]) ? node17039 : node17026;
												assign node17026 = (inp[10]) ? node17034 : node17027;
													assign node17027 = (inp[7]) ? node17031 : node17028;
														assign node17028 = (inp[8]) ? 4'b0001 : 4'b0000;
														assign node17031 = (inp[8]) ? 4'b0000 : 4'b0000;
													assign node17034 = (inp[7]) ? node17036 : 4'b0000;
														assign node17036 = (inp[2]) ? 4'b0001 : 4'b0000;
												assign node17039 = (inp[10]) ? node17045 : node17040;
													assign node17040 = (inp[2]) ? node17042 : 4'b0000;
														assign node17042 = (inp[8]) ? 4'b0001 : 4'b0000;
													assign node17045 = (inp[8]) ? 4'b0100 : node17046;
														assign node17046 = (inp[2]) ? 4'b0100 : 4'b0101;
										assign node17050 = (inp[4]) ? node17078 : node17051;
											assign node17051 = (inp[10]) ? node17067 : node17052;
												assign node17052 = (inp[2]) ? node17060 : node17053;
													assign node17053 = (inp[8]) ? node17057 : node17054;
														assign node17054 = (inp[12]) ? 4'b0001 : 4'b0000;
														assign node17057 = (inp[14]) ? 4'b0000 : 4'b0000;
													assign node17060 = (inp[12]) ? node17064 : node17061;
														assign node17061 = (inp[7]) ? 4'b0001 : 4'b0000;
														assign node17064 = (inp[14]) ? 4'b0000 : 4'b0000;
												assign node17067 = (inp[12]) ? node17073 : node17068;
													assign node17068 = (inp[7]) ? 4'b0001 : node17069;
														assign node17069 = (inp[8]) ? 4'b0001 : 4'b0000;
													assign node17073 = (inp[8]) ? 4'b0100 : node17074;
														assign node17074 = (inp[2]) ? 4'b0100 : 4'b0101;
											assign node17078 = (inp[10]) ? node17090 : node17079;
												assign node17079 = (inp[14]) ? node17085 : node17080;
													assign node17080 = (inp[2]) ? node17082 : 4'b0100;
														assign node17082 = (inp[8]) ? 4'b0100 : 4'b0100;
													assign node17085 = (inp[2]) ? node17087 : 4'b0101;
														assign node17087 = (inp[7]) ? 4'b0100 : 4'b0100;
												assign node17090 = (inp[12]) ? node17096 : node17091;
													assign node17091 = (inp[8]) ? 4'b0101 : node17092;
														assign node17092 = (inp[7]) ? 4'b0101 : 4'b0100;
													assign node17096 = (inp[7]) ? 4'b0001 : node17097;
														assign node17097 = (inp[14]) ? 4'b0001 : 4'b0000;
									assign node17101 = (inp[9]) ? node17151 : node17102;
										assign node17102 = (inp[4]) ? node17128 : node17103;
											assign node17103 = (inp[12]) ? node17117 : node17104;
												assign node17104 = (inp[2]) ? node17110 : node17105;
													assign node17105 = (inp[8]) ? 4'b0100 : node17106;
														assign node17106 = (inp[14]) ? 4'b0100 : 4'b0100;
													assign node17110 = (inp[14]) ? node17114 : node17111;
														assign node17111 = (inp[8]) ? 4'b0101 : 4'b0100;
														assign node17114 = (inp[8]) ? 4'b0100 : 4'b0101;
												assign node17117 = (inp[10]) ? node17121 : node17118;
													assign node17118 = (inp[7]) ? 4'b0101 : 4'b0100;
													assign node17121 = (inp[2]) ? node17125 : node17122;
														assign node17122 = (inp[8]) ? 4'b0000 : 4'b0000;
														assign node17125 = (inp[8]) ? 4'b0001 : 4'b0000;
											assign node17128 = (inp[12]) ? node17142 : node17129;
												assign node17129 = (inp[7]) ? node17135 : node17130;
													assign node17130 = (inp[8]) ? 4'b0001 : node17131;
														assign node17131 = (inp[2]) ? 4'b0000 : 4'b0001;
													assign node17135 = (inp[2]) ? node17139 : node17136;
														assign node17136 = (inp[8]) ? 4'b0000 : 4'b0000;
														assign node17139 = (inp[8]) ? 4'b0000 : 4'b0001;
												assign node17142 = (inp[10]) ? node17146 : node17143;
													assign node17143 = (inp[8]) ? 4'b0000 : 4'b0001;
													assign node17146 = (inp[8]) ? 4'b0111 : node17147;
														assign node17147 = (inp[14]) ? 4'b0110 : 4'b0110;
										assign node17151 = (inp[4]) ? node17171 : node17152;
											assign node17152 = (inp[10]) ? node17164 : node17153;
												assign node17153 = (inp[14]) ? node17159 : node17154;
													assign node17154 = (inp[8]) ? 4'b0000 : node17155;
														assign node17155 = (inp[7]) ? 4'b0000 : 4'b0000;
													assign node17159 = (inp[7]) ? node17161 : 4'b0001;
														assign node17161 = (inp[8]) ? 4'b0000 : 4'b0001;
												assign node17164 = (inp[12]) ? node17166 : 4'b0000;
													assign node17166 = (inp[7]) ? node17168 : 4'b0111;
														assign node17168 = (inp[2]) ? 4'b0110 : 4'b0111;
											assign node17171 = (inp[2]) ? node17181 : node17172;
												assign node17172 = (inp[10]) ? node17178 : node17173;
													assign node17173 = (inp[8]) ? 4'b0110 : node17174;
														assign node17174 = (inp[12]) ? 4'b0111 : 4'b0110;
													assign node17178 = (inp[12]) ? 4'b0011 : 4'b0111;
												assign node17181 = (inp[10]) ? node17189 : node17182;
													assign node17182 = (inp[8]) ? node17186 : node17183;
														assign node17183 = (inp[7]) ? 4'b0111 : 4'b0110;
														assign node17186 = (inp[7]) ? 4'b0110 : 4'b0111;
													assign node17189 = (inp[12]) ? 4'b0010 : 4'b0110;
								assign node17192 = (inp[5]) ? node17286 : node17193;
									assign node17193 = (inp[9]) ? node17233 : node17194;
										assign node17194 = (inp[4]) ? node17216 : node17195;
											assign node17195 = (inp[12]) ? node17207 : node17196;
												assign node17196 = (inp[8]) ? node17202 : node17197;
													assign node17197 = (inp[7]) ? node17199 : 4'b0100;
														assign node17199 = (inp[2]) ? 4'b0101 : 4'b0100;
													assign node17202 = (inp[7]) ? node17204 : 4'b0101;
														assign node17204 = (inp[2]) ? 4'b0100 : 4'b0100;
												assign node17207 = (inp[10]) ? 4'b0000 : node17208;
													assign node17208 = (inp[8]) ? node17212 : node17209;
														assign node17209 = (inp[7]) ? 4'b0101 : 4'b0100;
														assign node17212 = (inp[7]) ? 4'b0100 : 4'b0101;
											assign node17216 = (inp[12]) ? node17224 : node17217;
												assign node17217 = (inp[8]) ? 4'b0000 : node17218;
													assign node17218 = (inp[7]) ? 4'b0001 : node17219;
														assign node17219 = (inp[2]) ? 4'b0000 : 4'b0000;
												assign node17224 = (inp[10]) ? node17228 : node17225;
													assign node17225 = (inp[7]) ? 4'b0001 : 4'b0000;
													assign node17228 = (inp[7]) ? 4'b0110 : node17229;
														assign node17229 = (inp[2]) ? 4'b0110 : 4'b0111;
										assign node17233 = (inp[4]) ? node17259 : node17234;
											assign node17234 = (inp[12]) ? node17246 : node17235;
												assign node17235 = (inp[14]) ? node17241 : node17236;
													assign node17236 = (inp[10]) ? node17238 : 4'b0000;
														assign node17238 = (inp[8]) ? 4'b0001 : 4'b0001;
													assign node17241 = (inp[10]) ? 4'b0000 : node17242;
														assign node17242 = (inp[7]) ? 4'b0001 : 4'b0000;
												assign node17246 = (inp[10]) ? node17252 : node17247;
													assign node17247 = (inp[2]) ? node17249 : 4'b0001;
														assign node17249 = (inp[7]) ? 4'b0000 : 4'b0000;
													assign node17252 = (inp[7]) ? node17256 : node17253;
														assign node17253 = (inp[8]) ? 4'b0111 : 4'b0110;
														assign node17256 = (inp[14]) ? 4'b0110 : 4'b0110;
											assign node17259 = (inp[10]) ? node17273 : node17260;
												assign node17260 = (inp[8]) ? node17266 : node17261;
													assign node17261 = (inp[7]) ? 4'b0111 : node17262;
														assign node17262 = (inp[12]) ? 4'b0111 : 4'b0110;
													assign node17266 = (inp[7]) ? node17270 : node17267;
														assign node17267 = (inp[2]) ? 4'b0111 : 4'b0110;
														assign node17270 = (inp[2]) ? 4'b0110 : 4'b0110;
												assign node17273 = (inp[12]) ? node17279 : node17274;
													assign node17274 = (inp[8]) ? 4'b0111 : node17275;
														assign node17275 = (inp[7]) ? 4'b0110 : 4'b0110;
													assign node17279 = (inp[7]) ? node17283 : node17280;
														assign node17280 = (inp[8]) ? 4'b0011 : 4'b0010;
														assign node17283 = (inp[2]) ? 4'b0010 : 4'b0011;
									assign node17286 = (inp[8]) ? node17330 : node17287;
										assign node17287 = (inp[7]) ? node17317 : node17288;
											assign node17288 = (inp[2]) ? node17304 : node17289;
												assign node17289 = (inp[14]) ? node17297 : node17290;
													assign node17290 = (inp[9]) ? node17294 : node17291;
														assign node17291 = (inp[4]) ? 4'b0011 : 4'b0111;
														assign node17294 = (inp[4]) ? 4'b0111 : 4'b0011;
													assign node17297 = (inp[4]) ? node17301 : node17298;
														assign node17298 = (inp[9]) ? 4'b0010 : 4'b0110;
														assign node17301 = (inp[12]) ? 4'b0110 : 4'b0010;
												assign node17304 = (inp[10]) ? node17312 : node17305;
													assign node17305 = (inp[4]) ? node17309 : node17306;
														assign node17306 = (inp[9]) ? 4'b0010 : 4'b0110;
														assign node17309 = (inp[9]) ? 4'b0110 : 4'b0010;
													assign node17312 = (inp[4]) ? 4'b0110 : node17313;
														assign node17313 = (inp[9]) ? 4'b0010 : 4'b0110;
											assign node17317 = (inp[14]) ? node17325 : node17318;
												assign node17318 = (inp[2]) ? 4'b0011 : node17319;
													assign node17319 = (inp[10]) ? node17321 : 4'b0010;
														assign node17321 = (inp[4]) ? 4'b0110 : 4'b0010;
												assign node17325 = (inp[10]) ? 4'b0111 : node17326;
													assign node17326 = (inp[2]) ? 4'b0011 : 4'b0111;
										assign node17330 = (inp[7]) ? node17354 : node17331;
											assign node17331 = (inp[14]) ? node17343 : node17332;
												assign node17332 = (inp[2]) ? node17338 : node17333;
													assign node17333 = (inp[12]) ? node17335 : 4'b0010;
														assign node17335 = (inp[9]) ? 4'b0110 : 4'b0010;
													assign node17338 = (inp[4]) ? node17340 : 4'b0011;
														assign node17340 = (inp[9]) ? 4'b0111 : 4'b0011;
												assign node17343 = (inp[9]) ? node17349 : node17344;
													assign node17344 = (inp[2]) ? 4'b0011 : node17345;
														assign node17345 = (inp[12]) ? 4'b0011 : 4'b0111;
													assign node17349 = (inp[2]) ? node17351 : 4'b0111;
														assign node17351 = (inp[12]) ? 4'b0011 : 4'b0111;
											assign node17354 = (inp[2]) ? node17362 : node17355;
												assign node17355 = (inp[14]) ? 4'b0010 : node17356;
													assign node17356 = (inp[12]) ? node17358 : 4'b0111;
														assign node17358 = (inp[4]) ? 4'b0111 : 4'b0011;
												assign node17362 = (inp[10]) ? node17368 : node17363;
													assign node17363 = (inp[14]) ? 4'b0110 : node17364;
														assign node17364 = (inp[12]) ? 4'b0110 : 4'b0010;
													assign node17368 = (inp[9]) ? node17370 : 4'b0010;
														assign node17370 = (inp[4]) ? 4'b0110 : 4'b0010;
							assign node17373 = (inp[5]) ? node17567 : node17374;
								assign node17374 = (inp[3]) ? node17466 : node17375;
									assign node17375 = (inp[4]) ? node17423 : node17376;
										assign node17376 = (inp[9]) ? node17396 : node17377;
											assign node17377 = (inp[10]) ? node17389 : node17378;
												assign node17378 = (inp[12]) ? node17386 : node17379;
													assign node17379 = (inp[7]) ? node17383 : node17380;
														assign node17380 = (inp[8]) ? 4'b0111 : 4'b0110;
														assign node17383 = (inp[8]) ? 4'b0110 : 4'b0111;
													assign node17386 = (inp[8]) ? 4'b0111 : 4'b0110;
												assign node17389 = (inp[12]) ? 4'b0011 : node17390;
													assign node17390 = (inp[7]) ? 4'b0111 : node17391;
														assign node17391 = (inp[14]) ? 4'b0111 : 4'b0110;
											assign node17396 = (inp[10]) ? node17410 : node17397;
												assign node17397 = (inp[14]) ? node17403 : node17398;
													assign node17398 = (inp[8]) ? node17400 : 4'b0010;
														assign node17400 = (inp[12]) ? 4'b0010 : 4'b0011;
													assign node17403 = (inp[12]) ? node17407 : node17404;
														assign node17404 = (inp[8]) ? 4'b0010 : 4'b0011;
														assign node17407 = (inp[8]) ? 4'b0011 : 4'b0010;
												assign node17410 = (inp[12]) ? node17416 : node17411;
													assign node17411 = (inp[14]) ? 4'b0011 : node17412;
														assign node17412 = (inp[8]) ? 4'b0010 : 4'b0010;
													assign node17416 = (inp[7]) ? node17420 : node17417;
														assign node17417 = (inp[8]) ? 4'b0111 : 4'b0110;
														assign node17420 = (inp[8]) ? 4'b0110 : 4'b0111;
										assign node17423 = (inp[9]) ? node17449 : node17424;
											assign node17424 = (inp[10]) ? node17436 : node17425;
												assign node17425 = (inp[2]) ? node17431 : node17426;
													assign node17426 = (inp[14]) ? 4'b0011 : node17427;
														assign node17427 = (inp[12]) ? 4'b0011 : 4'b0010;
													assign node17431 = (inp[12]) ? node17433 : 4'b0011;
														assign node17433 = (inp[8]) ? 4'b0010 : 4'b0010;
												assign node17436 = (inp[12]) ? node17444 : node17437;
													assign node17437 = (inp[2]) ? node17441 : node17438;
														assign node17438 = (inp[8]) ? 4'b0010 : 4'b0010;
														assign node17441 = (inp[7]) ? 4'b0011 : 4'b0011;
													assign node17444 = (inp[2]) ? 4'b0110 : node17445;
														assign node17445 = (inp[7]) ? 4'b0110 : 4'b0111;
											assign node17449 = (inp[10]) ? node17455 : node17450;
												assign node17450 = (inp[8]) ? node17452 : 4'b0111;
													assign node17452 = (inp[7]) ? 4'b0110 : 4'b0111;
												assign node17455 = (inp[12]) ? node17461 : node17456;
													assign node17456 = (inp[8]) ? 4'b0110 : node17457;
														assign node17457 = (inp[7]) ? 4'b0110 : 4'b0110;
													assign node17461 = (inp[14]) ? node17463 : 4'b0010;
														assign node17463 = (inp[7]) ? 4'b0010 : 4'b0011;
									assign node17466 = (inp[9]) ? node17518 : node17467;
										assign node17467 = (inp[4]) ? node17493 : node17468;
											assign node17468 = (inp[10]) ? node17482 : node17469;
												assign node17469 = (inp[12]) ? node17477 : node17470;
													assign node17470 = (inp[2]) ? node17474 : node17471;
														assign node17471 = (inp[7]) ? 4'b0111 : 4'b0110;
														assign node17474 = (inp[7]) ? 4'b0110 : 4'b0111;
													assign node17477 = (inp[8]) ? 4'b0111 : node17478;
														assign node17478 = (inp[14]) ? 4'b0110 : 4'b0111;
												assign node17482 = (inp[12]) ? node17488 : node17483;
													assign node17483 = (inp[7]) ? 4'b0110 : node17484;
														assign node17484 = (inp[2]) ? 4'b0110 : 4'b0111;
													assign node17488 = (inp[14]) ? 4'b0010 : node17489;
														assign node17489 = (inp[7]) ? 4'b0010 : 4'b0011;
											assign node17493 = (inp[10]) ? node17507 : node17494;
												assign node17494 = (inp[2]) ? node17500 : node17495;
													assign node17495 = (inp[14]) ? node17497 : 4'b0010;
														assign node17497 = (inp[8]) ? 4'b0011 : 4'b0010;
													assign node17500 = (inp[12]) ? node17504 : node17501;
														assign node17501 = (inp[8]) ? 4'b0011 : 4'b0010;
														assign node17504 = (inp[8]) ? 4'b0010 : 4'b0011;
												assign node17507 = (inp[12]) ? node17513 : node17508;
													assign node17508 = (inp[8]) ? 4'b0011 : node17509;
														assign node17509 = (inp[14]) ? 4'b0010 : 4'b0010;
													assign node17513 = (inp[8]) ? 4'b0101 : node17514;
														assign node17514 = (inp[14]) ? 4'b0100 : 4'b0101;
										assign node17518 = (inp[4]) ? node17544 : node17519;
											assign node17519 = (inp[12]) ? node17533 : node17520;
												assign node17520 = (inp[14]) ? node17528 : node17521;
													assign node17521 = (inp[2]) ? node17525 : node17522;
														assign node17522 = (inp[8]) ? 4'b0010 : 4'b0010;
														assign node17525 = (inp[10]) ? 4'b0011 : 4'b0011;
													assign node17528 = (inp[8]) ? 4'b0010 : node17529;
														assign node17529 = (inp[10]) ? 4'b0011 : 4'b0010;
												assign node17533 = (inp[10]) ? node17539 : node17534;
													assign node17534 = (inp[2]) ? 4'b0011 : node17535;
														assign node17535 = (inp[14]) ? 4'b0011 : 4'b0010;
													assign node17539 = (inp[8]) ? 4'b0101 : node17540;
														assign node17540 = (inp[14]) ? 4'b0100 : 4'b0100;
											assign node17544 = (inp[10]) ? node17554 : node17545;
												assign node17545 = (inp[14]) ? node17549 : node17546;
													assign node17546 = (inp[8]) ? 4'b0101 : 4'b0100;
													assign node17549 = (inp[2]) ? node17551 : 4'b0100;
														assign node17551 = (inp[8]) ? 4'b0100 : 4'b0100;
												assign node17554 = (inp[12]) ? node17562 : node17555;
													assign node17555 = (inp[7]) ? node17559 : node17556;
														assign node17556 = (inp[8]) ? 4'b0101 : 4'b0100;
														assign node17559 = (inp[8]) ? 4'b0100 : 4'b0101;
													assign node17562 = (inp[7]) ? node17564 : 4'b0001;
														assign node17564 = (inp[14]) ? 4'b0000 : 4'b0000;
								assign node17567 = (inp[3]) ? node17649 : node17568;
									assign node17568 = (inp[4]) ? node17608 : node17569;
										assign node17569 = (inp[9]) ? node17591 : node17570;
											assign node17570 = (inp[12]) ? node17580 : node17571;
												assign node17571 = (inp[14]) ? node17573 : 4'b0110;
													assign node17573 = (inp[10]) ? node17577 : node17574;
														assign node17574 = (inp[8]) ? 4'b0110 : 4'b0110;
														assign node17577 = (inp[8]) ? 4'b0111 : 4'b0110;
												assign node17580 = (inp[10]) ? node17584 : node17581;
													assign node17581 = (inp[14]) ? 4'b0110 : 4'b0111;
													assign node17584 = (inp[14]) ? node17588 : node17585;
														assign node17585 = (inp[7]) ? 4'b0010 : 4'b0011;
														assign node17588 = (inp[7]) ? 4'b0010 : 4'b0010;
											assign node17591 = (inp[10]) ? node17597 : node17592;
												assign node17592 = (inp[7]) ? node17594 : 4'b0010;
													assign node17594 = (inp[8]) ? 4'b0010 : 4'b0011;
												assign node17597 = (inp[12]) ? node17603 : node17598;
													assign node17598 = (inp[14]) ? node17600 : 4'b0010;
														assign node17600 = (inp[8]) ? 4'b0011 : 4'b0010;
													assign node17603 = (inp[14]) ? node17605 : 4'b0101;
														assign node17605 = (inp[8]) ? 4'b0101 : 4'b0100;
										assign node17608 = (inp[9]) ? node17630 : node17609;
											assign node17609 = (inp[12]) ? node17621 : node17610;
												assign node17610 = (inp[8]) ? node17616 : node17611;
													assign node17611 = (inp[2]) ? 4'b0011 : node17612;
														assign node17612 = (inp[14]) ? 4'b0010 : 4'b0010;
													assign node17616 = (inp[7]) ? 4'b0010 : node17617;
														assign node17617 = (inp[2]) ? 4'b0011 : 4'b0010;
												assign node17621 = (inp[10]) ? node17625 : node17622;
													assign node17622 = (inp[8]) ? 4'b0010 : 4'b0011;
													assign node17625 = (inp[7]) ? 4'b0101 : node17626;
														assign node17626 = (inp[8]) ? 4'b0101 : 4'b0100;
											assign node17630 = (inp[10]) ? node17640 : node17631;
												assign node17631 = (inp[7]) ? node17633 : 4'b0100;
													assign node17633 = (inp[8]) ? node17637 : node17634;
														assign node17634 = (inp[14]) ? 4'b0101 : 4'b0100;
														assign node17637 = (inp[14]) ? 4'b0100 : 4'b0101;
												assign node17640 = (inp[12]) ? node17644 : node17641;
													assign node17641 = (inp[7]) ? 4'b0101 : 4'b0100;
													assign node17644 = (inp[7]) ? 4'b0001 : node17645;
														assign node17645 = (inp[8]) ? 4'b0001 : 4'b0000;
									assign node17649 = (inp[12]) ? node17693 : node17650;
										assign node17650 = (inp[7]) ? node17674 : node17651;
											assign node17651 = (inp[8]) ? node17661 : node17652;
												assign node17652 = (inp[2]) ? node17656 : node17653;
													assign node17653 = (inp[14]) ? 4'b0000 : 4'b0001;
													assign node17656 = (inp[14]) ? 4'b0100 : node17657;
														assign node17657 = (inp[9]) ? 4'b0000 : 4'b0100;
												assign node17661 = (inp[2]) ? node17669 : node17662;
													assign node17662 = (inp[9]) ? node17666 : node17663;
														assign node17663 = (inp[4]) ? 4'b0000 : 4'b0100;
														assign node17666 = (inp[10]) ? 4'b0001 : 4'b0101;
													assign node17669 = (inp[10]) ? node17671 : 4'b0001;
														assign node17671 = (inp[4]) ? 4'b0001 : 4'b0101;
											assign node17674 = (inp[8]) ? node17682 : node17675;
												assign node17675 = (inp[4]) ? node17677 : 4'b0101;
													assign node17677 = (inp[2]) ? node17679 : 4'b0000;
														assign node17679 = (inp[9]) ? 4'b0101 : 4'b0001;
												assign node17682 = (inp[2]) ? node17688 : node17683;
													assign node17683 = (inp[4]) ? node17685 : 4'b0101;
														assign node17685 = (inp[9]) ? 4'b0101 : 4'b0001;
													assign node17688 = (inp[10]) ? 4'b0000 : node17689;
														assign node17689 = (inp[9]) ? 4'b0000 : 4'b0100;
										assign node17693 = (inp[7]) ? node17719 : node17694;
											assign node17694 = (inp[8]) ? node17706 : node17695;
												assign node17695 = (inp[2]) ? node17701 : node17696;
													assign node17696 = (inp[4]) ? node17698 : 4'b0100;
														assign node17698 = (inp[10]) ? 4'b0001 : 4'b0101;
													assign node17701 = (inp[9]) ? 4'b0100 : node17702;
														assign node17702 = (inp[10]) ? 4'b0100 : 4'b0000;
												assign node17706 = (inp[14]) ? node17712 : node17707;
													assign node17707 = (inp[10]) ? node17709 : 4'b0001;
														assign node17709 = (inp[4]) ? 4'b0101 : 4'b0100;
													assign node17712 = (inp[10]) ? node17716 : node17713;
														assign node17713 = (inp[4]) ? 4'b0101 : 4'b0001;
														assign node17716 = (inp[4]) ? 4'b0001 : 4'b0001;
											assign node17719 = (inp[8]) ? node17733 : node17720;
												assign node17720 = (inp[2]) ? node17728 : node17721;
													assign node17721 = (inp[14]) ? node17725 : node17722;
														assign node17722 = (inp[4]) ? 4'b0000 : 4'b0100;
														assign node17725 = (inp[4]) ? 4'b0001 : 4'b0101;
													assign node17728 = (inp[14]) ? 4'b0001 : node17729;
														assign node17729 = (inp[4]) ? 4'b0101 : 4'b0001;
												assign node17733 = (inp[14]) ? 4'b0100 : node17734;
													assign node17734 = (inp[2]) ? node17738 : node17735;
														assign node17735 = (inp[10]) ? 4'b0101 : 4'b0001;
														assign node17738 = (inp[4]) ? 4'b0000 : 4'b0100;
						assign node17742 = (inp[7]) ? node18092 : node17743;
							assign node17743 = (inp[8]) ? node17915 : node17744;
								assign node17744 = (inp[14]) ? node17828 : node17745;
									assign node17745 = (inp[2]) ? node17783 : node17746;
										assign node17746 = (inp[15]) ? node17768 : node17747;
											assign node17747 = (inp[5]) ? node17761 : node17748;
												assign node17748 = (inp[3]) ? node17756 : node17749;
													assign node17749 = (inp[9]) ? node17753 : node17750;
														assign node17750 = (inp[4]) ? 4'b0001 : 4'b0101;
														assign node17753 = (inp[4]) ? 4'b0101 : 4'b0001;
													assign node17756 = (inp[12]) ? 4'b0111 : node17757;
														assign node17757 = (inp[9]) ? 4'b0001 : 4'b0101;
												assign node17761 = (inp[12]) ? node17763 : 4'b0111;
													assign node17763 = (inp[4]) ? 4'b0011 : node17764;
														assign node17764 = (inp[3]) ? 4'b0011 : 4'b0111;
											assign node17768 = (inp[5]) ? node17776 : node17769;
												assign node17769 = (inp[10]) ? node17771 : 4'b0111;
													assign node17771 = (inp[3]) ? 4'b0011 : node17772;
														assign node17772 = (inp[9]) ? 4'b0111 : 4'b0011;
												assign node17776 = (inp[3]) ? node17778 : 4'b0011;
													assign node17778 = (inp[10]) ? node17780 : 4'b0101;
														assign node17780 = (inp[9]) ? 4'b0001 : 4'b0001;
										assign node17783 = (inp[9]) ? node17809 : node17784;
											assign node17784 = (inp[4]) ? node17796 : node17785;
												assign node17785 = (inp[12]) ? node17791 : node17786;
													assign node17786 = (inp[5]) ? node17788 : 4'b0110;
														assign node17788 = (inp[3]) ? 4'b0100 : 4'b0110;
													assign node17791 = (inp[10]) ? node17793 : 4'b0100;
														assign node17793 = (inp[15]) ? 4'b0010 : 4'b0000;
												assign node17796 = (inp[12]) ? node17802 : node17797;
													assign node17797 = (inp[3]) ? node17799 : 4'b0000;
														assign node17799 = (inp[15]) ? 4'b0000 : 4'b0010;
													assign node17802 = (inp[10]) ? node17806 : node17803;
														assign node17803 = (inp[15]) ? 4'b0000 : 4'b0000;
														assign node17806 = (inp[5]) ? 4'b0100 : 4'b0110;
											assign node17809 = (inp[3]) ? node17821 : node17810;
												assign node17810 = (inp[12]) ? node17816 : node17811;
													assign node17811 = (inp[4]) ? node17813 : 4'b0010;
														assign node17813 = (inp[15]) ? 4'b0100 : 4'b0100;
													assign node17816 = (inp[4]) ? node17818 : 4'b0110;
														assign node17818 = (inp[10]) ? 4'b0010 : 4'b0110;
												assign node17821 = (inp[15]) ? 4'b0100 : node17822;
													assign node17822 = (inp[5]) ? node17824 : 4'b0000;
														assign node17824 = (inp[4]) ? 4'b0110 : 4'b0010;
									assign node17828 = (inp[15]) ? node17870 : node17829;
										assign node17829 = (inp[3]) ? node17849 : node17830;
											assign node17830 = (inp[2]) ? node17840 : node17831;
												assign node17831 = (inp[4]) ? node17837 : node17832;
													assign node17832 = (inp[9]) ? 4'b0000 : node17833;
														assign node17833 = (inp[12]) ? 4'b0000 : 4'b0100;
													assign node17837 = (inp[9]) ? 4'b0100 : 4'b0000;
												assign node17840 = (inp[12]) ? node17842 : 4'b0100;
													assign node17842 = (inp[9]) ? node17846 : node17843;
														assign node17843 = (inp[5]) ? 4'b0000 : 4'b0100;
														assign node17846 = (inp[5]) ? 4'b0110 : 4'b0000;
											assign node17849 = (inp[5]) ? node17861 : node17850;
												assign node17850 = (inp[9]) ? node17856 : node17851;
													assign node17851 = (inp[2]) ? node17853 : 4'b0000;
														assign node17853 = (inp[4]) ? 4'b0110 : 4'b0000;
													assign node17856 = (inp[4]) ? 4'b0110 : node17857;
														assign node17857 = (inp[10]) ? 4'b0110 : 4'b0000;
												assign node17861 = (inp[12]) ? 4'b0110 : node17862;
													assign node17862 = (inp[4]) ? node17866 : node17863;
														assign node17863 = (inp[9]) ? 4'b0010 : 4'b0110;
														assign node17866 = (inp[9]) ? 4'b0110 : 4'b0010;
										assign node17870 = (inp[3]) ? node17896 : node17871;
											assign node17871 = (inp[5]) ? node17883 : node17872;
												assign node17872 = (inp[10]) ? node17878 : node17873;
													assign node17873 = (inp[4]) ? node17875 : 4'b0110;
														assign node17875 = (inp[9]) ? 4'b0110 : 4'b0010;
													assign node17878 = (inp[9]) ? 4'b0010 : node17879;
														assign node17879 = (inp[2]) ? 4'b0110 : 4'b0010;
												assign node17883 = (inp[9]) ? node17889 : node17884;
													assign node17884 = (inp[2]) ? node17886 : 4'b0010;
														assign node17886 = (inp[4]) ? 4'b0100 : 4'b0010;
													assign node17889 = (inp[4]) ? node17893 : node17890;
														assign node17890 = (inp[10]) ? 4'b0000 : 4'b0010;
														assign node17893 = (inp[10]) ? 4'b0000 : 4'b0100;
											assign node17896 = (inp[5]) ? node17908 : node17897;
												assign node17897 = (inp[4]) ? node17903 : node17898;
													assign node17898 = (inp[10]) ? 4'b0010 : node17899;
														assign node17899 = (inp[9]) ? 4'b0010 : 4'b0110;
													assign node17903 = (inp[10]) ? node17905 : 4'b0100;
														assign node17905 = (inp[12]) ? 4'b0000 : 4'b0010;
												assign node17908 = (inp[10]) ? node17910 : 4'b0000;
													assign node17910 = (inp[9]) ? node17912 : 4'b0100;
														assign node17912 = (inp[4]) ? 4'b0100 : 4'b0000;
								assign node17915 = (inp[2]) ? node18011 : node17916;
									assign node17916 = (inp[14]) ? node17962 : node17917;
										assign node17917 = (inp[15]) ? node17939 : node17918;
											assign node17918 = (inp[5]) ? node17930 : node17919;
												assign node17919 = (inp[3]) ? node17925 : node17920;
													assign node17920 = (inp[4]) ? node17922 : 4'b0100;
														assign node17922 = (inp[9]) ? 4'b0100 : 4'b0000;
													assign node17925 = (inp[4]) ? 4'b0110 : node17926;
														assign node17926 = (inp[9]) ? 4'b0000 : 4'b0100;
												assign node17930 = (inp[12]) ? node17934 : node17931;
													assign node17931 = (inp[3]) ? 4'b0010 : 4'b0000;
													assign node17934 = (inp[4]) ? node17936 : 4'b0110;
														assign node17936 = (inp[3]) ? 4'b0010 : 4'b0110;
											assign node17939 = (inp[9]) ? node17951 : node17940;
												assign node17940 = (inp[5]) ? node17944 : node17941;
													assign node17941 = (inp[4]) ? 4'b0010 : 4'b0110;
													assign node17944 = (inp[3]) ? node17948 : node17945;
														assign node17945 = (inp[4]) ? 4'b0000 : 4'b0010;
														assign node17948 = (inp[4]) ? 4'b0000 : 4'b0100;
												assign node17951 = (inp[4]) ? node17959 : node17952;
													assign node17952 = (inp[12]) ? node17956 : node17953;
														assign node17953 = (inp[5]) ? 4'b0000 : 4'b0010;
														assign node17956 = (inp[10]) ? 4'b0100 : 4'b0000;
													assign node17959 = (inp[12]) ? 4'b0000 : 4'b0100;
										assign node17962 = (inp[12]) ? node17984 : node17963;
											assign node17963 = (inp[15]) ? node17977 : node17964;
												assign node17964 = (inp[4]) ? node17970 : node17965;
													assign node17965 = (inp[10]) ? node17967 : 4'b1001;
														assign node17967 = (inp[9]) ? 4'b1111 : 4'b1001;
													assign node17970 = (inp[3]) ? node17974 : node17971;
														assign node17971 = (inp[5]) ? 4'b1011 : 4'b1001;
														assign node17974 = (inp[10]) ? 4'b1011 : 4'b1111;
												assign node17977 = (inp[3]) ? 4'b1011 : node17978;
													assign node17978 = (inp[5]) ? node17980 : 4'b1111;
														assign node17980 = (inp[10]) ? 4'b1011 : 4'b1011;
											assign node17984 = (inp[15]) ? node17998 : node17985;
												assign node17985 = (inp[5]) ? node17993 : node17986;
													assign node17986 = (inp[3]) ? node17990 : node17987;
														assign node17987 = (inp[10]) ? 4'b1001 : 4'b1101;
														assign node17990 = (inp[10]) ? 4'b1001 : 4'b1011;
													assign node17993 = (inp[4]) ? node17995 : 4'b1011;
														assign node17995 = (inp[9]) ? 4'b1011 : 4'b1111;
												assign node17998 = (inp[3]) ? node18004 : node17999;
													assign node17999 = (inp[4]) ? node18001 : 4'b1011;
														assign node18001 = (inp[10]) ? 4'b1001 : 4'b1111;
													assign node18004 = (inp[5]) ? node18008 : node18005;
														assign node18005 = (inp[9]) ? 4'b1001 : 4'b1101;
														assign node18008 = (inp[9]) ? 4'b1101 : 4'b1001;
									assign node18011 = (inp[10]) ? node18053 : node18012;
										assign node18012 = (inp[9]) ? node18036 : node18013;
											assign node18013 = (inp[15]) ? node18023 : node18014;
												assign node18014 = (inp[12]) ? node18018 : node18015;
													assign node18015 = (inp[4]) ? 4'b1001 : 4'b1101;
													assign node18018 = (inp[4]) ? node18020 : 4'b1001;
														assign node18020 = (inp[14]) ? 4'b1111 : 4'b1101;
												assign node18023 = (inp[14]) ? node18031 : node18024;
													assign node18024 = (inp[12]) ? node18028 : node18025;
														assign node18025 = (inp[4]) ? 4'b1011 : 4'b1111;
														assign node18028 = (inp[4]) ? 4'b1111 : 4'b1011;
													assign node18031 = (inp[3]) ? 4'b1101 : node18032;
														assign node18032 = (inp[5]) ? 4'b1011 : 4'b1111;
											assign node18036 = (inp[3]) ? node18050 : node18037;
												assign node18037 = (inp[4]) ? node18043 : node18038;
													assign node18038 = (inp[14]) ? 4'b1001 : node18039;
														assign node18039 = (inp[15]) ? 4'b1101 : 4'b1111;
													assign node18043 = (inp[12]) ? node18047 : node18044;
														assign node18044 = (inp[15]) ? 4'b1111 : 4'b1101;
														assign node18047 = (inp[15]) ? 4'b1001 : 4'b1001;
												assign node18050 = (inp[15]) ? 4'b1101 : 4'b1111;
										assign node18053 = (inp[15]) ? node18071 : node18054;
											assign node18054 = (inp[4]) ? node18064 : node18055;
												assign node18055 = (inp[9]) ? node18061 : node18056;
													assign node18056 = (inp[14]) ? node18058 : 4'b1001;
														assign node18058 = (inp[3]) ? 4'b1001 : 4'b1001;
													assign node18061 = (inp[5]) ? 4'b1111 : 4'b1101;
												assign node18064 = (inp[9]) ? 4'b1011 : node18065;
													assign node18065 = (inp[5]) ? 4'b1111 : node18066;
														assign node18066 = (inp[3]) ? 4'b1111 : 4'b1101;
											assign node18071 = (inp[3]) ? node18085 : node18072;
												assign node18072 = (inp[5]) ? node18080 : node18073;
													assign node18073 = (inp[9]) ? node18077 : node18074;
														assign node18074 = (inp[4]) ? 4'b1111 : 4'b1011;
														assign node18077 = (inp[12]) ? 4'b1011 : 4'b1111;
													assign node18080 = (inp[4]) ? node18082 : 4'b1011;
														assign node18082 = (inp[9]) ? 4'b1001 : 4'b1101;
												assign node18085 = (inp[9]) ? node18089 : node18086;
													assign node18086 = (inp[4]) ? 4'b1101 : 4'b1001;
													assign node18089 = (inp[4]) ? 4'b1001 : 4'b1101;
							assign node18092 = (inp[8]) ? node18268 : node18093;
								assign node18093 = (inp[14]) ? node18183 : node18094;
									assign node18094 = (inp[2]) ? node18142 : node18095;
										assign node18095 = (inp[9]) ? node18123 : node18096;
											assign node18096 = (inp[15]) ? node18110 : node18097;
												assign node18097 = (inp[5]) ? node18105 : node18098;
													assign node18098 = (inp[10]) ? node18102 : node18099;
														assign node18099 = (inp[4]) ? 4'b0000 : 4'b0100;
														assign node18102 = (inp[3]) ? 4'b0000 : 4'b0100;
													assign node18105 = (inp[3]) ? node18107 : 4'b0000;
														assign node18107 = (inp[4]) ? 4'b0010 : 4'b0110;
												assign node18110 = (inp[3]) ? node18118 : node18111;
													assign node18111 = (inp[12]) ? node18115 : node18112;
														assign node18112 = (inp[4]) ? 4'b0010 : 4'b0110;
														assign node18115 = (inp[4]) ? 4'b0110 : 4'b0010;
													assign node18118 = (inp[12]) ? node18120 : 4'b0110;
														assign node18120 = (inp[10]) ? 4'b0000 : 4'b0100;
											assign node18123 = (inp[10]) ? node18131 : node18124;
												assign node18124 = (inp[3]) ? 4'b0110 : node18125;
													assign node18125 = (inp[12]) ? node18127 : 4'b0100;
														assign node18127 = (inp[5]) ? 4'b0110 : 4'b0100;
												assign node18131 = (inp[12]) ? node18137 : node18132;
													assign node18132 = (inp[4]) ? node18134 : 4'b0010;
														assign node18134 = (inp[5]) ? 4'b0100 : 4'b0110;
													assign node18137 = (inp[4]) ? node18139 : 4'b0100;
														assign node18139 = (inp[15]) ? 4'b0000 : 4'b0010;
										assign node18142 = (inp[3]) ? node18168 : node18143;
											assign node18143 = (inp[4]) ? node18157 : node18144;
												assign node18144 = (inp[12]) ? node18150 : node18145;
													assign node18145 = (inp[5]) ? 4'b1111 : node18146;
														assign node18146 = (inp[10]) ? 4'b1111 : 4'b1011;
													assign node18150 = (inp[9]) ? node18154 : node18151;
														assign node18151 = (inp[5]) ? 4'b1011 : 4'b1001;
														assign node18154 = (inp[5]) ? 4'b1101 : 4'b1111;
												assign node18157 = (inp[9]) ? node18163 : node18158;
													assign node18158 = (inp[10]) ? node18160 : 4'b1001;
														assign node18160 = (inp[15]) ? 4'b1101 : 4'b1111;
													assign node18163 = (inp[5]) ? node18165 : 4'b1011;
														assign node18165 = (inp[15]) ? 4'b1001 : 4'b1011;
											assign node18168 = (inp[15]) ? node18176 : node18169;
												assign node18169 = (inp[5]) ? 4'b1111 : node18170;
													assign node18170 = (inp[12]) ? node18172 : 4'b1001;
														assign node18172 = (inp[4]) ? 4'b1011 : 4'b1111;
												assign node18176 = (inp[5]) ? 4'b1001 : node18177;
													assign node18177 = (inp[4]) ? 4'b1001 : node18178;
														assign node18178 = (inp[12]) ? 4'b1011 : 4'b1111;
									assign node18183 = (inp[15]) ? node18227 : node18184;
										assign node18184 = (inp[3]) ? node18210 : node18185;
											assign node18185 = (inp[5]) ? node18197 : node18186;
												assign node18186 = (inp[12]) ? node18192 : node18187;
													assign node18187 = (inp[10]) ? node18189 : 4'b1101;
														assign node18189 = (inp[4]) ? 4'b1001 : 4'b1101;
													assign node18192 = (inp[4]) ? node18194 : 4'b1001;
														assign node18194 = (inp[9]) ? 4'b1001 : 4'b1101;
												assign node18197 = (inp[9]) ? node18205 : node18198;
													assign node18198 = (inp[4]) ? node18202 : node18199;
														assign node18199 = (inp[10]) ? 4'b1001 : 4'b1001;
														assign node18202 = (inp[12]) ? 4'b1111 : 4'b1001;
													assign node18205 = (inp[2]) ? 4'b1001 : node18206;
														assign node18206 = (inp[12]) ? 4'b1011 : 4'b1111;
											assign node18210 = (inp[10]) ? node18218 : node18211;
												assign node18211 = (inp[5]) ? node18213 : 4'b1001;
													assign node18213 = (inp[9]) ? node18215 : 4'b1011;
														assign node18215 = (inp[4]) ? 4'b1011 : 4'b1011;
												assign node18218 = (inp[9]) ? node18224 : node18219;
													assign node18219 = (inp[4]) ? 4'b1111 : node18220;
														assign node18220 = (inp[2]) ? 4'b1001 : 4'b1011;
													assign node18224 = (inp[4]) ? 4'b1011 : 4'b1111;
										assign node18227 = (inp[3]) ? node18249 : node18228;
											assign node18228 = (inp[5]) ? node18236 : node18229;
												assign node18229 = (inp[4]) ? 4'b1011 : node18230;
													assign node18230 = (inp[10]) ? 4'b1111 : node18231;
														assign node18231 = (inp[9]) ? 4'b1011 : 4'b1111;
												assign node18236 = (inp[9]) ? node18242 : node18237;
													assign node18237 = (inp[2]) ? node18239 : 4'b1011;
														assign node18239 = (inp[4]) ? 4'b1001 : 4'b1011;
													assign node18242 = (inp[12]) ? node18246 : node18243;
														assign node18243 = (inp[2]) ? 4'b1101 : 4'b1011;
														assign node18246 = (inp[4]) ? 4'b1001 : 4'b1101;
											assign node18249 = (inp[4]) ? node18261 : node18250;
												assign node18250 = (inp[5]) ? node18256 : node18251;
													assign node18251 = (inp[12]) ? 4'b1011 : node18252;
														assign node18252 = (inp[10]) ? 4'b1011 : 4'b1111;
													assign node18256 = (inp[10]) ? 4'b1001 : node18257;
														assign node18257 = (inp[12]) ? 4'b1101 : 4'b1001;
												assign node18261 = (inp[9]) ? node18263 : 4'b1101;
													assign node18263 = (inp[10]) ? 4'b1001 : node18264;
														assign node18264 = (inp[12]) ? 4'b1001 : 4'b1101;
								assign node18268 = (inp[14]) ? node18356 : node18269;
									assign node18269 = (inp[2]) ? node18315 : node18270;
										assign node18270 = (inp[5]) ? node18296 : node18271;
											assign node18271 = (inp[15]) ? node18283 : node18272;
												assign node18272 = (inp[3]) ? node18278 : node18273;
													assign node18273 = (inp[4]) ? 4'b1101 : node18274;
														assign node18274 = (inp[10]) ? 4'b1101 : 4'b1001;
													assign node18278 = (inp[4]) ? 4'b1111 : node18279;
														assign node18279 = (inp[10]) ? 4'b1111 : 4'b1001;
												assign node18283 = (inp[3]) ? node18289 : node18284;
													assign node18284 = (inp[4]) ? node18286 : 4'b1011;
														assign node18286 = (inp[9]) ? 4'b1011 : 4'b1111;
													assign node18289 = (inp[12]) ? node18293 : node18290;
														assign node18290 = (inp[9]) ? 4'b1011 : 4'b1111;
														assign node18293 = (inp[9]) ? 4'b1101 : 4'b1011;
											assign node18296 = (inp[15]) ? node18304 : node18297;
												assign node18297 = (inp[9]) ? 4'b1011 : node18298;
													assign node18298 = (inp[4]) ? 4'b1011 : node18299;
														assign node18299 = (inp[12]) ? 4'b1001 : 4'b1101;
												assign node18304 = (inp[4]) ? node18310 : node18305;
													assign node18305 = (inp[9]) ? 4'b1101 : node18306;
														assign node18306 = (inp[10]) ? 4'b1011 : 4'b1101;
													assign node18310 = (inp[3]) ? 4'b1001 : node18311;
														assign node18311 = (inp[9]) ? 4'b1001 : 4'b1101;
										assign node18315 = (inp[4]) ? node18337 : node18316;
											assign node18316 = (inp[9]) ? node18328 : node18317;
												assign node18317 = (inp[15]) ? node18323 : node18318;
													assign node18318 = (inp[5]) ? node18320 : 4'b1000;
														assign node18320 = (inp[3]) ? 4'b1010 : 4'b1000;
													assign node18323 = (inp[12]) ? 4'b1010 : node18324;
														assign node18324 = (inp[10]) ? 4'b1000 : 4'b1110;
												assign node18328 = (inp[12]) ? node18332 : node18329;
													assign node18329 = (inp[10]) ? 4'b1110 : 4'b1010;
													assign node18332 = (inp[15]) ? node18334 : 4'b1110;
														assign node18334 = (inp[3]) ? 4'b1100 : 4'b1100;
											assign node18337 = (inp[15]) ? node18345 : node18338;
												assign node18338 = (inp[12]) ? node18340 : 4'b1110;
													assign node18340 = (inp[9]) ? node18342 : 4'b1110;
														assign node18342 = (inp[5]) ? 4'b1010 : 4'b1000;
												assign node18345 = (inp[9]) ? node18351 : node18346;
													assign node18346 = (inp[10]) ? 4'b1100 : node18347;
														assign node18347 = (inp[12]) ? 4'b1100 : 4'b1000;
													assign node18351 = (inp[12]) ? 4'b1000 : node18352;
														assign node18352 = (inp[10]) ? 4'b1000 : 4'b1100;
									assign node18356 = (inp[10]) ? node18406 : node18357;
										assign node18357 = (inp[5]) ? node18383 : node18358;
											assign node18358 = (inp[15]) ? node18370 : node18359;
												assign node18359 = (inp[4]) ? node18365 : node18360;
													assign node18360 = (inp[2]) ? 4'b1100 : node18361;
														assign node18361 = (inp[12]) ? 4'b1000 : 4'b1000;
													assign node18365 = (inp[9]) ? node18367 : 4'b1000;
														assign node18367 = (inp[2]) ? 4'b1000 : 4'b1100;
												assign node18370 = (inp[3]) ? node18378 : node18371;
													assign node18371 = (inp[4]) ? node18375 : node18372;
														assign node18372 = (inp[2]) ? 4'b1110 : 4'b1010;
														assign node18375 = (inp[2]) ? 4'b1010 : 4'b1010;
													assign node18378 = (inp[4]) ? node18380 : 4'b1010;
														assign node18380 = (inp[12]) ? 4'b1100 : 4'b1000;
											assign node18383 = (inp[15]) ? node18395 : node18384;
												assign node18384 = (inp[3]) ? node18390 : node18385;
													assign node18385 = (inp[9]) ? node18387 : 4'b1000;
														assign node18387 = (inp[4]) ? 4'b1110 : 4'b1000;
													assign node18390 = (inp[2]) ? 4'b1010 : node18391;
														assign node18391 = (inp[9]) ? 4'b1110 : 4'b1010;
												assign node18395 = (inp[9]) ? node18401 : node18396;
													assign node18396 = (inp[2]) ? 4'b1010 : node18397;
														assign node18397 = (inp[12]) ? 4'b1100 : 4'b1010;
													assign node18401 = (inp[2]) ? 4'b1000 : node18402;
														assign node18402 = (inp[4]) ? 4'b1000 : 4'b1100;
										assign node18406 = (inp[15]) ? node18422 : node18407;
											assign node18407 = (inp[5]) ? node18413 : node18408;
												assign node18408 = (inp[4]) ? node18410 : 4'b1000;
													assign node18410 = (inp[9]) ? 4'b1010 : 4'b1110;
												assign node18413 = (inp[2]) ? node18415 : 4'b1110;
													assign node18415 = (inp[9]) ? node18419 : node18416;
														assign node18416 = (inp[4]) ? 4'b1110 : 4'b1000;
														assign node18419 = (inp[4]) ? 4'b1010 : 4'b1110;
											assign node18422 = (inp[5]) ? node18432 : node18423;
												assign node18423 = (inp[3]) ? node18429 : node18424;
													assign node18424 = (inp[2]) ? node18426 : 4'b1110;
														assign node18426 = (inp[9]) ? 4'b1110 : 4'b1010;
													assign node18429 = (inp[4]) ? 4'b1000 : 4'b1010;
												assign node18432 = (inp[3]) ? node18438 : node18433;
													assign node18433 = (inp[2]) ? 4'b1010 : node18434;
														assign node18434 = (inp[9]) ? 4'b1000 : 4'b1100;
													assign node18438 = (inp[12]) ? 4'b1100 : node18439;
														assign node18439 = (inp[9]) ? 4'b1100 : 4'b1000;
					assign node18443 = (inp[13]) ? node19173 : node18444;
						assign node18444 = (inp[7]) ? node18788 : node18445;
							assign node18445 = (inp[8]) ? node18629 : node18446;
								assign node18446 = (inp[2]) ? node18528 : node18447;
									assign node18447 = (inp[14]) ? node18487 : node18448;
										assign node18448 = (inp[5]) ? node18468 : node18449;
											assign node18449 = (inp[15]) ? node18459 : node18450;
												assign node18450 = (inp[12]) ? node18452 : 4'b0101;
													assign node18452 = (inp[4]) ? node18456 : node18453;
														assign node18453 = (inp[10]) ? 4'b0001 : 4'b0001;
														assign node18456 = (inp[3]) ? 4'b0001 : 4'b0101;
												assign node18459 = (inp[12]) ? node18465 : node18460;
													assign node18460 = (inp[4]) ? 4'b0011 : node18461;
														assign node18461 = (inp[9]) ? 4'b0011 : 4'b0111;
													assign node18465 = (inp[10]) ? 4'b0101 : 4'b0111;
											assign node18468 = (inp[15]) ? node18476 : node18469;
												assign node18469 = (inp[9]) ? node18471 : 4'b0011;
													assign node18471 = (inp[12]) ? node18473 : 4'b0111;
														assign node18473 = (inp[4]) ? 4'b0011 : 4'b0011;
												assign node18476 = (inp[3]) ? node18482 : node18477;
													assign node18477 = (inp[4]) ? node18479 : 4'b0011;
														assign node18479 = (inp[9]) ? 4'b0101 : 4'b0011;
													assign node18482 = (inp[10]) ? node18484 : 4'b0001;
														assign node18484 = (inp[12]) ? 4'b0001 : 4'b0101;
										assign node18487 = (inp[4]) ? node18511 : node18488;
											assign node18488 = (inp[9]) ? node18500 : node18489;
												assign node18489 = (inp[15]) ? node18495 : node18490;
													assign node18490 = (inp[5]) ? 4'b0010 : node18491;
														assign node18491 = (inp[12]) ? 4'b0000 : 4'b0100;
													assign node18495 = (inp[3]) ? node18497 : 4'b0110;
														assign node18497 = (inp[10]) ? 4'b0110 : 4'b0100;
												assign node18500 = (inp[10]) ? node18506 : node18501;
													assign node18501 = (inp[5]) ? node18503 : 4'b0010;
														assign node18503 = (inp[15]) ? 4'b0000 : 4'b0000;
													assign node18506 = (inp[12]) ? 4'b0100 : node18507;
														assign node18507 = (inp[15]) ? 4'b0000 : 4'b0000;
											assign node18511 = (inp[9]) ? node18519 : node18512;
												assign node18512 = (inp[10]) ? node18514 : 4'b0000;
													assign node18514 = (inp[12]) ? node18516 : 4'b0010;
														assign node18516 = (inp[5]) ? 4'b0110 : 4'b0100;
												assign node18519 = (inp[12]) ? node18525 : node18520;
													assign node18520 = (inp[15]) ? 4'b0100 : node18521;
														assign node18521 = (inp[3]) ? 4'b0110 : 4'b0100;
													assign node18525 = (inp[10]) ? 4'b0000 : 4'b0100;
									assign node18528 = (inp[14]) ? node18578 : node18529;
										assign node18529 = (inp[9]) ? node18555 : node18530;
											assign node18530 = (inp[4]) ? node18542 : node18531;
												assign node18531 = (inp[10]) ? node18537 : node18532;
													assign node18532 = (inp[15]) ? node18534 : 4'b0100;
														assign node18534 = (inp[12]) ? 4'b0110 : 4'b0100;
													assign node18537 = (inp[12]) ? node18539 : 4'b0100;
														assign node18539 = (inp[5]) ? 4'b0000 : 4'b0000;
												assign node18542 = (inp[3]) ? node18550 : node18543;
													assign node18543 = (inp[10]) ? node18547 : node18544;
														assign node18544 = (inp[15]) ? 4'b0010 : 4'b0000;
														assign node18547 = (inp[15]) ? 4'b0010 : 4'b0110;
													assign node18550 = (inp[12]) ? node18552 : 4'b0000;
														assign node18552 = (inp[10]) ? 4'b0100 : 4'b0000;
											assign node18555 = (inp[3]) ? node18563 : node18556;
												assign node18556 = (inp[12]) ? node18560 : node18557;
													assign node18557 = (inp[4]) ? 4'b0110 : 4'b0010;
													assign node18560 = (inp[4]) ? 4'b0010 : 4'b0110;
												assign node18563 = (inp[4]) ? node18571 : node18564;
													assign node18564 = (inp[12]) ? node18568 : node18565;
														assign node18565 = (inp[15]) ? 4'b0010 : 4'b0000;
														assign node18568 = (inp[5]) ? 4'b0100 : 4'b0010;
													assign node18571 = (inp[15]) ? node18575 : node18572;
														assign node18572 = (inp[12]) ? 4'b0010 : 4'b0110;
														assign node18575 = (inp[10]) ? 4'b0000 : 4'b0100;
										assign node18578 = (inp[5]) ? node18604 : node18579;
											assign node18579 = (inp[15]) ? node18591 : node18580;
												assign node18580 = (inp[3]) ? node18586 : node18581;
													assign node18581 = (inp[4]) ? 4'b0100 : node18582;
														assign node18582 = (inp[9]) ? 4'b0000 : 4'b0100;
													assign node18586 = (inp[12]) ? node18588 : 4'b0000;
														assign node18588 = (inp[4]) ? 4'b0010 : 4'b0110;
												assign node18591 = (inp[10]) ? node18599 : node18592;
													assign node18592 = (inp[9]) ? node18596 : node18593;
														assign node18593 = (inp[4]) ? 4'b0010 : 4'b0110;
														assign node18596 = (inp[4]) ? 4'b0100 : 4'b0010;
													assign node18599 = (inp[9]) ? node18601 : 4'b0110;
														assign node18601 = (inp[4]) ? 4'b0110 : 4'b0010;
											assign node18604 = (inp[15]) ? node18618 : node18605;
												assign node18605 = (inp[3]) ? node18613 : node18606;
													assign node18606 = (inp[4]) ? node18610 : node18607;
														assign node18607 = (inp[10]) ? 4'b0000 : 4'b0100;
														assign node18610 = (inp[10]) ? 4'b0110 : 4'b0000;
													assign node18613 = (inp[12]) ? 4'b0110 : node18614;
														assign node18614 = (inp[4]) ? 4'b0110 : 4'b0010;
												assign node18618 = (inp[3]) ? node18622 : node18619;
													assign node18619 = (inp[4]) ? 4'b0100 : 4'b0110;
													assign node18622 = (inp[9]) ? node18626 : node18623;
														assign node18623 = (inp[4]) ? 4'b0000 : 4'b0000;
														assign node18626 = (inp[4]) ? 4'b0100 : 4'b0000;
								assign node18629 = (inp[2]) ? node18713 : node18630;
									assign node18630 = (inp[14]) ? node18682 : node18631;
										assign node18631 = (inp[12]) ? node18655 : node18632;
											assign node18632 = (inp[5]) ? node18642 : node18633;
												assign node18633 = (inp[15]) ? node18639 : node18634;
													assign node18634 = (inp[9]) ? 4'b0100 : node18635;
														assign node18635 = (inp[4]) ? 4'b0000 : 4'b0100;
													assign node18639 = (inp[3]) ? 4'b0110 : 4'b0010;
												assign node18642 = (inp[15]) ? node18650 : node18643;
													assign node18643 = (inp[4]) ? node18647 : node18644;
														assign node18644 = (inp[3]) ? 4'b0110 : 4'b0100;
														assign node18647 = (inp[9]) ? 4'b0110 : 4'b0010;
													assign node18650 = (inp[9]) ? 4'b0100 : node18651;
														assign node18651 = (inp[3]) ? 4'b0100 : 4'b0110;
											assign node18655 = (inp[4]) ? node18671 : node18656;
												assign node18656 = (inp[10]) ? node18664 : node18657;
													assign node18657 = (inp[9]) ? node18661 : node18658;
														assign node18658 = (inp[5]) ? 4'b0100 : 4'b0100;
														assign node18661 = (inp[15]) ? 4'b0010 : 4'b0000;
													assign node18664 = (inp[9]) ? node18668 : node18665;
														assign node18665 = (inp[5]) ? 4'b0010 : 4'b0000;
														assign node18668 = (inp[3]) ? 4'b0110 : 4'b0100;
												assign node18671 = (inp[10]) ? node18677 : node18672;
													assign node18672 = (inp[9]) ? 4'b0110 : node18673;
														assign node18673 = (inp[5]) ? 4'b0010 : 4'b0010;
													assign node18677 = (inp[9]) ? node18679 : 4'b0100;
														assign node18679 = (inp[3]) ? 4'b0010 : 4'b0000;
										assign node18682 = (inp[15]) ? node18698 : node18683;
											assign node18683 = (inp[4]) ? node18691 : node18684;
												assign node18684 = (inp[9]) ? node18686 : 4'b1001;
													assign node18686 = (inp[10]) ? 4'b1111 : node18687;
														assign node18687 = (inp[3]) ? 4'b1011 : 4'b1001;
												assign node18691 = (inp[9]) ? 4'b1011 : node18692;
													assign node18692 = (inp[5]) ? 4'b1111 : node18693;
														assign node18693 = (inp[3]) ? 4'b1111 : 4'b1001;
											assign node18698 = (inp[4]) ? node18706 : node18699;
												assign node18699 = (inp[9]) ? node18701 : 4'b1011;
													assign node18701 = (inp[5]) ? 4'b1101 : node18702;
														assign node18702 = (inp[10]) ? 4'b1111 : 4'b1101;
												assign node18706 = (inp[9]) ? node18708 : 4'b1101;
													assign node18708 = (inp[12]) ? node18710 : 4'b1101;
														assign node18710 = (inp[5]) ? 4'b1001 : 4'b1011;
									assign node18713 = (inp[10]) ? node18749 : node18714;
										assign node18714 = (inp[12]) ? node18732 : node18715;
											assign node18715 = (inp[15]) ? node18723 : node18716;
												assign node18716 = (inp[5]) ? 4'b1111 : node18717;
													assign node18717 = (inp[4]) ? node18719 : 4'b1001;
														assign node18719 = (inp[3]) ? 4'b1111 : 4'b1101;
												assign node18723 = (inp[9]) ? node18729 : node18724;
													assign node18724 = (inp[4]) ? 4'b1011 : node18725;
														assign node18725 = (inp[3]) ? 4'b1111 : 4'b1111;
													assign node18729 = (inp[4]) ? 4'b1101 : 4'b1011;
											assign node18732 = (inp[9]) ? node18740 : node18733;
												assign node18733 = (inp[4]) ? 4'b1111 : node18734;
													assign node18734 = (inp[15]) ? 4'b1011 : node18735;
														assign node18735 = (inp[5]) ? 4'b1001 : 4'b1001;
												assign node18740 = (inp[4]) ? node18746 : node18741;
													assign node18741 = (inp[5]) ? 4'b1101 : node18742;
														assign node18742 = (inp[3]) ? 4'b1111 : 4'b1101;
													assign node18746 = (inp[3]) ? 4'b1001 : 4'b1011;
										assign node18749 = (inp[15]) ? node18769 : node18750;
											assign node18750 = (inp[3]) ? node18762 : node18751;
												assign node18751 = (inp[5]) ? node18757 : node18752;
													assign node18752 = (inp[9]) ? 4'b1101 : node18753;
														assign node18753 = (inp[4]) ? 4'b1101 : 4'b1001;
													assign node18757 = (inp[4]) ? node18759 : 4'b1001;
														assign node18759 = (inp[9]) ? 4'b1011 : 4'b1111;
												assign node18762 = (inp[9]) ? node18766 : node18763;
													assign node18763 = (inp[4]) ? 4'b1111 : 4'b1011;
													assign node18766 = (inp[4]) ? 4'b1011 : 4'b1111;
											assign node18769 = (inp[12]) ? node18781 : node18770;
												assign node18770 = (inp[5]) ? node18774 : node18771;
													assign node18771 = (inp[14]) ? 4'b1011 : 4'b1111;
													assign node18774 = (inp[4]) ? node18778 : node18775;
														assign node18775 = (inp[9]) ? 4'b1101 : 4'b1001;
														assign node18778 = (inp[9]) ? 4'b1001 : 4'b1101;
												assign node18781 = (inp[3]) ? 4'b1101 : node18782;
													assign node18782 = (inp[5]) ? node18784 : 4'b1111;
														assign node18784 = (inp[14]) ? 4'b1101 : 4'b1001;
							assign node18788 = (inp[8]) ? node18992 : node18789;
								assign node18789 = (inp[2]) ? node18899 : node18790;
									assign node18790 = (inp[14]) ? node18846 : node18791;
										assign node18791 = (inp[12]) ? node18817 : node18792;
											assign node18792 = (inp[5]) ? node18808 : node18793;
												assign node18793 = (inp[15]) ? node18801 : node18794;
													assign node18794 = (inp[9]) ? node18798 : node18795;
														assign node18795 = (inp[4]) ? 4'b0000 : 4'b0100;
														assign node18798 = (inp[3]) ? 4'b0110 : 4'b0000;
													assign node18801 = (inp[4]) ? node18805 : node18802;
														assign node18802 = (inp[9]) ? 4'b0010 : 4'b0110;
														assign node18805 = (inp[10]) ? 4'b0110 : 4'b0100;
												assign node18808 = (inp[10]) ? node18814 : node18809;
													assign node18809 = (inp[9]) ? 4'b0010 : node18810;
														assign node18810 = (inp[3]) ? 4'b0100 : 4'b0010;
													assign node18814 = (inp[3]) ? 4'b0000 : 4'b0100;
											assign node18817 = (inp[9]) ? node18833 : node18818;
												assign node18818 = (inp[5]) ? node18826 : node18819;
													assign node18819 = (inp[15]) ? node18823 : node18820;
														assign node18820 = (inp[4]) ? 4'b0100 : 4'b0000;
														assign node18823 = (inp[3]) ? 4'b0000 : 4'b0010;
													assign node18826 = (inp[4]) ? node18830 : node18827;
														assign node18827 = (inp[3]) ? 4'b0100 : 4'b0100;
														assign node18830 = (inp[15]) ? 4'b0100 : 4'b0110;
												assign node18833 = (inp[15]) ? node18839 : node18834;
													assign node18834 = (inp[3]) ? node18836 : 4'b0000;
														assign node18836 = (inp[4]) ? 4'b0010 : 4'b0010;
													assign node18839 = (inp[3]) ? node18843 : node18840;
														assign node18840 = (inp[10]) ? 4'b0110 : 4'b0010;
														assign node18843 = (inp[5]) ? 4'b0100 : 4'b0000;
										assign node18846 = (inp[4]) ? node18874 : node18847;
											assign node18847 = (inp[9]) ? node18861 : node18848;
												assign node18848 = (inp[10]) ? node18856 : node18849;
													assign node18849 = (inp[12]) ? node18853 : node18850;
														assign node18850 = (inp[3]) ? 4'b1101 : 4'b1111;
														assign node18853 = (inp[15]) ? 4'b1011 : 4'b1001;
													assign node18856 = (inp[3]) ? node18858 : 4'b1011;
														assign node18858 = (inp[12]) ? 4'b1001 : 4'b1001;
												assign node18861 = (inp[12]) ? node18869 : node18862;
													assign node18862 = (inp[10]) ? node18866 : node18863;
														assign node18863 = (inp[15]) ? 4'b1011 : 4'b1001;
														assign node18866 = (inp[3]) ? 4'b1101 : 4'b1111;
													assign node18869 = (inp[5]) ? 4'b1101 : node18870;
														assign node18870 = (inp[10]) ? 4'b1111 : 4'b1101;
											assign node18874 = (inp[9]) ? node18888 : node18875;
												assign node18875 = (inp[12]) ? node18883 : node18876;
													assign node18876 = (inp[10]) ? node18880 : node18877;
														assign node18877 = (inp[15]) ? 4'b1011 : 4'b1001;
														assign node18880 = (inp[3]) ? 4'b1111 : 4'b1101;
													assign node18883 = (inp[15]) ? 4'b1101 : node18884;
														assign node18884 = (inp[5]) ? 4'b1111 : 4'b1101;
												assign node18888 = (inp[10]) ? node18894 : node18889;
													assign node18889 = (inp[5]) ? 4'b1111 : node18890;
														assign node18890 = (inp[15]) ? 4'b1111 : 4'b1101;
													assign node18894 = (inp[15]) ? node18896 : 4'b1011;
														assign node18896 = (inp[3]) ? 4'b1001 : 4'b1011;
									assign node18899 = (inp[15]) ? node18945 : node18900;
										assign node18900 = (inp[3]) ? node18926 : node18901;
											assign node18901 = (inp[5]) ? node18915 : node18902;
												assign node18902 = (inp[14]) ? node18908 : node18903;
													assign node18903 = (inp[10]) ? node18905 : 4'b1001;
														assign node18905 = (inp[9]) ? 4'b1001 : 4'b1101;
													assign node18908 = (inp[10]) ? node18912 : node18909;
														assign node18909 = (inp[12]) ? 4'b1101 : 4'b1001;
														assign node18912 = (inp[4]) ? 4'b1001 : 4'b1001;
												assign node18915 = (inp[9]) ? node18923 : node18916;
													assign node18916 = (inp[12]) ? node18920 : node18917;
														assign node18917 = (inp[4]) ? 4'b1001 : 4'b1001;
														assign node18920 = (inp[4]) ? 4'b1111 : 4'b1001;
													assign node18923 = (inp[14]) ? 4'b1111 : 4'b1011;
											assign node18926 = (inp[5]) ? node18936 : node18927;
												assign node18927 = (inp[12]) ? node18929 : 4'b1001;
													assign node18929 = (inp[10]) ? node18933 : node18930;
														assign node18930 = (inp[14]) ? 4'b1111 : 4'b1011;
														assign node18933 = (inp[9]) ? 4'b1011 : 4'b1001;
												assign node18936 = (inp[4]) ? node18938 : 4'b1011;
													assign node18938 = (inp[12]) ? node18942 : node18939;
														assign node18939 = (inp[9]) ? 4'b1111 : 4'b1111;
														assign node18942 = (inp[9]) ? 4'b1011 : 4'b1111;
										assign node18945 = (inp[3]) ? node18967 : node18946;
											assign node18946 = (inp[5]) ? node18956 : node18947;
												assign node18947 = (inp[14]) ? node18951 : node18948;
													assign node18948 = (inp[9]) ? 4'b1111 : 4'b1011;
													assign node18951 = (inp[4]) ? 4'b1111 : node18952;
														assign node18952 = (inp[12]) ? 4'b1011 : 4'b1011;
												assign node18956 = (inp[9]) ? node18962 : node18957;
													assign node18957 = (inp[12]) ? node18959 : 4'b1011;
														assign node18959 = (inp[4]) ? 4'b1101 : 4'b1011;
													assign node18962 = (inp[12]) ? 4'b1001 : node18963;
														assign node18963 = (inp[4]) ? 4'b1101 : 4'b1001;
											assign node18967 = (inp[5]) ? node18979 : node18968;
												assign node18968 = (inp[4]) ? node18974 : node18969;
													assign node18969 = (inp[9]) ? 4'b1101 : node18970;
														assign node18970 = (inp[10]) ? 4'b1011 : 4'b1011;
													assign node18974 = (inp[9]) ? node18976 : 4'b1101;
														assign node18976 = (inp[12]) ? 4'b1001 : 4'b1101;
												assign node18979 = (inp[9]) ? node18987 : node18980;
													assign node18980 = (inp[10]) ? node18984 : node18981;
														assign node18981 = (inp[4]) ? 4'b1001 : 4'b1101;
														assign node18984 = (inp[4]) ? 4'b1101 : 4'b1001;
													assign node18987 = (inp[14]) ? 4'b1101 : node18988;
														assign node18988 = (inp[4]) ? 4'b1001 : 4'b1101;
								assign node18992 = (inp[2]) ? node19090 : node18993;
									assign node18993 = (inp[14]) ? node19047 : node18994;
										assign node18994 = (inp[3]) ? node19022 : node18995;
											assign node18995 = (inp[15]) ? node19011 : node18996;
												assign node18996 = (inp[9]) ? node19004 : node18997;
													assign node18997 = (inp[10]) ? node19001 : node18998;
														assign node18998 = (inp[4]) ? 4'b1001 : 4'b1101;
														assign node19001 = (inp[4]) ? 4'b1101 : 4'b1001;
													assign node19004 = (inp[5]) ? node19008 : node19005;
														assign node19005 = (inp[12]) ? 4'b1001 : 4'b1101;
														assign node19008 = (inp[4]) ? 4'b1011 : 4'b1111;
												assign node19011 = (inp[5]) ? node19017 : node19012;
													assign node19012 = (inp[4]) ? node19014 : 4'b1111;
														assign node19014 = (inp[9]) ? 4'b1011 : 4'b1111;
													assign node19017 = (inp[12]) ? 4'b1101 : node19018;
														assign node19018 = (inp[9]) ? 4'b1101 : 4'b1111;
											assign node19022 = (inp[15]) ? node19034 : node19023;
												assign node19023 = (inp[5]) ? node19029 : node19024;
													assign node19024 = (inp[4]) ? node19026 : 4'b1111;
														assign node19026 = (inp[10]) ? 4'b1011 : 4'b1001;
													assign node19029 = (inp[12]) ? 4'b1011 : node19030;
														assign node19030 = (inp[10]) ? 4'b1011 : 4'b1011;
												assign node19034 = (inp[5]) ? node19042 : node19035;
													assign node19035 = (inp[4]) ? node19039 : node19036;
														assign node19036 = (inp[12]) ? 4'b1011 : 4'b1111;
														assign node19039 = (inp[12]) ? 4'b1001 : 4'b1101;
													assign node19042 = (inp[9]) ? node19044 : 4'b1001;
														assign node19044 = (inp[4]) ? 4'b1001 : 4'b1101;
										assign node19047 = (inp[9]) ? node19067 : node19048;
											assign node19048 = (inp[4]) ? node19060 : node19049;
												assign node19049 = (inp[15]) ? node19055 : node19050;
													assign node19050 = (inp[5]) ? node19052 : 4'b1000;
														assign node19052 = (inp[10]) ? 4'b1000 : 4'b1100;
													assign node19055 = (inp[3]) ? 4'b1000 : node19056;
														assign node19056 = (inp[10]) ? 4'b1010 : 4'b1010;
												assign node19060 = (inp[15]) ? node19064 : node19061;
													assign node19061 = (inp[12]) ? 4'b1110 : 4'b1010;
													assign node19064 = (inp[10]) ? 4'b1100 : 4'b1000;
											assign node19067 = (inp[4]) ? node19077 : node19068;
												assign node19068 = (inp[3]) ? node19074 : node19069;
													assign node19069 = (inp[10]) ? node19071 : 4'b1110;
														assign node19071 = (inp[12]) ? 4'b1100 : 4'b1110;
													assign node19074 = (inp[15]) ? 4'b1100 : 4'b1110;
												assign node19077 = (inp[12]) ? node19083 : node19078;
													assign node19078 = (inp[15]) ? 4'b1100 : node19079;
														assign node19079 = (inp[3]) ? 4'b1110 : 4'b1010;
													assign node19083 = (inp[5]) ? node19087 : node19084;
														assign node19084 = (inp[15]) ? 4'b1010 : 4'b1000;
														assign node19087 = (inp[15]) ? 4'b1000 : 4'b1010;
									assign node19090 = (inp[15]) ? node19132 : node19091;
										assign node19091 = (inp[3]) ? node19115 : node19092;
											assign node19092 = (inp[5]) ? node19104 : node19093;
												assign node19093 = (inp[4]) ? node19099 : node19094;
													assign node19094 = (inp[14]) ? node19096 : 4'b1000;
														assign node19096 = (inp[12]) ? 4'b1000 : 4'b1100;
													assign node19099 = (inp[9]) ? node19101 : 4'b1100;
														assign node19101 = (inp[14]) ? 4'b1000 : 4'b1100;
												assign node19104 = (inp[9]) ? node19112 : node19105;
													assign node19105 = (inp[4]) ? node19109 : node19106;
														assign node19106 = (inp[14]) ? 4'b1100 : 4'b1000;
														assign node19109 = (inp[12]) ? 4'b1110 : 4'b1000;
													assign node19112 = (inp[4]) ? 4'b1010 : 4'b1110;
											assign node19115 = (inp[5]) ? node19123 : node19116;
												assign node19116 = (inp[9]) ? 4'b1110 : node19117;
													assign node19117 = (inp[4]) ? 4'b1110 : node19118;
														assign node19118 = (inp[10]) ? 4'b1000 : 4'b1100;
												assign node19123 = (inp[9]) ? node19129 : node19124;
													assign node19124 = (inp[4]) ? 4'b1110 : node19125;
														assign node19125 = (inp[12]) ? 4'b1010 : 4'b1110;
													assign node19129 = (inp[4]) ? 4'b1010 : 4'b1110;
										assign node19132 = (inp[3]) ? node19152 : node19133;
											assign node19133 = (inp[5]) ? node19141 : node19134;
												assign node19134 = (inp[14]) ? node19136 : 4'b1110;
													assign node19136 = (inp[9]) ? 4'b1010 : node19137;
														assign node19137 = (inp[4]) ? 4'b1110 : 4'b1010;
												assign node19141 = (inp[4]) ? node19147 : node19142;
													assign node19142 = (inp[9]) ? node19144 : 4'b1010;
														assign node19144 = (inp[10]) ? 4'b1100 : 4'b1010;
													assign node19147 = (inp[10]) ? 4'b1100 : node19148;
														assign node19148 = (inp[12]) ? 4'b1000 : 4'b1010;
											assign node19152 = (inp[5]) ? node19162 : node19153;
												assign node19153 = (inp[9]) ? node19159 : node19154;
													assign node19154 = (inp[14]) ? 4'b1010 : node19155;
														assign node19155 = (inp[12]) ? 4'b1100 : 4'b1110;
													assign node19159 = (inp[4]) ? 4'b1000 : 4'b1100;
												assign node19162 = (inp[9]) ? node19168 : node19163;
													assign node19163 = (inp[12]) ? 4'b1000 : node19164;
														assign node19164 = (inp[14]) ? 4'b1000 : 4'b1100;
													assign node19168 = (inp[4]) ? 4'b1000 : node19169;
														assign node19169 = (inp[12]) ? 4'b1100 : 4'b1000;
						assign node19173 = (inp[15]) ? node19537 : node19174;
							assign node19174 = (inp[3]) ? node19360 : node19175;
								assign node19175 = (inp[5]) ? node19271 : node19176;
									assign node19176 = (inp[7]) ? node19224 : node19177;
										assign node19177 = (inp[8]) ? node19199 : node19178;
											assign node19178 = (inp[14]) ? node19190 : node19179;
												assign node19179 = (inp[2]) ? node19187 : node19180;
													assign node19180 = (inp[4]) ? node19184 : node19181;
														assign node19181 = (inp[10]) ? 4'b1101 : 4'b1001;
														assign node19184 = (inp[9]) ? 4'b1001 : 4'b1101;
													assign node19187 = (inp[9]) ? 4'b1000 : 4'b1100;
												assign node19190 = (inp[2]) ? node19194 : node19191;
													assign node19191 = (inp[9]) ? 4'b1100 : 4'b1000;
													assign node19194 = (inp[4]) ? node19196 : 4'b1100;
														assign node19196 = (inp[9]) ? 4'b1000 : 4'b1100;
											assign node19199 = (inp[4]) ? node19213 : node19200;
												assign node19200 = (inp[14]) ? node19208 : node19201;
													assign node19201 = (inp[2]) ? node19205 : node19202;
														assign node19202 = (inp[10]) ? 4'b1000 : 4'b1000;
														assign node19205 = (inp[9]) ? 4'b1101 : 4'b1001;
													assign node19208 = (inp[12]) ? 4'b1001 : node19209;
														assign node19209 = (inp[2]) ? 4'b1001 : 4'b1001;
												assign node19213 = (inp[10]) ? node19219 : node19214;
													assign node19214 = (inp[2]) ? node19216 : 4'b1101;
														assign node19216 = (inp[14]) ? 4'b1001 : 4'b1001;
													assign node19219 = (inp[2]) ? 4'b1101 : node19220;
														assign node19220 = (inp[14]) ? 4'b1101 : 4'b1100;
										assign node19224 = (inp[8]) ? node19246 : node19225;
											assign node19225 = (inp[14]) ? node19239 : node19226;
												assign node19226 = (inp[2]) ? node19234 : node19227;
													assign node19227 = (inp[12]) ? node19231 : node19228;
														assign node19228 = (inp[9]) ? 4'b1000 : 4'b1000;
														assign node19231 = (inp[9]) ? 4'b1100 : 4'b1000;
													assign node19234 = (inp[9]) ? node19236 : 4'b1001;
														assign node19236 = (inp[4]) ? 4'b1001 : 4'b1101;
												assign node19239 = (inp[4]) ? node19241 : 4'b1101;
													assign node19241 = (inp[9]) ? 4'b1001 : node19242;
														assign node19242 = (inp[12]) ? 4'b1101 : 4'b1001;
											assign node19246 = (inp[2]) ? node19258 : node19247;
												assign node19247 = (inp[14]) ? node19253 : node19248;
													assign node19248 = (inp[12]) ? node19250 : 4'b1101;
														assign node19250 = (inp[10]) ? 4'b1101 : 4'b1001;
													assign node19253 = (inp[10]) ? node19255 : 4'b1000;
														assign node19255 = (inp[12]) ? 4'b1000 : 4'b1100;
												assign node19258 = (inp[12]) ? node19266 : node19259;
													assign node19259 = (inp[10]) ? node19263 : node19260;
														assign node19260 = (inp[4]) ? 4'b1000 : 4'b1000;
														assign node19263 = (inp[9]) ? 4'b1000 : 4'b1100;
													assign node19266 = (inp[10]) ? node19268 : 4'b1100;
														assign node19268 = (inp[14]) ? 4'b1100 : 4'b1000;
									assign node19271 = (inp[4]) ? node19317 : node19272;
										assign node19272 = (inp[9]) ? node19298 : node19273;
											assign node19273 = (inp[12]) ? node19285 : node19274;
												assign node19274 = (inp[10]) ? node19280 : node19275;
													assign node19275 = (inp[8]) ? node19277 : 4'b1101;
														assign node19277 = (inp[14]) ? 4'b1101 : 4'b1100;
													assign node19280 = (inp[7]) ? node19282 : 4'b1000;
														assign node19282 = (inp[8]) ? 4'b1000 : 4'b1001;
												assign node19285 = (inp[8]) ? node19291 : node19286;
													assign node19286 = (inp[2]) ? 4'b1001 : node19287;
														assign node19287 = (inp[14]) ? 4'b1001 : 4'b1000;
													assign node19291 = (inp[14]) ? node19295 : node19292;
														assign node19292 = (inp[7]) ? 4'b1001 : 4'b1000;
														assign node19295 = (inp[7]) ? 4'b1000 : 4'b1001;
											assign node19298 = (inp[10]) ? node19306 : node19299;
												assign node19299 = (inp[12]) ? 4'b1110 : node19300;
													assign node19300 = (inp[2]) ? node19302 : 4'b1000;
														assign node19302 = (inp[8]) ? 4'b1001 : 4'b1000;
												assign node19306 = (inp[14]) ? node19312 : node19307;
													assign node19307 = (inp[8]) ? 4'b1111 : node19308;
														assign node19308 = (inp[12]) ? 4'b1110 : 4'b1110;
													assign node19312 = (inp[7]) ? 4'b1110 : node19313;
														assign node19313 = (inp[8]) ? 4'b1111 : 4'b1110;
										assign node19317 = (inp[9]) ? node19341 : node19318;
											assign node19318 = (inp[10]) ? node19328 : node19319;
												assign node19319 = (inp[12]) ? node19323 : node19320;
													assign node19320 = (inp[8]) ? 4'b1000 : 4'b1001;
													assign node19323 = (inp[2]) ? node19325 : 4'b1110;
														assign node19325 = (inp[7]) ? 4'b1111 : 4'b1110;
												assign node19328 = (inp[14]) ? node19334 : node19329;
													assign node19329 = (inp[7]) ? 4'b1110 : node19330;
														assign node19330 = (inp[2]) ? 4'b1110 : 4'b1110;
													assign node19334 = (inp[2]) ? node19338 : node19335;
														assign node19335 = (inp[12]) ? 4'b1111 : 4'b1110;
														assign node19338 = (inp[8]) ? 4'b1110 : 4'b1111;
											assign node19341 = (inp[10]) ? node19351 : node19342;
												assign node19342 = (inp[8]) ? node19348 : node19343;
													assign node19343 = (inp[2]) ? 4'b1110 : node19344;
														assign node19344 = (inp[7]) ? 4'b1110 : 4'b1111;
													assign node19348 = (inp[7]) ? 4'b1011 : 4'b1010;
												assign node19351 = (inp[12]) ? node19357 : node19352;
													assign node19352 = (inp[8]) ? node19354 : 4'b1010;
														assign node19354 = (inp[7]) ? 4'b1010 : 4'b1011;
													assign node19357 = (inp[7]) ? 4'b1011 : 4'b1010;
								assign node19360 = (inp[5]) ? node19450 : node19361;
									assign node19361 = (inp[4]) ? node19405 : node19362;
										assign node19362 = (inp[9]) ? node19384 : node19363;
											assign node19363 = (inp[12]) ? node19371 : node19364;
												assign node19364 = (inp[10]) ? node19366 : 4'b1101;
													assign node19366 = (inp[8]) ? node19368 : 4'b1000;
														assign node19368 = (inp[7]) ? 4'b1000 : 4'b1001;
												assign node19371 = (inp[7]) ? node19377 : node19372;
													assign node19372 = (inp[8]) ? node19374 : 4'b1000;
														assign node19374 = (inp[2]) ? 4'b1001 : 4'b1000;
													assign node19377 = (inp[8]) ? node19381 : node19378;
														assign node19378 = (inp[2]) ? 4'b1001 : 4'b1000;
														assign node19381 = (inp[10]) ? 4'b1001 : 4'b1000;
											assign node19384 = (inp[10]) ? node19396 : node19385;
												assign node19385 = (inp[12]) ? node19391 : node19386;
													assign node19386 = (inp[14]) ? 4'b1001 : node19387;
														assign node19387 = (inp[7]) ? 4'b1000 : 4'b1001;
													assign node19391 = (inp[14]) ? 4'b1110 : node19392;
														assign node19392 = (inp[7]) ? 4'b1110 : 4'b1110;
												assign node19396 = (inp[8]) ? node19402 : node19397;
													assign node19397 = (inp[7]) ? 4'b1111 : node19398;
														assign node19398 = (inp[12]) ? 4'b1111 : 4'b1110;
													assign node19402 = (inp[7]) ? 4'b1110 : 4'b1111;
										assign node19405 = (inp[9]) ? node19425 : node19406;
											assign node19406 = (inp[10]) ? node19412 : node19407;
												assign node19407 = (inp[8]) ? node19409 : 4'b1111;
													assign node19409 = (inp[14]) ? 4'b1000 : 4'b1001;
												assign node19412 = (inp[14]) ? node19420 : node19413;
													assign node19413 = (inp[2]) ? node19417 : node19414;
														assign node19414 = (inp[7]) ? 4'b1110 : 4'b1111;
														assign node19417 = (inp[8]) ? 4'b1110 : 4'b1110;
													assign node19420 = (inp[12]) ? 4'b1111 : node19421;
														assign node19421 = (inp[2]) ? 4'b1111 : 4'b1110;
											assign node19425 = (inp[12]) ? node19437 : node19426;
												assign node19426 = (inp[10]) ? node19432 : node19427;
													assign node19427 = (inp[7]) ? node19429 : 4'b1111;
														assign node19429 = (inp[14]) ? 4'b1110 : 4'b1111;
													assign node19432 = (inp[7]) ? 4'b1010 : node19433;
														assign node19433 = (inp[8]) ? 4'b1011 : 4'b1010;
												assign node19437 = (inp[8]) ? node19443 : node19438;
													assign node19438 = (inp[7]) ? node19440 : 4'b1010;
														assign node19440 = (inp[2]) ? 4'b1011 : 4'b1010;
													assign node19443 = (inp[7]) ? node19447 : node19444;
														assign node19444 = (inp[2]) ? 4'b1011 : 4'b1010;
														assign node19447 = (inp[2]) ? 4'b1010 : 4'b1011;
									assign node19450 = (inp[4]) ? node19498 : node19451;
										assign node19451 = (inp[9]) ? node19481 : node19452;
											assign node19452 = (inp[10]) ? node19468 : node19453;
												assign node19453 = (inp[12]) ? node19461 : node19454;
													assign node19454 = (inp[8]) ? node19458 : node19455;
														assign node19455 = (inp[2]) ? 4'b1110 : 4'b1111;
														assign node19458 = (inp[7]) ? 4'b1110 : 4'b1111;
													assign node19461 = (inp[14]) ? node19465 : node19462;
														assign node19462 = (inp[2]) ? 4'b1010 : 4'b1011;
														assign node19465 = (inp[2]) ? 4'b1011 : 4'b1010;
												assign node19468 = (inp[7]) ? node19474 : node19469;
													assign node19469 = (inp[12]) ? 4'b1011 : node19470;
														assign node19470 = (inp[8]) ? 4'b1011 : 4'b1010;
													assign node19474 = (inp[8]) ? node19478 : node19475;
														assign node19475 = (inp[2]) ? 4'b1011 : 4'b1010;
														assign node19478 = (inp[14]) ? 4'b1010 : 4'b1010;
											assign node19481 = (inp[12]) ? node19487 : node19482;
												assign node19482 = (inp[10]) ? 4'b1111 : node19483;
													assign node19483 = (inp[7]) ? 4'b1011 : 4'b1010;
												assign node19487 = (inp[7]) ? node19493 : node19488;
													assign node19488 = (inp[8]) ? node19490 : 4'b1110;
														assign node19490 = (inp[2]) ? 4'b1111 : 4'b1110;
													assign node19493 = (inp[2]) ? 4'b1111 : node19494;
														assign node19494 = (inp[8]) ? 4'b1111 : 4'b1110;
										assign node19498 = (inp[9]) ? node19520 : node19499;
											assign node19499 = (inp[10]) ? node19511 : node19500;
												assign node19500 = (inp[12]) ? node19506 : node19501;
													assign node19501 = (inp[14]) ? 4'b1011 : node19502;
														assign node19502 = (inp[7]) ? 4'b1010 : 4'b1011;
													assign node19506 = (inp[8]) ? 4'b1111 : node19507;
														assign node19507 = (inp[2]) ? 4'b1110 : 4'b1110;
												assign node19511 = (inp[2]) ? node19513 : 4'b1111;
													assign node19513 = (inp[8]) ? node19517 : node19514;
														assign node19514 = (inp[7]) ? 4'b1111 : 4'b1110;
														assign node19517 = (inp[7]) ? 4'b1110 : 4'b1111;
											assign node19520 = (inp[12]) ? node19530 : node19521;
												assign node19521 = (inp[10]) ? node19527 : node19522;
													assign node19522 = (inp[14]) ? node19524 : 4'b1111;
														assign node19524 = (inp[2]) ? 4'b1110 : 4'b1110;
													assign node19527 = (inp[2]) ? 4'b1010 : 4'b1011;
												assign node19530 = (inp[10]) ? node19532 : 4'b1010;
													assign node19532 = (inp[7]) ? 4'b1011 : node19533;
														assign node19533 = (inp[14]) ? 4'b1011 : 4'b1010;
							assign node19537 = (inp[5]) ? node19713 : node19538;
								assign node19538 = (inp[3]) ? node19624 : node19539;
									assign node19539 = (inp[8]) ? node19581 : node19540;
										assign node19540 = (inp[7]) ? node19558 : node19541;
											assign node19541 = (inp[14]) ? node19549 : node19542;
												assign node19542 = (inp[4]) ? node19546 : node19543;
													assign node19543 = (inp[10]) ? 4'b1111 : 4'b1011;
													assign node19546 = (inp[9]) ? 4'b1010 : 4'b1110;
												assign node19549 = (inp[4]) ? node19551 : 4'b1110;
													assign node19551 = (inp[9]) ? node19555 : node19552;
														assign node19552 = (inp[12]) ? 4'b1110 : 4'b1110;
														assign node19555 = (inp[10]) ? 4'b1010 : 4'b1110;
											assign node19558 = (inp[2]) ? node19570 : node19559;
												assign node19559 = (inp[14]) ? node19565 : node19560;
													assign node19560 = (inp[9]) ? 4'b1110 : node19561;
														assign node19561 = (inp[4]) ? 4'b1010 : 4'b1010;
													assign node19565 = (inp[9]) ? 4'b1111 : node19566;
														assign node19566 = (inp[10]) ? 4'b1111 : 4'b1011;
												assign node19570 = (inp[4]) ? node19576 : node19571;
													assign node19571 = (inp[10]) ? 4'b1011 : node19572;
														assign node19572 = (inp[12]) ? 4'b1011 : 4'b1011;
													assign node19576 = (inp[9]) ? node19578 : 4'b1111;
														assign node19578 = (inp[10]) ? 4'b1011 : 4'b1111;
										assign node19581 = (inp[7]) ? node19601 : node19582;
											assign node19582 = (inp[4]) ? node19590 : node19583;
												assign node19583 = (inp[9]) ? 4'b1111 : node19584;
													assign node19584 = (inp[10]) ? 4'b1011 : node19585;
														assign node19585 = (inp[12]) ? 4'b1011 : 4'b1111;
												assign node19590 = (inp[9]) ? node19596 : node19591;
													assign node19591 = (inp[10]) ? 4'b1111 : node19592;
														assign node19592 = (inp[14]) ? 4'b1011 : 4'b1010;
													assign node19596 = (inp[2]) ? 4'b1011 : node19597;
														assign node19597 = (inp[14]) ? 4'b1011 : 4'b1010;
											assign node19601 = (inp[14]) ? node19613 : node19602;
												assign node19602 = (inp[2]) ? node19608 : node19603;
													assign node19603 = (inp[10]) ? node19605 : 4'b1111;
														assign node19605 = (inp[4]) ? 4'b1011 : 4'b1011;
													assign node19608 = (inp[9]) ? node19610 : 4'b1010;
														assign node19610 = (inp[4]) ? 4'b1010 : 4'b1010;
												assign node19613 = (inp[12]) ? node19619 : node19614;
													assign node19614 = (inp[10]) ? 4'b1110 : node19615;
														assign node19615 = (inp[4]) ? 4'b1010 : 4'b1010;
													assign node19619 = (inp[10]) ? node19621 : 4'b1110;
														assign node19621 = (inp[4]) ? 4'b1110 : 4'b1010;
									assign node19624 = (inp[9]) ? node19672 : node19625;
										assign node19625 = (inp[4]) ? node19645 : node19626;
											assign node19626 = (inp[12]) ? node19634 : node19627;
												assign node19627 = (inp[8]) ? node19631 : node19628;
													assign node19628 = (inp[10]) ? 4'b1010 : 4'b1110;
													assign node19631 = (inp[14]) ? 4'b1111 : 4'b1011;
												assign node19634 = (inp[7]) ? node19640 : node19635;
													assign node19635 = (inp[8]) ? node19637 : 4'b1010;
														assign node19637 = (inp[14]) ? 4'b1011 : 4'b1010;
													assign node19640 = (inp[14]) ? node19642 : 4'b1011;
														assign node19642 = (inp[8]) ? 4'b1010 : 4'b1011;
											assign node19645 = (inp[12]) ? node19659 : node19646;
												assign node19646 = (inp[10]) ? node19654 : node19647;
													assign node19647 = (inp[2]) ? node19651 : node19648;
														assign node19648 = (inp[14]) ? 4'b1010 : 4'b1011;
														assign node19651 = (inp[8]) ? 4'b1011 : 4'b1011;
													assign node19654 = (inp[14]) ? 4'b1100 : node19655;
														assign node19655 = (inp[7]) ? 4'b1100 : 4'b1101;
												assign node19659 = (inp[14]) ? node19667 : node19660;
													assign node19660 = (inp[7]) ? node19664 : node19661;
														assign node19661 = (inp[2]) ? 4'b1100 : 4'b1100;
														assign node19664 = (inp[8]) ? 4'b1100 : 4'b1101;
													assign node19667 = (inp[2]) ? node19669 : 4'b1100;
														assign node19669 = (inp[8]) ? 4'b1101 : 4'b1100;
										assign node19672 = (inp[4]) ? node19692 : node19673;
											assign node19673 = (inp[10]) ? node19683 : node19674;
												assign node19674 = (inp[12]) ? node19680 : node19675;
													assign node19675 = (inp[7]) ? 4'b1011 : node19676;
														assign node19676 = (inp[8]) ? 4'b1011 : 4'b1010;
													assign node19680 = (inp[2]) ? 4'b1101 : 4'b1100;
												assign node19683 = (inp[8]) ? node19687 : node19684;
													assign node19684 = (inp[7]) ? 4'b1101 : 4'b1100;
													assign node19687 = (inp[12]) ? node19689 : 4'b1101;
														assign node19689 = (inp[7]) ? 4'b1101 : 4'b1101;
											assign node19692 = (inp[12]) ? node19702 : node19693;
												assign node19693 = (inp[10]) ? node19699 : node19694;
													assign node19694 = (inp[7]) ? 4'b1100 : node19695;
														assign node19695 = (inp[8]) ? 4'b1101 : 4'b1100;
													assign node19699 = (inp[14]) ? 4'b1001 : 4'b1000;
												assign node19702 = (inp[10]) ? node19708 : node19703;
													assign node19703 = (inp[8]) ? node19705 : 4'b1000;
														assign node19705 = (inp[7]) ? 4'b1000 : 4'b1001;
													assign node19708 = (inp[14]) ? node19710 : 4'b1001;
														assign node19710 = (inp[8]) ? 4'b1000 : 4'b1000;
								assign node19713 = (inp[3]) ? node19801 : node19714;
									assign node19714 = (inp[4]) ? node19756 : node19715;
										assign node19715 = (inp[9]) ? node19735 : node19716;
											assign node19716 = (inp[12]) ? node19726 : node19717;
												assign node19717 = (inp[10]) ? node19723 : node19718;
													assign node19718 = (inp[7]) ? 4'b1111 : node19719;
														assign node19719 = (inp[14]) ? 4'b1110 : 4'b1111;
													assign node19723 = (inp[8]) ? 4'b1010 : 4'b1011;
												assign node19726 = (inp[10]) ? node19728 : 4'b1010;
													assign node19728 = (inp[2]) ? node19732 : node19729;
														assign node19729 = (inp[7]) ? 4'b1010 : 4'b1011;
														assign node19732 = (inp[8]) ? 4'b1010 : 4'b1010;
											assign node19735 = (inp[12]) ? node19747 : node19736;
												assign node19736 = (inp[10]) ? node19742 : node19737;
													assign node19737 = (inp[14]) ? node19739 : 4'b1011;
														assign node19739 = (inp[7]) ? 4'b1011 : 4'b1010;
													assign node19742 = (inp[14]) ? node19744 : 4'b1100;
														assign node19744 = (inp[7]) ? 4'b1101 : 4'b1100;
												assign node19747 = (inp[8]) ? node19749 : 4'b1100;
													assign node19749 = (inp[10]) ? node19753 : node19750;
														assign node19750 = (inp[2]) ? 4'b1100 : 4'b1100;
														assign node19753 = (inp[7]) ? 4'b1100 : 4'b1101;
										assign node19756 = (inp[9]) ? node19780 : node19757;
											assign node19757 = (inp[12]) ? node19769 : node19758;
												assign node19758 = (inp[10]) ? node19764 : node19759;
													assign node19759 = (inp[14]) ? 4'b1011 : node19760;
														assign node19760 = (inp[8]) ? 4'b1010 : 4'b1010;
													assign node19764 = (inp[14]) ? 4'b1100 : node19765;
														assign node19765 = (inp[7]) ? 4'b1101 : 4'b1100;
												assign node19769 = (inp[10]) ? node19775 : node19770;
													assign node19770 = (inp[14]) ? node19772 : 4'b1101;
														assign node19772 = (inp[7]) ? 4'b1100 : 4'b1100;
													assign node19775 = (inp[2]) ? 4'b1101 : node19776;
														assign node19776 = (inp[7]) ? 4'b1101 : 4'b1100;
											assign node19780 = (inp[10]) ? node19790 : node19781;
												assign node19781 = (inp[12]) ? node19785 : node19782;
													assign node19782 = (inp[2]) ? 4'b1101 : 4'b1100;
													assign node19785 = (inp[7]) ? 4'b1001 : node19786;
														assign node19786 = (inp[8]) ? 4'b1001 : 4'b1000;
												assign node19790 = (inp[8]) ? node19796 : node19791;
													assign node19791 = (inp[7]) ? node19793 : 4'b1000;
														assign node19793 = (inp[14]) ? 4'b1001 : 4'b1000;
													assign node19796 = (inp[7]) ? node19798 : 4'b1001;
														assign node19798 = (inp[14]) ? 4'b1000 : 4'b1001;
									assign node19801 = (inp[9]) ? node19841 : node19802;
										assign node19802 = (inp[4]) ? node19824 : node19803;
											assign node19803 = (inp[10]) ? node19815 : node19804;
												assign node19804 = (inp[12]) ? node19810 : node19805;
													assign node19805 = (inp[2]) ? node19807 : 4'b1100;
														assign node19807 = (inp[8]) ? 4'b1100 : 4'b1101;
													assign node19810 = (inp[2]) ? node19812 : 4'b1001;
														assign node19812 = (inp[7]) ? 4'b1000 : 4'b1000;
												assign node19815 = (inp[12]) ? 4'b1001 : node19816;
													assign node19816 = (inp[7]) ? node19820 : node19817;
														assign node19817 = (inp[8]) ? 4'b1001 : 4'b1000;
														assign node19820 = (inp[8]) ? 4'b1000 : 4'b1000;
											assign node19824 = (inp[10]) ? node19836 : node19825;
												assign node19825 = (inp[12]) ? node19833 : node19826;
													assign node19826 = (inp[2]) ? node19830 : node19827;
														assign node19827 = (inp[8]) ? 4'b1001 : 4'b1000;
														assign node19830 = (inp[7]) ? 4'b1000 : 4'b1000;
													assign node19833 = (inp[7]) ? 4'b1100 : 4'b1101;
												assign node19836 = (inp[12]) ? node19838 : 4'b1101;
													assign node19838 = (inp[2]) ? 4'b1101 : 4'b1100;
										assign node19841 = (inp[4]) ? node19861 : node19842;
											assign node19842 = (inp[12]) ? node19854 : node19843;
												assign node19843 = (inp[10]) ? node19849 : node19844;
													assign node19844 = (inp[7]) ? node19846 : 4'b1001;
														assign node19846 = (inp[14]) ? 4'b1001 : 4'b1000;
													assign node19849 = (inp[8]) ? 4'b1101 : node19850;
														assign node19850 = (inp[7]) ? 4'b1101 : 4'b1100;
												assign node19854 = (inp[7]) ? 4'b1100 : node19855;
													assign node19855 = (inp[10]) ? node19857 : 4'b1101;
														assign node19857 = (inp[8]) ? 4'b1100 : 4'b1100;
											assign node19861 = (inp[12]) ? node19867 : node19862;
												assign node19862 = (inp[10]) ? 4'b1001 : node19863;
													assign node19863 = (inp[7]) ? 4'b1101 : 4'b1100;
												assign node19867 = (inp[14]) ? node19869 : 4'b1001;
													assign node19869 = (inp[7]) ? 4'b1000 : node19870;
														assign node19870 = (inp[8]) ? 4'b1001 : 4'b1000;
				assign node19874 = (inp[1]) ? node21320 : node19875;
					assign node19875 = (inp[13]) ? node20597 : node19876;
						assign node19876 = (inp[15]) ? node20230 : node19877;
							assign node19877 = (inp[3]) ? node20055 : node19878;
								assign node19878 = (inp[5]) ? node19970 : node19879;
									assign node19879 = (inp[12]) ? node19925 : node19880;
										assign node19880 = (inp[2]) ? node19902 : node19881;
											assign node19881 = (inp[9]) ? node19891 : node19882;
												assign node19882 = (inp[7]) ? 4'b1100 : node19883;
													assign node19883 = (inp[10]) ? node19887 : node19884;
														assign node19884 = (inp[8]) ? 4'b1100 : 4'b1100;
														assign node19887 = (inp[14]) ? 4'b1101 : 4'b1100;
												assign node19891 = (inp[8]) ? node19899 : node19892;
													assign node19892 = (inp[7]) ? node19896 : node19893;
														assign node19893 = (inp[14]) ? 4'b1000 : 4'b1001;
														assign node19896 = (inp[14]) ? 4'b1101 : 4'b1100;
													assign node19899 = (inp[4]) ? 4'b1101 : 4'b1001;
											assign node19902 = (inp[14]) ? node19912 : node19903;
												assign node19903 = (inp[9]) ? node19905 : 4'b1001;
													assign node19905 = (inp[8]) ? node19909 : node19906;
														assign node19906 = (inp[7]) ? 4'b1001 : 4'b1000;
														assign node19909 = (inp[7]) ? 4'b1100 : 4'b1101;
												assign node19912 = (inp[4]) ? node19920 : node19913;
													assign node19913 = (inp[8]) ? node19917 : node19914;
														assign node19914 = (inp[7]) ? 4'b1001 : 4'b1000;
														assign node19917 = (inp[9]) ? 4'b1000 : 4'b1000;
													assign node19920 = (inp[8]) ? 4'b1001 : node19921;
														assign node19921 = (inp[7]) ? 4'b1001 : 4'b1100;
										assign node19925 = (inp[7]) ? node19951 : node19926;
											assign node19926 = (inp[8]) ? node19940 : node19927;
												assign node19927 = (inp[14]) ? node19933 : node19928;
													assign node19928 = (inp[4]) ? node19930 : 4'b1101;
														assign node19930 = (inp[2]) ? 4'b1000 : 4'b1001;
													assign node19933 = (inp[9]) ? node19937 : node19934;
														assign node19934 = (inp[4]) ? 4'b1100 : 4'b1000;
														assign node19937 = (inp[4]) ? 4'b1000 : 4'b1100;
												assign node19940 = (inp[2]) ? node19946 : node19941;
													assign node19941 = (inp[14]) ? 4'b1101 : node19942;
														assign node19942 = (inp[4]) ? 4'b1000 : 4'b1000;
													assign node19946 = (inp[4]) ? 4'b1001 : node19947;
														assign node19947 = (inp[9]) ? 4'b1101 : 4'b1001;
											assign node19951 = (inp[8]) ? node19961 : node19952;
												assign node19952 = (inp[14]) ? node19956 : node19953;
													assign node19953 = (inp[4]) ? 4'b1100 : 4'b1000;
													assign node19956 = (inp[4]) ? 4'b1001 : node19957;
														assign node19957 = (inp[9]) ? 4'b1101 : 4'b1001;
												assign node19961 = (inp[14]) ? node19965 : node19962;
													assign node19962 = (inp[2]) ? 4'b1000 : 4'b1001;
													assign node19965 = (inp[4]) ? 4'b1000 : node19966;
														assign node19966 = (inp[9]) ? 4'b1100 : 4'b1000;
									assign node19970 = (inp[4]) ? node20014 : node19971;
										assign node19971 = (inp[9]) ? node19995 : node19972;
											assign node19972 = (inp[10]) ? node19982 : node19973;
												assign node19973 = (inp[12]) ? node19979 : node19974;
													assign node19974 = (inp[8]) ? 4'b1100 : node19975;
														assign node19975 = (inp[7]) ? 4'b1101 : 4'b1100;
													assign node19979 = (inp[8]) ? 4'b1000 : 4'b1001;
												assign node19982 = (inp[14]) ? node19988 : node19983;
													assign node19983 = (inp[7]) ? 4'b1000 : node19984;
														assign node19984 = (inp[12]) ? 4'b1000 : 4'b1001;
													assign node19988 = (inp[7]) ? node19992 : node19989;
														assign node19989 = (inp[8]) ? 4'b1001 : 4'b1000;
														assign node19992 = (inp[12]) ? 4'b1001 : 4'b1000;
											assign node19995 = (inp[10]) ? node20005 : node19996;
												assign node19996 = (inp[12]) ? node20002 : node19997;
													assign node19997 = (inp[8]) ? 4'b1001 : node19998;
														assign node19998 = (inp[7]) ? 4'b1001 : 4'b1000;
													assign node20002 = (inp[14]) ? 4'b1111 : 4'b1110;
												assign node20005 = (inp[8]) ? node20007 : 4'b1110;
													assign node20007 = (inp[12]) ? node20011 : node20008;
														assign node20008 = (inp[7]) ? 4'b1110 : 4'b1111;
														assign node20011 = (inp[14]) ? 4'b1110 : 4'b1110;
										assign node20014 = (inp[9]) ? node20032 : node20015;
											assign node20015 = (inp[10]) ? node20023 : node20016;
												assign node20016 = (inp[12]) ? 4'b1110 : node20017;
													assign node20017 = (inp[2]) ? node20019 : 4'b1000;
														assign node20019 = (inp[7]) ? 4'b1000 : 4'b1000;
												assign node20023 = (inp[2]) ? node20027 : node20024;
													assign node20024 = (inp[8]) ? 4'b1110 : 4'b1111;
													assign node20027 = (inp[8]) ? 4'b1111 : node20028;
														assign node20028 = (inp[7]) ? 4'b1111 : 4'b1110;
											assign node20032 = (inp[12]) ? node20042 : node20033;
												assign node20033 = (inp[10]) ? node20039 : node20034;
													assign node20034 = (inp[2]) ? node20036 : 4'b1110;
														assign node20036 = (inp[14]) ? 4'b1110 : 4'b1111;
													assign node20039 = (inp[8]) ? 4'b1010 : 4'b1011;
												assign node20042 = (inp[10]) ? node20048 : node20043;
													assign node20043 = (inp[2]) ? node20045 : 4'b1011;
														assign node20045 = (inp[14]) ? 4'b1010 : 4'b1011;
													assign node20048 = (inp[7]) ? node20052 : node20049;
														assign node20049 = (inp[8]) ? 4'b1011 : 4'b1010;
														assign node20052 = (inp[8]) ? 4'b1010 : 4'b1011;
								assign node20055 = (inp[5]) ? node20141 : node20056;
									assign node20056 = (inp[9]) ? node20090 : node20057;
										assign node20057 = (inp[4]) ? node20079 : node20058;
											assign node20058 = (inp[10]) ? node20068 : node20059;
												assign node20059 = (inp[12]) ? node20065 : node20060;
													assign node20060 = (inp[2]) ? 4'b1101 : node20061;
														assign node20061 = (inp[7]) ? 4'b1101 : 4'b1100;
													assign node20065 = (inp[7]) ? 4'b1001 : 4'b1000;
												assign node20068 = (inp[7]) ? node20074 : node20069;
													assign node20069 = (inp[8]) ? 4'b1001 : node20070;
														assign node20070 = (inp[2]) ? 4'b1000 : 4'b1001;
													assign node20074 = (inp[8]) ? 4'b1000 : node20075;
														assign node20075 = (inp[2]) ? 4'b1001 : 4'b1000;
											assign node20079 = (inp[10]) ? node20085 : node20080;
												assign node20080 = (inp[12]) ? node20082 : 4'b1001;
													assign node20082 = (inp[14]) ? 4'b1110 : 4'b1111;
												assign node20085 = (inp[8]) ? node20087 : 4'b1111;
													assign node20087 = (inp[2]) ? 4'b1111 : 4'b1110;
										assign node20090 = (inp[4]) ? node20118 : node20091;
											assign node20091 = (inp[12]) ? node20105 : node20092;
												assign node20092 = (inp[10]) ? node20100 : node20093;
													assign node20093 = (inp[14]) ? node20097 : node20094;
														assign node20094 = (inp[8]) ? 4'b1000 : 4'b1000;
														assign node20097 = (inp[2]) ? 4'b1001 : 4'b1000;
													assign node20100 = (inp[14]) ? node20102 : 4'b1110;
														assign node20102 = (inp[8]) ? 4'b1111 : 4'b1110;
												assign node20105 = (inp[2]) ? node20111 : node20106;
													assign node20106 = (inp[8]) ? 4'b1111 : node20107;
														assign node20107 = (inp[14]) ? 4'b1111 : 4'b1110;
													assign node20111 = (inp[7]) ? node20115 : node20112;
														assign node20112 = (inp[8]) ? 4'b1111 : 4'b1110;
														assign node20115 = (inp[8]) ? 4'b1110 : 4'b1111;
											assign node20118 = (inp[12]) ? node20132 : node20119;
												assign node20119 = (inp[10]) ? node20127 : node20120;
													assign node20120 = (inp[2]) ? node20124 : node20121;
														assign node20121 = (inp[8]) ? 4'b1110 : 4'b1111;
														assign node20124 = (inp[7]) ? 4'b1110 : 4'b1110;
													assign node20127 = (inp[14]) ? 4'b1011 : node20128;
														assign node20128 = (inp[8]) ? 4'b1010 : 4'b1010;
												assign node20132 = (inp[7]) ? node20136 : node20133;
													assign node20133 = (inp[8]) ? 4'b1011 : 4'b1010;
													assign node20136 = (inp[8]) ? 4'b1010 : node20137;
														assign node20137 = (inp[2]) ? 4'b1011 : 4'b1010;
									assign node20141 = (inp[9]) ? node20185 : node20142;
										assign node20142 = (inp[4]) ? node20160 : node20143;
											assign node20143 = (inp[12]) ? node20151 : node20144;
												assign node20144 = (inp[10]) ? node20146 : 4'b1110;
													assign node20146 = (inp[7]) ? node20148 : 4'b1011;
														assign node20148 = (inp[8]) ? 4'b1010 : 4'b1011;
												assign node20151 = (inp[14]) ? node20153 : 4'b1010;
													assign node20153 = (inp[10]) ? node20157 : node20154;
														assign node20154 = (inp[2]) ? 4'b1010 : 4'b1010;
														assign node20157 = (inp[8]) ? 4'b1010 : 4'b1010;
											assign node20160 = (inp[12]) ? node20172 : node20161;
												assign node20161 = (inp[10]) ? node20167 : node20162;
													assign node20162 = (inp[14]) ? node20164 : 4'b1010;
														assign node20164 = (inp[8]) ? 4'b1010 : 4'b1011;
													assign node20167 = (inp[7]) ? node20169 : 4'b1110;
														assign node20169 = (inp[8]) ? 4'b1110 : 4'b1110;
												assign node20172 = (inp[8]) ? node20178 : node20173;
													assign node20173 = (inp[7]) ? 4'b1111 : node20174;
														assign node20174 = (inp[14]) ? 4'b1110 : 4'b1111;
													assign node20178 = (inp[10]) ? node20182 : node20179;
														assign node20179 = (inp[2]) ? 4'b1110 : 4'b1110;
														assign node20182 = (inp[14]) ? 4'b1111 : 4'b1110;
										assign node20185 = (inp[4]) ? node20205 : node20186;
											assign node20186 = (inp[10]) ? node20194 : node20187;
												assign node20187 = (inp[12]) ? node20189 : 4'b1011;
													assign node20189 = (inp[8]) ? 4'b1110 : node20190;
														assign node20190 = (inp[7]) ? 4'b1111 : 4'b1110;
												assign node20194 = (inp[14]) ? node20200 : node20195;
													assign node20195 = (inp[7]) ? 4'b1111 : node20196;
														assign node20196 = (inp[8]) ? 4'b1111 : 4'b1110;
													assign node20200 = (inp[12]) ? node20202 : 4'b1110;
														assign node20202 = (inp[2]) ? 4'b1111 : 4'b1110;
											assign node20205 = (inp[12]) ? node20217 : node20206;
												assign node20206 = (inp[10]) ? node20212 : node20207;
													assign node20207 = (inp[14]) ? node20209 : 4'b1110;
														assign node20209 = (inp[8]) ? 4'b1110 : 4'b1111;
													assign node20212 = (inp[14]) ? node20214 : 4'b1011;
														assign node20214 = (inp[8]) ? 4'b1010 : 4'b1011;
												assign node20217 = (inp[2]) ? node20223 : node20218;
													assign node20218 = (inp[14]) ? 4'b1011 : node20219;
														assign node20219 = (inp[7]) ? 4'b1010 : 4'b1011;
													assign node20223 = (inp[7]) ? node20227 : node20224;
														assign node20224 = (inp[8]) ? 4'b1011 : 4'b1010;
														assign node20227 = (inp[8]) ? 4'b1010 : 4'b1011;
							assign node20230 = (inp[3]) ? node20418 : node20231;
								assign node20231 = (inp[5]) ? node20327 : node20232;
									assign node20232 = (inp[14]) ? node20284 : node20233;
										assign node20233 = (inp[12]) ? node20263 : node20234;
											assign node20234 = (inp[8]) ? node20250 : node20235;
												assign node20235 = (inp[10]) ? node20243 : node20236;
													assign node20236 = (inp[7]) ? node20240 : node20237;
														assign node20237 = (inp[2]) ? 4'b1110 : 4'b1111;
														assign node20240 = (inp[2]) ? 4'b1011 : 4'b1010;
													assign node20243 = (inp[4]) ? node20247 : node20244;
														assign node20244 = (inp[9]) ? 4'b1111 : 4'b1011;
														assign node20247 = (inp[9]) ? 4'b1011 : 4'b1110;
												assign node20250 = (inp[7]) ? node20256 : node20251;
													assign node20251 = (inp[2]) ? 4'b1011 : node20252;
														assign node20252 = (inp[10]) ? 4'b1010 : 4'b1110;
													assign node20256 = (inp[2]) ? node20260 : node20257;
														assign node20257 = (inp[10]) ? 4'b1011 : 4'b1011;
														assign node20260 = (inp[9]) ? 4'b1010 : 4'b1110;
											assign node20263 = (inp[2]) ? node20273 : node20264;
												assign node20264 = (inp[8]) ? node20270 : node20265;
													assign node20265 = (inp[4]) ? 4'b1011 : node20266;
														assign node20266 = (inp[9]) ? 4'b1111 : 4'b1011;
													assign node20270 = (inp[7]) ? 4'b1011 : 4'b1010;
												assign node20273 = (inp[9]) ? node20281 : node20274;
													assign node20274 = (inp[4]) ? node20278 : node20275;
														assign node20275 = (inp[8]) ? 4'b1010 : 4'b1011;
														assign node20278 = (inp[7]) ? 4'b1110 : 4'b1111;
													assign node20281 = (inp[4]) ? 4'b1010 : 4'b1110;
										assign node20284 = (inp[12]) ? node20298 : node20285;
											assign node20285 = (inp[9]) ? node20293 : node20286;
												assign node20286 = (inp[4]) ? node20290 : node20287;
													assign node20287 = (inp[10]) ? 4'b1010 : 4'b1110;
													assign node20290 = (inp[7]) ? 4'b1110 : 4'b1111;
												assign node20293 = (inp[4]) ? 4'b1010 : node20294;
													assign node20294 = (inp[8]) ? 4'b1110 : 4'b1010;
											assign node20298 = (inp[8]) ? node20312 : node20299;
												assign node20299 = (inp[7]) ? node20307 : node20300;
													assign node20300 = (inp[2]) ? node20304 : node20301;
														assign node20301 = (inp[4]) ? 4'b1010 : 4'b1110;
														assign node20304 = (inp[4]) ? 4'b1110 : 4'b1010;
													assign node20307 = (inp[2]) ? node20309 : 4'b1011;
														assign node20309 = (inp[9]) ? 4'b1011 : 4'b1111;
												assign node20312 = (inp[7]) ? node20320 : node20313;
													assign node20313 = (inp[4]) ? node20317 : node20314;
														assign node20314 = (inp[9]) ? 4'b1111 : 4'b1011;
														assign node20317 = (inp[9]) ? 4'b1011 : 4'b1111;
													assign node20320 = (inp[9]) ? node20324 : node20321;
														assign node20321 = (inp[4]) ? 4'b1110 : 4'b1010;
														assign node20324 = (inp[2]) ? 4'b1110 : 4'b1010;
									assign node20327 = (inp[9]) ? node20369 : node20328;
										assign node20328 = (inp[4]) ? node20350 : node20329;
											assign node20329 = (inp[10]) ? node20341 : node20330;
												assign node20330 = (inp[12]) ? node20336 : node20331;
													assign node20331 = (inp[8]) ? node20333 : 4'b1110;
														assign node20333 = (inp[2]) ? 4'b1111 : 4'b1110;
													assign node20336 = (inp[7]) ? node20338 : 4'b1011;
														assign node20338 = (inp[14]) ? 4'b1011 : 4'b1010;
												assign node20341 = (inp[12]) ? 4'b1010 : node20342;
													assign node20342 = (inp[8]) ? node20346 : node20343;
														assign node20343 = (inp[7]) ? 4'b1011 : 4'b1010;
														assign node20346 = (inp[7]) ? 4'b1010 : 4'b1011;
											assign node20350 = (inp[10]) ? node20358 : node20351;
												assign node20351 = (inp[12]) ? 4'b1101 : node20352;
													assign node20352 = (inp[7]) ? 4'b1010 : node20353;
														assign node20353 = (inp[8]) ? 4'b1011 : 4'b1010;
												assign node20358 = (inp[8]) ? node20364 : node20359;
													assign node20359 = (inp[12]) ? 4'b1101 : node20360;
														assign node20360 = (inp[7]) ? 4'b1101 : 4'b1100;
													assign node20364 = (inp[14]) ? node20366 : 4'b1100;
														assign node20366 = (inp[2]) ? 4'b1101 : 4'b1100;
										assign node20369 = (inp[4]) ? node20395 : node20370;
											assign node20370 = (inp[10]) ? node20382 : node20371;
												assign node20371 = (inp[12]) ? node20377 : node20372;
													assign node20372 = (inp[8]) ? node20374 : 4'b1011;
														assign node20374 = (inp[7]) ? 4'b1010 : 4'b1011;
													assign node20377 = (inp[2]) ? node20379 : 4'b1101;
														assign node20379 = (inp[7]) ? 4'b1101 : 4'b1100;
												assign node20382 = (inp[14]) ? node20390 : node20383;
													assign node20383 = (inp[2]) ? node20387 : node20384;
														assign node20384 = (inp[12]) ? 4'b1100 : 4'b1100;
														assign node20387 = (inp[12]) ? 4'b1101 : 4'b1100;
													assign node20390 = (inp[7]) ? 4'b1101 : node20391;
														assign node20391 = (inp[8]) ? 4'b1101 : 4'b1100;
											assign node20395 = (inp[12]) ? node20405 : node20396;
												assign node20396 = (inp[10]) ? node20402 : node20397;
													assign node20397 = (inp[2]) ? 4'b1101 : node20398;
														assign node20398 = (inp[14]) ? 4'b1101 : 4'b1100;
													assign node20402 = (inp[7]) ? 4'b1000 : 4'b1001;
												assign node20405 = (inp[2]) ? node20413 : node20406;
													assign node20406 = (inp[10]) ? node20410 : node20407;
														assign node20407 = (inp[7]) ? 4'b1001 : 4'b1000;
														assign node20410 = (inp[7]) ? 4'b1000 : 4'b1001;
													assign node20413 = (inp[7]) ? node20415 : 4'b1000;
														assign node20415 = (inp[8]) ? 4'b1000 : 4'b1001;
								assign node20418 = (inp[5]) ? node20504 : node20419;
									assign node20419 = (inp[9]) ? node20459 : node20420;
										assign node20420 = (inp[4]) ? node20446 : node20421;
											assign node20421 = (inp[10]) ? node20435 : node20422;
												assign node20422 = (inp[12]) ? node20430 : node20423;
													assign node20423 = (inp[8]) ? node20427 : node20424;
														assign node20424 = (inp[14]) ? 4'b1110 : 4'b1111;
														assign node20427 = (inp[2]) ? 4'b1110 : 4'b1110;
													assign node20430 = (inp[2]) ? 4'b1011 : node20431;
														assign node20431 = (inp[8]) ? 4'b1010 : 4'b1011;
												assign node20435 = (inp[2]) ? node20441 : node20436;
													assign node20436 = (inp[7]) ? node20438 : 4'b1011;
														assign node20438 = (inp[8]) ? 4'b1010 : 4'b1010;
													assign node20441 = (inp[14]) ? node20443 : 4'b1010;
														assign node20443 = (inp[8]) ? 4'b1010 : 4'b1011;
											assign node20446 = (inp[10]) ? node20454 : node20447;
												assign node20447 = (inp[12]) ? node20451 : node20448;
													assign node20448 = (inp[7]) ? 4'b1011 : 4'b1010;
													assign node20451 = (inp[2]) ? 4'b1100 : 4'b1101;
												assign node20454 = (inp[7]) ? node20456 : 4'b1101;
													assign node20456 = (inp[8]) ? 4'b1100 : 4'b1101;
										assign node20459 = (inp[4]) ? node20487 : node20460;
											assign node20460 = (inp[12]) ? node20474 : node20461;
												assign node20461 = (inp[10]) ? node20467 : node20462;
													assign node20462 = (inp[14]) ? node20464 : 4'b1011;
														assign node20464 = (inp[8]) ? 4'b1010 : 4'b1010;
													assign node20467 = (inp[14]) ? node20471 : node20468;
														assign node20468 = (inp[2]) ? 4'b1100 : 4'b1100;
														assign node20471 = (inp[8]) ? 4'b1100 : 4'b1101;
												assign node20474 = (inp[10]) ? node20480 : node20475;
													assign node20475 = (inp[14]) ? node20477 : 4'b1101;
														assign node20477 = (inp[8]) ? 4'b1101 : 4'b1101;
													assign node20480 = (inp[7]) ? node20484 : node20481;
														assign node20481 = (inp[8]) ? 4'b1101 : 4'b1100;
														assign node20484 = (inp[8]) ? 4'b1100 : 4'b1101;
											assign node20487 = (inp[10]) ? node20495 : node20488;
												assign node20488 = (inp[12]) ? 4'b1001 : node20489;
													assign node20489 = (inp[7]) ? 4'b1100 : node20490;
														assign node20490 = (inp[2]) ? 4'b1100 : 4'b1101;
												assign node20495 = (inp[14]) ? node20497 : 4'b1000;
													assign node20497 = (inp[8]) ? node20501 : node20498;
														assign node20498 = (inp[7]) ? 4'b1001 : 4'b1000;
														assign node20501 = (inp[7]) ? 4'b1000 : 4'b1001;
									assign node20504 = (inp[12]) ? node20546 : node20505;
										assign node20505 = (inp[14]) ? node20527 : node20506;
											assign node20506 = (inp[8]) ? node20516 : node20507;
												assign node20507 = (inp[2]) ? node20511 : node20508;
													assign node20508 = (inp[7]) ? 4'b1100 : 4'b1101;
													assign node20511 = (inp[7]) ? 4'b1001 : node20512;
														assign node20512 = (inp[10]) ? 4'b1000 : 4'b1000;
												assign node20516 = (inp[7]) ? node20522 : node20517;
													assign node20517 = (inp[2]) ? 4'b1001 : node20518;
														assign node20518 = (inp[9]) ? 4'b1100 : 4'b1000;
													assign node20522 = (inp[2]) ? node20524 : 4'b1001;
														assign node20524 = (inp[9]) ? 4'b1100 : 4'b1000;
											assign node20527 = (inp[7]) ? node20535 : node20528;
												assign node20528 = (inp[8]) ? node20530 : 4'b1100;
													assign node20530 = (inp[9]) ? node20532 : 4'b1101;
														assign node20532 = (inp[4]) ? 4'b1101 : 4'b1001;
												assign node20535 = (inp[8]) ? node20541 : node20536;
													assign node20536 = (inp[9]) ? node20538 : 4'b1001;
														assign node20538 = (inp[10]) ? 4'b1101 : 4'b1001;
													assign node20541 = (inp[2]) ? 4'b1100 : node20542;
														assign node20542 = (inp[10]) ? 4'b1100 : 4'b1000;
										assign node20546 = (inp[2]) ? node20570 : node20547;
											assign node20547 = (inp[4]) ? node20557 : node20548;
												assign node20548 = (inp[9]) ? node20554 : node20549;
													assign node20549 = (inp[7]) ? node20551 : 4'b1001;
														assign node20551 = (inp[14]) ? 4'b1000 : 4'b1001;
													assign node20554 = (inp[14]) ? 4'b1100 : 4'b1101;
												assign node20557 = (inp[9]) ? node20563 : node20558;
													assign node20558 = (inp[7]) ? node20560 : 4'b1100;
														assign node20560 = (inp[14]) ? 4'b1100 : 4'b1101;
													assign node20563 = (inp[7]) ? node20567 : node20564;
														assign node20564 = (inp[14]) ? 4'b1000 : 4'b1000;
														assign node20567 = (inp[8]) ? 4'b1001 : 4'b1000;
											assign node20570 = (inp[14]) ? node20586 : node20571;
												assign node20571 = (inp[10]) ? node20579 : node20572;
													assign node20572 = (inp[8]) ? node20576 : node20573;
														assign node20573 = (inp[7]) ? 4'b1101 : 4'b1000;
														assign node20576 = (inp[7]) ? 4'b1000 : 4'b1001;
													assign node20579 = (inp[4]) ? node20583 : node20580;
														assign node20580 = (inp[9]) ? 4'b1100 : 4'b1000;
														assign node20583 = (inp[8]) ? 4'b1101 : 4'b1100;
												assign node20586 = (inp[7]) ? node20592 : node20587;
													assign node20587 = (inp[8]) ? node20589 : 4'b1000;
														assign node20589 = (inp[4]) ? 4'b1001 : 4'b1001;
													assign node20592 = (inp[9]) ? 4'b1101 : node20593;
														assign node20593 = (inp[4]) ? 4'b1101 : 4'b1001;
						assign node20597 = (inp[8]) ? node20963 : node20598;
							assign node20598 = (inp[7]) ? node20776 : node20599;
								assign node20599 = (inp[14]) ? node20699 : node20600;
									assign node20600 = (inp[2]) ? node20648 : node20601;
										assign node20601 = (inp[4]) ? node20625 : node20602;
											assign node20602 = (inp[15]) ? node20614 : node20603;
												assign node20603 = (inp[5]) ? node20609 : node20604;
													assign node20604 = (inp[12]) ? 4'b1001 : node20605;
														assign node20605 = (inp[10]) ? 4'b1101 : 4'b1001;
													assign node20609 = (inp[9]) ? 4'b1001 : node20610;
														assign node20610 = (inp[10]) ? 4'b1011 : 4'b1111;
												assign node20614 = (inp[3]) ? node20620 : node20615;
													assign node20615 = (inp[12]) ? 4'b1011 : node20616;
														assign node20616 = (inp[10]) ? 4'b1011 : 4'b1011;
													assign node20620 = (inp[12]) ? node20622 : 4'b1011;
														assign node20622 = (inp[9]) ? 4'b1101 : 4'b1001;
											assign node20625 = (inp[9]) ? node20637 : node20626;
												assign node20626 = (inp[10]) ? node20632 : node20627;
													assign node20627 = (inp[12]) ? 4'b1111 : node20628;
														assign node20628 = (inp[15]) ? 4'b1011 : 4'b1001;
													assign node20632 = (inp[15]) ? 4'b1101 : node20633;
														assign node20633 = (inp[3]) ? 4'b1111 : 4'b1101;
												assign node20637 = (inp[12]) ? node20643 : node20638;
													assign node20638 = (inp[10]) ? 4'b1011 : node20639;
														assign node20639 = (inp[5]) ? 4'b1111 : 4'b1101;
													assign node20643 = (inp[15]) ? 4'b1001 : node20644;
														assign node20644 = (inp[3]) ? 4'b1011 : 4'b1001;
										assign node20648 = (inp[15]) ? node20674 : node20649;
											assign node20649 = (inp[3]) ? node20663 : node20650;
												assign node20650 = (inp[5]) ? node20656 : node20651;
													assign node20651 = (inp[12]) ? 4'b1100 : node20652;
														assign node20652 = (inp[4]) ? 4'b1000 : 4'b1000;
													assign node20656 = (inp[4]) ? node20660 : node20657;
														assign node20657 = (inp[9]) ? 4'b1110 : 4'b1000;
														assign node20660 = (inp[10]) ? 4'b1010 : 4'b1110;
												assign node20663 = (inp[12]) ? node20669 : node20664;
													assign node20664 = (inp[9]) ? 4'b1110 : node20665;
														assign node20665 = (inp[5]) ? 4'b1010 : 4'b1000;
													assign node20669 = (inp[9]) ? node20671 : 4'b1110;
														assign node20671 = (inp[4]) ? 4'b1010 : 4'b1110;
											assign node20674 = (inp[3]) ? node20686 : node20675;
												assign node20675 = (inp[5]) ? node20679 : node20676;
													assign node20676 = (inp[4]) ? 4'b1110 : 4'b1010;
													assign node20679 = (inp[10]) ? node20683 : node20680;
														assign node20680 = (inp[4]) ? 4'b1000 : 4'b1010;
														assign node20683 = (inp[12]) ? 4'b1100 : 4'b1000;
												assign node20686 = (inp[12]) ? node20692 : node20687;
													assign node20687 = (inp[10]) ? 4'b1100 : node20688;
														assign node20688 = (inp[9]) ? 4'b1100 : 4'b1010;
													assign node20692 = (inp[4]) ? node20696 : node20693;
														assign node20693 = (inp[9]) ? 4'b1100 : 4'b1000;
														assign node20696 = (inp[9]) ? 4'b1000 : 4'b1100;
									assign node20699 = (inp[15]) ? node20739 : node20700;
										assign node20700 = (inp[5]) ? node20726 : node20701;
											assign node20701 = (inp[3]) ? node20715 : node20702;
												assign node20702 = (inp[4]) ? node20708 : node20703;
													assign node20703 = (inp[10]) ? 4'b1000 : node20704;
														assign node20704 = (inp[12]) ? 4'b1100 : 4'b1100;
													assign node20708 = (inp[10]) ? node20712 : node20709;
														assign node20709 = (inp[2]) ? 4'b1000 : 4'b1000;
														assign node20712 = (inp[9]) ? 4'b1000 : 4'b1100;
												assign node20715 = (inp[9]) ? node20723 : node20716;
													assign node20716 = (inp[4]) ? node20720 : node20717;
														assign node20717 = (inp[10]) ? 4'b1000 : 4'b1100;
														assign node20720 = (inp[10]) ? 4'b1110 : 4'b1000;
													assign node20723 = (inp[4]) ? 4'b1010 : 4'b1110;
											assign node20726 = (inp[4]) ? node20734 : node20727;
												assign node20727 = (inp[9]) ? 4'b1110 : node20728;
													assign node20728 = (inp[3]) ? node20730 : 4'b1000;
														assign node20730 = (inp[10]) ? 4'b1010 : 4'b1110;
												assign node20734 = (inp[9]) ? node20736 : 4'b1110;
													assign node20736 = (inp[10]) ? 4'b1010 : 4'b1110;
										assign node20739 = (inp[3]) ? node20755 : node20740;
											assign node20740 = (inp[5]) ? node20748 : node20741;
												assign node20741 = (inp[9]) ? node20743 : 4'b1110;
													assign node20743 = (inp[12]) ? 4'b1010 : node20744;
														assign node20744 = (inp[10]) ? 4'b1010 : 4'b1110;
												assign node20748 = (inp[10]) ? 4'b1100 : node20749;
													assign node20749 = (inp[4]) ? node20751 : 4'b1010;
														assign node20751 = (inp[9]) ? 4'b1100 : 4'b1000;
											assign node20755 = (inp[5]) ? node20767 : node20756;
												assign node20756 = (inp[4]) ? node20762 : node20757;
													assign node20757 = (inp[9]) ? node20759 : 4'b1010;
														assign node20759 = (inp[12]) ? 4'b1100 : 4'b1000;
													assign node20762 = (inp[9]) ? node20764 : 4'b1100;
														assign node20764 = (inp[10]) ? 4'b1000 : 4'b1100;
												assign node20767 = (inp[9]) ? node20773 : node20768;
													assign node20768 = (inp[4]) ? node20770 : 4'b1000;
														assign node20770 = (inp[12]) ? 4'b1100 : 4'b1000;
													assign node20773 = (inp[4]) ? 4'b1000 : 4'b1100;
								assign node20776 = (inp[14]) ? node20872 : node20777;
									assign node20777 = (inp[2]) ? node20827 : node20778;
										assign node20778 = (inp[15]) ? node20800 : node20779;
											assign node20779 = (inp[5]) ? node20787 : node20780;
												assign node20780 = (inp[9]) ? 4'b1110 : node20781;
													assign node20781 = (inp[3]) ? 4'b1000 : node20782;
														assign node20782 = (inp[10]) ? 4'b1100 : 4'b1000;
												assign node20787 = (inp[9]) ? node20793 : node20788;
													assign node20788 = (inp[4]) ? 4'b1110 : node20789;
														assign node20789 = (inp[12]) ? 4'b1010 : 4'b1110;
													assign node20793 = (inp[4]) ? node20797 : node20794;
														assign node20794 = (inp[12]) ? 4'b1110 : 4'b1000;
														assign node20797 = (inp[10]) ? 4'b1010 : 4'b1010;
											assign node20800 = (inp[5]) ? node20812 : node20801;
												assign node20801 = (inp[3]) ? node20807 : node20802;
													assign node20802 = (inp[12]) ? node20804 : 4'b1010;
														assign node20804 = (inp[4]) ? 4'b1010 : 4'b1010;
													assign node20807 = (inp[9]) ? 4'b1100 : node20808;
														assign node20808 = (inp[10]) ? 4'b1010 : 4'b1100;
												assign node20812 = (inp[12]) ? node20820 : node20813;
													assign node20813 = (inp[10]) ? node20817 : node20814;
														assign node20814 = (inp[3]) ? 4'b1100 : 4'b1010;
														assign node20817 = (inp[4]) ? 4'b1100 : 4'b1000;
													assign node20820 = (inp[3]) ? node20824 : node20821;
														assign node20821 = (inp[4]) ? 4'b1100 : 4'b1100;
														assign node20824 = (inp[9]) ? 4'b1000 : 4'b1000;
										assign node20827 = (inp[3]) ? node20851 : node20828;
											assign node20828 = (inp[15]) ? node20840 : node20829;
												assign node20829 = (inp[5]) ? node20835 : node20830;
													assign node20830 = (inp[10]) ? node20832 : 4'b0001;
														assign node20832 = (inp[4]) ? 4'b0001 : 4'b0001;
													assign node20835 = (inp[4]) ? node20837 : 4'b0111;
														assign node20837 = (inp[9]) ? 4'b0011 : 4'b0111;
												assign node20840 = (inp[5]) ? node20846 : node20841;
													assign node20841 = (inp[9]) ? 4'b0111 : node20842;
														assign node20842 = (inp[4]) ? 4'b0111 : 4'b0011;
													assign node20846 = (inp[9]) ? 4'b0001 : node20847;
														assign node20847 = (inp[10]) ? 4'b0001 : 4'b0011;
											assign node20851 = (inp[15]) ? node20859 : node20852;
												assign node20852 = (inp[9]) ? node20856 : node20853;
													assign node20853 = (inp[12]) ? 4'b0001 : 4'b0101;
													assign node20856 = (inp[4]) ? 4'b0011 : 4'b0111;
												assign node20859 = (inp[5]) ? node20867 : node20860;
													assign node20860 = (inp[12]) ? node20864 : node20861;
														assign node20861 = (inp[10]) ? 4'b0101 : 4'b0111;
														assign node20864 = (inp[4]) ? 4'b0001 : 4'b0011;
													assign node20867 = (inp[10]) ? node20869 : 4'b0101;
														assign node20869 = (inp[9]) ? 4'b0101 : 4'b0001;
									assign node20872 = (inp[2]) ? node20916 : node20873;
										assign node20873 = (inp[12]) ? node20893 : node20874;
											assign node20874 = (inp[9]) ? node20886 : node20875;
												assign node20875 = (inp[10]) ? node20881 : node20876;
													assign node20876 = (inp[4]) ? node20878 : 4'b0101;
														assign node20878 = (inp[15]) ? 4'b0011 : 4'b0001;
													assign node20881 = (inp[4]) ? 4'b0111 : node20882;
														assign node20882 = (inp[15]) ? 4'b0001 : 4'b0001;
												assign node20886 = (inp[15]) ? node20888 : 4'b0011;
													assign node20888 = (inp[10]) ? node20890 : 4'b0011;
														assign node20890 = (inp[3]) ? 4'b0001 : 4'b0011;
											assign node20893 = (inp[3]) ? node20907 : node20894;
												assign node20894 = (inp[15]) ? node20900 : node20895;
													assign node20895 = (inp[10]) ? node20897 : 4'b0001;
														assign node20897 = (inp[9]) ? 4'b0111 : 4'b0001;
													assign node20900 = (inp[9]) ? node20904 : node20901;
														assign node20901 = (inp[4]) ? 4'b0111 : 4'b0011;
														assign node20904 = (inp[5]) ? 4'b0101 : 4'b0011;
												assign node20907 = (inp[15]) ? node20913 : node20908;
													assign node20908 = (inp[4]) ? 4'b0111 : node20909;
														assign node20909 = (inp[9]) ? 4'b0111 : 4'b0001;
													assign node20913 = (inp[4]) ? 4'b0001 : 4'b0101;
										assign node20916 = (inp[10]) ? node20940 : node20917;
											assign node20917 = (inp[12]) ? node20929 : node20918;
												assign node20918 = (inp[4]) ? node20922 : node20919;
													assign node20919 = (inp[9]) ? 4'b0001 : 4'b0101;
													assign node20922 = (inp[9]) ? node20926 : node20923;
														assign node20923 = (inp[15]) ? 4'b0011 : 4'b0001;
														assign node20926 = (inp[15]) ? 4'b0101 : 4'b0101;
												assign node20929 = (inp[3]) ? node20937 : node20930;
													assign node20930 = (inp[9]) ? node20934 : node20931;
														assign node20931 = (inp[4]) ? 4'b0101 : 4'b0011;
														assign node20934 = (inp[4]) ? 4'b0001 : 4'b0101;
													assign node20937 = (inp[15]) ? 4'b0001 : 4'b0011;
											assign node20940 = (inp[4]) ? node20950 : node20941;
												assign node20941 = (inp[9]) ? node20945 : node20942;
													assign node20942 = (inp[15]) ? 4'b0011 : 4'b0001;
													assign node20945 = (inp[15]) ? node20947 : 4'b0111;
														assign node20947 = (inp[3]) ? 4'b0101 : 4'b0111;
												assign node20950 = (inp[9]) ? node20958 : node20951;
													assign node20951 = (inp[5]) ? node20955 : node20952;
														assign node20952 = (inp[12]) ? 4'b0101 : 4'b0101;
														assign node20955 = (inp[15]) ? 4'b0101 : 4'b0111;
													assign node20958 = (inp[5]) ? node20960 : 4'b0001;
														assign node20960 = (inp[3]) ? 4'b0011 : 4'b0001;
							assign node20963 = (inp[7]) ? node21139 : node20964;
								assign node20964 = (inp[14]) ? node21056 : node20965;
									assign node20965 = (inp[2]) ? node21015 : node20966;
										assign node20966 = (inp[5]) ? node20994 : node20967;
											assign node20967 = (inp[3]) ? node20981 : node20968;
												assign node20968 = (inp[10]) ? node20974 : node20969;
													assign node20969 = (inp[4]) ? node20971 : 4'b1010;
														assign node20971 = (inp[9]) ? 4'b1110 : 4'b1010;
													assign node20974 = (inp[4]) ? node20978 : node20975;
														assign node20975 = (inp[9]) ? 4'b1110 : 4'b1010;
														assign node20978 = (inp[9]) ? 4'b1010 : 4'b1110;
												assign node20981 = (inp[15]) ? node20987 : node20982;
													assign node20982 = (inp[4]) ? node20984 : 4'b1000;
														assign node20984 = (inp[12]) ? 4'b1010 : 4'b1110;
													assign node20987 = (inp[4]) ? node20991 : node20988;
														assign node20988 = (inp[9]) ? 4'b1100 : 4'b1010;
														assign node20991 = (inp[9]) ? 4'b1000 : 4'b1100;
											assign node20994 = (inp[10]) ? node21010 : node20995;
												assign node20995 = (inp[12]) ? node21003 : node20996;
													assign node20996 = (inp[9]) ? node21000 : node20997;
														assign node20997 = (inp[4]) ? 4'b1000 : 4'b1110;
														assign node21000 = (inp[15]) ? 4'b1000 : 4'b1110;
													assign node21003 = (inp[9]) ? node21007 : node21004;
														assign node21004 = (inp[4]) ? 4'b1100 : 4'b1010;
														assign node21007 = (inp[4]) ? 4'b1000 : 4'b1100;
												assign node21010 = (inp[3]) ? node21012 : 4'b1000;
													assign node21012 = (inp[15]) ? 4'b1000 : 4'b1010;
										assign node21015 = (inp[9]) ? node21041 : node21016;
											assign node21016 = (inp[3]) ? node21030 : node21017;
												assign node21017 = (inp[15]) ? node21023 : node21018;
													assign node21018 = (inp[4]) ? 4'b0111 : node21019;
														assign node21019 = (inp[10]) ? 4'b0001 : 4'b0101;
													assign node21023 = (inp[4]) ? node21027 : node21024;
														assign node21024 = (inp[5]) ? 4'b0011 : 4'b0011;
														assign node21027 = (inp[12]) ? 4'b0111 : 4'b0011;
												assign node21030 = (inp[5]) ? node21036 : node21031;
													assign node21031 = (inp[12]) ? 4'b0001 : node21032;
														assign node21032 = (inp[4]) ? 4'b0001 : 4'b0101;
													assign node21036 = (inp[10]) ? 4'b0111 : node21037;
														assign node21037 = (inp[12]) ? 4'b0101 : 4'b0001;
											assign node21041 = (inp[4]) ? node21053 : node21042;
												assign node21042 = (inp[10]) ? node21046 : node21043;
													assign node21043 = (inp[12]) ? 4'b0101 : 4'b0011;
													assign node21046 = (inp[15]) ? node21050 : node21047;
														assign node21047 = (inp[3]) ? 4'b0111 : 4'b0111;
														assign node21050 = (inp[5]) ? 4'b0101 : 4'b0111;
												assign node21053 = (inp[3]) ? 4'b0011 : 4'b0001;
									assign node21056 = (inp[4]) ? node21100 : node21057;
										assign node21057 = (inp[9]) ? node21081 : node21058;
											assign node21058 = (inp[10]) ? node21070 : node21059;
												assign node21059 = (inp[12]) ? node21065 : node21060;
													assign node21060 = (inp[2]) ? 4'b0101 : node21061;
														assign node21061 = (inp[15]) ? 4'b0111 : 4'b0101;
													assign node21065 = (inp[3]) ? node21067 : 4'b0001;
														assign node21067 = (inp[2]) ? 4'b0011 : 4'b0001;
												assign node21070 = (inp[15]) ? node21076 : node21071;
													assign node21071 = (inp[3]) ? node21073 : 4'b0001;
														assign node21073 = (inp[5]) ? 4'b0011 : 4'b0001;
													assign node21076 = (inp[5]) ? node21078 : 4'b0011;
														assign node21078 = (inp[2]) ? 4'b0011 : 4'b0001;
											assign node21081 = (inp[5]) ? node21093 : node21082;
												assign node21082 = (inp[2]) ? node21086 : node21083;
													assign node21083 = (inp[10]) ? 4'b0101 : 4'b0001;
													assign node21086 = (inp[10]) ? node21090 : node21087;
														assign node21087 = (inp[15]) ? 4'b0111 : 4'b0101;
														assign node21090 = (inp[12]) ? 4'b0101 : 4'b0101;
												assign node21093 = (inp[15]) ? node21095 : 4'b0111;
													assign node21095 = (inp[10]) ? 4'b0101 : node21096;
														assign node21096 = (inp[12]) ? 4'b0101 : 4'b0011;
										assign node21100 = (inp[9]) ? node21116 : node21101;
											assign node21101 = (inp[10]) ? 4'b0111 : node21102;
												assign node21102 = (inp[12]) ? node21110 : node21103;
													assign node21103 = (inp[3]) ? node21107 : node21104;
														assign node21104 = (inp[5]) ? 4'b0001 : 4'b0011;
														assign node21107 = (inp[15]) ? 4'b0001 : 4'b0001;
													assign node21110 = (inp[5]) ? 4'b0101 : node21111;
														assign node21111 = (inp[15]) ? 4'b0111 : 4'b0101;
											assign node21116 = (inp[10]) ? node21128 : node21117;
												assign node21117 = (inp[12]) ? node21123 : node21118;
													assign node21118 = (inp[15]) ? node21120 : 4'b0101;
														assign node21120 = (inp[5]) ? 4'b0101 : 4'b0111;
													assign node21123 = (inp[15]) ? node21125 : 4'b0011;
														assign node21125 = (inp[2]) ? 4'b0011 : 4'b0001;
												assign node21128 = (inp[15]) ? node21134 : node21129;
													assign node21129 = (inp[3]) ? 4'b0011 : node21130;
														assign node21130 = (inp[5]) ? 4'b0011 : 4'b0001;
													assign node21134 = (inp[5]) ? 4'b0001 : node21135;
														assign node21135 = (inp[3]) ? 4'b0001 : 4'b0011;
								assign node21139 = (inp[2]) ? node21219 : node21140;
									assign node21140 = (inp[14]) ? node21186 : node21141;
										assign node21141 = (inp[15]) ? node21163 : node21142;
											assign node21142 = (inp[3]) ? node21152 : node21143;
												assign node21143 = (inp[9]) ? node21149 : node21144;
													assign node21144 = (inp[10]) ? 4'b0001 : node21145;
														assign node21145 = (inp[5]) ? 4'b0001 : 4'b0101;
													assign node21149 = (inp[12]) ? 4'b0111 : 4'b0101;
												assign node21152 = (inp[10]) ? node21158 : node21153;
													assign node21153 = (inp[9]) ? 4'b0111 : node21154;
														assign node21154 = (inp[5]) ? 4'b0011 : 4'b0111;
													assign node21158 = (inp[12]) ? node21160 : 4'b0011;
														assign node21160 = (inp[5]) ? 4'b0011 : 4'b0011;
											assign node21163 = (inp[3]) ? node21175 : node21164;
												assign node21164 = (inp[5]) ? node21170 : node21165;
													assign node21165 = (inp[4]) ? 4'b0011 : node21166;
														assign node21166 = (inp[10]) ? 4'b0111 : 4'b0011;
													assign node21170 = (inp[4]) ? 4'b0101 : node21171;
														assign node21171 = (inp[9]) ? 4'b0101 : 4'b0011;
												assign node21175 = (inp[4]) ? node21181 : node21176;
													assign node21176 = (inp[5]) ? node21178 : 4'b0101;
														assign node21178 = (inp[9]) ? 4'b0001 : 4'b0001;
													assign node21181 = (inp[9]) ? 4'b0001 : node21182;
														assign node21182 = (inp[12]) ? 4'b0101 : 4'b0011;
										assign node21186 = (inp[15]) ? node21208 : node21187;
											assign node21187 = (inp[10]) ? node21199 : node21188;
												assign node21188 = (inp[12]) ? node21194 : node21189;
													assign node21189 = (inp[4]) ? 4'b0000 : node21190;
														assign node21190 = (inp[5]) ? 4'b0000 : 4'b0100;
													assign node21194 = (inp[9]) ? node21196 : 4'b0000;
														assign node21196 = (inp[4]) ? 4'b0010 : 4'b0110;
												assign node21199 = (inp[3]) ? node21201 : 4'b0110;
													assign node21201 = (inp[5]) ? node21205 : node21202;
														assign node21202 = (inp[4]) ? 4'b0110 : 4'b0110;
														assign node21205 = (inp[4]) ? 4'b0010 : 4'b0010;
											assign node21208 = (inp[9]) ? 4'b0100 : node21209;
												assign node21209 = (inp[10]) ? node21215 : node21210;
													assign node21210 = (inp[3]) ? 4'b0100 : node21211;
														assign node21211 = (inp[4]) ? 4'b0100 : 4'b0110;
													assign node21215 = (inp[3]) ? 4'b0000 : 4'b0010;
									assign node21219 = (inp[14]) ? node21267 : node21220;
										assign node21220 = (inp[15]) ? node21244 : node21221;
											assign node21221 = (inp[5]) ? node21235 : node21222;
												assign node21222 = (inp[12]) ? node21230 : node21223;
													assign node21223 = (inp[3]) ? node21227 : node21224;
														assign node21224 = (inp[9]) ? 4'b0100 : 4'b0100;
														assign node21227 = (inp[4]) ? 4'b0110 : 4'b0000;
													assign node21230 = (inp[9]) ? 4'b0000 : node21231;
														assign node21231 = (inp[4]) ? 4'b0100 : 4'b0000;
												assign node21235 = (inp[3]) ? node21241 : node21236;
													assign node21236 = (inp[12]) ? node21238 : 4'b0000;
														assign node21238 = (inp[4]) ? 4'b0010 : 4'b0110;
													assign node21241 = (inp[12]) ? 4'b0010 : 4'b0110;
											assign node21244 = (inp[5]) ? node21254 : node21245;
												assign node21245 = (inp[4]) ? node21251 : node21246;
													assign node21246 = (inp[9]) ? 4'b0110 : node21247;
														assign node21247 = (inp[10]) ? 4'b0010 : 4'b0010;
													assign node21251 = (inp[3]) ? 4'b0100 : 4'b0110;
												assign node21254 = (inp[9]) ? node21262 : node21255;
													assign node21255 = (inp[3]) ? node21259 : node21256;
														assign node21256 = (inp[4]) ? 4'b0010 : 4'b0110;
														assign node21259 = (inp[12]) ? 4'b0100 : 4'b0000;
													assign node21262 = (inp[10]) ? node21264 : 4'b0100;
														assign node21264 = (inp[4]) ? 4'b0000 : 4'b0100;
										assign node21267 = (inp[9]) ? node21293 : node21268;
											assign node21268 = (inp[4]) ? node21280 : node21269;
												assign node21269 = (inp[12]) ? node21275 : node21270;
													assign node21270 = (inp[10]) ? node21272 : 4'b0100;
														assign node21272 = (inp[3]) ? 4'b0010 : 4'b0000;
													assign node21275 = (inp[10]) ? node21277 : 4'b0010;
														assign node21277 = (inp[15]) ? 4'b0010 : 4'b0000;
												assign node21280 = (inp[10]) ? node21288 : node21281;
													assign node21281 = (inp[12]) ? node21285 : node21282;
														assign node21282 = (inp[3]) ? 4'b0000 : 4'b0010;
														assign node21285 = (inp[3]) ? 4'b0110 : 4'b0100;
													assign node21288 = (inp[15]) ? 4'b0100 : node21289;
														assign node21289 = (inp[12]) ? 4'b0110 : 4'b0100;
											assign node21293 = (inp[15]) ? node21307 : node21294;
												assign node21294 = (inp[4]) ? node21302 : node21295;
													assign node21295 = (inp[5]) ? node21299 : node21296;
														assign node21296 = (inp[3]) ? 4'b0110 : 4'b0100;
														assign node21299 = (inp[3]) ? 4'b0010 : 4'b0110;
													assign node21302 = (inp[10]) ? 4'b0010 : node21303;
														assign node21303 = (inp[12]) ? 4'b0010 : 4'b0110;
												assign node21307 = (inp[3]) ? node21315 : node21308;
													assign node21308 = (inp[5]) ? node21312 : node21309;
														assign node21309 = (inp[4]) ? 4'b0010 : 4'b0110;
														assign node21312 = (inp[4]) ? 4'b0000 : 4'b0010;
													assign node21315 = (inp[12]) ? 4'b0000 : node21316;
														assign node21316 = (inp[5]) ? 4'b0000 : 4'b0100;
					assign node21320 = (inp[13]) ? node22022 : node21321;
						assign node21321 = (inp[8]) ? node21693 : node21322;
							assign node21322 = (inp[7]) ? node21510 : node21323;
								assign node21323 = (inp[14]) ? node21419 : node21324;
									assign node21324 = (inp[2]) ? node21376 : node21325;
										assign node21325 = (inp[5]) ? node21351 : node21326;
											assign node21326 = (inp[4]) ? node21340 : node21327;
												assign node21327 = (inp[15]) ? node21333 : node21328;
													assign node21328 = (inp[3]) ? 4'b1111 : node21329;
														assign node21329 = (inp[10]) ? 4'b1101 : 4'b1001;
													assign node21333 = (inp[3]) ? node21337 : node21334;
														assign node21334 = (inp[9]) ? 4'b1111 : 4'b1011;
														assign node21337 = (inp[9]) ? 4'b1101 : 4'b1111;
												assign node21340 = (inp[9]) ? node21348 : node21341;
													assign node21341 = (inp[15]) ? node21345 : node21342;
														assign node21342 = (inp[3]) ? 4'b1111 : 4'b1101;
														assign node21345 = (inp[12]) ? 4'b1111 : 4'b1011;
													assign node21348 = (inp[15]) ? 4'b1001 : 4'b1011;
											assign node21351 = (inp[15]) ? node21361 : node21352;
												assign node21352 = (inp[4]) ? node21356 : node21353;
													assign node21353 = (inp[3]) ? 4'b1011 : 4'b1001;
													assign node21356 = (inp[9]) ? node21358 : 4'b1111;
														assign node21358 = (inp[12]) ? 4'b1011 : 4'b1111;
												assign node21361 = (inp[3]) ? node21369 : node21362;
													assign node21362 = (inp[4]) ? node21366 : node21363;
														assign node21363 = (inp[12]) ? 4'b1001 : 4'b1011;
														assign node21366 = (inp[9]) ? 4'b1001 : 4'b1101;
													assign node21369 = (inp[4]) ? node21373 : node21370;
														assign node21370 = (inp[10]) ? 4'b1001 : 4'b1001;
														assign node21373 = (inp[10]) ? 4'b1001 : 4'b1001;
										assign node21376 = (inp[5]) ? node21398 : node21377;
											assign node21377 = (inp[3]) ? node21385 : node21378;
												assign node21378 = (inp[15]) ? node21380 : 4'b1100;
													assign node21380 = (inp[10]) ? node21382 : 4'b1110;
														assign node21382 = (inp[12]) ? 4'b1010 : 4'b1010;
												assign node21385 = (inp[4]) ? node21393 : node21386;
													assign node21386 = (inp[12]) ? node21390 : node21387;
														assign node21387 = (inp[15]) ? 4'b1110 : 4'b1000;
														assign node21390 = (inp[9]) ? 4'b1110 : 4'b1010;
													assign node21393 = (inp[10]) ? 4'b1000 : node21394;
														assign node21394 = (inp[15]) ? 4'b1000 : 4'b1010;
											assign node21398 = (inp[15]) ? node21406 : node21399;
												assign node21399 = (inp[10]) ? 4'b1010 : node21400;
													assign node21400 = (inp[12]) ? 4'b1110 : node21401;
														assign node21401 = (inp[4]) ? 4'b1110 : 4'b1000;
												assign node21406 = (inp[10]) ? node21414 : node21407;
													assign node21407 = (inp[12]) ? node21411 : node21408;
														assign node21408 = (inp[4]) ? 4'b1010 : 4'b1110;
														assign node21411 = (inp[9]) ? 4'b1100 : 4'b1000;
													assign node21414 = (inp[9]) ? node21416 : 4'b1100;
														assign node21416 = (inp[4]) ? 4'b1000 : 4'b1100;
									assign node21419 = (inp[5]) ? node21463 : node21420;
										assign node21420 = (inp[15]) ? node21442 : node21421;
											assign node21421 = (inp[3]) ? node21431 : node21422;
												assign node21422 = (inp[12]) ? node21424 : 4'b1000;
													assign node21424 = (inp[4]) ? node21428 : node21425;
														assign node21425 = (inp[9]) ? 4'b1100 : 4'b1000;
														assign node21428 = (inp[9]) ? 4'b1000 : 4'b1100;
												assign node21431 = (inp[9]) ? node21437 : node21432;
													assign node21432 = (inp[4]) ? 4'b1110 : node21433;
														assign node21433 = (inp[12]) ? 4'b1000 : 4'b1100;
													assign node21437 = (inp[4]) ? node21439 : 4'b1110;
														assign node21439 = (inp[12]) ? 4'b1010 : 4'b1110;
											assign node21442 = (inp[4]) ? node21452 : node21443;
												assign node21443 = (inp[10]) ? node21449 : node21444;
													assign node21444 = (inp[12]) ? node21446 : 4'b1110;
														assign node21446 = (inp[9]) ? 4'b1110 : 4'b1010;
													assign node21449 = (inp[9]) ? 4'b1110 : 4'b1010;
												assign node21452 = (inp[3]) ? node21458 : node21453;
													assign node21453 = (inp[12]) ? node21455 : 4'b1010;
														assign node21455 = (inp[9]) ? 4'b1010 : 4'b1110;
													assign node21458 = (inp[2]) ? node21460 : 4'b1100;
														assign node21460 = (inp[10]) ? 4'b1000 : 4'b1010;
										assign node21463 = (inp[15]) ? node21485 : node21464;
											assign node21464 = (inp[3]) ? node21476 : node21465;
												assign node21465 = (inp[9]) ? node21471 : node21466;
													assign node21466 = (inp[4]) ? node21468 : 4'b1000;
														assign node21468 = (inp[10]) ? 4'b1110 : 4'b1000;
													assign node21471 = (inp[10]) ? node21473 : 4'b1110;
														assign node21473 = (inp[4]) ? 4'b1010 : 4'b1110;
												assign node21476 = (inp[10]) ? 4'b1010 : node21477;
													assign node21477 = (inp[9]) ? node21481 : node21478;
														assign node21478 = (inp[4]) ? 4'b1010 : 4'b1110;
														assign node21481 = (inp[4]) ? 4'b1010 : 4'b1010;
											assign node21485 = (inp[10]) ? node21497 : node21486;
												assign node21486 = (inp[3]) ? node21492 : node21487;
													assign node21487 = (inp[12]) ? 4'b1100 : node21488;
														assign node21488 = (inp[9]) ? 4'b1100 : 4'b1010;
													assign node21492 = (inp[2]) ? 4'b1100 : node21493;
														assign node21493 = (inp[12]) ? 4'b1000 : 4'b1100;
												assign node21497 = (inp[12]) ? node21503 : node21498;
													assign node21498 = (inp[4]) ? node21500 : 4'b1100;
														assign node21500 = (inp[9]) ? 4'b1000 : 4'b1100;
													assign node21503 = (inp[3]) ? node21507 : node21504;
														assign node21504 = (inp[9]) ? 4'b1000 : 4'b1100;
														assign node21507 = (inp[4]) ? 4'b1000 : 4'b1000;
								assign node21510 = (inp[14]) ? node21602 : node21511;
									assign node21511 = (inp[2]) ? node21559 : node21512;
										assign node21512 = (inp[15]) ? node21534 : node21513;
											assign node21513 = (inp[9]) ? node21523 : node21514;
												assign node21514 = (inp[10]) ? 4'b1000 : node21515;
													assign node21515 = (inp[3]) ? node21519 : node21516;
														assign node21516 = (inp[5]) ? 4'b1000 : 4'b1000;
														assign node21519 = (inp[4]) ? 4'b1110 : 4'b1000;
												assign node21523 = (inp[10]) ? node21531 : node21524;
													assign node21524 = (inp[12]) ? node21528 : node21525;
														assign node21525 = (inp[4]) ? 4'b1100 : 4'b1000;
														assign node21528 = (inp[4]) ? 4'b1010 : 4'b1110;
													assign node21531 = (inp[4]) ? 4'b1010 : 4'b1110;
											assign node21534 = (inp[5]) ? node21548 : node21535;
												assign node21535 = (inp[9]) ? node21541 : node21536;
													assign node21536 = (inp[12]) ? 4'b1110 : node21537;
														assign node21537 = (inp[4]) ? 4'b1010 : 4'b1010;
													assign node21541 = (inp[3]) ? node21545 : node21542;
														assign node21542 = (inp[4]) ? 4'b1110 : 4'b1010;
														assign node21545 = (inp[4]) ? 4'b1000 : 4'b1010;
												assign node21548 = (inp[9]) ? node21554 : node21549;
													assign node21549 = (inp[3]) ? node21551 : 4'b1010;
														assign node21551 = (inp[12]) ? 4'b1000 : 4'b1100;
													assign node21554 = (inp[4]) ? node21556 : 4'b1100;
														assign node21556 = (inp[10]) ? 4'b1000 : 4'b1100;
										assign node21559 = (inp[3]) ? node21583 : node21560;
											assign node21560 = (inp[15]) ? node21572 : node21561;
												assign node21561 = (inp[5]) ? node21567 : node21562;
													assign node21562 = (inp[10]) ? 4'b0001 : node21563;
														assign node21563 = (inp[4]) ? 4'b0101 : 4'b0001;
													assign node21567 = (inp[10]) ? 4'b0111 : node21568;
														assign node21568 = (inp[12]) ? 4'b0001 : 4'b0001;
												assign node21572 = (inp[5]) ? node21578 : node21573;
													assign node21573 = (inp[12]) ? node21575 : 4'b0111;
														assign node21575 = (inp[4]) ? 4'b0011 : 4'b0111;
													assign node21578 = (inp[4]) ? node21580 : 4'b0011;
														assign node21580 = (inp[12]) ? 4'b0101 : 4'b0001;
											assign node21583 = (inp[10]) ? node21595 : node21584;
												assign node21584 = (inp[5]) ? node21592 : node21585;
													assign node21585 = (inp[12]) ? node21589 : node21586;
														assign node21586 = (inp[15]) ? 4'b0011 : 4'b0001;
														assign node21589 = (inp[9]) ? 4'b0101 : 4'b0011;
													assign node21592 = (inp[15]) ? 4'b0001 : 4'b0011;
												assign node21595 = (inp[12]) ? 4'b0001 : node21596;
													assign node21596 = (inp[9]) ? node21598 : 4'b0101;
														assign node21598 = (inp[4]) ? 4'b0001 : 4'b0101;
									assign node21602 = (inp[3]) ? node21654 : node21603;
										assign node21603 = (inp[15]) ? node21629 : node21604;
											assign node21604 = (inp[5]) ? node21614 : node21605;
												assign node21605 = (inp[12]) ? node21607 : 4'b0101;
													assign node21607 = (inp[4]) ? node21611 : node21608;
														assign node21608 = (inp[9]) ? 4'b0101 : 4'b0001;
														assign node21611 = (inp[9]) ? 4'b0001 : 4'b0101;
												assign node21614 = (inp[9]) ? node21622 : node21615;
													assign node21615 = (inp[4]) ? node21619 : node21616;
														assign node21616 = (inp[10]) ? 4'b0001 : 4'b0101;
														assign node21619 = (inp[12]) ? 4'b0111 : 4'b0001;
													assign node21622 = (inp[4]) ? node21626 : node21623;
														assign node21623 = (inp[10]) ? 4'b0111 : 4'b0001;
														assign node21626 = (inp[12]) ? 4'b0011 : 4'b0011;
											assign node21629 = (inp[5]) ? node21641 : node21630;
												assign node21630 = (inp[12]) ? node21636 : node21631;
													assign node21631 = (inp[4]) ? node21633 : 4'b0111;
														assign node21633 = (inp[9]) ? 4'b0111 : 4'b0011;
													assign node21636 = (inp[10]) ? node21638 : 4'b0011;
														assign node21638 = (inp[2]) ? 4'b0111 : 4'b0011;
												assign node21641 = (inp[4]) ? node21649 : node21642;
													assign node21642 = (inp[10]) ? node21646 : node21643;
														assign node21643 = (inp[9]) ? 4'b0011 : 4'b0111;
														assign node21646 = (inp[9]) ? 4'b0101 : 4'b0011;
													assign node21649 = (inp[9]) ? node21651 : 4'b0101;
														assign node21651 = (inp[12]) ? 4'b0001 : 4'b0101;
										assign node21654 = (inp[15]) ? node21670 : node21655;
											assign node21655 = (inp[12]) ? node21663 : node21656;
												assign node21656 = (inp[2]) ? 4'b0001 : node21657;
													assign node21657 = (inp[9]) ? node21659 : 4'b0101;
														assign node21659 = (inp[4]) ? 4'b0011 : 4'b0011;
												assign node21663 = (inp[9]) ? node21667 : node21664;
													assign node21664 = (inp[4]) ? 4'b0111 : 4'b0011;
													assign node21667 = (inp[4]) ? 4'b0011 : 4'b0111;
											assign node21670 = (inp[5]) ? node21680 : node21671;
												assign node21671 = (inp[9]) ? node21677 : node21672;
													assign node21672 = (inp[2]) ? 4'b0011 : node21673;
														assign node21673 = (inp[12]) ? 4'b0011 : 4'b0111;
													assign node21677 = (inp[12]) ? 4'b0101 : 4'b0001;
												assign node21680 = (inp[12]) ? node21686 : node21681;
													assign node21681 = (inp[9]) ? 4'b0001 : node21682;
														assign node21682 = (inp[10]) ? 4'b0001 : 4'b0001;
													assign node21686 = (inp[10]) ? node21690 : node21687;
														assign node21687 = (inp[9]) ? 4'b0101 : 4'b0001;
														assign node21690 = (inp[4]) ? 4'b0001 : 4'b0001;
							assign node21693 = (inp[7]) ? node21857 : node21694;
								assign node21694 = (inp[14]) ? node21780 : node21695;
									assign node21695 = (inp[2]) ? node21737 : node21696;
										assign node21696 = (inp[15]) ? node21716 : node21697;
											assign node21697 = (inp[4]) ? node21707 : node21698;
												assign node21698 = (inp[3]) ? node21704 : node21699;
													assign node21699 = (inp[10]) ? node21701 : 4'b1000;
														assign node21701 = (inp[12]) ? 4'b1100 : 4'b1000;
													assign node21704 = (inp[12]) ? 4'b1010 : 4'b1000;
												assign node21707 = (inp[9]) ? node21713 : node21708;
													assign node21708 = (inp[5]) ? 4'b1110 : node21709;
														assign node21709 = (inp[12]) ? 4'b1100 : 4'b1000;
													assign node21713 = (inp[10]) ? 4'b1010 : 4'b1100;
											assign node21716 = (inp[5]) ? node21728 : node21717;
												assign node21717 = (inp[3]) ? node21723 : node21718;
													assign node21718 = (inp[10]) ? node21720 : 4'b1110;
														assign node21720 = (inp[9]) ? 4'b1010 : 4'b1110;
													assign node21723 = (inp[4]) ? 4'b1100 : node21724;
														assign node21724 = (inp[9]) ? 4'b1100 : 4'b1010;
												assign node21728 = (inp[9]) ? node21732 : node21729;
													assign node21729 = (inp[4]) ? 4'b1100 : 4'b1010;
													assign node21732 = (inp[4]) ? node21734 : 4'b1100;
														assign node21734 = (inp[12]) ? 4'b1000 : 4'b1100;
										assign node21737 = (inp[15]) ? node21759 : node21738;
											assign node21738 = (inp[5]) ? node21746 : node21739;
												assign node21739 = (inp[3]) ? 4'b0111 : node21740;
													assign node21740 = (inp[4]) ? node21742 : 4'b0001;
														assign node21742 = (inp[12]) ? 4'b0101 : 4'b0001;
												assign node21746 = (inp[4]) ? node21752 : node21747;
													assign node21747 = (inp[12]) ? 4'b0111 : node21748;
														assign node21748 = (inp[3]) ? 4'b0011 : 4'b0101;
													assign node21752 = (inp[9]) ? node21756 : node21753;
														assign node21753 = (inp[12]) ? 4'b0111 : 4'b0011;
														assign node21756 = (inp[12]) ? 4'b0011 : 4'b0011;
											assign node21759 = (inp[5]) ? node21771 : node21760;
												assign node21760 = (inp[3]) ? node21766 : node21761;
													assign node21761 = (inp[12]) ? node21763 : 4'b0011;
														assign node21763 = (inp[10]) ? 4'b0011 : 4'b0111;
													assign node21766 = (inp[12]) ? 4'b0101 : node21767;
														assign node21767 = (inp[4]) ? 4'b0101 : 4'b0011;
												assign node21771 = (inp[10]) ? 4'b0101 : node21772;
													assign node21772 = (inp[4]) ? node21776 : node21773;
														assign node21773 = (inp[12]) ? 4'b0001 : 4'b0011;
														assign node21776 = (inp[12]) ? 4'b0001 : 4'b0101;
									assign node21780 = (inp[15]) ? node21826 : node21781;
										assign node21781 = (inp[3]) ? node21807 : node21782;
											assign node21782 = (inp[5]) ? node21794 : node21783;
												assign node21783 = (inp[2]) ? node21789 : node21784;
													assign node21784 = (inp[9]) ? 4'b0101 : node21785;
														assign node21785 = (inp[4]) ? 4'b0001 : 4'b0001;
													assign node21789 = (inp[12]) ? node21791 : 4'b0001;
														assign node21791 = (inp[4]) ? 4'b0101 : 4'b0001;
												assign node21794 = (inp[9]) ? node21800 : node21795;
													assign node21795 = (inp[12]) ? node21797 : 4'b0001;
														assign node21797 = (inp[4]) ? 4'b0111 : 4'b0001;
													assign node21800 = (inp[4]) ? node21804 : node21801;
														assign node21801 = (inp[2]) ? 4'b0111 : 4'b0001;
														assign node21804 = (inp[12]) ? 4'b0011 : 4'b0011;
											assign node21807 = (inp[10]) ? node21817 : node21808;
												assign node21808 = (inp[9]) ? node21812 : node21809;
													assign node21809 = (inp[12]) ? 4'b0111 : 4'b0011;
													assign node21812 = (inp[2]) ? 4'b0111 : node21813;
														assign node21813 = (inp[4]) ? 4'b0011 : 4'b0111;
												assign node21817 = (inp[4]) ? node21823 : node21818;
													assign node21818 = (inp[9]) ? 4'b0111 : node21819;
														assign node21819 = (inp[5]) ? 4'b0011 : 4'b0001;
													assign node21823 = (inp[9]) ? 4'b0011 : 4'b0111;
										assign node21826 = (inp[3]) ? node21836 : node21827;
											assign node21827 = (inp[4]) ? 4'b0111 : node21828;
												assign node21828 = (inp[12]) ? 4'b0011 : node21829;
													assign node21829 = (inp[5]) ? node21831 : 4'b0111;
														assign node21831 = (inp[2]) ? 4'b0011 : 4'b0011;
											assign node21836 = (inp[5]) ? node21848 : node21837;
												assign node21837 = (inp[9]) ? node21843 : node21838;
													assign node21838 = (inp[4]) ? node21840 : 4'b0011;
														assign node21840 = (inp[10]) ? 4'b0101 : 4'b0001;
													assign node21843 = (inp[4]) ? node21845 : 4'b0101;
														assign node21845 = (inp[10]) ? 4'b0001 : 4'b0101;
												assign node21848 = (inp[12]) ? node21850 : 4'b0001;
													assign node21850 = (inp[9]) ? node21854 : node21851;
														assign node21851 = (inp[4]) ? 4'b0101 : 4'b0001;
														assign node21854 = (inp[4]) ? 4'b0001 : 4'b0101;
								assign node21857 = (inp[2]) ? node21947 : node21858;
									assign node21858 = (inp[14]) ? node21904 : node21859;
										assign node21859 = (inp[9]) ? node21883 : node21860;
											assign node21860 = (inp[4]) ? node21870 : node21861;
												assign node21861 = (inp[15]) ? node21863 : 4'b0001;
													assign node21863 = (inp[10]) ? node21867 : node21864;
														assign node21864 = (inp[5]) ? 4'b0001 : 4'b0111;
														assign node21867 = (inp[3]) ? 4'b0001 : 4'b0011;
												assign node21870 = (inp[12]) ? node21878 : node21871;
													assign node21871 = (inp[10]) ? node21875 : node21872;
														assign node21872 = (inp[5]) ? 4'b0001 : 4'b0011;
														assign node21875 = (inp[15]) ? 4'b0101 : 4'b0111;
													assign node21878 = (inp[15]) ? 4'b0101 : node21879;
														assign node21879 = (inp[3]) ? 4'b0111 : 4'b0101;
											assign node21883 = (inp[4]) ? node21895 : node21884;
												assign node21884 = (inp[5]) ? node21892 : node21885;
													assign node21885 = (inp[15]) ? node21889 : node21886;
														assign node21886 = (inp[3]) ? 4'b0001 : 4'b0101;
														assign node21889 = (inp[3]) ? 4'b0101 : 4'b0111;
													assign node21892 = (inp[15]) ? 4'b0101 : 4'b0111;
												assign node21895 = (inp[10]) ? node21901 : node21896;
													assign node21896 = (inp[12]) ? 4'b0011 : node21897;
														assign node21897 = (inp[3]) ? 4'b0101 : 4'b0101;
													assign node21901 = (inp[15]) ? 4'b0001 : 4'b0011;
										assign node21904 = (inp[15]) ? node21922 : node21905;
											assign node21905 = (inp[5]) ? node21913 : node21906;
												assign node21906 = (inp[3]) ? node21908 : 4'b0100;
													assign node21908 = (inp[4]) ? node21910 : 4'b0000;
														assign node21910 = (inp[12]) ? 4'b0110 : 4'b0010;
												assign node21913 = (inp[9]) ? node21917 : node21914;
													assign node21914 = (inp[3]) ? 4'b0010 : 4'b0000;
													assign node21917 = (inp[4]) ? node21919 : 4'b0110;
														assign node21919 = (inp[10]) ? 4'b0010 : 4'b0010;
											assign node21922 = (inp[5]) ? node21936 : node21923;
												assign node21923 = (inp[3]) ? node21929 : node21924;
													assign node21924 = (inp[10]) ? 4'b0010 : node21925;
														assign node21925 = (inp[4]) ? 4'b0110 : 4'b0010;
													assign node21929 = (inp[4]) ? node21933 : node21930;
														assign node21930 = (inp[10]) ? 4'b0100 : 4'b0010;
														assign node21933 = (inp[9]) ? 4'b0000 : 4'b0100;
												assign node21936 = (inp[12]) ? node21940 : node21937;
													assign node21937 = (inp[3]) ? 4'b0000 : 4'b0100;
													assign node21940 = (inp[9]) ? node21944 : node21941;
														assign node21941 = (inp[4]) ? 4'b0100 : 4'b0010;
														assign node21944 = (inp[4]) ? 4'b0000 : 4'b0100;
									assign node21947 = (inp[9]) ? node21985 : node21948;
										assign node21948 = (inp[4]) ? node21968 : node21949;
											assign node21949 = (inp[10]) ? node21961 : node21950;
												assign node21950 = (inp[12]) ? node21956 : node21951;
													assign node21951 = (inp[15]) ? 4'b0110 : node21952;
														assign node21952 = (inp[5]) ? 4'b0100 : 4'b0100;
													assign node21956 = (inp[5]) ? 4'b0000 : node21957;
														assign node21957 = (inp[15]) ? 4'b0010 : 4'b0000;
												assign node21961 = (inp[15]) ? 4'b0010 : node21962;
													assign node21962 = (inp[3]) ? node21964 : 4'b0000;
														assign node21964 = (inp[5]) ? 4'b0010 : 4'b0000;
											assign node21968 = (inp[10]) ? node21978 : node21969;
												assign node21969 = (inp[12]) ? node21973 : node21970;
													assign node21970 = (inp[5]) ? 4'b0000 : 4'b0010;
													assign node21973 = (inp[15]) ? node21975 : 4'b0110;
														assign node21975 = (inp[5]) ? 4'b0100 : 4'b0100;
												assign node21978 = (inp[14]) ? 4'b0100 : node21979;
													assign node21979 = (inp[3]) ? 4'b0110 : node21980;
														assign node21980 = (inp[12]) ? 4'b0100 : 4'b0110;
										assign node21985 = (inp[12]) ? node22007 : node21986;
											assign node21986 = (inp[15]) ? node21996 : node21987;
												assign node21987 = (inp[4]) ? node21993 : node21988;
													assign node21988 = (inp[10]) ? 4'b0110 : node21989;
														assign node21989 = (inp[5]) ? 4'b0000 : 4'b0000;
													assign node21993 = (inp[10]) ? 4'b0010 : 4'b0110;
												assign node21996 = (inp[3]) ? node22004 : node21997;
													assign node21997 = (inp[5]) ? node22001 : node21998;
														assign node21998 = (inp[14]) ? 4'b0110 : 4'b0010;
														assign node22001 = (inp[4]) ? 4'b0100 : 4'b0010;
													assign node22004 = (inp[10]) ? 4'b0000 : 4'b0100;
											assign node22007 = (inp[4]) ? node22017 : node22008;
												assign node22008 = (inp[3]) ? node22014 : node22009;
													assign node22009 = (inp[5]) ? 4'b0100 : node22010;
														assign node22010 = (inp[15]) ? 4'b0110 : 4'b0100;
													assign node22014 = (inp[15]) ? 4'b0100 : 4'b0110;
												assign node22017 = (inp[15]) ? node22019 : 4'b0010;
													assign node22019 = (inp[3]) ? 4'b0000 : 4'b0010;
						assign node22022 = (inp[15]) ? node22386 : node22023;
							assign node22023 = (inp[5]) ? node22183 : node22024;
								assign node22024 = (inp[3]) ? node22100 : node22025;
									assign node22025 = (inp[9]) ? node22067 : node22026;
										assign node22026 = (inp[4]) ? node22048 : node22027;
											assign node22027 = (inp[12]) ? node22037 : node22028;
												assign node22028 = (inp[10]) ? 4'b0000 : node22029;
													assign node22029 = (inp[14]) ? node22033 : node22030;
														assign node22030 = (inp[2]) ? 4'b0100 : 4'b0100;
														assign node22033 = (inp[8]) ? 4'b0100 : 4'b0100;
												assign node22037 = (inp[7]) ? node22043 : node22038;
													assign node22038 = (inp[8]) ? node22040 : 4'b0000;
														assign node22040 = (inp[2]) ? 4'b0001 : 4'b0000;
													assign node22043 = (inp[8]) ? node22045 : 4'b0001;
														assign node22045 = (inp[2]) ? 4'b0000 : 4'b0001;
											assign node22048 = (inp[10]) ? node22058 : node22049;
												assign node22049 = (inp[12]) ? node22053 : node22050;
													assign node22050 = (inp[2]) ? 4'b0000 : 4'b0001;
													assign node22053 = (inp[8]) ? node22055 : 4'b0100;
														assign node22055 = (inp[7]) ? 4'b0100 : 4'b0101;
												assign node22058 = (inp[8]) ? node22062 : node22059;
													assign node22059 = (inp[7]) ? 4'b0101 : 4'b0100;
													assign node22062 = (inp[7]) ? 4'b0100 : node22063;
														assign node22063 = (inp[14]) ? 4'b0101 : 4'b0100;
										assign node22067 = (inp[4]) ? node22083 : node22068;
											assign node22068 = (inp[10]) ? node22076 : node22069;
												assign node22069 = (inp[12]) ? 4'b0100 : node22070;
													assign node22070 = (inp[2]) ? 4'b0000 : node22071;
														assign node22071 = (inp[7]) ? 4'b0000 : 4'b0000;
												assign node22076 = (inp[2]) ? node22078 : 4'b0100;
													assign node22078 = (inp[8]) ? node22080 : 4'b0101;
														assign node22080 = (inp[7]) ? 4'b0100 : 4'b0101;
											assign node22083 = (inp[7]) ? node22091 : node22084;
												assign node22084 = (inp[12]) ? 4'b0001 : node22085;
													assign node22085 = (inp[8]) ? node22087 : 4'b0000;
														assign node22087 = (inp[14]) ? 4'b0001 : 4'b0000;
												assign node22091 = (inp[10]) ? node22095 : node22092;
													assign node22092 = (inp[12]) ? 4'b0000 : 4'b0100;
													assign node22095 = (inp[8]) ? 4'b0000 : node22096;
														assign node22096 = (inp[2]) ? 4'b0001 : 4'b0000;
									assign node22100 = (inp[9]) ? node22146 : node22101;
										assign node22101 = (inp[4]) ? node22125 : node22102;
											assign node22102 = (inp[10]) ? node22116 : node22103;
												assign node22103 = (inp[12]) ? node22111 : node22104;
													assign node22104 = (inp[8]) ? node22108 : node22105;
														assign node22105 = (inp[2]) ? 4'b0100 : 4'b0101;
														assign node22108 = (inp[7]) ? 4'b0100 : 4'b0101;
													assign node22111 = (inp[8]) ? node22113 : 4'b0000;
														assign node22113 = (inp[7]) ? 4'b0000 : 4'b0001;
												assign node22116 = (inp[2]) ? node22118 : 4'b0000;
													assign node22118 = (inp[8]) ? node22122 : node22119;
														assign node22119 = (inp[7]) ? 4'b0001 : 4'b0000;
														assign node22122 = (inp[7]) ? 4'b0000 : 4'b0001;
											assign node22125 = (inp[12]) ? node22135 : node22126;
												assign node22126 = (inp[10]) ? node22130 : node22127;
													assign node22127 = (inp[8]) ? 4'b0001 : 4'b0000;
													assign node22130 = (inp[14]) ? 4'b0111 : node22131;
														assign node22131 = (inp[7]) ? 4'b0111 : 4'b0110;
												assign node22135 = (inp[2]) ? node22141 : node22136;
													assign node22136 = (inp[10]) ? node22138 : 4'b0110;
														assign node22138 = (inp[7]) ? 4'b0111 : 4'b0110;
													assign node22141 = (inp[7]) ? 4'b0111 : node22142;
														assign node22142 = (inp[8]) ? 4'b0111 : 4'b0110;
										assign node22146 = (inp[4]) ? node22166 : node22147;
											assign node22147 = (inp[10]) ? node22155 : node22148;
												assign node22148 = (inp[12]) ? node22152 : node22149;
													assign node22149 = (inp[14]) ? 4'b0001 : 4'b0000;
													assign node22152 = (inp[2]) ? 4'b0111 : 4'b0110;
												assign node22155 = (inp[12]) ? node22161 : node22156;
													assign node22156 = (inp[8]) ? node22158 : 4'b0111;
														assign node22158 = (inp[14]) ? 4'b0110 : 4'b0110;
													assign node22161 = (inp[7]) ? node22163 : 4'b0110;
														assign node22163 = (inp[14]) ? 4'b0111 : 4'b0110;
											assign node22166 = (inp[10]) ? node22174 : node22167;
												assign node22167 = (inp[12]) ? 4'b0011 : node22168;
													assign node22168 = (inp[14]) ? node22170 : 4'b0110;
														assign node22170 = (inp[2]) ? 4'b0110 : 4'b0110;
												assign node22174 = (inp[2]) ? node22180 : node22175;
													assign node22175 = (inp[7]) ? 4'b0011 : node22176;
														assign node22176 = (inp[14]) ? 4'b0010 : 4'b0010;
													assign node22180 = (inp[12]) ? 4'b0010 : 4'b0011;
								assign node22183 = (inp[3]) ? node22273 : node22184;
									assign node22184 = (inp[4]) ? node22232 : node22185;
										assign node22185 = (inp[9]) ? node22211 : node22186;
											assign node22186 = (inp[10]) ? node22198 : node22187;
												assign node22187 = (inp[12]) ? node22193 : node22188;
													assign node22188 = (inp[2]) ? node22190 : 4'b0100;
														assign node22190 = (inp[7]) ? 4'b0101 : 4'b0100;
													assign node22193 = (inp[8]) ? 4'b0000 : node22194;
														assign node22194 = (inp[7]) ? 4'b0000 : 4'b0000;
												assign node22198 = (inp[14]) ? node22204 : node22199;
													assign node22199 = (inp[8]) ? node22201 : 4'b0001;
														assign node22201 = (inp[7]) ? 4'b0001 : 4'b0000;
													assign node22204 = (inp[7]) ? node22208 : node22205;
														assign node22205 = (inp[8]) ? 4'b0001 : 4'b0000;
														assign node22208 = (inp[8]) ? 4'b0000 : 4'b0001;
											assign node22211 = (inp[12]) ? node22223 : node22212;
												assign node22212 = (inp[10]) ? node22218 : node22213;
													assign node22213 = (inp[7]) ? 4'b0000 : node22214;
														assign node22214 = (inp[8]) ? 4'b0001 : 4'b0000;
													assign node22218 = (inp[8]) ? node22220 : 4'b0110;
														assign node22220 = (inp[14]) ? 4'b0111 : 4'b0110;
												assign node22223 = (inp[8]) ? 4'b0110 : node22224;
													assign node22224 = (inp[10]) ? node22228 : node22225;
														assign node22225 = (inp[14]) ? 4'b0111 : 4'b0111;
														assign node22228 = (inp[2]) ? 4'b0110 : 4'b0111;
										assign node22232 = (inp[9]) ? node22248 : node22233;
											assign node22233 = (inp[7]) ? node22243 : node22234;
												assign node22234 = (inp[10]) ? node22236 : 4'b0110;
													assign node22236 = (inp[12]) ? node22240 : node22237;
														assign node22237 = (inp[8]) ? 4'b0111 : 4'b0110;
														assign node22240 = (inp[2]) ? 4'b0111 : 4'b0110;
												assign node22243 = (inp[10]) ? 4'b0110 : node22244;
													assign node22244 = (inp[12]) ? 4'b0111 : 4'b0000;
											assign node22248 = (inp[12]) ? node22260 : node22249;
												assign node22249 = (inp[10]) ? node22255 : node22250;
													assign node22250 = (inp[8]) ? node22252 : 4'b0110;
														assign node22252 = (inp[7]) ? 4'b0110 : 4'b0111;
													assign node22255 = (inp[8]) ? node22257 : 4'b0011;
														assign node22257 = (inp[7]) ? 4'b0010 : 4'b0011;
												assign node22260 = (inp[10]) ? node22266 : node22261;
													assign node22261 = (inp[7]) ? 4'b0010 : node22262;
														assign node22262 = (inp[2]) ? 4'b0010 : 4'b0010;
													assign node22266 = (inp[2]) ? node22270 : node22267;
														assign node22267 = (inp[14]) ? 4'b0010 : 4'b0011;
														assign node22270 = (inp[7]) ? 4'b0011 : 4'b0010;
									assign node22273 = (inp[14]) ? node22327 : node22274;
										assign node22274 = (inp[12]) ? node22302 : node22275;
											assign node22275 = (inp[4]) ? node22291 : node22276;
												assign node22276 = (inp[7]) ? node22284 : node22277;
													assign node22277 = (inp[2]) ? node22281 : node22278;
														assign node22278 = (inp[8]) ? 4'b0010 : 4'b0011;
														assign node22281 = (inp[8]) ? 4'b0111 : 4'b0010;
													assign node22284 = (inp[2]) ? node22288 : node22285;
														assign node22285 = (inp[10]) ? 4'b0110 : 4'b0111;
														assign node22288 = (inp[8]) ? 4'b0010 : 4'b0011;
												assign node22291 = (inp[9]) ? node22297 : node22292;
													assign node22292 = (inp[10]) ? node22294 : 4'b0011;
														assign node22294 = (inp[7]) ? 4'b0111 : 4'b0110;
													assign node22297 = (inp[10]) ? 4'b0010 : node22298;
														assign node22298 = (inp[7]) ? 4'b0110 : 4'b0111;
											assign node22302 = (inp[8]) ? node22316 : node22303;
												assign node22303 = (inp[7]) ? node22309 : node22304;
													assign node22304 = (inp[2]) ? 4'b0110 : node22305;
														assign node22305 = (inp[10]) ? 4'b0111 : 4'b0011;
													assign node22309 = (inp[9]) ? node22313 : node22310;
														assign node22310 = (inp[4]) ? 4'b0111 : 4'b0011;
														assign node22313 = (inp[4]) ? 4'b0011 : 4'b0111;
												assign node22316 = (inp[10]) ? node22320 : node22317;
													assign node22317 = (inp[7]) ? 4'b0111 : 4'b0010;
													assign node22320 = (inp[7]) ? node22324 : node22321;
														assign node22321 = (inp[9]) ? 4'b0111 : 4'b0011;
														assign node22324 = (inp[2]) ? 4'b0010 : 4'b0011;
										assign node22327 = (inp[10]) ? node22357 : node22328;
											assign node22328 = (inp[4]) ? node22342 : node22329;
												assign node22329 = (inp[2]) ? node22337 : node22330;
													assign node22330 = (inp[12]) ? node22334 : node22331;
														assign node22331 = (inp[8]) ? 4'b0110 : 4'b0011;
														assign node22334 = (inp[9]) ? 4'b0111 : 4'b0010;
													assign node22337 = (inp[9]) ? 4'b0011 : node22338;
														assign node22338 = (inp[12]) ? 4'b0011 : 4'b0111;
												assign node22342 = (inp[7]) ? node22350 : node22343;
													assign node22343 = (inp[8]) ? node22347 : node22344;
														assign node22344 = (inp[2]) ? 4'b0010 : 4'b0110;
														assign node22347 = (inp[2]) ? 4'b0011 : 4'b0111;
													assign node22350 = (inp[8]) ? node22354 : node22351;
														assign node22351 = (inp[12]) ? 4'b0011 : 4'b0111;
														assign node22354 = (inp[12]) ? 4'b0010 : 4'b0110;
											assign node22357 = (inp[2]) ? node22373 : node22358;
												assign node22358 = (inp[12]) ? node22366 : node22359;
													assign node22359 = (inp[4]) ? node22363 : node22360;
														assign node22360 = (inp[8]) ? 4'b0010 : 4'b0010;
														assign node22363 = (inp[9]) ? 4'b0011 : 4'b0111;
													assign node22366 = (inp[9]) ? node22370 : node22367;
														assign node22367 = (inp[4]) ? 4'b0111 : 4'b0011;
														assign node22370 = (inp[4]) ? 4'b0010 : 4'b0111;
												assign node22373 = (inp[12]) ? node22379 : node22374;
													assign node22374 = (inp[8]) ? 4'b0110 : node22375;
														assign node22375 = (inp[7]) ? 4'b0011 : 4'b0010;
													assign node22379 = (inp[4]) ? node22383 : node22380;
														assign node22380 = (inp[8]) ? 4'b0110 : 4'b0110;
														assign node22383 = (inp[9]) ? 4'b0011 : 4'b0111;
							assign node22386 = (inp[5]) ? node22584 : node22387;
								assign node22387 = (inp[3]) ? node22489 : node22388;
									assign node22388 = (inp[9]) ? node22434 : node22389;
										assign node22389 = (inp[4]) ? node22411 : node22390;
											assign node22390 = (inp[12]) ? node22400 : node22391;
												assign node22391 = (inp[10]) ? node22395 : node22392;
													assign node22392 = (inp[14]) ? 4'b0111 : 4'b0110;
													assign node22395 = (inp[14]) ? 4'b0010 : node22396;
														assign node22396 = (inp[7]) ? 4'b0010 : 4'b0010;
												assign node22400 = (inp[14]) ? node22406 : node22401;
													assign node22401 = (inp[10]) ? node22403 : 4'b0010;
														assign node22403 = (inp[7]) ? 4'b0010 : 4'b0010;
													assign node22406 = (inp[10]) ? 4'b0010 : node22407;
														assign node22407 = (inp[8]) ? 4'b0010 : 4'b0010;
											assign node22411 = (inp[2]) ? node22421 : node22412;
												assign node22412 = (inp[8]) ? 4'b0110 : node22413;
													assign node22413 = (inp[12]) ? node22417 : node22414;
														assign node22414 = (inp[7]) ? 4'b0111 : 4'b0110;
														assign node22417 = (inp[7]) ? 4'b0110 : 4'b0111;
												assign node22421 = (inp[10]) ? node22429 : node22422;
													assign node22422 = (inp[12]) ? node22426 : node22423;
														assign node22423 = (inp[7]) ? 4'b0011 : 4'b0010;
														assign node22426 = (inp[7]) ? 4'b0110 : 4'b0110;
													assign node22429 = (inp[8]) ? 4'b0111 : node22430;
														assign node22430 = (inp[7]) ? 4'b0111 : 4'b0110;
										assign node22434 = (inp[4]) ? node22460 : node22435;
											assign node22435 = (inp[10]) ? node22449 : node22436;
												assign node22436 = (inp[12]) ? node22442 : node22437;
													assign node22437 = (inp[14]) ? 4'b0011 : node22438;
														assign node22438 = (inp[2]) ? 4'b0010 : 4'b0011;
													assign node22442 = (inp[2]) ? node22446 : node22443;
														assign node22443 = (inp[14]) ? 4'b0110 : 4'b0111;
														assign node22446 = (inp[7]) ? 4'b0110 : 4'b0110;
												assign node22449 = (inp[12]) ? node22455 : node22450;
													assign node22450 = (inp[8]) ? 4'b0110 : node22451;
														assign node22451 = (inp[7]) ? 4'b0111 : 4'b0110;
													assign node22455 = (inp[7]) ? 4'b0110 : node22456;
														assign node22456 = (inp[8]) ? 4'b0111 : 4'b0110;
											assign node22460 = (inp[12]) ? node22474 : node22461;
												assign node22461 = (inp[10]) ? node22467 : node22462;
													assign node22462 = (inp[2]) ? 4'b0111 : node22463;
														assign node22463 = (inp[8]) ? 4'b0110 : 4'b0111;
													assign node22467 = (inp[8]) ? node22471 : node22468;
														assign node22468 = (inp[14]) ? 4'b0010 : 4'b0010;
														assign node22471 = (inp[7]) ? 4'b0010 : 4'b0011;
												assign node22474 = (inp[14]) ? node22482 : node22475;
													assign node22475 = (inp[10]) ? node22479 : node22476;
														assign node22476 = (inp[8]) ? 4'b0011 : 4'b0010;
														assign node22479 = (inp[8]) ? 4'b0010 : 4'b0010;
													assign node22482 = (inp[8]) ? node22486 : node22483;
														assign node22483 = (inp[7]) ? 4'b0011 : 4'b0010;
														assign node22486 = (inp[7]) ? 4'b0010 : 4'b0011;
									assign node22489 = (inp[4]) ? node22537 : node22490;
										assign node22490 = (inp[9]) ? node22510 : node22491;
											assign node22491 = (inp[10]) ? node22501 : node22492;
												assign node22492 = (inp[12]) ? node22498 : node22493;
													assign node22493 = (inp[14]) ? node22495 : 4'b0111;
														assign node22495 = (inp[7]) ? 4'b0111 : 4'b0110;
													assign node22498 = (inp[2]) ? 4'b0011 : 4'b0010;
												assign node22501 = (inp[8]) ? node22503 : 4'b0011;
													assign node22503 = (inp[14]) ? node22507 : node22504;
														assign node22504 = (inp[12]) ? 4'b0010 : 4'b0010;
														assign node22507 = (inp[7]) ? 4'b0010 : 4'b0011;
											assign node22510 = (inp[10]) ? node22524 : node22511;
												assign node22511 = (inp[12]) ? node22519 : node22512;
													assign node22512 = (inp[7]) ? node22516 : node22513;
														assign node22513 = (inp[8]) ? 4'b0011 : 4'b0010;
														assign node22516 = (inp[8]) ? 4'b0010 : 4'b0011;
													assign node22519 = (inp[8]) ? node22521 : 4'b0100;
														assign node22521 = (inp[2]) ? 4'b0100 : 4'b0100;
												assign node22524 = (inp[7]) ? node22530 : node22525;
													assign node22525 = (inp[2]) ? 4'b0101 : node22526;
														assign node22526 = (inp[8]) ? 4'b0100 : 4'b0101;
													assign node22530 = (inp[12]) ? node22534 : node22531;
														assign node22531 = (inp[2]) ? 4'b0100 : 4'b0100;
														assign node22534 = (inp[14]) ? 4'b0101 : 4'b0100;
										assign node22537 = (inp[9]) ? node22563 : node22538;
											assign node22538 = (inp[12]) ? node22550 : node22539;
												assign node22539 = (inp[10]) ? node22545 : node22540;
													assign node22540 = (inp[7]) ? node22542 : 4'b0010;
														assign node22542 = (inp[8]) ? 4'b0010 : 4'b0011;
													assign node22545 = (inp[14]) ? 4'b0100 : node22546;
														assign node22546 = (inp[2]) ? 4'b0101 : 4'b0100;
												assign node22550 = (inp[8]) ? node22556 : node22551;
													assign node22551 = (inp[10]) ? node22553 : 4'b0100;
														assign node22553 = (inp[2]) ? 4'b0100 : 4'b0100;
													assign node22556 = (inp[14]) ? node22560 : node22557;
														assign node22557 = (inp[2]) ? 4'b0100 : 4'b0100;
														assign node22560 = (inp[7]) ? 4'b0100 : 4'b0101;
											assign node22563 = (inp[10]) ? node22577 : node22564;
												assign node22564 = (inp[12]) ? node22572 : node22565;
													assign node22565 = (inp[7]) ? node22569 : node22566;
														assign node22566 = (inp[14]) ? 4'b0100 : 4'b0100;
														assign node22569 = (inp[14]) ? 4'b0100 : 4'b0101;
													assign node22572 = (inp[2]) ? node22574 : 4'b0000;
														assign node22574 = (inp[7]) ? 4'b0001 : 4'b0000;
												assign node22577 = (inp[7]) ? 4'b0000 : node22578;
													assign node22578 = (inp[8]) ? node22580 : 4'b0000;
														assign node22580 = (inp[12]) ? 4'b0001 : 4'b0001;
								assign node22584 = (inp[3]) ? node22668 : node22585;
									assign node22585 = (inp[4]) ? node22627 : node22586;
										assign node22586 = (inp[9]) ? node22606 : node22587;
											assign node22587 = (inp[10]) ? node22599 : node22588;
												assign node22588 = (inp[12]) ? node22594 : node22589;
													assign node22589 = (inp[2]) ? node22591 : 4'b0111;
														assign node22591 = (inp[8]) ? 4'b0110 : 4'b0110;
													assign node22594 = (inp[14]) ? 4'b0011 : node22595;
														assign node22595 = (inp[8]) ? 4'b0011 : 4'b0010;
												assign node22599 = (inp[12]) ? 4'b0010 : node22600;
													assign node22600 = (inp[14]) ? node22602 : 4'b0010;
														assign node22602 = (inp[8]) ? 4'b0010 : 4'b0011;
											assign node22606 = (inp[10]) ? node22614 : node22607;
												assign node22607 = (inp[12]) ? node22609 : 4'b0010;
													assign node22609 = (inp[14]) ? 4'b0100 : node22610;
														assign node22610 = (inp[8]) ? 4'b0100 : 4'b0101;
												assign node22614 = (inp[12]) ? node22622 : node22615;
													assign node22615 = (inp[2]) ? node22619 : node22616;
														assign node22616 = (inp[14]) ? 4'b0100 : 4'b0101;
														assign node22619 = (inp[8]) ? 4'b0100 : 4'b0100;
													assign node22622 = (inp[7]) ? 4'b0101 : node22623;
														assign node22623 = (inp[2]) ? 4'b0101 : 4'b0100;
										assign node22627 = (inp[9]) ? node22641 : node22628;
											assign node22628 = (inp[10]) ? node22632 : node22629;
												assign node22629 = (inp[12]) ? 4'b0101 : 4'b0011;
												assign node22632 = (inp[12]) ? node22634 : 4'b0101;
													assign node22634 = (inp[7]) ? node22638 : node22635;
														assign node22635 = (inp[8]) ? 4'b0101 : 4'b0100;
														assign node22638 = (inp[2]) ? 4'b0100 : 4'b0100;
											assign node22641 = (inp[10]) ? node22655 : node22642;
												assign node22642 = (inp[12]) ? node22650 : node22643;
													assign node22643 = (inp[2]) ? node22647 : node22644;
														assign node22644 = (inp[7]) ? 4'b0101 : 4'b0100;
														assign node22647 = (inp[14]) ? 4'b0100 : 4'b0100;
													assign node22650 = (inp[8]) ? 4'b0001 : node22651;
														assign node22651 = (inp[7]) ? 4'b0001 : 4'b0000;
												assign node22655 = (inp[12]) ? node22661 : node22656;
													assign node22656 = (inp[7]) ? 4'b0001 : node22657;
														assign node22657 = (inp[8]) ? 4'b0001 : 4'b0000;
													assign node22661 = (inp[8]) ? node22665 : node22662;
														assign node22662 = (inp[2]) ? 4'b0001 : 4'b0000;
														assign node22665 = (inp[2]) ? 4'b0000 : 4'b0000;
									assign node22668 = (inp[10]) ? node22722 : node22669;
										assign node22669 = (inp[4]) ? node22699 : node22670;
											assign node22670 = (inp[7]) ? node22686 : node22671;
												assign node22671 = (inp[8]) ? node22679 : node22672;
													assign node22672 = (inp[9]) ? node22676 : node22673;
														assign node22673 = (inp[12]) ? 4'b0000 : 4'b0100;
														assign node22676 = (inp[12]) ? 4'b0100 : 4'b0000;
													assign node22679 = (inp[14]) ? node22683 : node22680;
														assign node22680 = (inp[12]) ? 4'b0000 : 4'b0100;
														assign node22683 = (inp[12]) ? 4'b0101 : 4'b0001;
												assign node22686 = (inp[8]) ? node22692 : node22687;
													assign node22687 = (inp[2]) ? node22689 : 4'b0000;
														assign node22689 = (inp[12]) ? 4'b0001 : 4'b0001;
													assign node22692 = (inp[2]) ? node22696 : node22693;
														assign node22693 = (inp[14]) ? 4'b0000 : 4'b0001;
														assign node22696 = (inp[12]) ? 4'b0000 : 4'b0000;
											assign node22699 = (inp[14]) ? node22711 : node22700;
												assign node22700 = (inp[9]) ? node22706 : node22701;
													assign node22701 = (inp[12]) ? node22703 : 4'b0001;
														assign node22703 = (inp[2]) ? 4'b0101 : 4'b0100;
													assign node22706 = (inp[7]) ? 4'b0100 : node22707;
														assign node22707 = (inp[2]) ? 4'b0100 : 4'b0100;
												assign node22711 = (inp[7]) ? node22717 : node22712;
													assign node22712 = (inp[8]) ? node22714 : 4'b0100;
														assign node22714 = (inp[9]) ? 4'b0101 : 4'b0001;
													assign node22717 = (inp[8]) ? node22719 : 4'b0001;
														assign node22719 = (inp[2]) ? 4'b0000 : 4'b0000;
										assign node22722 = (inp[7]) ? node22750 : node22723;
											assign node22723 = (inp[12]) ? node22737 : node22724;
												assign node22724 = (inp[8]) ? node22730 : node22725;
													assign node22725 = (inp[2]) ? 4'b0100 : node22726;
														assign node22726 = (inp[14]) ? 4'b0100 : 4'b0001;
													assign node22730 = (inp[14]) ? node22734 : node22731;
														assign node22731 = (inp[4]) ? 4'b0101 : 4'b0000;
														assign node22734 = (inp[2]) ? 4'b0001 : 4'b0101;
												assign node22737 = (inp[14]) ? node22745 : node22738;
													assign node22738 = (inp[8]) ? node22742 : node22739;
														assign node22739 = (inp[2]) ? 4'b0000 : 4'b0101;
														assign node22742 = (inp[9]) ? 4'b0100 : 4'b0000;
													assign node22745 = (inp[4]) ? node22747 : 4'b0000;
														assign node22747 = (inp[9]) ? 4'b0000 : 4'b0100;
											assign node22750 = (inp[8]) ? node22760 : node22751;
												assign node22751 = (inp[9]) ? node22757 : node22752;
													assign node22752 = (inp[4]) ? 4'b0101 : node22753;
														assign node22753 = (inp[2]) ? 4'b0001 : 4'b0000;
													assign node22757 = (inp[4]) ? 4'b0001 : 4'b0101;
												assign node22760 = (inp[14]) ? node22766 : node22761;
													assign node22761 = (inp[9]) ? 4'b0101 : node22762;
														assign node22762 = (inp[4]) ? 4'b0101 : 4'b0001;
													assign node22766 = (inp[12]) ? node22770 : node22767;
														assign node22767 = (inp[4]) ? 4'b0100 : 4'b0000;
														assign node22770 = (inp[4]) ? 4'b0000 : 4'b0100;

endmodule