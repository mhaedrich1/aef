module dtc_split66_bm60 (
	input  wire [12-1:0] inp,
	output wire [3-1:0] outp
);

	wire [3-1:0] node1;
	wire [3-1:0] node2;
	wire [3-1:0] node3;
	wire [3-1:0] node4;
	wire [3-1:0] node6;
	wire [3-1:0] node8;
	wire [3-1:0] node10;
	wire [3-1:0] node13;
	wire [3-1:0] node14;
	wire [3-1:0] node16;
	wire [3-1:0] node18;
	wire [3-1:0] node20;
	wire [3-1:0] node22;
	wire [3-1:0] node26;
	wire [3-1:0] node27;
	wire [3-1:0] node29;
	wire [3-1:0] node31;
	wire [3-1:0] node33;
	wire [3-1:0] node36;
	wire [3-1:0] node37;
	wire [3-1:0] node38;
	wire [3-1:0] node39;
	wire [3-1:0] node41;
	wire [3-1:0] node43;
	wire [3-1:0] node48;
	wire [3-1:0] node51;
	wire [3-1:0] node52;
	wire [3-1:0] node53;
	wire [3-1:0] node55;
	wire [3-1:0] node57;
	wire [3-1:0] node58;
	wire [3-1:0] node60;
	wire [3-1:0] node62;
	wire [3-1:0] node66;
	wire [3-1:0] node68;
	wire [3-1:0] node71;
	wire [3-1:0] node72;
	wire [3-1:0] node74;
	wire [3-1:0] node75;
	wire [3-1:0] node76;
	wire [3-1:0] node78;
	wire [3-1:0] node80;
	wire [3-1:0] node84;
	wire [3-1:0] node86;
	wire [3-1:0] node88;
	wire [3-1:0] node90;
	wire [3-1:0] node93;
	wire [3-1:0] node95;
	wire [3-1:0] node97;
	wire [3-1:0] node98;
	wire [3-1:0] node102;
	wire [3-1:0] node103;
	wire [3-1:0] node104;
	wire [3-1:0] node105;
	wire [3-1:0] node107;
	wire [3-1:0] node108;
	wire [3-1:0] node110;
	wire [3-1:0] node112;
	wire [3-1:0] node114;
	wire [3-1:0] node118;
	wire [3-1:0] node119;
	wire [3-1:0] node120;
	wire [3-1:0] node121;
	wire [3-1:0] node123;
	wire [3-1:0] node124;
	wire [3-1:0] node126;
	wire [3-1:0] node133;
	wire [3-1:0] node134;
	wire [3-1:0] node135;
	wire [3-1:0] node137;
	wire [3-1:0] node139;
	wire [3-1:0] node143;
	wire [3-1:0] node145;
	wire [3-1:0] node146;
	wire [3-1:0] node148;
	wire [3-1:0] node150;
	wire [3-1:0] node152;
	wire [3-1:0] node156;
	wire [3-1:0] node157;
	wire [3-1:0] node158;
	wire [3-1:0] node160;
	wire [3-1:0] node161;
	wire [3-1:0] node163;
	wire [3-1:0] node165;
	wire [3-1:0] node167;
	wire [3-1:0] node170;
	wire [3-1:0] node171;
	wire [3-1:0] node173;
	wire [3-1:0] node175;
	wire [3-1:0] node179;
	wire [3-1:0] node181;
	wire [3-1:0] node182;
	wire [3-1:0] node184;
	wire [3-1:0] node188;
	wire [3-1:0] node189;
	wire [3-1:0] node190;
	wire [3-1:0] node191;
	wire [3-1:0] node192;
	wire [3-1:0] node194;
	wire [3-1:0] node196;
	wire [3-1:0] node200;
	wire [3-1:0] node202;
	wire [3-1:0] node204;
	wire [3-1:0] node206;
	wire [3-1:0] node209;
	wire [3-1:0] node211;
	wire [3-1:0] node213;
	wire [3-1:0] node216;
	wire [3-1:0] node217;
	wire [3-1:0] node218;
	wire [3-1:0] node220;
	wire [3-1:0] node222;
	wire [3-1:0] node224;
	wire [3-1:0] node227;
	wire [3-1:0] node228;
	wire [3-1:0] node230;
	wire [3-1:0] node232;
	wire [3-1:0] node236;
	wire [3-1:0] node237;
	wire [3-1:0] node239;
	wire [3-1:0] node242;
	wire [3-1:0] node243;
	wire [3-1:0] node245;
	wire [3-1:0] node247;
	wire [3-1:0] node250;
	wire [3-1:0] node252;
	wire [3-1:0] node254;

	assign outp = (inp[2]) ? node102 : node1;
		assign node1 = (inp[3]) ? node51 : node2;
			assign node2 = (inp[10]) ? node26 : node3;
				assign node3 = (inp[5]) ? node13 : node4;
					assign node4 = (inp[4]) ? node6 : 3'b111;
						assign node6 = (inp[7]) ? node8 : 3'b110;
							assign node8 = (inp[8]) ? node10 : 3'b110;
								assign node10 = (inp[9]) ? 3'b111 : 3'b110;
					assign node13 = (inp[4]) ? 3'b111 : node14;
						assign node14 = (inp[7]) ? node16 : 3'b111;
							assign node16 = (inp[9]) ? node18 : 3'b111;
								assign node18 = (inp[11]) ? node20 : 3'b111;
									assign node20 = (inp[6]) ? node22 : 3'b111;
										assign node22 = (inp[8]) ? 3'b110 : 3'b111;
				assign node26 = (inp[4]) ? node36 : node27;
					assign node27 = (inp[8]) ? node29 : 3'b110;
						assign node29 = (inp[9]) ? node31 : 3'b110;
							assign node31 = (inp[5]) ? node33 : 3'b110;
								assign node33 = (inp[7]) ? 3'b111 : 3'b110;
					assign node36 = (inp[5]) ? node48 : node37;
						assign node37 = (inp[9]) ? 3'b110 : node38;
							assign node38 = (inp[7]) ? 3'b110 : node39;
								assign node39 = (inp[8]) ? node41 : 3'b111;
									assign node41 = (inp[11]) ? node43 : 3'b111;
										assign node43 = (inp[6]) ? 3'b110 : 3'b111;
						assign node48 = (inp[9]) ? 3'b011 : 3'b110;
			assign node51 = (inp[4]) ? node71 : node52;
				assign node52 = (inp[10]) ? node66 : node53;
					assign node53 = (inp[9]) ? node55 : 3'b111;
						assign node55 = (inp[5]) ? node57 : 3'b111;
							assign node57 = (inp[7]) ? 3'b110 : node58;
								assign node58 = (inp[6]) ? node60 : 3'b111;
									assign node60 = (inp[8]) ? node62 : 3'b111;
										assign node62 = (inp[11]) ? 3'b110 : 3'b111;
					assign node66 = (inp[9]) ? node68 : 3'b110;
						assign node68 = (inp[5]) ? 3'b011 : 3'b110;
				assign node71 = (inp[5]) ? node93 : node72;
					assign node72 = (inp[9]) ? node74 : 3'b011;
						assign node74 = (inp[10]) ? node84 : node75;
							assign node75 = (inp[7]) ? 3'b010 : node76;
								assign node76 = (inp[8]) ? node78 : 3'b011;
									assign node78 = (inp[6]) ? node80 : 3'b011;
										assign node80 = (inp[11]) ? 3'b010 : 3'b011;
							assign node84 = (inp[8]) ? node86 : 3'b011;
								assign node86 = (inp[11]) ? node88 : 3'b011;
									assign node88 = (inp[7]) ? node90 : 3'b011;
										assign node90 = (inp[6]) ? 3'b010 : 3'b011;
					assign node93 = (inp[8]) ? node95 : 3'b010;
						assign node95 = (inp[9]) ? node97 : 3'b010;
							assign node97 = (inp[10]) ? 3'b010 : node98;
								assign node98 = (inp[7]) ? 3'b011 : 3'b010;
		assign node102 = (inp[4]) ? node156 : node103;
			assign node103 = (inp[10]) ? node133 : node104;
				assign node104 = (inp[5]) ? node118 : node105;
					assign node105 = (inp[3]) ? node107 : 3'b011;
						assign node107 = (inp[9]) ? 3'b010 : node108;
							assign node108 = (inp[6]) ? node110 : 3'b011;
								assign node110 = (inp[8]) ? node112 : 3'b011;
									assign node112 = (inp[11]) ? node114 : 3'b011;
										assign node114 = (inp[7]) ? 3'b010 : 3'b011;
					assign node118 = (inp[3]) ? 3'b010 : node119;
						assign node119 = (inp[9]) ? 3'b010 : node120;
							assign node120 = (inp[7]) ? 3'b010 : node121;
								assign node121 = (inp[11]) ? node123 : 3'b011;
									assign node123 = (inp[0]) ? 3'b011 : node124;
										assign node124 = (inp[8]) ? node126 : 3'b011;
											assign node126 = (inp[6]) ? 3'b010 : 3'b011;
				assign node133 = (inp[3]) ? node143 : node134;
					assign node134 = (inp[5]) ? 3'b011 : node135;
						assign node135 = (inp[7]) ? node137 : 3'b010;
							assign node137 = (inp[9]) ? node139 : 3'b010;
								assign node139 = (inp[8]) ? 3'b011 : 3'b010;
					assign node143 = (inp[5]) ? node145 : 3'b111;
						assign node145 = (inp[9]) ? 3'b110 : node146;
							assign node146 = (inp[8]) ? node148 : 3'b111;
								assign node148 = (inp[11]) ? node150 : 3'b111;
									assign node150 = (inp[6]) ? node152 : 3'b111;
										assign node152 = (inp[7]) ? 3'b110 : 3'b111;
			assign node156 = (inp[3]) ? node188 : node157;
				assign node157 = (inp[5]) ? node179 : node158;
					assign node158 = (inp[9]) ? node160 : 3'b101;
						assign node160 = (inp[7]) ? node170 : node161;
							assign node161 = (inp[10]) ? node163 : 3'b101;
								assign node163 = (inp[11]) ? node165 : 3'b101;
									assign node165 = (inp[6]) ? node167 : 3'b101;
										assign node167 = (inp[8]) ? 3'b100 : 3'b101;
							assign node170 = (inp[10]) ? 3'b100 : node171;
								assign node171 = (inp[6]) ? node173 : 3'b101;
									assign node173 = (inp[11]) ? node175 : 3'b101;
										assign node175 = (inp[8]) ? 3'b100 : 3'b101;
					assign node179 = (inp[9]) ? node181 : 3'b100;
						assign node181 = (inp[10]) ? 3'b001 : node182;
							assign node182 = (inp[8]) ? node184 : 3'b100;
								assign node184 = (inp[7]) ? 3'b101 : 3'b100;
				assign node188 = (inp[10]) ? node216 : node189;
					assign node189 = (inp[9]) ? node209 : node190;
						assign node190 = (inp[5]) ? node200 : node191;
							assign node191 = (inp[7]) ? 3'b000 : node192;
								assign node192 = (inp[8]) ? node194 : 3'b001;
									assign node194 = (inp[6]) ? node196 : 3'b001;
										assign node196 = (inp[11]) ? 3'b000 : 3'b001;
							assign node200 = (inp[6]) ? node202 : 3'b001;
								assign node202 = (inp[11]) ? node204 : 3'b001;
									assign node204 = (inp[8]) ? node206 : 3'b001;
										assign node206 = (inp[7]) ? 3'b000 : 3'b001;
						assign node209 = (inp[8]) ? node211 : 3'b000;
							assign node211 = (inp[7]) ? node213 : 3'b000;
								assign node213 = (inp[5]) ? 3'b000 : 3'b001;
					assign node216 = (inp[9]) ? node236 : node217;
						assign node217 = (inp[7]) ? node227 : node218;
							assign node218 = (inp[8]) ? node220 : 3'b101;
								assign node220 = (inp[11]) ? node222 : 3'b101;
									assign node222 = (inp[5]) ? node224 : 3'b101;
										assign node224 = (inp[1]) ? 3'b101 : 3'b100;
							assign node227 = (inp[5]) ? 3'b100 : node228;
								assign node228 = (inp[11]) ? node230 : 3'b101;
									assign node230 = (inp[6]) ? node232 : 3'b101;
										assign node232 = (inp[8]) ? 3'b100 : 3'b101;
						assign node236 = (inp[5]) ? node242 : node237;
							assign node237 = (inp[7]) ? node239 : 3'b100;
								assign node239 = (inp[8]) ? 3'b101 : 3'b100;
							assign node242 = (inp[7]) ? node250 : node243;
								assign node243 = (inp[6]) ? node245 : 3'b001;
									assign node245 = (inp[11]) ? node247 : 3'b001;
										assign node247 = (inp[8]) ? 3'b000 : 3'b001;
								assign node250 = (inp[8]) ? node252 : 3'b000;
									assign node252 = (inp[11]) ? node254 : 3'b001;
										assign node254 = (inp[6]) ? 3'b000 : 3'b001;

endmodule