module dtc_split125_bm59 (
	input  wire [12-1:0] inp,
	output wire [3-1:0] outp
);

	wire [3-1:0] node1;
	wire [3-1:0] node2;
	wire [3-1:0] node3;
	wire [3-1:0] node4;
	wire [3-1:0] node5;
	wire [3-1:0] node6;
	wire [3-1:0] node7;
	wire [3-1:0] node8;
	wire [3-1:0] node12;
	wire [3-1:0] node15;
	wire [3-1:0] node16;
	wire [3-1:0] node19;
	wire [3-1:0] node22;
	wire [3-1:0] node24;
	wire [3-1:0] node25;
	wire [3-1:0] node26;
	wire [3-1:0] node27;
	wire [3-1:0] node31;
	wire [3-1:0] node34;
	wire [3-1:0] node38;
	wire [3-1:0] node39;
	wire [3-1:0] node40;
	wire [3-1:0] node41;
	wire [3-1:0] node42;
	wire [3-1:0] node43;
	wire [3-1:0] node47;
	wire [3-1:0] node49;
	wire [3-1:0] node52;
	wire [3-1:0] node53;
	wire [3-1:0] node56;
	wire [3-1:0] node58;
	wire [3-1:0] node60;
	wire [3-1:0] node63;
	wire [3-1:0] node64;
	wire [3-1:0] node66;
	wire [3-1:0] node70;
	wire [3-1:0] node71;
	wire [3-1:0] node72;
	wire [3-1:0] node73;
	wire [3-1:0] node74;
	wire [3-1:0] node78;
	wire [3-1:0] node79;
	wire [3-1:0] node83;
	wire [3-1:0] node86;
	wire [3-1:0] node87;
	wire [3-1:0] node88;
	wire [3-1:0] node91;
	wire [3-1:0] node93;
	wire [3-1:0] node94;
	wire [3-1:0] node98;
	wire [3-1:0] node99;
	wire [3-1:0] node101;
	wire [3-1:0] node104;
	wire [3-1:0] node107;
	wire [3-1:0] node108;
	wire [3-1:0] node109;
	wire [3-1:0] node110;
	wire [3-1:0] node112;
	wire [3-1:0] node114;
	wire [3-1:0] node117;
	wire [3-1:0] node118;
	wire [3-1:0] node119;
	wire [3-1:0] node120;
	wire [3-1:0] node125;
	wire [3-1:0] node127;
	wire [3-1:0] node128;
	wire [3-1:0] node132;
	wire [3-1:0] node133;
	wire [3-1:0] node134;
	wire [3-1:0] node135;
	wire [3-1:0] node139;
	wire [3-1:0] node140;
	wire [3-1:0] node144;
	wire [3-1:0] node145;
	wire [3-1:0] node146;
	wire [3-1:0] node147;
	wire [3-1:0] node152;
	wire [3-1:0] node153;
	wire [3-1:0] node154;
	wire [3-1:0] node158;
	wire [3-1:0] node161;
	wire [3-1:0] node163;
	wire [3-1:0] node165;
	wire [3-1:0] node166;
	wire [3-1:0] node167;
	wire [3-1:0] node168;
	wire [3-1:0] node172;
	wire [3-1:0] node173;
	wire [3-1:0] node177;
	wire [3-1:0] node180;
	wire [3-1:0] node181;
	wire [3-1:0] node182;
	wire [3-1:0] node183;
	wire [3-1:0] node184;
	wire [3-1:0] node185;
	wire [3-1:0] node187;
	wire [3-1:0] node189;
	wire [3-1:0] node193;
	wire [3-1:0] node194;
	wire [3-1:0] node195;
	wire [3-1:0] node196;
	wire [3-1:0] node197;
	wire [3-1:0] node201;
	wire [3-1:0] node205;
	wire [3-1:0] node207;
	wire [3-1:0] node211;
	wire [3-1:0] node212;
	wire [3-1:0] node213;
	wire [3-1:0] node214;
	wire [3-1:0] node215;
	wire [3-1:0] node218;
	wire [3-1:0] node219;
	wire [3-1:0] node220;
	wire [3-1:0] node225;
	wire [3-1:0] node228;
	wire [3-1:0] node229;
	wire [3-1:0] node230;
	wire [3-1:0] node232;
	wire [3-1:0] node235;
	wire [3-1:0] node237;
	wire [3-1:0] node241;
	wire [3-1:0] node242;
	wire [3-1:0] node244;
	wire [3-1:0] node246;
	wire [3-1:0] node247;
	wire [3-1:0] node250;
	wire [3-1:0] node253;
	wire [3-1:0] node254;
	wire [3-1:0] node256;
	wire [3-1:0] node257;
	wire [3-1:0] node262;
	wire [3-1:0] node263;
	wire [3-1:0] node264;
	wire [3-1:0] node266;
	wire [3-1:0] node267;
	wire [3-1:0] node270;
	wire [3-1:0] node272;
	wire [3-1:0] node273;
	wire [3-1:0] node276;
	wire [3-1:0] node278;
	wire [3-1:0] node282;
	wire [3-1:0] node283;
	wire [3-1:0] node284;
	wire [3-1:0] node285;
	wire [3-1:0] node286;
	wire [3-1:0] node289;
	wire [3-1:0] node290;
	wire [3-1:0] node292;
	wire [3-1:0] node295;
	wire [3-1:0] node298;
	wire [3-1:0] node299;
	wire [3-1:0] node301;
	wire [3-1:0] node304;
	wire [3-1:0] node305;
	wire [3-1:0] node309;
	wire [3-1:0] node310;
	wire [3-1:0] node311;
	wire [3-1:0] node312;
	wire [3-1:0] node314;
	wire [3-1:0] node320;
	wire [3-1:0] node322;
	wire [3-1:0] node323;
	wire [3-1:0] node324;
	wire [3-1:0] node325;
	wire [3-1:0] node328;
	wire [3-1:0] node329;
	wire [3-1:0] node333;

	assign outp = (inp[10]) ? node180 : node1;
		assign node1 = (inp[9]) ? node107 : node2;
			assign node2 = (inp[2]) ? node38 : node3;
				assign node3 = (inp[0]) ? 3'b110 : node4;
					assign node4 = (inp[3]) ? node22 : node5;
						assign node5 = (inp[7]) ? node15 : node6;
							assign node6 = (inp[5]) ? node12 : node7;
								assign node7 = (inp[11]) ? 3'b000 : node8;
									assign node8 = (inp[8]) ? 3'b100 : 3'b111;
								assign node12 = (inp[4]) ? 3'b010 : 3'b000;
							assign node15 = (inp[6]) ? node19 : node16;
								assign node16 = (inp[5]) ? 3'b110 : 3'b100;
								assign node19 = (inp[5]) ? 3'b100 : 3'b010;
						assign node22 = (inp[1]) ? node24 : 3'b111;
							assign node24 = (inp[4]) ? node34 : node25;
								assign node25 = (inp[7]) ? node31 : node26;
									assign node26 = (inp[8]) ? 3'b111 : node27;
										assign node27 = (inp[6]) ? 3'b111 : 3'b000;
									assign node31 = (inp[11]) ? 3'b010 : 3'b100;
								assign node34 = (inp[7]) ? 3'b100 : 3'b000;
				assign node38 = (inp[1]) ? node70 : node39;
					assign node39 = (inp[3]) ? node63 : node40;
						assign node40 = (inp[11]) ? node52 : node41;
							assign node41 = (inp[5]) ? node47 : node42;
								assign node42 = (inp[4]) ? 3'b010 : node43;
									assign node43 = (inp[7]) ? 3'b000 : 3'b110;
								assign node47 = (inp[0]) ? node49 : 3'b000;
									assign node49 = (inp[4]) ? 3'b000 : 3'b110;
							assign node52 = (inp[8]) ? node56 : node53;
								assign node53 = (inp[5]) ? 3'b010 : 3'b000;
								assign node56 = (inp[0]) ? node58 : 3'b010;
									assign node58 = (inp[7]) ? node60 : 3'b110;
										assign node60 = (inp[4]) ? 3'b110 : 3'b010;
						assign node63 = (inp[0]) ? 3'b110 : node64;
							assign node64 = (inp[11]) ? node66 : 3'b100;
								assign node66 = (inp[4]) ? 3'b110 : 3'b010;
					assign node70 = (inp[0]) ? node86 : node71;
						assign node71 = (inp[7]) ? node83 : node72;
							assign node72 = (inp[11]) ? node78 : node73;
								assign node73 = (inp[5]) ? 3'b010 : node74;
									assign node74 = (inp[6]) ? 3'b100 : 3'b010;
								assign node78 = (inp[6]) ? 3'b010 : node79;
									assign node79 = (inp[4]) ? 3'b010 : 3'b110;
							assign node83 = (inp[4]) ? 3'b000 : 3'b010;
						assign node86 = (inp[11]) ? node98 : node87;
							assign node87 = (inp[4]) ? node91 : node88;
								assign node88 = (inp[3]) ? 3'b010 : 3'b000;
								assign node91 = (inp[6]) ? node93 : 3'b000;
									assign node93 = (inp[7]) ? 3'b000 : node94;
										assign node94 = (inp[3]) ? 3'b000 : 3'b100;
							assign node98 = (inp[4]) ? node104 : node99;
								assign node99 = (inp[6]) ? node101 : 3'b010;
									assign node101 = (inp[3]) ? 3'b010 : 3'b000;
								assign node104 = (inp[6]) ? 3'b010 : 3'b000;
			assign node107 = (inp[0]) ? node161 : node108;
				assign node108 = (inp[2]) ? node132 : node109;
					assign node109 = (inp[1]) ? node117 : node110;
						assign node110 = (inp[7]) ? node112 : 3'b011;
							assign node112 = (inp[4]) ? node114 : 3'b011;
								assign node114 = (inp[5]) ? 3'b010 : 3'b011;
						assign node117 = (inp[4]) ? node125 : node118;
							assign node118 = (inp[3]) ? 3'b011 : node119;
								assign node119 = (inp[7]) ? 3'b100 : node120;
									assign node120 = (inp[5]) ? 3'b100 : 3'b010;
							assign node125 = (inp[6]) ? node127 : 3'b010;
								assign node127 = (inp[8]) ? 3'b000 : node128;
									assign node128 = (inp[5]) ? 3'b000 : 3'b010;
					assign node132 = (inp[8]) ? node144 : node133;
						assign node133 = (inp[7]) ? node139 : node134;
							assign node134 = (inp[6]) ? 3'b100 : node135;
								assign node135 = (inp[1]) ? 3'b000 : 3'b100;
							assign node139 = (inp[3]) ? 3'b000 : node140;
								assign node140 = (inp[11]) ? 3'b000 : 3'b010;
						assign node144 = (inp[3]) ? node152 : node145;
							assign node145 = (inp[4]) ? 3'b000 : node146;
								assign node146 = (inp[5]) ? 3'b000 : node147;
									assign node147 = (inp[1]) ? 3'b010 : 3'b000;
							assign node152 = (inp[7]) ? node158 : node153;
								assign node153 = (inp[6]) ? 3'b010 : node154;
									assign node154 = (inp[11]) ? 3'b110 : 3'b010;
								assign node158 = (inp[11]) ? 3'b010 : 3'b000;
				assign node161 = (inp[2]) ? node163 : 3'b010;
					assign node163 = (inp[7]) ? node165 : 3'b010;
						assign node165 = (inp[4]) ? node177 : node166;
							assign node166 = (inp[3]) ? node172 : node167;
								assign node167 = (inp[6]) ? 3'b000 : node168;
									assign node168 = (inp[5]) ? 3'b000 : 3'b010;
								assign node172 = (inp[8]) ? 3'b010 : node173;
									assign node173 = (inp[6]) ? 3'b000 : 3'b010;
							assign node177 = (inp[1]) ? 3'b000 : 3'b010;
		assign node180 = (inp[9]) ? node262 : node181;
			assign node181 = (inp[2]) ? node211 : node182;
				assign node182 = (inp[0]) ? 3'b100 : node183;
					assign node183 = (inp[1]) ? node193 : node184;
						assign node184 = (inp[3]) ? 3'b101 : node185;
							assign node185 = (inp[7]) ? node187 : 3'b101;
								assign node187 = (inp[4]) ? node189 : 3'b010;
									assign node189 = (inp[8]) ? 3'b000 : 3'b100;
						assign node193 = (inp[5]) ? node205 : node194;
							assign node194 = (inp[3]) ? 3'b010 : node195;
								assign node195 = (inp[8]) ? node201 : node196;
									assign node196 = (inp[11]) ? 3'b110 : node197;
										assign node197 = (inp[4]) ? 3'b110 : 3'b010;
									assign node201 = (inp[6]) ? 3'b100 : 3'b110;
							assign node205 = (inp[6]) ? node207 : 3'b100;
								assign node207 = (inp[11]) ? 3'b000 : 3'b010;
				assign node211 = (inp[1]) ? node241 : node212;
					assign node212 = (inp[0]) ? node228 : node213;
						assign node213 = (inp[11]) ? node225 : node214;
							assign node214 = (inp[4]) ? node218 : node215;
								assign node215 = (inp[5]) ? 3'b110 : 3'b100;
								assign node218 = (inp[5]) ? 3'b110 : node219;
									assign node219 = (inp[7]) ? 3'b010 : node220;
										assign node220 = (inp[8]) ? 3'b110 : 3'b010;
							assign node225 = (inp[3]) ? 3'b000 : 3'b110;
						assign node228 = (inp[3]) ? 3'b100 : node229;
							assign node229 = (inp[6]) ? node235 : node230;
								assign node230 = (inp[7]) ? node232 : 3'b100;
									assign node232 = (inp[4]) ? 3'b100 : 3'b000;
								assign node235 = (inp[4]) ? node237 : 3'b010;
									assign node237 = (inp[7]) ? 3'b100 : 3'b000;
					assign node241 = (inp[11]) ? node253 : node242;
						assign node242 = (inp[0]) ? node244 : 3'b000;
							assign node244 = (inp[4]) ? node246 : 3'b010;
								assign node246 = (inp[3]) ? node250 : node247;
									assign node247 = (inp[6]) ? 3'b000 : 3'b010;
									assign node250 = (inp[8]) ? 3'b100 : 3'b000;
						assign node253 = (inp[5]) ? 3'b000 : node254;
							assign node254 = (inp[7]) ? node256 : 3'b010;
								assign node256 = (inp[6]) ? 3'b000 : node257;
									assign node257 = (inp[8]) ? 3'b000 : 3'b010;
			assign node262 = (inp[2]) ? node282 : node263;
				assign node263 = (inp[0]) ? 3'b000 : node264;
					assign node264 = (inp[1]) ? node266 : 3'b001;
						assign node266 = (inp[3]) ? node270 : node267;
							assign node267 = (inp[8]) ? 3'b000 : 3'b010;
							assign node270 = (inp[7]) ? node272 : 3'b001;
								assign node272 = (inp[8]) ? node276 : node273;
									assign node273 = (inp[11]) ? 3'b000 : 3'b010;
									assign node276 = (inp[4]) ? node278 : 3'b001;
										assign node278 = (inp[11]) ? 3'b000 : 3'b001;
				assign node282 = (inp[0]) ? node320 : node283;
					assign node283 = (inp[11]) ? node309 : node284;
						assign node284 = (inp[1]) ? node298 : node285;
							assign node285 = (inp[3]) ? node289 : node286;
								assign node286 = (inp[4]) ? 3'b110 : 3'b010;
								assign node289 = (inp[8]) ? node295 : node290;
									assign node290 = (inp[7]) ? node292 : 3'b110;
										assign node292 = (inp[5]) ? 3'b110 : 3'b100;
									assign node295 = (inp[7]) ? 3'b110 : 3'b100;
							assign node298 = (inp[7]) ? node304 : node299;
								assign node299 = (inp[5]) ? node301 : 3'b010;
									assign node301 = (inp[4]) ? 3'b010 : 3'b110;
								assign node304 = (inp[4]) ? 3'b000 : node305;
									assign node305 = (inp[6]) ? 3'b010 : 3'b000;
						assign node309 = (inp[6]) ? 3'b000 : node310;
							assign node310 = (inp[1]) ? 3'b000 : node311;
								assign node311 = (inp[3]) ? 3'b100 : node312;
									assign node312 = (inp[8]) ? node314 : 3'b000;
										assign node314 = (inp[5]) ? 3'b000 : 3'b100;
					assign node320 = (inp[1]) ? node322 : 3'b000;
						assign node322 = (inp[3]) ? 3'b000 : node323;
							assign node323 = (inp[8]) ? node333 : node324;
								assign node324 = (inp[4]) ? node328 : node325;
									assign node325 = (inp[7]) ? 3'b000 : 3'b010;
									assign node328 = (inp[5]) ? 3'b000 : node329;
										assign node329 = (inp[7]) ? 3'b000 : 3'b100;
								assign node333 = (inp[5]) ? 3'b000 : 3'b010;

endmodule