module dtc_split125_bm34 (
	input  wire [9-1:0] inp,
	output wire [5-1:0] outp
);

	wire [5-1:0] node1;
	wire [5-1:0] node2;
	wire [5-1:0] node3;
	wire [5-1:0] node4;
	wire [5-1:0] node7;
	wire [5-1:0] node8;
	wire [5-1:0] node11;
	wire [5-1:0] node14;
	wire [5-1:0] node15;
	wire [5-1:0] node17;
	wire [5-1:0] node20;
	wire [5-1:0] node22;
	wire [5-1:0] node23;
	wire [5-1:0] node27;
	wire [5-1:0] node28;
	wire [5-1:0] node29;
	wire [5-1:0] node30;
	wire [5-1:0] node31;
	wire [5-1:0] node36;
	wire [5-1:0] node37;
	wire [5-1:0] node40;
	wire [5-1:0] node43;
	wire [5-1:0] node44;
	wire [5-1:0] node47;
	wire [5-1:0] node48;
	wire [5-1:0] node50;
	wire [5-1:0] node54;
	wire [5-1:0] node55;
	wire [5-1:0] node56;
	wire [5-1:0] node57;
	wire [5-1:0] node60;
	wire [5-1:0] node61;
	wire [5-1:0] node63;
	wire [5-1:0] node66;
	wire [5-1:0] node67;
	wire [5-1:0] node71;
	wire [5-1:0] node73;
	wire [5-1:0] node75;
	wire [5-1:0] node77;
	wire [5-1:0] node80;
	wire [5-1:0] node81;
	wire [5-1:0] node82;
	wire [5-1:0] node85;
	wire [5-1:0] node87;
	wire [5-1:0] node90;
	wire [5-1:0] node91;
	wire [5-1:0] node94;
	wire [5-1:0] node95;
	wire [5-1:0] node97;

	assign outp = (inp[2]) ? node54 : node1;
		assign node1 = (inp[7]) ? node27 : node2;
			assign node2 = (inp[0]) ? node14 : node3;
				assign node3 = (inp[8]) ? node7 : node4;
					assign node4 = (inp[5]) ? 5'b01010 : 5'b00111;
					assign node7 = (inp[4]) ? node11 : node8;
						assign node8 = (inp[1]) ? 5'b01000 : 5'b00000;
						assign node11 = (inp[5]) ? 5'b00000 : 5'b00001;
				assign node14 = (inp[8]) ? node20 : node15;
					assign node15 = (inp[6]) ? node17 : 5'b00010;
						assign node17 = (inp[5]) ? 5'b00010 : 5'b10011;
					assign node20 = (inp[5]) ? node22 : 5'b00110;
						assign node22 = (inp[6]) ? 5'b01011 : node23;
							assign node23 = (inp[1]) ? 5'b11010 : 5'b01011;
			assign node27 = (inp[0]) ? node43 : node28;
				assign node28 = (inp[1]) ? node36 : node29;
					assign node29 = (inp[4]) ? 5'b11110 : node30;
						assign node30 = (inp[3]) ? 5'b10111 : node31;
							assign node31 = (inp[8]) ? 5'b11110 : 5'b10110;
					assign node36 = (inp[6]) ? node40 : node37;
						assign node37 = (inp[8]) ? 5'b11111 : 5'b10110;
						assign node40 = (inp[5]) ? 5'b01011 : 5'b01110;
				assign node43 = (inp[8]) ? node47 : node44;
					assign node44 = (inp[3]) ? 5'b10011 : 5'b00010;
					assign node47 = (inp[4]) ? 5'b11010 : node48;
						assign node48 = (inp[3]) ? node50 : 5'b11010;
							assign node50 = (inp[1]) ? 5'b11011 : 5'b10011;
		assign node54 = (inp[8]) ? node80 : node55;
			assign node55 = (inp[7]) ? node71 : node56;
				assign node56 = (inp[0]) ? node60 : node57;
					assign node57 = (inp[5]) ? 5'b01001 : 5'b11001;
					assign node60 = (inp[5]) ? node66 : node61;
						assign node61 = (inp[3]) ? node63 : 5'b01111;
							assign node63 = (inp[6]) ? 5'b00001 : 5'b00000;
						assign node66 = (inp[1]) ? 5'b10111 : node67;
							assign node67 = (inp[4]) ? 5'b01110 : 5'b01111;
				assign node71 = (inp[6]) ? node73 : 5'b00100;
					assign node73 = (inp[5]) ? node75 : 5'b11101;
						assign node75 = (inp[0]) ? node77 : 5'b10100;
							assign node77 = (inp[3]) ? 5'b10000 : 5'b11111;
			assign node80 = (inp[7]) ? node90 : node81;
				assign node81 = (inp[5]) ? node85 : node82;
					assign node82 = (inp[0]) ? 5'b01100 : 5'b11101;
					assign node85 = (inp[6]) ? node87 : 5'b11100;
						assign node87 = (inp[1]) ? 5'b01100 : 5'b11100;
				assign node90 = (inp[1]) ? node94 : node91;
					assign node91 = (inp[5]) ? 5'b01001 : 5'b11001;
					assign node94 = (inp[6]) ? 5'b01100 : node95;
						assign node95 = (inp[0]) ? node97 : 5'b10100;
							assign node97 = (inp[4]) ? 5'b11000 : 5'b10100;

endmodule