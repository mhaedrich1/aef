module dtc_split125_bm32 (
	input  wire [15-1:0] inp,
	output wire [9-1:0] outp
);

	wire [9-1:0] node1;
	wire [9-1:0] node2;
	wire [9-1:0] node5;
	wire [9-1:0] node6;
	wire [9-1:0] node7;
	wire [9-1:0] node9;
	wire [9-1:0] node11;
	wire [9-1:0] node13;
	wire [9-1:0] node14;
	wire [9-1:0] node18;
	wire [9-1:0] node21;
	wire [9-1:0] node22;
	wire [9-1:0] node24;
	wire [9-1:0] node26;
	wire [9-1:0] node29;
	wire [9-1:0] node30;
	wire [9-1:0] node32;
	wire [9-1:0] node34;
	wire [9-1:0] node35;
	wire [9-1:0] node39;
	wire [9-1:0] node41;
	wire [9-1:0] node43;
	wire [9-1:0] node46;
	wire [9-1:0] node47;
	wire [9-1:0] node48;
	wire [9-1:0] node49;
	wire [9-1:0] node50;
	wire [9-1:0] node51;
	wire [9-1:0] node52;
	wire [9-1:0] node53;
	wire [9-1:0] node58;
	wire [9-1:0] node59;
	wire [9-1:0] node60;
	wire [9-1:0] node61;
	wire [9-1:0] node62;
	wire [9-1:0] node66;
	wire [9-1:0] node70;
	wire [9-1:0] node73;
	wire [9-1:0] node74;
	wire [9-1:0] node75;
	wire [9-1:0] node76;
	wire [9-1:0] node81;
	wire [9-1:0] node82;
	wire [9-1:0] node83;
	wire [9-1:0] node84;
	wire [9-1:0] node89;
	wire [9-1:0] node92;
	wire [9-1:0] node93;
	wire [9-1:0] node94;
	wire [9-1:0] node95;
	wire [9-1:0] node97;
	wire [9-1:0] node99;
	wire [9-1:0] node102;
	wire [9-1:0] node104;
	wire [9-1:0] node107;
	wire [9-1:0] node108;
	wire [9-1:0] node111;
	wire [9-1:0] node114;
	wire [9-1:0] node115;
	wire [9-1:0] node116;
	wire [9-1:0] node117;
	wire [9-1:0] node118;
	wire [9-1:0] node119;
	wire [9-1:0] node122;
	wire [9-1:0] node125;
	wire [9-1:0] node129;
	wire [9-1:0] node130;
	wire [9-1:0] node131;
	wire [9-1:0] node132;
	wire [9-1:0] node135;
	wire [9-1:0] node139;
	wire [9-1:0] node140;
	wire [9-1:0] node144;
	wire [9-1:0] node145;
	wire [9-1:0] node146;
	wire [9-1:0] node147;
	wire [9-1:0] node148;
	wire [9-1:0] node152;
	wire [9-1:0] node153;
	wire [9-1:0] node156;
	wire [9-1:0] node159;
	wire [9-1:0] node160;
	wire [9-1:0] node163;
	wire [9-1:0] node165;
	wire [9-1:0] node168;
	wire [9-1:0] node170;
	wire [9-1:0] node173;
	wire [9-1:0] node174;
	wire [9-1:0] node175;
	wire [9-1:0] node176;
	wire [9-1:0] node177;
	wire [9-1:0] node178;
	wire [9-1:0] node183;
	wire [9-1:0] node184;
	wire [9-1:0] node186;
	wire [9-1:0] node187;
	wire [9-1:0] node189;
	wire [9-1:0] node193;
	wire [9-1:0] node196;
	wire [9-1:0] node197;
	wire [9-1:0] node198;
	wire [9-1:0] node199;
	wire [9-1:0] node204;
	wire [9-1:0] node205;
	wire [9-1:0] node206;
	wire [9-1:0] node207;
	wire [9-1:0] node212;
	wire [9-1:0] node215;
	wire [9-1:0] node216;
	wire [9-1:0] node217;
	wire [9-1:0] node218;
	wire [9-1:0] node219;
	wire [9-1:0] node224;
	wire [9-1:0] node225;
	wire [9-1:0] node226;
	wire [9-1:0] node227;
	wire [9-1:0] node232;
	wire [9-1:0] node235;
	wire [9-1:0] node236;
	wire [9-1:0] node237;
	wire [9-1:0] node238;
	wire [9-1:0] node239;
	wire [9-1:0] node240;
	wire [9-1:0] node243;
	wire [9-1:0] node247;
	wire [9-1:0] node248;
	wire [9-1:0] node249;
	wire [9-1:0] node250;
	wire [9-1:0] node255;
	wire [9-1:0] node256;
	wire [9-1:0] node260;
	wire [9-1:0] node261;
	wire [9-1:0] node262;
	wire [9-1:0] node263;
	wire [9-1:0] node265;
	wire [9-1:0] node267;
	wire [9-1:0] node271;
	wire [9-1:0] node274;
	wire [9-1:0] node276;
	wire [9-1:0] node279;
	wire [9-1:0] node280;
	wire [9-1:0] node281;
	wire [9-1:0] node282;
	wire [9-1:0] node283;
	wire [9-1:0] node286;
	wire [9-1:0] node290;
	wire [9-1:0] node291;
	wire [9-1:0] node292;
	wire [9-1:0] node293;
	wire [9-1:0] node298;
	wire [9-1:0] node301;
	wire [9-1:0] node302;
	wire [9-1:0] node303;
	wire [9-1:0] node304;
	wire [9-1:0] node305;
	wire [9-1:0] node309;
	wire [9-1:0] node310;
	wire [9-1:0] node314;
	wire [9-1:0] node315;
	wire [9-1:0] node316;
	wire [9-1:0] node321;
	wire [9-1:0] node322;
	wire [9-1:0] node325;
	wire [9-1:0] node328;
	wire [9-1:0] node329;
	wire [9-1:0] node330;
	wire [9-1:0] node331;
	wire [9-1:0] node332;
	wire [9-1:0] node335;
	wire [9-1:0] node337;
	wire [9-1:0] node340;
	wire [9-1:0] node341;
	wire [9-1:0] node344;
	wire [9-1:0] node346;
	wire [9-1:0] node347;
	wire [9-1:0] node350;
	wire [9-1:0] node353;
	wire [9-1:0] node354;
	wire [9-1:0] node356;
	wire [9-1:0] node359;
	wire [9-1:0] node360;
	wire [9-1:0] node363;
	wire [9-1:0] node364;
	wire [9-1:0] node367;
	wire [9-1:0] node368;
	wire [9-1:0] node371;
	wire [9-1:0] node374;
	wire [9-1:0] node375;
	wire [9-1:0] node376;
	wire [9-1:0] node377;
	wire [9-1:0] node380;
	wire [9-1:0] node381;
	wire [9-1:0] node384;
	wire [9-1:0] node387;
	wire [9-1:0] node388;
	wire [9-1:0] node391;
	wire [9-1:0] node393;
	wire [9-1:0] node394;
	wire [9-1:0] node397;
	wire [9-1:0] node400;
	wire [9-1:0] node401;
	wire [9-1:0] node402;
	wire [9-1:0] node405;
	wire [9-1:0] node408;
	wire [9-1:0] node409;
	wire [9-1:0] node412;
	wire [9-1:0] node413;
	wire [9-1:0] node414;
	wire [9-1:0] node417;
	wire [9-1:0] node418;
	wire [9-1:0] node421;
	wire [9-1:0] node424;
	wire [9-1:0] node425;
	wire [9-1:0] node428;
	wire [9-1:0] node429;
	wire [9-1:0] node432;

	assign outp = (inp[12]) ? node46 : node1;
		assign node1 = (inp[13]) ? node5 : node2;
			assign node2 = (inp[11]) ? 9'b101010101 : 9'b101010000;
			assign node5 = (inp[14]) ? node21 : node6;
				assign node6 = (inp[0]) ? node18 : node7;
					assign node7 = (inp[3]) ? node9 : 9'b101010001;
						assign node9 = (inp[8]) ? node11 : 9'b100010001;
							assign node11 = (inp[9]) ? node13 : 9'b100010001;
								assign node13 = (inp[4]) ? 9'b100010001 : node14;
									assign node14 = (inp[6]) ? 9'b001010001 : 9'b101010001;
					assign node18 = (inp[3]) ? 9'b000010101 : 9'b101010101;
				assign node21 = (inp[3]) ? node29 : node22;
					assign node22 = (inp[8]) ? node24 : 9'b111010101;
						assign node24 = (inp[9]) ? node26 : 9'b101010101;
							assign node26 = (inp[4]) ? 9'b111010101 : 9'b101010101;
					assign node29 = (inp[0]) ? node39 : node30;
						assign node30 = (inp[8]) ? node32 : 9'b111010111;
							assign node32 = (inp[9]) ? node34 : 9'b101010111;
								assign node34 = (inp[4]) ? 9'b111010111 : node35;
									assign node35 = (inp[6]) ? 9'b011010101 : 9'b111010101;
						assign node39 = (inp[8]) ? node41 : 9'b011010111;
							assign node41 = (inp[9]) ? node43 : 9'b001010111;
								assign node43 = (inp[4]) ? 9'b001010101 : 9'b000010111;
		assign node46 = (inp[8]) ? node328 : node47;
			assign node47 = (inp[6]) ? node173 : node48;
				assign node48 = (inp[13]) ? node92 : node49;
					assign node49 = (inp[11]) ? node73 : node50;
						assign node50 = (inp[7]) ? node58 : node51;
							assign node51 = (inp[1]) ? 9'b111011000 : node52;
								assign node52 = (inp[9]) ? 9'b111011000 : node53;
									assign node53 = (inp[2]) ? 9'b111111000 : 9'b111110000;
							assign node58 = (inp[4]) ? node70 : node59;
								assign node59 = (inp[9]) ? 9'b111111000 : node60;
									assign node60 = (inp[3]) ? node66 : node61;
										assign node61 = (inp[2]) ? 9'b111111000 : node62;
											assign node62 = (inp[1]) ? 9'b111111000 : 9'b111110000;
										assign node66 = (inp[1]) ? 9'b111111000 : 9'b111110000;
								assign node70 = (inp[9]) ? 9'b111010000 : 9'b111110000;
						assign node73 = (inp[7]) ? node81 : node74;
							assign node74 = (inp[9]) ? 9'b111011100 : node75;
								assign node75 = (inp[1]) ? 9'b111011100 : node76;
									assign node76 = (inp[2]) ? 9'b111111100 : 9'b111110100;
							assign node81 = (inp[4]) ? node89 : node82;
								assign node82 = (inp[2]) ? 9'b111111100 : node83;
									assign node83 = (inp[9]) ? 9'b111111100 : node84;
										assign node84 = (inp[1]) ? 9'b111111100 : 9'b111110100;
								assign node89 = (inp[9]) ? 9'b111010100 : 9'b111110100;
					assign node92 = (inp[3]) ? node114 : node93;
						assign node93 = (inp[9]) ? node107 : node94;
							assign node94 = (inp[1]) ? node102 : node95;
								assign node95 = (inp[2]) ? node97 : 9'b111110100;
									assign node97 = (inp[7]) ? node99 : 9'b111111100;
										assign node99 = (inp[4]) ? 9'b111110100 : 9'b111111100;
								assign node102 = (inp[7]) ? node104 : 9'b111011100;
									assign node104 = (inp[4]) ? 9'b111110100 : 9'b111111100;
							assign node107 = (inp[4]) ? node111 : node108;
								assign node108 = (inp[7]) ? 9'b111111100 : 9'b111011100;
								assign node111 = (inp[7]) ? 9'b111010100 : 9'b111011100;
						assign node114 = (inp[14]) ? node144 : node115;
							assign node115 = (inp[7]) ? node129 : node116;
								assign node116 = (inp[9]) ? 9'b110011110 : node117;
									assign node117 = (inp[1]) ? node125 : node118;
										assign node118 = (inp[10]) ? node122 : node119;
											assign node119 = (inp[2]) ? 9'b110111100 : 9'b110110100;
											assign node122 = (inp[2]) ? 9'b110111110 : 9'b110110110;
										assign node125 = (inp[10]) ? 9'b110011110 : 9'b110011100;
								assign node129 = (inp[4]) ? node139 : node130;
									assign node130 = (inp[9]) ? 9'b110111110 : node131;
										assign node131 = (inp[10]) ? node135 : node132;
											assign node132 = (inp[2]) ? 9'b110111100 : 9'b110110100;
											assign node135 = (inp[5]) ? 9'b110111110 : 9'b110110110;
									assign node139 = (inp[9]) ? 9'b110010110 : node140;
										assign node140 = (inp[11]) ? 9'b110110110 : 9'b110110100;
							assign node144 = (inp[9]) ? node168 : node145;
								assign node145 = (inp[10]) ? node159 : node146;
									assign node146 = (inp[11]) ? node152 : node147;
										assign node147 = (inp[7]) ? 9'b111111100 : node148;
											assign node148 = (inp[1]) ? 9'b111011100 : 9'b111111100;
										assign node152 = (inp[7]) ? node156 : node153;
											assign node153 = (inp[1]) ? 9'b111011100 : 9'b111110100;
											assign node156 = (inp[4]) ? 9'b111110100 : 9'b111111100;
									assign node159 = (inp[1]) ? node163 : node160;
										assign node160 = (inp[2]) ? 9'b111111110 : 9'b111110110;
										assign node163 = (inp[7]) ? node165 : 9'b111011110;
											assign node165 = (inp[5]) ? 9'b111110110 : 9'b111111110;
								assign node168 = (inp[7]) ? node170 : 9'b111011110;
									assign node170 = (inp[4]) ? 9'b111010110 : 9'b111111110;
				assign node173 = (inp[13]) ? node215 : node174;
					assign node174 = (inp[11]) ? node196 : node175;
						assign node175 = (inp[7]) ? node183 : node176;
							assign node176 = (inp[9]) ? 9'b111011000 : node177;
								assign node177 = (inp[1]) ? 9'b111011000 : node178;
									assign node178 = (inp[2]) ? 9'b111111000 : 9'b111110000;
							assign node183 = (inp[4]) ? node193 : node184;
								assign node184 = (inp[0]) ? node186 : 9'b111111000;
									assign node186 = (inp[1]) ? 9'b111111000 : node187;
										assign node187 = (inp[10]) ? node189 : 9'b111110000;
											assign node189 = (inp[3]) ? 9'b111110000 : 9'b111111000;
								assign node193 = (inp[9]) ? 9'b111010000 : 9'b111110000;
						assign node196 = (inp[7]) ? node204 : node197;
							assign node197 = (inp[9]) ? 9'b111011101 : node198;
								assign node198 = (inp[1]) ? 9'b111011101 : node199;
									assign node199 = (inp[2]) ? 9'b111111101 : 9'b111110101;
							assign node204 = (inp[4]) ? node212 : node205;
								assign node205 = (inp[9]) ? 9'b111111101 : node206;
									assign node206 = (inp[1]) ? 9'b111111101 : node207;
										assign node207 = (inp[0]) ? 9'b111111101 : 9'b111110101;
								assign node212 = (inp[9]) ? 9'b111010101 : 9'b111110101;
					assign node215 = (inp[3]) ? node235 : node216;
						assign node216 = (inp[7]) ? node224 : node217;
							assign node217 = (inp[9]) ? 9'b111011101 : node218;
								assign node218 = (inp[1]) ? 9'b111011101 : node219;
									assign node219 = (inp[2]) ? 9'b111111101 : 9'b111110101;
							assign node224 = (inp[4]) ? node232 : node225;
								assign node225 = (inp[2]) ? 9'b111111101 : node226;
									assign node226 = (inp[1]) ? 9'b111111101 : node227;
										assign node227 = (inp[9]) ? 9'b111111101 : 9'b111110101;
								assign node232 = (inp[9]) ? 9'b111010101 : 9'b111110101;
						assign node235 = (inp[14]) ? node279 : node236;
							assign node236 = (inp[5]) ? node260 : node237;
								assign node237 = (inp[7]) ? node247 : node238;
									assign node238 = (inp[9]) ? 9'b110001111 : node239;
										assign node239 = (inp[1]) ? node243 : node240;
											assign node240 = (inp[2]) ? 9'b110101101 : 9'b110100101;
											assign node243 = (inp[10]) ? 9'b110001111 : 9'b110001101;
									assign node247 = (inp[4]) ? node255 : node248;
										assign node248 = (inp[1]) ? 9'b110101111 : node249;
											assign node249 = (inp[9]) ? 9'b110101111 : node250;
												assign node250 = (inp[2]) ? 9'b110101101 : 9'b110100101;
										assign node255 = (inp[9]) ? 9'b110000111 : node256;
											assign node256 = (inp[10]) ? 9'b110100111 : 9'b110100101;
								assign node260 = (inp[9]) ? node274 : node261;
									assign node261 = (inp[10]) ? node271 : node262;
										assign node262 = (inp[2]) ? 9'b110111101 : node263;
											assign node263 = (inp[1]) ? node265 : 9'b110110101;
												assign node265 = (inp[7]) ? node267 : 9'b110011101;
													assign node267 = (inp[0]) ? 9'b110111101 : 9'b110110101;
										assign node271 = (inp[7]) ? 9'b110110111 : 9'b110011111;
									assign node274 = (inp[7]) ? node276 : 9'b110011111;
										assign node276 = (inp[4]) ? 9'b110010111 : 9'b110111111;
							assign node279 = (inp[5]) ? node301 : node280;
								assign node280 = (inp[7]) ? node290 : node281;
									assign node281 = (inp[9]) ? 9'b111001111 : node282;
										assign node282 = (inp[10]) ? node286 : node283;
											assign node283 = (inp[1]) ? 9'b111001101 : 9'b111100101;
											assign node286 = (inp[11]) ? 9'b111001111 : 9'b111101111;
									assign node290 = (inp[4]) ? node298 : node291;
										assign node291 = (inp[9]) ? 9'b111101111 : node292;
											assign node292 = (inp[0]) ? 9'b111100111 : node293;
												assign node293 = (inp[10]) ? 9'b111101111 : 9'b111101101;
										assign node298 = (inp[9]) ? 9'b111000111 : 9'b111100111;
								assign node301 = (inp[9]) ? node321 : node302;
									assign node302 = (inp[10]) ? node314 : node303;
										assign node303 = (inp[7]) ? node309 : node304;
											assign node304 = (inp[1]) ? 9'b111011101 : node305;
												assign node305 = (inp[4]) ? 9'b111111101 : 9'b111110101;
											assign node309 = (inp[4]) ? 9'b111110101 : node310;
												assign node310 = (inp[2]) ? 9'b111111101 : 9'b111110101;
										assign node314 = (inp[1]) ? 9'b111011111 : node315;
											assign node315 = (inp[7]) ? 9'b111110111 : node316;
												assign node316 = (inp[2]) ? 9'b111111111 : 9'b111110111;
									assign node321 = (inp[4]) ? node325 : node322;
										assign node322 = (inp[7]) ? 9'b111111111 : 9'b111011111;
										assign node325 = (inp[7]) ? 9'b111010111 : 9'b111011111;
			assign node328 = (inp[9]) ? node374 : node329;
				assign node329 = (inp[4]) ? node353 : node330;
					assign node330 = (inp[6]) ? node340 : node331;
						assign node331 = (inp[13]) ? node335 : node332;
							assign node332 = (inp[11]) ? 9'b101111100 : 9'b101111000;
							assign node335 = (inp[3]) ? node337 : 9'b101111100;
								assign node337 = (inp[14]) ? 9'b101111110 : 9'b100111110;
						assign node340 = (inp[13]) ? node344 : node341;
							assign node341 = (inp[11]) ? 9'b101111101 : 9'b101111000;
							assign node344 = (inp[3]) ? node346 : 9'b101111101;
								assign node346 = (inp[14]) ? node350 : node347;
									assign node347 = (inp[5]) ? 9'b100111111 : 9'b100101111;
									assign node350 = (inp[5]) ? 9'b101111111 : 9'b101101111;
					assign node353 = (inp[13]) ? node359 : node354;
						assign node354 = (inp[11]) ? node356 : 9'b101010000;
							assign node356 = (inp[6]) ? 9'b101010101 : 9'b101010100;
						assign node359 = (inp[3]) ? node363 : node360;
							assign node360 = (inp[6]) ? 9'b101010101 : 9'b101010100;
							assign node363 = (inp[6]) ? node367 : node364;
								assign node364 = (inp[14]) ? 9'b101010110 : 9'b100010110;
								assign node367 = (inp[5]) ? node371 : node368;
									assign node368 = (inp[14]) ? 9'b101000111 : 9'b100000111;
									assign node371 = (inp[14]) ? 9'b101010111 : 9'b100010111;
				assign node374 = (inp[6]) ? node400 : node375;
					assign node375 = (inp[4]) ? node387 : node376;
						assign node376 = (inp[13]) ? node380 : node377;
							assign node377 = (inp[11]) ? 9'b101010100 : 9'b101010000;
							assign node380 = (inp[0]) ? node384 : node381;
								assign node381 = (inp[3]) ? 9'b111010100 : 9'b101010100;
								assign node384 = (inp[3]) ? 9'b100010110 : 9'b101010100;
						assign node387 = (inp[13]) ? node391 : node388;
							assign node388 = (inp[11]) ? 9'b111010100 : 9'b111010000;
							assign node391 = (inp[3]) ? node393 : 9'b111010100;
								assign node393 = (inp[0]) ? node397 : node394;
									assign node394 = (inp[14]) ? 9'b111010110 : 9'b110010110;
									assign node397 = (inp[14]) ? 9'b101010100 : 9'b100010100;
					assign node400 = (inp[13]) ? node408 : node401;
						assign node401 = (inp[11]) ? node405 : node402;
							assign node402 = (inp[4]) ? 9'b111010000 : 9'b101010000;
							assign node405 = (inp[4]) ? 9'b111010101 : 9'b101010101;
						assign node408 = (inp[3]) ? node412 : node409;
							assign node409 = (inp[4]) ? 9'b111010101 : 9'b101010101;
							assign node412 = (inp[0]) ? node424 : node413;
								assign node413 = (inp[4]) ? node417 : node414;
									assign node414 = (inp[5]) ? 9'b011010101 : 9'b011000101;
									assign node417 = (inp[14]) ? node421 : node418;
										assign node418 = (inp[5]) ? 9'b110010111 : 9'b110000111;
										assign node421 = (inp[5]) ? 9'b111010111 : 9'b111000111;
								assign node424 = (inp[4]) ? node428 : node425;
									assign node425 = (inp[5]) ? 9'b100010111 : 9'b100000111;
									assign node428 = (inp[14]) ? node432 : node429;
										assign node429 = (inp[5]) ? 9'b100010101 : 9'b100000101;
										assign node432 = (inp[5]) ? 9'b101010101 : 9'b101000101;

endmodule