module dtc_split05_bm26 (
	input  wire [15-1:0] inp,
	output wire [15-1:0] outp
);

	wire [15-1:0] node1;
	wire [15-1:0] node2;
	wire [15-1:0] node3;
	wire [15-1:0] node4;
	wire [15-1:0] node5;
	wire [15-1:0] node6;
	wire [15-1:0] node7;
	wire [15-1:0] node8;
	wire [15-1:0] node9;
	wire [15-1:0] node12;
	wire [15-1:0] node13;
	wire [15-1:0] node17;
	wire [15-1:0] node18;
	wire [15-1:0] node22;
	wire [15-1:0] node23;
	wire [15-1:0] node24;
	wire [15-1:0] node26;
	wire [15-1:0] node29;
	wire [15-1:0] node32;
	wire [15-1:0] node34;
	wire [15-1:0] node37;
	wire [15-1:0] node38;
	wire [15-1:0] node39;
	wire [15-1:0] node41;
	wire [15-1:0] node44;
	wire [15-1:0] node45;
	wire [15-1:0] node46;
	wire [15-1:0] node47;
	wire [15-1:0] node50;
	wire [15-1:0] node53;
	wire [15-1:0] node55;
	wire [15-1:0] node56;
	wire [15-1:0] node61;
	wire [15-1:0] node64;
	wire [15-1:0] node65;
	wire [15-1:0] node66;
	wire [15-1:0] node67;
	wire [15-1:0] node68;
	wire [15-1:0] node69;
	wire [15-1:0] node73;
	wire [15-1:0] node74;
	wire [15-1:0] node75;
	wire [15-1:0] node80;
	wire [15-1:0] node81;
	wire [15-1:0] node83;
	wire [15-1:0] node86;
	wire [15-1:0] node87;
	wire [15-1:0] node91;
	wire [15-1:0] node92;
	wire [15-1:0] node93;
	wire [15-1:0] node96;
	wire [15-1:0] node99;
	wire [15-1:0] node102;
	wire [15-1:0] node103;
	wire [15-1:0] node104;
	wire [15-1:0] node106;
	wire [15-1:0] node109;
	wire [15-1:0] node112;
	wire [15-1:0] node113;
	wire [15-1:0] node114;
	wire [15-1:0] node118;
	wire [15-1:0] node121;
	wire [15-1:0] node122;
	wire [15-1:0] node123;
	wire [15-1:0] node124;
	wire [15-1:0] node125;
	wire [15-1:0] node127;
	wire [15-1:0] node128;
	wire [15-1:0] node129;
	wire [15-1:0] node134;
	wire [15-1:0] node135;
	wire [15-1:0] node139;
	wire [15-1:0] node140;
	wire [15-1:0] node141;
	wire [15-1:0] node142;
	wire [15-1:0] node144;
	wire [15-1:0] node145;
	wire [15-1:0] node149;
	wire [15-1:0] node150;
	wire [15-1:0] node154;
	wire [15-1:0] node157;
	wire [15-1:0] node158;
	wire [15-1:0] node161;
	wire [15-1:0] node164;
	wire [15-1:0] node165;
	wire [15-1:0] node166;
	wire [15-1:0] node167;
	wire [15-1:0] node168;
	wire [15-1:0] node172;
	wire [15-1:0] node175;
	wire [15-1:0] node176;
	wire [15-1:0] node177;
	wire [15-1:0] node180;
	wire [15-1:0] node182;
	wire [15-1:0] node185;
	wire [15-1:0] node188;
	wire [15-1:0] node189;
	wire [15-1:0] node190;
	wire [15-1:0] node194;
	wire [15-1:0] node195;
	wire [15-1:0] node196;
	wire [15-1:0] node201;
	wire [15-1:0] node202;
	wire [15-1:0] node203;
	wire [15-1:0] node204;
	wire [15-1:0] node205;
	wire [15-1:0] node206;
	wire [15-1:0] node209;
	wire [15-1:0] node212;
	wire [15-1:0] node215;
	wire [15-1:0] node216;
	wire [15-1:0] node219;
	wire [15-1:0] node220;
	wire [15-1:0] node223;
	wire [15-1:0] node226;
	wire [15-1:0] node227;
	wire [15-1:0] node228;
	wire [15-1:0] node230;
	wire [15-1:0] node233;
	wire [15-1:0] node236;
	wire [15-1:0] node237;
	wire [15-1:0] node241;
	wire [15-1:0] node242;
	wire [15-1:0] node243;
	wire [15-1:0] node245;
	wire [15-1:0] node248;
	wire [15-1:0] node251;
	wire [15-1:0] node252;
	wire [15-1:0] node253;
	wire [15-1:0] node255;
	wire [15-1:0] node257;
	wire [15-1:0] node260;
	wire [15-1:0] node263;
	wire [15-1:0] node264;
	wire [15-1:0] node266;
	wire [15-1:0] node269;
	wire [15-1:0] node271;
	wire [15-1:0] node272;
	wire [15-1:0] node275;
	wire [15-1:0] node278;
	wire [15-1:0] node279;
	wire [15-1:0] node280;
	wire [15-1:0] node281;
	wire [15-1:0] node282;
	wire [15-1:0] node283;
	wire [15-1:0] node284;
	wire [15-1:0] node286;
	wire [15-1:0] node290;
	wire [15-1:0] node293;
	wire [15-1:0] node294;
	wire [15-1:0] node295;
	wire [15-1:0] node296;
	wire [15-1:0] node299;
	wire [15-1:0] node302;
	wire [15-1:0] node305;
	wire [15-1:0] node307;
	wire [15-1:0] node310;
	wire [15-1:0] node311;
	wire [15-1:0] node312;
	wire [15-1:0] node313;
	wire [15-1:0] node316;
	wire [15-1:0] node319;
	wire [15-1:0] node320;
	wire [15-1:0] node323;
	wire [15-1:0] node324;
	wire [15-1:0] node328;
	wire [15-1:0] node329;
	wire [15-1:0] node331;
	wire [15-1:0] node332;
	wire [15-1:0] node336;
	wire [15-1:0] node339;
	wire [15-1:0] node340;
	wire [15-1:0] node341;
	wire [15-1:0] node342;
	wire [15-1:0] node343;
	wire [15-1:0] node347;
	wire [15-1:0] node348;
	wire [15-1:0] node352;
	wire [15-1:0] node353;
	wire [15-1:0] node354;
	wire [15-1:0] node358;
	wire [15-1:0] node361;
	wire [15-1:0] node362;
	wire [15-1:0] node363;
	wire [15-1:0] node364;
	wire [15-1:0] node367;
	wire [15-1:0] node368;
	wire [15-1:0] node372;
	wire [15-1:0] node373;
	wire [15-1:0] node375;
	wire [15-1:0] node377;
	wire [15-1:0] node381;
	wire [15-1:0] node382;
	wire [15-1:0] node383;
	wire [15-1:0] node385;
	wire [15-1:0] node388;
	wire [15-1:0] node389;
	wire [15-1:0] node391;
	wire [15-1:0] node395;
	wire [15-1:0] node396;
	wire [15-1:0] node399;
	wire [15-1:0] node401;
	wire [15-1:0] node403;
	wire [15-1:0] node406;
	wire [15-1:0] node407;
	wire [15-1:0] node408;
	wire [15-1:0] node409;
	wire [15-1:0] node410;
	wire [15-1:0] node411;
	wire [15-1:0] node415;
	wire [15-1:0] node416;
	wire [15-1:0] node419;
	wire [15-1:0] node422;
	wire [15-1:0] node423;
	wire [15-1:0] node424;
	wire [15-1:0] node425;
	wire [15-1:0] node426;
	wire [15-1:0] node431;
	wire [15-1:0] node432;
	wire [15-1:0] node436;
	wire [15-1:0] node437;
	wire [15-1:0] node440;
	wire [15-1:0] node443;
	wire [15-1:0] node444;
	wire [15-1:0] node445;
	wire [15-1:0] node446;
	wire [15-1:0] node447;
	wire [15-1:0] node450;
	wire [15-1:0] node454;
	wire [15-1:0] node456;
	wire [15-1:0] node459;
	wire [15-1:0] node460;
	wire [15-1:0] node461;
	wire [15-1:0] node465;
	wire [15-1:0] node466;
	wire [15-1:0] node467;
	wire [15-1:0] node470;
	wire [15-1:0] node473;
	wire [15-1:0] node475;
	wire [15-1:0] node478;
	wire [15-1:0] node479;
	wire [15-1:0] node480;
	wire [15-1:0] node481;
	wire [15-1:0] node482;
	wire [15-1:0] node483;
	wire [15-1:0] node487;
	wire [15-1:0] node490;
	wire [15-1:0] node492;
	wire [15-1:0] node493;
	wire [15-1:0] node497;
	wire [15-1:0] node498;
	wire [15-1:0] node499;
	wire [15-1:0] node502;
	wire [15-1:0] node505;
	wire [15-1:0] node506;
	wire [15-1:0] node507;
	wire [15-1:0] node510;
	wire [15-1:0] node514;
	wire [15-1:0] node515;
	wire [15-1:0] node516;
	wire [15-1:0] node517;
	wire [15-1:0] node521;
	wire [15-1:0] node524;
	wire [15-1:0] node525;
	wire [15-1:0] node527;
	wire [15-1:0] node530;
	wire [15-1:0] node531;
	wire [15-1:0] node535;
	wire [15-1:0] node536;
	wire [15-1:0] node537;
	wire [15-1:0] node538;
	wire [15-1:0] node539;
	wire [15-1:0] node540;
	wire [15-1:0] node541;
	wire [15-1:0] node542;
	wire [15-1:0] node545;
	wire [15-1:0] node548;
	wire [15-1:0] node549;
	wire [15-1:0] node550;
	wire [15-1:0] node553;
	wire [15-1:0] node554;
	wire [15-1:0] node558;
	wire [15-1:0] node559;
	wire [15-1:0] node563;
	wire [15-1:0] node564;
	wire [15-1:0] node565;
	wire [15-1:0] node568;
	wire [15-1:0] node569;
	wire [15-1:0] node573;
	wire [15-1:0] node574;
	wire [15-1:0] node578;
	wire [15-1:0] node579;
	wire [15-1:0] node580;
	wire [15-1:0] node582;
	wire [15-1:0] node583;
	wire [15-1:0] node585;
	wire [15-1:0] node586;
	wire [15-1:0] node590;
	wire [15-1:0] node592;
	wire [15-1:0] node595;
	wire [15-1:0] node596;
	wire [15-1:0] node599;
	wire [15-1:0] node600;
	wire [15-1:0] node604;
	wire [15-1:0] node605;
	wire [15-1:0] node608;
	wire [15-1:0] node610;
	wire [15-1:0] node612;
	wire [15-1:0] node615;
	wire [15-1:0] node616;
	wire [15-1:0] node617;
	wire [15-1:0] node618;
	wire [15-1:0] node619;
	wire [15-1:0] node623;
	wire [15-1:0] node624;
	wire [15-1:0] node625;
	wire [15-1:0] node627;
	wire [15-1:0] node630;
	wire [15-1:0] node632;
	wire [15-1:0] node636;
	wire [15-1:0] node637;
	wire [15-1:0] node638;
	wire [15-1:0] node640;
	wire [15-1:0] node645;
	wire [15-1:0] node646;
	wire [15-1:0] node647;
	wire [15-1:0] node648;
	wire [15-1:0] node650;
	wire [15-1:0] node653;
	wire [15-1:0] node655;
	wire [15-1:0] node658;
	wire [15-1:0] node660;
	wire [15-1:0] node661;
	wire [15-1:0] node665;
	wire [15-1:0] node666;
	wire [15-1:0] node669;
	wire [15-1:0] node671;
	wire [15-1:0] node672;
	wire [15-1:0] node676;
	wire [15-1:0] node677;
	wire [15-1:0] node678;
	wire [15-1:0] node679;
	wire [15-1:0] node680;
	wire [15-1:0] node681;
	wire [15-1:0] node682;
	wire [15-1:0] node685;
	wire [15-1:0] node687;
	wire [15-1:0] node691;
	wire [15-1:0] node693;
	wire [15-1:0] node696;
	wire [15-1:0] node697;
	wire [15-1:0] node698;
	wire [15-1:0] node701;
	wire [15-1:0] node702;
	wire [15-1:0] node704;
	wire [15-1:0] node708;
	wire [15-1:0] node709;
	wire [15-1:0] node710;
	wire [15-1:0] node714;
	wire [15-1:0] node717;
	wire [15-1:0] node718;
	wire [15-1:0] node719;
	wire [15-1:0] node720;
	wire [15-1:0] node723;
	wire [15-1:0] node726;
	wire [15-1:0] node729;
	wire [15-1:0] node731;
	wire [15-1:0] node732;
	wire [15-1:0] node733;
	wire [15-1:0] node738;
	wire [15-1:0] node739;
	wire [15-1:0] node740;
	wire [15-1:0] node741;
	wire [15-1:0] node742;
	wire [15-1:0] node745;
	wire [15-1:0] node746;
	wire [15-1:0] node750;
	wire [15-1:0] node752;
	wire [15-1:0] node755;
	wire [15-1:0] node756;
	wire [15-1:0] node757;
	wire [15-1:0] node759;
	wire [15-1:0] node762;
	wire [15-1:0] node765;
	wire [15-1:0] node767;
	wire [15-1:0] node769;
	wire [15-1:0] node770;
	wire [15-1:0] node774;
	wire [15-1:0] node775;
	wire [15-1:0] node776;
	wire [15-1:0] node778;
	wire [15-1:0] node779;
	wire [15-1:0] node783;
	wire [15-1:0] node784;
	wire [15-1:0] node785;
	wire [15-1:0] node789;
	wire [15-1:0] node790;
	wire [15-1:0] node793;
	wire [15-1:0] node795;
	wire [15-1:0] node798;
	wire [15-1:0] node799;
	wire [15-1:0] node800;
	wire [15-1:0] node804;
	wire [15-1:0] node805;
	wire [15-1:0] node809;
	wire [15-1:0] node810;
	wire [15-1:0] node811;
	wire [15-1:0] node812;
	wire [15-1:0] node813;
	wire [15-1:0] node814;
	wire [15-1:0] node815;
	wire [15-1:0] node818;
	wire [15-1:0] node819;
	wire [15-1:0] node823;
	wire [15-1:0] node824;
	wire [15-1:0] node827;
	wire [15-1:0] node829;
	wire [15-1:0] node832;
	wire [15-1:0] node833;
	wire [15-1:0] node834;
	wire [15-1:0] node837;
	wire [15-1:0] node839;
	wire [15-1:0] node842;
	wire [15-1:0] node843;
	wire [15-1:0] node847;
	wire [15-1:0] node848;
	wire [15-1:0] node849;
	wire [15-1:0] node850;
	wire [15-1:0] node853;
	wire [15-1:0] node856;
	wire [15-1:0] node857;
	wire [15-1:0] node858;
	wire [15-1:0] node862;
	wire [15-1:0] node863;
	wire [15-1:0] node865;
	wire [15-1:0] node869;
	wire [15-1:0] node870;
	wire [15-1:0] node873;
	wire [15-1:0] node874;
	wire [15-1:0] node877;
	wire [15-1:0] node878;
	wire [15-1:0] node881;
	wire [15-1:0] node884;
	wire [15-1:0] node885;
	wire [15-1:0] node886;
	wire [15-1:0] node887;
	wire [15-1:0] node888;
	wire [15-1:0] node889;
	wire [15-1:0] node890;
	wire [15-1:0] node894;
	wire [15-1:0] node897;
	wire [15-1:0] node900;
	wire [15-1:0] node901;
	wire [15-1:0] node904;
	wire [15-1:0] node907;
	wire [15-1:0] node908;
	wire [15-1:0] node909;
	wire [15-1:0] node913;
	wire [15-1:0] node914;
	wire [15-1:0] node917;
	wire [15-1:0] node920;
	wire [15-1:0] node921;
	wire [15-1:0] node922;
	wire [15-1:0] node923;
	wire [15-1:0] node926;
	wire [15-1:0] node929;
	wire [15-1:0] node930;
	wire [15-1:0] node933;
	wire [15-1:0] node934;
	wire [15-1:0] node938;
	wire [15-1:0] node939;
	wire [15-1:0] node940;
	wire [15-1:0] node943;
	wire [15-1:0] node946;
	wire [15-1:0] node948;
	wire [15-1:0] node949;
	wire [15-1:0] node953;
	wire [15-1:0] node954;
	wire [15-1:0] node955;
	wire [15-1:0] node956;
	wire [15-1:0] node957;
	wire [15-1:0] node958;
	wire [15-1:0] node960;
	wire [15-1:0] node964;
	wire [15-1:0] node965;
	wire [15-1:0] node966;
	wire [15-1:0] node970;
	wire [15-1:0] node971;
	wire [15-1:0] node975;
	wire [15-1:0] node976;
	wire [15-1:0] node977;
	wire [15-1:0] node979;
	wire [15-1:0] node982;
	wire [15-1:0] node984;
	wire [15-1:0] node985;
	wire [15-1:0] node986;
	wire [15-1:0] node990;
	wire [15-1:0] node993;
	wire [15-1:0] node995;
	wire [15-1:0] node997;
	wire [15-1:0] node1000;
	wire [15-1:0] node1001;
	wire [15-1:0] node1002;
	wire [15-1:0] node1005;
	wire [15-1:0] node1007;
	wire [15-1:0] node1008;
	wire [15-1:0] node1009;
	wire [15-1:0] node1013;
	wire [15-1:0] node1016;
	wire [15-1:0] node1017;
	wire [15-1:0] node1019;
	wire [15-1:0] node1020;
	wire [15-1:0] node1023;
	wire [15-1:0] node1026;
	wire [15-1:0] node1028;
	wire [15-1:0] node1030;
	wire [15-1:0] node1033;
	wire [15-1:0] node1034;
	wire [15-1:0] node1035;
	wire [15-1:0] node1036;
	wire [15-1:0] node1039;
	wire [15-1:0] node1041;
	wire [15-1:0] node1042;
	wire [15-1:0] node1045;
	wire [15-1:0] node1048;
	wire [15-1:0] node1049;
	wire [15-1:0] node1050;
	wire [15-1:0] node1053;
	wire [15-1:0] node1054;
	wire [15-1:0] node1058;
	wire [15-1:0] node1059;
	wire [15-1:0] node1063;
	wire [15-1:0] node1064;
	wire [15-1:0] node1065;
	wire [15-1:0] node1066;
	wire [15-1:0] node1068;
	wire [15-1:0] node1071;
	wire [15-1:0] node1072;
	wire [15-1:0] node1073;
	wire [15-1:0] node1075;
	wire [15-1:0] node1080;
	wire [15-1:0] node1081;
	wire [15-1:0] node1083;
	wire [15-1:0] node1085;
	wire [15-1:0] node1089;
	wire [15-1:0] node1090;
	wire [15-1:0] node1091;
	wire [15-1:0] node1094;
	wire [15-1:0] node1097;
	wire [15-1:0] node1099;
	wire [15-1:0] node1101;
	wire [15-1:0] node1103;
	wire [15-1:0] node1106;
	wire [15-1:0] node1107;
	wire [15-1:0] node1108;
	wire [15-1:0] node1109;
	wire [15-1:0] node1110;
	wire [15-1:0] node1111;
	wire [15-1:0] node1112;
	wire [15-1:0] node1113;
	wire [15-1:0] node1115;
	wire [15-1:0] node1118;
	wire [15-1:0] node1119;
	wire [15-1:0] node1120;
	wire [15-1:0] node1122;
	wire [15-1:0] node1125;
	wire [15-1:0] node1128;
	wire [15-1:0] node1129;
	wire [15-1:0] node1133;
	wire [15-1:0] node1134;
	wire [15-1:0] node1135;
	wire [15-1:0] node1136;
	wire [15-1:0] node1139;
	wire [15-1:0] node1143;
	wire [15-1:0] node1145;
	wire [15-1:0] node1148;
	wire [15-1:0] node1149;
	wire [15-1:0] node1150;
	wire [15-1:0] node1151;
	wire [15-1:0] node1152;
	wire [15-1:0] node1155;
	wire [15-1:0] node1157;
	wire [15-1:0] node1158;
	wire [15-1:0] node1162;
	wire [15-1:0] node1164;
	wire [15-1:0] node1165;
	wire [15-1:0] node1169;
	wire [15-1:0] node1170;
	wire [15-1:0] node1173;
	wire [15-1:0] node1176;
	wire [15-1:0] node1177;
	wire [15-1:0] node1179;
	wire [15-1:0] node1181;
	wire [15-1:0] node1184;
	wire [15-1:0] node1187;
	wire [15-1:0] node1188;
	wire [15-1:0] node1189;
	wire [15-1:0] node1190;
	wire [15-1:0] node1191;
	wire [15-1:0] node1193;
	wire [15-1:0] node1196;
	wire [15-1:0] node1199;
	wire [15-1:0] node1202;
	wire [15-1:0] node1203;
	wire [15-1:0] node1204;
	wire [15-1:0] node1206;
	wire [15-1:0] node1209;
	wire [15-1:0] node1212;
	wire [15-1:0] node1214;
	wire [15-1:0] node1215;
	wire [15-1:0] node1218;
	wire [15-1:0] node1220;
	wire [15-1:0] node1223;
	wire [15-1:0] node1224;
	wire [15-1:0] node1225;
	wire [15-1:0] node1227;
	wire [15-1:0] node1230;
	wire [15-1:0] node1231;
	wire [15-1:0] node1232;
	wire [15-1:0] node1237;
	wire [15-1:0] node1238;
	wire [15-1:0] node1239;
	wire [15-1:0] node1242;
	wire [15-1:0] node1243;
	wire [15-1:0] node1245;
	wire [15-1:0] node1248;
	wire [15-1:0] node1251;
	wire [15-1:0] node1253;
	wire [15-1:0] node1256;
	wire [15-1:0] node1257;
	wire [15-1:0] node1258;
	wire [15-1:0] node1259;
	wire [15-1:0] node1260;
	wire [15-1:0] node1262;
	wire [15-1:0] node1265;
	wire [15-1:0] node1267;
	wire [15-1:0] node1270;
	wire [15-1:0] node1271;
	wire [15-1:0] node1273;
	wire [15-1:0] node1276;
	wire [15-1:0] node1279;
	wire [15-1:0] node1280;
	wire [15-1:0] node1281;
	wire [15-1:0] node1282;
	wire [15-1:0] node1285;
	wire [15-1:0] node1288;
	wire [15-1:0] node1289;
	wire [15-1:0] node1292;
	wire [15-1:0] node1293;
	wire [15-1:0] node1295;
	wire [15-1:0] node1298;
	wire [15-1:0] node1301;
	wire [15-1:0] node1303;
	wire [15-1:0] node1304;
	wire [15-1:0] node1306;
	wire [15-1:0] node1308;
	wire [15-1:0] node1311;
	wire [15-1:0] node1314;
	wire [15-1:0] node1315;
	wire [15-1:0] node1316;
	wire [15-1:0] node1317;
	wire [15-1:0] node1319;
	wire [15-1:0] node1322;
	wire [15-1:0] node1323;
	wire [15-1:0] node1327;
	wire [15-1:0] node1328;
	wire [15-1:0] node1329;
	wire [15-1:0] node1333;
	wire [15-1:0] node1335;
	wire [15-1:0] node1336;
	wire [15-1:0] node1337;
	wire [15-1:0] node1341;
	wire [15-1:0] node1342;
	wire [15-1:0] node1346;
	wire [15-1:0] node1347;
	wire [15-1:0] node1348;
	wire [15-1:0] node1351;
	wire [15-1:0] node1352;
	wire [15-1:0] node1356;
	wire [15-1:0] node1357;
	wire [15-1:0] node1358;
	wire [15-1:0] node1361;
	wire [15-1:0] node1364;
	wire [15-1:0] node1365;
	wire [15-1:0] node1366;
	wire [15-1:0] node1370;
	wire [15-1:0] node1372;
	wire [15-1:0] node1375;
	wire [15-1:0] node1376;
	wire [15-1:0] node1377;
	wire [15-1:0] node1378;
	wire [15-1:0] node1379;
	wire [15-1:0] node1380;
	wire [15-1:0] node1382;
	wire [15-1:0] node1383;
	wire [15-1:0] node1387;
	wire [15-1:0] node1388;
	wire [15-1:0] node1389;
	wire [15-1:0] node1391;
	wire [15-1:0] node1392;
	wire [15-1:0] node1397;
	wire [15-1:0] node1399;
	wire [15-1:0] node1402;
	wire [15-1:0] node1403;
	wire [15-1:0] node1404;
	wire [15-1:0] node1406;
	wire [15-1:0] node1407;
	wire [15-1:0] node1411;
	wire [15-1:0] node1412;
	wire [15-1:0] node1413;
	wire [15-1:0] node1418;
	wire [15-1:0] node1420;
	wire [15-1:0] node1423;
	wire [15-1:0] node1424;
	wire [15-1:0] node1425;
	wire [15-1:0] node1426;
	wire [15-1:0] node1427;
	wire [15-1:0] node1430;
	wire [15-1:0] node1433;
	wire [15-1:0] node1436;
	wire [15-1:0] node1438;
	wire [15-1:0] node1441;
	wire [15-1:0] node1442;
	wire [15-1:0] node1445;
	wire [15-1:0] node1447;
	wire [15-1:0] node1449;
	wire [15-1:0] node1451;
	wire [15-1:0] node1454;
	wire [15-1:0] node1455;
	wire [15-1:0] node1456;
	wire [15-1:0] node1458;
	wire [15-1:0] node1459;
	wire [15-1:0] node1461;
	wire [15-1:0] node1463;
	wire [15-1:0] node1466;
	wire [15-1:0] node1469;
	wire [15-1:0] node1470;
	wire [15-1:0] node1472;
	wire [15-1:0] node1473;
	wire [15-1:0] node1477;
	wire [15-1:0] node1478;
	wire [15-1:0] node1481;
	wire [15-1:0] node1484;
	wire [15-1:0] node1485;
	wire [15-1:0] node1486;
	wire [15-1:0] node1488;
	wire [15-1:0] node1491;
	wire [15-1:0] node1492;
	wire [15-1:0] node1493;
	wire [15-1:0] node1497;
	wire [15-1:0] node1499;
	wire [15-1:0] node1502;
	wire [15-1:0] node1503;
	wire [15-1:0] node1505;
	wire [15-1:0] node1507;
	wire [15-1:0] node1510;
	wire [15-1:0] node1512;
	wire [15-1:0] node1513;
	wire [15-1:0] node1517;
	wire [15-1:0] node1518;
	wire [15-1:0] node1519;
	wire [15-1:0] node1520;
	wire [15-1:0] node1521;
	wire [15-1:0] node1522;
	wire [15-1:0] node1524;
	wire [15-1:0] node1528;
	wire [15-1:0] node1529;
	wire [15-1:0] node1531;
	wire [15-1:0] node1534;
	wire [15-1:0] node1537;
	wire [15-1:0] node1538;
	wire [15-1:0] node1539;
	wire [15-1:0] node1542;
	wire [15-1:0] node1544;
	wire [15-1:0] node1547;
	wire [15-1:0] node1548;
	wire [15-1:0] node1551;
	wire [15-1:0] node1553;
	wire [15-1:0] node1555;
	wire [15-1:0] node1558;
	wire [15-1:0] node1559;
	wire [15-1:0] node1560;
	wire [15-1:0] node1561;
	wire [15-1:0] node1565;
	wire [15-1:0] node1566;
	wire [15-1:0] node1569;
	wire [15-1:0] node1572;
	wire [15-1:0] node1573;
	wire [15-1:0] node1574;
	wire [15-1:0] node1577;
	wire [15-1:0] node1580;
	wire [15-1:0] node1581;
	wire [15-1:0] node1582;
	wire [15-1:0] node1586;
	wire [15-1:0] node1587;
	wire [15-1:0] node1590;
	wire [15-1:0] node1593;
	wire [15-1:0] node1594;
	wire [15-1:0] node1595;
	wire [15-1:0] node1596;
	wire [15-1:0] node1597;
	wire [15-1:0] node1599;
	wire [15-1:0] node1602;
	wire [15-1:0] node1603;
	wire [15-1:0] node1605;
	wire [15-1:0] node1609;
	wire [15-1:0] node1610;
	wire [15-1:0] node1612;
	wire [15-1:0] node1615;
	wire [15-1:0] node1616;
	wire [15-1:0] node1617;
	wire [15-1:0] node1622;
	wire [15-1:0] node1623;
	wire [15-1:0] node1624;
	wire [15-1:0] node1625;
	wire [15-1:0] node1629;
	wire [15-1:0] node1631;
	wire [15-1:0] node1634;
	wire [15-1:0] node1636;
	wire [15-1:0] node1637;
	wire [15-1:0] node1638;
	wire [15-1:0] node1640;
	wire [15-1:0] node1644;
	wire [15-1:0] node1647;
	wire [15-1:0] node1648;
	wire [15-1:0] node1649;
	wire [15-1:0] node1651;
	wire [15-1:0] node1654;
	wire [15-1:0] node1655;
	wire [15-1:0] node1656;
	wire [15-1:0] node1660;
	wire [15-1:0] node1661;
	wire [15-1:0] node1665;
	wire [15-1:0] node1666;
	wire [15-1:0] node1667;
	wire [15-1:0] node1669;
	wire [15-1:0] node1672;
	wire [15-1:0] node1675;
	wire [15-1:0] node1676;
	wire [15-1:0] node1678;
	wire [15-1:0] node1681;
	wire [15-1:0] node1682;
	wire [15-1:0] node1686;
	wire [15-1:0] node1687;
	wire [15-1:0] node1688;
	wire [15-1:0] node1689;
	wire [15-1:0] node1690;
	wire [15-1:0] node1691;
	wire [15-1:0] node1692;
	wire [15-1:0] node1693;
	wire [15-1:0] node1694;
	wire [15-1:0] node1698;
	wire [15-1:0] node1699;
	wire [15-1:0] node1701;
	wire [15-1:0] node1705;
	wire [15-1:0] node1706;
	wire [15-1:0] node1709;
	wire [15-1:0] node1710;
	wire [15-1:0] node1714;
	wire [15-1:0] node1715;
	wire [15-1:0] node1716;
	wire [15-1:0] node1720;
	wire [15-1:0] node1722;
	wire [15-1:0] node1724;
	wire [15-1:0] node1725;
	wire [15-1:0] node1726;
	wire [15-1:0] node1731;
	wire [15-1:0] node1732;
	wire [15-1:0] node1733;
	wire [15-1:0] node1734;
	wire [15-1:0] node1735;
	wire [15-1:0] node1739;
	wire [15-1:0] node1740;
	wire [15-1:0] node1745;
	wire [15-1:0] node1746;
	wire [15-1:0] node1748;
	wire [15-1:0] node1750;
	wire [15-1:0] node1753;
	wire [15-1:0] node1754;
	wire [15-1:0] node1757;
	wire [15-1:0] node1760;
	wire [15-1:0] node1761;
	wire [15-1:0] node1762;
	wire [15-1:0] node1763;
	wire [15-1:0] node1764;
	wire [15-1:0] node1768;
	wire [15-1:0] node1770;
	wire [15-1:0] node1773;
	wire [15-1:0] node1774;
	wire [15-1:0] node1775;
	wire [15-1:0] node1776;
	wire [15-1:0] node1781;
	wire [15-1:0] node1783;
	wire [15-1:0] node1784;
	wire [15-1:0] node1788;
	wire [15-1:0] node1789;
	wire [15-1:0] node1790;
	wire [15-1:0] node1791;
	wire [15-1:0] node1793;
	wire [15-1:0] node1796;
	wire [15-1:0] node1798;
	wire [15-1:0] node1801;
	wire [15-1:0] node1802;
	wire [15-1:0] node1804;
	wire [15-1:0] node1805;
	wire [15-1:0] node1806;
	wire [15-1:0] node1812;
	wire [15-1:0] node1813;
	wire [15-1:0] node1816;
	wire [15-1:0] node1818;
	wire [15-1:0] node1819;
	wire [15-1:0] node1822;
	wire [15-1:0] node1825;
	wire [15-1:0] node1826;
	wire [15-1:0] node1827;
	wire [15-1:0] node1828;
	wire [15-1:0] node1829;
	wire [15-1:0] node1830;
	wire [15-1:0] node1833;
	wire [15-1:0] node1836;
	wire [15-1:0] node1837;
	wire [15-1:0] node1841;
	wire [15-1:0] node1842;
	wire [15-1:0] node1845;
	wire [15-1:0] node1848;
	wire [15-1:0] node1849;
	wire [15-1:0] node1850;
	wire [15-1:0] node1852;
	wire [15-1:0] node1853;
	wire [15-1:0] node1857;
	wire [15-1:0] node1858;
	wire [15-1:0] node1859;
	wire [15-1:0] node1864;
	wire [15-1:0] node1865;
	wire [15-1:0] node1867;
	wire [15-1:0] node1869;
	wire [15-1:0] node1872;
	wire [15-1:0] node1873;
	wire [15-1:0] node1875;
	wire [15-1:0] node1878;
	wire [15-1:0] node1881;
	wire [15-1:0] node1882;
	wire [15-1:0] node1883;
	wire [15-1:0] node1884;
	wire [15-1:0] node1886;
	wire [15-1:0] node1889;
	wire [15-1:0] node1890;
	wire [15-1:0] node1892;
	wire [15-1:0] node1893;
	wire [15-1:0] node1895;
	wire [15-1:0] node1900;
	wire [15-1:0] node1901;
	wire [15-1:0] node1904;
	wire [15-1:0] node1905;
	wire [15-1:0] node1909;
	wire [15-1:0] node1910;
	wire [15-1:0] node1911;
	wire [15-1:0] node1912;
	wire [15-1:0] node1915;
	wire [15-1:0] node1918;
	wire [15-1:0] node1919;
	wire [15-1:0] node1922;
	wire [15-1:0] node1923;
	wire [15-1:0] node1927;
	wire [15-1:0] node1928;
	wire [15-1:0] node1929;
	wire [15-1:0] node1931;
	wire [15-1:0] node1934;
	wire [15-1:0] node1937;
	wire [15-1:0] node1938;
	wire [15-1:0] node1939;
	wire [15-1:0] node1941;
	wire [15-1:0] node1945;
	wire [15-1:0] node1947;
	wire [15-1:0] node1950;
	wire [15-1:0] node1951;
	wire [15-1:0] node1952;
	wire [15-1:0] node1953;
	wire [15-1:0] node1954;
	wire [15-1:0] node1955;
	wire [15-1:0] node1956;
	wire [15-1:0] node1958;
	wire [15-1:0] node1961;
	wire [15-1:0] node1964;
	wire [15-1:0] node1965;
	wire [15-1:0] node1967;
	wire [15-1:0] node1970;
	wire [15-1:0] node1971;
	wire [15-1:0] node1975;
	wire [15-1:0] node1976;
	wire [15-1:0] node1978;
	wire [15-1:0] node1981;
	wire [15-1:0] node1984;
	wire [15-1:0] node1985;
	wire [15-1:0] node1986;
	wire [15-1:0] node1987;
	wire [15-1:0] node1990;
	wire [15-1:0] node1992;
	wire [15-1:0] node1995;
	wire [15-1:0] node1997;
	wire [15-1:0] node1998;
	wire [15-1:0] node2001;
	wire [15-1:0] node2002;
	wire [15-1:0] node2006;
	wire [15-1:0] node2007;
	wire [15-1:0] node2008;
	wire [15-1:0] node2011;
	wire [15-1:0] node2012;
	wire [15-1:0] node2016;
	wire [15-1:0] node2017;
	wire [15-1:0] node2021;
	wire [15-1:0] node2022;
	wire [15-1:0] node2023;
	wire [15-1:0] node2025;
	wire [15-1:0] node2028;
	wire [15-1:0] node2029;
	wire [15-1:0] node2030;
	wire [15-1:0] node2032;
	wire [15-1:0] node2035;
	wire [15-1:0] node2036;
	wire [15-1:0] node2037;
	wire [15-1:0] node2042;
	wire [15-1:0] node2043;
	wire [15-1:0] node2044;
	wire [15-1:0] node2046;
	wire [15-1:0] node2049;
	wire [15-1:0] node2052;
	wire [15-1:0] node2055;
	wire [15-1:0] node2056;
	wire [15-1:0] node2057;
	wire [15-1:0] node2060;
	wire [15-1:0] node2061;
	wire [15-1:0] node2064;
	wire [15-1:0] node2066;
	wire [15-1:0] node2069;
	wire [15-1:0] node2071;
	wire [15-1:0] node2072;
	wire [15-1:0] node2074;
	wire [15-1:0] node2078;
	wire [15-1:0] node2079;
	wire [15-1:0] node2080;
	wire [15-1:0] node2081;
	wire [15-1:0] node2082;
	wire [15-1:0] node2083;
	wire [15-1:0] node2087;
	wire [15-1:0] node2088;
	wire [15-1:0] node2089;
	wire [15-1:0] node2093;
	wire [15-1:0] node2095;
	wire [15-1:0] node2098;
	wire [15-1:0] node2099;
	wire [15-1:0] node2100;
	wire [15-1:0] node2104;
	wire [15-1:0] node2107;
	wire [15-1:0] node2108;
	wire [15-1:0] node2109;
	wire [15-1:0] node2110;
	wire [15-1:0] node2111;
	wire [15-1:0] node2113;
	wire [15-1:0] node2117;
	wire [15-1:0] node2120;
	wire [15-1:0] node2121;
	wire [15-1:0] node2124;
	wire [15-1:0] node2126;
	wire [15-1:0] node2127;
	wire [15-1:0] node2131;
	wire [15-1:0] node2132;
	wire [15-1:0] node2134;
	wire [15-1:0] node2137;
	wire [15-1:0] node2138;
	wire [15-1:0] node2140;
	wire [15-1:0] node2143;
	wire [15-1:0] node2145;
	wire [15-1:0] node2148;
	wire [15-1:0] node2149;
	wire [15-1:0] node2150;
	wire [15-1:0] node2151;
	wire [15-1:0] node2152;
	wire [15-1:0] node2154;
	wire [15-1:0] node2157;
	wire [15-1:0] node2158;
	wire [15-1:0] node2161;
	wire [15-1:0] node2165;
	wire [15-1:0] node2166;
	wire [15-1:0] node2167;
	wire [15-1:0] node2170;
	wire [15-1:0] node2171;
	wire [15-1:0] node2175;
	wire [15-1:0] node2176;
	wire [15-1:0] node2180;
	wire [15-1:0] node2181;
	wire [15-1:0] node2182;
	wire [15-1:0] node2183;
	wire [15-1:0] node2186;
	wire [15-1:0] node2188;
	wire [15-1:0] node2189;
	wire [15-1:0] node2193;
	wire [15-1:0] node2194;
	wire [15-1:0] node2196;
	wire [15-1:0] node2199;
	wire [15-1:0] node2201;
	wire [15-1:0] node2204;
	wire [15-1:0] node2205;
	wire [15-1:0] node2207;
	wire [15-1:0] node2208;
	wire [15-1:0] node2211;
	wire [15-1:0] node2214;
	wire [15-1:0] node2215;
	wire [15-1:0] node2216;
	wire [15-1:0] node2220;

	assign outp = (inp[4]) ? node1106 : node1;
		assign node1 = (inp[2]) ? node535 : node2;
			assign node2 = (inp[11]) ? node278 : node3;
				assign node3 = (inp[9]) ? node121 : node4;
					assign node4 = (inp[1]) ? node64 : node5;
						assign node5 = (inp[3]) ? node37 : node6;
							assign node6 = (inp[7]) ? node22 : node7;
								assign node7 = (inp[13]) ? node17 : node8;
									assign node8 = (inp[10]) ? node12 : node9;
										assign node9 = (inp[8]) ? 15'b000011111111111 : 15'b000111111111111;
										assign node12 = (inp[0]) ? 15'b000011111111111 : node13;
											assign node13 = (inp[12]) ? 15'b000011111111111 : 15'b000111111111111;
									assign node17 = (inp[10]) ? 15'b000001111111111 : node18;
										assign node18 = (inp[12]) ? 15'b000011111111111 : 15'b000001111111111;
								assign node22 = (inp[6]) ? node32 : node23;
									assign node23 = (inp[12]) ? node29 : node24;
										assign node24 = (inp[14]) ? node26 : 15'b000111111111111;
											assign node26 = (inp[10]) ? 15'b000011111111111 : 15'b000111111111111;
										assign node29 = (inp[5]) ? 15'b000001111111111 : 15'b000011111111111;
									assign node32 = (inp[14]) ? node34 : 15'b000001111111111;
										assign node34 = (inp[12]) ? 15'b000000011111111 : 15'b000001111111111;
							assign node37 = (inp[10]) ? node61 : node38;
								assign node38 = (inp[5]) ? node44 : node39;
									assign node39 = (inp[0]) ? node41 : 15'b000111111111111;
										assign node41 = (inp[12]) ? 15'b000001111111111 : 15'b000011111111111;
									assign node44 = (inp[7]) ? 15'b000000011111111 : node45;
										assign node45 = (inp[0]) ? node53 : node46;
											assign node46 = (inp[13]) ? node50 : node47;
												assign node47 = (inp[8]) ? 15'b000011111111111 : 15'b000111111111111;
												assign node50 = (inp[8]) ? 15'b000001111111111 : 15'b000011111111111;
											assign node53 = (inp[14]) ? node55 : 15'b000011111111111;
												assign node55 = (inp[13]) ? 15'b000000111111111 : node56;
													assign node56 = (inp[8]) ? 15'b000000111111111 : 15'b000001111111111;
								assign node61 = (inp[12]) ? 15'b000000011111111 : 15'b000000111111111;
						assign node64 = (inp[0]) ? node102 : node65;
							assign node65 = (inp[7]) ? node91 : node66;
								assign node66 = (inp[8]) ? node80 : node67;
									assign node67 = (inp[6]) ? node73 : node68;
										assign node68 = (inp[3]) ? 15'b000001111111111 : node69;
											assign node69 = (inp[13]) ? 15'b000011111111111 : 15'b000111111111111;
										assign node73 = (inp[12]) ? 15'b000001111111111 : node74;
											assign node74 = (inp[13]) ? 15'b000011111111111 : node75;
												assign node75 = (inp[5]) ? 15'b000001111111111 : 15'b000011111111111;
									assign node80 = (inp[13]) ? node86 : node81;
										assign node81 = (inp[5]) ? node83 : 15'b000011111111111;
											assign node83 = (inp[6]) ? 15'b000000111111111 : 15'b000001111111111;
										assign node86 = (inp[12]) ? 15'b000000011111111 : node87;
											assign node87 = (inp[6]) ? 15'b000000111111111 : 15'b000001111111111;
								assign node91 = (inp[3]) ? node99 : node92;
									assign node92 = (inp[6]) ? node96 : node93;
										assign node93 = (inp[12]) ? 15'b000001111111111 : 15'b000111111111111;
										assign node96 = (inp[14]) ? 15'b000000111111111 : 15'b000001111111111;
									assign node99 = (inp[12]) ? 15'b000000011111111 : 15'b000000111111111;
							assign node102 = (inp[3]) ? node112 : node103;
								assign node103 = (inp[14]) ? node109 : node104;
									assign node104 = (inp[6]) ? node106 : 15'b000001111111111;
										assign node106 = (inp[5]) ? 15'b000000111111111 : 15'b000001111111111;
									assign node109 = (inp[7]) ? 15'b000000011111111 : 15'b000000111111111;
								assign node112 = (inp[8]) ? node118 : node113;
									assign node113 = (inp[10]) ? 15'b000000001111111 : node114;
										assign node114 = (inp[6]) ? 15'b000000111111111 : 15'b000001111111111;
									assign node118 = (inp[10]) ? 15'b000000011111111 : 15'b000000001111111;
					assign node121 = (inp[14]) ? node201 : node122;
						assign node122 = (inp[5]) ? node164 : node123;
							assign node123 = (inp[8]) ? node139 : node124;
								assign node124 = (inp[12]) ? node134 : node125;
									assign node125 = (inp[0]) ? node127 : 15'b001111111111111;
										assign node127 = (inp[6]) ? 15'b000001111111111 : node128;
											assign node128 = (inp[3]) ? 15'b000011111111111 : node129;
												assign node129 = (inp[10]) ? 15'b000011111111111 : 15'b000111111111111;
									assign node134 = (inp[3]) ? 15'b000000111111111 : node135;
										assign node135 = (inp[0]) ? 15'b000001111111111 : 15'b000011111111111;
								assign node139 = (inp[6]) ? node157 : node140;
									assign node140 = (inp[13]) ? node154 : node141;
										assign node141 = (inp[3]) ? node149 : node142;
											assign node142 = (inp[12]) ? node144 : 15'b000011111111111;
												assign node144 = (inp[1]) ? 15'b000001111111111 : node145;
													assign node145 = (inp[0]) ? 15'b000001111111111 : 15'b000011111111111;
											assign node149 = (inp[0]) ? 15'b000001111111111 : node150;
												assign node150 = (inp[12]) ? 15'b000001111111111 : 15'b000011111111111;
										assign node154 = (inp[7]) ? 15'b000000111111111 : 15'b000001111111111;
									assign node157 = (inp[12]) ? node161 : node158;
										assign node158 = (inp[0]) ? 15'b000000111111111 : 15'b000001111111111;
										assign node161 = (inp[0]) ? 15'b000000001111111 : 15'b000000011111111;
							assign node164 = (inp[8]) ? node188 : node165;
								assign node165 = (inp[1]) ? node175 : node166;
									assign node166 = (inp[12]) ? node172 : node167;
										assign node167 = (inp[13]) ? 15'b000001111111111 : node168;
											assign node168 = (inp[3]) ? 15'b000011111111111 : 15'b000111111111111;
										assign node172 = (inp[0]) ? 15'b000000111111111 : 15'b000001111111111;
									assign node175 = (inp[13]) ? node185 : node176;
										assign node176 = (inp[12]) ? node180 : node177;
											assign node177 = (inp[10]) ? 15'b000000111111111 : 15'b000001111111111;
											assign node180 = (inp[6]) ? node182 : 15'b000000111111111;
												assign node182 = (inp[7]) ? 15'b000000001111111 : 15'b000000111111111;
										assign node185 = (inp[6]) ? 15'b000000001111111 : 15'b000000011111111;
								assign node188 = (inp[6]) ? node194 : node189;
									assign node189 = (inp[0]) ? 15'b000000011111111 : node190;
										assign node190 = (inp[10]) ? 15'b000000111111111 : 15'b000001111111111;
									assign node194 = (inp[0]) ? 15'b000000001111111 : node195;
										assign node195 = (inp[1]) ? 15'b000000001111111 : node196;
											assign node196 = (inp[7]) ? 15'b000000111111111 : 15'b000000011111111;
						assign node201 = (inp[10]) ? node241 : node202;
							assign node202 = (inp[1]) ? node226 : node203;
								assign node203 = (inp[6]) ? node215 : node204;
									assign node204 = (inp[5]) ? node212 : node205;
										assign node205 = (inp[12]) ? node209 : node206;
											assign node206 = (inp[13]) ? 15'b000111111111111 : 15'b000011111111111;
											assign node209 = (inp[8]) ? 15'b000000111111111 : 15'b000001111111111;
										assign node212 = (inp[13]) ? 15'b000000111111111 : 15'b000001111111111;
									assign node215 = (inp[13]) ? node219 : node216;
										assign node216 = (inp[7]) ? 15'b000000111111111 : 15'b000001111111111;
										assign node219 = (inp[8]) ? node223 : node220;
											assign node220 = (inp[7]) ? 15'b000000011111111 : 15'b000000111111111;
											assign node223 = (inp[5]) ? 15'b000000000111111 : 15'b000000001111111;
								assign node226 = (inp[13]) ? node236 : node227;
									assign node227 = (inp[5]) ? node233 : node228;
										assign node228 = (inp[7]) ? node230 : 15'b000011111111111;
											assign node230 = (inp[6]) ? 15'b000000111111111 : 15'b000000011111111;
										assign node233 = (inp[3]) ? 15'b000000001111111 : 15'b000000011111111;
									assign node236 = (inp[7]) ? 15'b000000001111111 : node237;
										assign node237 = (inp[8]) ? 15'b000000000111111 : 15'b000000011111111;
							assign node241 = (inp[12]) ? node251 : node242;
								assign node242 = (inp[3]) ? node248 : node243;
									assign node243 = (inp[0]) ? node245 : 15'b000000111111111;
										assign node245 = (inp[6]) ? 15'b000000000111111 : 15'b000001111111111;
									assign node248 = (inp[8]) ? 15'b000000001111111 : 15'b000000000111111;
								assign node251 = (inp[13]) ? node263 : node252;
									assign node252 = (inp[0]) ? node260 : node253;
										assign node253 = (inp[1]) ? node255 : 15'b000000001111111;
											assign node255 = (inp[5]) ? node257 : 15'b000000001111111;
												assign node257 = (inp[7]) ? 15'b000000000011111 : 15'b000000000111111;
										assign node260 = (inp[8]) ? 15'b000000001111111 : 15'b000000011111111;
									assign node263 = (inp[0]) ? node269 : node264;
										assign node264 = (inp[5]) ? node266 : 15'b000000011111111;
											assign node266 = (inp[7]) ? 15'b000000000111111 : 15'b000000001111111;
										assign node269 = (inp[6]) ? node271 : 15'b000000000111111;
											assign node271 = (inp[1]) ? node275 : node272;
												assign node272 = (inp[3]) ? 15'b000000000011111 : 15'b000000000111111;
												assign node275 = (inp[7]) ? 15'b000000000001111 : 15'b000000000011111;
				assign node278 = (inp[8]) ? node406 : node279;
					assign node279 = (inp[10]) ? node339 : node280;
						assign node280 = (inp[13]) ? node310 : node281;
							assign node281 = (inp[0]) ? node293 : node282;
								assign node282 = (inp[3]) ? node290 : node283;
									assign node283 = (inp[6]) ? 15'b000001111111111 : node284;
										assign node284 = (inp[14]) ? node286 : 15'b000011111111111;
											assign node286 = (inp[7]) ? 15'b000001111111111 : 15'b000011111111111;
									assign node290 = (inp[6]) ? 15'b000001111111111 : 15'b000000111111111;
								assign node293 = (inp[9]) ? node305 : node294;
									assign node294 = (inp[7]) ? node302 : node295;
										assign node295 = (inp[3]) ? node299 : node296;
											assign node296 = (inp[12]) ? 15'b000001111111111 : 15'b000111111111111;
											assign node299 = (inp[6]) ? 15'b000000111111111 : 15'b000001111111111;
										assign node302 = (inp[14]) ? 15'b000000111111111 : 15'b000001111111111;
									assign node305 = (inp[1]) ? node307 : 15'b000000111111111;
										assign node307 = (inp[3]) ? 15'b000000011111111 : 15'b000000001111111;
							assign node310 = (inp[1]) ? node328 : node311;
								assign node311 = (inp[0]) ? node319 : node312;
									assign node312 = (inp[3]) ? node316 : node313;
										assign node313 = (inp[6]) ? 15'b000011111111111 : 15'b000111111111111;
										assign node316 = (inp[7]) ? 15'b000000111111111 : 15'b000001111111111;
									assign node319 = (inp[6]) ? node323 : node320;
										assign node320 = (inp[7]) ? 15'b000001111111111 : 15'b000000111111111;
										assign node323 = (inp[9]) ? 15'b000000111111111 : node324;
											assign node324 = (inp[3]) ? 15'b000000011111111 : 15'b000000111111111;
								assign node328 = (inp[3]) ? node336 : node329;
									assign node329 = (inp[7]) ? node331 : 15'b000000111111111;
										assign node331 = (inp[9]) ? 15'b000000001111111 : node332;
											assign node332 = (inp[5]) ? 15'b000000011111111 : 15'b000000111111111;
									assign node336 = (inp[9]) ? 15'b000000011111111 : 15'b000000001111111;
						assign node339 = (inp[0]) ? node361 : node340;
							assign node340 = (inp[9]) ? node352 : node341;
								assign node341 = (inp[12]) ? node347 : node342;
									assign node342 = (inp[7]) ? 15'b000001111111111 : node343;
										assign node343 = (inp[6]) ? 15'b000001111111111 : 15'b000011111111111;
									assign node347 = (inp[7]) ? 15'b000000011111111 : node348;
										assign node348 = (inp[5]) ? 15'b000000111111111 : 15'b000001111111111;
								assign node352 = (inp[12]) ? node358 : node353;
									assign node353 = (inp[3]) ? 15'b000000001111111 : node354;
										assign node354 = (inp[14]) ? 15'b000000111111111 : 15'b000001111111111;
									assign node358 = (inp[14]) ? 15'b000000001111111 : 15'b000000111111111;
							assign node361 = (inp[6]) ? node381 : node362;
								assign node362 = (inp[5]) ? node372 : node363;
									assign node363 = (inp[3]) ? node367 : node364;
										assign node364 = (inp[12]) ? 15'b000000111111111 : 15'b000001111111111;
										assign node367 = (inp[12]) ? 15'b000000011111111 : node368;
											assign node368 = (inp[1]) ? 15'b000000011111111 : 15'b000000111111111;
									assign node372 = (inp[12]) ? 15'b000000000111111 : node373;
										assign node373 = (inp[13]) ? node375 : 15'b000000011111111;
											assign node375 = (inp[3]) ? node377 : 15'b000000011111111;
												assign node377 = (inp[9]) ? 15'b000000000111111 : 15'b000000001111111;
								assign node381 = (inp[3]) ? node395 : node382;
									assign node382 = (inp[9]) ? node388 : node383;
										assign node383 = (inp[13]) ? node385 : 15'b000000111111111;
											assign node385 = (inp[5]) ? 15'b000000001111111 : 15'b000000011111111;
										assign node388 = (inp[14]) ? 15'b000000000111111 : node389;
											assign node389 = (inp[13]) ? node391 : 15'b000000011111111;
												assign node391 = (inp[7]) ? 15'b000000000111111 : 15'b000000001111111;
									assign node395 = (inp[13]) ? node399 : node396;
										assign node396 = (inp[14]) ? 15'b000000000111111 : 15'b000000001111111;
										assign node399 = (inp[9]) ? node401 : 15'b000000000011111;
											assign node401 = (inp[1]) ? node403 : 15'b000000000111111;
												assign node403 = (inp[7]) ? 15'b000000000011111 : 15'b000000000111111;
					assign node406 = (inp[7]) ? node478 : node407;
						assign node407 = (inp[14]) ? node443 : node408;
							assign node408 = (inp[3]) ? node422 : node409;
								assign node409 = (inp[5]) ? node415 : node410;
									assign node410 = (inp[1]) ? 15'b000001111111111 : node411;
										assign node411 = (inp[9]) ? 15'b000011111111111 : 15'b000111111111111;
									assign node415 = (inp[1]) ? node419 : node416;
										assign node416 = (inp[0]) ? 15'b000001111111111 : 15'b000000111111111;
										assign node419 = (inp[13]) ? 15'b000000001111111 : 15'b000000011111111;
								assign node422 = (inp[10]) ? node436 : node423;
									assign node423 = (inp[9]) ? node431 : node424;
										assign node424 = (inp[12]) ? 15'b000000011111111 : node425;
											assign node425 = (inp[13]) ? 15'b000000111111111 : node426;
												assign node426 = (inp[0]) ? 15'b000000111111111 : 15'b000001111111111;
										assign node431 = (inp[5]) ? 15'b000000011111111 : node432;
											assign node432 = (inp[6]) ? 15'b000000011111111 : 15'b000000111111111;
									assign node436 = (inp[6]) ? node440 : node437;
										assign node437 = (inp[9]) ? 15'b000000111111111 : 15'b000000011111111;
										assign node440 = (inp[5]) ? 15'b000000001111111 : 15'b000000011111111;
							assign node443 = (inp[9]) ? node459 : node444;
								assign node444 = (inp[3]) ? node454 : node445;
									assign node445 = (inp[5]) ? 15'b000000001111111 : node446;
										assign node446 = (inp[6]) ? node450 : node447;
											assign node447 = (inp[13]) ? 15'b000000111111111 : 15'b000001111111111;
											assign node450 = (inp[10]) ? 15'b000000011111111 : 15'b000000111111111;
									assign node454 = (inp[6]) ? node456 : 15'b000000011111111;
										assign node456 = (inp[12]) ? 15'b000000011111111 : 15'b000000001111111;
								assign node459 = (inp[1]) ? node465 : node460;
									assign node460 = (inp[3]) ? 15'b000000001111111 : node461;
										assign node461 = (inp[12]) ? 15'b000000011111111 : 15'b000000001111111;
									assign node465 = (inp[10]) ? node473 : node466;
										assign node466 = (inp[5]) ? node470 : node467;
											assign node467 = (inp[13]) ? 15'b000000001111111 : 15'b000000111111111;
											assign node470 = (inp[3]) ? 15'b000000000011111 : 15'b000000001111111;
										assign node473 = (inp[3]) ? node475 : 15'b000000000111111;
											assign node475 = (inp[12]) ? 15'b000000000001111 : 15'b000000000111111;
						assign node478 = (inp[1]) ? node514 : node479;
							assign node479 = (inp[3]) ? node497 : node480;
								assign node480 = (inp[13]) ? node490 : node481;
									assign node481 = (inp[0]) ? node487 : node482;
										assign node482 = (inp[14]) ? 15'b000000111111111 : node483;
											assign node483 = (inp[12]) ? 15'b000011111111111 : 15'b000000111111111;
										assign node487 = (inp[5]) ? 15'b000000011111111 : 15'b000000111111111;
									assign node490 = (inp[12]) ? node492 : 15'b000000111111111;
										assign node492 = (inp[9]) ? 15'b000000001111111 : node493;
											assign node493 = (inp[14]) ? 15'b000000000111111 : 15'b000000001111111;
								assign node497 = (inp[10]) ? node505 : node498;
									assign node498 = (inp[13]) ? node502 : node499;
										assign node499 = (inp[14]) ? 15'b000000111111111 : 15'b000000011111111;
										assign node502 = (inp[5]) ? 15'b000000001111111 : 15'b000000000111111;
									assign node505 = (inp[0]) ? 15'b000000000111111 : node506;
										assign node506 = (inp[5]) ? node510 : node507;
											assign node507 = (inp[12]) ? 15'b000000011111111 : 15'b000000001111111;
											assign node510 = (inp[9]) ? 15'b000000000011111 : 15'b000000000111111;
							assign node514 = (inp[10]) ? node524 : node515;
								assign node515 = (inp[5]) ? node521 : node516;
									assign node516 = (inp[14]) ? 15'b000000001111111 : node517;
										assign node517 = (inp[12]) ? 15'b000000001111111 : 15'b000000111111111;
									assign node521 = (inp[6]) ? 15'b000000000011111 : 15'b000000001111111;
								assign node524 = (inp[13]) ? node530 : node525;
									assign node525 = (inp[5]) ? node527 : 15'b000000001111111;
										assign node527 = (inp[12]) ? 15'b000000000001111 : 15'b000000000111111;
									assign node530 = (inp[9]) ? 15'b000000000011111 : node531;
										assign node531 = (inp[5]) ? 15'b000000000011111 : 15'b000000001111111;
			assign node535 = (inp[5]) ? node809 : node536;
				assign node536 = (inp[0]) ? node676 : node537;
					assign node537 = (inp[3]) ? node615 : node538;
						assign node538 = (inp[14]) ? node578 : node539;
							assign node539 = (inp[10]) ? node563 : node540;
								assign node540 = (inp[8]) ? node548 : node541;
									assign node541 = (inp[1]) ? node545 : node542;
										assign node542 = (inp[7]) ? 15'b000011111111111 : 15'b000111111111111;
										assign node545 = (inp[12]) ? 15'b000001111111111 : 15'b000011111111111;
									assign node548 = (inp[13]) ? node558 : node549;
										assign node549 = (inp[12]) ? node553 : node550;
											assign node550 = (inp[1]) ? 15'b000011111111111 : 15'b001111111111111;
											assign node553 = (inp[7]) ? 15'b000011111111111 : node554;
												assign node554 = (inp[6]) ? 15'b000001111111111 : 15'b000000111111111;
										assign node558 = (inp[9]) ? 15'b000000111111111 : node559;
											assign node559 = (inp[6]) ? 15'b000000011111111 : 15'b000001111111111;
								assign node563 = (inp[7]) ? node573 : node564;
									assign node564 = (inp[11]) ? node568 : node565;
										assign node565 = (inp[6]) ? 15'b000001111111111 : 15'b000011111111111;
										assign node568 = (inp[1]) ? 15'b000000111111111 : node569;
											assign node569 = (inp[12]) ? 15'b000000111111111 : 15'b000001111111111;
									assign node573 = (inp[12]) ? 15'b000000011111111 : node574;
										assign node574 = (inp[11]) ? 15'b000000111111111 : 15'b000001111111111;
							assign node578 = (inp[1]) ? node604 : node579;
								assign node579 = (inp[12]) ? node595 : node580;
									assign node580 = (inp[7]) ? node582 : 15'b000001111111111;
										assign node582 = (inp[8]) ? node590 : node583;
											assign node583 = (inp[10]) ? node585 : 15'b000001111111111;
												assign node585 = (inp[6]) ? 15'b000000011111111 : node586;
													assign node586 = (inp[11]) ? 15'b000000111111111 : 15'b000001111111111;
											assign node590 = (inp[6]) ? node592 : 15'b000000111111111;
												assign node592 = (inp[11]) ? 15'b000000011111111 : 15'b000000111111111;
									assign node595 = (inp[9]) ? node599 : node596;
										assign node596 = (inp[10]) ? 15'b000000111111111 : 15'b000001111111111;
										assign node599 = (inp[7]) ? 15'b000000001111111 : node600;
											assign node600 = (inp[8]) ? 15'b000000011111111 : 15'b000000111111111;
								assign node604 = (inp[13]) ? node608 : node605;
									assign node605 = (inp[7]) ? 15'b000000111111111 : 15'b000000011111111;
									assign node608 = (inp[12]) ? node610 : 15'b000000001111111;
										assign node610 = (inp[8]) ? node612 : 15'b000000111111111;
											assign node612 = (inp[6]) ? 15'b000000000111111 : 15'b000000000011111;
						assign node615 = (inp[9]) ? node645 : node616;
							assign node616 = (inp[12]) ? node636 : node617;
								assign node617 = (inp[8]) ? node623 : node618;
									assign node618 = (inp[1]) ? 15'b000000111111111 : node619;
										assign node619 = (inp[14]) ? 15'b000001111111111 : 15'b000011111111111;
									assign node623 = (inp[14]) ? 15'b000000011111111 : node624;
										assign node624 = (inp[13]) ? node630 : node625;
											assign node625 = (inp[7]) ? node627 : 15'b000001111111111;
												assign node627 = (inp[6]) ? 15'b000000111111111 : 15'b000001111111111;
											assign node630 = (inp[6]) ? node632 : 15'b000000111111111;
												assign node632 = (inp[7]) ? 15'b000000001111111 : 15'b000000011111111;
								assign node636 = (inp[1]) ? 15'b000000001111111 : node637;
									assign node637 = (inp[14]) ? 15'b000000011111111 : node638;
										assign node638 = (inp[8]) ? node640 : 15'b000000111111111;
											assign node640 = (inp[13]) ? 15'b000000001111111 : 15'b000000011111111;
							assign node645 = (inp[11]) ? node665 : node646;
								assign node646 = (inp[7]) ? node658 : node647;
									assign node647 = (inp[14]) ? node653 : node648;
										assign node648 = (inp[6]) ? node650 : 15'b000001111111111;
											assign node650 = (inp[10]) ? 15'b000000011111111 : 15'b000001111111111;
										assign node653 = (inp[13]) ? node655 : 15'b000000011111111;
											assign node655 = (inp[8]) ? 15'b000000000111111 : 15'b000000011111111;
									assign node658 = (inp[1]) ? node660 : 15'b000000111111111;
										assign node660 = (inp[13]) ? 15'b000000001111111 : node661;
											assign node661 = (inp[14]) ? 15'b000000000111111 : 15'b000000001111111;
								assign node665 = (inp[12]) ? node669 : node666;
									assign node666 = (inp[1]) ? 15'b000000001111111 : 15'b000001111111111;
									assign node669 = (inp[13]) ? node671 : 15'b000000001111111;
										assign node671 = (inp[14]) ? 15'b000000000011111 : node672;
											assign node672 = (inp[10]) ? 15'b000000000111111 : 15'b000000001111111;
					assign node676 = (inp[13]) ? node738 : node677;
						assign node677 = (inp[7]) ? node717 : node678;
							assign node678 = (inp[9]) ? node696 : node679;
								assign node679 = (inp[11]) ? node691 : node680;
									assign node680 = (inp[6]) ? 15'b000111111111111 : node681;
										assign node681 = (inp[8]) ? node685 : node682;
											assign node682 = (inp[1]) ? 15'b000001111111111 : 15'b000011111111111;
											assign node685 = (inp[3]) ? node687 : 15'b000001111111111;
												assign node687 = (inp[12]) ? 15'b000000011111111 : 15'b000000111111111;
									assign node691 = (inp[3]) ? node693 : 15'b000000001111111;
										assign node693 = (inp[10]) ? 15'b000000111111111 : 15'b000000011111111;
								assign node696 = (inp[10]) ? node708 : node697;
									assign node697 = (inp[1]) ? node701 : node698;
										assign node698 = (inp[14]) ? 15'b000000111111111 : 15'b000011111111111;
										assign node701 = (inp[8]) ? 15'b000000011111111 : node702;
											assign node702 = (inp[11]) ? node704 : 15'b000000111111111;
												assign node704 = (inp[3]) ? 15'b000000011111111 : 15'b000000111111111;
									assign node708 = (inp[6]) ? node714 : node709;
										assign node709 = (inp[14]) ? 15'b000000011111111 : node710;
											assign node710 = (inp[3]) ? 15'b000000011111111 : 15'b000000111111111;
										assign node714 = (inp[12]) ? 15'b000000011111111 : 15'b000000001111111;
							assign node717 = (inp[14]) ? node729 : node718;
								assign node718 = (inp[10]) ? node726 : node719;
									assign node719 = (inp[1]) ? node723 : node720;
										assign node720 = (inp[6]) ? 15'b000000011111111 : 15'b000000111111111;
										assign node723 = (inp[3]) ? 15'b000000011111111 : 15'b000000111111111;
									assign node726 = (inp[6]) ? 15'b000000001111111 : 15'b000000011111111;
								assign node729 = (inp[11]) ? node731 : 15'b000000001111111;
									assign node731 = (inp[10]) ? 15'b000000000111111 : node732;
										assign node732 = (inp[8]) ? 15'b000000000111111 : node733;
											assign node733 = (inp[12]) ? 15'b000000001111111 : 15'b000000011111111;
						assign node738 = (inp[12]) ? node774 : node739;
							assign node739 = (inp[1]) ? node755 : node740;
								assign node740 = (inp[10]) ? node750 : node741;
									assign node741 = (inp[9]) ? node745 : node742;
										assign node742 = (inp[3]) ? 15'b000000111111111 : 15'b000001111111111;
										assign node745 = (inp[3]) ? 15'b000000011111111 : node746;
											assign node746 = (inp[7]) ? 15'b000000001111111 : 15'b000000011111111;
									assign node750 = (inp[14]) ? node752 : 15'b000000011111111;
										assign node752 = (inp[11]) ? 15'b000000001111111 : 15'b000000011111111;
								assign node755 = (inp[6]) ? node765 : node756;
									assign node756 = (inp[11]) ? node762 : node757;
										assign node757 = (inp[8]) ? node759 : 15'b000000011111111;
											assign node759 = (inp[3]) ? 15'b000000000111111 : 15'b000000011111111;
										assign node762 = (inp[9]) ? 15'b000000000011111 : 15'b000000001111111;
									assign node765 = (inp[14]) ? node767 : 15'b000000000111111;
										assign node767 = (inp[3]) ? node769 : 15'b000000001111111;
											assign node769 = (inp[11]) ? 15'b000000000111111 : node770;
												assign node770 = (inp[7]) ? 15'b000000000111111 : 15'b000000001111111;
							assign node774 = (inp[3]) ? node798 : node775;
								assign node775 = (inp[8]) ? node783 : node776;
									assign node776 = (inp[14]) ? node778 : 15'b000000111111111;
										assign node778 = (inp[1]) ? 15'b000000001111111 : node779;
											assign node779 = (inp[7]) ? 15'b000000001111111 : 15'b000000111111111;
									assign node783 = (inp[9]) ? node789 : node784;
										assign node784 = (inp[10]) ? 15'b000000001111111 : node785;
											assign node785 = (inp[14]) ? 15'b000000011111111 : 15'b000000001111111;
										assign node789 = (inp[11]) ? node793 : node790;
											assign node790 = (inp[6]) ? 15'b000000000111111 : 15'b000000001111111;
											assign node793 = (inp[6]) ? node795 : 15'b000000000111111;
												assign node795 = (inp[10]) ? 15'b000000000111111 : 15'b000000000011111;
								assign node798 = (inp[14]) ? node804 : node799;
									assign node799 = (inp[1]) ? 15'b000000000111111 : node800;
										assign node800 = (inp[6]) ? 15'b000000000111111 : 15'b000000001111111;
									assign node804 = (inp[6]) ? 15'b000000000001111 : node805;
										assign node805 = (inp[10]) ? 15'b000000000011111 : 15'b000000001111111;
				assign node809 = (inp[12]) ? node953 : node810;
					assign node810 = (inp[8]) ? node884 : node811;
						assign node811 = (inp[10]) ? node847 : node812;
							assign node812 = (inp[1]) ? node832 : node813;
								assign node813 = (inp[0]) ? node823 : node814;
									assign node814 = (inp[14]) ? node818 : node815;
										assign node815 = (inp[11]) ? 15'b000001111111111 : 15'b000011111111111;
										assign node818 = (inp[9]) ? 15'b000000011111111 : node819;
											assign node819 = (inp[11]) ? 15'b000000111111111 : 15'b000001111111111;
									assign node823 = (inp[9]) ? node827 : node824;
										assign node824 = (inp[14]) ? 15'b000000111111111 : 15'b000001111111111;
										assign node827 = (inp[3]) ? node829 : 15'b000001111111111;
											assign node829 = (inp[13]) ? 15'b000000001111111 : 15'b000000011111111;
								assign node832 = (inp[11]) ? node842 : node833;
									assign node833 = (inp[9]) ? node837 : node834;
										assign node834 = (inp[3]) ? 15'b000000111111111 : 15'b000001111111111;
										assign node837 = (inp[14]) ? node839 : 15'b000000111111111;
											assign node839 = (inp[7]) ? 15'b000000001111111 : 15'b000000011111111;
									assign node842 = (inp[9]) ? 15'b000000011111111 : node843;
										assign node843 = (inp[14]) ? 15'b000000001111111 : 15'b000000000111111;
							assign node847 = (inp[11]) ? node869 : node848;
								assign node848 = (inp[0]) ? node856 : node849;
									assign node849 = (inp[14]) ? node853 : node850;
										assign node850 = (inp[7]) ? 15'b000001111111111 : 15'b000000111111111;
										assign node853 = (inp[1]) ? 15'b000000111111111 : 15'b000000011111111;
									assign node856 = (inp[14]) ? node862 : node857;
										assign node857 = (inp[6]) ? 15'b000000011111111 : node858;
											assign node858 = (inp[13]) ? 15'b000000011111111 : 15'b000000111111111;
										assign node862 = (inp[9]) ? 15'b000000001111111 : node863;
											assign node863 = (inp[13]) ? node865 : 15'b000000011111111;
												assign node865 = (inp[3]) ? 15'b000000001111111 : 15'b000000011111111;
								assign node869 = (inp[7]) ? node873 : node870;
									assign node870 = (inp[6]) ? 15'b000000011111111 : 15'b000000111111111;
									assign node873 = (inp[9]) ? node877 : node874;
										assign node874 = (inp[14]) ? 15'b000000011111111 : 15'b000000001111111;
										assign node877 = (inp[0]) ? node881 : node878;
											assign node878 = (inp[1]) ? 15'b000000000111111 : 15'b000000001111111;
											assign node881 = (inp[1]) ? 15'b000000000011111 : 15'b000000000111111;
						assign node884 = (inp[6]) ? node920 : node885;
							assign node885 = (inp[14]) ? node907 : node886;
								assign node886 = (inp[10]) ? node900 : node887;
									assign node887 = (inp[7]) ? node897 : node888;
										assign node888 = (inp[9]) ? node894 : node889;
											assign node889 = (inp[3]) ? 15'b000001111111111 : node890;
												assign node890 = (inp[11]) ? 15'b000001111111111 : 15'b000011111111111;
											assign node894 = (inp[1]) ? 15'b000001111111111 : 15'b000000111111111;
										assign node897 = (inp[13]) ? 15'b000000111111111 : 15'b000000011111111;
									assign node900 = (inp[0]) ? node904 : node901;
										assign node901 = (inp[3]) ? 15'b000000011111111 : 15'b000000111111111;
										assign node904 = (inp[3]) ? 15'b000000000011111 : 15'b000000011111111;
								assign node907 = (inp[3]) ? node913 : node908;
									assign node908 = (inp[7]) ? 15'b000000111111111 : node909;
										assign node909 = (inp[13]) ? 15'b000000001111111 : 15'b000000011111111;
									assign node913 = (inp[1]) ? node917 : node914;
										assign node914 = (inp[0]) ? 15'b000000000111111 : 15'b000000001111111;
										assign node917 = (inp[0]) ? 15'b000000000011111 : 15'b000000000111111;
							assign node920 = (inp[3]) ? node938 : node921;
								assign node921 = (inp[0]) ? node929 : node922;
									assign node922 = (inp[14]) ? node926 : node923;
										assign node923 = (inp[1]) ? 15'b000000011111111 : 15'b000000001111111;
										assign node926 = (inp[10]) ? 15'b000000011111111 : 15'b000000111111111;
									assign node929 = (inp[7]) ? node933 : node930;
										assign node930 = (inp[11]) ? 15'b000000000111111 : 15'b000000001111111;
										assign node933 = (inp[1]) ? 15'b000000000011111 : node934;
											assign node934 = (inp[11]) ? 15'b000000000011111 : 15'b000000001111111;
								assign node938 = (inp[0]) ? node946 : node939;
									assign node939 = (inp[14]) ? node943 : node940;
										assign node940 = (inp[1]) ? 15'b000000000111111 : 15'b000000001111111;
										assign node943 = (inp[13]) ? 15'b000000000011111 : 15'b000000000111111;
									assign node946 = (inp[13]) ? node948 : 15'b000000000001111;
										assign node948 = (inp[14]) ? 15'b000000000011111 : node949;
											assign node949 = (inp[9]) ? 15'b000000000111111 : 15'b000000000011111;
					assign node953 = (inp[10]) ? node1033 : node954;
						assign node954 = (inp[11]) ? node1000 : node955;
							assign node955 = (inp[7]) ? node975 : node956;
								assign node956 = (inp[1]) ? node964 : node957;
									assign node957 = (inp[3]) ? 15'b000000011111111 : node958;
										assign node958 = (inp[6]) ? node960 : 15'b000001111111111;
											assign node960 = (inp[14]) ? 15'b000000011111111 : 15'b000000111111111;
									assign node964 = (inp[14]) ? node970 : node965;
										assign node965 = (inp[13]) ? 15'b000000001111111 : node966;
											assign node966 = (inp[9]) ? 15'b000000111111111 : 15'b000001111111111;
										assign node970 = (inp[8]) ? 15'b000000000111111 : node971;
											assign node971 = (inp[13]) ? 15'b000000001111111 : 15'b000000011111111;
								assign node975 = (inp[1]) ? node993 : node976;
									assign node976 = (inp[14]) ? node982 : node977;
										assign node977 = (inp[9]) ? node979 : 15'b000000011111111;
											assign node979 = (inp[6]) ? 15'b000000001111111 : 15'b000000011111111;
										assign node982 = (inp[13]) ? node984 : 15'b000000001111111;
											assign node984 = (inp[9]) ? node990 : node985;
												assign node985 = (inp[6]) ? 15'b000000001111111 : node986;
													assign node986 = (inp[3]) ? 15'b000000000111111 : 15'b000000001111111;
												assign node990 = (inp[8]) ? 15'b000000000011111 : 15'b000000000111111;
									assign node993 = (inp[8]) ? node995 : 15'b000000011111111;
										assign node995 = (inp[14]) ? node997 : 15'b000000000111111;
											assign node997 = (inp[9]) ? 15'b000000000001111 : 15'b000000000111111;
							assign node1000 = (inp[13]) ? node1016 : node1001;
								assign node1001 = (inp[1]) ? node1005 : node1002;
									assign node1002 = (inp[9]) ? 15'b000000000111111 : 15'b000000011111111;
									assign node1005 = (inp[14]) ? node1007 : 15'b000000001111111;
										assign node1007 = (inp[0]) ? node1013 : node1008;
											assign node1008 = (inp[3]) ? 15'b000000001111111 : node1009;
												assign node1009 = (inp[9]) ? 15'b000000000111111 : 15'b000000001111111;
											assign node1013 = (inp[6]) ? 15'b000000000011111 : 15'b000000000111111;
								assign node1016 = (inp[8]) ? node1026 : node1017;
									assign node1017 = (inp[7]) ? node1019 : 15'b000000001111111;
										assign node1019 = (inp[0]) ? node1023 : node1020;
											assign node1020 = (inp[14]) ? 15'b000000000111111 : 15'b000000001111111;
											assign node1023 = (inp[1]) ? 15'b000000000011111 : 15'b000000000111111;
									assign node1026 = (inp[3]) ? node1028 : 15'b000000000111111;
										assign node1028 = (inp[0]) ? node1030 : 15'b000000000011111;
											assign node1030 = (inp[14]) ? 15'b000000000000111 : 15'b000000000001111;
						assign node1033 = (inp[9]) ? node1063 : node1034;
							assign node1034 = (inp[3]) ? node1048 : node1035;
								assign node1035 = (inp[13]) ? node1039 : node1036;
									assign node1036 = (inp[14]) ? 15'b000000001111111 : 15'b000000011111111;
									assign node1039 = (inp[6]) ? node1041 : 15'b000000011111111;
										assign node1041 = (inp[1]) ? node1045 : node1042;
											assign node1042 = (inp[8]) ? 15'b000000000111111 : 15'b000000001111111;
											assign node1045 = (inp[14]) ? 15'b000000000001111 : 15'b000000000111111;
								assign node1048 = (inp[6]) ? node1058 : node1049;
									assign node1049 = (inp[0]) ? node1053 : node1050;
										assign node1050 = (inp[1]) ? 15'b000000000111111 : 15'b000000001111111;
										assign node1053 = (inp[14]) ? 15'b000000000111111 : node1054;
											assign node1054 = (inp[1]) ? 15'b000000000011111 : 15'b000000000111111;
									assign node1058 = (inp[11]) ? 15'b000000000001111 : node1059;
										assign node1059 = (inp[0]) ? 15'b000000000001111 : 15'b000000000111111;
							assign node1063 = (inp[11]) ? node1089 : node1064;
								assign node1064 = (inp[1]) ? node1080 : node1065;
									assign node1065 = (inp[13]) ? node1071 : node1066;
										assign node1066 = (inp[0]) ? node1068 : 15'b000000011111111;
											assign node1068 = (inp[6]) ? 15'b000000000111111 : 15'b000000001111111;
										assign node1071 = (inp[6]) ? 15'b000000000011111 : node1072;
											assign node1072 = (inp[3]) ? 15'b000000000001111 : node1073;
												assign node1073 = (inp[7]) ? node1075 : 15'b000000001111111;
													assign node1075 = (inp[14]) ? 15'b000000001111111 : 15'b000000000111111;
									assign node1080 = (inp[3]) ? 15'b000000000001111 : node1081;
										assign node1081 = (inp[13]) ? node1083 : 15'b000000000111111;
											assign node1083 = (inp[8]) ? node1085 : 15'b000000000111111;
												assign node1085 = (inp[0]) ? 15'b000000000001111 : 15'b000000000011111;
								assign node1089 = (inp[6]) ? node1097 : node1090;
									assign node1090 = (inp[1]) ? node1094 : node1091;
										assign node1091 = (inp[3]) ? 15'b000000000001111 : 15'b000000000011111;
										assign node1094 = (inp[13]) ? 15'b000000000011111 : 15'b000000000111111;
									assign node1097 = (inp[1]) ? node1099 : 15'b000000000011111;
										assign node1099 = (inp[8]) ? node1101 : 15'b000000000001111;
											assign node1101 = (inp[3]) ? node1103 : 15'b000000000000111;
												assign node1103 = (inp[0]) ? 15'b000000000000011 : 15'b000000000000111;
		assign node1106 = (inp[10]) ? node1686 : node1107;
			assign node1107 = (inp[5]) ? node1375 : node1108;
				assign node1108 = (inp[14]) ? node1256 : node1109;
					assign node1109 = (inp[7]) ? node1187 : node1110;
						assign node1110 = (inp[9]) ? node1148 : node1111;
							assign node1111 = (inp[6]) ? node1133 : node1112;
								assign node1112 = (inp[0]) ? node1118 : node1113;
									assign node1113 = (inp[12]) ? node1115 : 15'b000111111111111;
										assign node1115 = (inp[11]) ? 15'b000001111111111 : 15'b000011111111111;
									assign node1118 = (inp[1]) ? node1128 : node1119;
										assign node1119 = (inp[3]) ? node1125 : node1120;
											assign node1120 = (inp[12]) ? node1122 : 15'b000011111111111;
												assign node1122 = (inp[8]) ? 15'b000001111111111 : 15'b000011111111111;
											assign node1125 = (inp[2]) ? 15'b000000111111111 : 15'b000011111111111;
										assign node1128 = (inp[8]) ? 15'b000000011111111 : node1129;
											assign node1129 = (inp[13]) ? 15'b000000111111111 : 15'b000001111111111;
								assign node1133 = (inp[2]) ? node1143 : node1134;
									assign node1134 = (inp[1]) ? 15'b000000111111111 : node1135;
										assign node1135 = (inp[8]) ? node1139 : node1136;
											assign node1136 = (inp[11]) ? 15'b000001111111111 : 15'b000011111111111;
											assign node1139 = (inp[3]) ? 15'b000000111111111 : 15'b000001111111111;
									assign node1143 = (inp[8]) ? node1145 : 15'b000000111111111;
										assign node1145 = (inp[1]) ? 15'b000000001111111 : 15'b000000011111111;
							assign node1148 = (inp[13]) ? node1176 : node1149;
								assign node1149 = (inp[2]) ? node1169 : node1150;
									assign node1150 = (inp[3]) ? node1162 : node1151;
										assign node1151 = (inp[11]) ? node1155 : node1152;
											assign node1152 = (inp[6]) ? 15'b000011111111111 : 15'b000111111111111;
											assign node1155 = (inp[6]) ? node1157 : 15'b000001111111111;
												assign node1157 = (inp[8]) ? 15'b000000111111111 : node1158;
													assign node1158 = (inp[1]) ? 15'b000000111111111 : 15'b000001111111111;
										assign node1162 = (inp[8]) ? node1164 : 15'b000001111111111;
											assign node1164 = (inp[11]) ? 15'b000000011111111 : node1165;
												assign node1165 = (inp[1]) ? 15'b000000011111111 : 15'b000000111111111;
									assign node1169 = (inp[12]) ? node1173 : node1170;
										assign node1170 = (inp[11]) ? 15'b000000111111111 : 15'b000000011111111;
										assign node1173 = (inp[11]) ? 15'b000000011111111 : 15'b000000111111111;
								assign node1176 = (inp[6]) ? node1184 : node1177;
									assign node1177 = (inp[0]) ? node1179 : 15'b000001111111111;
										assign node1179 = (inp[3]) ? node1181 : 15'b000000011111111;
											assign node1181 = (inp[2]) ? 15'b000000001111111 : 15'b000000011111111;
									assign node1184 = (inp[3]) ? 15'b000000000111111 : 15'b000000001111111;
						assign node1187 = (inp[3]) ? node1223 : node1188;
							assign node1188 = (inp[11]) ? node1202 : node1189;
								assign node1189 = (inp[12]) ? node1199 : node1190;
									assign node1190 = (inp[0]) ? node1196 : node1191;
										assign node1191 = (inp[6]) ? node1193 : 15'b000011111111111;
											assign node1193 = (inp[1]) ? 15'b000001111111111 : 15'b000011111111111;
										assign node1196 = (inp[1]) ? 15'b000001111111111 : 15'b000000111111111;
									assign node1199 = (inp[2]) ? 15'b000000001111111 : 15'b000000111111111;
								assign node1202 = (inp[6]) ? node1212 : node1203;
									assign node1203 = (inp[8]) ? node1209 : node1204;
										assign node1204 = (inp[2]) ? node1206 : 15'b000000111111111;
											assign node1206 = (inp[0]) ? 15'b000000011111111 : 15'b000000111111111;
										assign node1209 = (inp[13]) ? 15'b000000111111111 : 15'b000001111111111;
									assign node1212 = (inp[0]) ? node1214 : 15'b000000011111111;
										assign node1214 = (inp[1]) ? node1218 : node1215;
											assign node1215 = (inp[12]) ? 15'b000000001111111 : 15'b000000111111111;
											assign node1218 = (inp[12]) ? node1220 : 15'b000000001111111;
												assign node1220 = (inp[9]) ? 15'b000000000111111 : 15'b000000001111111;
							assign node1223 = (inp[8]) ? node1237 : node1224;
								assign node1224 = (inp[0]) ? node1230 : node1225;
									assign node1225 = (inp[12]) ? node1227 : 15'b000000111111111;
										assign node1227 = (inp[9]) ? 15'b000000011111111 : 15'b000001111111111;
									assign node1230 = (inp[1]) ? 15'b000000000111111 : node1231;
										assign node1231 = (inp[13]) ? 15'b000000011111111 : node1232;
											assign node1232 = (inp[9]) ? 15'b000000011111111 : 15'b000000111111111;
								assign node1237 = (inp[6]) ? node1251 : node1238;
									assign node1238 = (inp[9]) ? node1242 : node1239;
										assign node1239 = (inp[1]) ? 15'b000000011111111 : 15'b000000111111111;
										assign node1242 = (inp[12]) ? node1248 : node1243;
											assign node1243 = (inp[2]) ? node1245 : 15'b000000011111111;
												assign node1245 = (inp[1]) ? 15'b000000001111111 : 15'b000000011111111;
											assign node1248 = (inp[11]) ? 15'b000000000111111 : 15'b000000001111111;
									assign node1251 = (inp[2]) ? node1253 : 15'b000000001111111;
										assign node1253 = (inp[0]) ? 15'b000000000111111 : 15'b000000001111111;
					assign node1256 = (inp[9]) ? node1314 : node1257;
						assign node1257 = (inp[11]) ? node1279 : node1258;
							assign node1258 = (inp[1]) ? node1270 : node1259;
								assign node1259 = (inp[8]) ? node1265 : node1260;
									assign node1260 = (inp[13]) ? node1262 : 15'b000001111111111;
										assign node1262 = (inp[7]) ? 15'b000000011111111 : 15'b000000111111111;
									assign node1265 = (inp[12]) ? node1267 : 15'b000000111111111;
										assign node1267 = (inp[3]) ? 15'b000000001111111 : 15'b000001111111111;
								assign node1270 = (inp[6]) ? node1276 : node1271;
									assign node1271 = (inp[8]) ? node1273 : 15'b000000111111111;
										assign node1273 = (inp[0]) ? 15'b000000011111111 : 15'b000000111111111;
									assign node1276 = (inp[3]) ? 15'b000000001111111 : 15'b000000011111111;
							assign node1279 = (inp[12]) ? node1301 : node1280;
								assign node1280 = (inp[8]) ? node1288 : node1281;
									assign node1281 = (inp[0]) ? node1285 : node1282;
										assign node1282 = (inp[1]) ? 15'b000000111111111 : 15'b000001111111111;
										assign node1285 = (inp[2]) ? 15'b000000011111111 : 15'b000000111111111;
									assign node1288 = (inp[1]) ? node1292 : node1289;
										assign node1289 = (inp[7]) ? 15'b000000111111111 : 15'b000000011111111;
										assign node1292 = (inp[13]) ? node1298 : node1293;
											assign node1293 = (inp[7]) ? node1295 : 15'b000000001111111;
												assign node1295 = (inp[6]) ? 15'b000000001111111 : 15'b000000011111111;
											assign node1298 = (inp[2]) ? 15'b000000000011111 : 15'b000000001111111;
								assign node1301 = (inp[1]) ? node1303 : 15'b000000001111111;
									assign node1303 = (inp[3]) ? node1311 : node1304;
										assign node1304 = (inp[7]) ? node1306 : 15'b000000011111111;
											assign node1306 = (inp[0]) ? node1308 : 15'b000000001111111;
												assign node1308 = (inp[2]) ? 15'b000000000111111 : 15'b000000001111111;
										assign node1311 = (inp[7]) ? 15'b000000000011111 : 15'b000000000111111;
						assign node1314 = (inp[2]) ? node1346 : node1315;
							assign node1315 = (inp[3]) ? node1327 : node1316;
								assign node1316 = (inp[7]) ? node1322 : node1317;
									assign node1317 = (inp[11]) ? node1319 : 15'b000001111111111;
										assign node1319 = (inp[13]) ? 15'b000000001111111 : 15'b000000011111111;
									assign node1322 = (inp[8]) ? 15'b000000011111111 : node1323;
										assign node1323 = (inp[1]) ? 15'b000000001111111 : 15'b000000011111111;
								assign node1327 = (inp[6]) ? node1333 : node1328;
									assign node1328 = (inp[1]) ? 15'b000000011111111 : node1329;
										assign node1329 = (inp[11]) ? 15'b000000000111111 : 15'b000000001111111;
									assign node1333 = (inp[8]) ? node1335 : 15'b000000011111111;
										assign node1335 = (inp[1]) ? node1341 : node1336;
											assign node1336 = (inp[11]) ? 15'b000000000111111 : node1337;
												assign node1337 = (inp[7]) ? 15'b000000000111111 : 15'b000000011111111;
											assign node1341 = (inp[11]) ? 15'b000000000011111 : node1342;
												assign node1342 = (inp[7]) ? 15'b000000000011111 : 15'b000000000111111;
							assign node1346 = (inp[7]) ? node1356 : node1347;
								assign node1347 = (inp[6]) ? node1351 : node1348;
									assign node1348 = (inp[13]) ? 15'b000000011111111 : 15'b000000001111111;
									assign node1351 = (inp[0]) ? 15'b000000000111111 : node1352;
										assign node1352 = (inp[8]) ? 15'b000000000111111 : 15'b000000001111111;
								assign node1356 = (inp[3]) ? node1364 : node1357;
									assign node1357 = (inp[0]) ? node1361 : node1358;
										assign node1358 = (inp[13]) ? 15'b000000000111111 : 15'b000000001111111;
										assign node1361 = (inp[8]) ? 15'b000000000000111 : 15'b000000000111111;
									assign node1364 = (inp[8]) ? node1370 : node1365;
										assign node1365 = (inp[0]) ? 15'b000000000011111 : node1366;
											assign node1366 = (inp[11]) ? 15'b000000000011111 : 15'b000000011111111;
										assign node1370 = (inp[6]) ? node1372 : 15'b000000000011111;
											assign node1372 = (inp[0]) ? 15'b000000000000111 : 15'b000000000011111;
				assign node1375 = (inp[12]) ? node1517 : node1376;
					assign node1376 = (inp[3]) ? node1454 : node1377;
						assign node1377 = (inp[8]) ? node1423 : node1378;
							assign node1378 = (inp[7]) ? node1402 : node1379;
								assign node1379 = (inp[2]) ? node1387 : node1380;
									assign node1380 = (inp[14]) ? node1382 : 15'b000001111111111;
										assign node1382 = (inp[9]) ? 15'b000000111111111 : node1383;
											assign node1383 = (inp[11]) ? 15'b000011111111111 : 15'b000001111111111;
									assign node1387 = (inp[13]) ? node1397 : node1388;
										assign node1388 = (inp[0]) ? 15'b000000111111111 : node1389;
											assign node1389 = (inp[1]) ? node1391 : 15'b000001111111111;
												assign node1391 = (inp[9]) ? 15'b000000111111111 : node1392;
													assign node1392 = (inp[11]) ? 15'b000000111111111 : 15'b000001111111111;
										assign node1397 = (inp[9]) ? node1399 : 15'b000000111111111;
											assign node1399 = (inp[0]) ? 15'b000000001111111 : 15'b000000011111111;
								assign node1402 = (inp[14]) ? node1418 : node1403;
									assign node1403 = (inp[6]) ? node1411 : node1404;
										assign node1404 = (inp[1]) ? node1406 : 15'b000000111111111;
											assign node1406 = (inp[13]) ? 15'b000000111111111 : node1407;
												assign node1407 = (inp[11]) ? 15'b000000111111111 : 15'b000001111111111;
										assign node1411 = (inp[1]) ? 15'b000000001111111 : node1412;
											assign node1412 = (inp[11]) ? 15'b000000011111111 : node1413;
												assign node1413 = (inp[0]) ? 15'b000000111111111 : 15'b000000011111111;
									assign node1418 = (inp[0]) ? node1420 : 15'b000000111111111;
										assign node1420 = (inp[9]) ? 15'b000000000111111 : 15'b000000001111111;
							assign node1423 = (inp[9]) ? node1441 : node1424;
								assign node1424 = (inp[14]) ? node1436 : node1425;
									assign node1425 = (inp[11]) ? node1433 : node1426;
										assign node1426 = (inp[2]) ? node1430 : node1427;
											assign node1427 = (inp[1]) ? 15'b000011111111111 : 15'b000001111111111;
											assign node1430 = (inp[6]) ? 15'b000000111111111 : 15'b000000011111111;
										assign node1433 = (inp[7]) ? 15'b000000011111111 : 15'b000000001111111;
									assign node1436 = (inp[11]) ? node1438 : 15'b000000011111111;
										assign node1438 = (inp[6]) ? 15'b000000011111111 : 15'b000000111111111;
								assign node1441 = (inp[6]) ? node1445 : node1442;
									assign node1442 = (inp[1]) ? 15'b000000001111111 : 15'b000000011111111;
									assign node1445 = (inp[2]) ? node1447 : 15'b000000001111111;
										assign node1447 = (inp[13]) ? node1449 : 15'b000000000111111;
											assign node1449 = (inp[11]) ? node1451 : 15'b000000000111111;
												assign node1451 = (inp[14]) ? 15'b000000000001111 : 15'b000000000011111;
						assign node1454 = (inp[1]) ? node1484 : node1455;
							assign node1455 = (inp[8]) ? node1469 : node1456;
								assign node1456 = (inp[9]) ? node1458 : 15'b000001111111111;
									assign node1458 = (inp[6]) ? node1466 : node1459;
										assign node1459 = (inp[11]) ? node1461 : 15'b000000111111111;
											assign node1461 = (inp[14]) ? node1463 : 15'b000000011111111;
												assign node1463 = (inp[13]) ? 15'b000000011111111 : 15'b000000111111111;
										assign node1466 = (inp[11]) ? 15'b000000000111111 : 15'b000000011111111;
								assign node1469 = (inp[0]) ? node1477 : node1470;
									assign node1470 = (inp[11]) ? node1472 : 15'b000000011111111;
										assign node1472 = (inp[9]) ? 15'b000000001111111 : node1473;
											assign node1473 = (inp[6]) ? 15'b000000000111111 : 15'b000000001111111;
									assign node1477 = (inp[14]) ? node1481 : node1478;
										assign node1478 = (inp[9]) ? 15'b000000000111111 : 15'b000000001111111;
										assign node1481 = (inp[7]) ? 15'b000000000011111 : 15'b000000000111111;
							assign node1484 = (inp[9]) ? node1502 : node1485;
								assign node1485 = (inp[11]) ? node1491 : node1486;
									assign node1486 = (inp[7]) ? node1488 : 15'b000000011111111;
										assign node1488 = (inp[8]) ? 15'b000000011111111 : 15'b000000001111111;
									assign node1491 = (inp[6]) ? node1497 : node1492;
										assign node1492 = (inp[14]) ? 15'b000000000111111 : node1493;
											assign node1493 = (inp[2]) ? 15'b000000001111111 : 15'b000000011111111;
										assign node1497 = (inp[13]) ? node1499 : 15'b000000000111111;
											assign node1499 = (inp[2]) ? 15'b000000000001111 : 15'b000000000011111;
								assign node1502 = (inp[8]) ? node1510 : node1503;
									assign node1503 = (inp[13]) ? node1505 : 15'b000000000111111;
										assign node1505 = (inp[6]) ? node1507 : 15'b000000000111111;
											assign node1507 = (inp[0]) ? 15'b000000000011111 : 15'b000000000111111;
									assign node1510 = (inp[14]) ? node1512 : 15'b000000001111111;
										assign node1512 = (inp[0]) ? 15'b000000000001111 : node1513;
											assign node1513 = (inp[11]) ? 15'b000000000111111 : 15'b000000000011111;
					assign node1517 = (inp[7]) ? node1593 : node1518;
						assign node1518 = (inp[14]) ? node1558 : node1519;
							assign node1519 = (inp[9]) ? node1537 : node1520;
								assign node1520 = (inp[11]) ? node1528 : node1521;
									assign node1521 = (inp[8]) ? 15'b000000011111111 : node1522;
										assign node1522 = (inp[3]) ? node1524 : 15'b000001111111111;
											assign node1524 = (inp[13]) ? 15'b000001111111111 : 15'b000000111111111;
									assign node1528 = (inp[0]) ? node1534 : node1529;
										assign node1529 = (inp[1]) ? node1531 : 15'b000000111111111;
											assign node1531 = (inp[2]) ? 15'b000000011111111 : 15'b000000111111111;
										assign node1534 = (inp[1]) ? 15'b000000001111111 : 15'b000000011111111;
								assign node1537 = (inp[11]) ? node1547 : node1538;
									assign node1538 = (inp[13]) ? node1542 : node1539;
										assign node1539 = (inp[2]) ? 15'b000000011111111 : 15'b000000111111111;
										assign node1542 = (inp[1]) ? node1544 : 15'b000000011111111;
											assign node1544 = (inp[3]) ? 15'b000000000111111 : 15'b000000001111111;
									assign node1547 = (inp[8]) ? node1551 : node1548;
										assign node1548 = (inp[6]) ? 15'b000000000111111 : 15'b000000011111111;
										assign node1551 = (inp[6]) ? node1553 : 15'b000000000111111;
											assign node1553 = (inp[3]) ? node1555 : 15'b000000000011111;
												assign node1555 = (inp[13]) ? 15'b000000000011111 : 15'b000000000111111;
							assign node1558 = (inp[2]) ? node1572 : node1559;
								assign node1559 = (inp[8]) ? node1565 : node1560;
									assign node1560 = (inp[9]) ? 15'b000000001111111 : node1561;
										assign node1561 = (inp[13]) ? 15'b000000001111111 : 15'b000000011111111;
									assign node1565 = (inp[3]) ? node1569 : node1566;
										assign node1566 = (inp[11]) ? 15'b000000000111111 : 15'b000000001111111;
										assign node1569 = (inp[1]) ? 15'b000000000111111 : 15'b000000000011111;
								assign node1572 = (inp[0]) ? node1580 : node1573;
									assign node1573 = (inp[13]) ? node1577 : node1574;
										assign node1574 = (inp[11]) ? 15'b000000001111111 : 15'b000000000111111;
										assign node1577 = (inp[9]) ? 15'b000000000111111 : 15'b000000000011111;
									assign node1580 = (inp[1]) ? node1586 : node1581;
										assign node1581 = (inp[11]) ? 15'b000000000111111 : node1582;
											assign node1582 = (inp[13]) ? 15'b000000000111111 : 15'b000000000011111;
										assign node1586 = (inp[3]) ? node1590 : node1587;
											assign node1587 = (inp[13]) ? 15'b000000000011111 : 15'b000000001111111;
											assign node1590 = (inp[13]) ? 15'b000000000001111 : 15'b000000000011111;
						assign node1593 = (inp[13]) ? node1647 : node1594;
							assign node1594 = (inp[2]) ? node1622 : node1595;
								assign node1595 = (inp[0]) ? node1609 : node1596;
									assign node1596 = (inp[8]) ? node1602 : node1597;
										assign node1597 = (inp[9]) ? node1599 : 15'b000000111111111;
											assign node1599 = (inp[3]) ? 15'b000000001111111 : 15'b000000011111111;
										assign node1602 = (inp[11]) ? 15'b000000011111111 : node1603;
											assign node1603 = (inp[9]) ? node1605 : 15'b000000001111111;
												assign node1605 = (inp[14]) ? 15'b000000000111111 : 15'b000000001111111;
									assign node1609 = (inp[8]) ? node1615 : node1610;
										assign node1610 = (inp[9]) ? node1612 : 15'b000000001111111;
											assign node1612 = (inp[3]) ? 15'b000000000111111 : 15'b000000001111111;
										assign node1615 = (inp[6]) ? 15'b000000000011111 : node1616;
											assign node1616 = (inp[1]) ? 15'b000000000011111 : node1617;
												assign node1617 = (inp[9]) ? 15'b000000000111111 : 15'b000000001111111;
								assign node1622 = (inp[3]) ? node1634 : node1623;
									assign node1623 = (inp[11]) ? node1629 : node1624;
										assign node1624 = (inp[8]) ? 15'b000000000111111 : node1625;
											assign node1625 = (inp[14]) ? 15'b000000000111111 : 15'b000000001111111;
										assign node1629 = (inp[14]) ? node1631 : 15'b000000011111111;
											assign node1631 = (inp[8]) ? 15'b000000000111111 : 15'b000000001111111;
									assign node1634 = (inp[9]) ? node1636 : 15'b000000000111111;
										assign node1636 = (inp[8]) ? node1644 : node1637;
											assign node1637 = (inp[14]) ? 15'b000000000011111 : node1638;
												assign node1638 = (inp[11]) ? node1640 : 15'b000000000111111;
													assign node1640 = (inp[1]) ? 15'b000000000011111 : 15'b000000000111111;
											assign node1644 = (inp[14]) ? 15'b000000000000111 : 15'b000000000011111;
							assign node1647 = (inp[2]) ? node1665 : node1648;
								assign node1648 = (inp[3]) ? node1654 : node1649;
									assign node1649 = (inp[14]) ? node1651 : 15'b000000001111111;
										assign node1651 = (inp[6]) ? 15'b000000000111111 : 15'b000000000011111;
									assign node1654 = (inp[0]) ? node1660 : node1655;
										assign node1655 = (inp[11]) ? 15'b000000000011111 : node1656;
											assign node1656 = (inp[14]) ? 15'b000000000111111 : 15'b000000011111111;
										assign node1660 = (inp[14]) ? 15'b000000000011111 : node1661;
											assign node1661 = (inp[1]) ? 15'b000000000001111 : 15'b000000000011111;
								assign node1665 = (inp[8]) ? node1675 : node1666;
									assign node1666 = (inp[3]) ? node1672 : node1667;
										assign node1667 = (inp[0]) ? node1669 : 15'b000000000111111;
											assign node1669 = (inp[1]) ? 15'b000000000111111 : 15'b000000000011111;
										assign node1672 = (inp[0]) ? 15'b000000000011111 : 15'b000000000001111;
									assign node1675 = (inp[14]) ? node1681 : node1676;
										assign node1676 = (inp[1]) ? node1678 : 15'b000000000011111;
											assign node1678 = (inp[9]) ? 15'b000000000000111 : 15'b000000000011111;
										assign node1681 = (inp[0]) ? 15'b000000000000111 : node1682;
											assign node1682 = (inp[3]) ? 15'b000000000000111 : 15'b000000000001111;
			assign node1686 = (inp[8]) ? node1950 : node1687;
				assign node1687 = (inp[0]) ? node1825 : node1688;
					assign node1688 = (inp[6]) ? node1760 : node1689;
						assign node1689 = (inp[11]) ? node1731 : node1690;
							assign node1690 = (inp[13]) ? node1714 : node1691;
								assign node1691 = (inp[2]) ? node1705 : node1692;
									assign node1692 = (inp[12]) ? node1698 : node1693;
										assign node1693 = (inp[9]) ? 15'b000001111111111 : node1694;
											assign node1694 = (inp[5]) ? 15'b000111111111111 : 15'b000011111111111;
										assign node1698 = (inp[1]) ? 15'b000000111111111 : node1699;
											assign node1699 = (inp[14]) ? node1701 : 15'b000001111111111;
												assign node1701 = (inp[5]) ? 15'b000000111111111 : 15'b000001111111111;
									assign node1705 = (inp[7]) ? node1709 : node1706;
										assign node1706 = (inp[12]) ? 15'b000011111111111 : 15'b000000111111111;
										assign node1709 = (inp[14]) ? 15'b000000001111111 : node1710;
											assign node1710 = (inp[12]) ? 15'b000000011111111 : 15'b000000111111111;
								assign node1714 = (inp[3]) ? node1720 : node1715;
									assign node1715 = (inp[12]) ? 15'b000000011111111 : node1716;
										assign node1716 = (inp[14]) ? 15'b000001111111111 : 15'b000000111111111;
									assign node1720 = (inp[5]) ? node1722 : 15'b000000111111111;
										assign node1722 = (inp[9]) ? node1724 : 15'b000000011111111;
											assign node1724 = (inp[12]) ? 15'b000000000011111 : node1725;
												assign node1725 = (inp[1]) ? 15'b000000001111111 : node1726;
													assign node1726 = (inp[7]) ? 15'b000000001111111 : 15'b000000011111111;
							assign node1731 = (inp[9]) ? node1745 : node1732;
								assign node1732 = (inp[5]) ? 15'b000000011111111 : node1733;
									assign node1733 = (inp[14]) ? node1739 : node1734;
										assign node1734 = (inp[3]) ? 15'b000000011111111 : node1735;
											assign node1735 = (inp[13]) ? 15'b000000111111111 : 15'b000001111111111;
										assign node1739 = (inp[3]) ? 15'b000000001111111 : node1740;
											assign node1740 = (inp[12]) ? 15'b000000001111111 : 15'b000000111111111;
								assign node1745 = (inp[2]) ? node1753 : node1746;
									assign node1746 = (inp[1]) ? node1748 : 15'b000000011111111;
										assign node1748 = (inp[3]) ? node1750 : 15'b000000001111111;
											assign node1750 = (inp[5]) ? 15'b000000001111111 : 15'b000000011111111;
									assign node1753 = (inp[1]) ? node1757 : node1754;
										assign node1754 = (inp[3]) ? 15'b000000000111111 : 15'b000000001111111;
										assign node1757 = (inp[7]) ? 15'b000000000111111 : 15'b000000000011111;
						assign node1760 = (inp[5]) ? node1788 : node1761;
							assign node1761 = (inp[1]) ? node1773 : node1762;
								assign node1762 = (inp[9]) ? node1768 : node1763;
									assign node1763 = (inp[14]) ? 15'b000000001111111 : node1764;
										assign node1764 = (inp[11]) ? 15'b000001111111111 : 15'b000011111111111;
									assign node1768 = (inp[7]) ? node1770 : 15'b000000011111111;
										assign node1770 = (inp[13]) ? 15'b000000001111111 : 15'b000000011111111;
								assign node1773 = (inp[2]) ? node1781 : node1774;
									assign node1774 = (inp[7]) ? 15'b000000001111111 : node1775;
										assign node1775 = (inp[11]) ? 15'b000000001111111 : node1776;
											assign node1776 = (inp[12]) ? 15'b000000011111111 : 15'b000000111111111;
									assign node1781 = (inp[12]) ? node1783 : 15'b000000001111111;
										assign node1783 = (inp[3]) ? 15'b000000000111111 : node1784;
											assign node1784 = (inp[9]) ? 15'b000000000111111 : 15'b000000001111111;
							assign node1788 = (inp[13]) ? node1812 : node1789;
								assign node1789 = (inp[12]) ? node1801 : node1790;
									assign node1790 = (inp[11]) ? node1796 : node1791;
										assign node1791 = (inp[3]) ? node1793 : 15'b000000111111111;
											assign node1793 = (inp[7]) ? 15'b000000001111111 : 15'b000000011111111;
										assign node1796 = (inp[7]) ? node1798 : 15'b000000001111111;
											assign node1798 = (inp[2]) ? 15'b000000001111111 : 15'b000000011111111;
									assign node1801 = (inp[9]) ? 15'b000000000111111 : node1802;
										assign node1802 = (inp[3]) ? node1804 : 15'b000000001111111;
											assign node1804 = (inp[2]) ? 15'b000000000111111 : node1805;
												assign node1805 = (inp[14]) ? 15'b000000001111111 : node1806;
													assign node1806 = (inp[7]) ? 15'b000000000111111 : 15'b000000001111111;
								assign node1812 = (inp[11]) ? node1816 : node1813;
									assign node1813 = (inp[9]) ? 15'b000000000111111 : 15'b000000001111111;
									assign node1816 = (inp[7]) ? node1818 : 15'b000000000111111;
										assign node1818 = (inp[12]) ? node1822 : node1819;
											assign node1819 = (inp[1]) ? 15'b000000000001111 : 15'b000000000011111;
											assign node1822 = (inp[1]) ? 15'b000000000000111 : 15'b000000000001111;
					assign node1825 = (inp[7]) ? node1881 : node1826;
						assign node1826 = (inp[14]) ? node1848 : node1827;
							assign node1827 = (inp[3]) ? node1841 : node1828;
								assign node1828 = (inp[5]) ? node1836 : node1829;
									assign node1829 = (inp[11]) ? node1833 : node1830;
										assign node1830 = (inp[9]) ? 15'b000000111111111 : 15'b000001111111111;
										assign node1833 = (inp[9]) ? 15'b000000011111111 : 15'b000000111111111;
									assign node1836 = (inp[1]) ? 15'b000000001111111 : node1837;
										assign node1837 = (inp[2]) ? 15'b000000001111111 : 15'b000000111111111;
								assign node1841 = (inp[6]) ? node1845 : node1842;
									assign node1842 = (inp[5]) ? 15'b000000001111111 : 15'b000000011111111;
									assign node1845 = (inp[11]) ? 15'b000000000111111 : 15'b000000000011111;
							assign node1848 = (inp[11]) ? node1864 : node1849;
								assign node1849 = (inp[9]) ? node1857 : node1850;
									assign node1850 = (inp[13]) ? node1852 : 15'b000001111111111;
										assign node1852 = (inp[6]) ? 15'b000000001111111 : node1853;
											assign node1853 = (inp[1]) ? 15'b000000001111111 : 15'b000000011111111;
									assign node1857 = (inp[5]) ? 15'b000000000111111 : node1858;
										assign node1858 = (inp[1]) ? 15'b000000001111111 : node1859;
											assign node1859 = (inp[13]) ? 15'b000000000111111 : 15'b000000001111111;
								assign node1864 = (inp[13]) ? node1872 : node1865;
									assign node1865 = (inp[12]) ? node1867 : 15'b000000011111111;
										assign node1867 = (inp[9]) ? node1869 : 15'b000000000111111;
											assign node1869 = (inp[6]) ? 15'b000000000111111 : 15'b000000001111111;
									assign node1872 = (inp[1]) ? node1878 : node1873;
										assign node1873 = (inp[6]) ? node1875 : 15'b000000000111111;
											assign node1875 = (inp[9]) ? 15'b000000000011111 : 15'b000000000111111;
										assign node1878 = (inp[3]) ? 15'b000000000000111 : 15'b000000000011111;
						assign node1881 = (inp[11]) ? node1909 : node1882;
							assign node1882 = (inp[13]) ? node1900 : node1883;
								assign node1883 = (inp[2]) ? node1889 : node1884;
									assign node1884 = (inp[1]) ? node1886 : 15'b000000011111111;
										assign node1886 = (inp[3]) ? 15'b000000000111111 : 15'b000000001111111;
									assign node1889 = (inp[1]) ? 15'b000000000111111 : node1890;
										assign node1890 = (inp[3]) ? node1892 : 15'b000000001111111;
											assign node1892 = (inp[5]) ? 15'b000000000111111 : node1893;
												assign node1893 = (inp[9]) ? node1895 : 15'b000000001111111;
													assign node1895 = (inp[12]) ? 15'b000000000111111 : 15'b000000001111111;
								assign node1900 = (inp[12]) ? node1904 : node1901;
									assign node1901 = (inp[14]) ? 15'b000000001111111 : 15'b000000000111111;
									assign node1904 = (inp[9]) ? 15'b000000000001111 : node1905;
										assign node1905 = (inp[3]) ? 15'b000000000011111 : 15'b000000000111111;
							assign node1909 = (inp[2]) ? node1927 : node1910;
								assign node1910 = (inp[9]) ? node1918 : node1911;
									assign node1911 = (inp[3]) ? node1915 : node1912;
										assign node1912 = (inp[12]) ? 15'b000000001111111 : 15'b000000011111111;
										assign node1915 = (inp[1]) ? 15'b000000000111111 : 15'b000000001111111;
									assign node1918 = (inp[13]) ? node1922 : node1919;
										assign node1919 = (inp[6]) ? 15'b000000000011111 : 15'b000000001111111;
										assign node1922 = (inp[6]) ? 15'b000000000011111 : node1923;
											assign node1923 = (inp[3]) ? 15'b000000000001111 : 15'b000000000011111;
								assign node1927 = (inp[14]) ? node1937 : node1928;
									assign node1928 = (inp[1]) ? node1934 : node1929;
										assign node1929 = (inp[6]) ? node1931 : 15'b000000001111111;
											assign node1931 = (inp[13]) ? 15'b000000000011111 : 15'b000000000111111;
										assign node1934 = (inp[13]) ? 15'b000000000001111 : 15'b000000000011111;
									assign node1937 = (inp[5]) ? node1945 : node1938;
										assign node1938 = (inp[9]) ? 15'b000000000001111 : node1939;
											assign node1939 = (inp[3]) ? node1941 : 15'b000000000011111;
												assign node1941 = (inp[12]) ? 15'b000000000001111 : 15'b000000000011111;
										assign node1945 = (inp[3]) ? node1947 : 15'b000000000001111;
											assign node1947 = (inp[6]) ? 15'b000000000001111 : 15'b000000000000111;
				assign node1950 = (inp[13]) ? node2078 : node1951;
					assign node1951 = (inp[2]) ? node2021 : node1952;
						assign node1952 = (inp[12]) ? node1984 : node1953;
							assign node1953 = (inp[7]) ? node1975 : node1954;
								assign node1954 = (inp[11]) ? node1964 : node1955;
									assign node1955 = (inp[0]) ? node1961 : node1956;
										assign node1956 = (inp[3]) ? node1958 : 15'b000001111111111;
											assign node1958 = (inp[14]) ? 15'b000000111111111 : 15'b000001111111111;
										assign node1961 = (inp[14]) ? 15'b000000011111111 : 15'b000000111111111;
									assign node1964 = (inp[5]) ? node1970 : node1965;
										assign node1965 = (inp[3]) ? node1967 : 15'b000000111111111;
											assign node1967 = (inp[1]) ? 15'b000000001111111 : 15'b000000011111111;
										assign node1970 = (inp[0]) ? 15'b000000001111111 : node1971;
											assign node1971 = (inp[6]) ? 15'b000000001111111 : 15'b000000011111111;
								assign node1975 = (inp[9]) ? node1981 : node1976;
									assign node1976 = (inp[14]) ? node1978 : 15'b000000111111111;
										assign node1978 = (inp[3]) ? 15'b000000011111111 : 15'b000000001111111;
									assign node1981 = (inp[0]) ? 15'b000000000011111 : 15'b000000001111111;
							assign node1984 = (inp[6]) ? node2006 : node1985;
								assign node1985 = (inp[7]) ? node1995 : node1986;
									assign node1986 = (inp[14]) ? node1990 : node1987;
										assign node1987 = (inp[3]) ? 15'b000000001111111 : 15'b000000011111111;
										assign node1990 = (inp[3]) ? node1992 : 15'b000000001111111;
											assign node1992 = (inp[5]) ? 15'b000000001111111 : 15'b000000000111111;
									assign node1995 = (inp[9]) ? node1997 : 15'b000000011111111;
										assign node1997 = (inp[5]) ? node2001 : node1998;
											assign node1998 = (inp[11]) ? 15'b000000000111111 : 15'b000000001111111;
											assign node2001 = (inp[14]) ? 15'b000000000011111 : node2002;
												assign node2002 = (inp[11]) ? 15'b000000000111111 : 15'b000000000011111;
								assign node2006 = (inp[14]) ? node2016 : node2007;
									assign node2007 = (inp[3]) ? node2011 : node2008;
										assign node2008 = (inp[9]) ? 15'b000000000111111 : 15'b000000001111111;
										assign node2011 = (inp[9]) ? 15'b000000000011111 : node2012;
											assign node2012 = (inp[1]) ? 15'b000000000111111 : 15'b000000000011111;
									assign node2016 = (inp[0]) ? 15'b000000000111111 : node2017;
										assign node2017 = (inp[9]) ? 15'b000000000111111 : 15'b000000000011111;
						assign node2021 = (inp[12]) ? node2055 : node2022;
							assign node2022 = (inp[14]) ? node2028 : node2023;
								assign node2023 = (inp[1]) ? node2025 : 15'b000000001111111;
									assign node2025 = (inp[3]) ? 15'b000000000111111 : 15'b000000001111111;
								assign node2028 = (inp[9]) ? node2042 : node2029;
									assign node2029 = (inp[0]) ? node2035 : node2030;
										assign node2030 = (inp[5]) ? node2032 : 15'b000000000111111;
											assign node2032 = (inp[1]) ? 15'b000000000111111 : 15'b000000001111111;
										assign node2035 = (inp[6]) ? 15'b000000000001111 : node2036;
											assign node2036 = (inp[3]) ? 15'b000000000111111 : node2037;
												assign node2037 = (inp[1]) ? 15'b000000000011111 : 15'b000000000111111;
									assign node2042 = (inp[7]) ? node2052 : node2043;
										assign node2043 = (inp[5]) ? node2049 : node2044;
											assign node2044 = (inp[0]) ? node2046 : 15'b000000000111111;
												assign node2046 = (inp[6]) ? 15'b000000000011111 : 15'b000000000111111;
											assign node2049 = (inp[0]) ? 15'b000000000001111 : 15'b000000000011111;
										assign node2052 = (inp[1]) ? 15'b000000000000111 : 15'b000000000001111;
							assign node2055 = (inp[7]) ? node2069 : node2056;
								assign node2056 = (inp[3]) ? node2060 : node2057;
									assign node2057 = (inp[6]) ? 15'b000000000111111 : 15'b000000011111111;
									assign node2060 = (inp[6]) ? node2064 : node2061;
										assign node2061 = (inp[11]) ? 15'b000000000011111 : 15'b000000000111111;
										assign node2064 = (inp[14]) ? node2066 : 15'b000000000001111;
											assign node2066 = (inp[11]) ? 15'b000000000111111 : 15'b000000000011111;
								assign node2069 = (inp[1]) ? node2071 : 15'b000000000011111;
									assign node2071 = (inp[3]) ? 15'b000000000011111 : node2072;
										assign node2072 = (inp[5]) ? node2074 : 15'b000000000001111;
											assign node2074 = (inp[0]) ? 15'b000000000000011 : 15'b000000000000111;
					assign node2078 = (inp[11]) ? node2148 : node2079;
						assign node2079 = (inp[5]) ? node2107 : node2080;
							assign node2080 = (inp[6]) ? node2098 : node2081;
								assign node2081 = (inp[14]) ? node2087 : node2082;
									assign node2082 = (inp[2]) ? 15'b000000001111111 : node2083;
										assign node2083 = (inp[3]) ? 15'b000000011111111 : 15'b000000001111111;
									assign node2087 = (inp[3]) ? node2093 : node2088;
										assign node2088 = (inp[2]) ? 15'b000000001111111 : node2089;
											assign node2089 = (inp[12]) ? 15'b000000011111111 : 15'b000000111111111;
										assign node2093 = (inp[7]) ? node2095 : 15'b000000000111111;
											assign node2095 = (inp[1]) ? 15'b000000000001111 : 15'b000000000011111;
								assign node2098 = (inp[14]) ? node2104 : node2099;
									assign node2099 = (inp[0]) ? 15'b000000000111111 : node2100;
										assign node2100 = (inp[7]) ? 15'b000000000011111 : 15'b000000000111111;
									assign node2104 = (inp[1]) ? 15'b000000000001111 : 15'b000000001111111;
							assign node2107 = (inp[9]) ? node2131 : node2108;
								assign node2108 = (inp[7]) ? node2120 : node2109;
									assign node2109 = (inp[2]) ? node2117 : node2110;
										assign node2110 = (inp[14]) ? 15'b000000000111111 : node2111;
											assign node2111 = (inp[1]) ? node2113 : 15'b000000011111111;
												assign node2113 = (inp[0]) ? 15'b000000000111111 : 15'b000000001111111;
										assign node2117 = (inp[12]) ? 15'b000000000011111 : 15'b000000000111111;
									assign node2120 = (inp[0]) ? node2124 : node2121;
										assign node2121 = (inp[3]) ? 15'b000000000111111 : 15'b000000000011111;
										assign node2124 = (inp[6]) ? node2126 : 15'b000000000011111;
											assign node2126 = (inp[2]) ? 15'b000000000000111 : node2127;
												assign node2127 = (inp[12]) ? 15'b000000000001111 : 15'b000000000011111;
								assign node2131 = (inp[0]) ? node2137 : node2132;
									assign node2132 = (inp[6]) ? node2134 : 15'b000000000011111;
										assign node2134 = (inp[14]) ? 15'b000000000001111 : 15'b000000000011111;
									assign node2137 = (inp[2]) ? node2143 : node2138;
										assign node2138 = (inp[12]) ? node2140 : 15'b000000000011111;
											assign node2140 = (inp[14]) ? 15'b000000000000111 : 15'b000000000011111;
										assign node2143 = (inp[7]) ? node2145 : 15'b000000000000111;
											assign node2145 = (inp[12]) ? 15'b000000000000111 : 15'b000000000001111;
						assign node2148 = (inp[3]) ? node2180 : node2149;
							assign node2149 = (inp[0]) ? node2165 : node2150;
								assign node2150 = (inp[12]) ? 15'b000000000011111 : node2151;
									assign node2151 = (inp[9]) ? node2157 : node2152;
										assign node2152 = (inp[14]) ? node2154 : 15'b000000011111111;
											assign node2154 = (inp[7]) ? 15'b000000000111111 : 15'b000000001111111;
										assign node2157 = (inp[2]) ? node2161 : node2158;
											assign node2158 = (inp[1]) ? 15'b000000000111111 : 15'b000000001111111;
											assign node2161 = (inp[7]) ? 15'b000000000011111 : 15'b000000000001111;
								assign node2165 = (inp[1]) ? node2175 : node2166;
									assign node2166 = (inp[9]) ? node2170 : node2167;
										assign node2167 = (inp[5]) ? 15'b000000000111111 : 15'b000000011111111;
										assign node2170 = (inp[7]) ? 15'b000000000001111 : node2171;
											assign node2171 = (inp[14]) ? 15'b000000000011111 : 15'b000000000111111;
									assign node2175 = (inp[12]) ? 15'b000000000001111 : node2176;
										assign node2176 = (inp[5]) ? 15'b000000000001111 : 15'b000000000011111;
							assign node2180 = (inp[5]) ? node2204 : node2181;
								assign node2181 = (inp[7]) ? node2193 : node2182;
									assign node2182 = (inp[14]) ? node2186 : node2183;
										assign node2183 = (inp[2]) ? 15'b000000011111111 : 15'b000000000111111;
										assign node2186 = (inp[6]) ? node2188 : 15'b000000000011111;
											assign node2188 = (inp[9]) ? 15'b000000000001111 : node2189;
												assign node2189 = (inp[1]) ? 15'b000000000001111 : 15'b000000000011111;
									assign node2193 = (inp[9]) ? node2199 : node2194;
										assign node2194 = (inp[0]) ? node2196 : 15'b000000000001111;
											assign node2196 = (inp[1]) ? 15'b000000000011111 : 15'b000000000111111;
										assign node2199 = (inp[1]) ? node2201 : 15'b000000000001111;
											assign node2201 = (inp[12]) ? 15'b000000000000111 : 15'b000000000001111;
								assign node2204 = (inp[2]) ? node2214 : node2205;
									assign node2205 = (inp[0]) ? node2207 : 15'b000000000001111;
										assign node2207 = (inp[6]) ? node2211 : node2208;
											assign node2208 = (inp[14]) ? 15'b000000000000111 : 15'b000000000011111;
											assign node2211 = (inp[14]) ? 15'b000000000000111 : 15'b000000000000011;
									assign node2214 = (inp[14]) ? node2220 : node2215;
										assign node2215 = (inp[7]) ? 15'b000000000000111 : node2216;
											assign node2216 = (inp[6]) ? 15'b000000000000011 : 15'b000000000000111;
										assign node2220 = (inp[7]) ? 15'b000000000000111 : 15'b000000000011111;

endmodule