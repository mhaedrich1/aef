module dtc_split66_bm32 (
	input  wire [15-1:0] inp,
	output wire [9-1:0] outp
);

	wire [9-1:0] node1;
	wire [9-1:0] node2;
	wire [9-1:0] node5;
	wire [9-1:0] node6;
	wire [9-1:0] node7;
	wire [9-1:0] node9;
	wire [9-1:0] node11;
	wire [9-1:0] node12;
	wire [9-1:0] node14;
	wire [9-1:0] node18;
	wire [9-1:0] node21;
	wire [9-1:0] node22;
	wire [9-1:0] node24;
	wire [9-1:0] node26;
	wire [9-1:0] node29;
	wire [9-1:0] node30;
	wire [9-1:0] node31;
	wire [9-1:0] node34;
	wire [9-1:0] node35;
	wire [9-1:0] node37;
	wire [9-1:0] node41;
	wire [9-1:0] node43;
	wire [9-1:0] node45;
	wire [9-1:0] node48;
	wire [9-1:0] node49;
	wire [9-1:0] node50;
	wire [9-1:0] node51;
	wire [9-1:0] node52;
	wire [9-1:0] node53;
	wire [9-1:0] node54;
	wire [9-1:0] node55;
	wire [9-1:0] node60;
	wire [9-1:0] node61;
	wire [9-1:0] node62;
	wire [9-1:0] node63;
	wire [9-1:0] node68;
	wire [9-1:0] node71;
	wire [9-1:0] node72;
	wire [9-1:0] node73;
	wire [9-1:0] node74;
	wire [9-1:0] node79;
	wire [9-1:0] node80;
	wire [9-1:0] node81;
	wire [9-1:0] node82;
	wire [9-1:0] node87;
	wire [9-1:0] node90;
	wire [9-1:0] node91;
	wire [9-1:0] node92;
	wire [9-1:0] node93;
	wire [9-1:0] node94;
	wire [9-1:0] node99;
	wire [9-1:0] node100;
	wire [9-1:0] node101;
	wire [9-1:0] node102;
	wire [9-1:0] node107;
	wire [9-1:0] node110;
	wire [9-1:0] node111;
	wire [9-1:0] node112;
	wire [9-1:0] node113;
	wire [9-1:0] node114;
	wire [9-1:0] node116;
	wire [9-1:0] node118;
	wire [9-1:0] node121;
	wire [9-1:0] node123;
	wire [9-1:0] node126;
	wire [9-1:0] node127;
	wire [9-1:0] node128;
	wire [9-1:0] node132;
	wire [9-1:0] node133;
	wire [9-1:0] node134;
	wire [9-1:0] node139;
	wire [9-1:0] node140;
	wire [9-1:0] node143;
	wire [9-1:0] node146;
	wire [9-1:0] node147;
	wire [9-1:0] node148;
	wire [9-1:0] node149;
	wire [9-1:0] node150;
	wire [9-1:0] node153;
	wire [9-1:0] node156;
	wire [9-1:0] node157;
	wire [9-1:0] node158;
	wire [9-1:0] node163;
	wire [9-1:0] node164;
	wire [9-1:0] node166;
	wire [9-1:0] node168;
	wire [9-1:0] node171;
	wire [9-1:0] node173;
	wire [9-1:0] node176;
	wire [9-1:0] node177;
	wire [9-1:0] node180;
	wire [9-1:0] node183;
	wire [9-1:0] node184;
	wire [9-1:0] node185;
	wire [9-1:0] node186;
	wire [9-1:0] node187;
	wire [9-1:0] node188;
	wire [9-1:0] node193;
	wire [9-1:0] node194;
	wire [9-1:0] node195;
	wire [9-1:0] node196;
	wire [9-1:0] node201;
	wire [9-1:0] node204;
	wire [9-1:0] node205;
	wire [9-1:0] node206;
	wire [9-1:0] node207;
	wire [9-1:0] node212;
	wire [9-1:0] node213;
	wire [9-1:0] node214;
	wire [9-1:0] node215;
	wire [9-1:0] node220;
	wire [9-1:0] node223;
	wire [9-1:0] node224;
	wire [9-1:0] node225;
	wire [9-1:0] node226;
	wire [9-1:0] node227;
	wire [9-1:0] node232;
	wire [9-1:0] node233;
	wire [9-1:0] node234;
	wire [9-1:0] node235;
	wire [9-1:0] node240;
	wire [9-1:0] node243;
	wire [9-1:0] node244;
	wire [9-1:0] node245;
	wire [9-1:0] node246;
	wire [9-1:0] node247;
	wire [9-1:0] node248;
	wire [9-1:0] node249;
	wire [9-1:0] node253;
	wire [9-1:0] node254;
	wire [9-1:0] node255;
	wire [9-1:0] node260;
	wire [9-1:0] node261;
	wire [9-1:0] node262;
	wire [9-1:0] node265;
	wire [9-1:0] node268;
	wire [9-1:0] node269;
	wire [9-1:0] node270;
	wire [9-1:0] node275;
	wire [9-1:0] node277;
	wire [9-1:0] node280;
	wire [9-1:0] node281;
	wire [9-1:0] node282;
	wire [9-1:0] node283;
	wire [9-1:0] node285;
	wire [9-1:0] node287;
	wire [9-1:0] node290;
	wire [9-1:0] node292;
	wire [9-1:0] node295;
	wire [9-1:0] node296;
	wire [9-1:0] node298;
	wire [9-1:0] node300;
	wire [9-1:0] node303;
	wire [9-1:0] node305;
	wire [9-1:0] node308;
	wire [9-1:0] node310;
	wire [9-1:0] node313;
	wire [9-1:0] node314;
	wire [9-1:0] node315;
	wire [9-1:0] node316;
	wire [9-1:0] node317;
	wire [9-1:0] node319;
	wire [9-1:0] node321;
	wire [9-1:0] node324;
	wire [9-1:0] node326;
	wire [9-1:0] node329;
	wire [9-1:0] node330;
	wire [9-1:0] node331;
	wire [9-1:0] node332;
	wire [9-1:0] node336;
	wire [9-1:0] node337;
	wire [9-1:0] node341;
	wire [9-1:0] node342;
	wire [9-1:0] node343;
	wire [9-1:0] node348;
	wire [9-1:0] node350;
	wire [9-1:0] node353;
	wire [9-1:0] node354;
	wire [9-1:0] node355;
	wire [9-1:0] node356;
	wire [9-1:0] node358;
	wire [9-1:0] node360;
	wire [9-1:0] node363;
	wire [9-1:0] node365;
	wire [9-1:0] node368;
	wire [9-1:0] node369;
	wire [9-1:0] node371;
	wire [9-1:0] node373;
	wire [9-1:0] node376;
	wire [9-1:0] node378;
	wire [9-1:0] node381;
	wire [9-1:0] node382;
	wire [9-1:0] node385;
	wire [9-1:0] node388;
	wire [9-1:0] node389;
	wire [9-1:0] node390;
	wire [9-1:0] node391;
	wire [9-1:0] node393;
	wire [9-1:0] node396;
	wire [9-1:0] node397;
	wire [9-1:0] node400;
	wire [9-1:0] node401;
	wire [9-1:0] node404;
	wire [9-1:0] node405;
	wire [9-1:0] node408;
	wire [9-1:0] node411;
	wire [9-1:0] node412;
	wire [9-1:0] node414;
	wire [9-1:0] node417;
	wire [9-1:0] node418;
	wire [9-1:0] node421;
	wire [9-1:0] node422;
	wire [9-1:0] node425;
	wire [9-1:0] node426;
	wire [9-1:0] node429;
	wire [9-1:0] node432;
	wire [9-1:0] node433;
	wire [9-1:0] node434;
	wire [9-1:0] node435;
	wire [9-1:0] node438;
	wire [9-1:0] node440;
	wire [9-1:0] node443;
	wire [9-1:0] node444;
	wire [9-1:0] node447;
	wire [9-1:0] node449;
	wire [9-1:0] node450;
	wire [9-1:0] node453;
	wire [9-1:0] node456;
	wire [9-1:0] node457;
	wire [9-1:0] node458;
	wire [9-1:0] node461;
	wire [9-1:0] node464;
	wire [9-1:0] node465;
	wire [9-1:0] node468;
	wire [9-1:0] node469;
	wire [9-1:0] node470;
	wire [9-1:0] node473;
	wire [9-1:0] node474;
	wire [9-1:0] node477;
	wire [9-1:0] node480;
	wire [9-1:0] node481;
	wire [9-1:0] node484;
	wire [9-1:0] node485;
	wire [9-1:0] node488;

	assign outp = (inp[12]) ? node48 : node1;
		assign node1 = (inp[13]) ? node5 : node2;
			assign node2 = (inp[11]) ? 9'b101010101 : 9'b101010000;
			assign node5 = (inp[14]) ? node21 : node6;
				assign node6 = (inp[0]) ? node18 : node7;
					assign node7 = (inp[3]) ? node9 : 9'b101010001;
						assign node9 = (inp[8]) ? node11 : 9'b100010001;
							assign node11 = (inp[4]) ? 9'b100010001 : node12;
								assign node12 = (inp[9]) ? node14 : 9'b100010001;
									assign node14 = (inp[6]) ? 9'b001010001 : 9'b101010001;
					assign node18 = (inp[3]) ? 9'b000010101 : 9'b101010101;
				assign node21 = (inp[3]) ? node29 : node22;
					assign node22 = (inp[8]) ? node24 : 9'b111010101;
						assign node24 = (inp[9]) ? node26 : 9'b101010101;
							assign node26 = (inp[4]) ? 9'b111010101 : 9'b101010101;
					assign node29 = (inp[0]) ? node41 : node30;
						assign node30 = (inp[9]) ? node34 : node31;
							assign node31 = (inp[8]) ? 9'b101010111 : 9'b111010111;
							assign node34 = (inp[4]) ? 9'b111010111 : node35;
								assign node35 = (inp[8]) ? node37 : 9'b111010111;
									assign node37 = (inp[6]) ? 9'b011010101 : 9'b111010101;
						assign node41 = (inp[8]) ? node43 : 9'b011010111;
							assign node43 = (inp[9]) ? node45 : 9'b001010111;
								assign node45 = (inp[4]) ? 9'b001010101 : 9'b000010111;
		assign node48 = (inp[8]) ? node388 : node49;
			assign node49 = (inp[6]) ? node183 : node50;
				assign node50 = (inp[13]) ? node90 : node51;
					assign node51 = (inp[11]) ? node71 : node52;
						assign node52 = (inp[7]) ? node60 : node53;
							assign node53 = (inp[1]) ? 9'b111011000 : node54;
								assign node54 = (inp[9]) ? 9'b111011000 : node55;
									assign node55 = (inp[2]) ? 9'b111111000 : 9'b111110000;
							assign node60 = (inp[4]) ? node68 : node61;
								assign node61 = (inp[2]) ? 9'b111111000 : node62;
									assign node62 = (inp[9]) ? 9'b111111000 : node63;
										assign node63 = (inp[1]) ? 9'b111111000 : 9'b111110000;
								assign node68 = (inp[9]) ? 9'b111010000 : 9'b111110000;
						assign node71 = (inp[7]) ? node79 : node72;
							assign node72 = (inp[1]) ? 9'b111011100 : node73;
								assign node73 = (inp[9]) ? 9'b111011100 : node74;
									assign node74 = (inp[2]) ? 9'b111111100 : 9'b111110100;
							assign node79 = (inp[4]) ? node87 : node80;
								assign node80 = (inp[1]) ? 9'b111111100 : node81;
									assign node81 = (inp[2]) ? 9'b111111100 : node82;
										assign node82 = (inp[9]) ? 9'b111111100 : 9'b111110100;
								assign node87 = (inp[9]) ? 9'b111010100 : 9'b111110100;
					assign node90 = (inp[3]) ? node110 : node91;
						assign node91 = (inp[7]) ? node99 : node92;
							assign node92 = (inp[1]) ? 9'b111011100 : node93;
								assign node93 = (inp[9]) ? 9'b111011100 : node94;
									assign node94 = (inp[2]) ? 9'b111111100 : 9'b111110100;
							assign node99 = (inp[4]) ? node107 : node100;
								assign node100 = (inp[2]) ? 9'b111111100 : node101;
									assign node101 = (inp[9]) ? 9'b111111100 : node102;
										assign node102 = (inp[1]) ? 9'b111111100 : 9'b111110100;
								assign node107 = (inp[9]) ? 9'b111010100 : 9'b111110100;
						assign node110 = (inp[14]) ? node146 : node111;
							assign node111 = (inp[9]) ? node139 : node112;
								assign node112 = (inp[10]) ? node126 : node113;
									assign node113 = (inp[1]) ? node121 : node114;
										assign node114 = (inp[2]) ? node116 : 9'b110110100;
											assign node116 = (inp[7]) ? node118 : 9'b110111100;
												assign node118 = (inp[4]) ? 9'b110110100 : 9'b110111100;
										assign node121 = (inp[7]) ? node123 : 9'b110011100;
											assign node123 = (inp[4]) ? 9'b110110100 : 9'b110111100;
									assign node126 = (inp[7]) ? node132 : node127;
										assign node127 = (inp[1]) ? 9'b110011110 : node128;
											assign node128 = (inp[2]) ? 9'b110111110 : 9'b110110110;
										assign node132 = (inp[4]) ? 9'b110110110 : node133;
											assign node133 = (inp[2]) ? 9'b110111110 : node134;
												assign node134 = (inp[1]) ? 9'b110111110 : 9'b110110110;
								assign node139 = (inp[4]) ? node143 : node140;
									assign node140 = (inp[7]) ? 9'b110111110 : 9'b110011110;
									assign node143 = (inp[7]) ? 9'b110010110 : 9'b110011110;
							assign node146 = (inp[9]) ? node176 : node147;
								assign node147 = (inp[10]) ? node163 : node148;
									assign node148 = (inp[4]) ? node156 : node149;
										assign node149 = (inp[1]) ? node153 : node150;
											assign node150 = (inp[2]) ? 9'b111111100 : 9'b111110100;
											assign node153 = (inp[7]) ? 9'b111111100 : 9'b111011100;
										assign node156 = (inp[7]) ? 9'b111110100 : node157;
											assign node157 = (inp[1]) ? 9'b111011100 : node158;
												assign node158 = (inp[2]) ? 9'b111111100 : 9'b111110100;
									assign node163 = (inp[1]) ? node171 : node164;
										assign node164 = (inp[2]) ? node166 : 9'b111110110;
											assign node166 = (inp[7]) ? node168 : 9'b111111110;
												assign node168 = (inp[4]) ? 9'b111110110 : 9'b111111110;
										assign node171 = (inp[7]) ? node173 : 9'b111011110;
											assign node173 = (inp[4]) ? 9'b111110110 : 9'b111111110;
								assign node176 = (inp[4]) ? node180 : node177;
									assign node177 = (inp[7]) ? 9'b111111110 : 9'b111011110;
									assign node180 = (inp[7]) ? 9'b111010110 : 9'b111011110;
				assign node183 = (inp[13]) ? node223 : node184;
					assign node184 = (inp[11]) ? node204 : node185;
						assign node185 = (inp[7]) ? node193 : node186;
							assign node186 = (inp[1]) ? 9'b111011000 : node187;
								assign node187 = (inp[9]) ? 9'b111011000 : node188;
									assign node188 = (inp[2]) ? 9'b111111000 : 9'b111110000;
							assign node193 = (inp[4]) ? node201 : node194;
								assign node194 = (inp[2]) ? 9'b111111000 : node195;
									assign node195 = (inp[1]) ? 9'b111111000 : node196;
										assign node196 = (inp[9]) ? 9'b111111000 : 9'b111110000;
								assign node201 = (inp[9]) ? 9'b111010000 : 9'b111110000;
						assign node204 = (inp[7]) ? node212 : node205;
							assign node205 = (inp[9]) ? 9'b111011101 : node206;
								assign node206 = (inp[1]) ? 9'b111011101 : node207;
									assign node207 = (inp[2]) ? 9'b111111101 : 9'b111110101;
							assign node212 = (inp[4]) ? node220 : node213;
								assign node213 = (inp[9]) ? 9'b111111101 : node214;
									assign node214 = (inp[1]) ? 9'b111111101 : node215;
										assign node215 = (inp[2]) ? 9'b111111101 : 9'b111110101;
								assign node220 = (inp[9]) ? 9'b111010101 : 9'b111110101;
					assign node223 = (inp[3]) ? node243 : node224;
						assign node224 = (inp[7]) ? node232 : node225;
							assign node225 = (inp[1]) ? 9'b111011101 : node226;
								assign node226 = (inp[9]) ? 9'b111011101 : node227;
									assign node227 = (inp[2]) ? 9'b111111101 : 9'b111110101;
							assign node232 = (inp[4]) ? node240 : node233;
								assign node233 = (inp[2]) ? 9'b111111101 : node234;
									assign node234 = (inp[1]) ? 9'b111111101 : node235;
										assign node235 = (inp[9]) ? 9'b111111101 : 9'b111110101;
								assign node240 = (inp[9]) ? 9'b111010101 : 9'b111110101;
						assign node243 = (inp[14]) ? node313 : node244;
							assign node244 = (inp[5]) ? node280 : node245;
								assign node245 = (inp[9]) ? node275 : node246;
									assign node246 = (inp[10]) ? node260 : node247;
										assign node247 = (inp[7]) ? node253 : node248;
											assign node248 = (inp[1]) ? 9'b110001101 : node249;
												assign node249 = (inp[2]) ? 9'b110101101 : 9'b110100101;
											assign node253 = (inp[4]) ? 9'b110100101 : node254;
												assign node254 = (inp[2]) ? 9'b110101101 : node255;
													assign node255 = (inp[1]) ? 9'b110101101 : 9'b110100101;
										assign node260 = (inp[4]) ? node268 : node261;
											assign node261 = (inp[1]) ? node265 : node262;
												assign node262 = (inp[2]) ? 9'b110101111 : 9'b110100111;
												assign node265 = (inp[7]) ? 9'b110101111 : 9'b110001111;
											assign node268 = (inp[7]) ? 9'b110100111 : node269;
												assign node269 = (inp[1]) ? 9'b110001111 : node270;
													assign node270 = (inp[2]) ? 9'b110101111 : 9'b110100111;
									assign node275 = (inp[7]) ? node277 : 9'b110001111;
										assign node277 = (inp[4]) ? 9'b110000111 : 9'b110101111;
								assign node280 = (inp[9]) ? node308 : node281;
									assign node281 = (inp[10]) ? node295 : node282;
										assign node282 = (inp[1]) ? node290 : node283;
											assign node283 = (inp[2]) ? node285 : 9'b110110101;
												assign node285 = (inp[7]) ? node287 : 9'b110111101;
													assign node287 = (inp[4]) ? 9'b110110101 : 9'b110111101;
											assign node290 = (inp[7]) ? node292 : 9'b110011101;
												assign node292 = (inp[4]) ? 9'b110110101 : 9'b110111101;
										assign node295 = (inp[1]) ? node303 : node296;
											assign node296 = (inp[2]) ? node298 : 9'b110110111;
												assign node298 = (inp[7]) ? node300 : 9'b110111111;
													assign node300 = (inp[4]) ? 9'b110110111 : 9'b110111111;
											assign node303 = (inp[7]) ? node305 : 9'b110011111;
												assign node305 = (inp[4]) ? 9'b110110111 : 9'b110111111;
									assign node308 = (inp[7]) ? node310 : 9'b110011111;
										assign node310 = (inp[4]) ? 9'b110010111 : 9'b110111111;
							assign node313 = (inp[5]) ? node353 : node314;
								assign node314 = (inp[9]) ? node348 : node315;
									assign node315 = (inp[10]) ? node329 : node316;
										assign node316 = (inp[1]) ? node324 : node317;
											assign node317 = (inp[2]) ? node319 : 9'b111100101;
												assign node319 = (inp[7]) ? node321 : 9'b111101101;
													assign node321 = (inp[4]) ? 9'b111100101 : 9'b111101101;
											assign node324 = (inp[7]) ? node326 : 9'b111001101;
												assign node326 = (inp[4]) ? 9'b111100101 : 9'b111101101;
										assign node329 = (inp[4]) ? node341 : node330;
											assign node330 = (inp[7]) ? node336 : node331;
												assign node331 = (inp[1]) ? 9'b111001111 : node332;
													assign node332 = (inp[2]) ? 9'b111101111 : 9'b111100111;
												assign node336 = (inp[1]) ? 9'b111101111 : node337;
													assign node337 = (inp[2]) ? 9'b111101111 : 9'b111100111;
											assign node341 = (inp[7]) ? 9'b111100111 : node342;
												assign node342 = (inp[1]) ? 9'b111001111 : node343;
													assign node343 = (inp[2]) ? 9'b111101111 : 9'b111100111;
									assign node348 = (inp[7]) ? node350 : 9'b111001111;
										assign node350 = (inp[4]) ? 9'b111000111 : 9'b111101111;
								assign node353 = (inp[9]) ? node381 : node354;
									assign node354 = (inp[10]) ? node368 : node355;
										assign node355 = (inp[1]) ? node363 : node356;
											assign node356 = (inp[2]) ? node358 : 9'b111110101;
												assign node358 = (inp[4]) ? node360 : 9'b111111101;
													assign node360 = (inp[7]) ? 9'b111110101 : 9'b111111101;
											assign node363 = (inp[7]) ? node365 : 9'b111011101;
												assign node365 = (inp[4]) ? 9'b111110101 : 9'b111111101;
										assign node368 = (inp[1]) ? node376 : node369;
											assign node369 = (inp[2]) ? node371 : 9'b111110111;
												assign node371 = (inp[7]) ? node373 : 9'b111111111;
													assign node373 = (inp[4]) ? 9'b111110111 : 9'b111111111;
											assign node376 = (inp[7]) ? node378 : 9'b111011111;
												assign node378 = (inp[4]) ? 9'b111110111 : 9'b111111111;
									assign node381 = (inp[4]) ? node385 : node382;
										assign node382 = (inp[7]) ? 9'b111111111 : 9'b111011111;
										assign node385 = (inp[7]) ? 9'b111010111 : 9'b111011111;
			assign node388 = (inp[9]) ? node432 : node389;
				assign node389 = (inp[4]) ? node411 : node390;
					assign node390 = (inp[13]) ? node396 : node391;
						assign node391 = (inp[11]) ? node393 : 9'b101111000;
							assign node393 = (inp[6]) ? 9'b101111101 : 9'b101111100;
						assign node396 = (inp[3]) ? node400 : node397;
							assign node397 = (inp[6]) ? 9'b101111101 : 9'b101111100;
							assign node400 = (inp[6]) ? node404 : node401;
								assign node401 = (inp[14]) ? 9'b101111110 : 9'b100111110;
								assign node404 = (inp[14]) ? node408 : node405;
									assign node405 = (inp[5]) ? 9'b100111111 : 9'b100101111;
									assign node408 = (inp[5]) ? 9'b101111111 : 9'b101101111;
					assign node411 = (inp[13]) ? node417 : node412;
						assign node412 = (inp[11]) ? node414 : 9'b101010000;
							assign node414 = (inp[6]) ? 9'b101010101 : 9'b101010100;
						assign node417 = (inp[3]) ? node421 : node418;
							assign node418 = (inp[6]) ? 9'b101010101 : 9'b101010100;
							assign node421 = (inp[6]) ? node425 : node422;
								assign node422 = (inp[14]) ? 9'b101010110 : 9'b100010110;
								assign node425 = (inp[14]) ? node429 : node426;
									assign node426 = (inp[5]) ? 9'b100010111 : 9'b100000111;
									assign node429 = (inp[5]) ? 9'b101010111 : 9'b101000111;
				assign node432 = (inp[6]) ? node456 : node433;
					assign node433 = (inp[4]) ? node443 : node434;
						assign node434 = (inp[13]) ? node438 : node435;
							assign node435 = (inp[11]) ? 9'b101010100 : 9'b101010000;
							assign node438 = (inp[3]) ? node440 : 9'b101010100;
								assign node440 = (inp[0]) ? 9'b100010110 : 9'b111010100;
						assign node443 = (inp[13]) ? node447 : node444;
							assign node444 = (inp[11]) ? 9'b111010100 : 9'b111010000;
							assign node447 = (inp[3]) ? node449 : 9'b111010100;
								assign node449 = (inp[0]) ? node453 : node450;
									assign node450 = (inp[14]) ? 9'b111010110 : 9'b110010110;
									assign node453 = (inp[14]) ? 9'b101010100 : 9'b100010100;
					assign node456 = (inp[13]) ? node464 : node457;
						assign node457 = (inp[11]) ? node461 : node458;
							assign node458 = (inp[4]) ? 9'b111010000 : 9'b101010000;
							assign node461 = (inp[4]) ? 9'b111010101 : 9'b101010101;
						assign node464 = (inp[3]) ? node468 : node465;
							assign node465 = (inp[4]) ? 9'b111010101 : 9'b101010101;
							assign node468 = (inp[0]) ? node480 : node469;
								assign node469 = (inp[4]) ? node473 : node470;
									assign node470 = (inp[5]) ? 9'b011010101 : 9'b011000101;
									assign node473 = (inp[5]) ? node477 : node474;
										assign node474 = (inp[14]) ? 9'b111000111 : 9'b110000111;
										assign node477 = (inp[14]) ? 9'b111010111 : 9'b110010111;
								assign node480 = (inp[4]) ? node484 : node481;
									assign node481 = (inp[5]) ? 9'b100010111 : 9'b100000111;
									assign node484 = (inp[5]) ? node488 : node485;
										assign node485 = (inp[14]) ? 9'b101000101 : 9'b100000101;
										assign node488 = (inp[14]) ? 9'b101010101 : 9'b100010101;

endmodule