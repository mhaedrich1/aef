module dtc_split5_bm21 (
	input  wire [10-1:0] inp,
	output wire [10-1:0] outp
);

	wire [10-1:0] node1;
	wire [10-1:0] node2;
	wire [10-1:0] node3;
	wire [10-1:0] node4;
	wire [10-1:0] node5;
	wire [10-1:0] node6;
	wire [10-1:0] node7;
	wire [10-1:0] node10;
	wire [10-1:0] node13;
	wire [10-1:0] node14;
	wire [10-1:0] node17;
	wire [10-1:0] node20;
	wire [10-1:0] node21;
	wire [10-1:0] node22;
	wire [10-1:0] node25;
	wire [10-1:0] node28;
	wire [10-1:0] node29;
	wire [10-1:0] node32;
	wire [10-1:0] node35;
	wire [10-1:0] node36;
	wire [10-1:0] node37;
	wire [10-1:0] node39;
	wire [10-1:0] node42;
	wire [10-1:0] node43;
	wire [10-1:0] node46;
	wire [10-1:0] node49;
	wire [10-1:0] node50;
	wire [10-1:0] node51;
	wire [10-1:0] node54;
	wire [10-1:0] node57;
	wire [10-1:0] node58;
	wire [10-1:0] node61;
	wire [10-1:0] node64;
	wire [10-1:0] node65;
	wire [10-1:0] node66;
	wire [10-1:0] node67;
	wire [10-1:0] node68;
	wire [10-1:0] node71;
	wire [10-1:0] node74;
	wire [10-1:0] node75;
	wire [10-1:0] node78;
	wire [10-1:0] node81;
	wire [10-1:0] node82;
	wire [10-1:0] node83;
	wire [10-1:0] node86;
	wire [10-1:0] node89;
	wire [10-1:0] node90;
	wire [10-1:0] node93;
	wire [10-1:0] node96;
	wire [10-1:0] node97;
	wire [10-1:0] node98;
	wire [10-1:0] node99;
	wire [10-1:0] node102;
	wire [10-1:0] node105;
	wire [10-1:0] node106;
	wire [10-1:0] node109;
	wire [10-1:0] node112;
	wire [10-1:0] node113;
	wire [10-1:0] node115;
	wire [10-1:0] node118;
	wire [10-1:0] node119;
	wire [10-1:0] node122;
	wire [10-1:0] node125;
	wire [10-1:0] node126;
	wire [10-1:0] node127;
	wire [10-1:0] node128;
	wire [10-1:0] node129;
	wire [10-1:0] node130;
	wire [10-1:0] node133;
	wire [10-1:0] node136;
	wire [10-1:0] node137;
	wire [10-1:0] node140;
	wire [10-1:0] node143;
	wire [10-1:0] node144;
	wire [10-1:0] node146;
	wire [10-1:0] node149;
	wire [10-1:0] node150;
	wire [10-1:0] node153;
	wire [10-1:0] node156;
	wire [10-1:0] node157;
	wire [10-1:0] node158;
	wire [10-1:0] node159;
	wire [10-1:0] node162;
	wire [10-1:0] node165;
	wire [10-1:0] node166;
	wire [10-1:0] node169;
	wire [10-1:0] node172;
	wire [10-1:0] node173;
	wire [10-1:0] node174;
	wire [10-1:0] node177;
	wire [10-1:0] node180;
	wire [10-1:0] node181;
	wire [10-1:0] node184;
	wire [10-1:0] node187;
	wire [10-1:0] node188;
	wire [10-1:0] node189;
	wire [10-1:0] node190;
	wire [10-1:0] node191;
	wire [10-1:0] node194;
	wire [10-1:0] node197;
	wire [10-1:0] node198;
	wire [10-1:0] node201;
	wire [10-1:0] node204;
	wire [10-1:0] node205;
	wire [10-1:0] node206;
	wire [10-1:0] node209;
	wire [10-1:0] node212;
	wire [10-1:0] node213;
	wire [10-1:0] node216;
	wire [10-1:0] node219;
	wire [10-1:0] node220;
	wire [10-1:0] node221;
	wire [10-1:0] node222;
	wire [10-1:0] node225;
	wire [10-1:0] node228;
	wire [10-1:0] node229;
	wire [10-1:0] node232;
	wire [10-1:0] node235;
	wire [10-1:0] node236;
	wire [10-1:0] node237;
	wire [10-1:0] node240;
	wire [10-1:0] node243;
	wire [10-1:0] node244;
	wire [10-1:0] node247;
	wire [10-1:0] node250;
	wire [10-1:0] node251;
	wire [10-1:0] node252;
	wire [10-1:0] node253;
	wire [10-1:0] node254;
	wire [10-1:0] node255;
	wire [10-1:0] node256;
	wire [10-1:0] node259;
	wire [10-1:0] node262;
	wire [10-1:0] node263;
	wire [10-1:0] node266;
	wire [10-1:0] node269;
	wire [10-1:0] node270;
	wire [10-1:0] node271;
	wire [10-1:0] node274;
	wire [10-1:0] node277;
	wire [10-1:0] node278;
	wire [10-1:0] node281;
	wire [10-1:0] node284;
	wire [10-1:0] node285;
	wire [10-1:0] node286;
	wire [10-1:0] node287;
	wire [10-1:0] node290;
	wire [10-1:0] node293;
	wire [10-1:0] node294;
	wire [10-1:0] node297;
	wire [10-1:0] node300;
	wire [10-1:0] node301;
	wire [10-1:0] node302;
	wire [10-1:0] node305;
	wire [10-1:0] node308;
	wire [10-1:0] node309;
	wire [10-1:0] node313;
	wire [10-1:0] node314;
	wire [10-1:0] node315;
	wire [10-1:0] node316;
	wire [10-1:0] node317;
	wire [10-1:0] node320;
	wire [10-1:0] node323;
	wire [10-1:0] node324;
	wire [10-1:0] node327;
	wire [10-1:0] node330;
	wire [10-1:0] node331;
	wire [10-1:0] node332;
	wire [10-1:0] node335;
	wire [10-1:0] node338;
	wire [10-1:0] node339;
	wire [10-1:0] node342;
	wire [10-1:0] node345;
	wire [10-1:0] node346;
	wire [10-1:0] node347;
	wire [10-1:0] node348;
	wire [10-1:0] node351;
	wire [10-1:0] node354;
	wire [10-1:0] node355;
	wire [10-1:0] node358;
	wire [10-1:0] node361;
	wire [10-1:0] node362;
	wire [10-1:0] node364;
	wire [10-1:0] node367;
	wire [10-1:0] node368;
	wire [10-1:0] node371;
	wire [10-1:0] node374;
	wire [10-1:0] node375;
	wire [10-1:0] node376;
	wire [10-1:0] node377;
	wire [10-1:0] node378;
	wire [10-1:0] node379;
	wire [10-1:0] node382;
	wire [10-1:0] node385;
	wire [10-1:0] node386;
	wire [10-1:0] node389;
	wire [10-1:0] node392;
	wire [10-1:0] node393;
	wire [10-1:0] node395;
	wire [10-1:0] node398;
	wire [10-1:0] node399;
	wire [10-1:0] node402;
	wire [10-1:0] node405;
	wire [10-1:0] node406;
	wire [10-1:0] node407;
	wire [10-1:0] node409;
	wire [10-1:0] node412;
	wire [10-1:0] node413;
	wire [10-1:0] node416;
	wire [10-1:0] node419;
	wire [10-1:0] node420;
	wire [10-1:0] node421;
	wire [10-1:0] node424;
	wire [10-1:0] node427;
	wire [10-1:0] node428;
	wire [10-1:0] node431;
	wire [10-1:0] node434;
	wire [10-1:0] node435;
	wire [10-1:0] node436;
	wire [10-1:0] node437;
	wire [10-1:0] node438;
	wire [10-1:0] node441;
	wire [10-1:0] node444;
	wire [10-1:0] node445;
	wire [10-1:0] node448;
	wire [10-1:0] node451;
	wire [10-1:0] node452;
	wire [10-1:0] node453;
	wire [10-1:0] node456;
	wire [10-1:0] node459;
	wire [10-1:0] node461;
	wire [10-1:0] node464;
	wire [10-1:0] node465;
	wire [10-1:0] node466;
	wire [10-1:0] node468;
	wire [10-1:0] node471;
	wire [10-1:0] node472;
	wire [10-1:0] node475;
	wire [10-1:0] node478;
	wire [10-1:0] node479;
	wire [10-1:0] node480;
	wire [10-1:0] node483;
	wire [10-1:0] node486;
	wire [10-1:0] node487;
	wire [10-1:0] node490;

	assign outp = (inp[3]) ? node250 : node1;
		assign node1 = (inp[4]) ? node125 : node2;
			assign node2 = (inp[2]) ? node64 : node3;
				assign node3 = (inp[5]) ? node35 : node4;
					assign node4 = (inp[6]) ? node20 : node5;
						assign node5 = (inp[1]) ? node13 : node6;
							assign node6 = (inp[9]) ? node10 : node7;
								assign node7 = (inp[0]) ? 10'b0011111111 : 10'b0111111111;
								assign node10 = (inp[8]) ? 10'b0001111111 : 10'b0011111111;
							assign node13 = (inp[0]) ? node17 : node14;
								assign node14 = (inp[9]) ? 10'b0001111111 : 10'b0011111111;
								assign node17 = (inp[7]) ? 10'b0000111111 : 10'b0001111111;
						assign node20 = (inp[9]) ? node28 : node21;
							assign node21 = (inp[7]) ? node25 : node22;
								assign node22 = (inp[0]) ? 10'b0001111111 : 10'b0011111111;
								assign node25 = (inp[8]) ? 10'b0000111111 : 10'b0001111111;
							assign node28 = (inp[8]) ? node32 : node29;
								assign node29 = (inp[7]) ? 10'b0000011111 : 10'b0001111111;
								assign node32 = (inp[1]) ? 10'b0000011111 : 10'b0000111111;
					assign node35 = (inp[0]) ? node49 : node36;
						assign node36 = (inp[8]) ? node42 : node37;
							assign node37 = (inp[9]) ? node39 : 10'b0011111111;
								assign node39 = (inp[7]) ? 10'b0000111111 : 10'b0001111111;
							assign node42 = (inp[9]) ? node46 : node43;
								assign node43 = (inp[1]) ? 10'b0000111111 : 10'b0001111111;
								assign node46 = (inp[6]) ? 10'b0000011111 : 10'b0000111111;
						assign node49 = (inp[7]) ? node57 : node50;
							assign node50 = (inp[9]) ? node54 : node51;
								assign node51 = (inp[8]) ? 10'b0000111111 : 10'b0001111111;
								assign node54 = (inp[8]) ? 10'b0000011111 : 10'b0000111111;
							assign node57 = (inp[8]) ? node61 : node58;
								assign node58 = (inp[1]) ? 10'b0000011111 : 10'b0000111111;
								assign node61 = (inp[9]) ? 10'b0000011111 : 10'b0000001111;
				assign node64 = (inp[8]) ? node96 : node65;
					assign node65 = (inp[1]) ? node81 : node66;
						assign node66 = (inp[0]) ? node74 : node67;
							assign node67 = (inp[5]) ? node71 : node68;
								assign node68 = (inp[7]) ? 10'b0001111111 : 10'b0011111111;
								assign node71 = (inp[6]) ? 10'b0000111111 : 10'b0001111111;
							assign node74 = (inp[9]) ? node78 : node75;
								assign node75 = (inp[6]) ? 10'b0000111111 : 10'b0001111111;
								assign node78 = (inp[6]) ? 10'b0000001111 : 10'b0000111111;
						assign node81 = (inp[0]) ? node89 : node82;
							assign node82 = (inp[9]) ? node86 : node83;
								assign node83 = (inp[7]) ? 10'b0000111111 : 10'b0011111111;
								assign node86 = (inp[6]) ? 10'b0000011111 : 10'b0000111111;
							assign node89 = (inp[5]) ? node93 : node90;
								assign node90 = (inp[9]) ? 10'b0000001111 : 10'b0000111111;
								assign node93 = (inp[6]) ? 10'b0000001111 : 10'b0000011111;
					assign node96 = (inp[7]) ? node112 : node97;
						assign node97 = (inp[9]) ? node105 : node98;
							assign node98 = (inp[1]) ? node102 : node99;
								assign node99 = (inp[0]) ? 10'b0000111111 : 10'b0001111111;
								assign node102 = (inp[0]) ? 10'b0000011111 : 10'b0000111111;
							assign node105 = (inp[5]) ? node109 : node106;
								assign node106 = (inp[1]) ? 10'b0000011111 : 10'b0000011111;
								assign node109 = (inp[0]) ? 10'b0000000111 : 10'b0000011111;
						assign node112 = (inp[6]) ? node118 : node113;
							assign node113 = (inp[9]) ? node115 : 10'b0000111111;
								assign node115 = (inp[5]) ? 10'b0000001111 : 10'b0000011111;
							assign node118 = (inp[5]) ? node122 : node119;
								assign node119 = (inp[9]) ? 10'b0000000111 : 10'b0000011111;
								assign node122 = (inp[0]) ? 10'b0000000111 : 10'b0000001111;
			assign node125 = (inp[6]) ? node187 : node126;
				assign node126 = (inp[8]) ? node156 : node127;
					assign node127 = (inp[7]) ? node143 : node128;
						assign node128 = (inp[0]) ? node136 : node129;
							assign node129 = (inp[1]) ? node133 : node130;
								assign node130 = (inp[5]) ? 10'b0001111111 : 10'b0011111111;
								assign node133 = (inp[9]) ? 10'b0000111111 : 10'b0001111111;
							assign node136 = (inp[5]) ? node140 : node137;
								assign node137 = (inp[1]) ? 10'b0000111111 : 10'b0001111111;
								assign node140 = (inp[1]) ? 10'b0000001111 : 10'b0000011111;
						assign node143 = (inp[9]) ? node149 : node144;
							assign node144 = (inp[2]) ? node146 : 10'b0000111111;
								assign node146 = (inp[1]) ? 10'b0000011111 : 10'b0000111111;
							assign node149 = (inp[1]) ? node153 : node150;
								assign node150 = (inp[5]) ? 10'b0000011111 : 10'b0000111111;
								assign node153 = (inp[5]) ? 10'b0000001111 : 10'b0000011111;
					assign node156 = (inp[1]) ? node172 : node157;
						assign node157 = (inp[5]) ? node165 : node158;
							assign node158 = (inp[0]) ? node162 : node159;
								assign node159 = (inp[9]) ? 10'b0000111111 : 10'b0001111111;
								assign node162 = (inp[2]) ? 10'b0000011111 : 10'b0000111111;
							assign node165 = (inp[0]) ? node169 : node166;
								assign node166 = (inp[2]) ? 10'b0000011111 : 10'b0000111111;
								assign node169 = (inp[2]) ? 10'b0000001111 : 10'b0000011111;
						assign node172 = (inp[9]) ? node180 : node173;
							assign node173 = (inp[0]) ? node177 : node174;
								assign node174 = (inp[2]) ? 10'b0000011111 : 10'b0000111111;
								assign node177 = (inp[5]) ? 10'b0000001111 : 10'b0000011111;
							assign node180 = (inp[7]) ? node184 : node181;
								assign node181 = (inp[5]) ? 10'b0000001111 : 10'b0000011111;
								assign node184 = (inp[0]) ? 10'b0000000111 : 10'b0000001111;
				assign node187 = (inp[0]) ? node219 : node188;
					assign node188 = (inp[7]) ? node204 : node189;
						assign node189 = (inp[5]) ? node197 : node190;
							assign node190 = (inp[1]) ? node194 : node191;
								assign node191 = (inp[9]) ? 10'b0000111111 : 10'b0001111111;
								assign node194 = (inp[2]) ? 10'b0000011111 : 10'b0000011111;
							assign node197 = (inp[1]) ? node201 : node198;
								assign node198 = (inp[8]) ? 10'b0000011111 : 10'b0000111111;
								assign node201 = (inp[8]) ? 10'b0000001111 : 10'b0000011111;
						assign node204 = (inp[2]) ? node212 : node205;
							assign node205 = (inp[1]) ? node209 : node206;
								assign node206 = (inp[5]) ? 10'b0000011111 : 10'b0000011111;
								assign node209 = (inp[8]) ? 10'b0000011111 : 10'b0000001111;
							assign node212 = (inp[8]) ? node216 : node213;
								assign node213 = (inp[5]) ? 10'b0000001111 : 10'b0000011111;
								assign node216 = (inp[5]) ? 10'b0000000111 : 10'b0000001111;
					assign node219 = (inp[5]) ? node235 : node220;
						assign node220 = (inp[7]) ? node228 : node221;
							assign node221 = (inp[2]) ? node225 : node222;
								assign node222 = (inp[9]) ? 10'b0000011111 : 10'b0000111111;
								assign node225 = (inp[9]) ? 10'b0000001111 : 10'b0000001111;
							assign node228 = (inp[8]) ? node232 : node229;
								assign node229 = (inp[1]) ? 10'b0000001111 : 10'b0000011111;
								assign node232 = (inp[9]) ? 10'b0000000111 : 10'b0000001111;
						assign node235 = (inp[2]) ? node243 : node236;
							assign node236 = (inp[9]) ? node240 : node237;
								assign node237 = (inp[7]) ? 10'b0000001111 : 10'b0000001111;
								assign node240 = (inp[1]) ? 10'b0000000111 : 10'b0000001111;
							assign node243 = (inp[7]) ? node247 : node244;
								assign node244 = (inp[9]) ? 10'b0000000111 : 10'b0000001111;
								assign node247 = (inp[8]) ? 10'b0000000011 : 10'b0000000111;
		assign node250 = (inp[1]) ? node374 : node251;
			assign node251 = (inp[5]) ? node313 : node252;
				assign node252 = (inp[8]) ? node284 : node253;
					assign node253 = (inp[4]) ? node269 : node254;
						assign node254 = (inp[0]) ? node262 : node255;
							assign node255 = (inp[6]) ? node259 : node256;
								assign node256 = (inp[9]) ? 10'b0001111111 : 10'b0011111111;
								assign node259 = (inp[9]) ? 10'b0000111111 : 10'b0001111111;
							assign node262 = (inp[6]) ? node266 : node263;
								assign node263 = (inp[7]) ? 10'b0000111111 : 10'b0001111111;
								assign node266 = (inp[9]) ? 10'b0000011111 : 10'b0000111111;
						assign node269 = (inp[2]) ? node277 : node270;
							assign node270 = (inp[6]) ? node274 : node271;
								assign node271 = (inp[7]) ? 10'b0000111111 : 10'b0001111111;
								assign node274 = (inp[9]) ? 10'b0000011111 : 10'b0000111111;
							assign node277 = (inp[0]) ? node281 : node278;
								assign node278 = (inp[6]) ? 10'b0000011111 : 10'b0000011111;
								assign node281 = (inp[7]) ? 10'b0000001111 : 10'b0000011111;
					assign node284 = (inp[0]) ? node300 : node285;
						assign node285 = (inp[6]) ? node293 : node286;
							assign node286 = (inp[2]) ? node290 : node287;
								assign node287 = (inp[9]) ? 10'b0000111111 : 10'b0001111111;
								assign node290 = (inp[9]) ? 10'b0000001111 : 10'b0000111111;
							assign node293 = (inp[4]) ? node297 : node294;
								assign node294 = (inp[9]) ? 10'b0000011111 : 10'b0000111111;
								assign node297 = (inp[2]) ? 10'b0000000111 : 10'b0000011111;
						assign node300 = (inp[4]) ? node308 : node301;
							assign node301 = (inp[9]) ? node305 : node302;
								assign node302 = (inp[7]) ? 10'b0000011111 : 10'b0000011111;
								assign node305 = (inp[2]) ? 10'b0000001111 : 10'b0000011111;
							assign node308 = (inp[7]) ? 10'b0000000111 : node309;
								assign node309 = (inp[6]) ? 10'b0000000111 : 10'b0000011111;
				assign node313 = (inp[2]) ? node345 : node314;
					assign node314 = (inp[0]) ? node330 : node315;
						assign node315 = (inp[4]) ? node323 : node316;
							assign node316 = (inp[8]) ? node320 : node317;
								assign node317 = (inp[6]) ? 10'b0000111111 : 10'b0001111111;
								assign node320 = (inp[9]) ? 10'b0000011111 : 10'b0000111111;
							assign node323 = (inp[6]) ? node327 : node324;
								assign node324 = (inp[9]) ? 10'b0000011111 : 10'b0000111111;
								assign node327 = (inp[7]) ? 10'b0000001111 : 10'b0000011111;
						assign node330 = (inp[4]) ? node338 : node331;
							assign node331 = (inp[9]) ? node335 : node332;
								assign node332 = (inp[8]) ? 10'b0000011111 : 10'b0001111111;
								assign node335 = (inp[6]) ? 10'b0000001111 : 10'b0000011111;
							assign node338 = (inp[7]) ? node342 : node339;
								assign node339 = (inp[6]) ? 10'b0000001111 : 10'b0000001111;
								assign node342 = (inp[8]) ? 10'b0000000111 : 10'b0000001111;
					assign node345 = (inp[6]) ? node361 : node346;
						assign node346 = (inp[8]) ? node354 : node347;
							assign node347 = (inp[7]) ? node351 : node348;
								assign node348 = (inp[4]) ? 10'b0000011111 : 10'b0000111111;
								assign node351 = (inp[4]) ? 10'b0000001111 : 10'b0000011111;
							assign node354 = (inp[7]) ? node358 : node355;
								assign node355 = (inp[9]) ? 10'b0000001111 : 10'b0000011111;
								assign node358 = (inp[4]) ? 10'b0000000111 : 10'b0000001111;
						assign node361 = (inp[9]) ? node367 : node362;
							assign node362 = (inp[8]) ? node364 : 10'b0000001111;
								assign node364 = (inp[0]) ? 10'b0000000111 : 10'b0000001111;
							assign node367 = (inp[0]) ? node371 : node368;
								assign node368 = (inp[8]) ? 10'b0000000111 : 10'b0000001111;
								assign node371 = (inp[8]) ? 10'b0000000011 : 10'b0000000011;
			assign node374 = (inp[7]) ? node434 : node375;
				assign node375 = (inp[2]) ? node405 : node376;
					assign node376 = (inp[0]) ? node392 : node377;
						assign node377 = (inp[5]) ? node385 : node378;
							assign node378 = (inp[4]) ? node382 : node379;
								assign node379 = (inp[8]) ? 10'b0000111111 : 10'b0001111111;
								assign node382 = (inp[9]) ? 10'b0000011111 : 10'b0000111111;
							assign node385 = (inp[8]) ? node389 : node386;
								assign node386 = (inp[6]) ? 10'b0000011111 : 10'b0000111111;
								assign node389 = (inp[4]) ? 10'b0000001111 : 10'b0000011111;
						assign node392 = (inp[9]) ? node398 : node393;
							assign node393 = (inp[6]) ? node395 : 10'b0000111111;
								assign node395 = (inp[8]) ? 10'b0000001111 : 10'b0000011111;
							assign node398 = (inp[5]) ? node402 : node399;
								assign node399 = (inp[8]) ? 10'b0000001111 : 10'b0000011111;
								assign node402 = (inp[8]) ? 10'b0000000011 : 10'b0000001111;
					assign node405 = (inp[5]) ? node419 : node406;
						assign node406 = (inp[0]) ? node412 : node407;
							assign node407 = (inp[4]) ? node409 : 10'b0000111111;
								assign node409 = (inp[8]) ? 10'b0000001111 : 10'b0000011111;
							assign node412 = (inp[9]) ? node416 : node413;
								assign node413 = (inp[6]) ? 10'b0000001111 : 10'b0000011111;
								assign node416 = (inp[6]) ? 10'b0000000111 : 10'b0000001111;
						assign node419 = (inp[4]) ? node427 : node420;
							assign node420 = (inp[0]) ? node424 : node421;
								assign node421 = (inp[8]) ? 10'b0000001111 : 10'b0000011111;
								assign node424 = (inp[8]) ? 10'b0000000111 : 10'b0000001111;
							assign node427 = (inp[0]) ? node431 : node428;
								assign node428 = (inp[6]) ? 10'b0000000111 : 10'b0000001111;
								assign node431 = (inp[8]) ? 10'b0000000011 : 10'b0000000011;
				assign node434 = (inp[6]) ? node464 : node435;
					assign node435 = (inp[2]) ? node451 : node436;
						assign node436 = (inp[0]) ? node444 : node437;
							assign node437 = (inp[8]) ? node441 : node438;
								assign node438 = (inp[5]) ? 10'b0000001111 : 10'b0000111111;
								assign node441 = (inp[5]) ? 10'b0000001111 : 10'b0000011111;
							assign node444 = (inp[9]) ? node448 : node445;
								assign node445 = (inp[8]) ? 10'b0000001111 : 10'b0000001111;
								assign node448 = (inp[5]) ? 10'b0000000111 : 10'b0000001111;
						assign node451 = (inp[9]) ? node459 : node452;
							assign node452 = (inp[8]) ? node456 : node453;
								assign node453 = (inp[5]) ? 10'b0000001111 : 10'b0000001111;
								assign node456 = (inp[0]) ? 10'b0000000111 : 10'b0000001111;
							assign node459 = (inp[5]) ? node461 : 10'b0000000111;
								assign node461 = (inp[0]) ? 10'b0000000001 : 10'b0000000111;
					assign node464 = (inp[4]) ? node478 : node465;
						assign node465 = (inp[5]) ? node471 : node466;
							assign node466 = (inp[2]) ? node468 : 10'b0000001111;
								assign node468 = (inp[0]) ? 10'b0000000111 : 10'b0000001111;
							assign node471 = (inp[9]) ? node475 : node472;
								assign node472 = (inp[8]) ? 10'b0000000111 : 10'b0000001111;
								assign node475 = (inp[0]) ? 10'b0000000011 : 10'b0000000111;
						assign node478 = (inp[0]) ? node486 : node479;
							assign node479 = (inp[2]) ? node483 : node480;
								assign node480 = (inp[5]) ? 10'b0000000111 : 10'b0000001111;
								assign node483 = (inp[8]) ? 10'b0000000011 : 10'b0000000111;
							assign node486 = (inp[5]) ? node490 : node487;
								assign node487 = (inp[9]) ? 10'b0000000011 : 10'b0000000111;
								assign node490 = (inp[2]) ? 10'b0000000001 : 10'b0000000011;

endmodule