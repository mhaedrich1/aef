module dtc_split25_bm48 (
	input  wire [14-1:0] inp,
	output wire [14-1:0] outp
);

	wire [14-1:0] node1;
	wire [14-1:0] node2;
	wire [14-1:0] node3;
	wire [14-1:0] node4;
	wire [14-1:0] node6;
	wire [14-1:0] node7;
	wire [14-1:0] node8;
	wire [14-1:0] node9;
	wire [14-1:0] node13;
	wire [14-1:0] node15;
	wire [14-1:0] node16;
	wire [14-1:0] node20;
	wire [14-1:0] node22;
	wire [14-1:0] node23;
	wire [14-1:0] node25;
	wire [14-1:0] node27;
	wire [14-1:0] node31;
	wire [14-1:0] node32;
	wire [14-1:0] node33;
	wire [14-1:0] node35;
	wire [14-1:0] node36;
	wire [14-1:0] node38;
	wire [14-1:0] node39;
	wire [14-1:0] node43;
	wire [14-1:0] node44;
	wire [14-1:0] node45;
	wire [14-1:0] node50;
	wire [14-1:0] node52;
	wire [14-1:0] node53;
	wire [14-1:0] node54;
	wire [14-1:0] node56;
	wire [14-1:0] node60;
	wire [14-1:0] node61;
	wire [14-1:0] node63;
	wire [14-1:0] node66;
	wire [14-1:0] node67;
	wire [14-1:0] node71;
	wire [14-1:0] node72;
	wire [14-1:0] node74;
	wire [14-1:0] node75;
	wire [14-1:0] node76;
	wire [14-1:0] node82;
	wire [14-1:0] node83;
	wire [14-1:0] node85;
	wire [14-1:0] node87;
	wire [14-1:0] node89;
	wire [14-1:0] node90;
	wire [14-1:0] node94;
	wire [14-1:0] node95;
	wire [14-1:0] node96;
	wire [14-1:0] node97;
	wire [14-1:0] node98;
	wire [14-1:0] node101;
	wire [14-1:0] node102;
	wire [14-1:0] node104;
	wire [14-1:0] node108;
	wire [14-1:0] node110;
	wire [14-1:0] node111;
	wire [14-1:0] node112;
	wire [14-1:0] node117;
	wire [14-1:0] node118;
	wire [14-1:0] node119;
	wire [14-1:0] node121;
	wire [14-1:0] node122;
	wire [14-1:0] node128;
	wire [14-1:0] node129;
	wire [14-1:0] node131;
	wire [14-1:0] node133;
	wire [14-1:0] node134;
	wire [14-1:0] node138;
	wire [14-1:0] node139;
	wire [14-1:0] node140;
	wire [14-1:0] node142;
	wire [14-1:0] node143;
	wire [14-1:0] node146;
	wire [14-1:0] node149;
	wire [14-1:0] node150;
	wire [14-1:0] node151;
	wire [14-1:0] node154;
	wire [14-1:0] node158;
	wire [14-1:0] node160;
	wire [14-1:0] node161;
	wire [14-1:0] node163;
	wire [14-1:0] node167;
	wire [14-1:0] node168;
	wire [14-1:0] node169;
	wire [14-1:0] node170;
	wire [14-1:0] node171;
	wire [14-1:0] node173;
	wire [14-1:0] node174;
	wire [14-1:0] node176;
	wire [14-1:0] node182;
	wire [14-1:0] node183;
	wire [14-1:0] node184;
	wire [14-1:0] node185;
	wire [14-1:0] node186;
	wire [14-1:0] node188;
	wire [14-1:0] node189;
	wire [14-1:0] node195;
	wire [14-1:0] node196;
	wire [14-1:0] node197;
	wire [14-1:0] node200;
	wire [14-1:0] node203;
	wire [14-1:0] node204;
	wire [14-1:0] node205;
	wire [14-1:0] node209;
	wire [14-1:0] node210;
	wire [14-1:0] node214;
	wire [14-1:0] node215;
	wire [14-1:0] node217;
	wire [14-1:0] node219;
	wire [14-1:0] node221;
	wire [14-1:0] node225;
	wire [14-1:0] node226;
	wire [14-1:0] node227;
	wire [14-1:0] node228;
	wire [14-1:0] node229;
	wire [14-1:0] node230;
	wire [14-1:0] node231;
	wire [14-1:0] node235;
	wire [14-1:0] node236;
	wire [14-1:0] node237;
	wire [14-1:0] node241;
	wire [14-1:0] node243;
	wire [14-1:0] node248;
	wire [14-1:0] node249;
	wire [14-1:0] node251;
	wire [14-1:0] node253;
	wire [14-1:0] node256;
	wire [14-1:0] node257;
	wire [14-1:0] node258;
	wire [14-1:0] node260;
	wire [14-1:0] node261;
	wire [14-1:0] node264;
	wire [14-1:0] node268;
	wire [14-1:0] node270;
	wire [14-1:0] node272;
	wire [14-1:0] node274;
	wire [14-1:0] node277;
	wire [14-1:0] node278;
	wire [14-1:0] node279;
	wire [14-1:0] node280;
	wire [14-1:0] node281;
	wire [14-1:0] node284;
	wire [14-1:0] node288;
	wire [14-1:0] node290;
	wire [14-1:0] node291;
	wire [14-1:0] node294;
	wire [14-1:0] node296;
	wire [14-1:0] node298;
	wire [14-1:0] node302;
	wire [14-1:0] node303;
	wire [14-1:0] node304;
	wire [14-1:0] node305;
	wire [14-1:0] node307;
	wire [14-1:0] node309;
	wire [14-1:0] node310;
	wire [14-1:0] node311;
	wire [14-1:0] node312;
	wire [14-1:0] node314;
	wire [14-1:0] node319;
	wire [14-1:0] node321;
	wire [14-1:0] node323;
	wire [14-1:0] node325;
	wire [14-1:0] node328;
	wire [14-1:0] node330;
	wire [14-1:0] node331;
	wire [14-1:0] node332;
	wire [14-1:0] node333;
	wire [14-1:0] node334;
	wire [14-1:0] node335;
	wire [14-1:0] node339;
	wire [14-1:0] node340;
	wire [14-1:0] node343;
	wire [14-1:0] node346;
	wire [14-1:0] node347;
	wire [14-1:0] node348;
	wire [14-1:0] node353;
	wire [14-1:0] node355;
	wire [14-1:0] node357;
	wire [14-1:0] node358;
	wire [14-1:0] node362;
	wire [14-1:0] node364;
	wire [14-1:0] node365;
	wire [14-1:0] node367;
	wire [14-1:0] node369;
	wire [14-1:0] node373;
	wire [14-1:0] node374;
	wire [14-1:0] node376;
	wire [14-1:0] node378;
	wire [14-1:0] node379;
	wire [14-1:0] node381;
	wire [14-1:0] node382;
	wire [14-1:0] node383;
	wire [14-1:0] node389;
	wire [14-1:0] node390;
	wire [14-1:0] node391;
	wire [14-1:0] node392;
	wire [14-1:0] node393;
	wire [14-1:0] node394;
	wire [14-1:0] node397;
	wire [14-1:0] node400;
	wire [14-1:0] node401;
	wire [14-1:0] node403;
	wire [14-1:0] node408;
	wire [14-1:0] node409;
	wire [14-1:0] node410;
	wire [14-1:0] node411;
	wire [14-1:0] node412;
	wire [14-1:0] node417;
	wire [14-1:0] node418;
	wire [14-1:0] node420;
	wire [14-1:0] node423;
	wire [14-1:0] node424;
	wire [14-1:0] node428;
	wire [14-1:0] node429;
	wire [14-1:0] node430;
	wire [14-1:0] node432;
	wire [14-1:0] node435;
	wire [14-1:0] node436;
	wire [14-1:0] node441;
	wire [14-1:0] node443;
	wire [14-1:0] node445;
	wire [14-1:0] node446;
	wire [14-1:0] node448;
	wire [14-1:0] node450;
	wire [14-1:0] node453;
	wire [14-1:0] node454;
	wire [14-1:0] node455;
	wire [14-1:0] node460;
	wire [14-1:0] node461;
	wire [14-1:0] node462;
	wire [14-1:0] node463;
	wire [14-1:0] node464;
	wire [14-1:0] node466;
	wire [14-1:0] node467;
	wire [14-1:0] node468;
	wire [14-1:0] node473;
	wire [14-1:0] node474;
	wire [14-1:0] node476;
	wire [14-1:0] node478;
	wire [14-1:0] node479;
	wire [14-1:0] node483;
	wire [14-1:0] node484;
	wire [14-1:0] node485;
	wire [14-1:0] node486;
	wire [14-1:0] node491;
	wire [14-1:0] node492;
	wire [14-1:0] node494;
	wire [14-1:0] node498;
	wire [14-1:0] node499;
	wire [14-1:0] node501;
	wire [14-1:0] node502;
	wire [14-1:0] node503;
	wire [14-1:0] node504;
	wire [14-1:0] node508;
	wire [14-1:0] node509;
	wire [14-1:0] node514;
	wire [14-1:0] node516;
	wire [14-1:0] node517;
	wire [14-1:0] node520;
	wire [14-1:0] node521;
	wire [14-1:0] node523;
	wire [14-1:0] node527;
	wire [14-1:0] node528;
	wire [14-1:0] node529;
	wire [14-1:0] node530;
	wire [14-1:0] node532;
	wire [14-1:0] node536;
	wire [14-1:0] node537;
	wire [14-1:0] node538;
	wire [14-1:0] node539;
	wire [14-1:0] node541;
	wire [14-1:0] node544;
	wire [14-1:0] node546;
	wire [14-1:0] node549;
	wire [14-1:0] node550;
	wire [14-1:0] node551;
	wire [14-1:0] node555;
	wire [14-1:0] node558;
	wire [14-1:0] node560;
	wire [14-1:0] node562;
	wire [14-1:0] node564;
	wire [14-1:0] node568;
	wire [14-1:0] node569;
	wire [14-1:0] node570;
	wire [14-1:0] node572;
	wire [14-1:0] node573;
	wire [14-1:0] node574;
	wire [14-1:0] node575;
	wire [14-1:0] node576;
	wire [14-1:0] node582;
	wire [14-1:0] node584;
	wire [14-1:0] node587;
	wire [14-1:0] node588;
	wire [14-1:0] node589;
	wire [14-1:0] node590;
	wire [14-1:0] node592;
	wire [14-1:0] node593;
	wire [14-1:0] node597;
	wire [14-1:0] node601;
	wire [14-1:0] node603;
	wire [14-1:0] node604;
	wire [14-1:0] node605;
	wire [14-1:0] node606;
	wire [14-1:0] node609;
	wire [14-1:0] node612;
	wire [14-1:0] node613;
	wire [14-1:0] node617;
	wire [14-1:0] node619;
	wire [14-1:0] node621;
	wire [14-1:0] node624;
	wire [14-1:0] node625;
	wire [14-1:0] node626;
	wire [14-1:0] node627;
	wire [14-1:0] node629;
	wire [14-1:0] node630;
	wire [14-1:0] node634;
	wire [14-1:0] node635;
	wire [14-1:0] node639;
	wire [14-1:0] node641;
	wire [14-1:0] node643;
	wire [14-1:0] node645;
	wire [14-1:0] node646;

	assign outp = (inp[10]) ? node302 : node1;
		assign node1 = (inp[8]) ? node167 : node2;
			assign node2 = (inp[11]) ? node82 : node3;
				assign node3 = (inp[12]) ? node31 : node4;
					assign node4 = (inp[13]) ? node6 : 14'b00000100000011;
						assign node6 = (inp[9]) ? node20 : node7;
							assign node7 = (inp[6]) ? node13 : node8;
								assign node8 = (inp[3]) ? 14'b00000000000000 : node9;
									assign node9 = (inp[1]) ? 14'b11000000000100 : 14'b00000000000000;
								assign node13 = (inp[3]) ? node15 : 14'b00000000000000;
									assign node15 = (inp[7]) ? 14'b00000000000000 : node16;
										assign node16 = (inp[1]) ? 14'b00000000000000 : 14'b11000000000100;
							assign node20 = (inp[1]) ? node22 : 14'b00000000000000;
								assign node22 = (inp[5]) ? 14'b00000000000000 : node23;
									assign node23 = (inp[6]) ? node25 : 14'b00000000000000;
										assign node25 = (inp[3]) ? node27 : 14'b00000000000000;
											assign node27 = (inp[2]) ? 14'b01100000000110 : 14'b00000000000000;
					assign node31 = (inp[0]) ? node71 : node32;
						assign node32 = (inp[1]) ? node50 : node33;
							assign node33 = (inp[3]) ? node35 : 14'b00000000000000;
								assign node35 = (inp[5]) ? node43 : node36;
									assign node36 = (inp[13]) ? node38 : 14'b00000000000000;
										assign node38 = (inp[7]) ? 14'b00000000000000 : node39;
											assign node39 = (inp[9]) ? 14'b00000000000000 : 14'b00000000000000;
									assign node43 = (inp[13]) ? 14'b00000000000000 : node44;
										assign node44 = (inp[2]) ? 14'b00000000000000 : node45;
											assign node45 = (inp[9]) ? 14'b00000000000000 : 14'b00000000000000;
							assign node50 = (inp[5]) ? node52 : 14'b00000000000000;
								assign node52 = (inp[13]) ? node60 : node53;
									assign node53 = (inp[2]) ? 14'b00000000000000 : node54;
										assign node54 = (inp[6]) ? node56 : 14'b00000000000000;
											assign node56 = (inp[7]) ? 14'b00001000000101 : 14'b00000000000000;
									assign node60 = (inp[7]) ? node66 : node61;
										assign node61 = (inp[3]) ? node63 : 14'b00000000000000;
											assign node63 = (inp[6]) ? 14'b00000000011101 : 14'b00000000000000;
										assign node66 = (inp[2]) ? 14'b00000000000000 : node67;
											assign node67 = (inp[6]) ? 14'b00000000000000 : 14'b11110111110010;
						assign node71 = (inp[4]) ? 14'b00000000000000 : node72;
							assign node72 = (inp[1]) ? node74 : 14'b00000000000000;
								assign node74 = (inp[3]) ? 14'b00000000000000 : node75;
									assign node75 = (inp[5]) ? 14'b00000000000000 : node76;
										assign node76 = (inp[2]) ? 14'b00000000000000 : 14'b00100000000011;
				assign node82 = (inp[1]) ? node94 : node83;
					assign node83 = (inp[12]) ? node85 : 14'b00000000000000;
						assign node85 = (inp[6]) ? node87 : 14'b00000000000000;
							assign node87 = (inp[3]) ? node89 : 14'b00000000000000;
								assign node89 = (inp[9]) ? 14'b00000000000000 : node90;
									assign node90 = (inp[13]) ? 14'b00100100001101 : 14'b01100000001010;
					assign node94 = (inp[6]) ? node128 : node95;
						assign node95 = (inp[9]) ? node117 : node96;
							assign node96 = (inp[3]) ? node108 : node97;
								assign node97 = (inp[13]) ? node101 : node98;
									assign node98 = (inp[12]) ? 14'b10000100011000 : 14'b00000000000000;
									assign node101 = (inp[12]) ? 14'b00000000000000 : node102;
										assign node102 = (inp[2]) ? node104 : 14'b00000000000000;
											assign node104 = (inp[7]) ? 14'b10110101111111 : 14'b00000000000000;
								assign node108 = (inp[13]) ? node110 : 14'b00000000000000;
									assign node110 = (inp[2]) ? 14'b00000000000000 : node111;
										assign node111 = (inp[0]) ? 14'b00000000000000 : node112;
											assign node112 = (inp[12]) ? 14'b10010101111110 : 14'b10000100101010;
							assign node117 = (inp[2]) ? 14'b00000000000000 : node118;
								assign node118 = (inp[0]) ? 14'b00000000000000 : node119;
									assign node119 = (inp[7]) ? node121 : 14'b00000000000000;
										assign node121 = (inp[12]) ? 14'b10100010001100 : node122;
											assign node122 = (inp[13]) ? 14'b00000000000000 : 14'b10010000001101;
						assign node128 = (inp[7]) ? node138 : node129;
							assign node129 = (inp[5]) ? node131 : 14'b00000000000000;
								assign node131 = (inp[3]) ? node133 : 14'b00000000000000;
									assign node133 = (inp[0]) ? 14'b00000000000000 : node134;
										assign node134 = (inp[12]) ? 14'b00000000011100 : 14'b00000000000000;
							assign node138 = (inp[2]) ? node158 : node139;
								assign node139 = (inp[9]) ? node149 : node140;
									assign node140 = (inp[12]) ? node142 : 14'b00000000000000;
										assign node142 = (inp[13]) ? node146 : node143;
											assign node143 = (inp[4]) ? 14'b00000000000000 : 14'b00000000000000;
											assign node146 = (inp[5]) ? 14'b00001000000001 : 14'b00000000000000;
									assign node149 = (inp[12]) ? 14'b00000000000000 : node150;
										assign node150 = (inp[5]) ? node154 : node151;
											assign node151 = (inp[0]) ? 14'b00000000000000 : 14'b10100000111010;
											assign node154 = (inp[0]) ? 14'b01001000000101 : 14'b00000000000000;
								assign node158 = (inp[5]) ? node160 : 14'b00000000000000;
									assign node160 = (inp[12]) ? 14'b00000000000000 : node161;
										assign node161 = (inp[3]) ? node163 : 14'b00000000000000;
											assign node163 = (inp[13]) ? 14'b01001000000101 : 14'b00000000000000;
			assign node167 = (inp[12]) ? node225 : node168;
				assign node168 = (inp[1]) ? node182 : node169;
					assign node169 = (inp[0]) ? 14'b00000000000000 : node170;
						assign node170 = (inp[7]) ? 14'b00000000000000 : node171;
							assign node171 = (inp[11]) ? node173 : 14'b00000000000000;
								assign node173 = (inp[9]) ? 14'b00000000000000 : node174;
									assign node174 = (inp[3]) ? node176 : 14'b00000000000000;
										assign node176 = (inp[13]) ? 14'b00100000000011 : 14'b00000000000000;
					assign node182 = (inp[6]) ? node214 : node183;
						assign node183 = (inp[11]) ? node195 : node184;
							assign node184 = (inp[13]) ? 14'b00000000000000 : node185;
								assign node185 = (inp[0]) ? 14'b00000000000000 : node186;
									assign node186 = (inp[3]) ? node188 : 14'b00000000000000;
										assign node188 = (inp[2]) ? 14'b00000000000000 : node189;
											assign node189 = (inp[4]) ? 14'b10100100101000 : 14'b10100100111000;
							assign node195 = (inp[3]) ? node203 : node196;
								assign node196 = (inp[13]) ? node200 : node197;
									assign node197 = (inp[9]) ? 14'b00000000000000 : 14'b01001000000100;
									assign node200 = (inp[9]) ? 14'b00000000000000 : 14'b00000000011100;
								assign node203 = (inp[13]) ? node209 : node204;
									assign node204 = (inp[7]) ? 14'b00000000000000 : node205;
										assign node205 = (inp[2]) ? 14'b00000000000000 : 14'b00000100000001;
									assign node209 = (inp[4]) ? 14'b00000000000000 : node210;
										assign node210 = (inp[5]) ? 14'b00000000000000 : 14'b00000000011100;
						assign node214 = (inp[13]) ? 14'b00000000000000 : node215;
							assign node215 = (inp[7]) ? node217 : 14'b00000000000000;
								assign node217 = (inp[3]) ? node219 : 14'b00000000000000;
									assign node219 = (inp[9]) ? node221 : 14'b00000000000000;
										assign node221 = (inp[4]) ? 14'b00000000000000 : 14'b00000000011100;
				assign node225 = (inp[11]) ? node277 : node226;
					assign node226 = (inp[6]) ? node248 : node227;
						assign node227 = (inp[0]) ? 14'b00000000000000 : node228;
							assign node228 = (inp[2]) ? 14'b00000000000000 : node229;
								assign node229 = (inp[5]) ? node235 : node230;
									assign node230 = (inp[7]) ? 14'b00000000000000 : node231;
										assign node231 = (inp[4]) ? 14'b00001000000101 : 14'b00000000000000;
									assign node235 = (inp[4]) ? node241 : node236;
										assign node236 = (inp[3]) ? 14'b10000100111010 : node237;
											assign node237 = (inp[9]) ? 14'b00000000000000 : 14'b00000000011100;
										assign node241 = (inp[1]) ? node243 : 14'b00000000000000;
											assign node243 = (inp[7]) ? 14'b00000000000000 : 14'b10000100101010;
						assign node248 = (inp[13]) ? node256 : node249;
							assign node249 = (inp[9]) ? node251 : 14'b00000000000000;
								assign node251 = (inp[3]) ? node253 : 14'b00000000000000;
									assign node253 = (inp[1]) ? 14'b00000000000000 : 14'b11110111110010;
							assign node256 = (inp[9]) ? node268 : node257;
								assign node257 = (inp[3]) ? 14'b00000000000000 : node258;
									assign node258 = (inp[1]) ? node260 : 14'b00000000000000;
										assign node260 = (inp[5]) ? node264 : node261;
											assign node261 = (inp[7]) ? 14'b00000000000000 : 14'b10010100011100;
											assign node264 = (inp[0]) ? 14'b11100100010100 : 14'b11100100000100;
								assign node268 = (inp[3]) ? node270 : 14'b00000000000000;
									assign node270 = (inp[1]) ? node272 : 14'b01001000000100;
										assign node272 = (inp[7]) ? node274 : 14'b00000000000000;
											assign node274 = (inp[5]) ? 14'b01001000001001 : 14'b00000000000000;
					assign node277 = (inp[13]) ? 14'b01000000010100 : node278;
						assign node278 = (inp[3]) ? node288 : node279;
							assign node279 = (inp[9]) ? 14'b00000000000000 : node280;
								assign node280 = (inp[6]) ? node284 : node281;
									assign node281 = (inp[1]) ? 14'b00100100011111 : 14'b00000000000000;
									assign node284 = (inp[1]) ? 14'b01000100000100 : 14'b00000000000000;
							assign node288 = (inp[9]) ? node290 : 14'b00000000000000;
								assign node290 = (inp[1]) ? node294 : node291;
									assign node291 = (inp[6]) ? 14'b10100010001100 : 14'b00000000000000;
									assign node294 = (inp[5]) ? node296 : 14'b00000000000000;
										assign node296 = (inp[7]) ? node298 : 14'b00000000000000;
											assign node298 = (inp[4]) ? 14'b00000000000000 : 14'b10000000011010;
		assign node302 = (inp[12]) ? node460 : node303;
			assign node303 = (inp[13]) ? node373 : node304;
				assign node304 = (inp[11]) ? node328 : node305;
					assign node305 = (inp[8]) ? node307 : 14'b10000100001000;
						assign node307 = (inp[1]) ? node309 : 14'b00000000000000;
							assign node309 = (inp[6]) ? node319 : node310;
								assign node310 = (inp[9]) ? 14'b00000000000000 : node311;
									assign node311 = (inp[3]) ? 14'b00000000000000 : node312;
										assign node312 = (inp[5]) ? node314 : 14'b00100000000011;
											assign node314 = (inp[7]) ? 14'b00100000000011 : 14'b00000000000000;
								assign node319 = (inp[7]) ? node321 : 14'b00000000000000;
									assign node321 = (inp[3]) ? node323 : 14'b00000000000000;
										assign node323 = (inp[9]) ? node325 : 14'b00000000000000;
											assign node325 = (inp[5]) ? 14'b10100000001000 : 14'b00000000000000;
					assign node328 = (inp[1]) ? node330 : 14'b00000000000000;
						assign node330 = (inp[6]) ? node362 : node331;
							assign node331 = (inp[9]) ? node353 : node332;
								assign node332 = (inp[3]) ? node346 : node333;
									assign node333 = (inp[8]) ? node339 : node334;
										assign node334 = (inp[5]) ? 14'b00000000000000 : node335;
											assign node335 = (inp[2]) ? 14'b01001000000101 : 14'b00000000000000;
										assign node339 = (inp[4]) ? node343 : node340;
											assign node340 = (inp[5]) ? 14'b00000000000000 : 14'b10000001001101;
											assign node343 = (inp[2]) ? 14'b10000100001101 : 14'b10000010001101;
									assign node346 = (inp[2]) ? 14'b00000000000000 : node347;
										assign node347 = (inp[0]) ? 14'b00000000000000 : node348;
											assign node348 = (inp[7]) ? 14'b00100000000011 : 14'b00100000001010;
								assign node353 = (inp[4]) ? node355 : 14'b00000000000000;
									assign node355 = (inp[3]) ? node357 : 14'b00000000000000;
										assign node357 = (inp[7]) ? 14'b00000000000000 : node358;
											assign node358 = (inp[0]) ? 14'b00000000000000 : 14'b00100000001010;
							assign node362 = (inp[9]) ? node364 : 14'b00000000000000;
								assign node364 = (inp[5]) ? 14'b00000000000000 : node365;
									assign node365 = (inp[7]) ? node367 : 14'b00000000000000;
										assign node367 = (inp[3]) ? node369 : 14'b00000000000000;
											assign node369 = (inp[8]) ? 14'b01001000000100 : 14'b00000100001111;
				assign node373 = (inp[1]) ? node389 : node374;
					assign node374 = (inp[8]) ? node376 : 14'b00000000000000;
						assign node376 = (inp[3]) ? node378 : 14'b00000000000000;
							assign node378 = (inp[2]) ? 14'b00000000000000 : node379;
								assign node379 = (inp[11]) ? node381 : 14'b00000000000000;
									assign node381 = (inp[7]) ? 14'b00000000000000 : node382;
										assign node382 = (inp[0]) ? 14'b00000000000000 : node383;
											assign node383 = (inp[6]) ? 14'b10000100111010 : 14'b00000000000000;
					assign node389 = (inp[2]) ? node441 : node390;
						assign node390 = (inp[11]) ? node408 : node391;
							assign node391 = (inp[6]) ? 14'b00000000000000 : node392;
								assign node392 = (inp[0]) ? node400 : node393;
									assign node393 = (inp[7]) ? node397 : node394;
										assign node394 = (inp[8]) ? 14'b00001000001001 : 14'b00000000000000;
										assign node397 = (inp[8]) ? 14'b00000000000000 : 14'b00001000000100;
									assign node400 = (inp[3]) ? 14'b00000000000000 : node401;
										assign node401 = (inp[7]) ? node403 : 14'b00000000000000;
											assign node403 = (inp[5]) ? 14'b00000000000000 : 14'b00000000000000;
							assign node408 = (inp[8]) ? node428 : node409;
								assign node409 = (inp[3]) ? node417 : node410;
									assign node410 = (inp[5]) ? 14'b00000000000000 : node411;
										assign node411 = (inp[4]) ? 14'b00000000000000 : node412;
											assign node412 = (inp[0]) ? 14'b00000000000000 : 14'b00000000000000;
									assign node417 = (inp[6]) ? node423 : node418;
										assign node418 = (inp[4]) ? node420 : 14'b00000000000000;
											assign node420 = (inp[9]) ? 14'b00000000000000 : 14'b00100000000011;
										assign node423 = (inp[5]) ? 14'b10100101111111 : node424;
											assign node424 = (inp[7]) ? 14'b00001000001001 : 14'b00000000000000;
								assign node428 = (inp[6]) ? 14'b00000000000000 : node429;
									assign node429 = (inp[9]) ? node435 : node430;
										assign node430 = (inp[0]) ? node432 : 14'b10000000001010;
											assign node432 = (inp[3]) ? 14'b00000000000000 : 14'b10100100011000;
										assign node435 = (inp[5]) ? 14'b00000000000000 : node436;
											assign node436 = (inp[0]) ? 14'b00000000000000 : 14'b10100100111000;
						assign node441 = (inp[11]) ? node443 : 14'b00000000000000;
							assign node443 = (inp[7]) ? node445 : 14'b00000000000000;
								assign node445 = (inp[8]) ? node453 : node446;
									assign node446 = (inp[3]) ? node448 : 14'b00000000000000;
										assign node448 = (inp[6]) ? node450 : 14'b00000000000000;
											assign node450 = (inp[9]) ? 14'b01000100000010 : 14'b00000000000000;
									assign node453 = (inp[3]) ? 14'b00000000000000 : node454;
										assign node454 = (inp[6]) ? 14'b00000000000000 : node455;
											assign node455 = (inp[9]) ? 14'b00000000000000 : 14'b10100100011000;
			assign node460 = (inp[13]) ? node568 : node461;
				assign node461 = (inp[11]) ? node527 : node462;
					assign node462 = (inp[8]) ? node498 : node463;
						assign node463 = (inp[6]) ? node473 : node464;
							assign node464 = (inp[0]) ? node466 : 14'b00000000000000;
								assign node466 = (inp[7]) ? 14'b00000000000000 : node467;
									assign node467 = (inp[9]) ? 14'b00000000000000 : node468;
										assign node468 = (inp[4]) ? 14'b00000000000000 : 14'b01001000000100;
							assign node473 = (inp[3]) ? node483 : node474;
								assign node474 = (inp[5]) ? node476 : 14'b00000000000000;
									assign node476 = (inp[7]) ? node478 : 14'b00000000000000;
										assign node478 = (inp[9]) ? 14'b00000000000000 : node479;
											assign node479 = (inp[4]) ? 14'b00000000000000 : 14'b00000000000000;
								assign node483 = (inp[9]) ? node491 : node484;
									assign node484 = (inp[2]) ? 14'b00000000000000 : node485;
										assign node485 = (inp[1]) ? 14'b00000000000000 : node486;
											assign node486 = (inp[7]) ? 14'b00000000000000 : 14'b10100100101000;
									assign node491 = (inp[7]) ? 14'b00000000000000 : node492;
										assign node492 = (inp[5]) ? node494 : 14'b00000000000000;
											assign node494 = (inp[1]) ? 14'b00001000001100 : 14'b00000000000000;
						assign node498 = (inp[9]) ? node514 : node499;
							assign node499 = (inp[1]) ? node501 : 14'b00000000000000;
								assign node501 = (inp[6]) ? 14'b00000000000000 : node502;
									assign node502 = (inp[3]) ? node508 : node503;
										assign node503 = (inp[0]) ? 14'b00000000000000 : node504;
											assign node504 = (inp[2]) ? 14'b00000000000000 : 14'b10100100101000;
										assign node508 = (inp[0]) ? 14'b00000000000000 : node509;
											assign node509 = (inp[7]) ? 14'b00000000000000 : 14'b00000000011100;
							assign node514 = (inp[3]) ? node516 : 14'b00000000000000;
								assign node516 = (inp[1]) ? node520 : node517;
									assign node517 = (inp[6]) ? 14'b01100000001010 : 14'b00000000000000;
									assign node520 = (inp[0]) ? 14'b00000000000000 : node521;
										assign node521 = (inp[6]) ? node523 : 14'b00000000011100;
											assign node523 = (inp[7]) ? 14'b00000000000000 : 14'b00000000000000;
					assign node527 = (inp[8]) ? 14'b00000000000000 : node528;
						assign node528 = (inp[1]) ? node536 : node529;
							assign node529 = (inp[9]) ? 14'b00000000000000 : node530;
								assign node530 = (inp[6]) ? node532 : 14'b00000000000000;
									assign node532 = (inp[3]) ? 14'b01001000000101 : 14'b00000000000000;
							assign node536 = (inp[2]) ? node558 : node537;
								assign node537 = (inp[0]) ? node549 : node538;
									assign node538 = (inp[9]) ? node544 : node539;
										assign node539 = (inp[3]) ? node541 : 14'b00000000000000;
											assign node541 = (inp[4]) ? 14'b00100100001101 : 14'b00000000000000;
										assign node544 = (inp[3]) ? node546 : 14'b00100100001101;
											assign node546 = (inp[7]) ? 14'b00000000000000 : 14'b00000100001111;
									assign node549 = (inp[4]) ? node555 : node550;
										assign node550 = (inp[3]) ? 14'b00000000000000 : node551;
											assign node551 = (inp[9]) ? 14'b00000000000000 : 14'b00001000000101;
										assign node555 = (inp[6]) ? 14'b00000100001111 : 14'b00000000000000;
								assign node558 = (inp[4]) ? node560 : 14'b00000000000000;
									assign node560 = (inp[3]) ? node562 : 14'b00000000000000;
										assign node562 = (inp[9]) ? node564 : 14'b00000000000000;
											assign node564 = (inp[6]) ? 14'b00000100001111 : 14'b00000000000000;
				assign node568 = (inp[11]) ? node624 : node569;
					assign node569 = (inp[1]) ? node587 : node570;
						assign node570 = (inp[3]) ? node572 : 14'b00000000000000;
							assign node572 = (inp[9]) ? node582 : node573;
								assign node573 = (inp[7]) ? 14'b00000000000000 : node574;
									assign node574 = (inp[2]) ? 14'b00000000000000 : node575;
										assign node575 = (inp[5]) ? 14'b00000000000000 : node576;
											assign node576 = (inp[4]) ? 14'b00000000000000 : 14'b10000000111000;
								assign node582 = (inp[8]) ? node584 : 14'b00000000000000;
									assign node584 = (inp[6]) ? 14'b00100100001101 : 14'b00000000000000;
						assign node587 = (inp[3]) ? node601 : node588;
							assign node588 = (inp[9]) ? 14'b00000000000000 : node589;
								assign node589 = (inp[6]) ? node597 : node590;
									assign node590 = (inp[8]) ? node592 : 14'b00000000011101;
										assign node592 = (inp[2]) ? 14'b00001000000100 : node593;
											assign node593 = (inp[0]) ? 14'b00001000000100 : 14'b10000000101000;
									assign node597 = (inp[8]) ? 14'b00000100001110 : 14'b00000000000000;
							assign node601 = (inp[9]) ? node603 : 14'b00000000000000;
								assign node603 = (inp[2]) ? node617 : node604;
									assign node604 = (inp[0]) ? node612 : node605;
										assign node605 = (inp[5]) ? node609 : node606;
											assign node606 = (inp[6]) ? 14'b00000000000000 : 14'b01100000001010;
											assign node609 = (inp[7]) ? 14'b00000000011100 : 14'b00000000011101;
										assign node612 = (inp[8]) ? 14'b00000000000000 : node613;
											assign node613 = (inp[5]) ? 14'b00000000000000 : 14'b00000000000000;
									assign node617 = (inp[5]) ? node619 : 14'b00000000000000;
										assign node619 = (inp[6]) ? node621 : 14'b00000000000000;
											assign node621 = (inp[4]) ? 14'b00000000000000 : 14'b00000000000000;
					assign node624 = (inp[8]) ? 14'b10000100001000 : node625;
						assign node625 = (inp[9]) ? node639 : node626;
							assign node626 = (inp[3]) ? node634 : node627;
								assign node627 = (inp[1]) ? node629 : 14'b00000000000000;
									assign node629 = (inp[0]) ? 14'b00000000000000 : node630;
										assign node630 = (inp[7]) ? 14'b01001000000101 : 14'b00000000000000;
								assign node634 = (inp[1]) ? 14'b00000000000000 : node635;
									assign node635 = (inp[6]) ? 14'b10010101111110 : 14'b00000000000000;
							assign node639 = (inp[2]) ? node641 : 14'b00000000000000;
								assign node641 = (inp[1]) ? node643 : 14'b00000000000000;
									assign node643 = (inp[6]) ? node645 : 14'b00000000000000;
										assign node645 = (inp[4]) ? 14'b00000000000000 : node646;
											assign node646 = (inp[5]) ? 14'b10100100001000 : 14'b00000000000000;

endmodule